magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< poly >>
rect -50 50 0 66
rect -50 16 -34 50
rect -50 0 0 16
rect 31246 -274 31297 -258
rect 31280 -308 31297 -274
rect 31246 -324 31297 -308
<< polycont >>
rect -34 16 0 50
rect 31246 -308 31280 -274
<< npolyres >>
rect 0 0 31297 66
rect 31231 -96 31297 0
rect -50 -162 31297 -96
rect -50 -258 16 -162
rect -50 -324 31246 -258
<< locali >>
rect -34 50 0 66
rect -34 0 0 16
rect 31246 -274 31281 -258
rect 31280 -308 31281 -274
rect 31246 -324 31281 -308
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_0
timestamp 1701704242
transform 1 0 31230 0 1 -324
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_1
timestamp 1701704242
transform 1 0 -50 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 34450354
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 34449298
<< end >>
