magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -89 -36 245 1036
<< pmos >>
rect 0 0 50 1000
rect 106 0 156 1000
<< pdiff >>
rect -50 0 0 1000
rect 156 0 206 1000
<< poly >>
rect 0 1000 50 1026
rect 0 -26 50 0
rect 106 1000 156 1026
rect 106 -26 156 0
<< locali >>
rect -45 -4 -11 946
rect 61 -4 95 946
rect 167 -4 201 946
use DFL1sd2_CDNS_52468879185113  DFL1sd2_CDNS_52468879185113_0
timestamp 1701704242
transform 1 0 50 0 1 0
box -36 -36 92 1036
use DFL1sd_CDNS_52468879185122  DFL1sd_CDNS_52468879185122_0
timestamp 1701704242
transform -1 0 0 0 1 0
box -36 -36 89 1036
use DFL1sd_CDNS_52468879185122  DFL1sd_CDNS_52468879185122_1
timestamp 1701704242
transform 1 0 156 0 1 0
box -36 -36 89 1036
<< labels >>
flabel comment s -28 471 -28 471 0 FreeSans 300 0 0 0 S
flabel comment s 78 471 78 471 0 FreeSans 300 0 0 0 D
flabel comment s 184 471 184 471 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 80363740
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 80362164
<< end >>
