magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -74 825 1614 2035
<< pwell >>
rect 788 61 874 735
rect 1488 61 1574 735
rect 788 -25 1574 61
<< mvpsubdiff >>
rect 814 685 848 709
rect 814 615 848 651
rect 1514 685 1548 709
rect 814 545 848 581
rect 814 475 848 511
rect 814 405 848 441
rect 814 336 848 371
rect 814 267 848 302
rect 814 198 848 233
rect 814 129 848 164
rect 814 35 848 95
rect 1514 616 1548 651
rect 1514 547 1548 582
rect 1514 478 1548 513
rect 1514 409 1548 444
rect 1514 339 1548 375
rect 1514 269 1548 305
rect 1514 199 1548 235
rect 1514 129 1548 165
rect 1514 59 1548 95
rect 814 1 838 35
rect 872 1 910 35
rect 944 1 982 35
rect 1016 1 1054 35
rect 1088 1 1126 35
rect 1160 1 1198 35
rect 1232 1 1270 35
rect 1304 1 1342 35
rect 1376 1 1414 35
rect 1448 25 1514 35
rect 1448 1 1548 25
<< mvnsubdiff >>
rect 0 1935 34 1969
rect 68 1935 103 1969
rect 137 1935 172 1969
rect 206 1935 241 1969
rect 275 1935 310 1969
rect 344 1935 379 1969
rect 413 1935 448 1969
rect 482 1935 517 1969
rect 551 1935 586 1969
rect 620 1935 655 1969
rect 689 1935 724 1969
rect 758 1935 793 1969
rect 827 1935 862 1969
rect 896 1935 931 1969
rect 965 1935 1000 1969
rect 1034 1935 1069 1969
rect 1103 1935 1138 1969
rect 1172 1935 1207 1969
rect 1241 1935 1275 1969
rect 1309 1935 1343 1969
rect 1377 1935 1411 1969
rect 1445 1935 1479 1969
rect 1513 1935 1547 1969
<< mvpsubdiffcont >>
rect 814 651 848 685
rect 1514 651 1548 685
rect 814 581 848 615
rect 814 511 848 545
rect 814 441 848 475
rect 814 371 848 405
rect 814 302 848 336
rect 814 233 848 267
rect 814 164 848 198
rect 814 95 848 129
rect 1514 582 1548 616
rect 1514 513 1548 547
rect 1514 444 1548 478
rect 1514 375 1548 409
rect 1514 305 1548 339
rect 1514 235 1548 269
rect 1514 165 1548 199
rect 1514 95 1548 129
rect 838 1 872 35
rect 910 1 944 35
rect 982 1 1016 35
rect 1054 1 1088 35
rect 1126 1 1160 35
rect 1198 1 1232 35
rect 1270 1 1304 35
rect 1342 1 1376 35
rect 1414 1 1448 35
rect 1514 25 1548 59
<< mvnsubdiffcont >>
rect 34 1935 68 1969
rect 103 1935 137 1969
rect 172 1935 206 1969
rect 241 1935 275 1969
rect 310 1935 344 1969
rect 379 1935 413 1969
rect 448 1935 482 1969
rect 517 1935 551 1969
rect 586 1935 620 1969
rect 655 1935 689 1969
rect 724 1935 758 1969
rect 793 1935 827 1969
rect 862 1935 896 1969
rect 931 1935 965 1969
rect 1000 1935 1034 1969
rect 1069 1935 1103 1969
rect 1138 1935 1172 1969
rect 1207 1935 1241 1969
rect 1275 1935 1309 1969
rect 1343 1935 1377 1969
rect 1411 1935 1445 1969
rect 1479 1935 1513 1969
<< poly >>
rect 45 829 145 835
rect 201 829 301 835
rect 357 829 457 835
rect 513 763 613 835
rect 669 797 769 835
rect 935 829 1035 835
rect 1091 829 1191 899
rect 1247 829 1347 899
rect 1403 829 1503 899
rect 669 763 685 797
rect 719 763 769 797
rect 914 813 1503 829
rect 914 779 930 813
rect 964 779 998 813
rect 1032 779 1066 813
rect 1100 779 1134 813
rect 1168 779 1503 813
rect 914 763 1503 779
rect 669 729 769 763
rect 669 695 685 729
rect 719 695 769 729
rect 669 679 769 695
rect 975 655 1075 763
rect 1131 655 1231 763
rect 1287 644 1387 763
<< polycont >>
rect 685 763 719 797
rect 930 779 964 813
rect 998 779 1032 813
rect 1066 779 1100 813
rect 1134 779 1168 813
rect 685 695 719 729
<< locali >>
rect 0 1865 34 1969
rect 68 1935 103 1969
rect 137 1935 172 1969
rect 206 1935 241 1969
rect 275 1935 310 1969
rect 344 1935 379 1969
rect 413 1935 448 1969
rect 482 1935 517 1969
rect 551 1935 586 1969
rect 620 1935 655 1969
rect 689 1935 724 1969
rect 758 1935 793 1969
rect 827 1935 862 1969
rect 896 1935 931 1969
rect 965 1935 1000 1969
rect 1034 1935 1069 1969
rect 1103 1935 1138 1969
rect 1172 1935 1207 1969
rect 1241 1935 1275 1969
rect 1309 1935 1343 1969
rect 1377 1935 1411 1969
rect 1445 1935 1479 1969
rect 1513 1935 1547 1969
rect 312 1865 346 1935
rect 624 1865 658 1935
rect 0 1474 34 1512
rect 0 1402 34 1440
rect 312 1474 346 1512
rect 312 1402 346 1440
rect 624 1474 658 1512
rect 624 1402 658 1440
rect 190 1068 228 1102
rect 430 1068 468 1102
rect 924 1068 962 1102
rect 1164 1068 1202 1102
rect 1476 1068 1514 1102
rect 1080 994 1118 1028
rect 1319 994 1357 1028
rect 780 813 814 915
rect 1358 869 1392 915
rect 1242 835 1392 869
rect 333 779 367 813
rect 685 797 719 813
rect 780 779 930 813
rect 964 779 998 813
rect 1032 779 1066 813
rect 1100 779 1134 813
rect 1168 779 1184 813
rect 685 729 719 763
rect 1242 713 1276 835
rect 685 679 719 695
rect 814 685 848 701
rect 814 615 848 651
rect 1514 685 1548 701
rect 1514 616 1548 651
rect 814 545 848 581
rect 964 566 1002 600
rect 1204 566 1242 600
rect 1514 547 1548 582
rect 814 475 848 511
rect 814 405 848 441
rect 814 336 848 371
rect 1086 448 1120 486
rect 1086 376 1120 414
rect 1398 448 1432 486
rect 1398 376 1432 414
rect 1514 478 1548 513
rect 1514 409 1548 444
rect 814 296 848 302
rect 814 224 848 233
rect 814 152 848 164
rect 814 35 848 95
rect 1514 339 1548 375
rect 1514 296 1548 305
rect 1514 224 1548 235
rect 1514 152 1548 165
rect 1514 59 1548 95
rect 814 1 838 35
rect 874 1 910 35
rect 953 1 982 35
rect 1033 1 1054 35
rect 1113 1 1126 35
rect 1193 1 1198 35
rect 1232 1 1239 35
rect 1304 1 1319 35
rect 1376 1 1399 35
rect 1448 1 1479 35
rect 1513 25 1514 35
rect 1513 1 1548 25
<< viali >>
rect 0 1512 34 1546
rect 0 1440 34 1474
rect 0 1368 34 1402
rect 312 1512 346 1546
rect 312 1440 346 1474
rect 312 1368 346 1402
rect 624 1512 658 1546
rect 624 1440 658 1474
rect 624 1368 658 1402
rect 156 1068 190 1102
rect 228 1068 262 1102
rect 396 1068 430 1102
rect 468 1068 502 1102
rect 890 1068 924 1102
rect 962 1068 996 1102
rect 1130 1068 1164 1102
rect 1202 1068 1236 1102
rect 1442 1068 1476 1102
rect 1514 1068 1548 1102
rect 1046 994 1080 1028
rect 1118 994 1152 1028
rect 1285 994 1319 1028
rect 1357 994 1391 1028
rect 930 566 964 600
rect 1002 566 1036 600
rect 1170 566 1204 600
rect 1242 566 1276 600
rect 1086 486 1120 520
rect 1086 414 1120 448
rect 1086 342 1120 376
rect 1398 486 1432 520
rect 1398 414 1432 448
rect 1398 342 1432 376
rect 814 267 848 296
rect 814 262 848 267
rect 814 198 848 224
rect 814 190 848 198
rect 814 129 848 152
rect 814 118 848 129
rect 1514 269 1548 296
rect 1514 262 1548 269
rect 1514 199 1548 224
rect 1514 190 1548 199
rect 1514 129 1548 152
rect 1514 118 1548 129
rect 840 1 872 35
rect 872 1 874 35
rect 919 1 944 35
rect 944 1 953 35
rect 999 1 1016 35
rect 1016 1 1033 35
rect 1079 1 1088 35
rect 1088 1 1113 35
rect 1159 1 1160 35
rect 1160 1 1193 35
rect 1239 1 1270 35
rect 1270 1 1273 35
rect 1319 1 1342 35
rect 1342 1 1353 35
rect 1399 1 1414 35
rect 1414 1 1433 35
rect 1479 1 1513 35
<< metal1 >>
rect -6 1546 667 1558
rect -6 1512 0 1546
rect 34 1512 312 1546
rect 346 1512 624 1546
rect 658 1512 667 1546
rect -6 1474 667 1512
rect -6 1440 0 1474
rect 34 1440 312 1474
rect 346 1440 624 1474
rect 658 1440 667 1474
rect -6 1402 667 1440
rect -6 1368 0 1402
rect 34 1368 312 1402
rect 346 1368 624 1402
rect 658 1368 667 1402
rect -6 1356 667 1368
rect 144 1102 1560 1108
rect 144 1068 156 1102
rect 190 1068 228 1102
rect 262 1068 396 1102
rect 430 1068 468 1102
rect 502 1068 890 1102
rect 924 1068 962 1102
rect 996 1068 1130 1102
rect 1164 1068 1202 1102
rect 1236 1068 1442 1102
rect 1476 1068 1514 1102
rect 1548 1068 1560 1102
rect 144 1062 1560 1068
rect 1034 1028 1403 1034
rect 1034 994 1046 1028
rect 1080 994 1118 1028
rect 1152 994 1285 1028
rect 1319 994 1357 1028
rect 1391 994 1403 1028
rect 1034 988 1403 994
rect 918 600 1288 606
rect 918 566 930 600
rect 964 566 1002 600
rect 1036 566 1170 600
rect 1204 566 1242 600
rect 1276 566 1288 600
rect 918 560 1288 566
rect 1078 520 1438 532
rect 1078 486 1086 520
rect 1120 486 1398 520
rect 1432 486 1438 520
rect 1078 448 1438 486
rect 1078 414 1086 448
rect 1120 414 1398 448
rect 1432 414 1438 448
rect 1078 376 1438 414
rect 1078 342 1086 376
rect 1120 342 1398 376
rect 1432 342 1438 376
rect 1078 330 1438 342
rect 802 296 860 302
rect 802 262 814 296
rect 848 269 860 296
rect 1502 296 1560 302
rect 1502 269 1514 296
rect 848 262 1514 269
rect 1548 262 1560 296
rect 802 224 1560 262
rect 802 190 814 224
rect 848 190 1514 224
rect 1548 190 1560 224
rect 802 152 1560 190
rect 802 118 814 152
rect 848 118 1514 152
rect 1548 118 1560 152
rect 802 35 1560 118
rect 802 1 840 35
rect 874 1 919 35
rect 953 1 999 35
rect 1033 1 1079 35
rect 1113 1 1159 35
rect 1193 1 1239 35
rect 1273 1 1319 35
rect 1353 1 1399 35
rect 1433 1 1479 35
rect 1513 1 1560 35
rect 802 -5 1560 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1701704242
transform -1 0 262 0 -1 1102
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1701704242
transform 1 0 396 0 -1 1102
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1701704242
transform 1 0 890 0 -1 1102
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_3
timestamp 1701704242
transform 1 0 1130 0 -1 1102
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_4
timestamp 1701704242
transform 1 0 1442 0 -1 1102
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_5
timestamp 1701704242
transform 1 0 1285 0 -1 1028
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_6
timestamp 1701704242
transform 1 0 1046 0 -1 1028
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_7
timestamp 1701704242
transform 1 0 1170 0 -1 600
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_8
timestamp 1701704242
transform 1 0 930 0 -1 600
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_0
timestamp 1701704242
transform 0 -1 658 -1 0 1546
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_1
timestamp 1701704242
transform 0 -1 34 -1 0 1546
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_2
timestamp 1701704242
transform 0 -1 346 -1 0 1546
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_3
timestamp 1701704242
transform 0 -1 1120 -1 0 520
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_4
timestamp 1701704242
transform 0 -1 1432 -1 0 520
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_0
timestamp 1701704242
transform 1 0 814 0 -1 296
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_1
timestamp 1701704242
transform 1 0 1514 0 -1 296
box 0 0 1 1
use nfet_CDNS_524688791851195  nfet_CDNS_524688791851195_0
timestamp 1701704242
transform -1 0 1387 0 -1 709
box -79 -26 491 626
use pfet_CDNS_52468879185352  pfet_CDNS_52468879185352_0
timestamp 1701704242
transform 1 0 669 0 -1 1861
box -119 -66 219 1066
use pfet_CDNS_52468879185355  pfet_CDNS_52468879185355_0
timestamp 1701704242
transform 1 0 935 0 -1 1861
box -119 -66 687 1066
use pfet_CDNS_52468879185355  pfet_CDNS_52468879185355_1
timestamp 1701704242
transform 1 0 45 0 -1 1861
box -119 -66 687 1066
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_0
timestamp 1701704242
transform -1 0 735 0 1 679
box 0 0 1 1
use PYL1_CDNS_52468879185309  PYL1_CDNS_52468879185309_0
timestamp 1701704242
transform 0 1 914 1 0 763
box 0 0 1 1
use PYL1_CDNS_52468879185318  PYL1_CDNS_52468879185318_0
timestamp 1701704242
transform 0 -1 602 1 0 763
box 0 0 66 542
<< labels >>
flabel metal1 s 911 1087 911 1087 0 FreeSans 600 0 0 0 n<0>
flabel metal1 s 1085 483 1116 515 0 FreeSans 600 0 0 0 vgnd
port 1 nsew
flabel metal1 s 312 1441 343 1472 0 FreeSans 600 0 0 0 vcc_io
port 2 nsew
flabel locali s 978 779 1012 813 0 FreeSans 600 0 0 0 din
port 4 nsew
flabel locali s 333 779 367 813 0 FreeSans 600 0 0 0 ctl_in
port 5 nsew
flabel locali s 1242 779 1276 813 0 FreeSans 600 0 0 0 out
port 6 nsew
flabel locali s 685 779 719 813 0 FreeSans 600 0 0 0 ctl_in_n
port 7 nsew
<< properties >>
string GDS_END 85824686
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85816088
string path -0.650 48.800 39.325 48.800 
<< end >>
