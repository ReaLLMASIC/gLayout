magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< metal3 >>
rect 99 6053 4879 6096
rect 99 5817 4887 6053
rect 99 5447 4879 5817
rect 99 5211 4887 5447
rect 99 5168 4879 5211
rect 10078 5168 14858 6096
<< obsm3 >>
rect 99 11648 14858 40000
<< metal4 >>
rect 0 39983 254 40000
rect 0 39919 269 39983
rect 285 39919 349 39983
rect 365 39919 429 39983
rect 445 39919 509 39983
rect 525 39919 589 39983
rect 605 39919 669 39983
rect 685 39919 749 39983
rect 765 39919 829 39983
rect 845 39919 909 39983
rect 925 39919 989 39983
rect 1005 39919 1069 39983
rect 1085 39919 1149 39983
rect 1165 39919 1229 39983
rect 1245 39919 1309 39983
rect 1325 39919 1389 39983
rect 1405 39919 1469 39983
rect 1485 39919 1549 39983
rect 1565 39919 1629 39983
rect 1645 39919 1709 39983
rect 1725 39919 1789 39983
rect 1805 39919 1869 39983
rect 1885 39919 1949 39983
rect 1965 39919 2029 39983
rect 2045 39919 2109 39983
rect 2125 39919 2189 39983
rect 2205 39919 2269 39983
rect 2285 39919 2349 39983
rect 2365 39919 2429 39983
rect 2445 39919 2509 39983
rect 2525 39919 2589 39983
rect 2605 39919 2669 39983
rect 0 39902 254 39919
rect 0 39838 269 39902
rect 285 39838 349 39902
rect 365 39838 429 39902
rect 445 39838 509 39902
rect 525 39838 589 39902
rect 605 39838 669 39902
rect 685 39838 749 39902
rect 765 39838 829 39902
rect 845 39838 909 39902
rect 925 39838 989 39902
rect 1005 39838 1069 39902
rect 1085 39838 1149 39902
rect 1165 39838 1229 39902
rect 1245 39838 1309 39902
rect 1325 39838 1389 39902
rect 1405 39838 1469 39902
rect 1485 39838 1549 39902
rect 1565 39838 1629 39902
rect 1645 39838 1709 39902
rect 1725 39838 1789 39902
rect 1805 39838 1869 39902
rect 1885 39838 1949 39902
rect 1965 39838 2029 39902
rect 2045 39838 2109 39902
rect 2125 39838 2189 39902
rect 2205 39838 2269 39902
rect 2285 39838 2349 39902
rect 2365 39838 2429 39902
rect 2445 39838 2509 39902
rect 2525 39838 2589 39902
rect 2605 39838 2669 39902
rect 0 39821 254 39838
rect 0 39757 269 39821
rect 285 39757 349 39821
rect 365 39757 429 39821
rect 445 39757 509 39821
rect 525 39757 589 39821
rect 605 39757 669 39821
rect 685 39757 749 39821
rect 765 39757 829 39821
rect 845 39757 909 39821
rect 925 39757 989 39821
rect 1005 39757 1069 39821
rect 1085 39757 1149 39821
rect 1165 39757 1229 39821
rect 1245 39757 1309 39821
rect 1325 39757 1389 39821
rect 1405 39757 1469 39821
rect 1485 39757 1549 39821
rect 1565 39757 1629 39821
rect 1645 39757 1709 39821
rect 1725 39757 1789 39821
rect 1805 39757 1869 39821
rect 1885 39757 1949 39821
rect 1965 39757 2029 39821
rect 2045 39757 2109 39821
rect 2125 39757 2189 39821
rect 2205 39757 2269 39821
rect 2285 39757 2349 39821
rect 2365 39757 2429 39821
rect 2445 39757 2509 39821
rect 2525 39757 2589 39821
rect 2605 39757 2669 39821
rect 0 39740 254 39757
rect 0 39676 269 39740
rect 285 39676 349 39740
rect 365 39676 429 39740
rect 445 39676 509 39740
rect 525 39676 589 39740
rect 605 39676 669 39740
rect 685 39676 749 39740
rect 765 39676 829 39740
rect 845 39676 909 39740
rect 925 39676 989 39740
rect 1005 39676 1069 39740
rect 1085 39676 1149 39740
rect 1165 39676 1229 39740
rect 1245 39676 1309 39740
rect 1325 39676 1389 39740
rect 1405 39676 1469 39740
rect 1485 39676 1549 39740
rect 1565 39676 1629 39740
rect 1645 39676 1709 39740
rect 1725 39676 1789 39740
rect 1805 39676 1869 39740
rect 1885 39676 1949 39740
rect 1965 39676 2029 39740
rect 2045 39676 2109 39740
rect 2125 39676 2189 39740
rect 2205 39676 2269 39740
rect 2285 39676 2349 39740
rect 2365 39676 2429 39740
rect 2445 39676 2509 39740
rect 2525 39676 2589 39740
rect 2605 39676 2669 39740
rect 0 39659 254 39676
rect 0 39595 269 39659
rect 285 39595 349 39659
rect 365 39595 429 39659
rect 445 39595 509 39659
rect 525 39595 589 39659
rect 605 39595 669 39659
rect 685 39595 749 39659
rect 765 39595 829 39659
rect 845 39595 909 39659
rect 925 39595 989 39659
rect 1005 39595 1069 39659
rect 1085 39595 1149 39659
rect 1165 39595 1229 39659
rect 1245 39595 1309 39659
rect 1325 39595 1389 39659
rect 1405 39595 1469 39659
rect 1485 39595 1549 39659
rect 1565 39595 1629 39659
rect 1645 39595 1709 39659
rect 1725 39595 1789 39659
rect 1805 39595 1869 39659
rect 1885 39595 1949 39659
rect 1965 39595 2029 39659
rect 2045 39595 2109 39659
rect 2125 39595 2189 39659
rect 2205 39595 2269 39659
rect 2285 39595 2349 39659
rect 2365 39595 2429 39659
rect 2445 39595 2509 39659
rect 2525 39595 2589 39659
rect 2605 39595 2669 39659
rect 0 39578 254 39595
rect 0 39514 269 39578
rect 285 39514 349 39578
rect 365 39514 429 39578
rect 445 39514 509 39578
rect 525 39514 589 39578
rect 605 39514 669 39578
rect 685 39514 749 39578
rect 765 39514 829 39578
rect 845 39514 909 39578
rect 925 39514 989 39578
rect 1005 39514 1069 39578
rect 1085 39514 1149 39578
rect 1165 39514 1229 39578
rect 1245 39514 1309 39578
rect 1325 39514 1389 39578
rect 1405 39514 1469 39578
rect 1485 39514 1549 39578
rect 1565 39514 1629 39578
rect 1645 39514 1709 39578
rect 1725 39514 1789 39578
rect 1805 39514 1869 39578
rect 1885 39514 1949 39578
rect 1965 39514 2029 39578
rect 2045 39514 2109 39578
rect 2125 39514 2189 39578
rect 2205 39514 2269 39578
rect 2285 39514 2349 39578
rect 2365 39514 2429 39578
rect 2445 39514 2509 39578
rect 2525 39514 2589 39578
rect 2605 39514 2669 39578
rect 0 39497 254 39514
rect 0 39433 269 39497
rect 285 39433 349 39497
rect 365 39433 429 39497
rect 445 39433 509 39497
rect 525 39433 589 39497
rect 605 39433 669 39497
rect 685 39433 749 39497
rect 765 39433 829 39497
rect 845 39433 909 39497
rect 925 39433 989 39497
rect 1005 39433 1069 39497
rect 1085 39433 1149 39497
rect 1165 39433 1229 39497
rect 1245 39433 1309 39497
rect 1325 39433 1389 39497
rect 1405 39433 1469 39497
rect 1485 39433 1549 39497
rect 1565 39433 1629 39497
rect 1645 39433 1709 39497
rect 1725 39433 1789 39497
rect 1805 39433 1869 39497
rect 1885 39433 1949 39497
rect 1965 39433 2029 39497
rect 2045 39433 2109 39497
rect 2125 39433 2189 39497
rect 2205 39433 2269 39497
rect 2285 39433 2349 39497
rect 2365 39433 2429 39497
rect 2445 39433 2509 39497
rect 2525 39433 2589 39497
rect 2605 39433 2669 39497
rect 2726 39434 12265 39986
rect 14746 39983 15000 40000
rect 12306 39919 12370 39983
rect 12386 39919 12450 39983
rect 12466 39919 12530 39983
rect 12546 39919 12610 39983
rect 12626 39919 12690 39983
rect 12706 39919 12770 39983
rect 12786 39919 12850 39983
rect 12866 39919 12930 39983
rect 12946 39919 13010 39983
rect 13026 39919 13090 39983
rect 13106 39919 13170 39983
rect 13186 39919 13250 39983
rect 13266 39919 13330 39983
rect 13346 39919 13410 39983
rect 13426 39919 13490 39983
rect 13506 39919 13570 39983
rect 13586 39919 13650 39983
rect 13666 39919 13730 39983
rect 13746 39919 13810 39983
rect 13826 39919 13890 39983
rect 13906 39919 13970 39983
rect 13986 39919 14050 39983
rect 14066 39919 14130 39983
rect 14146 39919 14210 39983
rect 14226 39919 14290 39983
rect 14306 39919 14370 39983
rect 14386 39919 14450 39983
rect 14466 39919 14530 39983
rect 14546 39919 14610 39983
rect 14626 39919 14690 39983
rect 14706 39919 15000 39983
rect 14746 39902 15000 39919
rect 12306 39838 12370 39902
rect 12386 39838 12450 39902
rect 12466 39838 12530 39902
rect 12546 39838 12610 39902
rect 12626 39838 12690 39902
rect 12706 39838 12770 39902
rect 12786 39838 12850 39902
rect 12866 39838 12930 39902
rect 12946 39838 13010 39902
rect 13026 39838 13090 39902
rect 13106 39838 13170 39902
rect 13186 39838 13250 39902
rect 13266 39838 13330 39902
rect 13346 39838 13410 39902
rect 13426 39838 13490 39902
rect 13506 39838 13570 39902
rect 13586 39838 13650 39902
rect 13666 39838 13730 39902
rect 13746 39838 13810 39902
rect 13826 39838 13890 39902
rect 13906 39838 13970 39902
rect 13986 39838 14050 39902
rect 14066 39838 14130 39902
rect 14146 39838 14210 39902
rect 14226 39838 14290 39902
rect 14306 39838 14370 39902
rect 14386 39838 14450 39902
rect 14466 39838 14530 39902
rect 14546 39838 14610 39902
rect 14626 39838 14690 39902
rect 14706 39838 15000 39902
rect 14746 39821 15000 39838
rect 12306 39757 12370 39821
rect 12386 39757 12450 39821
rect 12466 39757 12530 39821
rect 12546 39757 12610 39821
rect 12626 39757 12690 39821
rect 12706 39757 12770 39821
rect 12786 39757 12850 39821
rect 12866 39757 12930 39821
rect 12946 39757 13010 39821
rect 13026 39757 13090 39821
rect 13106 39757 13170 39821
rect 13186 39757 13250 39821
rect 13266 39757 13330 39821
rect 13346 39757 13410 39821
rect 13426 39757 13490 39821
rect 13506 39757 13570 39821
rect 13586 39757 13650 39821
rect 13666 39757 13730 39821
rect 13746 39757 13810 39821
rect 13826 39757 13890 39821
rect 13906 39757 13970 39821
rect 13986 39757 14050 39821
rect 14066 39757 14130 39821
rect 14146 39757 14210 39821
rect 14226 39757 14290 39821
rect 14306 39757 14370 39821
rect 14386 39757 14450 39821
rect 14466 39757 14530 39821
rect 14546 39757 14610 39821
rect 14626 39757 14690 39821
rect 14706 39757 15000 39821
rect 14746 39740 15000 39757
rect 12306 39676 12370 39740
rect 12386 39676 12450 39740
rect 12466 39676 12530 39740
rect 12546 39676 12610 39740
rect 12626 39676 12690 39740
rect 12706 39676 12770 39740
rect 12786 39676 12850 39740
rect 12866 39676 12930 39740
rect 12946 39676 13010 39740
rect 13026 39676 13090 39740
rect 13106 39676 13170 39740
rect 13186 39676 13250 39740
rect 13266 39676 13330 39740
rect 13346 39676 13410 39740
rect 13426 39676 13490 39740
rect 13506 39676 13570 39740
rect 13586 39676 13650 39740
rect 13666 39676 13730 39740
rect 13746 39676 13810 39740
rect 13826 39676 13890 39740
rect 13906 39676 13970 39740
rect 13986 39676 14050 39740
rect 14066 39676 14130 39740
rect 14146 39676 14210 39740
rect 14226 39676 14290 39740
rect 14306 39676 14370 39740
rect 14386 39676 14450 39740
rect 14466 39676 14530 39740
rect 14546 39676 14610 39740
rect 14626 39676 14690 39740
rect 14706 39676 15000 39740
rect 14746 39659 15000 39676
rect 12306 39595 12370 39659
rect 12386 39595 12450 39659
rect 12466 39595 12530 39659
rect 12546 39595 12610 39659
rect 12626 39595 12690 39659
rect 12706 39595 12770 39659
rect 12786 39595 12850 39659
rect 12866 39595 12930 39659
rect 12946 39595 13010 39659
rect 13026 39595 13090 39659
rect 13106 39595 13170 39659
rect 13186 39595 13250 39659
rect 13266 39595 13330 39659
rect 13346 39595 13410 39659
rect 13426 39595 13490 39659
rect 13506 39595 13570 39659
rect 13586 39595 13650 39659
rect 13666 39595 13730 39659
rect 13746 39595 13810 39659
rect 13826 39595 13890 39659
rect 13906 39595 13970 39659
rect 13986 39595 14050 39659
rect 14066 39595 14130 39659
rect 14146 39595 14210 39659
rect 14226 39595 14290 39659
rect 14306 39595 14370 39659
rect 14386 39595 14450 39659
rect 14466 39595 14530 39659
rect 14546 39595 14610 39659
rect 14626 39595 14690 39659
rect 14706 39595 15000 39659
rect 14746 39578 15000 39595
rect 12306 39514 12370 39578
rect 12386 39514 12450 39578
rect 12466 39514 12530 39578
rect 12546 39514 12610 39578
rect 12626 39514 12690 39578
rect 12706 39514 12770 39578
rect 12786 39514 12850 39578
rect 12866 39514 12930 39578
rect 12946 39514 13010 39578
rect 13026 39514 13090 39578
rect 13106 39514 13170 39578
rect 13186 39514 13250 39578
rect 13266 39514 13330 39578
rect 13346 39514 13410 39578
rect 13426 39514 13490 39578
rect 13506 39514 13570 39578
rect 13586 39514 13650 39578
rect 13666 39514 13730 39578
rect 13746 39514 13810 39578
rect 13826 39514 13890 39578
rect 13906 39514 13970 39578
rect 13986 39514 14050 39578
rect 14066 39514 14130 39578
rect 14146 39514 14210 39578
rect 14226 39514 14290 39578
rect 14306 39514 14370 39578
rect 14386 39514 14450 39578
rect 14466 39514 14530 39578
rect 14546 39514 14610 39578
rect 14626 39514 14690 39578
rect 14706 39514 15000 39578
rect 14746 39497 15000 39514
rect 12306 39433 12370 39497
rect 12386 39433 12450 39497
rect 12466 39433 12530 39497
rect 12546 39433 12610 39497
rect 12626 39433 12690 39497
rect 12706 39433 12770 39497
rect 12786 39433 12850 39497
rect 12866 39433 12930 39497
rect 12946 39433 13010 39497
rect 13026 39433 13090 39497
rect 13106 39433 13170 39497
rect 13186 39433 13250 39497
rect 13266 39433 13330 39497
rect 13346 39433 13410 39497
rect 13426 39433 13490 39497
rect 13506 39433 13570 39497
rect 13586 39433 13650 39497
rect 13666 39433 13730 39497
rect 13746 39433 13810 39497
rect 13826 39433 13890 39497
rect 13906 39433 13970 39497
rect 13986 39433 14050 39497
rect 14066 39433 14130 39497
rect 14146 39433 14210 39497
rect 14226 39433 14290 39497
rect 14306 39433 14370 39497
rect 14386 39433 14450 39497
rect 14466 39433 14530 39497
rect 14546 39433 14610 39497
rect 14626 39433 14690 39497
rect 14706 39433 15000 39497
rect 0 39416 254 39433
rect 14746 39416 15000 39433
rect 0 39352 269 39416
rect 285 39352 349 39416
rect 365 39352 429 39416
rect 445 39352 509 39416
rect 525 39352 589 39416
rect 605 39352 669 39416
rect 685 39352 749 39416
rect 765 39352 829 39416
rect 845 39352 909 39416
rect 925 39352 989 39416
rect 1005 39352 1069 39416
rect 1085 39352 1149 39416
rect 1165 39352 1229 39416
rect 1245 39352 1309 39416
rect 1325 39352 1389 39416
rect 1405 39352 1469 39416
rect 1485 39352 1549 39416
rect 1565 39352 1629 39416
rect 1645 39352 1709 39416
rect 1725 39352 1789 39416
rect 1805 39352 1869 39416
rect 1885 39352 1949 39416
rect 1965 39352 2029 39416
rect 2045 39352 2109 39416
rect 2125 39352 2189 39416
rect 2205 39352 2269 39416
rect 2285 39352 2349 39416
rect 2365 39352 2429 39416
rect 2445 39352 2509 39416
rect 2525 39352 2589 39416
rect 2605 39352 2669 39416
rect 0 39335 254 39352
rect 0 39271 269 39335
rect 285 39271 349 39335
rect 365 39271 429 39335
rect 445 39271 509 39335
rect 525 39271 589 39335
rect 605 39271 669 39335
rect 685 39271 749 39335
rect 765 39271 829 39335
rect 845 39271 909 39335
rect 925 39271 989 39335
rect 1005 39271 1069 39335
rect 1085 39271 1149 39335
rect 1165 39271 1229 39335
rect 1245 39271 1309 39335
rect 1325 39271 1389 39335
rect 1405 39271 1469 39335
rect 1485 39271 1549 39335
rect 1565 39271 1629 39335
rect 1645 39271 1709 39335
rect 1725 39271 1789 39335
rect 1805 39271 1869 39335
rect 1885 39271 1949 39335
rect 1965 39271 2029 39335
rect 2045 39271 2109 39335
rect 2125 39271 2189 39335
rect 2205 39271 2269 39335
rect 2285 39271 2349 39335
rect 2365 39271 2429 39335
rect 2445 39271 2509 39335
rect 2525 39271 2589 39335
rect 2605 39271 2669 39335
rect 0 39254 254 39271
rect 0 39190 269 39254
rect 285 39190 349 39254
rect 365 39190 429 39254
rect 445 39190 509 39254
rect 525 39190 589 39254
rect 605 39190 669 39254
rect 685 39190 749 39254
rect 765 39190 829 39254
rect 845 39190 909 39254
rect 925 39190 989 39254
rect 1005 39190 1069 39254
rect 1085 39190 1149 39254
rect 1165 39190 1229 39254
rect 1245 39190 1309 39254
rect 1325 39190 1389 39254
rect 1405 39190 1469 39254
rect 1485 39190 1549 39254
rect 1565 39190 1629 39254
rect 1645 39190 1709 39254
rect 1725 39190 1789 39254
rect 1805 39190 1869 39254
rect 1885 39190 1949 39254
rect 1965 39190 2029 39254
rect 2045 39190 2109 39254
rect 2125 39190 2189 39254
rect 2205 39190 2269 39254
rect 2285 39190 2349 39254
rect 2365 39190 2429 39254
rect 2445 39190 2509 39254
rect 2525 39190 2589 39254
rect 2605 39190 2669 39254
rect 2719 39246 2851 39394
rect 0 39173 254 39190
rect 0 39109 269 39173
rect 285 39109 349 39173
rect 365 39109 429 39173
rect 445 39109 509 39173
rect 525 39109 589 39173
rect 605 39109 669 39173
rect 685 39109 749 39173
rect 765 39109 829 39173
rect 845 39109 909 39173
rect 925 39109 989 39173
rect 1005 39109 1069 39173
rect 1085 39109 1149 39173
rect 1165 39109 1229 39173
rect 1245 39109 1309 39173
rect 1325 39109 1389 39173
rect 1405 39109 1469 39173
rect 1485 39109 1549 39173
rect 1565 39109 1629 39173
rect 1645 39109 1709 39173
rect 1725 39109 1789 39173
rect 1805 39109 1869 39173
rect 1885 39109 1949 39173
rect 1965 39109 2029 39173
rect 2045 39109 2109 39173
rect 2125 39109 2189 39173
rect 2205 39109 2269 39173
rect 2285 39109 2349 39173
rect 2365 39109 2429 39173
rect 2445 39109 2509 39173
rect 2525 39109 2589 39173
rect 2605 39109 2669 39173
rect 12136 39246 12268 39394
rect 12306 39352 12370 39416
rect 12386 39352 12450 39416
rect 12466 39352 12530 39416
rect 12546 39352 12610 39416
rect 12626 39352 12690 39416
rect 12706 39352 12770 39416
rect 12786 39352 12850 39416
rect 12866 39352 12930 39416
rect 12946 39352 13010 39416
rect 13026 39352 13090 39416
rect 13106 39352 13170 39416
rect 13186 39352 13250 39416
rect 13266 39352 13330 39416
rect 13346 39352 13410 39416
rect 13426 39352 13490 39416
rect 13506 39352 13570 39416
rect 13586 39352 13650 39416
rect 13666 39352 13730 39416
rect 13746 39352 13810 39416
rect 13826 39352 13890 39416
rect 13906 39352 13970 39416
rect 13986 39352 14050 39416
rect 14066 39352 14130 39416
rect 14146 39352 14210 39416
rect 14226 39352 14290 39416
rect 14306 39352 14370 39416
rect 14386 39352 14450 39416
rect 14466 39352 14530 39416
rect 14546 39352 14610 39416
rect 14626 39352 14690 39416
rect 14706 39352 15000 39416
rect 14746 39335 15000 39352
rect 12306 39271 12370 39335
rect 12386 39271 12450 39335
rect 12466 39271 12530 39335
rect 12546 39271 12610 39335
rect 12626 39271 12690 39335
rect 12706 39271 12770 39335
rect 12786 39271 12850 39335
rect 12866 39271 12930 39335
rect 12946 39271 13010 39335
rect 13026 39271 13090 39335
rect 13106 39271 13170 39335
rect 13186 39271 13250 39335
rect 13266 39271 13330 39335
rect 13346 39271 13410 39335
rect 13426 39271 13490 39335
rect 13506 39271 13570 39335
rect 13586 39271 13650 39335
rect 13666 39271 13730 39335
rect 13746 39271 13810 39335
rect 13826 39271 13890 39335
rect 13906 39271 13970 39335
rect 13986 39271 14050 39335
rect 14066 39271 14130 39335
rect 14146 39271 14210 39335
rect 14226 39271 14290 39335
rect 14306 39271 14370 39335
rect 14386 39271 14450 39335
rect 14466 39271 14530 39335
rect 14546 39271 14610 39335
rect 14626 39271 14690 39335
rect 14706 39271 15000 39335
rect 14746 39254 15000 39271
rect 12306 39190 12370 39254
rect 12386 39190 12450 39254
rect 12466 39190 12530 39254
rect 12546 39190 12610 39254
rect 12626 39190 12690 39254
rect 12706 39190 12770 39254
rect 12786 39190 12850 39254
rect 12866 39190 12930 39254
rect 12946 39190 13010 39254
rect 13026 39190 13090 39254
rect 13106 39190 13170 39254
rect 13186 39190 13250 39254
rect 13266 39190 13330 39254
rect 13346 39190 13410 39254
rect 13426 39190 13490 39254
rect 13506 39190 13570 39254
rect 13586 39190 13650 39254
rect 13666 39190 13730 39254
rect 13746 39190 13810 39254
rect 13826 39190 13890 39254
rect 13906 39190 13970 39254
rect 13986 39190 14050 39254
rect 14066 39190 14130 39254
rect 14146 39190 14210 39254
rect 14226 39190 14290 39254
rect 14306 39190 14370 39254
rect 14386 39190 14450 39254
rect 14466 39190 14530 39254
rect 14546 39190 14610 39254
rect 14626 39190 14690 39254
rect 14706 39190 15000 39254
rect 14746 39173 15000 39190
rect 12306 39109 12370 39173
rect 12386 39109 12450 39173
rect 12466 39109 12530 39173
rect 12546 39109 12610 39173
rect 12626 39109 12690 39173
rect 12706 39109 12770 39173
rect 12786 39109 12850 39173
rect 12866 39109 12930 39173
rect 12946 39109 13010 39173
rect 13026 39109 13090 39173
rect 13106 39109 13170 39173
rect 13186 39109 13250 39173
rect 13266 39109 13330 39173
rect 13346 39109 13410 39173
rect 13426 39109 13490 39173
rect 13506 39109 13570 39173
rect 13586 39109 13650 39173
rect 13666 39109 13730 39173
rect 13746 39109 13810 39173
rect 13826 39109 13890 39173
rect 13906 39109 13970 39173
rect 13986 39109 14050 39173
rect 14066 39109 14130 39173
rect 14146 39109 14210 39173
rect 14226 39109 14290 39173
rect 14306 39109 14370 39173
rect 14386 39109 14450 39173
rect 14466 39109 14530 39173
rect 14546 39109 14610 39173
rect 14626 39109 14690 39173
rect 14706 39109 15000 39173
rect 0 39092 254 39109
rect 14746 39092 15000 39109
rect 0 39028 269 39092
rect 285 39028 349 39092
rect 365 39028 429 39092
rect 445 39028 509 39092
rect 525 39028 589 39092
rect 605 39028 669 39092
rect 685 39028 749 39092
rect 765 39028 829 39092
rect 845 39028 909 39092
rect 925 39028 989 39092
rect 1005 39028 1069 39092
rect 1085 39028 1149 39092
rect 1165 39028 1229 39092
rect 1245 39028 1309 39092
rect 1325 39028 1389 39092
rect 1405 39028 1469 39092
rect 1485 39028 1549 39092
rect 1565 39028 1629 39092
rect 1645 39028 1709 39092
rect 1725 39028 1789 39092
rect 1805 39028 1869 39092
rect 1885 39028 1949 39092
rect 1965 39028 2029 39092
rect 2045 39028 2109 39092
rect 2125 39028 2189 39092
rect 2205 39028 2269 39092
rect 2285 39028 2349 39092
rect 2365 39028 2429 39092
rect 2445 39028 2509 39092
rect 2525 39028 2589 39092
rect 2605 39028 2669 39092
rect 12306 39028 12370 39092
rect 12386 39028 12450 39092
rect 12466 39028 12530 39092
rect 12546 39028 12610 39092
rect 12626 39028 12690 39092
rect 12706 39028 12770 39092
rect 12786 39028 12850 39092
rect 12866 39028 12930 39092
rect 12946 39028 13010 39092
rect 13026 39028 13090 39092
rect 13106 39028 13170 39092
rect 13186 39028 13250 39092
rect 13266 39028 13330 39092
rect 13346 39028 13410 39092
rect 13426 39028 13490 39092
rect 13506 39028 13570 39092
rect 13586 39028 13650 39092
rect 13666 39028 13730 39092
rect 13746 39028 13810 39092
rect 13826 39028 13890 39092
rect 13906 39028 13970 39092
rect 13986 39028 14050 39092
rect 14066 39028 14130 39092
rect 14146 39028 14210 39092
rect 14226 39028 14290 39092
rect 14306 39028 14370 39092
rect 14386 39028 14450 39092
rect 14466 39028 14530 39092
rect 14546 39028 14610 39092
rect 14626 39028 14690 39092
rect 14706 39028 15000 39092
rect 0 39011 254 39028
rect 14746 39011 15000 39028
rect 0 35187 2669 39011
rect 12306 35187 15000 39011
rect 0 35157 254 35187
rect 14746 35157 15000 35187
rect 0 14007 254 19000
rect 14746 14007 15000 19000
rect 0 12817 254 13707
rect 14746 12817 15000 13707
rect 0 11647 254 12537
rect 14746 12534 15000 12537
rect 269 12470 333 12534
rect 351 12470 415 12534
rect 433 12470 497 12534
rect 515 12470 579 12534
rect 597 12470 661 12534
rect 678 12470 742 12534
rect 759 12470 823 12534
rect 840 12470 904 12534
rect 921 12470 985 12534
rect 1002 12470 1066 12534
rect 1083 12470 1147 12534
rect 1164 12470 1228 12534
rect 1245 12470 1309 12534
rect 1326 12470 1390 12534
rect 1407 12470 1471 12534
rect 1488 12470 1552 12534
rect 1569 12470 1633 12534
rect 1650 12470 1714 12534
rect 1731 12470 1795 12534
rect 1812 12470 1876 12534
rect 1893 12470 1957 12534
rect 1974 12470 2038 12534
rect 2055 12470 2119 12534
rect 2136 12470 2200 12534
rect 2217 12470 2281 12534
rect 2298 12470 2362 12534
rect 2379 12470 2443 12534
rect 2460 12470 2524 12534
rect 2541 12470 2605 12534
rect 2622 12470 2686 12534
rect 2703 12470 2767 12534
rect 2784 12470 2848 12534
rect 2865 12470 2929 12534
rect 2946 12470 3010 12534
rect 3027 12470 3091 12534
rect 3108 12470 3172 12534
rect 3189 12470 3253 12534
rect 3270 12470 3334 12534
rect 3351 12470 3415 12534
rect 3432 12470 3496 12534
rect 3513 12470 3577 12534
rect 3594 12470 3658 12534
rect 3675 12470 3739 12534
rect 3756 12470 3820 12534
rect 3837 12470 3901 12534
rect 3918 12470 3982 12534
rect 3999 12470 4063 12534
rect 4080 12470 4144 12534
rect 4161 12470 4225 12534
rect 4242 12470 4306 12534
rect 4323 12470 4387 12534
rect 4404 12470 4468 12534
rect 4485 12470 4549 12534
rect 4566 12470 4630 12534
rect 4647 12470 4711 12534
rect 4728 12470 4792 12534
rect 4809 12470 4873 12534
rect 10084 12470 10148 12534
rect 10166 12470 10230 12534
rect 10248 12470 10312 12534
rect 10330 12470 10394 12534
rect 10412 12470 10476 12534
rect 10494 12470 10558 12534
rect 10576 12470 10640 12534
rect 10657 12470 10721 12534
rect 10738 12470 10802 12534
rect 10819 12470 10883 12534
rect 10900 12470 10964 12534
rect 10981 12470 11045 12534
rect 11062 12470 11126 12534
rect 11143 12470 11207 12534
rect 11224 12470 11288 12534
rect 11305 12470 11369 12534
rect 11386 12470 11450 12534
rect 11467 12470 11531 12534
rect 11548 12470 11612 12534
rect 11629 12470 11693 12534
rect 11710 12470 11774 12534
rect 11791 12470 11855 12534
rect 11872 12470 11936 12534
rect 11953 12470 12017 12534
rect 12034 12470 12098 12534
rect 12115 12470 12179 12534
rect 12196 12470 12260 12534
rect 12277 12470 12341 12534
rect 12358 12470 12422 12534
rect 12439 12470 12503 12534
rect 12520 12470 12584 12534
rect 12601 12470 12665 12534
rect 12682 12470 12746 12534
rect 12763 12470 12827 12534
rect 12844 12470 12908 12534
rect 12925 12470 12989 12534
rect 13006 12470 13070 12534
rect 13087 12470 13151 12534
rect 13168 12470 13232 12534
rect 13249 12470 13313 12534
rect 13330 12470 13394 12534
rect 13411 12470 13475 12534
rect 13492 12470 13556 12534
rect 13573 12470 13637 12534
rect 13654 12470 13718 12534
rect 13735 12470 13799 12534
rect 13816 12470 13880 12534
rect 13897 12470 13961 12534
rect 13978 12470 14042 12534
rect 14059 12470 14123 12534
rect 14140 12470 14204 12534
rect 14221 12470 14285 12534
rect 14302 12470 14366 12534
rect 14383 12470 14447 12534
rect 14464 12470 14528 12534
rect 14545 12470 14609 12534
rect 14626 12470 14690 12534
rect 14707 12470 15000 12534
rect 14746 12452 15000 12470
rect 269 12388 333 12452
rect 351 12388 415 12452
rect 433 12388 497 12452
rect 515 12388 579 12452
rect 597 12388 661 12452
rect 678 12388 742 12452
rect 759 12388 823 12452
rect 840 12388 904 12452
rect 921 12388 985 12452
rect 1002 12388 1066 12452
rect 1083 12388 1147 12452
rect 1164 12388 1228 12452
rect 1245 12388 1309 12452
rect 1326 12388 1390 12452
rect 1407 12388 1471 12452
rect 1488 12388 1552 12452
rect 1569 12388 1633 12452
rect 1650 12388 1714 12452
rect 1731 12388 1795 12452
rect 1812 12388 1876 12452
rect 1893 12388 1957 12452
rect 1974 12388 2038 12452
rect 2055 12388 2119 12452
rect 2136 12388 2200 12452
rect 2217 12388 2281 12452
rect 2298 12388 2362 12452
rect 2379 12388 2443 12452
rect 2460 12388 2524 12452
rect 2541 12388 2605 12452
rect 2622 12388 2686 12452
rect 2703 12388 2767 12452
rect 2784 12388 2848 12452
rect 2865 12388 2929 12452
rect 2946 12388 3010 12452
rect 3027 12388 3091 12452
rect 3108 12388 3172 12452
rect 3189 12388 3253 12452
rect 3270 12388 3334 12452
rect 3351 12388 3415 12452
rect 3432 12388 3496 12452
rect 3513 12388 3577 12452
rect 3594 12388 3658 12452
rect 3675 12388 3739 12452
rect 3756 12388 3820 12452
rect 3837 12388 3901 12452
rect 3918 12388 3982 12452
rect 3999 12388 4063 12452
rect 4080 12388 4144 12452
rect 4161 12388 4225 12452
rect 4242 12388 4306 12452
rect 4323 12388 4387 12452
rect 4404 12388 4468 12452
rect 4485 12388 4549 12452
rect 4566 12388 4630 12452
rect 4647 12388 4711 12452
rect 4728 12388 4792 12452
rect 4809 12388 4873 12452
rect 10084 12388 10148 12452
rect 10166 12388 10230 12452
rect 10248 12388 10312 12452
rect 10330 12388 10394 12452
rect 10412 12388 10476 12452
rect 10494 12388 10558 12452
rect 10576 12388 10640 12452
rect 10657 12388 10721 12452
rect 10738 12388 10802 12452
rect 10819 12388 10883 12452
rect 10900 12388 10964 12452
rect 10981 12388 11045 12452
rect 11062 12388 11126 12452
rect 11143 12388 11207 12452
rect 11224 12388 11288 12452
rect 11305 12388 11369 12452
rect 11386 12388 11450 12452
rect 11467 12388 11531 12452
rect 11548 12388 11612 12452
rect 11629 12388 11693 12452
rect 11710 12388 11774 12452
rect 11791 12388 11855 12452
rect 11872 12388 11936 12452
rect 11953 12388 12017 12452
rect 12034 12388 12098 12452
rect 12115 12388 12179 12452
rect 12196 12388 12260 12452
rect 12277 12388 12341 12452
rect 12358 12388 12422 12452
rect 12439 12388 12503 12452
rect 12520 12388 12584 12452
rect 12601 12388 12665 12452
rect 12682 12388 12746 12452
rect 12763 12388 12827 12452
rect 12844 12388 12908 12452
rect 12925 12388 12989 12452
rect 13006 12388 13070 12452
rect 13087 12388 13151 12452
rect 13168 12388 13232 12452
rect 13249 12388 13313 12452
rect 13330 12388 13394 12452
rect 13411 12388 13475 12452
rect 13492 12388 13556 12452
rect 13573 12388 13637 12452
rect 13654 12388 13718 12452
rect 13735 12388 13799 12452
rect 13816 12388 13880 12452
rect 13897 12388 13961 12452
rect 13978 12388 14042 12452
rect 14059 12388 14123 12452
rect 14140 12388 14204 12452
rect 14221 12388 14285 12452
rect 14302 12388 14366 12452
rect 14383 12388 14447 12452
rect 14464 12388 14528 12452
rect 14545 12388 14609 12452
rect 14626 12388 14690 12452
rect 14707 12388 15000 12452
rect 14746 12370 15000 12388
rect 269 12306 333 12370
rect 351 12306 415 12370
rect 433 12306 497 12370
rect 515 12306 579 12370
rect 597 12306 661 12370
rect 678 12306 742 12370
rect 759 12306 823 12370
rect 840 12306 904 12370
rect 921 12306 985 12370
rect 1002 12306 1066 12370
rect 1083 12306 1147 12370
rect 1164 12306 1228 12370
rect 1245 12306 1309 12370
rect 1326 12306 1390 12370
rect 1407 12306 1471 12370
rect 1488 12306 1552 12370
rect 1569 12306 1633 12370
rect 1650 12306 1714 12370
rect 1731 12306 1795 12370
rect 1812 12306 1876 12370
rect 1893 12306 1957 12370
rect 1974 12306 2038 12370
rect 2055 12306 2119 12370
rect 2136 12306 2200 12370
rect 2217 12306 2281 12370
rect 2298 12306 2362 12370
rect 2379 12306 2443 12370
rect 2460 12306 2524 12370
rect 2541 12306 2605 12370
rect 2622 12306 2686 12370
rect 2703 12306 2767 12370
rect 2784 12306 2848 12370
rect 2865 12306 2929 12370
rect 2946 12306 3010 12370
rect 3027 12306 3091 12370
rect 3108 12306 3172 12370
rect 3189 12306 3253 12370
rect 3270 12306 3334 12370
rect 3351 12306 3415 12370
rect 3432 12306 3496 12370
rect 3513 12306 3577 12370
rect 3594 12306 3658 12370
rect 3675 12306 3739 12370
rect 3756 12306 3820 12370
rect 3837 12306 3901 12370
rect 3918 12306 3982 12370
rect 3999 12306 4063 12370
rect 4080 12306 4144 12370
rect 4161 12306 4225 12370
rect 4242 12306 4306 12370
rect 4323 12306 4387 12370
rect 4404 12306 4468 12370
rect 4485 12306 4549 12370
rect 4566 12306 4630 12370
rect 4647 12306 4711 12370
rect 4728 12306 4792 12370
rect 4809 12306 4873 12370
rect 10084 12306 10148 12370
rect 10166 12306 10230 12370
rect 10248 12306 10312 12370
rect 10330 12306 10394 12370
rect 10412 12306 10476 12370
rect 10494 12306 10558 12370
rect 10576 12306 10640 12370
rect 10657 12306 10721 12370
rect 10738 12306 10802 12370
rect 10819 12306 10883 12370
rect 10900 12306 10964 12370
rect 10981 12306 11045 12370
rect 11062 12306 11126 12370
rect 11143 12306 11207 12370
rect 11224 12306 11288 12370
rect 11305 12306 11369 12370
rect 11386 12306 11450 12370
rect 11467 12306 11531 12370
rect 11548 12306 11612 12370
rect 11629 12306 11693 12370
rect 11710 12306 11774 12370
rect 11791 12306 11855 12370
rect 11872 12306 11936 12370
rect 11953 12306 12017 12370
rect 12034 12306 12098 12370
rect 12115 12306 12179 12370
rect 12196 12306 12260 12370
rect 12277 12306 12341 12370
rect 12358 12306 12422 12370
rect 12439 12306 12503 12370
rect 12520 12306 12584 12370
rect 12601 12306 12665 12370
rect 12682 12306 12746 12370
rect 12763 12306 12827 12370
rect 12844 12306 12908 12370
rect 12925 12306 12989 12370
rect 13006 12306 13070 12370
rect 13087 12306 13151 12370
rect 13168 12306 13232 12370
rect 13249 12306 13313 12370
rect 13330 12306 13394 12370
rect 13411 12306 13475 12370
rect 13492 12306 13556 12370
rect 13573 12306 13637 12370
rect 13654 12306 13718 12370
rect 13735 12306 13799 12370
rect 13816 12306 13880 12370
rect 13897 12306 13961 12370
rect 13978 12306 14042 12370
rect 14059 12306 14123 12370
rect 14140 12306 14204 12370
rect 14221 12306 14285 12370
rect 14302 12306 14366 12370
rect 14383 12306 14447 12370
rect 14464 12306 14528 12370
rect 14545 12306 14609 12370
rect 14626 12306 14690 12370
rect 14707 12306 15000 12370
rect 14746 12288 15000 12306
rect 269 12224 333 12288
rect 351 12224 415 12288
rect 433 12224 497 12288
rect 515 12224 579 12288
rect 597 12224 661 12288
rect 678 12224 742 12288
rect 759 12224 823 12288
rect 840 12224 904 12288
rect 921 12224 985 12288
rect 1002 12224 1066 12288
rect 1083 12224 1147 12288
rect 1164 12224 1228 12288
rect 1245 12224 1309 12288
rect 1326 12224 1390 12288
rect 1407 12224 1471 12288
rect 1488 12224 1552 12288
rect 1569 12224 1633 12288
rect 1650 12224 1714 12288
rect 1731 12224 1795 12288
rect 1812 12224 1876 12288
rect 1893 12224 1957 12288
rect 1974 12224 2038 12288
rect 2055 12224 2119 12288
rect 2136 12224 2200 12288
rect 2217 12224 2281 12288
rect 2298 12224 2362 12288
rect 2379 12224 2443 12288
rect 2460 12224 2524 12288
rect 2541 12224 2605 12288
rect 2622 12224 2686 12288
rect 2703 12224 2767 12288
rect 2784 12224 2848 12288
rect 2865 12224 2929 12288
rect 2946 12224 3010 12288
rect 3027 12224 3091 12288
rect 3108 12224 3172 12288
rect 3189 12224 3253 12288
rect 3270 12224 3334 12288
rect 3351 12224 3415 12288
rect 3432 12224 3496 12288
rect 3513 12224 3577 12288
rect 3594 12224 3658 12288
rect 3675 12224 3739 12288
rect 3756 12224 3820 12288
rect 3837 12224 3901 12288
rect 3918 12224 3982 12288
rect 3999 12224 4063 12288
rect 4080 12224 4144 12288
rect 4161 12224 4225 12288
rect 4242 12224 4306 12288
rect 4323 12224 4387 12288
rect 4404 12224 4468 12288
rect 4485 12224 4549 12288
rect 4566 12224 4630 12288
rect 4647 12224 4711 12288
rect 4728 12224 4792 12288
rect 4809 12224 4873 12288
rect 10084 12224 10148 12288
rect 10166 12224 10230 12288
rect 10248 12224 10312 12288
rect 10330 12224 10394 12288
rect 10412 12224 10476 12288
rect 10494 12224 10558 12288
rect 10576 12224 10640 12288
rect 10657 12224 10721 12288
rect 10738 12224 10802 12288
rect 10819 12224 10883 12288
rect 10900 12224 10964 12288
rect 10981 12224 11045 12288
rect 11062 12224 11126 12288
rect 11143 12224 11207 12288
rect 11224 12224 11288 12288
rect 11305 12224 11369 12288
rect 11386 12224 11450 12288
rect 11467 12224 11531 12288
rect 11548 12224 11612 12288
rect 11629 12224 11693 12288
rect 11710 12224 11774 12288
rect 11791 12224 11855 12288
rect 11872 12224 11936 12288
rect 11953 12224 12017 12288
rect 12034 12224 12098 12288
rect 12115 12224 12179 12288
rect 12196 12224 12260 12288
rect 12277 12224 12341 12288
rect 12358 12224 12422 12288
rect 12439 12224 12503 12288
rect 12520 12224 12584 12288
rect 12601 12224 12665 12288
rect 12682 12224 12746 12288
rect 12763 12224 12827 12288
rect 12844 12224 12908 12288
rect 12925 12224 12989 12288
rect 13006 12224 13070 12288
rect 13087 12224 13151 12288
rect 13168 12224 13232 12288
rect 13249 12224 13313 12288
rect 13330 12224 13394 12288
rect 13411 12224 13475 12288
rect 13492 12224 13556 12288
rect 13573 12224 13637 12288
rect 13654 12224 13718 12288
rect 13735 12224 13799 12288
rect 13816 12224 13880 12288
rect 13897 12224 13961 12288
rect 13978 12224 14042 12288
rect 14059 12224 14123 12288
rect 14140 12224 14204 12288
rect 14221 12224 14285 12288
rect 14302 12224 14366 12288
rect 14383 12224 14447 12288
rect 14464 12224 14528 12288
rect 14545 12224 14609 12288
rect 14626 12224 14690 12288
rect 14707 12224 15000 12288
rect 14746 12206 15000 12224
rect 269 12142 333 12206
rect 351 12142 415 12206
rect 433 12142 497 12206
rect 515 12142 579 12206
rect 597 12142 661 12206
rect 678 12142 742 12206
rect 759 12142 823 12206
rect 840 12142 904 12206
rect 921 12142 985 12206
rect 1002 12142 1066 12206
rect 1083 12142 1147 12206
rect 1164 12142 1228 12206
rect 1245 12142 1309 12206
rect 1326 12142 1390 12206
rect 1407 12142 1471 12206
rect 1488 12142 1552 12206
rect 1569 12142 1633 12206
rect 1650 12142 1714 12206
rect 1731 12142 1795 12206
rect 1812 12142 1876 12206
rect 1893 12142 1957 12206
rect 1974 12142 2038 12206
rect 2055 12142 2119 12206
rect 2136 12142 2200 12206
rect 2217 12142 2281 12206
rect 2298 12142 2362 12206
rect 2379 12142 2443 12206
rect 2460 12142 2524 12206
rect 2541 12142 2605 12206
rect 2622 12142 2686 12206
rect 2703 12142 2767 12206
rect 2784 12142 2848 12206
rect 2865 12142 2929 12206
rect 2946 12142 3010 12206
rect 3027 12142 3091 12206
rect 3108 12142 3172 12206
rect 3189 12142 3253 12206
rect 3270 12142 3334 12206
rect 3351 12142 3415 12206
rect 3432 12142 3496 12206
rect 3513 12142 3577 12206
rect 3594 12142 3658 12206
rect 3675 12142 3739 12206
rect 3756 12142 3820 12206
rect 3837 12142 3901 12206
rect 3918 12142 3982 12206
rect 3999 12142 4063 12206
rect 4080 12142 4144 12206
rect 4161 12142 4225 12206
rect 4242 12142 4306 12206
rect 4323 12142 4387 12206
rect 4404 12142 4468 12206
rect 4485 12142 4549 12206
rect 4566 12142 4630 12206
rect 4647 12142 4711 12206
rect 4728 12142 4792 12206
rect 4809 12142 4873 12206
rect 10084 12142 10148 12206
rect 10166 12142 10230 12206
rect 10248 12142 10312 12206
rect 10330 12142 10394 12206
rect 10412 12142 10476 12206
rect 10494 12142 10558 12206
rect 10576 12142 10640 12206
rect 10657 12142 10721 12206
rect 10738 12142 10802 12206
rect 10819 12142 10883 12206
rect 10900 12142 10964 12206
rect 10981 12142 11045 12206
rect 11062 12142 11126 12206
rect 11143 12142 11207 12206
rect 11224 12142 11288 12206
rect 11305 12142 11369 12206
rect 11386 12142 11450 12206
rect 11467 12142 11531 12206
rect 11548 12142 11612 12206
rect 11629 12142 11693 12206
rect 11710 12142 11774 12206
rect 11791 12142 11855 12206
rect 11872 12142 11936 12206
rect 11953 12142 12017 12206
rect 12034 12142 12098 12206
rect 12115 12142 12179 12206
rect 12196 12142 12260 12206
rect 12277 12142 12341 12206
rect 12358 12142 12422 12206
rect 12439 12142 12503 12206
rect 12520 12142 12584 12206
rect 12601 12142 12665 12206
rect 12682 12142 12746 12206
rect 12763 12142 12827 12206
rect 12844 12142 12908 12206
rect 12925 12142 12989 12206
rect 13006 12142 13070 12206
rect 13087 12142 13151 12206
rect 13168 12142 13232 12206
rect 13249 12142 13313 12206
rect 13330 12142 13394 12206
rect 13411 12142 13475 12206
rect 13492 12142 13556 12206
rect 13573 12142 13637 12206
rect 13654 12142 13718 12206
rect 13735 12142 13799 12206
rect 13816 12142 13880 12206
rect 13897 12142 13961 12206
rect 13978 12142 14042 12206
rect 14059 12142 14123 12206
rect 14140 12142 14204 12206
rect 14221 12142 14285 12206
rect 14302 12142 14366 12206
rect 14383 12142 14447 12206
rect 14464 12142 14528 12206
rect 14545 12142 14609 12206
rect 14626 12142 14690 12206
rect 14707 12142 15000 12206
rect 14746 12124 15000 12142
rect 269 12060 333 12124
rect 351 12060 415 12124
rect 433 12060 497 12124
rect 515 12060 579 12124
rect 597 12060 661 12124
rect 678 12060 742 12124
rect 759 12060 823 12124
rect 840 12060 904 12124
rect 921 12060 985 12124
rect 1002 12060 1066 12124
rect 1083 12060 1147 12124
rect 1164 12060 1228 12124
rect 1245 12060 1309 12124
rect 1326 12060 1390 12124
rect 1407 12060 1471 12124
rect 1488 12060 1552 12124
rect 1569 12060 1633 12124
rect 1650 12060 1714 12124
rect 1731 12060 1795 12124
rect 1812 12060 1876 12124
rect 1893 12060 1957 12124
rect 1974 12060 2038 12124
rect 2055 12060 2119 12124
rect 2136 12060 2200 12124
rect 2217 12060 2281 12124
rect 2298 12060 2362 12124
rect 2379 12060 2443 12124
rect 2460 12060 2524 12124
rect 2541 12060 2605 12124
rect 2622 12060 2686 12124
rect 2703 12060 2767 12124
rect 2784 12060 2848 12124
rect 2865 12060 2929 12124
rect 2946 12060 3010 12124
rect 3027 12060 3091 12124
rect 3108 12060 3172 12124
rect 3189 12060 3253 12124
rect 3270 12060 3334 12124
rect 3351 12060 3415 12124
rect 3432 12060 3496 12124
rect 3513 12060 3577 12124
rect 3594 12060 3658 12124
rect 3675 12060 3739 12124
rect 3756 12060 3820 12124
rect 3837 12060 3901 12124
rect 3918 12060 3982 12124
rect 3999 12060 4063 12124
rect 4080 12060 4144 12124
rect 4161 12060 4225 12124
rect 4242 12060 4306 12124
rect 4323 12060 4387 12124
rect 4404 12060 4468 12124
rect 4485 12060 4549 12124
rect 4566 12060 4630 12124
rect 4647 12060 4711 12124
rect 4728 12060 4792 12124
rect 4809 12060 4873 12124
rect 10084 12060 10148 12124
rect 10166 12060 10230 12124
rect 10248 12060 10312 12124
rect 10330 12060 10394 12124
rect 10412 12060 10476 12124
rect 10494 12060 10558 12124
rect 10576 12060 10640 12124
rect 10657 12060 10721 12124
rect 10738 12060 10802 12124
rect 10819 12060 10883 12124
rect 10900 12060 10964 12124
rect 10981 12060 11045 12124
rect 11062 12060 11126 12124
rect 11143 12060 11207 12124
rect 11224 12060 11288 12124
rect 11305 12060 11369 12124
rect 11386 12060 11450 12124
rect 11467 12060 11531 12124
rect 11548 12060 11612 12124
rect 11629 12060 11693 12124
rect 11710 12060 11774 12124
rect 11791 12060 11855 12124
rect 11872 12060 11936 12124
rect 11953 12060 12017 12124
rect 12034 12060 12098 12124
rect 12115 12060 12179 12124
rect 12196 12060 12260 12124
rect 12277 12060 12341 12124
rect 12358 12060 12422 12124
rect 12439 12060 12503 12124
rect 12520 12060 12584 12124
rect 12601 12060 12665 12124
rect 12682 12060 12746 12124
rect 12763 12060 12827 12124
rect 12844 12060 12908 12124
rect 12925 12060 12989 12124
rect 13006 12060 13070 12124
rect 13087 12060 13151 12124
rect 13168 12060 13232 12124
rect 13249 12060 13313 12124
rect 13330 12060 13394 12124
rect 13411 12060 13475 12124
rect 13492 12060 13556 12124
rect 13573 12060 13637 12124
rect 13654 12060 13718 12124
rect 13735 12060 13799 12124
rect 13816 12060 13880 12124
rect 13897 12060 13961 12124
rect 13978 12060 14042 12124
rect 14059 12060 14123 12124
rect 14140 12060 14204 12124
rect 14221 12060 14285 12124
rect 14302 12060 14366 12124
rect 14383 12060 14447 12124
rect 14464 12060 14528 12124
rect 14545 12060 14609 12124
rect 14626 12060 14690 12124
rect 14707 12060 15000 12124
rect 14746 12042 15000 12060
rect 269 11978 333 12042
rect 351 11978 415 12042
rect 433 11978 497 12042
rect 515 11978 579 12042
rect 597 11978 661 12042
rect 678 11978 742 12042
rect 759 11978 823 12042
rect 840 11978 904 12042
rect 921 11978 985 12042
rect 1002 11978 1066 12042
rect 1083 11978 1147 12042
rect 1164 11978 1228 12042
rect 1245 11978 1309 12042
rect 1326 11978 1390 12042
rect 1407 11978 1471 12042
rect 1488 11978 1552 12042
rect 1569 11978 1633 12042
rect 1650 11978 1714 12042
rect 1731 11978 1795 12042
rect 1812 11978 1876 12042
rect 1893 11978 1957 12042
rect 1974 11978 2038 12042
rect 2055 11978 2119 12042
rect 2136 11978 2200 12042
rect 2217 11978 2281 12042
rect 2298 11978 2362 12042
rect 2379 11978 2443 12042
rect 2460 11978 2524 12042
rect 2541 11978 2605 12042
rect 2622 11978 2686 12042
rect 2703 11978 2767 12042
rect 2784 11978 2848 12042
rect 2865 11978 2929 12042
rect 2946 11978 3010 12042
rect 3027 11978 3091 12042
rect 3108 11978 3172 12042
rect 3189 11978 3253 12042
rect 3270 11978 3334 12042
rect 3351 11978 3415 12042
rect 3432 11978 3496 12042
rect 3513 11978 3577 12042
rect 3594 11978 3658 12042
rect 3675 11978 3739 12042
rect 3756 11978 3820 12042
rect 3837 11978 3901 12042
rect 3918 11978 3982 12042
rect 3999 11978 4063 12042
rect 4080 11978 4144 12042
rect 4161 11978 4225 12042
rect 4242 11978 4306 12042
rect 4323 11978 4387 12042
rect 4404 11978 4468 12042
rect 4485 11978 4549 12042
rect 4566 11978 4630 12042
rect 4647 11978 4711 12042
rect 4728 11978 4792 12042
rect 4809 11978 4873 12042
rect 10084 11978 10148 12042
rect 10166 11978 10230 12042
rect 10248 11978 10312 12042
rect 10330 11978 10394 12042
rect 10412 11978 10476 12042
rect 10494 11978 10558 12042
rect 10576 11978 10640 12042
rect 10657 11978 10721 12042
rect 10738 11978 10802 12042
rect 10819 11978 10883 12042
rect 10900 11978 10964 12042
rect 10981 11978 11045 12042
rect 11062 11978 11126 12042
rect 11143 11978 11207 12042
rect 11224 11978 11288 12042
rect 11305 11978 11369 12042
rect 11386 11978 11450 12042
rect 11467 11978 11531 12042
rect 11548 11978 11612 12042
rect 11629 11978 11693 12042
rect 11710 11978 11774 12042
rect 11791 11978 11855 12042
rect 11872 11978 11936 12042
rect 11953 11978 12017 12042
rect 12034 11978 12098 12042
rect 12115 11978 12179 12042
rect 12196 11978 12260 12042
rect 12277 11978 12341 12042
rect 12358 11978 12422 12042
rect 12439 11978 12503 12042
rect 12520 11978 12584 12042
rect 12601 11978 12665 12042
rect 12682 11978 12746 12042
rect 12763 11978 12827 12042
rect 12844 11978 12908 12042
rect 12925 11978 12989 12042
rect 13006 11978 13070 12042
rect 13087 11978 13151 12042
rect 13168 11978 13232 12042
rect 13249 11978 13313 12042
rect 13330 11978 13394 12042
rect 13411 11978 13475 12042
rect 13492 11978 13556 12042
rect 13573 11978 13637 12042
rect 13654 11978 13718 12042
rect 13735 11978 13799 12042
rect 13816 11978 13880 12042
rect 13897 11978 13961 12042
rect 13978 11978 14042 12042
rect 14059 11978 14123 12042
rect 14140 11978 14204 12042
rect 14221 11978 14285 12042
rect 14302 11978 14366 12042
rect 14383 11978 14447 12042
rect 14464 11978 14528 12042
rect 14545 11978 14609 12042
rect 14626 11978 14690 12042
rect 14707 11978 15000 12042
rect 14746 11960 15000 11978
rect 269 11896 333 11960
rect 351 11896 415 11960
rect 433 11896 497 11960
rect 515 11896 579 11960
rect 597 11896 661 11960
rect 678 11896 742 11960
rect 759 11896 823 11960
rect 840 11896 904 11960
rect 921 11896 985 11960
rect 1002 11896 1066 11960
rect 1083 11896 1147 11960
rect 1164 11896 1228 11960
rect 1245 11896 1309 11960
rect 1326 11896 1390 11960
rect 1407 11896 1471 11960
rect 1488 11896 1552 11960
rect 1569 11896 1633 11960
rect 1650 11896 1714 11960
rect 1731 11896 1795 11960
rect 1812 11896 1876 11960
rect 1893 11896 1957 11960
rect 1974 11896 2038 11960
rect 2055 11896 2119 11960
rect 2136 11896 2200 11960
rect 2217 11896 2281 11960
rect 2298 11896 2362 11960
rect 2379 11896 2443 11960
rect 2460 11896 2524 11960
rect 2541 11896 2605 11960
rect 2622 11896 2686 11960
rect 2703 11896 2767 11960
rect 2784 11896 2848 11960
rect 2865 11896 2929 11960
rect 2946 11896 3010 11960
rect 3027 11896 3091 11960
rect 3108 11896 3172 11960
rect 3189 11896 3253 11960
rect 3270 11896 3334 11960
rect 3351 11896 3415 11960
rect 3432 11896 3496 11960
rect 3513 11896 3577 11960
rect 3594 11896 3658 11960
rect 3675 11896 3739 11960
rect 3756 11896 3820 11960
rect 3837 11896 3901 11960
rect 3918 11896 3982 11960
rect 3999 11896 4063 11960
rect 4080 11896 4144 11960
rect 4161 11896 4225 11960
rect 4242 11896 4306 11960
rect 4323 11896 4387 11960
rect 4404 11896 4468 11960
rect 4485 11896 4549 11960
rect 4566 11896 4630 11960
rect 4647 11896 4711 11960
rect 4728 11896 4792 11960
rect 4809 11896 4873 11960
rect 10084 11896 10148 11960
rect 10166 11896 10230 11960
rect 10248 11896 10312 11960
rect 10330 11896 10394 11960
rect 10412 11896 10476 11960
rect 10494 11896 10558 11960
rect 10576 11896 10640 11960
rect 10657 11896 10721 11960
rect 10738 11896 10802 11960
rect 10819 11896 10883 11960
rect 10900 11896 10964 11960
rect 10981 11896 11045 11960
rect 11062 11896 11126 11960
rect 11143 11896 11207 11960
rect 11224 11896 11288 11960
rect 11305 11896 11369 11960
rect 11386 11896 11450 11960
rect 11467 11896 11531 11960
rect 11548 11896 11612 11960
rect 11629 11896 11693 11960
rect 11710 11896 11774 11960
rect 11791 11896 11855 11960
rect 11872 11896 11936 11960
rect 11953 11896 12017 11960
rect 12034 11896 12098 11960
rect 12115 11896 12179 11960
rect 12196 11896 12260 11960
rect 12277 11896 12341 11960
rect 12358 11896 12422 11960
rect 12439 11896 12503 11960
rect 12520 11896 12584 11960
rect 12601 11896 12665 11960
rect 12682 11896 12746 11960
rect 12763 11896 12827 11960
rect 12844 11896 12908 11960
rect 12925 11896 12989 11960
rect 13006 11896 13070 11960
rect 13087 11896 13151 11960
rect 13168 11896 13232 11960
rect 13249 11896 13313 11960
rect 13330 11896 13394 11960
rect 13411 11896 13475 11960
rect 13492 11896 13556 11960
rect 13573 11896 13637 11960
rect 13654 11896 13718 11960
rect 13735 11896 13799 11960
rect 13816 11896 13880 11960
rect 13897 11896 13961 11960
rect 13978 11896 14042 11960
rect 14059 11896 14123 11960
rect 14140 11896 14204 11960
rect 14221 11896 14285 11960
rect 14302 11896 14366 11960
rect 14383 11896 14447 11960
rect 14464 11896 14528 11960
rect 14545 11896 14609 11960
rect 14626 11896 14690 11960
rect 14707 11896 15000 11960
rect 14746 11878 15000 11896
rect 269 11814 333 11878
rect 351 11814 415 11878
rect 433 11814 497 11878
rect 515 11814 579 11878
rect 597 11814 661 11878
rect 678 11814 742 11878
rect 759 11814 823 11878
rect 840 11814 904 11878
rect 921 11814 985 11878
rect 1002 11814 1066 11878
rect 1083 11814 1147 11878
rect 1164 11814 1228 11878
rect 1245 11814 1309 11878
rect 1326 11814 1390 11878
rect 1407 11814 1471 11878
rect 1488 11814 1552 11878
rect 1569 11814 1633 11878
rect 1650 11814 1714 11878
rect 1731 11814 1795 11878
rect 1812 11814 1876 11878
rect 1893 11814 1957 11878
rect 1974 11814 2038 11878
rect 2055 11814 2119 11878
rect 2136 11814 2200 11878
rect 2217 11814 2281 11878
rect 2298 11814 2362 11878
rect 2379 11814 2443 11878
rect 2460 11814 2524 11878
rect 2541 11814 2605 11878
rect 2622 11814 2686 11878
rect 2703 11814 2767 11878
rect 2784 11814 2848 11878
rect 2865 11814 2929 11878
rect 2946 11814 3010 11878
rect 3027 11814 3091 11878
rect 3108 11814 3172 11878
rect 3189 11814 3253 11878
rect 3270 11814 3334 11878
rect 3351 11814 3415 11878
rect 3432 11814 3496 11878
rect 3513 11814 3577 11878
rect 3594 11814 3658 11878
rect 3675 11814 3739 11878
rect 3756 11814 3820 11878
rect 3837 11814 3901 11878
rect 3918 11814 3982 11878
rect 3999 11814 4063 11878
rect 4080 11814 4144 11878
rect 4161 11814 4225 11878
rect 4242 11814 4306 11878
rect 4323 11814 4387 11878
rect 4404 11814 4468 11878
rect 4485 11814 4549 11878
rect 4566 11814 4630 11878
rect 4647 11814 4711 11878
rect 4728 11814 4792 11878
rect 4809 11814 4873 11878
rect 10084 11814 10148 11878
rect 10166 11814 10230 11878
rect 10248 11814 10312 11878
rect 10330 11814 10394 11878
rect 10412 11814 10476 11878
rect 10494 11814 10558 11878
rect 10576 11814 10640 11878
rect 10657 11814 10721 11878
rect 10738 11814 10802 11878
rect 10819 11814 10883 11878
rect 10900 11814 10964 11878
rect 10981 11814 11045 11878
rect 11062 11814 11126 11878
rect 11143 11814 11207 11878
rect 11224 11814 11288 11878
rect 11305 11814 11369 11878
rect 11386 11814 11450 11878
rect 11467 11814 11531 11878
rect 11548 11814 11612 11878
rect 11629 11814 11693 11878
rect 11710 11814 11774 11878
rect 11791 11814 11855 11878
rect 11872 11814 11936 11878
rect 11953 11814 12017 11878
rect 12034 11814 12098 11878
rect 12115 11814 12179 11878
rect 12196 11814 12260 11878
rect 12277 11814 12341 11878
rect 12358 11814 12422 11878
rect 12439 11814 12503 11878
rect 12520 11814 12584 11878
rect 12601 11814 12665 11878
rect 12682 11814 12746 11878
rect 12763 11814 12827 11878
rect 12844 11814 12908 11878
rect 12925 11814 12989 11878
rect 13006 11814 13070 11878
rect 13087 11814 13151 11878
rect 13168 11814 13232 11878
rect 13249 11814 13313 11878
rect 13330 11814 13394 11878
rect 13411 11814 13475 11878
rect 13492 11814 13556 11878
rect 13573 11814 13637 11878
rect 13654 11814 13718 11878
rect 13735 11814 13799 11878
rect 13816 11814 13880 11878
rect 13897 11814 13961 11878
rect 13978 11814 14042 11878
rect 14059 11814 14123 11878
rect 14140 11814 14204 11878
rect 14221 11814 14285 11878
rect 14302 11814 14366 11878
rect 14383 11814 14447 11878
rect 14464 11814 14528 11878
rect 14545 11814 14609 11878
rect 14626 11814 14690 11878
rect 14707 11814 15000 11878
rect 14746 11796 15000 11814
rect 269 11732 333 11796
rect 351 11732 415 11796
rect 433 11732 497 11796
rect 515 11732 579 11796
rect 597 11732 661 11796
rect 678 11732 742 11796
rect 759 11732 823 11796
rect 840 11732 904 11796
rect 921 11732 985 11796
rect 1002 11732 1066 11796
rect 1083 11732 1147 11796
rect 1164 11732 1228 11796
rect 1245 11732 1309 11796
rect 1326 11732 1390 11796
rect 1407 11732 1471 11796
rect 1488 11732 1552 11796
rect 1569 11732 1633 11796
rect 1650 11732 1714 11796
rect 1731 11732 1795 11796
rect 1812 11732 1876 11796
rect 1893 11732 1957 11796
rect 1974 11732 2038 11796
rect 2055 11732 2119 11796
rect 2136 11732 2200 11796
rect 2217 11732 2281 11796
rect 2298 11732 2362 11796
rect 2379 11732 2443 11796
rect 2460 11732 2524 11796
rect 2541 11732 2605 11796
rect 2622 11732 2686 11796
rect 2703 11732 2767 11796
rect 2784 11732 2848 11796
rect 2865 11732 2929 11796
rect 2946 11732 3010 11796
rect 3027 11732 3091 11796
rect 3108 11732 3172 11796
rect 3189 11732 3253 11796
rect 3270 11732 3334 11796
rect 3351 11732 3415 11796
rect 3432 11732 3496 11796
rect 3513 11732 3577 11796
rect 3594 11732 3658 11796
rect 3675 11732 3739 11796
rect 3756 11732 3820 11796
rect 3837 11732 3901 11796
rect 3918 11732 3982 11796
rect 3999 11732 4063 11796
rect 4080 11732 4144 11796
rect 4161 11732 4225 11796
rect 4242 11732 4306 11796
rect 4323 11732 4387 11796
rect 4404 11732 4468 11796
rect 4485 11732 4549 11796
rect 4566 11732 4630 11796
rect 4647 11732 4711 11796
rect 4728 11732 4792 11796
rect 4809 11732 4873 11796
rect 10084 11732 10148 11796
rect 10166 11732 10230 11796
rect 10248 11732 10312 11796
rect 10330 11732 10394 11796
rect 10412 11732 10476 11796
rect 10494 11732 10558 11796
rect 10576 11732 10640 11796
rect 10657 11732 10721 11796
rect 10738 11732 10802 11796
rect 10819 11732 10883 11796
rect 10900 11732 10964 11796
rect 10981 11732 11045 11796
rect 11062 11732 11126 11796
rect 11143 11732 11207 11796
rect 11224 11732 11288 11796
rect 11305 11732 11369 11796
rect 11386 11732 11450 11796
rect 11467 11732 11531 11796
rect 11548 11732 11612 11796
rect 11629 11732 11693 11796
rect 11710 11732 11774 11796
rect 11791 11732 11855 11796
rect 11872 11732 11936 11796
rect 11953 11732 12017 11796
rect 12034 11732 12098 11796
rect 12115 11732 12179 11796
rect 12196 11732 12260 11796
rect 12277 11732 12341 11796
rect 12358 11732 12422 11796
rect 12439 11732 12503 11796
rect 12520 11732 12584 11796
rect 12601 11732 12665 11796
rect 12682 11732 12746 11796
rect 12763 11732 12827 11796
rect 12844 11732 12908 11796
rect 12925 11732 12989 11796
rect 13006 11732 13070 11796
rect 13087 11732 13151 11796
rect 13168 11732 13232 11796
rect 13249 11732 13313 11796
rect 13330 11732 13394 11796
rect 13411 11732 13475 11796
rect 13492 11732 13556 11796
rect 13573 11732 13637 11796
rect 13654 11732 13718 11796
rect 13735 11732 13799 11796
rect 13816 11732 13880 11796
rect 13897 11732 13961 11796
rect 13978 11732 14042 11796
rect 14059 11732 14123 11796
rect 14140 11732 14204 11796
rect 14221 11732 14285 11796
rect 14302 11732 14366 11796
rect 14383 11732 14447 11796
rect 14464 11732 14528 11796
rect 14545 11732 14609 11796
rect 14626 11732 14690 11796
rect 14707 11732 15000 11796
rect 14746 11714 15000 11732
rect 269 11650 333 11714
rect 351 11650 415 11714
rect 433 11650 497 11714
rect 515 11650 579 11714
rect 597 11650 661 11714
rect 678 11650 742 11714
rect 759 11650 823 11714
rect 840 11650 904 11714
rect 921 11650 985 11714
rect 1002 11650 1066 11714
rect 1083 11650 1147 11714
rect 1164 11650 1228 11714
rect 1245 11650 1309 11714
rect 1326 11650 1390 11714
rect 1407 11650 1471 11714
rect 1488 11650 1552 11714
rect 1569 11650 1633 11714
rect 1650 11650 1714 11714
rect 1731 11650 1795 11714
rect 1812 11650 1876 11714
rect 1893 11650 1957 11714
rect 1974 11650 2038 11714
rect 2055 11650 2119 11714
rect 2136 11650 2200 11714
rect 2217 11650 2281 11714
rect 2298 11650 2362 11714
rect 2379 11650 2443 11714
rect 2460 11650 2524 11714
rect 2541 11650 2605 11714
rect 2622 11650 2686 11714
rect 2703 11650 2767 11714
rect 2784 11650 2848 11714
rect 2865 11650 2929 11714
rect 2946 11650 3010 11714
rect 3027 11650 3091 11714
rect 3108 11650 3172 11714
rect 3189 11650 3253 11714
rect 3270 11650 3334 11714
rect 3351 11650 3415 11714
rect 3432 11650 3496 11714
rect 3513 11650 3577 11714
rect 3594 11650 3658 11714
rect 3675 11650 3739 11714
rect 3756 11650 3820 11714
rect 3837 11650 3901 11714
rect 3918 11650 3982 11714
rect 3999 11650 4063 11714
rect 4080 11650 4144 11714
rect 4161 11650 4225 11714
rect 4242 11650 4306 11714
rect 4323 11650 4387 11714
rect 4404 11650 4468 11714
rect 4485 11650 4549 11714
rect 4566 11650 4630 11714
rect 4647 11650 4711 11714
rect 4728 11650 4792 11714
rect 4809 11650 4873 11714
rect 10084 11650 10148 11714
rect 10166 11650 10230 11714
rect 10248 11650 10312 11714
rect 10330 11650 10394 11714
rect 10412 11650 10476 11714
rect 10494 11650 10558 11714
rect 10576 11650 10640 11714
rect 10657 11650 10721 11714
rect 10738 11650 10802 11714
rect 10819 11650 10883 11714
rect 10900 11650 10964 11714
rect 10981 11650 11045 11714
rect 11062 11650 11126 11714
rect 11143 11650 11207 11714
rect 11224 11650 11288 11714
rect 11305 11650 11369 11714
rect 11386 11650 11450 11714
rect 11467 11650 11531 11714
rect 11548 11650 11612 11714
rect 11629 11650 11693 11714
rect 11710 11650 11774 11714
rect 11791 11650 11855 11714
rect 11872 11650 11936 11714
rect 11953 11650 12017 11714
rect 12034 11650 12098 11714
rect 12115 11650 12179 11714
rect 12196 11650 12260 11714
rect 12277 11650 12341 11714
rect 12358 11650 12422 11714
rect 12439 11650 12503 11714
rect 12520 11650 12584 11714
rect 12601 11650 12665 11714
rect 12682 11650 12746 11714
rect 12763 11650 12827 11714
rect 12844 11650 12908 11714
rect 12925 11650 12989 11714
rect 13006 11650 13070 11714
rect 13087 11650 13151 11714
rect 13168 11650 13232 11714
rect 13249 11650 13313 11714
rect 13330 11650 13394 11714
rect 13411 11650 13475 11714
rect 13492 11650 13556 11714
rect 13573 11650 13637 11714
rect 13654 11650 13718 11714
rect 13735 11650 13799 11714
rect 13816 11650 13880 11714
rect 13897 11650 13961 11714
rect 13978 11650 14042 11714
rect 14059 11650 14123 11714
rect 14140 11650 14204 11714
rect 14221 11650 14285 11714
rect 14302 11650 14366 11714
rect 14383 11650 14447 11714
rect 14464 11650 14528 11714
rect 14545 11650 14609 11714
rect 14626 11650 14690 11714
rect 14707 11650 15000 11714
rect 14746 11647 15000 11650
rect 0 11281 15000 11347
rect 0 10625 15000 11221
rect 0 10329 254 10565
rect 14746 10329 15000 10565
rect 0 9673 15000 10269
rect 0 9547 15000 9613
rect 0 8317 254 9247
rect 14746 8317 15000 9247
rect 0 7347 254 8037
rect 14746 7347 15000 8037
rect 0 6377 254 7067
rect 14746 6377 15000 7067
rect 0 6053 254 6097
rect 14746 6053 15000 6097
rect 0 5817 379 6053
rect 465 5817 701 6053
rect 787 5817 1023 6053
rect 1109 5817 1345 6053
rect 1431 5817 1667 6053
rect 1753 5817 1989 6053
rect 2075 5817 2311 6053
rect 2397 5817 2633 6053
rect 2719 5817 2955 6053
rect 3041 5817 3277 6053
rect 3363 5817 3599 6053
rect 3685 5817 3921 6053
rect 4007 5817 4243 6053
rect 4329 5817 4565 6053
rect 4651 5817 4887 6053
rect 10111 5817 10347 6053
rect 10432 5817 10668 6053
rect 10753 5817 10989 6053
rect 11074 5817 11310 6053
rect 11395 5817 11631 6053
rect 11716 5817 11952 6053
rect 12037 5817 12273 6053
rect 12358 5817 12594 6053
rect 12679 5817 12915 6053
rect 13000 5817 13236 6053
rect 13321 5817 13557 6053
rect 13642 5817 13878 6053
rect 13963 5817 14199 6053
rect 14284 5817 14520 6053
rect 14605 5817 15000 6053
rect 0 5447 254 5817
rect 14746 5447 15000 5817
rect 0 5211 379 5447
rect 465 5211 701 5447
rect 787 5211 1023 5447
rect 1109 5211 1345 5447
rect 1431 5211 1667 5447
rect 1753 5211 1989 5447
rect 2075 5211 2311 5447
rect 2397 5211 2633 5447
rect 2719 5211 2955 5447
rect 3041 5211 3277 5447
rect 3363 5211 3599 5447
rect 3685 5211 3921 5447
rect 4007 5211 4243 5447
rect 4329 5211 4565 5447
rect 4651 5211 4887 5447
rect 10111 5211 10347 5447
rect 10432 5211 10668 5447
rect 10753 5211 10989 5447
rect 11074 5211 11310 5447
rect 11395 5211 11631 5447
rect 11716 5211 11952 5447
rect 12037 5211 12273 5447
rect 12358 5211 12594 5447
rect 12679 5211 12915 5447
rect 13000 5211 13236 5447
rect 13321 5211 13557 5447
rect 13642 5211 13878 5447
rect 13963 5211 14199 5447
rect 14284 5211 14520 5447
rect 14605 5211 15000 5447
rect 0 5167 254 5211
rect 14746 5167 15000 5211
rect 0 3957 254 4887
rect 14746 3957 15000 4887
rect 0 2987 193 3677
rect 14807 2987 15000 3677
rect 0 1777 254 2707
rect 14746 1777 15000 2707
rect 0 407 254 1497
rect 14746 407 15000 1497
<< obsm4 >>
rect 334 39983 2646 40000
rect 349 39919 365 39983
rect 429 39919 445 39983
rect 509 39919 525 39983
rect 589 39919 605 39983
rect 669 39919 685 39983
rect 749 39919 765 39983
rect 829 39919 845 39983
rect 909 39919 925 39983
rect 989 39919 1005 39983
rect 1069 39919 1085 39983
rect 1149 39919 1165 39983
rect 1229 39919 1245 39983
rect 1309 39919 1325 39983
rect 1389 39919 1405 39983
rect 1469 39919 1485 39983
rect 1549 39919 1565 39983
rect 1629 39919 1645 39983
rect 1709 39919 1725 39983
rect 1789 39919 1805 39983
rect 1869 39919 1885 39983
rect 1949 39919 1965 39983
rect 2029 39919 2045 39983
rect 2109 39919 2125 39983
rect 2189 39919 2205 39983
rect 2269 39919 2285 39983
rect 2349 39919 2365 39983
rect 2429 39919 2445 39983
rect 2509 39919 2525 39983
rect 2589 39919 2605 39983
rect 334 39902 2646 39919
rect 349 39838 365 39902
rect 429 39838 445 39902
rect 509 39838 525 39902
rect 589 39838 605 39902
rect 669 39838 685 39902
rect 749 39838 765 39902
rect 829 39838 845 39902
rect 909 39838 925 39902
rect 989 39838 1005 39902
rect 1069 39838 1085 39902
rect 1149 39838 1165 39902
rect 1229 39838 1245 39902
rect 1309 39838 1325 39902
rect 1389 39838 1405 39902
rect 1469 39838 1485 39902
rect 1549 39838 1565 39902
rect 1629 39838 1645 39902
rect 1709 39838 1725 39902
rect 1789 39838 1805 39902
rect 1869 39838 1885 39902
rect 1949 39838 1965 39902
rect 2029 39838 2045 39902
rect 2109 39838 2125 39902
rect 2189 39838 2205 39902
rect 2269 39838 2285 39902
rect 2349 39838 2365 39902
rect 2429 39838 2445 39902
rect 2509 39838 2525 39902
rect 2589 39838 2605 39902
rect 334 39821 2646 39838
rect 349 39757 365 39821
rect 429 39757 445 39821
rect 509 39757 525 39821
rect 589 39757 605 39821
rect 669 39757 685 39821
rect 749 39757 765 39821
rect 829 39757 845 39821
rect 909 39757 925 39821
rect 989 39757 1005 39821
rect 1069 39757 1085 39821
rect 1149 39757 1165 39821
rect 1229 39757 1245 39821
rect 1309 39757 1325 39821
rect 1389 39757 1405 39821
rect 1469 39757 1485 39821
rect 1549 39757 1565 39821
rect 1629 39757 1645 39821
rect 1709 39757 1725 39821
rect 1789 39757 1805 39821
rect 1869 39757 1885 39821
rect 1949 39757 1965 39821
rect 2029 39757 2045 39821
rect 2109 39757 2125 39821
rect 2189 39757 2205 39821
rect 2269 39757 2285 39821
rect 2349 39757 2365 39821
rect 2429 39757 2445 39821
rect 2509 39757 2525 39821
rect 2589 39757 2605 39821
rect 334 39740 2646 39757
rect 349 39676 365 39740
rect 429 39676 445 39740
rect 509 39676 525 39740
rect 589 39676 605 39740
rect 669 39676 685 39740
rect 749 39676 765 39740
rect 829 39676 845 39740
rect 909 39676 925 39740
rect 989 39676 1005 39740
rect 1069 39676 1085 39740
rect 1149 39676 1165 39740
rect 1229 39676 1245 39740
rect 1309 39676 1325 39740
rect 1389 39676 1405 39740
rect 1469 39676 1485 39740
rect 1549 39676 1565 39740
rect 1629 39676 1645 39740
rect 1709 39676 1725 39740
rect 1789 39676 1805 39740
rect 1869 39676 1885 39740
rect 1949 39676 1965 39740
rect 2029 39676 2045 39740
rect 2109 39676 2125 39740
rect 2189 39676 2205 39740
rect 2269 39676 2285 39740
rect 2349 39676 2365 39740
rect 2429 39676 2445 39740
rect 2509 39676 2525 39740
rect 2589 39676 2605 39740
rect 334 39659 2646 39676
rect 349 39595 365 39659
rect 429 39595 445 39659
rect 509 39595 525 39659
rect 589 39595 605 39659
rect 669 39595 685 39659
rect 749 39595 765 39659
rect 829 39595 845 39659
rect 909 39595 925 39659
rect 989 39595 1005 39659
rect 1069 39595 1085 39659
rect 1149 39595 1165 39659
rect 1229 39595 1245 39659
rect 1309 39595 1325 39659
rect 1389 39595 1405 39659
rect 1469 39595 1485 39659
rect 1549 39595 1565 39659
rect 1629 39595 1645 39659
rect 1709 39595 1725 39659
rect 1789 39595 1805 39659
rect 1869 39595 1885 39659
rect 1949 39595 1965 39659
rect 2029 39595 2045 39659
rect 2109 39595 2125 39659
rect 2189 39595 2205 39659
rect 2269 39595 2285 39659
rect 2349 39595 2365 39659
rect 2429 39595 2445 39659
rect 2509 39595 2525 39659
rect 2589 39595 2605 39659
rect 334 39578 2646 39595
rect 349 39514 365 39578
rect 429 39514 445 39578
rect 509 39514 525 39578
rect 589 39514 605 39578
rect 669 39514 685 39578
rect 749 39514 765 39578
rect 829 39514 845 39578
rect 909 39514 925 39578
rect 989 39514 1005 39578
rect 1069 39514 1085 39578
rect 1149 39514 1165 39578
rect 1229 39514 1245 39578
rect 1309 39514 1325 39578
rect 1389 39514 1405 39578
rect 1469 39514 1485 39578
rect 1549 39514 1565 39578
rect 1629 39514 1645 39578
rect 1709 39514 1725 39578
rect 1789 39514 1805 39578
rect 1869 39514 1885 39578
rect 1949 39514 1965 39578
rect 2029 39514 2045 39578
rect 2109 39514 2125 39578
rect 2189 39514 2205 39578
rect 2269 39514 2285 39578
rect 2349 39514 2365 39578
rect 2429 39514 2445 39578
rect 2509 39514 2525 39578
rect 2589 39514 2605 39578
rect 334 39497 2646 39514
rect 349 39433 365 39497
rect 429 39433 445 39497
rect 509 39433 525 39497
rect 589 39433 605 39497
rect 669 39433 685 39497
rect 749 39433 765 39497
rect 829 39433 845 39497
rect 909 39433 925 39497
rect 989 39433 1005 39497
rect 1069 39433 1085 39497
rect 1149 39433 1165 39497
rect 1229 39433 1245 39497
rect 1309 39433 1325 39497
rect 1389 39433 1405 39497
rect 1469 39433 1485 39497
rect 1549 39433 1565 39497
rect 1629 39433 1645 39497
rect 1709 39433 1725 39497
rect 1789 39433 1805 39497
rect 1869 39433 1885 39497
rect 1949 39433 1965 39497
rect 2029 39433 2045 39497
rect 2109 39433 2125 39497
rect 2189 39433 2205 39497
rect 2269 39433 2285 39497
rect 2349 39433 2365 39497
rect 2429 39433 2445 39497
rect 2509 39433 2525 39497
rect 2589 39433 2605 39497
rect 12345 39983 14666 40000
rect 12370 39919 12386 39983
rect 12450 39919 12466 39983
rect 12530 39919 12546 39983
rect 12610 39919 12626 39983
rect 12690 39919 12706 39983
rect 12770 39919 12786 39983
rect 12850 39919 12866 39983
rect 12930 39919 12946 39983
rect 13010 39919 13026 39983
rect 13090 39919 13106 39983
rect 13170 39919 13186 39983
rect 13250 39919 13266 39983
rect 13330 39919 13346 39983
rect 13410 39919 13426 39983
rect 13490 39919 13506 39983
rect 13570 39919 13586 39983
rect 13650 39919 13666 39983
rect 13730 39919 13746 39983
rect 13810 39919 13826 39983
rect 13890 39919 13906 39983
rect 13970 39919 13986 39983
rect 14050 39919 14066 39983
rect 14130 39919 14146 39983
rect 14210 39919 14226 39983
rect 14290 39919 14306 39983
rect 14370 39919 14386 39983
rect 14450 39919 14466 39983
rect 14530 39919 14546 39983
rect 14610 39919 14626 39983
rect 12345 39902 14666 39919
rect 12370 39838 12386 39902
rect 12450 39838 12466 39902
rect 12530 39838 12546 39902
rect 12610 39838 12626 39902
rect 12690 39838 12706 39902
rect 12770 39838 12786 39902
rect 12850 39838 12866 39902
rect 12930 39838 12946 39902
rect 13010 39838 13026 39902
rect 13090 39838 13106 39902
rect 13170 39838 13186 39902
rect 13250 39838 13266 39902
rect 13330 39838 13346 39902
rect 13410 39838 13426 39902
rect 13490 39838 13506 39902
rect 13570 39838 13586 39902
rect 13650 39838 13666 39902
rect 13730 39838 13746 39902
rect 13810 39838 13826 39902
rect 13890 39838 13906 39902
rect 13970 39838 13986 39902
rect 14050 39838 14066 39902
rect 14130 39838 14146 39902
rect 14210 39838 14226 39902
rect 14290 39838 14306 39902
rect 14370 39838 14386 39902
rect 14450 39838 14466 39902
rect 14530 39838 14546 39902
rect 14610 39838 14626 39902
rect 12345 39821 14666 39838
rect 12370 39757 12386 39821
rect 12450 39757 12466 39821
rect 12530 39757 12546 39821
rect 12610 39757 12626 39821
rect 12690 39757 12706 39821
rect 12770 39757 12786 39821
rect 12850 39757 12866 39821
rect 12930 39757 12946 39821
rect 13010 39757 13026 39821
rect 13090 39757 13106 39821
rect 13170 39757 13186 39821
rect 13250 39757 13266 39821
rect 13330 39757 13346 39821
rect 13410 39757 13426 39821
rect 13490 39757 13506 39821
rect 13570 39757 13586 39821
rect 13650 39757 13666 39821
rect 13730 39757 13746 39821
rect 13810 39757 13826 39821
rect 13890 39757 13906 39821
rect 13970 39757 13986 39821
rect 14050 39757 14066 39821
rect 14130 39757 14146 39821
rect 14210 39757 14226 39821
rect 14290 39757 14306 39821
rect 14370 39757 14386 39821
rect 14450 39757 14466 39821
rect 14530 39757 14546 39821
rect 14610 39757 14626 39821
rect 12345 39740 14666 39757
rect 12370 39676 12386 39740
rect 12450 39676 12466 39740
rect 12530 39676 12546 39740
rect 12610 39676 12626 39740
rect 12690 39676 12706 39740
rect 12770 39676 12786 39740
rect 12850 39676 12866 39740
rect 12930 39676 12946 39740
rect 13010 39676 13026 39740
rect 13090 39676 13106 39740
rect 13170 39676 13186 39740
rect 13250 39676 13266 39740
rect 13330 39676 13346 39740
rect 13410 39676 13426 39740
rect 13490 39676 13506 39740
rect 13570 39676 13586 39740
rect 13650 39676 13666 39740
rect 13730 39676 13746 39740
rect 13810 39676 13826 39740
rect 13890 39676 13906 39740
rect 13970 39676 13986 39740
rect 14050 39676 14066 39740
rect 14130 39676 14146 39740
rect 14210 39676 14226 39740
rect 14290 39676 14306 39740
rect 14370 39676 14386 39740
rect 14450 39676 14466 39740
rect 14530 39676 14546 39740
rect 14610 39676 14626 39740
rect 12345 39659 14666 39676
rect 12370 39595 12386 39659
rect 12450 39595 12466 39659
rect 12530 39595 12546 39659
rect 12610 39595 12626 39659
rect 12690 39595 12706 39659
rect 12770 39595 12786 39659
rect 12850 39595 12866 39659
rect 12930 39595 12946 39659
rect 13010 39595 13026 39659
rect 13090 39595 13106 39659
rect 13170 39595 13186 39659
rect 13250 39595 13266 39659
rect 13330 39595 13346 39659
rect 13410 39595 13426 39659
rect 13490 39595 13506 39659
rect 13570 39595 13586 39659
rect 13650 39595 13666 39659
rect 13730 39595 13746 39659
rect 13810 39595 13826 39659
rect 13890 39595 13906 39659
rect 13970 39595 13986 39659
rect 14050 39595 14066 39659
rect 14130 39595 14146 39659
rect 14210 39595 14226 39659
rect 14290 39595 14306 39659
rect 14370 39595 14386 39659
rect 14450 39595 14466 39659
rect 14530 39595 14546 39659
rect 14610 39595 14626 39659
rect 12345 39578 14666 39595
rect 12370 39514 12386 39578
rect 12450 39514 12466 39578
rect 12530 39514 12546 39578
rect 12610 39514 12626 39578
rect 12690 39514 12706 39578
rect 12770 39514 12786 39578
rect 12850 39514 12866 39578
rect 12930 39514 12946 39578
rect 13010 39514 13026 39578
rect 13090 39514 13106 39578
rect 13170 39514 13186 39578
rect 13250 39514 13266 39578
rect 13330 39514 13346 39578
rect 13410 39514 13426 39578
rect 13490 39514 13506 39578
rect 13570 39514 13586 39578
rect 13650 39514 13666 39578
rect 13730 39514 13746 39578
rect 13810 39514 13826 39578
rect 13890 39514 13906 39578
rect 13970 39514 13986 39578
rect 14050 39514 14066 39578
rect 14130 39514 14146 39578
rect 14210 39514 14226 39578
rect 14290 39514 14306 39578
rect 14370 39514 14386 39578
rect 14450 39514 14466 39578
rect 14530 39514 14546 39578
rect 14610 39514 14626 39578
rect 12345 39497 14666 39514
rect 12370 39433 12386 39497
rect 12450 39433 12466 39497
rect 12530 39433 12546 39497
rect 12610 39433 12626 39497
rect 12690 39433 12706 39497
rect 12770 39433 12786 39497
rect 12850 39433 12866 39497
rect 12930 39433 12946 39497
rect 13010 39433 13026 39497
rect 13090 39433 13106 39497
rect 13170 39433 13186 39497
rect 13250 39433 13266 39497
rect 13330 39433 13346 39497
rect 13410 39433 13426 39497
rect 13490 39433 13506 39497
rect 13570 39433 13586 39497
rect 13650 39433 13666 39497
rect 13730 39433 13746 39497
rect 13810 39433 13826 39497
rect 13890 39433 13906 39497
rect 13970 39433 13986 39497
rect 14050 39433 14066 39497
rect 14130 39433 14146 39497
rect 14210 39433 14226 39497
rect 14290 39433 14306 39497
rect 14370 39433 14386 39497
rect 14450 39433 14466 39497
rect 14530 39433 14546 39497
rect 14610 39433 14626 39497
rect 334 39416 2639 39433
rect 12348 39416 14666 39433
rect 349 39352 365 39416
rect 429 39352 445 39416
rect 509 39352 525 39416
rect 589 39352 605 39416
rect 669 39352 685 39416
rect 749 39352 765 39416
rect 829 39352 845 39416
rect 909 39352 925 39416
rect 989 39352 1005 39416
rect 1069 39352 1085 39416
rect 1149 39352 1165 39416
rect 1229 39352 1245 39416
rect 1309 39352 1325 39416
rect 1389 39352 1405 39416
rect 1469 39352 1485 39416
rect 1549 39352 1565 39416
rect 1629 39352 1645 39416
rect 1709 39352 1725 39416
rect 1789 39352 1805 39416
rect 1869 39352 1885 39416
rect 1949 39352 1965 39416
rect 2029 39352 2045 39416
rect 2109 39352 2125 39416
rect 2189 39352 2205 39416
rect 2269 39352 2285 39416
rect 2349 39352 2365 39416
rect 2429 39352 2445 39416
rect 2509 39352 2525 39416
rect 2589 39352 2605 39416
rect 334 39335 2639 39352
rect 349 39271 365 39335
rect 429 39271 445 39335
rect 509 39271 525 39335
rect 589 39271 605 39335
rect 669 39271 685 39335
rect 749 39271 765 39335
rect 829 39271 845 39335
rect 909 39271 925 39335
rect 989 39271 1005 39335
rect 1069 39271 1085 39335
rect 1149 39271 1165 39335
rect 1229 39271 1245 39335
rect 1309 39271 1325 39335
rect 1389 39271 1405 39335
rect 1469 39271 1485 39335
rect 1549 39271 1565 39335
rect 1629 39271 1645 39335
rect 1709 39271 1725 39335
rect 1789 39271 1805 39335
rect 1869 39271 1885 39335
rect 1949 39271 1965 39335
rect 2029 39271 2045 39335
rect 2109 39271 2125 39335
rect 2189 39271 2205 39335
rect 2269 39271 2285 39335
rect 2349 39271 2365 39335
rect 2429 39271 2445 39335
rect 2509 39271 2525 39335
rect 2589 39271 2605 39335
rect 334 39254 2639 39271
rect 349 39190 365 39254
rect 429 39190 445 39254
rect 509 39190 525 39254
rect 589 39190 605 39254
rect 669 39190 685 39254
rect 749 39190 765 39254
rect 829 39190 845 39254
rect 909 39190 925 39254
rect 989 39190 1005 39254
rect 1069 39190 1085 39254
rect 1149 39190 1165 39254
rect 1229 39190 1245 39254
rect 1309 39190 1325 39254
rect 1389 39190 1405 39254
rect 1469 39190 1485 39254
rect 1549 39190 1565 39254
rect 1629 39190 1645 39254
rect 1709 39190 1725 39254
rect 1789 39190 1805 39254
rect 1869 39190 1885 39254
rect 1949 39190 1965 39254
rect 2029 39190 2045 39254
rect 2109 39190 2125 39254
rect 2189 39190 2205 39254
rect 2269 39190 2285 39254
rect 2349 39190 2365 39254
rect 2429 39190 2445 39254
rect 2509 39190 2525 39254
rect 2589 39190 2605 39254
rect 334 39173 2639 39190
rect 349 39109 365 39173
rect 429 39109 445 39173
rect 509 39109 525 39173
rect 589 39109 605 39173
rect 669 39109 685 39173
rect 749 39109 765 39173
rect 829 39109 845 39173
rect 909 39109 925 39173
rect 989 39109 1005 39173
rect 1069 39109 1085 39173
rect 1149 39109 1165 39173
rect 1229 39109 1245 39173
rect 1309 39109 1325 39173
rect 1389 39109 1405 39173
rect 1469 39109 1485 39173
rect 1549 39109 1565 39173
rect 1629 39109 1645 39173
rect 1709 39109 1725 39173
rect 1789 39109 1805 39173
rect 1869 39109 1885 39173
rect 1949 39109 1965 39173
rect 2029 39109 2045 39173
rect 2109 39109 2125 39173
rect 2189 39109 2205 39173
rect 2269 39109 2285 39173
rect 2349 39109 2365 39173
rect 2429 39109 2445 39173
rect 2509 39109 2525 39173
rect 2589 39109 2605 39173
rect 2931 39166 12056 39354
rect 12370 39352 12386 39416
rect 12450 39352 12466 39416
rect 12530 39352 12546 39416
rect 12610 39352 12626 39416
rect 12690 39352 12706 39416
rect 12770 39352 12786 39416
rect 12850 39352 12866 39416
rect 12930 39352 12946 39416
rect 13010 39352 13026 39416
rect 13090 39352 13106 39416
rect 13170 39352 13186 39416
rect 13250 39352 13266 39416
rect 13330 39352 13346 39416
rect 13410 39352 13426 39416
rect 13490 39352 13506 39416
rect 13570 39352 13586 39416
rect 13650 39352 13666 39416
rect 13730 39352 13746 39416
rect 13810 39352 13826 39416
rect 13890 39352 13906 39416
rect 13970 39352 13986 39416
rect 14050 39352 14066 39416
rect 14130 39352 14146 39416
rect 14210 39352 14226 39416
rect 14290 39352 14306 39416
rect 14370 39352 14386 39416
rect 14450 39352 14466 39416
rect 14530 39352 14546 39416
rect 14610 39352 14626 39416
rect 12348 39335 14666 39352
rect 12370 39271 12386 39335
rect 12450 39271 12466 39335
rect 12530 39271 12546 39335
rect 12610 39271 12626 39335
rect 12690 39271 12706 39335
rect 12770 39271 12786 39335
rect 12850 39271 12866 39335
rect 12930 39271 12946 39335
rect 13010 39271 13026 39335
rect 13090 39271 13106 39335
rect 13170 39271 13186 39335
rect 13250 39271 13266 39335
rect 13330 39271 13346 39335
rect 13410 39271 13426 39335
rect 13490 39271 13506 39335
rect 13570 39271 13586 39335
rect 13650 39271 13666 39335
rect 13730 39271 13746 39335
rect 13810 39271 13826 39335
rect 13890 39271 13906 39335
rect 13970 39271 13986 39335
rect 14050 39271 14066 39335
rect 14130 39271 14146 39335
rect 14210 39271 14226 39335
rect 14290 39271 14306 39335
rect 14370 39271 14386 39335
rect 14450 39271 14466 39335
rect 14530 39271 14546 39335
rect 14610 39271 14626 39335
rect 12348 39254 14666 39271
rect 12370 39190 12386 39254
rect 12450 39190 12466 39254
rect 12530 39190 12546 39254
rect 12610 39190 12626 39254
rect 12690 39190 12706 39254
rect 12770 39190 12786 39254
rect 12850 39190 12866 39254
rect 12930 39190 12946 39254
rect 13010 39190 13026 39254
rect 13090 39190 13106 39254
rect 13170 39190 13186 39254
rect 13250 39190 13266 39254
rect 13330 39190 13346 39254
rect 13410 39190 13426 39254
rect 13490 39190 13506 39254
rect 13570 39190 13586 39254
rect 13650 39190 13666 39254
rect 13730 39190 13746 39254
rect 13810 39190 13826 39254
rect 13890 39190 13906 39254
rect 13970 39190 13986 39254
rect 14050 39190 14066 39254
rect 14130 39190 14146 39254
rect 14210 39190 14226 39254
rect 14290 39190 14306 39254
rect 14370 39190 14386 39254
rect 14450 39190 14466 39254
rect 14530 39190 14546 39254
rect 14610 39190 14626 39254
rect 12348 39173 14666 39190
rect 2669 39109 12306 39166
rect 12370 39109 12386 39173
rect 12450 39109 12466 39173
rect 12530 39109 12546 39173
rect 12610 39109 12626 39173
rect 12690 39109 12706 39173
rect 12770 39109 12786 39173
rect 12850 39109 12866 39173
rect 12930 39109 12946 39173
rect 13010 39109 13026 39173
rect 13090 39109 13106 39173
rect 13170 39109 13186 39173
rect 13250 39109 13266 39173
rect 13330 39109 13346 39173
rect 13410 39109 13426 39173
rect 13490 39109 13506 39173
rect 13570 39109 13586 39173
rect 13650 39109 13666 39173
rect 13730 39109 13746 39173
rect 13810 39109 13826 39173
rect 13890 39109 13906 39173
rect 13970 39109 13986 39173
rect 14050 39109 14066 39173
rect 14130 39109 14146 39173
rect 14210 39109 14226 39173
rect 14290 39109 14306 39173
rect 14370 39109 14386 39173
rect 14450 39109 14466 39173
rect 14530 39109 14546 39173
rect 14610 39109 14626 39173
rect 334 39092 14666 39109
rect 349 39028 365 39092
rect 429 39028 445 39092
rect 509 39028 525 39092
rect 589 39028 605 39092
rect 669 39028 685 39092
rect 749 39028 765 39092
rect 829 39028 845 39092
rect 909 39028 925 39092
rect 989 39028 1005 39092
rect 1069 39028 1085 39092
rect 1149 39028 1165 39092
rect 1229 39028 1245 39092
rect 1309 39028 1325 39092
rect 1389 39028 1405 39092
rect 1469 39028 1485 39092
rect 1549 39028 1565 39092
rect 1629 39028 1645 39092
rect 1709 39028 1725 39092
rect 1789 39028 1805 39092
rect 1869 39028 1885 39092
rect 1949 39028 1965 39092
rect 2029 39028 2045 39092
rect 2109 39028 2125 39092
rect 2189 39028 2205 39092
rect 2269 39028 2285 39092
rect 2349 39028 2365 39092
rect 2429 39028 2445 39092
rect 2509 39028 2525 39092
rect 2589 39028 2605 39092
rect 2669 39028 12306 39092
rect 12370 39028 12386 39092
rect 12450 39028 12466 39092
rect 12530 39028 12546 39092
rect 12610 39028 12626 39092
rect 12690 39028 12706 39092
rect 12770 39028 12786 39092
rect 12850 39028 12866 39092
rect 12930 39028 12946 39092
rect 13010 39028 13026 39092
rect 13090 39028 13106 39092
rect 13170 39028 13186 39092
rect 13250 39028 13266 39092
rect 13330 39028 13346 39092
rect 13410 39028 13426 39092
rect 13490 39028 13506 39092
rect 13570 39028 13586 39092
rect 13650 39028 13666 39092
rect 13730 39028 13746 39092
rect 13810 39028 13826 39092
rect 13890 39028 13906 39092
rect 13970 39028 13986 39092
rect 14050 39028 14066 39092
rect 14130 39028 14146 39092
rect 14210 39028 14226 39092
rect 14290 39028 14306 39092
rect 14370 39028 14386 39092
rect 14450 39028 14466 39092
rect 14530 39028 14546 39092
rect 14610 39028 14626 39092
rect 334 39011 14666 39028
rect 2669 35187 12306 39011
rect 334 35077 14666 35187
rect 193 19080 14807 35077
rect 334 13927 14666 19080
rect 193 13787 14807 13927
rect 334 12737 14666 13787
rect 193 12617 14807 12737
rect 334 12534 14666 12617
rect 334 12470 351 12534
rect 415 12470 433 12534
rect 497 12470 515 12534
rect 579 12470 597 12534
rect 661 12470 678 12534
rect 742 12470 759 12534
rect 823 12470 840 12534
rect 904 12470 921 12534
rect 985 12470 1002 12534
rect 1066 12470 1083 12534
rect 1147 12470 1164 12534
rect 1228 12470 1245 12534
rect 1309 12470 1326 12534
rect 1390 12470 1407 12534
rect 1471 12470 1488 12534
rect 1552 12470 1569 12534
rect 1633 12470 1650 12534
rect 1714 12470 1731 12534
rect 1795 12470 1812 12534
rect 1876 12470 1893 12534
rect 1957 12470 1974 12534
rect 2038 12470 2055 12534
rect 2119 12470 2136 12534
rect 2200 12470 2217 12534
rect 2281 12470 2298 12534
rect 2362 12470 2379 12534
rect 2443 12470 2460 12534
rect 2524 12470 2541 12534
rect 2605 12470 2622 12534
rect 2686 12470 2703 12534
rect 2767 12470 2784 12534
rect 2848 12470 2865 12534
rect 2929 12470 2946 12534
rect 3010 12470 3027 12534
rect 3091 12470 3108 12534
rect 3172 12470 3189 12534
rect 3253 12470 3270 12534
rect 3334 12470 3351 12534
rect 3415 12470 3432 12534
rect 3496 12470 3513 12534
rect 3577 12470 3594 12534
rect 3658 12470 3675 12534
rect 3739 12470 3756 12534
rect 3820 12470 3837 12534
rect 3901 12470 3918 12534
rect 3982 12470 3999 12534
rect 4063 12470 4080 12534
rect 4144 12470 4161 12534
rect 4225 12470 4242 12534
rect 4306 12470 4323 12534
rect 4387 12470 4404 12534
rect 4468 12470 4485 12534
rect 4549 12470 4566 12534
rect 4630 12470 4647 12534
rect 4711 12470 4728 12534
rect 4792 12470 4809 12534
rect 4873 12470 10084 12534
rect 10148 12470 10166 12534
rect 10230 12470 10248 12534
rect 10312 12470 10330 12534
rect 10394 12470 10412 12534
rect 10476 12470 10494 12534
rect 10558 12470 10576 12534
rect 10640 12470 10657 12534
rect 10721 12470 10738 12534
rect 10802 12470 10819 12534
rect 10883 12470 10900 12534
rect 10964 12470 10981 12534
rect 11045 12470 11062 12534
rect 11126 12470 11143 12534
rect 11207 12470 11224 12534
rect 11288 12470 11305 12534
rect 11369 12470 11386 12534
rect 11450 12470 11467 12534
rect 11531 12470 11548 12534
rect 11612 12470 11629 12534
rect 11693 12470 11710 12534
rect 11774 12470 11791 12534
rect 11855 12470 11872 12534
rect 11936 12470 11953 12534
rect 12017 12470 12034 12534
rect 12098 12470 12115 12534
rect 12179 12470 12196 12534
rect 12260 12470 12277 12534
rect 12341 12470 12358 12534
rect 12422 12470 12439 12534
rect 12503 12470 12520 12534
rect 12584 12470 12601 12534
rect 12665 12470 12682 12534
rect 12746 12470 12763 12534
rect 12827 12470 12844 12534
rect 12908 12470 12925 12534
rect 12989 12470 13006 12534
rect 13070 12470 13087 12534
rect 13151 12470 13168 12534
rect 13232 12470 13249 12534
rect 13313 12470 13330 12534
rect 13394 12470 13411 12534
rect 13475 12470 13492 12534
rect 13556 12470 13573 12534
rect 13637 12470 13654 12534
rect 13718 12470 13735 12534
rect 13799 12470 13816 12534
rect 13880 12470 13897 12534
rect 13961 12470 13978 12534
rect 14042 12470 14059 12534
rect 14123 12470 14140 12534
rect 14204 12470 14221 12534
rect 14285 12470 14302 12534
rect 14366 12470 14383 12534
rect 14447 12470 14464 12534
rect 14528 12470 14545 12534
rect 14609 12470 14626 12534
rect 334 12452 14666 12470
rect 334 12388 351 12452
rect 415 12388 433 12452
rect 497 12388 515 12452
rect 579 12388 597 12452
rect 661 12388 678 12452
rect 742 12388 759 12452
rect 823 12388 840 12452
rect 904 12388 921 12452
rect 985 12388 1002 12452
rect 1066 12388 1083 12452
rect 1147 12388 1164 12452
rect 1228 12388 1245 12452
rect 1309 12388 1326 12452
rect 1390 12388 1407 12452
rect 1471 12388 1488 12452
rect 1552 12388 1569 12452
rect 1633 12388 1650 12452
rect 1714 12388 1731 12452
rect 1795 12388 1812 12452
rect 1876 12388 1893 12452
rect 1957 12388 1974 12452
rect 2038 12388 2055 12452
rect 2119 12388 2136 12452
rect 2200 12388 2217 12452
rect 2281 12388 2298 12452
rect 2362 12388 2379 12452
rect 2443 12388 2460 12452
rect 2524 12388 2541 12452
rect 2605 12388 2622 12452
rect 2686 12388 2703 12452
rect 2767 12388 2784 12452
rect 2848 12388 2865 12452
rect 2929 12388 2946 12452
rect 3010 12388 3027 12452
rect 3091 12388 3108 12452
rect 3172 12388 3189 12452
rect 3253 12388 3270 12452
rect 3334 12388 3351 12452
rect 3415 12388 3432 12452
rect 3496 12388 3513 12452
rect 3577 12388 3594 12452
rect 3658 12388 3675 12452
rect 3739 12388 3756 12452
rect 3820 12388 3837 12452
rect 3901 12388 3918 12452
rect 3982 12388 3999 12452
rect 4063 12388 4080 12452
rect 4144 12388 4161 12452
rect 4225 12388 4242 12452
rect 4306 12388 4323 12452
rect 4387 12388 4404 12452
rect 4468 12388 4485 12452
rect 4549 12388 4566 12452
rect 4630 12388 4647 12452
rect 4711 12388 4728 12452
rect 4792 12388 4809 12452
rect 4873 12388 10084 12452
rect 10148 12388 10166 12452
rect 10230 12388 10248 12452
rect 10312 12388 10330 12452
rect 10394 12388 10412 12452
rect 10476 12388 10494 12452
rect 10558 12388 10576 12452
rect 10640 12388 10657 12452
rect 10721 12388 10738 12452
rect 10802 12388 10819 12452
rect 10883 12388 10900 12452
rect 10964 12388 10981 12452
rect 11045 12388 11062 12452
rect 11126 12388 11143 12452
rect 11207 12388 11224 12452
rect 11288 12388 11305 12452
rect 11369 12388 11386 12452
rect 11450 12388 11467 12452
rect 11531 12388 11548 12452
rect 11612 12388 11629 12452
rect 11693 12388 11710 12452
rect 11774 12388 11791 12452
rect 11855 12388 11872 12452
rect 11936 12388 11953 12452
rect 12017 12388 12034 12452
rect 12098 12388 12115 12452
rect 12179 12388 12196 12452
rect 12260 12388 12277 12452
rect 12341 12388 12358 12452
rect 12422 12388 12439 12452
rect 12503 12388 12520 12452
rect 12584 12388 12601 12452
rect 12665 12388 12682 12452
rect 12746 12388 12763 12452
rect 12827 12388 12844 12452
rect 12908 12388 12925 12452
rect 12989 12388 13006 12452
rect 13070 12388 13087 12452
rect 13151 12388 13168 12452
rect 13232 12388 13249 12452
rect 13313 12388 13330 12452
rect 13394 12388 13411 12452
rect 13475 12388 13492 12452
rect 13556 12388 13573 12452
rect 13637 12388 13654 12452
rect 13718 12388 13735 12452
rect 13799 12388 13816 12452
rect 13880 12388 13897 12452
rect 13961 12388 13978 12452
rect 14042 12388 14059 12452
rect 14123 12388 14140 12452
rect 14204 12388 14221 12452
rect 14285 12388 14302 12452
rect 14366 12388 14383 12452
rect 14447 12388 14464 12452
rect 14528 12388 14545 12452
rect 14609 12388 14626 12452
rect 334 12370 14666 12388
rect 334 12306 351 12370
rect 415 12306 433 12370
rect 497 12306 515 12370
rect 579 12306 597 12370
rect 661 12306 678 12370
rect 742 12306 759 12370
rect 823 12306 840 12370
rect 904 12306 921 12370
rect 985 12306 1002 12370
rect 1066 12306 1083 12370
rect 1147 12306 1164 12370
rect 1228 12306 1245 12370
rect 1309 12306 1326 12370
rect 1390 12306 1407 12370
rect 1471 12306 1488 12370
rect 1552 12306 1569 12370
rect 1633 12306 1650 12370
rect 1714 12306 1731 12370
rect 1795 12306 1812 12370
rect 1876 12306 1893 12370
rect 1957 12306 1974 12370
rect 2038 12306 2055 12370
rect 2119 12306 2136 12370
rect 2200 12306 2217 12370
rect 2281 12306 2298 12370
rect 2362 12306 2379 12370
rect 2443 12306 2460 12370
rect 2524 12306 2541 12370
rect 2605 12306 2622 12370
rect 2686 12306 2703 12370
rect 2767 12306 2784 12370
rect 2848 12306 2865 12370
rect 2929 12306 2946 12370
rect 3010 12306 3027 12370
rect 3091 12306 3108 12370
rect 3172 12306 3189 12370
rect 3253 12306 3270 12370
rect 3334 12306 3351 12370
rect 3415 12306 3432 12370
rect 3496 12306 3513 12370
rect 3577 12306 3594 12370
rect 3658 12306 3675 12370
rect 3739 12306 3756 12370
rect 3820 12306 3837 12370
rect 3901 12306 3918 12370
rect 3982 12306 3999 12370
rect 4063 12306 4080 12370
rect 4144 12306 4161 12370
rect 4225 12306 4242 12370
rect 4306 12306 4323 12370
rect 4387 12306 4404 12370
rect 4468 12306 4485 12370
rect 4549 12306 4566 12370
rect 4630 12306 4647 12370
rect 4711 12306 4728 12370
rect 4792 12306 4809 12370
rect 4873 12306 10084 12370
rect 10148 12306 10166 12370
rect 10230 12306 10248 12370
rect 10312 12306 10330 12370
rect 10394 12306 10412 12370
rect 10476 12306 10494 12370
rect 10558 12306 10576 12370
rect 10640 12306 10657 12370
rect 10721 12306 10738 12370
rect 10802 12306 10819 12370
rect 10883 12306 10900 12370
rect 10964 12306 10981 12370
rect 11045 12306 11062 12370
rect 11126 12306 11143 12370
rect 11207 12306 11224 12370
rect 11288 12306 11305 12370
rect 11369 12306 11386 12370
rect 11450 12306 11467 12370
rect 11531 12306 11548 12370
rect 11612 12306 11629 12370
rect 11693 12306 11710 12370
rect 11774 12306 11791 12370
rect 11855 12306 11872 12370
rect 11936 12306 11953 12370
rect 12017 12306 12034 12370
rect 12098 12306 12115 12370
rect 12179 12306 12196 12370
rect 12260 12306 12277 12370
rect 12341 12306 12358 12370
rect 12422 12306 12439 12370
rect 12503 12306 12520 12370
rect 12584 12306 12601 12370
rect 12665 12306 12682 12370
rect 12746 12306 12763 12370
rect 12827 12306 12844 12370
rect 12908 12306 12925 12370
rect 12989 12306 13006 12370
rect 13070 12306 13087 12370
rect 13151 12306 13168 12370
rect 13232 12306 13249 12370
rect 13313 12306 13330 12370
rect 13394 12306 13411 12370
rect 13475 12306 13492 12370
rect 13556 12306 13573 12370
rect 13637 12306 13654 12370
rect 13718 12306 13735 12370
rect 13799 12306 13816 12370
rect 13880 12306 13897 12370
rect 13961 12306 13978 12370
rect 14042 12306 14059 12370
rect 14123 12306 14140 12370
rect 14204 12306 14221 12370
rect 14285 12306 14302 12370
rect 14366 12306 14383 12370
rect 14447 12306 14464 12370
rect 14528 12306 14545 12370
rect 14609 12306 14626 12370
rect 334 12288 14666 12306
rect 334 12224 351 12288
rect 415 12224 433 12288
rect 497 12224 515 12288
rect 579 12224 597 12288
rect 661 12224 678 12288
rect 742 12224 759 12288
rect 823 12224 840 12288
rect 904 12224 921 12288
rect 985 12224 1002 12288
rect 1066 12224 1083 12288
rect 1147 12224 1164 12288
rect 1228 12224 1245 12288
rect 1309 12224 1326 12288
rect 1390 12224 1407 12288
rect 1471 12224 1488 12288
rect 1552 12224 1569 12288
rect 1633 12224 1650 12288
rect 1714 12224 1731 12288
rect 1795 12224 1812 12288
rect 1876 12224 1893 12288
rect 1957 12224 1974 12288
rect 2038 12224 2055 12288
rect 2119 12224 2136 12288
rect 2200 12224 2217 12288
rect 2281 12224 2298 12288
rect 2362 12224 2379 12288
rect 2443 12224 2460 12288
rect 2524 12224 2541 12288
rect 2605 12224 2622 12288
rect 2686 12224 2703 12288
rect 2767 12224 2784 12288
rect 2848 12224 2865 12288
rect 2929 12224 2946 12288
rect 3010 12224 3027 12288
rect 3091 12224 3108 12288
rect 3172 12224 3189 12288
rect 3253 12224 3270 12288
rect 3334 12224 3351 12288
rect 3415 12224 3432 12288
rect 3496 12224 3513 12288
rect 3577 12224 3594 12288
rect 3658 12224 3675 12288
rect 3739 12224 3756 12288
rect 3820 12224 3837 12288
rect 3901 12224 3918 12288
rect 3982 12224 3999 12288
rect 4063 12224 4080 12288
rect 4144 12224 4161 12288
rect 4225 12224 4242 12288
rect 4306 12224 4323 12288
rect 4387 12224 4404 12288
rect 4468 12224 4485 12288
rect 4549 12224 4566 12288
rect 4630 12224 4647 12288
rect 4711 12224 4728 12288
rect 4792 12224 4809 12288
rect 4873 12224 10084 12288
rect 10148 12224 10166 12288
rect 10230 12224 10248 12288
rect 10312 12224 10330 12288
rect 10394 12224 10412 12288
rect 10476 12224 10494 12288
rect 10558 12224 10576 12288
rect 10640 12224 10657 12288
rect 10721 12224 10738 12288
rect 10802 12224 10819 12288
rect 10883 12224 10900 12288
rect 10964 12224 10981 12288
rect 11045 12224 11062 12288
rect 11126 12224 11143 12288
rect 11207 12224 11224 12288
rect 11288 12224 11305 12288
rect 11369 12224 11386 12288
rect 11450 12224 11467 12288
rect 11531 12224 11548 12288
rect 11612 12224 11629 12288
rect 11693 12224 11710 12288
rect 11774 12224 11791 12288
rect 11855 12224 11872 12288
rect 11936 12224 11953 12288
rect 12017 12224 12034 12288
rect 12098 12224 12115 12288
rect 12179 12224 12196 12288
rect 12260 12224 12277 12288
rect 12341 12224 12358 12288
rect 12422 12224 12439 12288
rect 12503 12224 12520 12288
rect 12584 12224 12601 12288
rect 12665 12224 12682 12288
rect 12746 12224 12763 12288
rect 12827 12224 12844 12288
rect 12908 12224 12925 12288
rect 12989 12224 13006 12288
rect 13070 12224 13087 12288
rect 13151 12224 13168 12288
rect 13232 12224 13249 12288
rect 13313 12224 13330 12288
rect 13394 12224 13411 12288
rect 13475 12224 13492 12288
rect 13556 12224 13573 12288
rect 13637 12224 13654 12288
rect 13718 12224 13735 12288
rect 13799 12224 13816 12288
rect 13880 12224 13897 12288
rect 13961 12224 13978 12288
rect 14042 12224 14059 12288
rect 14123 12224 14140 12288
rect 14204 12224 14221 12288
rect 14285 12224 14302 12288
rect 14366 12224 14383 12288
rect 14447 12224 14464 12288
rect 14528 12224 14545 12288
rect 14609 12224 14626 12288
rect 334 12206 14666 12224
rect 334 12142 351 12206
rect 415 12142 433 12206
rect 497 12142 515 12206
rect 579 12142 597 12206
rect 661 12142 678 12206
rect 742 12142 759 12206
rect 823 12142 840 12206
rect 904 12142 921 12206
rect 985 12142 1002 12206
rect 1066 12142 1083 12206
rect 1147 12142 1164 12206
rect 1228 12142 1245 12206
rect 1309 12142 1326 12206
rect 1390 12142 1407 12206
rect 1471 12142 1488 12206
rect 1552 12142 1569 12206
rect 1633 12142 1650 12206
rect 1714 12142 1731 12206
rect 1795 12142 1812 12206
rect 1876 12142 1893 12206
rect 1957 12142 1974 12206
rect 2038 12142 2055 12206
rect 2119 12142 2136 12206
rect 2200 12142 2217 12206
rect 2281 12142 2298 12206
rect 2362 12142 2379 12206
rect 2443 12142 2460 12206
rect 2524 12142 2541 12206
rect 2605 12142 2622 12206
rect 2686 12142 2703 12206
rect 2767 12142 2784 12206
rect 2848 12142 2865 12206
rect 2929 12142 2946 12206
rect 3010 12142 3027 12206
rect 3091 12142 3108 12206
rect 3172 12142 3189 12206
rect 3253 12142 3270 12206
rect 3334 12142 3351 12206
rect 3415 12142 3432 12206
rect 3496 12142 3513 12206
rect 3577 12142 3594 12206
rect 3658 12142 3675 12206
rect 3739 12142 3756 12206
rect 3820 12142 3837 12206
rect 3901 12142 3918 12206
rect 3982 12142 3999 12206
rect 4063 12142 4080 12206
rect 4144 12142 4161 12206
rect 4225 12142 4242 12206
rect 4306 12142 4323 12206
rect 4387 12142 4404 12206
rect 4468 12142 4485 12206
rect 4549 12142 4566 12206
rect 4630 12142 4647 12206
rect 4711 12142 4728 12206
rect 4792 12142 4809 12206
rect 4873 12142 10084 12206
rect 10148 12142 10166 12206
rect 10230 12142 10248 12206
rect 10312 12142 10330 12206
rect 10394 12142 10412 12206
rect 10476 12142 10494 12206
rect 10558 12142 10576 12206
rect 10640 12142 10657 12206
rect 10721 12142 10738 12206
rect 10802 12142 10819 12206
rect 10883 12142 10900 12206
rect 10964 12142 10981 12206
rect 11045 12142 11062 12206
rect 11126 12142 11143 12206
rect 11207 12142 11224 12206
rect 11288 12142 11305 12206
rect 11369 12142 11386 12206
rect 11450 12142 11467 12206
rect 11531 12142 11548 12206
rect 11612 12142 11629 12206
rect 11693 12142 11710 12206
rect 11774 12142 11791 12206
rect 11855 12142 11872 12206
rect 11936 12142 11953 12206
rect 12017 12142 12034 12206
rect 12098 12142 12115 12206
rect 12179 12142 12196 12206
rect 12260 12142 12277 12206
rect 12341 12142 12358 12206
rect 12422 12142 12439 12206
rect 12503 12142 12520 12206
rect 12584 12142 12601 12206
rect 12665 12142 12682 12206
rect 12746 12142 12763 12206
rect 12827 12142 12844 12206
rect 12908 12142 12925 12206
rect 12989 12142 13006 12206
rect 13070 12142 13087 12206
rect 13151 12142 13168 12206
rect 13232 12142 13249 12206
rect 13313 12142 13330 12206
rect 13394 12142 13411 12206
rect 13475 12142 13492 12206
rect 13556 12142 13573 12206
rect 13637 12142 13654 12206
rect 13718 12142 13735 12206
rect 13799 12142 13816 12206
rect 13880 12142 13897 12206
rect 13961 12142 13978 12206
rect 14042 12142 14059 12206
rect 14123 12142 14140 12206
rect 14204 12142 14221 12206
rect 14285 12142 14302 12206
rect 14366 12142 14383 12206
rect 14447 12142 14464 12206
rect 14528 12142 14545 12206
rect 14609 12142 14626 12206
rect 334 12124 14666 12142
rect 334 12060 351 12124
rect 415 12060 433 12124
rect 497 12060 515 12124
rect 579 12060 597 12124
rect 661 12060 678 12124
rect 742 12060 759 12124
rect 823 12060 840 12124
rect 904 12060 921 12124
rect 985 12060 1002 12124
rect 1066 12060 1083 12124
rect 1147 12060 1164 12124
rect 1228 12060 1245 12124
rect 1309 12060 1326 12124
rect 1390 12060 1407 12124
rect 1471 12060 1488 12124
rect 1552 12060 1569 12124
rect 1633 12060 1650 12124
rect 1714 12060 1731 12124
rect 1795 12060 1812 12124
rect 1876 12060 1893 12124
rect 1957 12060 1974 12124
rect 2038 12060 2055 12124
rect 2119 12060 2136 12124
rect 2200 12060 2217 12124
rect 2281 12060 2298 12124
rect 2362 12060 2379 12124
rect 2443 12060 2460 12124
rect 2524 12060 2541 12124
rect 2605 12060 2622 12124
rect 2686 12060 2703 12124
rect 2767 12060 2784 12124
rect 2848 12060 2865 12124
rect 2929 12060 2946 12124
rect 3010 12060 3027 12124
rect 3091 12060 3108 12124
rect 3172 12060 3189 12124
rect 3253 12060 3270 12124
rect 3334 12060 3351 12124
rect 3415 12060 3432 12124
rect 3496 12060 3513 12124
rect 3577 12060 3594 12124
rect 3658 12060 3675 12124
rect 3739 12060 3756 12124
rect 3820 12060 3837 12124
rect 3901 12060 3918 12124
rect 3982 12060 3999 12124
rect 4063 12060 4080 12124
rect 4144 12060 4161 12124
rect 4225 12060 4242 12124
rect 4306 12060 4323 12124
rect 4387 12060 4404 12124
rect 4468 12060 4485 12124
rect 4549 12060 4566 12124
rect 4630 12060 4647 12124
rect 4711 12060 4728 12124
rect 4792 12060 4809 12124
rect 4873 12060 10084 12124
rect 10148 12060 10166 12124
rect 10230 12060 10248 12124
rect 10312 12060 10330 12124
rect 10394 12060 10412 12124
rect 10476 12060 10494 12124
rect 10558 12060 10576 12124
rect 10640 12060 10657 12124
rect 10721 12060 10738 12124
rect 10802 12060 10819 12124
rect 10883 12060 10900 12124
rect 10964 12060 10981 12124
rect 11045 12060 11062 12124
rect 11126 12060 11143 12124
rect 11207 12060 11224 12124
rect 11288 12060 11305 12124
rect 11369 12060 11386 12124
rect 11450 12060 11467 12124
rect 11531 12060 11548 12124
rect 11612 12060 11629 12124
rect 11693 12060 11710 12124
rect 11774 12060 11791 12124
rect 11855 12060 11872 12124
rect 11936 12060 11953 12124
rect 12017 12060 12034 12124
rect 12098 12060 12115 12124
rect 12179 12060 12196 12124
rect 12260 12060 12277 12124
rect 12341 12060 12358 12124
rect 12422 12060 12439 12124
rect 12503 12060 12520 12124
rect 12584 12060 12601 12124
rect 12665 12060 12682 12124
rect 12746 12060 12763 12124
rect 12827 12060 12844 12124
rect 12908 12060 12925 12124
rect 12989 12060 13006 12124
rect 13070 12060 13087 12124
rect 13151 12060 13168 12124
rect 13232 12060 13249 12124
rect 13313 12060 13330 12124
rect 13394 12060 13411 12124
rect 13475 12060 13492 12124
rect 13556 12060 13573 12124
rect 13637 12060 13654 12124
rect 13718 12060 13735 12124
rect 13799 12060 13816 12124
rect 13880 12060 13897 12124
rect 13961 12060 13978 12124
rect 14042 12060 14059 12124
rect 14123 12060 14140 12124
rect 14204 12060 14221 12124
rect 14285 12060 14302 12124
rect 14366 12060 14383 12124
rect 14447 12060 14464 12124
rect 14528 12060 14545 12124
rect 14609 12060 14626 12124
rect 334 12042 14666 12060
rect 334 11978 351 12042
rect 415 11978 433 12042
rect 497 11978 515 12042
rect 579 11978 597 12042
rect 661 11978 678 12042
rect 742 11978 759 12042
rect 823 11978 840 12042
rect 904 11978 921 12042
rect 985 11978 1002 12042
rect 1066 11978 1083 12042
rect 1147 11978 1164 12042
rect 1228 11978 1245 12042
rect 1309 11978 1326 12042
rect 1390 11978 1407 12042
rect 1471 11978 1488 12042
rect 1552 11978 1569 12042
rect 1633 11978 1650 12042
rect 1714 11978 1731 12042
rect 1795 11978 1812 12042
rect 1876 11978 1893 12042
rect 1957 11978 1974 12042
rect 2038 11978 2055 12042
rect 2119 11978 2136 12042
rect 2200 11978 2217 12042
rect 2281 11978 2298 12042
rect 2362 11978 2379 12042
rect 2443 11978 2460 12042
rect 2524 11978 2541 12042
rect 2605 11978 2622 12042
rect 2686 11978 2703 12042
rect 2767 11978 2784 12042
rect 2848 11978 2865 12042
rect 2929 11978 2946 12042
rect 3010 11978 3027 12042
rect 3091 11978 3108 12042
rect 3172 11978 3189 12042
rect 3253 11978 3270 12042
rect 3334 11978 3351 12042
rect 3415 11978 3432 12042
rect 3496 11978 3513 12042
rect 3577 11978 3594 12042
rect 3658 11978 3675 12042
rect 3739 11978 3756 12042
rect 3820 11978 3837 12042
rect 3901 11978 3918 12042
rect 3982 11978 3999 12042
rect 4063 11978 4080 12042
rect 4144 11978 4161 12042
rect 4225 11978 4242 12042
rect 4306 11978 4323 12042
rect 4387 11978 4404 12042
rect 4468 11978 4485 12042
rect 4549 11978 4566 12042
rect 4630 11978 4647 12042
rect 4711 11978 4728 12042
rect 4792 11978 4809 12042
rect 4873 11978 10084 12042
rect 10148 11978 10166 12042
rect 10230 11978 10248 12042
rect 10312 11978 10330 12042
rect 10394 11978 10412 12042
rect 10476 11978 10494 12042
rect 10558 11978 10576 12042
rect 10640 11978 10657 12042
rect 10721 11978 10738 12042
rect 10802 11978 10819 12042
rect 10883 11978 10900 12042
rect 10964 11978 10981 12042
rect 11045 11978 11062 12042
rect 11126 11978 11143 12042
rect 11207 11978 11224 12042
rect 11288 11978 11305 12042
rect 11369 11978 11386 12042
rect 11450 11978 11467 12042
rect 11531 11978 11548 12042
rect 11612 11978 11629 12042
rect 11693 11978 11710 12042
rect 11774 11978 11791 12042
rect 11855 11978 11872 12042
rect 11936 11978 11953 12042
rect 12017 11978 12034 12042
rect 12098 11978 12115 12042
rect 12179 11978 12196 12042
rect 12260 11978 12277 12042
rect 12341 11978 12358 12042
rect 12422 11978 12439 12042
rect 12503 11978 12520 12042
rect 12584 11978 12601 12042
rect 12665 11978 12682 12042
rect 12746 11978 12763 12042
rect 12827 11978 12844 12042
rect 12908 11978 12925 12042
rect 12989 11978 13006 12042
rect 13070 11978 13087 12042
rect 13151 11978 13168 12042
rect 13232 11978 13249 12042
rect 13313 11978 13330 12042
rect 13394 11978 13411 12042
rect 13475 11978 13492 12042
rect 13556 11978 13573 12042
rect 13637 11978 13654 12042
rect 13718 11978 13735 12042
rect 13799 11978 13816 12042
rect 13880 11978 13897 12042
rect 13961 11978 13978 12042
rect 14042 11978 14059 12042
rect 14123 11978 14140 12042
rect 14204 11978 14221 12042
rect 14285 11978 14302 12042
rect 14366 11978 14383 12042
rect 14447 11978 14464 12042
rect 14528 11978 14545 12042
rect 14609 11978 14626 12042
rect 334 11960 14666 11978
rect 334 11896 351 11960
rect 415 11896 433 11960
rect 497 11896 515 11960
rect 579 11896 597 11960
rect 661 11896 678 11960
rect 742 11896 759 11960
rect 823 11896 840 11960
rect 904 11896 921 11960
rect 985 11896 1002 11960
rect 1066 11896 1083 11960
rect 1147 11896 1164 11960
rect 1228 11896 1245 11960
rect 1309 11896 1326 11960
rect 1390 11896 1407 11960
rect 1471 11896 1488 11960
rect 1552 11896 1569 11960
rect 1633 11896 1650 11960
rect 1714 11896 1731 11960
rect 1795 11896 1812 11960
rect 1876 11896 1893 11960
rect 1957 11896 1974 11960
rect 2038 11896 2055 11960
rect 2119 11896 2136 11960
rect 2200 11896 2217 11960
rect 2281 11896 2298 11960
rect 2362 11896 2379 11960
rect 2443 11896 2460 11960
rect 2524 11896 2541 11960
rect 2605 11896 2622 11960
rect 2686 11896 2703 11960
rect 2767 11896 2784 11960
rect 2848 11896 2865 11960
rect 2929 11896 2946 11960
rect 3010 11896 3027 11960
rect 3091 11896 3108 11960
rect 3172 11896 3189 11960
rect 3253 11896 3270 11960
rect 3334 11896 3351 11960
rect 3415 11896 3432 11960
rect 3496 11896 3513 11960
rect 3577 11896 3594 11960
rect 3658 11896 3675 11960
rect 3739 11896 3756 11960
rect 3820 11896 3837 11960
rect 3901 11896 3918 11960
rect 3982 11896 3999 11960
rect 4063 11896 4080 11960
rect 4144 11896 4161 11960
rect 4225 11896 4242 11960
rect 4306 11896 4323 11960
rect 4387 11896 4404 11960
rect 4468 11896 4485 11960
rect 4549 11896 4566 11960
rect 4630 11896 4647 11960
rect 4711 11896 4728 11960
rect 4792 11896 4809 11960
rect 4873 11896 10084 11960
rect 10148 11896 10166 11960
rect 10230 11896 10248 11960
rect 10312 11896 10330 11960
rect 10394 11896 10412 11960
rect 10476 11896 10494 11960
rect 10558 11896 10576 11960
rect 10640 11896 10657 11960
rect 10721 11896 10738 11960
rect 10802 11896 10819 11960
rect 10883 11896 10900 11960
rect 10964 11896 10981 11960
rect 11045 11896 11062 11960
rect 11126 11896 11143 11960
rect 11207 11896 11224 11960
rect 11288 11896 11305 11960
rect 11369 11896 11386 11960
rect 11450 11896 11467 11960
rect 11531 11896 11548 11960
rect 11612 11896 11629 11960
rect 11693 11896 11710 11960
rect 11774 11896 11791 11960
rect 11855 11896 11872 11960
rect 11936 11896 11953 11960
rect 12017 11896 12034 11960
rect 12098 11896 12115 11960
rect 12179 11896 12196 11960
rect 12260 11896 12277 11960
rect 12341 11896 12358 11960
rect 12422 11896 12439 11960
rect 12503 11896 12520 11960
rect 12584 11896 12601 11960
rect 12665 11896 12682 11960
rect 12746 11896 12763 11960
rect 12827 11896 12844 11960
rect 12908 11896 12925 11960
rect 12989 11896 13006 11960
rect 13070 11896 13087 11960
rect 13151 11896 13168 11960
rect 13232 11896 13249 11960
rect 13313 11896 13330 11960
rect 13394 11896 13411 11960
rect 13475 11896 13492 11960
rect 13556 11896 13573 11960
rect 13637 11896 13654 11960
rect 13718 11896 13735 11960
rect 13799 11896 13816 11960
rect 13880 11896 13897 11960
rect 13961 11896 13978 11960
rect 14042 11896 14059 11960
rect 14123 11896 14140 11960
rect 14204 11896 14221 11960
rect 14285 11896 14302 11960
rect 14366 11896 14383 11960
rect 14447 11896 14464 11960
rect 14528 11896 14545 11960
rect 14609 11896 14626 11960
rect 334 11878 14666 11896
rect 334 11814 351 11878
rect 415 11814 433 11878
rect 497 11814 515 11878
rect 579 11814 597 11878
rect 661 11814 678 11878
rect 742 11814 759 11878
rect 823 11814 840 11878
rect 904 11814 921 11878
rect 985 11814 1002 11878
rect 1066 11814 1083 11878
rect 1147 11814 1164 11878
rect 1228 11814 1245 11878
rect 1309 11814 1326 11878
rect 1390 11814 1407 11878
rect 1471 11814 1488 11878
rect 1552 11814 1569 11878
rect 1633 11814 1650 11878
rect 1714 11814 1731 11878
rect 1795 11814 1812 11878
rect 1876 11814 1893 11878
rect 1957 11814 1974 11878
rect 2038 11814 2055 11878
rect 2119 11814 2136 11878
rect 2200 11814 2217 11878
rect 2281 11814 2298 11878
rect 2362 11814 2379 11878
rect 2443 11814 2460 11878
rect 2524 11814 2541 11878
rect 2605 11814 2622 11878
rect 2686 11814 2703 11878
rect 2767 11814 2784 11878
rect 2848 11814 2865 11878
rect 2929 11814 2946 11878
rect 3010 11814 3027 11878
rect 3091 11814 3108 11878
rect 3172 11814 3189 11878
rect 3253 11814 3270 11878
rect 3334 11814 3351 11878
rect 3415 11814 3432 11878
rect 3496 11814 3513 11878
rect 3577 11814 3594 11878
rect 3658 11814 3675 11878
rect 3739 11814 3756 11878
rect 3820 11814 3837 11878
rect 3901 11814 3918 11878
rect 3982 11814 3999 11878
rect 4063 11814 4080 11878
rect 4144 11814 4161 11878
rect 4225 11814 4242 11878
rect 4306 11814 4323 11878
rect 4387 11814 4404 11878
rect 4468 11814 4485 11878
rect 4549 11814 4566 11878
rect 4630 11814 4647 11878
rect 4711 11814 4728 11878
rect 4792 11814 4809 11878
rect 4873 11814 10084 11878
rect 10148 11814 10166 11878
rect 10230 11814 10248 11878
rect 10312 11814 10330 11878
rect 10394 11814 10412 11878
rect 10476 11814 10494 11878
rect 10558 11814 10576 11878
rect 10640 11814 10657 11878
rect 10721 11814 10738 11878
rect 10802 11814 10819 11878
rect 10883 11814 10900 11878
rect 10964 11814 10981 11878
rect 11045 11814 11062 11878
rect 11126 11814 11143 11878
rect 11207 11814 11224 11878
rect 11288 11814 11305 11878
rect 11369 11814 11386 11878
rect 11450 11814 11467 11878
rect 11531 11814 11548 11878
rect 11612 11814 11629 11878
rect 11693 11814 11710 11878
rect 11774 11814 11791 11878
rect 11855 11814 11872 11878
rect 11936 11814 11953 11878
rect 12017 11814 12034 11878
rect 12098 11814 12115 11878
rect 12179 11814 12196 11878
rect 12260 11814 12277 11878
rect 12341 11814 12358 11878
rect 12422 11814 12439 11878
rect 12503 11814 12520 11878
rect 12584 11814 12601 11878
rect 12665 11814 12682 11878
rect 12746 11814 12763 11878
rect 12827 11814 12844 11878
rect 12908 11814 12925 11878
rect 12989 11814 13006 11878
rect 13070 11814 13087 11878
rect 13151 11814 13168 11878
rect 13232 11814 13249 11878
rect 13313 11814 13330 11878
rect 13394 11814 13411 11878
rect 13475 11814 13492 11878
rect 13556 11814 13573 11878
rect 13637 11814 13654 11878
rect 13718 11814 13735 11878
rect 13799 11814 13816 11878
rect 13880 11814 13897 11878
rect 13961 11814 13978 11878
rect 14042 11814 14059 11878
rect 14123 11814 14140 11878
rect 14204 11814 14221 11878
rect 14285 11814 14302 11878
rect 14366 11814 14383 11878
rect 14447 11814 14464 11878
rect 14528 11814 14545 11878
rect 14609 11814 14626 11878
rect 334 11796 14666 11814
rect 334 11732 351 11796
rect 415 11732 433 11796
rect 497 11732 515 11796
rect 579 11732 597 11796
rect 661 11732 678 11796
rect 742 11732 759 11796
rect 823 11732 840 11796
rect 904 11732 921 11796
rect 985 11732 1002 11796
rect 1066 11732 1083 11796
rect 1147 11732 1164 11796
rect 1228 11732 1245 11796
rect 1309 11732 1326 11796
rect 1390 11732 1407 11796
rect 1471 11732 1488 11796
rect 1552 11732 1569 11796
rect 1633 11732 1650 11796
rect 1714 11732 1731 11796
rect 1795 11732 1812 11796
rect 1876 11732 1893 11796
rect 1957 11732 1974 11796
rect 2038 11732 2055 11796
rect 2119 11732 2136 11796
rect 2200 11732 2217 11796
rect 2281 11732 2298 11796
rect 2362 11732 2379 11796
rect 2443 11732 2460 11796
rect 2524 11732 2541 11796
rect 2605 11732 2622 11796
rect 2686 11732 2703 11796
rect 2767 11732 2784 11796
rect 2848 11732 2865 11796
rect 2929 11732 2946 11796
rect 3010 11732 3027 11796
rect 3091 11732 3108 11796
rect 3172 11732 3189 11796
rect 3253 11732 3270 11796
rect 3334 11732 3351 11796
rect 3415 11732 3432 11796
rect 3496 11732 3513 11796
rect 3577 11732 3594 11796
rect 3658 11732 3675 11796
rect 3739 11732 3756 11796
rect 3820 11732 3837 11796
rect 3901 11732 3918 11796
rect 3982 11732 3999 11796
rect 4063 11732 4080 11796
rect 4144 11732 4161 11796
rect 4225 11732 4242 11796
rect 4306 11732 4323 11796
rect 4387 11732 4404 11796
rect 4468 11732 4485 11796
rect 4549 11732 4566 11796
rect 4630 11732 4647 11796
rect 4711 11732 4728 11796
rect 4792 11732 4809 11796
rect 4873 11732 10084 11796
rect 10148 11732 10166 11796
rect 10230 11732 10248 11796
rect 10312 11732 10330 11796
rect 10394 11732 10412 11796
rect 10476 11732 10494 11796
rect 10558 11732 10576 11796
rect 10640 11732 10657 11796
rect 10721 11732 10738 11796
rect 10802 11732 10819 11796
rect 10883 11732 10900 11796
rect 10964 11732 10981 11796
rect 11045 11732 11062 11796
rect 11126 11732 11143 11796
rect 11207 11732 11224 11796
rect 11288 11732 11305 11796
rect 11369 11732 11386 11796
rect 11450 11732 11467 11796
rect 11531 11732 11548 11796
rect 11612 11732 11629 11796
rect 11693 11732 11710 11796
rect 11774 11732 11791 11796
rect 11855 11732 11872 11796
rect 11936 11732 11953 11796
rect 12017 11732 12034 11796
rect 12098 11732 12115 11796
rect 12179 11732 12196 11796
rect 12260 11732 12277 11796
rect 12341 11732 12358 11796
rect 12422 11732 12439 11796
rect 12503 11732 12520 11796
rect 12584 11732 12601 11796
rect 12665 11732 12682 11796
rect 12746 11732 12763 11796
rect 12827 11732 12844 11796
rect 12908 11732 12925 11796
rect 12989 11732 13006 11796
rect 13070 11732 13087 11796
rect 13151 11732 13168 11796
rect 13232 11732 13249 11796
rect 13313 11732 13330 11796
rect 13394 11732 13411 11796
rect 13475 11732 13492 11796
rect 13556 11732 13573 11796
rect 13637 11732 13654 11796
rect 13718 11732 13735 11796
rect 13799 11732 13816 11796
rect 13880 11732 13897 11796
rect 13961 11732 13978 11796
rect 14042 11732 14059 11796
rect 14123 11732 14140 11796
rect 14204 11732 14221 11796
rect 14285 11732 14302 11796
rect 14366 11732 14383 11796
rect 14447 11732 14464 11796
rect 14528 11732 14545 11796
rect 14609 11732 14626 11796
rect 334 11714 14666 11732
rect 334 11650 351 11714
rect 415 11650 433 11714
rect 497 11650 515 11714
rect 579 11650 597 11714
rect 661 11650 678 11714
rect 742 11650 759 11714
rect 823 11650 840 11714
rect 904 11650 921 11714
rect 985 11650 1002 11714
rect 1066 11650 1083 11714
rect 1147 11650 1164 11714
rect 1228 11650 1245 11714
rect 1309 11650 1326 11714
rect 1390 11650 1407 11714
rect 1471 11650 1488 11714
rect 1552 11650 1569 11714
rect 1633 11650 1650 11714
rect 1714 11650 1731 11714
rect 1795 11650 1812 11714
rect 1876 11650 1893 11714
rect 1957 11650 1974 11714
rect 2038 11650 2055 11714
rect 2119 11650 2136 11714
rect 2200 11650 2217 11714
rect 2281 11650 2298 11714
rect 2362 11650 2379 11714
rect 2443 11650 2460 11714
rect 2524 11650 2541 11714
rect 2605 11650 2622 11714
rect 2686 11650 2703 11714
rect 2767 11650 2784 11714
rect 2848 11650 2865 11714
rect 2929 11650 2946 11714
rect 3010 11650 3027 11714
rect 3091 11650 3108 11714
rect 3172 11650 3189 11714
rect 3253 11650 3270 11714
rect 3334 11650 3351 11714
rect 3415 11650 3432 11714
rect 3496 11650 3513 11714
rect 3577 11650 3594 11714
rect 3658 11650 3675 11714
rect 3739 11650 3756 11714
rect 3820 11650 3837 11714
rect 3901 11650 3918 11714
rect 3982 11650 3999 11714
rect 4063 11650 4080 11714
rect 4144 11650 4161 11714
rect 4225 11650 4242 11714
rect 4306 11650 4323 11714
rect 4387 11650 4404 11714
rect 4468 11650 4485 11714
rect 4549 11650 4566 11714
rect 4630 11650 4647 11714
rect 4711 11650 4728 11714
rect 4792 11650 4809 11714
rect 4873 11650 10084 11714
rect 10148 11650 10166 11714
rect 10230 11650 10248 11714
rect 10312 11650 10330 11714
rect 10394 11650 10412 11714
rect 10476 11650 10494 11714
rect 10558 11650 10576 11714
rect 10640 11650 10657 11714
rect 10721 11650 10738 11714
rect 10802 11650 10819 11714
rect 10883 11650 10900 11714
rect 10964 11650 10981 11714
rect 11045 11650 11062 11714
rect 11126 11650 11143 11714
rect 11207 11650 11224 11714
rect 11288 11650 11305 11714
rect 11369 11650 11386 11714
rect 11450 11650 11467 11714
rect 11531 11650 11548 11714
rect 11612 11650 11629 11714
rect 11693 11650 11710 11714
rect 11774 11650 11791 11714
rect 11855 11650 11872 11714
rect 11936 11650 11953 11714
rect 12017 11650 12034 11714
rect 12098 11650 12115 11714
rect 12179 11650 12196 11714
rect 12260 11650 12277 11714
rect 12341 11650 12358 11714
rect 12422 11650 12439 11714
rect 12503 11650 12520 11714
rect 12584 11650 12601 11714
rect 12665 11650 12682 11714
rect 12746 11650 12763 11714
rect 12827 11650 12844 11714
rect 12908 11650 12925 11714
rect 12989 11650 13006 11714
rect 13070 11650 13087 11714
rect 13151 11650 13168 11714
rect 13232 11650 13249 11714
rect 13313 11650 13330 11714
rect 13394 11650 13411 11714
rect 13475 11650 13492 11714
rect 13556 11650 13573 11714
rect 13637 11650 13654 11714
rect 13718 11650 13735 11714
rect 13799 11650 13816 11714
rect 13880 11650 13897 11714
rect 13961 11650 13978 11714
rect 14042 11650 14059 11714
rect 14123 11650 14140 11714
rect 14204 11650 14221 11714
rect 14285 11650 14302 11714
rect 14366 11650 14383 11714
rect 14447 11650 14464 11714
rect 14528 11650 14545 11714
rect 14609 11650 14626 11714
rect 334 11567 14666 11650
rect 193 11427 14807 11567
rect 334 10349 14666 10545
rect 193 9327 14807 9467
rect 334 8237 14666 9327
rect 193 8117 14807 8237
rect 334 7267 14666 8117
rect 193 7147 14807 7267
rect 334 6297 14666 7147
rect 193 6177 14807 6297
rect 334 6053 14666 6177
rect 379 5817 465 6053
rect 701 5817 787 6053
rect 1023 5817 1109 6053
rect 1345 5817 1431 6053
rect 1667 5817 1753 6053
rect 1989 5817 2075 6053
rect 2311 5817 2397 6053
rect 2633 5817 2719 6053
rect 2955 5817 3041 6053
rect 3277 5817 3363 6053
rect 3599 5817 3685 6053
rect 3921 5817 4007 6053
rect 4243 5817 4329 6053
rect 4565 5817 4651 6053
rect 4887 5817 10111 6053
rect 10347 5817 10432 6053
rect 10668 5817 10753 6053
rect 10989 5817 11074 6053
rect 11310 5817 11395 6053
rect 11631 5817 11716 6053
rect 11952 5817 12037 6053
rect 12273 5817 12358 6053
rect 12594 5817 12679 6053
rect 12915 5817 13000 6053
rect 13236 5817 13321 6053
rect 13557 5817 13642 6053
rect 13878 5817 13963 6053
rect 14199 5817 14284 6053
rect 14520 5817 14605 6053
rect 334 5447 14666 5817
rect 379 5211 465 5447
rect 701 5211 787 5447
rect 1023 5211 1109 5447
rect 1345 5211 1431 5447
rect 1667 5211 1753 5447
rect 1989 5211 2075 5447
rect 2311 5211 2397 5447
rect 2633 5211 2719 5447
rect 2955 5211 3041 5447
rect 3277 5211 3363 5447
rect 3599 5211 3685 5447
rect 3921 5211 4007 5447
rect 4243 5211 4329 5447
rect 4565 5211 4651 5447
rect 4887 5211 10111 5447
rect 10347 5211 10432 5447
rect 10668 5211 10753 5447
rect 10989 5211 11074 5447
rect 11310 5211 11395 5447
rect 11631 5211 11716 5447
rect 11952 5211 12037 5447
rect 12273 5211 12358 5447
rect 12594 5211 12679 5447
rect 12915 5211 13000 5447
rect 13236 5211 13321 5447
rect 13557 5211 13642 5447
rect 13878 5211 13963 5447
rect 14199 5211 14284 5447
rect 14520 5211 14605 5447
rect 334 5087 14666 5211
rect 193 4967 14807 5087
rect 334 3877 14666 4967
rect 193 3757 14807 3877
rect 273 2907 14727 3757
rect 193 2787 14807 2907
rect 334 1697 14666 2787
rect 193 1577 14807 1697
rect 334 407 14666 1577
<< metal5 >>
rect 0 35157 254 40000
rect 14746 35157 15000 40000
rect 0 14007 254 18997
rect 0 12837 254 13687
rect 0 11667 254 12517
rect 0 9547 254 11347
rect 0 8337 254 9227
rect 0 7368 254 8017
rect 14746 14007 15000 18997
rect 14746 12837 15000 13687
rect 14746 11667 15000 12517
rect 14746 9547 15000 11347
rect 14746 8337 15000 9227
rect 14746 7368 15000 8017
rect 0 6397 254 7047
rect 0 6053 254 6077
rect 14746 6397 15000 7047
rect 14746 6053 15000 6077
rect 0 5817 379 6053
rect 465 5817 701 6053
rect 787 5817 1023 6053
rect 1109 5817 1345 6053
rect 1431 5817 1667 6053
rect 1753 5817 1989 6053
rect 2075 5817 2311 6053
rect 2397 5817 2633 6053
rect 2719 5817 2955 6053
rect 3041 5817 3277 6053
rect 3363 5817 3599 6053
rect 3685 5817 3921 6053
rect 4007 5817 4243 6053
rect 4329 5817 4565 6053
rect 4651 5817 4887 6053
rect 10111 5817 10347 6053
rect 10432 5817 10668 6053
rect 10753 5817 10989 6053
rect 11074 5817 11310 6053
rect 11395 5817 11631 6053
rect 11716 5817 11952 6053
rect 12037 5817 12273 6053
rect 12358 5817 12594 6053
rect 12679 5817 12915 6053
rect 13000 5817 13236 6053
rect 13321 5817 13557 6053
rect 13642 5817 13878 6053
rect 13963 5817 14199 6053
rect 14284 5817 14520 6053
rect 14605 5817 15000 6053
rect 0 5447 254 5817
rect 14746 5447 15000 5817
rect 0 5211 379 5447
rect 465 5211 701 5447
rect 787 5211 1023 5447
rect 1109 5211 1345 5447
rect 1431 5211 1667 5447
rect 1753 5211 1989 5447
rect 2075 5211 2311 5447
rect 2397 5211 2633 5447
rect 2719 5211 2955 5447
rect 3041 5211 3277 5447
rect 3363 5211 3599 5447
rect 3685 5211 3921 5447
rect 4007 5211 4243 5447
rect 4329 5211 4565 5447
rect 4651 5211 4887 5447
rect 10111 5211 10347 5447
rect 10432 5211 10668 5447
rect 10753 5211 10989 5447
rect 11074 5211 11310 5447
rect 11395 5211 11631 5447
rect 11716 5211 11952 5447
rect 12037 5211 12273 5447
rect 12358 5211 12594 5447
rect 12679 5211 12915 5447
rect 13000 5211 13236 5447
rect 13321 5211 13557 5447
rect 13642 5211 13878 5447
rect 13963 5211 14199 5447
rect 14284 5211 14520 5447
rect 14605 5211 15000 5447
rect 0 5187 254 5211
rect 0 3977 254 4867
rect 14746 5187 15000 5211
rect 14746 3977 15000 4867
rect 0 3007 193 3657
rect 14807 3007 15000 3657
rect 0 1797 254 2687
rect 0 427 254 1477
rect 14746 1797 15000 2687
rect 14746 427 15000 1477
<< obsm5 >>
rect 574 34837 14426 40000
rect 0 19317 15000 34837
rect 574 7368 14426 19317
rect 0 7367 15000 7368
rect 574 6053 14426 7367
rect 701 5817 787 6053
rect 1023 5817 1109 6053
rect 1345 5817 1431 6053
rect 1667 5817 1753 6053
rect 1989 5817 2075 6053
rect 2311 5817 2397 6053
rect 2633 5817 2719 6053
rect 2955 5817 3041 6053
rect 3277 5817 3363 6053
rect 3599 5817 3685 6053
rect 3921 5817 4007 6053
rect 4243 5817 4329 6053
rect 4565 5817 4651 6053
rect 4887 5817 10111 6053
rect 10347 5817 10432 6053
rect 10668 5817 10753 6053
rect 10989 5817 11074 6053
rect 11310 5817 11395 6053
rect 11631 5817 11716 6053
rect 11952 5817 12037 6053
rect 12273 5817 12358 6053
rect 12594 5817 12679 6053
rect 12915 5817 13000 6053
rect 13236 5817 13321 6053
rect 13557 5817 13642 6053
rect 13878 5817 13963 6053
rect 14199 5817 14284 6053
rect 574 5447 14426 5817
rect 701 5211 787 5447
rect 1023 5211 1109 5447
rect 1345 5211 1431 5447
rect 1667 5211 1753 5447
rect 1989 5211 2075 5447
rect 2311 5211 2397 5447
rect 2633 5211 2719 5447
rect 2955 5211 3041 5447
rect 3277 5211 3363 5447
rect 3599 5211 3685 5447
rect 3921 5211 4007 5447
rect 4243 5211 4329 5447
rect 4565 5211 4651 5447
rect 4887 5211 10111 5447
rect 10347 5211 10432 5447
rect 10668 5211 10753 5447
rect 10989 5211 11074 5447
rect 11310 5211 11395 5447
rect 11631 5211 11716 5447
rect 11952 5211 12037 5447
rect 12273 5211 12358 5447
rect 12594 5211 12679 5447
rect 12915 5211 13000 5447
rect 13236 5211 13321 5447
rect 13557 5211 13642 5447
rect 13878 5211 13963 5447
rect 14199 5211 14284 5447
rect 574 3657 14426 5211
rect 513 3007 14487 3657
rect 574 427 14426 3007
<< labels >>
rlabel metal5 s 0 9547 254 11347 6 VSSA
port 1 nsew ground bidirectional
rlabel metal5 s 0 7368 254 8017 6 VSSA
port 1 nsew ground bidirectional
rlabel metal5 s 14746 9547 15000 11347 6 VSSA
port 1 nsew ground bidirectional
rlabel metal5 s 14746 7368 15000 8017 6 VSSA
port 1 nsew ground bidirectional
rlabel metal4 s 0 11281 15000 11347 6 VSSA
port 1 nsew ground bidirectional
rlabel metal4 s 0 9547 15000 9613 6 VSSA
port 1 nsew ground bidirectional
rlabel metal4 s 0 10329 254 10565 6 VSSA
port 1 nsew ground bidirectional
rlabel metal4 s 0 7347 254 8037 6 VSSA
port 1 nsew ground bidirectional
rlabel metal4 s 14746 10329 15000 10565 6 VSSA
port 1 nsew ground bidirectional
rlabel metal4 s 14746 7347 15000 8037 6 VSSA
port 1 nsew ground bidirectional
rlabel metal5 s 0 14007 254 18997 6 VDDIO
port 2 nsew power bidirectional
rlabel metal5 s 0 3977 254 4867 6 VDDIO
port 2 nsew power bidirectional
rlabel metal5 s 14746 14007 15000 18997 6 VDDIO
port 2 nsew power bidirectional
rlabel metal5 s 14746 3977 15000 4867 6 VDDIO
port 2 nsew power bidirectional
rlabel metal4 s 0 3957 254 4887 6 VDDIO
port 2 nsew power bidirectional
rlabel metal4 s 0 14007 254 19000 6 VDDIO
port 2 nsew power bidirectional
rlabel metal4 s 14746 3957 15000 4887 6 VDDIO
port 2 nsew power bidirectional
rlabel metal4 s 14746 14007 15000 19000 6 VDDIO
port 2 nsew power bidirectional
rlabel metal5 s 0 12837 254 13687 6 VDDIO_Q
port 3 nsew power bidirectional
rlabel metal5 s 14746 12837 15000 13687 6 VDDIO_Q
port 3 nsew power bidirectional
rlabel metal4 s 0 12817 254 13707 6 VDDIO_Q
port 3 nsew power bidirectional
rlabel metal4 s 14746 12817 15000 13707 6 VDDIO_Q
port 3 nsew power bidirectional
rlabel metal5 s 0 8337 254 9227 6 VSSD
port 4 nsew ground bidirectional
rlabel metal5 s 14746 8337 15000 9227 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 0 8317 254 9247 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 14746 8317 15000 9247 6 VSSD
port 4 nsew ground bidirectional
rlabel metal5 s 0 5187 254 6077 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 14746 5187 15000 6077 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 14746 35157 15000 40000 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 0 35157 254 40000 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 0 5167 254 6097 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14746 5167 15000 6097 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14746 35157 15000 40000 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 0 35157 254 40000 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 99 5168 4879 6096 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10078 5168 14858 6096 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2719 39246 2851 39394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2726 39434 12265 39986 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12136 39246 12268 39394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14800 6042 14840 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14800 5956 14840 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14800 5870 14840 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14800 5784 14840 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14800 5698 14840 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14800 5612 14840 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14800 5526 14840 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14800 5440 14840 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14800 5354 14840 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14800 5268 14840 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14800 5182 14840 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14786 39919 14850 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14786 39838 14850 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14786 39757 14850 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14786 39676 14850 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14786 39595 14850 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14786 39514 14850 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14786 39433 14850 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14786 39352 14850 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14786 39271 14850 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14786 39190 14850 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14786 39109 14850 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14786 39028 14850 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12306 35187 14746 39011 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12306 35187 14850 39011 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14719 6042 14759 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14719 5956 14759 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14719 5870 14759 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14719 5784 14759 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14719 5698 14759 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14719 5612 14759 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14719 5526 14759 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14719 5440 14759 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14719 5354 14759 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14719 5268 14759 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14719 5182 14759 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14706 39919 14746 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14706 39919 14770 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14706 39838 14746 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14706 39838 14770 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14706 39757 14746 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14706 39757 14770 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14706 39676 14746 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14706 39676 14770 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14706 39595 14746 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14706 39595 14770 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14706 39514 14746 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14706 39514 14770 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14706 39433 14746 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14706 39433 14770 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14706 39352 14746 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14706 39352 14770 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14706 39271 14746 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14706 39271 14770 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14706 39190 14746 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14706 39190 14770 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14706 39109 14746 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14706 39109 14770 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14706 39028 14746 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14706 39028 14770 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14626 39919 14690 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14626 39919 14690 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14626 39838 14690 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14626 39838 14690 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14626 39757 14690 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14626 39757 14690 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14626 39676 14690 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14626 39676 14690 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14626 39595 14690 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14626 39595 14690 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14626 39514 14690 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14626 39514 14690 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14626 39433 14690 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14626 39433 14690 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14626 39352 14690 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14626 39352 14690 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14626 39271 14690 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14626 39271 14690 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14626 39190 14690 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14626 39190 14690 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14626 39109 14690 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14626 39109 14690 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14626 39028 14690 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14626 39028 14690 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 6042 14678 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 14605 5817 14746 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14605 5817 14746 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14605 5817 14746 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 5698 14678 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 5612 14678 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 5526 14678 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 5440 14678 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 14605 5211 14746 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14605 5211 14746 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14605 5211 14746 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14546 39919 14610 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14546 39919 14610 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14546 39838 14610 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14546 39838 14610 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14546 39757 14610 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14546 39757 14610 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14546 39676 14610 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14546 39676 14610 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14546 39595 14610 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14546 39595 14610 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14546 39514 14610 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14546 39514 14610 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14546 39433 14610 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14546 39433 14610 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14546 39352 14610 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14546 39352 14610 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14546 39271 14610 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14546 39271 14610 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14546 39190 14610 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14546 39190 14610 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14546 39109 14610 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14546 39109 14610 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14546 39028 14610 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14546 39028 14610 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14557 6042 14597 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14557 5956 14597 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14557 5870 14597 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14557 5784 14597 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14557 5698 14597 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14557 5612 14597 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14557 5526 14597 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14557 5440 14597 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14557 5354 14597 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14557 5268 14597 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14557 5182 14597 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14466 39919 14530 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14466 39919 14530 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14466 39838 14530 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14466 39838 14530 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14466 39757 14530 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14466 39757 14530 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14466 39676 14530 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14466 39676 14530 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14466 39595 14530 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14466 39595 14530 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14466 39514 14530 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14466 39514 14530 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14466 39433 14530 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14466 39433 14530 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14466 39352 14530 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14466 39352 14530 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14466 39271 14530 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14466 39271 14530 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14466 39190 14530 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14466 39190 14530 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14466 39109 14530 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14466 39109 14530 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14466 39028 14530 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14466 39028 14530 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14476 6042 14516 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 14284 5817 14520 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14284 5817 14520 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14284 5817 14520 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14476 5698 14516 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14476 5612 14516 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14476 5526 14516 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14476 5440 14516 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 14284 5211 14520 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14284 5211 14520 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14284 5211 14520 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14386 39919 14450 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14386 39919 14450 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14386 39838 14450 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14386 39838 14450 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14386 39757 14450 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14386 39757 14450 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14386 39676 14450 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14386 39676 14450 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14386 39595 14450 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14386 39595 14450 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14386 39514 14450 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14386 39514 14450 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14386 39433 14450 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14386 39433 14450 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14386 39352 14450 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14386 39352 14450 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14386 39271 14450 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14386 39271 14450 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14386 39190 14450 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14386 39190 14450 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14386 39109 14450 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14386 39109 14450 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14386 39028 14450 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14386 39028 14450 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14395 5698 14435 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14395 5612 14435 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14395 5526 14435 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14306 39919 14370 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14306 39919 14370 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14306 39838 14370 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14306 39838 14370 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14306 39757 14370 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14306 39757 14370 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14306 39676 14370 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14306 39676 14370 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14306 39595 14370 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14306 39595 14370 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14306 39514 14370 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14306 39514 14370 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14306 39433 14370 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14306 39433 14370 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14306 39352 14370 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14306 39352 14370 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14306 39271 14370 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14306 39271 14370 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14306 39190 14370 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14306 39190 14370 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14306 39109 14370 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14306 39109 14370 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14306 39028 14370 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14306 39028 14370 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14314 5698 14354 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14314 5612 14354 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14314 5526 14354 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14226 39919 14290 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14226 39919 14290 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14226 39838 14290 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14226 39838 14290 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14226 39757 14290 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14226 39757 14290 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14226 39676 14290 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14226 39676 14290 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14226 39595 14290 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14226 39595 14290 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14226 39514 14290 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14226 39514 14290 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14226 39433 14290 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14226 39433 14290 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14226 39352 14290 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14226 39352 14290 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14226 39271 14290 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14226 39271 14290 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14226 39190 14290 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14226 39190 14290 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14226 39109 14290 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14226 39109 14290 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14226 39028 14290 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14226 39028 14290 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14233 6042 14273 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14233 5956 14273 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14233 5870 14273 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14233 5784 14273 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14233 5698 14273 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14233 5612 14273 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14233 5526 14273 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14233 5440 14273 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14233 5354 14273 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14233 5268 14273 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14233 5182 14273 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14146 39919 14210 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14146 39919 14210 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14146 39838 14210 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14146 39838 14210 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14146 39757 14210 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14146 39757 14210 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14146 39676 14210 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14146 39676 14210 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14146 39595 14210 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14146 39595 14210 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14146 39514 14210 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14146 39514 14210 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14146 39433 14210 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14146 39433 14210 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14146 39352 14210 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14146 39352 14210 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14146 39271 14210 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14146 39271 14210 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14146 39190 14210 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14146 39190 14210 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14146 39109 14210 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14146 39109 14210 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14146 39028 14210 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14146 39028 14210 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14152 6042 14192 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 13963 5817 14199 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13963 5817 14199 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13963 5817 14199 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14152 5698 14192 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14152 5612 14192 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14152 5526 14192 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14152 5440 14192 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 13963 5211 14199 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13963 5211 14199 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13963 5211 14199 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14066 39919 14130 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14066 39919 14130 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14066 39838 14130 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14066 39838 14130 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14066 39757 14130 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14066 39757 14130 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14066 39676 14130 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14066 39676 14130 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14066 39595 14130 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14066 39595 14130 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14066 39514 14130 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14066 39514 14130 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14066 39433 14130 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14066 39433 14130 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14066 39352 14130 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14066 39352 14130 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14066 39271 14130 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14066 39271 14130 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14066 39190 14130 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14066 39190 14130 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14066 39109 14130 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14066 39109 14130 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14066 39028 14130 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14066 39028 14130 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14071 5698 14111 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14071 5612 14111 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14071 5526 14111 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13986 39919 14050 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13986 39919 14050 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13986 39838 14050 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13986 39838 14050 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13986 39757 14050 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13986 39757 14050 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13986 39676 14050 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13986 39676 14050 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13986 39595 14050 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13986 39595 14050 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13986 39514 14050 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13986 39514 14050 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13986 39433 14050 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13986 39433 14050 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13986 39352 14050 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13986 39352 14050 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13986 39271 14050 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13986 39271 14050 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13986 39190 14050 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13986 39190 14050 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13986 39109 14050 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13986 39109 14050 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13986 39028 14050 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13986 39028 14050 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13990 5698 14030 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13990 5612 14030 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13990 5526 14030 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13906 39919 13970 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13906 39919 13970 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13906 39838 13970 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13906 39838 13970 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13906 39757 13970 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13906 39757 13970 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13906 39676 13970 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13906 39676 13970 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13906 39595 13970 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13906 39595 13970 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13906 39514 13970 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13906 39514 13970 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13906 39433 13970 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13906 39433 13970 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13906 39352 13970 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13906 39352 13970 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13906 39271 13970 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13906 39271 13970 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13906 39190 13970 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13906 39190 13970 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13906 39109 13970 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13906 39109 13970 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13906 39028 13970 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13906 39028 13970 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13909 6042 13949 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13909 5956 13949 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13909 5870 13949 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13909 5784 13949 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13909 5698 13949 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13909 5612 13949 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13909 5526 13949 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13909 5440 13949 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13909 5354 13949 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13909 5268 13949 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13909 5182 13949 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13826 39919 13890 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13826 39919 13890 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13826 39838 13890 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13826 39838 13890 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13826 39757 13890 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13826 39757 13890 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13826 39676 13890 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13826 39676 13890 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13826 39595 13890 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13826 39595 13890 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13826 39514 13890 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13826 39514 13890 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13826 39433 13890 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13826 39433 13890 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13826 39352 13890 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13826 39352 13890 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13826 39271 13890 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13826 39271 13890 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13826 39190 13890 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13826 39190 13890 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13826 39109 13890 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13826 39109 13890 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13826 39028 13890 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13826 39028 13890 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13828 6042 13868 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 13642 5817 13878 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13642 5817 13878 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13642 5817 13878 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13828 5698 13868 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13828 5612 13868 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13828 5526 13868 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13828 5440 13868 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 13642 5211 13878 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13642 5211 13878 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13642 5211 13878 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13746 39919 13810 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13746 39919 13810 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13746 39838 13810 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13746 39838 13810 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13746 39757 13810 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13746 39757 13810 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13746 39676 13810 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13746 39676 13810 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13746 39595 13810 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13746 39595 13810 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13746 39514 13810 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13746 39514 13810 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13746 39433 13810 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13746 39433 13810 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13746 39352 13810 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13746 39352 13810 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13746 39271 13810 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13746 39271 13810 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13746 39190 13810 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13746 39190 13810 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13746 39109 13810 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13746 39109 13810 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13746 39028 13810 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13746 39028 13810 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13747 5698 13787 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13747 5612 13787 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13747 5526 13787 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13666 39919 13730 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13666 39919 13730 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13666 39838 13730 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13666 39838 13730 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13666 39757 13730 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13666 39757 13730 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13666 39676 13730 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13666 39676 13730 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13666 39595 13730 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13666 39595 13730 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13666 39514 13730 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13666 39514 13730 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13666 39433 13730 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13666 39433 13730 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13666 39352 13730 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13666 39352 13730 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13666 39271 13730 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13666 39271 13730 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13666 39190 13730 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13666 39190 13730 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13666 39109 13730 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13666 39109 13730 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13666 39028 13730 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13666 39028 13730 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13666 5698 13706 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13666 5612 13706 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13666 5526 13706 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13586 39919 13650 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13586 39919 13650 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13586 39838 13650 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13586 39838 13650 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13586 39757 13650 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13586 39757 13650 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13586 39676 13650 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13586 39676 13650 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13586 39595 13650 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13586 39595 13650 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13586 39514 13650 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13586 39514 13650 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13586 39433 13650 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13586 39433 13650 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13586 39352 13650 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13586 39352 13650 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13586 39271 13650 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13586 39271 13650 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13586 39190 13650 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13586 39190 13650 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13586 39109 13650 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13586 39109 13650 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13586 39028 13650 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13586 39028 13650 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13585 6042 13625 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13585 5956 13625 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13585 5870 13625 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13585 5784 13625 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13585 5698 13625 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13585 5612 13625 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13585 5526 13625 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13585 5440 13625 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13585 5354 13625 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13585 5268 13625 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13585 5182 13625 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13506 39919 13570 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13506 39919 13570 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13506 39838 13570 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13506 39838 13570 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13506 39757 13570 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13506 39757 13570 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13506 39676 13570 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13506 39676 13570 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13506 39595 13570 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13506 39595 13570 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13506 39514 13570 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13506 39514 13570 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13506 39433 13570 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13506 39433 13570 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13506 39352 13570 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13506 39352 13570 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13506 39271 13570 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13506 39271 13570 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13506 39190 13570 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13506 39190 13570 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13506 39109 13570 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13506 39109 13570 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13506 39028 13570 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13506 39028 13570 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13504 6042 13544 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 13321 5817 13557 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13321 5817 13557 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13321 5817 13557 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13504 5698 13544 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13504 5612 13544 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13504 5526 13544 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13504 5440 13544 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 13321 5211 13557 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13321 5211 13557 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13321 5211 13557 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13426 39919 13490 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13426 39919 13490 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13426 39838 13490 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13426 39838 13490 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13426 39757 13490 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13426 39757 13490 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13426 39676 13490 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13426 39676 13490 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13426 39595 13490 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13426 39595 13490 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13426 39514 13490 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13426 39514 13490 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13426 39433 13490 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13426 39433 13490 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13426 39352 13490 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13426 39352 13490 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13426 39271 13490 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13426 39271 13490 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13426 39190 13490 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13426 39190 13490 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13426 39109 13490 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13426 39109 13490 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13426 39028 13490 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13426 39028 13490 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13423 5698 13463 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13423 5612 13463 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13423 5526 13463 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13346 39919 13410 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13346 39919 13410 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13346 39838 13410 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13346 39838 13410 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13346 39757 13410 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13346 39757 13410 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13346 39676 13410 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13346 39676 13410 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13346 39595 13410 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13346 39595 13410 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13346 39514 13410 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13346 39514 13410 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13346 39433 13410 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13346 39433 13410 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13346 39352 13410 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13346 39352 13410 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13346 39271 13410 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13346 39271 13410 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13346 39190 13410 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13346 39190 13410 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13346 39109 13410 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13346 39109 13410 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13346 39028 13410 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13346 39028 13410 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13342 5698 13382 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13342 5612 13382 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13342 5526 13382 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13266 39919 13330 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13266 39919 13330 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13266 39838 13330 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13266 39838 13330 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13266 39757 13330 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13266 39757 13330 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13266 39676 13330 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13266 39676 13330 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13266 39595 13330 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13266 39595 13330 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13266 39514 13330 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13266 39514 13330 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13266 39433 13330 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13266 39433 13330 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13266 39352 13330 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13266 39352 13330 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13266 39271 13330 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13266 39271 13330 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13266 39190 13330 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13266 39190 13330 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13266 39109 13330 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13266 39109 13330 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13266 39028 13330 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13266 39028 13330 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13261 6042 13301 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13261 5956 13301 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13261 5870 13301 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13261 5784 13301 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13261 5698 13301 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13261 5612 13301 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13261 5526 13301 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13261 5440 13301 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13261 5354 13301 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13261 5268 13301 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13261 5182 13301 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13186 39919 13250 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13186 39919 13250 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13186 39838 13250 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13186 39838 13250 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13186 39757 13250 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13186 39757 13250 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13186 39676 13250 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13186 39676 13250 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13186 39595 13250 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13186 39595 13250 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13186 39514 13250 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13186 39514 13250 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13186 39433 13250 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13186 39433 13250 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13186 39352 13250 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13186 39352 13250 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13186 39271 13250 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13186 39271 13250 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13186 39190 13250 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13186 39190 13250 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13186 39109 13250 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13186 39109 13250 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13186 39028 13250 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13186 39028 13250 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13180 6042 13220 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 13000 5817 13236 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13000 5817 13236 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13000 5817 13236 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13180 5698 13220 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13180 5612 13220 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13180 5526 13220 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13180 5440 13220 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 13000 5211 13236 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13000 5211 13236 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13000 5211 13236 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13106 39919 13170 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13106 39919 13170 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13106 39838 13170 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13106 39838 13170 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13106 39757 13170 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13106 39757 13170 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13106 39676 13170 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13106 39676 13170 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13106 39595 13170 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13106 39595 13170 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13106 39514 13170 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13106 39514 13170 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13106 39433 13170 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13106 39433 13170 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13106 39352 13170 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13106 39352 13170 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13106 39271 13170 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13106 39271 13170 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13106 39190 13170 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13106 39190 13170 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13106 39109 13170 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13106 39109 13170 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13106 39028 13170 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13106 39028 13170 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13099 5698 13139 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13099 5612 13139 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13099 5526 13139 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13026 39919 13090 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13026 39919 13090 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13026 39838 13090 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13026 39838 13090 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13026 39757 13090 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13026 39757 13090 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13026 39676 13090 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13026 39676 13090 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13026 39595 13090 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13026 39595 13090 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13026 39514 13090 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13026 39514 13090 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13026 39433 13090 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13026 39433 13090 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13026 39352 13090 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13026 39352 13090 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13026 39271 13090 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13026 39271 13090 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13026 39190 13090 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13026 39190 13090 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13026 39109 13090 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13026 39109 13090 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 13026 39028 13090 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13026 39028 13090 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13018 5698 13058 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13018 5612 13058 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13018 5526 13058 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12946 39919 13010 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12946 39919 13010 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12946 39838 13010 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12946 39838 13010 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12946 39757 13010 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12946 39757 13010 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12946 39676 13010 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12946 39676 13010 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12946 39595 13010 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12946 39595 13010 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12946 39514 13010 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12946 39514 13010 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12946 39433 13010 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12946 39433 13010 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12946 39352 13010 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12946 39352 13010 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12946 39271 13010 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12946 39271 13010 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12946 39190 13010 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12946 39190 13010 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12946 39109 13010 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12946 39109 13010 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12946 39028 13010 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12946 39028 13010 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12937 6042 12977 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12937 5956 12977 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12937 5870 12977 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12937 5784 12977 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12937 5698 12977 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12937 5612 12977 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12937 5526 12977 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12937 5440 12977 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12937 5354 12977 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12937 5268 12977 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12937 5182 12977 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12866 39919 12930 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12866 39919 12930 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12866 39838 12930 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12866 39838 12930 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12866 39757 12930 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12866 39757 12930 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12866 39676 12930 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12866 39676 12930 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12866 39595 12930 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12866 39595 12930 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12866 39514 12930 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12866 39514 12930 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12866 39433 12930 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12866 39433 12930 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12866 39352 12930 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12866 39352 12930 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12866 39271 12930 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12866 39271 12930 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12866 39190 12930 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12866 39190 12930 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12866 39109 12930 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12866 39109 12930 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12866 39028 12930 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12866 39028 12930 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12856 6042 12896 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 12679 5817 12915 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12679 5817 12915 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12679 5817 12915 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12856 5698 12896 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12856 5612 12896 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12856 5526 12896 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12856 5440 12896 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 12679 5211 12915 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12679 5211 12915 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12679 5211 12915 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12786 39919 12850 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12786 39919 12850 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12786 39838 12850 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12786 39838 12850 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12786 39757 12850 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12786 39757 12850 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12786 39676 12850 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12786 39676 12850 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12786 39595 12850 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12786 39595 12850 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12786 39514 12850 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12786 39514 12850 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12786 39433 12850 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12786 39433 12850 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12786 39352 12850 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12786 39352 12850 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12786 39271 12850 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12786 39271 12850 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12786 39190 12850 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12786 39190 12850 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12786 39109 12850 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12786 39109 12850 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12786 39028 12850 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12786 39028 12850 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12775 5698 12815 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12775 5612 12815 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12775 5526 12815 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12706 39919 12770 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12706 39919 12770 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12706 39838 12770 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12706 39838 12770 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12706 39757 12770 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12706 39757 12770 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12706 39676 12770 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12706 39676 12770 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12706 39595 12770 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12706 39595 12770 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12706 39514 12770 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12706 39514 12770 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12706 39433 12770 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12706 39433 12770 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12706 39352 12770 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12706 39352 12770 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12706 39271 12770 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12706 39271 12770 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12706 39190 12770 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12706 39190 12770 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12706 39109 12770 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12706 39109 12770 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12706 39028 12770 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12706 39028 12770 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12694 5698 12734 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12694 5612 12734 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12694 5526 12734 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12626 39919 12690 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12626 39919 12690 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12626 39838 12690 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12626 39838 12690 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12626 39757 12690 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12626 39757 12690 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12626 39676 12690 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12626 39676 12690 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12626 39595 12690 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12626 39595 12690 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12626 39514 12690 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12626 39514 12690 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12626 39433 12690 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12626 39433 12690 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12626 39352 12690 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12626 39352 12690 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12626 39271 12690 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12626 39271 12690 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12626 39190 12690 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12626 39190 12690 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12626 39109 12690 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12626 39109 12690 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12626 39028 12690 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12626 39028 12690 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12613 6042 12653 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12613 5956 12653 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12613 5870 12653 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12613 5784 12653 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12613 5698 12653 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12613 5612 12653 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12613 5526 12653 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12613 5440 12653 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12613 5354 12653 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12613 5268 12653 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12613 5182 12653 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12546 39919 12610 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12546 39919 12610 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12546 39838 12610 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12546 39838 12610 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12546 39757 12610 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12546 39757 12610 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12546 39676 12610 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12546 39676 12610 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12546 39595 12610 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12546 39595 12610 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12546 39514 12610 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12546 39514 12610 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12546 39433 12610 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12546 39433 12610 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12546 39352 12610 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12546 39352 12610 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12546 39271 12610 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12546 39271 12610 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12546 39190 12610 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12546 39190 12610 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12546 39109 12610 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12546 39109 12610 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12546 39028 12610 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12546 39028 12610 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12532 6042 12572 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 12358 5817 12594 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12358 5817 12594 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12358 5817 12594 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12532 5698 12572 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12532 5612 12572 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12532 5526 12572 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12532 5440 12572 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 12358 5211 12594 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12358 5211 12594 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12358 5211 12594 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12466 39919 12530 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12466 39919 12530 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12466 39838 12530 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12466 39838 12530 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12466 39757 12530 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12466 39757 12530 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12466 39676 12530 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12466 39676 12530 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12466 39595 12530 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12466 39595 12530 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12466 39514 12530 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12466 39514 12530 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12466 39433 12530 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12466 39433 12530 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12466 39352 12530 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12466 39352 12530 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12466 39271 12530 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12466 39271 12530 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12466 39190 12530 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12466 39190 12530 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12466 39109 12530 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12466 39109 12530 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12466 39028 12530 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12466 39028 12530 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12451 5698 12491 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12451 5612 12491 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12451 5526 12491 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12386 39919 12450 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12386 39919 12450 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12386 39838 12450 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12386 39838 12450 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12386 39757 12450 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12386 39757 12450 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12386 39676 12450 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12386 39676 12450 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12386 39595 12450 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12386 39595 12450 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12386 39514 12450 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12386 39514 12450 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12386 39433 12450 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12386 39433 12450 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12386 39352 12450 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12386 39352 12450 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12386 39271 12450 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12386 39271 12450 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12386 39190 12450 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12386 39190 12450 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12386 39109 12450 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12386 39109 12450 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12386 39028 12450 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12386 39028 12450 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12370 5698 12410 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12370 5612 12410 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12370 5526 12410 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12306 39919 12370 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12306 39919 12370 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12306 39838 12370 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12306 39838 12370 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12306 39757 12370 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12306 39757 12370 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12306 39676 12370 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12306 39676 12370 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12306 39595 12370 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12306 39595 12370 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12306 39514 12370 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12306 39514 12370 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12306 39433 12370 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12306 39433 12370 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12306 39352 12370 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12306 39352 12370 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12306 39271 12370 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12306 39271 12370 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12306 39190 12370 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12306 39190 12370 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12306 39109 12370 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12306 39109 12370 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12306 39028 12370 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12306 39028 12370 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12289 6042 12329 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12289 5956 12329 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12289 5870 12329 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12289 5784 12329 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12289 5698 12329 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12289 5612 12329 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12289 5526 12329 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12289 5440 12329 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12289 5354 12329 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12289 5268 12329 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12289 5182 12329 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7417 39438 12264 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12208 6042 12248 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 12037 5817 12273 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12037 5817 12273 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12037 5817 12273 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12208 5698 12248 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12208 5612 12248 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12208 5526 12248 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12208 5440 12248 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 12037 5211 12273 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12037 5211 12273 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12037 5211 12273 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12170 39329 12234 39393 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12170 39247 12234 39311 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12127 5698 12167 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12127 5612 12167 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12127 5526 12167 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12046 5698 12086 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12046 5612 12086 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12046 5526 12086 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11965 6042 12005 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11965 5956 12005 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11965 5870 12005 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11965 5784 12005 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11965 5698 12005 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11965 5612 12005 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11965 5526 12005 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11965 5440 12005 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11965 5354 12005 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11965 5268 12005 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11965 5182 12005 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11884 6042 11924 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 11716 5817 11952 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 11716 5817 11952 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11716 5817 11952 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11884 5698 11924 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11884 5612 11924 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11884 5526 11924 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11884 5440 11924 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 11716 5211 11952 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 11716 5211 11952 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11716 5211 11952 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11803 5698 11843 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11803 5612 11843 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11803 5526 11843 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11722 5698 11762 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11722 5612 11762 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11722 5526 11762 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11641 6042 11681 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11641 5956 11681 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11641 5870 11681 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11641 5784 11681 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11641 5698 11681 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11641 5612 11681 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11641 5526 11681 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11641 5440 11681 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11641 5354 11681 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11641 5268 11681 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11641 5182 11681 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11560 6042 11600 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 11395 5817 11631 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 11395 5817 11631 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11395 5817 11631 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11560 5698 11600 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11560 5612 11600 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11560 5526 11600 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11560 5440 11600 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 11395 5211 11631 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 11395 5211 11631 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11395 5211 11631 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11479 5698 11519 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11479 5612 11519 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11479 5526 11519 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11398 5698 11438 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11398 5612 11438 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11398 5526 11438 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11317 6042 11357 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11317 5956 11357 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11317 5870 11357 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11317 5784 11357 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11317 5698 11357 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11317 5612 11357 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11317 5526 11357 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11317 5440 11357 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11317 5354 11357 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11317 5268 11357 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11317 5182 11357 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11236 6042 11276 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 11074 5817 11310 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 11074 5817 11310 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11074 5817 11310 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11236 5698 11276 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11236 5612 11276 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11236 5526 11276 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11236 5440 11276 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 11074 5211 11310 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 11074 5211 11310 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11074 5211 11310 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11155 5698 11195 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11155 5612 11195 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11155 5526 11195 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11074 5698 11114 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11074 5612 11114 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11074 5526 11114 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10993 6042 11033 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10993 5956 11033 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10993 5870 11033 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10993 5784 11033 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10993 5698 11033 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10993 5612 11033 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10993 5526 11033 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10993 5440 11033 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10993 5354 11033 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10993 5268 11033 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10993 5182 11033 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10912 6042 10952 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 10753 5817 10989 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 10753 5817 10989 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10753 5817 10989 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10912 5698 10952 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10912 5612 10952 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10912 5526 10952 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10912 5440 10952 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 10753 5211 10989 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 10753 5211 10989 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10753 5211 10989 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10831 5698 10871 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10831 5612 10871 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10831 5526 10871 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10750 5698 10790 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10750 5612 10790 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10750 5526 10790 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10669 6042 10709 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10669 5956 10709 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10669 5870 10709 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10669 5784 10709 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10669 5698 10709 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10669 5612 10709 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10669 5526 10709 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10669 5440 10709 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10669 5354 10709 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10669 5268 10709 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10669 5182 10709 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10588 6042 10628 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 10432 5817 10668 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 10432 5817 10668 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10432 5817 10668 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10588 5698 10628 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10588 5612 10628 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10588 5526 10628 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10588 5440 10628 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 10432 5211 10668 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 10432 5211 10668 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10432 5211 10668 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10506 5698 10546 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10506 5612 10546 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10506 5526 10546 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10424 5698 10464 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10424 5612 10464 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10424 5526 10464 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10342 6042 10382 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10342 5956 10382 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10342 5870 10382 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10342 5784 10382 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10342 5698 10382 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10342 5612 10382 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10342 5526 10382 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10342 5440 10382 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10342 5354 10382 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10342 5268 10382 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10342 5182 10382 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10260 6042 10300 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 10111 5817 10347 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 10111 5817 10347 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10111 5817 10347 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10260 5698 10300 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10260 5612 10300 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10260 5526 10300 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10260 5440 10300 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 10111 5211 10347 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 10111 5211 10347 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10111 5211 10347 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10178 5698 10218 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10178 5612 10218 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10178 5526 10218 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10096 5698 10136 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10096 5612 10136 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10096 5526 10136 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5400 39438 7417 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5319 39918 5383 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5319 39838 5383 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5319 39758 5383 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5319 39678 5383 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5319 39598 5383 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5319 39518 5383 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5319 39438 5383 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5238 39918 5302 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5238 39838 5302 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5238 39758 5302 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5238 39678 5302 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5238 39598 5302 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5238 39518 5302 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5238 39438 5302 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5157 39918 5221 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5157 39838 5221 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5157 39758 5221 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5157 39678 5221 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5157 39598 5221 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5157 39518 5221 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5157 39438 5221 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5076 39918 5140 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5076 39838 5140 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5076 39758 5140 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5076 39678 5140 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5076 39598 5140 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5076 39518 5140 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5076 39438 5140 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4995 39918 5059 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4995 39838 5059 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4995 39758 5059 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4995 39678 5059 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4995 39598 5059 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4995 39518 5059 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4995 39438 5059 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4914 39918 4978 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4914 39838 4978 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4914 39758 4978 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4914 39678 4978 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4914 39598 4978 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4914 39518 4978 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4914 39438 4978 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4833 39918 4897 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4833 39838 4897 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4833 39758 4897 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4833 39678 4897 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4833 39598 4897 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4833 39518 4897 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4833 39438 4897 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4821 6042 4861 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 4651 5817 4887 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 4651 5817 4887 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4651 5817 4887 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4821 5698 4861 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4821 5612 4861 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4821 5526 4861 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4821 5440 4861 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 4651 5211 4887 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 4651 5211 4887 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4651 5211 4887 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4752 39918 4816 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4752 39838 4816 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4752 39758 4816 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4752 39678 4816 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4752 39598 4816 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4752 39518 4816 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4752 39438 4816 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4740 5698 4780 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4740 5612 4780 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4740 5526 4780 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4671 39918 4735 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4671 39838 4735 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4671 39758 4735 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4671 39678 4735 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4671 39598 4735 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4671 39518 4735 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4671 39438 4735 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4659 5698 4699 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4659 5612 4699 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4659 5526 4699 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4590 39918 4654 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4590 39838 4654 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4590 39758 4654 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4590 39678 4654 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4590 39598 4654 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4590 39518 4654 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4590 39438 4654 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4578 6042 4618 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4578 5956 4618 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4578 5870 4618 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4578 5784 4618 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4578 5698 4618 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4578 5612 4618 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4578 5526 4618 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4578 5440 4618 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4578 5354 4618 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4578 5268 4618 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4578 5182 4618 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4509 39918 4573 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4509 39838 4573 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4509 39758 4573 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4509 39678 4573 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4509 39598 4573 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4509 39518 4573 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4509 39438 4573 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4497 6042 4537 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 4329 5817 4565 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 4329 5817 4565 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4329 5817 4565 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4497 5698 4537 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4497 5612 4537 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4497 5526 4537 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4497 5440 4537 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 4329 5211 4565 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 4329 5211 4565 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4329 5211 4565 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4428 39918 4492 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4428 39838 4492 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4428 39758 4492 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4428 39678 4492 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4428 39598 4492 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4428 39518 4492 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4428 39438 4492 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4416 5698 4456 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4416 5612 4456 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4416 5526 4456 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4347 39918 4411 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4347 39838 4411 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4347 39758 4411 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4347 39678 4411 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4347 39598 4411 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4347 39518 4411 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4347 39438 4411 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4335 5698 4375 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4335 5612 4375 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4335 5526 4375 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4266 39918 4330 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4266 39838 4330 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4266 39758 4330 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4266 39678 4330 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4266 39598 4330 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4266 39518 4330 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4266 39438 4330 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4254 6042 4294 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4254 5956 4294 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4254 5870 4294 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4254 5784 4294 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4254 5698 4294 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4254 5612 4294 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4254 5526 4294 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4254 5440 4294 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4254 5354 4294 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4254 5268 4294 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4254 5182 4294 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4185 39918 4249 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4185 39838 4249 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4185 39758 4249 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4185 39678 4249 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4185 39598 4249 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4185 39518 4249 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4185 39438 4249 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4173 6042 4213 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 4007 5817 4243 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 4007 5817 4243 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4007 5817 4243 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4173 5698 4213 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4173 5612 4213 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4173 5526 4213 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4173 5440 4213 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 4007 5211 4243 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 4007 5211 4243 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4007 5211 4243 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4104 39918 4168 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4104 39838 4168 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4104 39758 4168 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4104 39678 4168 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4104 39598 4168 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4104 39518 4168 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4104 39438 4168 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4092 5698 4132 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4092 5612 4132 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4092 5526 4132 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4023 39918 4087 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4023 39838 4087 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4023 39758 4087 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4023 39678 4087 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4023 39598 4087 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4023 39518 4087 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4023 39438 4087 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4011 5698 4051 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4011 5612 4051 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4011 5526 4051 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3942 39918 4006 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3942 39838 4006 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3942 39758 4006 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3942 39678 4006 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3942 39598 4006 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3942 39518 4006 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3942 39438 4006 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3930 6042 3970 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3930 5956 3970 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3930 5870 3970 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3930 5784 3970 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3930 5698 3970 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3930 5612 3970 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3930 5526 3970 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3930 5440 3970 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3930 5354 3970 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3930 5268 3970 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3930 5182 3970 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3861 39918 3925 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3861 39838 3925 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3861 39758 3925 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3861 39678 3925 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3861 39598 3925 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3861 39518 3925 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3861 39438 3925 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3849 6042 3889 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 3685 5817 3921 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 3685 5817 3921 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3685 5817 3921 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3849 5698 3889 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3849 5612 3889 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3849 5526 3889 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3849 5440 3889 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 3685 5211 3921 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 3685 5211 3921 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3685 5211 3921 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3780 39918 3844 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3780 39838 3844 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3780 39758 3844 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3780 39678 3844 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3780 39598 3844 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3780 39518 3844 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3780 39438 3844 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3768 5698 3808 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3768 5612 3808 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3768 5526 3808 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3699 39918 3763 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3699 39838 3763 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3699 39758 3763 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3699 39678 3763 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3699 39598 3763 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3699 39518 3763 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3699 39438 3763 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3687 5698 3727 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3687 5612 3727 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3687 5526 3727 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3618 39918 3682 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3618 39838 3682 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3618 39758 3682 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3618 39678 3682 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3618 39598 3682 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3618 39518 3682 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3618 39438 3682 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3606 6042 3646 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3606 5956 3646 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3606 5870 3646 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3606 5784 3646 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3606 5698 3646 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3606 5612 3646 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3606 5526 3646 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3606 5440 3646 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3606 5354 3646 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3606 5268 3646 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3606 5182 3646 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3537 39918 3601 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3537 39838 3601 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3537 39758 3601 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3537 39678 3601 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3537 39598 3601 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3537 39518 3601 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3537 39438 3601 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3525 6042 3565 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 3363 5817 3599 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 3363 5817 3599 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3363 5817 3599 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3525 5698 3565 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3525 5612 3565 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3525 5526 3565 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3525 5440 3565 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 3363 5211 3599 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 3363 5211 3599 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3363 5211 3599 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3456 39918 3520 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3456 39838 3520 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3456 39758 3520 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3456 39678 3520 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3456 39598 3520 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3456 39518 3520 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3456 39438 3520 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3444 5698 3484 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3444 5612 3484 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3444 5526 3484 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3375 39918 3439 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3375 39838 3439 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3375 39758 3439 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3375 39678 3439 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3375 39598 3439 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3375 39518 3439 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3375 39438 3439 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3363 5698 3403 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3363 5612 3403 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3363 5526 3403 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3294 39918 3358 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3294 39838 3358 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3294 39758 3358 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3294 39678 3358 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3294 39598 3358 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3294 39518 3358 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3294 39438 3358 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3282 6042 3322 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3282 5956 3322 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3282 5870 3322 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3282 5784 3322 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3282 5698 3322 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3282 5612 3322 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3282 5526 3322 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3282 5440 3322 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3282 5354 3322 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3282 5268 3322 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3282 5182 3322 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3213 39918 3277 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3213 39838 3277 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3213 39758 3277 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3213 39678 3277 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3213 39598 3277 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3213 39518 3277 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3213 39438 3277 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3201 6042 3241 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 3041 5817 3277 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 3041 5817 3277 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3041 5817 3277 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3201 5698 3241 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3201 5612 3241 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3201 5526 3241 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3201 5440 3241 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 3041 5211 3277 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 3041 5211 3277 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3041 5211 3277 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3132 39918 3196 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3132 39838 3196 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3132 39758 3196 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3132 39678 3196 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3132 39598 3196 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3132 39518 3196 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3132 39438 3196 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3120 5698 3160 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3120 5612 3160 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3120 5526 3160 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3051 39918 3115 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3051 39838 3115 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3051 39758 3115 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3051 39678 3115 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3051 39598 3115 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3051 39518 3115 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3051 39438 3115 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3039 5698 3079 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3039 5612 3079 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3039 5526 3079 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2970 39918 3034 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2970 39838 3034 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2970 39758 3034 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2970 39678 3034 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2970 39598 3034 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2970 39518 3034 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2970 39438 3034 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2958 6042 2998 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2958 5956 2998 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2958 5870 2998 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2958 5784 2998 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2958 5698 2998 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2958 5612 2998 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2958 5526 2998 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2958 5440 2998 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2958 5354 2998 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2958 5268 2998 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2958 5182 2998 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2889 39918 2953 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2889 39838 2953 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2889 39758 2953 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2889 39678 2953 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2889 39598 2953 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2889 39518 2953 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2889 39438 2953 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2877 6042 2917 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 2719 5817 2955 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2719 5817 2955 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2719 5817 2955 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2877 5698 2917 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2877 5612 2917 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2877 5526 2917 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2877 5440 2917 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 2719 5211 2955 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2719 5211 2955 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2719 5211 2955 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2808 39918 2872 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2808 39838 2872 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2808 39758 2872 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2808 39678 2872 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2808 39598 2872 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2808 39518 2872 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2808 39438 2872 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2796 5698 2836 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2796 5612 2836 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2796 5526 2836 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2753 39329 2817 39393 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2753 39247 2817 39311 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2727 39918 2791 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2727 39838 2791 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2727 39758 2791 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2727 39678 2791 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2727 39598 2791 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2727 39518 2791 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2727 39438 2791 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2715 5698 2755 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2715 5612 2755 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2715 5526 2755 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2634 6042 2674 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2634 5956 2674 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2634 5870 2674 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2634 5784 2674 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2634 5698 2674 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2634 5612 2674 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2634 5526 2674 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2634 5440 2674 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2634 5354 2674 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2634 5268 2674 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2634 5182 2674 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2605 39919 2669 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2605 39919 2669 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2605 39838 2669 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2605 39838 2669 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2605 39757 2669 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2605 39757 2669 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2605 39676 2669 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2605 39676 2669 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2605 39595 2669 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2605 39595 2669 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2605 39514 2669 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2605 39514 2669 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2605 39433 2669 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2605 39433 2669 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2605 39352 2669 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2605 39352 2669 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2605 39271 2669 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2605 39271 2669 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2605 39190 2669 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2605 39190 2669 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2605 39109 2669 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2605 39109 2669 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2605 39028 2669 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2605 39028 2669 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 254 35187 2669 39011 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 125 35187 2669 39011 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2553 6042 2593 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 2397 5817 2633 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2397 5817 2633 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2397 5817 2633 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2553 5698 2593 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2553 5612 2593 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2553 5526 2593 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2553 5440 2593 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 2397 5211 2633 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2397 5211 2633 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2397 5211 2633 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2525 39919 2589 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2525 39919 2589 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2525 39838 2589 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2525 39838 2589 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2525 39757 2589 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2525 39757 2589 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2525 39676 2589 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2525 39676 2589 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2525 39595 2589 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2525 39595 2589 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2525 39514 2589 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2525 39514 2589 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2525 39433 2589 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2525 39433 2589 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2525 39352 2589 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2525 39352 2589 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2525 39271 2589 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2525 39271 2589 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2525 39190 2589 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2525 39190 2589 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2525 39109 2589 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2525 39109 2589 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2525 39028 2589 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2525 39028 2589 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2472 5698 2512 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2472 5612 2512 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2472 5526 2512 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2445 39919 2509 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2445 39919 2509 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2445 39838 2509 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2445 39838 2509 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2445 39757 2509 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2445 39757 2509 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2445 39676 2509 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2445 39676 2509 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2445 39595 2509 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2445 39595 2509 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2445 39514 2509 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2445 39514 2509 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2445 39433 2509 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2445 39433 2509 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2445 39352 2509 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2445 39352 2509 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2445 39271 2509 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2445 39271 2509 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2445 39190 2509 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2445 39190 2509 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2445 39109 2509 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2445 39109 2509 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2445 39028 2509 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2445 39028 2509 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2391 5698 2431 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2391 5612 2431 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2391 5526 2431 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2365 39919 2429 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2365 39919 2429 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2365 39838 2429 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2365 39838 2429 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2365 39757 2429 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2365 39757 2429 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2365 39676 2429 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2365 39676 2429 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2365 39595 2429 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2365 39595 2429 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2365 39514 2429 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2365 39514 2429 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2365 39433 2429 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2365 39433 2429 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2365 39352 2429 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2365 39352 2429 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2365 39271 2429 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2365 39271 2429 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2365 39190 2429 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2365 39190 2429 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2365 39109 2429 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2365 39109 2429 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2365 39028 2429 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2365 39028 2429 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2310 6042 2350 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2310 5956 2350 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2310 5870 2350 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2310 5784 2350 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2310 5698 2350 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2310 5612 2350 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2310 5526 2350 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2310 5440 2350 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2310 5354 2350 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2310 5268 2350 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2310 5182 2350 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2285 39919 2349 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2285 39919 2349 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2285 39838 2349 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2285 39838 2349 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2285 39757 2349 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2285 39757 2349 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2285 39676 2349 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2285 39676 2349 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2285 39595 2349 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2285 39595 2349 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2285 39514 2349 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2285 39514 2349 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2285 39433 2349 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2285 39433 2349 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2285 39352 2349 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2285 39352 2349 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2285 39271 2349 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2285 39271 2349 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2285 39190 2349 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2285 39190 2349 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2285 39109 2349 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2285 39109 2349 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2285 39028 2349 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2285 39028 2349 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2229 6042 2269 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 2075 5817 2311 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2075 5817 2311 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2075 5817 2311 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2229 5698 2269 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2229 5612 2269 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2229 5526 2269 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2229 5440 2269 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 2075 5211 2311 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2075 5211 2311 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2075 5211 2311 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2205 39919 2269 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2205 39919 2269 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2205 39838 2269 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2205 39838 2269 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2205 39757 2269 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2205 39757 2269 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2205 39676 2269 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2205 39676 2269 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2205 39595 2269 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2205 39595 2269 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2205 39514 2269 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2205 39514 2269 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2205 39433 2269 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2205 39433 2269 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2205 39352 2269 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2205 39352 2269 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2205 39271 2269 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2205 39271 2269 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2205 39190 2269 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2205 39190 2269 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2205 39109 2269 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2205 39109 2269 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2205 39028 2269 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2205 39028 2269 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2148 5698 2188 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2148 5612 2188 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2148 5526 2188 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2125 39919 2189 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2125 39919 2189 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2125 39838 2189 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2125 39838 2189 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2125 39757 2189 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2125 39757 2189 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2125 39676 2189 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2125 39676 2189 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2125 39595 2189 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2125 39595 2189 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2125 39514 2189 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2125 39514 2189 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2125 39433 2189 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2125 39433 2189 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2125 39352 2189 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2125 39352 2189 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2125 39271 2189 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2125 39271 2189 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2125 39190 2189 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2125 39190 2189 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2125 39109 2189 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2125 39109 2189 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2125 39028 2189 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2125 39028 2189 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2067 5698 2107 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2067 5612 2107 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2067 5526 2107 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2045 39919 2109 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2045 39919 2109 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2045 39838 2109 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2045 39838 2109 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2045 39757 2109 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2045 39757 2109 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2045 39676 2109 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2045 39676 2109 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2045 39595 2109 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2045 39595 2109 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2045 39514 2109 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2045 39514 2109 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2045 39433 2109 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2045 39433 2109 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2045 39352 2109 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2045 39352 2109 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2045 39271 2109 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2045 39271 2109 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2045 39190 2109 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2045 39190 2109 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2045 39109 2109 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2045 39109 2109 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2045 39028 2109 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2045 39028 2109 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1986 6042 2026 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1986 5956 2026 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1986 5870 2026 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1986 5784 2026 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1986 5698 2026 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1986 5612 2026 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1986 5526 2026 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1986 5440 2026 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1986 5354 2026 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1986 5268 2026 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1986 5182 2026 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1965 39919 2029 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1965 39919 2029 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1965 39838 2029 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1965 39838 2029 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1965 39757 2029 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1965 39757 2029 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1965 39676 2029 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1965 39676 2029 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1965 39595 2029 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1965 39595 2029 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1965 39514 2029 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1965 39514 2029 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1965 39433 2029 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1965 39433 2029 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1965 39352 2029 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1965 39352 2029 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1965 39271 2029 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1965 39271 2029 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1965 39190 2029 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1965 39190 2029 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1965 39109 2029 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1965 39109 2029 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1965 39028 2029 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1965 39028 2029 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1905 6042 1945 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 1753 5817 1989 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1753 5817 1989 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1753 5817 1989 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1905 5698 1945 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1905 5612 1945 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1905 5526 1945 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1905 5440 1945 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 1753 5211 1989 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1753 5211 1989 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1753 5211 1989 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1885 39919 1949 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1885 39919 1949 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1885 39838 1949 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1885 39838 1949 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1885 39757 1949 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1885 39757 1949 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1885 39676 1949 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1885 39676 1949 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1885 39595 1949 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1885 39595 1949 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1885 39514 1949 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1885 39514 1949 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1885 39433 1949 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1885 39433 1949 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1885 39352 1949 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1885 39352 1949 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1885 39271 1949 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1885 39271 1949 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1885 39190 1949 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1885 39190 1949 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1885 39109 1949 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1885 39109 1949 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1885 39028 1949 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1885 39028 1949 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1824 5698 1864 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1824 5612 1864 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1824 5526 1864 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1805 39919 1869 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1805 39919 1869 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1805 39838 1869 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1805 39838 1869 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1805 39757 1869 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1805 39757 1869 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1805 39676 1869 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1805 39676 1869 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1805 39595 1869 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1805 39595 1869 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1805 39514 1869 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1805 39514 1869 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1805 39433 1869 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1805 39433 1869 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1805 39352 1869 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1805 39352 1869 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1805 39271 1869 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1805 39271 1869 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1805 39190 1869 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1805 39190 1869 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1805 39109 1869 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1805 39109 1869 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1805 39028 1869 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1805 39028 1869 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1743 5698 1783 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1743 5612 1783 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1743 5526 1783 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1725 39919 1789 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1725 39919 1789 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1725 39838 1789 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1725 39838 1789 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1725 39757 1789 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1725 39757 1789 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1725 39676 1789 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1725 39676 1789 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1725 39595 1789 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1725 39595 1789 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1725 39514 1789 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1725 39514 1789 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1725 39433 1789 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1725 39433 1789 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1725 39352 1789 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1725 39352 1789 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1725 39271 1789 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1725 39271 1789 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1725 39190 1789 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1725 39190 1789 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1725 39109 1789 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1725 39109 1789 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1725 39028 1789 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1725 39028 1789 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1662 6042 1702 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1662 5956 1702 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1662 5870 1702 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1662 5784 1702 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1662 5698 1702 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1662 5612 1702 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1662 5526 1702 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1662 5440 1702 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1662 5354 1702 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1662 5268 1702 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1662 5182 1702 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1645 39919 1709 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1645 39919 1709 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1645 39838 1709 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1645 39838 1709 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1645 39757 1709 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1645 39757 1709 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1645 39676 1709 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1645 39676 1709 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1645 39595 1709 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1645 39595 1709 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1645 39514 1709 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1645 39514 1709 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1645 39433 1709 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1645 39433 1709 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1645 39352 1709 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1645 39352 1709 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1645 39271 1709 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1645 39271 1709 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1645 39190 1709 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1645 39190 1709 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1645 39109 1709 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1645 39109 1709 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1645 39028 1709 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1645 39028 1709 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1581 6042 1621 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 1431 5817 1667 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1431 5817 1667 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1431 5817 1667 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1581 5698 1621 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1581 5612 1621 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1581 5526 1621 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1581 5440 1621 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 1431 5211 1667 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1431 5211 1667 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1431 5211 1667 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1565 39919 1629 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1565 39919 1629 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1565 39838 1629 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1565 39838 1629 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1565 39757 1629 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1565 39757 1629 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1565 39676 1629 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1565 39676 1629 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1565 39595 1629 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1565 39595 1629 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1565 39514 1629 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1565 39514 1629 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1565 39433 1629 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1565 39433 1629 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1565 39352 1629 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1565 39352 1629 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1565 39271 1629 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1565 39271 1629 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1565 39190 1629 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1565 39190 1629 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1565 39109 1629 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1565 39109 1629 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1565 39028 1629 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1565 39028 1629 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1500 5698 1540 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1500 5612 1540 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1500 5526 1540 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1485 39919 1549 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1485 39919 1549 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1485 39838 1549 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1485 39838 1549 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1485 39757 1549 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1485 39757 1549 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1485 39676 1549 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1485 39676 1549 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1485 39595 1549 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1485 39595 1549 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1485 39514 1549 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1485 39514 1549 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1485 39433 1549 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1485 39433 1549 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1485 39352 1549 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1485 39352 1549 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1485 39271 1549 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1485 39271 1549 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1485 39190 1549 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1485 39190 1549 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1485 39109 1549 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1485 39109 1549 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1485 39028 1549 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1485 39028 1549 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1419 5698 1459 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1419 5612 1459 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1419 5526 1459 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1405 39919 1469 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1405 39919 1469 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1405 39838 1469 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1405 39838 1469 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1405 39757 1469 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1405 39757 1469 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1405 39676 1469 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1405 39676 1469 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1405 39595 1469 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1405 39595 1469 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1405 39514 1469 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1405 39514 1469 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1405 39433 1469 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1405 39433 1469 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1405 39352 1469 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1405 39352 1469 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1405 39271 1469 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1405 39271 1469 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1405 39190 1469 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1405 39190 1469 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1405 39109 1469 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1405 39109 1469 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1405 39028 1469 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1405 39028 1469 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1338 6042 1378 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1338 5956 1378 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1338 5870 1378 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1338 5784 1378 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1338 5698 1378 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1338 5612 1378 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1338 5526 1378 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1338 5440 1378 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1338 5354 1378 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1338 5268 1378 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1338 5182 1378 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1325 39919 1389 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1325 39919 1389 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1325 39838 1389 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1325 39838 1389 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1325 39757 1389 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1325 39757 1389 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1325 39676 1389 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1325 39676 1389 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1325 39595 1389 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1325 39595 1389 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1325 39514 1389 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1325 39514 1389 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1325 39433 1389 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1325 39433 1389 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1325 39352 1389 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1325 39352 1389 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1325 39271 1389 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1325 39271 1389 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1325 39190 1389 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1325 39190 1389 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1325 39109 1389 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1325 39109 1389 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1325 39028 1389 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1325 39028 1389 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1245 39919 1309 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1245 39919 1309 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1245 39838 1309 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1245 39838 1309 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1245 39757 1309 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1245 39757 1309 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1245 39676 1309 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1245 39676 1309 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1245 39595 1309 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1245 39595 1309 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1245 39514 1309 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1245 39514 1309 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1245 39433 1309 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1245 39433 1309 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1245 39352 1309 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1245 39352 1309 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1245 39271 1309 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1245 39271 1309 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1245 39190 1309 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1245 39190 1309 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1245 39109 1309 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1245 39109 1309 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1245 39028 1309 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1245 39028 1309 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 6042 1297 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 1109 5817 1345 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1109 5817 1345 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1109 5817 1345 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 5698 1297 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 5612 1297 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 5526 1297 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 5440 1297 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 1109 5211 1345 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1109 5211 1345 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1109 5211 1345 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1165 39919 1229 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1165 39919 1229 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1165 39838 1229 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1165 39838 1229 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1165 39757 1229 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1165 39757 1229 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1165 39676 1229 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1165 39676 1229 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1165 39595 1229 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1165 39595 1229 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1165 39514 1229 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1165 39514 1229 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1165 39433 1229 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1165 39433 1229 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1165 39352 1229 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1165 39352 1229 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1165 39271 1229 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1165 39271 1229 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1165 39190 1229 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1165 39190 1229 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1165 39109 1229 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1165 39109 1229 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1165 39028 1229 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1165 39028 1229 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1176 5698 1216 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1176 5612 1216 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1176 5526 1216 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1085 39919 1149 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1085 39919 1149 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1085 39838 1149 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1085 39838 1149 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1085 39757 1149 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1085 39757 1149 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1085 39676 1149 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1085 39676 1149 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1085 39595 1149 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1085 39595 1149 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1085 39514 1149 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1085 39514 1149 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1085 39433 1149 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1085 39433 1149 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1085 39352 1149 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1085 39352 1149 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1085 39271 1149 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1085 39271 1149 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1085 39190 1149 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1085 39190 1149 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1085 39109 1149 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1085 39109 1149 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1085 39028 1149 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1085 39028 1149 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1095 5698 1135 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1095 5612 1135 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1095 5526 1135 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1005 39919 1069 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1005 39919 1069 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1005 39838 1069 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1005 39838 1069 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1005 39757 1069 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1005 39757 1069 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1005 39676 1069 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1005 39676 1069 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1005 39595 1069 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1005 39595 1069 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1005 39514 1069 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1005 39514 1069 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1005 39433 1069 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1005 39433 1069 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1005 39352 1069 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1005 39352 1069 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1005 39271 1069 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1005 39271 1069 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1005 39190 1069 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1005 39190 1069 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1005 39109 1069 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1005 39109 1069 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 1005 39028 1069 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1005 39028 1069 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1014 6042 1054 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1014 5956 1054 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1014 5870 1054 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1014 5784 1054 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1014 5698 1054 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1014 5612 1054 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1014 5526 1054 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1014 5440 1054 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1014 5354 1054 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1014 5268 1054 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1014 5182 1054 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 925 39919 989 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 925 39919 989 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 925 39838 989 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 925 39838 989 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 925 39757 989 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 925 39757 989 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 925 39676 989 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 925 39676 989 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 925 39595 989 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 925 39595 989 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 925 39514 989 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 925 39514 989 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 925 39433 989 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 925 39433 989 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 925 39352 989 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 925 39352 989 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 925 39271 989 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 925 39271 989 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 925 39190 989 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 925 39190 989 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 925 39109 989 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 925 39109 989 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 925 39028 989 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 925 39028 989 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 933 6042 973 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 787 5817 1023 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 787 5817 1023 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 787 5817 1023 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 933 5698 973 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 933 5612 973 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 933 5526 973 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 933 5440 973 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 787 5211 1023 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 787 5211 1023 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 787 5211 1023 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 845 39919 909 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 845 39919 909 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 845 39838 909 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 845 39838 909 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 845 39757 909 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 845 39757 909 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 845 39676 909 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 845 39676 909 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 845 39595 909 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 845 39595 909 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 845 39514 909 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 845 39514 909 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 845 39433 909 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 845 39433 909 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 845 39352 909 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 845 39352 909 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 845 39271 909 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 845 39271 909 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 845 39190 909 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 845 39190 909 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 845 39109 909 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 845 39109 909 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 845 39028 909 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 845 39028 909 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 852 5698 892 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 852 5612 892 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 852 5526 892 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 765 39919 829 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 765 39919 829 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 765 39838 829 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 765 39838 829 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 765 39757 829 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 765 39757 829 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 765 39676 829 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 765 39676 829 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 765 39595 829 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 765 39595 829 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 765 39514 829 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 765 39514 829 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 765 39433 829 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 765 39433 829 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 765 39352 829 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 765 39352 829 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 765 39271 829 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 765 39271 829 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 765 39190 829 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 765 39190 829 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 765 39109 829 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 765 39109 829 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 765 39028 829 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 765 39028 829 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 771 5698 811 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 771 5612 811 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 771 5526 811 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 685 39919 749 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 685 39919 749 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 685 39838 749 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 685 39838 749 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 685 39757 749 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 685 39757 749 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 685 39676 749 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 685 39676 749 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 685 39595 749 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 685 39595 749 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 685 39514 749 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 685 39514 749 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 685 39433 749 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 685 39433 749 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 685 39352 749 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 685 39352 749 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 685 39271 749 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 685 39271 749 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 685 39190 749 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 685 39190 749 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 685 39109 749 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 685 39109 749 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 685 39028 749 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 685 39028 749 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 690 6042 730 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 690 5956 730 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 690 5870 730 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 690 5784 730 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 690 5698 730 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 690 5612 730 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 690 5526 730 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 690 5440 730 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 690 5354 730 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 690 5268 730 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 690 5182 730 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 605 39919 669 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 605 39919 669 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 605 39838 669 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 605 39838 669 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 605 39757 669 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 605 39757 669 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 605 39676 669 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 605 39676 669 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 605 39595 669 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 605 39595 669 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 605 39514 669 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 605 39514 669 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 605 39433 669 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 605 39433 669 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 605 39352 669 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 605 39352 669 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 605 39271 669 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 605 39271 669 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 605 39190 669 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 605 39190 669 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 605 39109 669 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 605 39109 669 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 605 39028 669 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 605 39028 669 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 609 6042 649 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 465 5817 701 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 465 5817 701 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 465 5817 701 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 609 5698 649 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 609 5612 649 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 609 5526 649 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 609 5440 649 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 465 5211 701 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 465 5211 701 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 465 5211 701 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 525 39919 589 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 525 39919 589 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 525 39838 589 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 525 39838 589 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 525 39757 589 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 525 39757 589 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 525 39676 589 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 525 39676 589 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 525 39595 589 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 525 39595 589 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 525 39514 589 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 525 39514 589 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 525 39433 589 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 525 39433 589 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 525 39352 589 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 525 39352 589 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 525 39271 589 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 525 39271 589 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 525 39190 589 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 525 39190 589 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 525 39109 589 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 525 39109 589 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 525 39028 589 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 525 39028 589 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 527 5698 567 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 527 5612 567 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 527 5526 567 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 445 39919 509 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 445 39919 509 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 445 39838 509 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 445 39838 509 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 445 39757 509 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 445 39757 509 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 445 39676 509 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 445 39676 509 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 445 39595 509 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 445 39595 509 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 445 39514 509 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 445 39514 509 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 445 39433 509 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 445 39433 509 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 445 39352 509 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 445 39352 509 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 445 39271 509 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 445 39271 509 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 445 39190 509 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 445 39190 509 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 445 39109 509 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 445 39109 509 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 445 39028 509 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 445 39028 509 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 445 5698 485 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 445 5612 485 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 445 5526 485 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 365 39919 429 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 365 39919 429 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 365 39838 429 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 365 39838 429 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 365 39757 429 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 365 39757 429 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 365 39676 429 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 365 39676 429 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 365 39595 429 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 365 39595 429 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 365 39514 429 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 365 39514 429 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 365 39433 429 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 365 39433 429 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 365 39352 429 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 365 39352 429 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 365 39271 429 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 365 39271 429 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 365 39190 429 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 365 39190 429 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 365 39109 429 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 365 39109 429 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 365 39028 429 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 365 39028 429 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 363 6042 403 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 363 5956 403 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 363 5870 403 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 363 5784 403 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 363 5698 403 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 363 5612 403 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 363 5526 403 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 363 5440 403 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 363 5354 403 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 363 5268 403 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 363 5182 403 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 285 39919 349 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 285 39919 349 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 285 39838 349 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 285 39838 349 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 285 39757 349 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 285 39757 349 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 285 39676 349 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 285 39676 349 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 285 39595 349 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 285 39595 349 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 285 39514 349 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 285 39514 349 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 285 39433 349 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 285 39433 349 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 285 39352 349 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 285 39352 349 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 285 39271 349 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 285 39271 349 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 285 39190 349 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 285 39190 349 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 285 39109 349 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 285 39109 349 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 285 39028 349 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 285 39028 349 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 281 6042 321 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 254 5817 379 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 254 5817 379 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 254 5817 379 6053 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 281 5698 321 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 281 5612 321 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 281 5526 321 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 281 5440 321 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 254 5211 379 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 254 5211 379 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 254 5211 379 5447 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 254 39919 269 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 205 39919 269 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 254 39838 269 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 205 39838 269 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 254 39757 269 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 205 39757 269 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 254 39676 269 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 205 39676 269 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 254 39595 269 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 205 39595 269 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 254 39514 269 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 205 39514 269 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 254 39433 269 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 205 39433 269 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 254 39352 269 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 205 39352 269 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 254 39271 269 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 205 39271 269 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 254 39190 269 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 205 39190 269 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 254 39109 269 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 205 39109 269 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 254 39028 269 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 205 39028 269 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 199 6042 239 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 199 5956 239 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 199 5870 239 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 199 5784 239 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 199 5698 239 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 199 5612 239 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 199 5526 239 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 199 5440 239 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 199 5354 239 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 199 5268 239 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 199 5182 239 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 125 39919 189 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 125 39838 189 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 125 39757 189 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 125 39676 189 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 125 39595 189 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 125 39514 189 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 125 39433 189 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 125 39352 189 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 125 39271 189 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 125 39190 189 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 125 39109 189 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 125 39028 189 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 117 6042 157 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 117 5956 157 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 117 5870 157 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 117 5784 157 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 117 5698 157 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 117 5612 157 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 117 5526 157 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 117 5440 157 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 117 5354 157 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 117 5268 157 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 117 5182 157 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 0 6397 254 7047 6 VSWITCH
port 6 nsew power bidirectional
rlabel metal5 s 14746 6397 15000 7047 6 VSWITCH
port 6 nsew power bidirectional
rlabel metal4 s 0 6377 254 7067 6 VSWITCH
port 6 nsew power bidirectional
rlabel metal4 s 14746 6377 15000 7067 6 VSWITCH
port 6 nsew power bidirectional
rlabel metal5 s 0 11667 254 12517 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal5 s 14746 11667 15000 12517 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 0 11647 254 12537 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14746 11647 15000 12537 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14788 12470 14852 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14788 12388 14852 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14788 12306 14852 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14788 12224 14852 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14788 12142 14852 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14788 12060 14852 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14788 11978 14852 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14788 11896 14852 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14788 11814 14852 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14788 11732 14852 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14788 11650 14852 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14707 12470 14746 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14707 12470 14771 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14707 12388 14746 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14707 12388 14771 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14707 12306 14746 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14707 12306 14771 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14707 12224 14746 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14707 12224 14771 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14707 12142 14746 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14707 12142 14771 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14707 12060 14746 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14707 12060 14771 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14707 11978 14746 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14707 11978 14771 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14707 11896 14746 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14707 11896 14771 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14707 11814 14746 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14707 11814 14771 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14707 11732 14746 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14707 11732 14771 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14707 11650 14746 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14707 11650 14771 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14626 12470 14690 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14626 12470 14690 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14626 12388 14690 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14626 12388 14690 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14626 12306 14690 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14626 12306 14690 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14626 12224 14690 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14626 12224 14690 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14626 12142 14690 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14626 12142 14690 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14626 12060 14690 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14626 12060 14690 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14626 11978 14690 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14626 11978 14690 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14626 11896 14690 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14626 11896 14690 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14626 11814 14690 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14626 11814 14690 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14626 11732 14690 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14626 11732 14690 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14626 11650 14690 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14626 11650 14690 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14545 12470 14609 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14545 12470 14609 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14545 12388 14609 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14545 12388 14609 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14545 12306 14609 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14545 12306 14609 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14545 12224 14609 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14545 12224 14609 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14545 12142 14609 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14545 12142 14609 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14545 12060 14609 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14545 12060 14609 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14545 11978 14609 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14545 11978 14609 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14545 11896 14609 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14545 11896 14609 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14545 11814 14609 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14545 11814 14609 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14545 11732 14609 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14545 11732 14609 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14545 11650 14609 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14545 11650 14609 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14464 12470 14528 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14464 12470 14528 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14464 12388 14528 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14464 12388 14528 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14464 12306 14528 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14464 12306 14528 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14464 12224 14528 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14464 12224 14528 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14464 12142 14528 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14464 12142 14528 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14464 12060 14528 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14464 12060 14528 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14464 11978 14528 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14464 11978 14528 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14464 11896 14528 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14464 11896 14528 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14464 11814 14528 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14464 11814 14528 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14464 11732 14528 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14464 11732 14528 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14464 11650 14528 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14464 11650 14528 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14383 12470 14447 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14383 12470 14447 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14383 12388 14447 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14383 12388 14447 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14383 12306 14447 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14383 12306 14447 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14383 12224 14447 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14383 12224 14447 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14383 12142 14447 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14383 12142 14447 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14383 12060 14447 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14383 12060 14447 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14383 11978 14447 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14383 11978 14447 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14383 11896 14447 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14383 11896 14447 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14383 11814 14447 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14383 11814 14447 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14383 11732 14447 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14383 11732 14447 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14383 11650 14447 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14383 11650 14447 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14302 12470 14366 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14302 12470 14366 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14302 12388 14366 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14302 12388 14366 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14302 12306 14366 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14302 12306 14366 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14302 12224 14366 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14302 12224 14366 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14302 12142 14366 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14302 12142 14366 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14302 12060 14366 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14302 12060 14366 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14302 11978 14366 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14302 11978 14366 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14302 11896 14366 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14302 11896 14366 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14302 11814 14366 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14302 11814 14366 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14302 11732 14366 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14302 11732 14366 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14302 11650 14366 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14302 11650 14366 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14221 12470 14285 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14221 12470 14285 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14221 12388 14285 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14221 12388 14285 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14221 12306 14285 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14221 12306 14285 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14221 12224 14285 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14221 12224 14285 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14221 12142 14285 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14221 12142 14285 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14221 12060 14285 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14221 12060 14285 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14221 11978 14285 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14221 11978 14285 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14221 11896 14285 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14221 11896 14285 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14221 11814 14285 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14221 11814 14285 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14221 11732 14285 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14221 11732 14285 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14221 11650 14285 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14221 11650 14285 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14140 12470 14204 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14140 12470 14204 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14140 12388 14204 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14140 12388 14204 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14140 12306 14204 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14140 12306 14204 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14140 12224 14204 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14140 12224 14204 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14140 12142 14204 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14140 12142 14204 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14140 12060 14204 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14140 12060 14204 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14140 11978 14204 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14140 11978 14204 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14140 11896 14204 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14140 11896 14204 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14140 11814 14204 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14140 11814 14204 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14140 11732 14204 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14140 11732 14204 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14140 11650 14204 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14140 11650 14204 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14059 12470 14123 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14059 12470 14123 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14059 12388 14123 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14059 12388 14123 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14059 12306 14123 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14059 12306 14123 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14059 12224 14123 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14059 12224 14123 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14059 12142 14123 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14059 12142 14123 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14059 12060 14123 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14059 12060 14123 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14059 11978 14123 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14059 11978 14123 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14059 11896 14123 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14059 11896 14123 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14059 11814 14123 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14059 11814 14123 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14059 11732 14123 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14059 11732 14123 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14059 11650 14123 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14059 11650 14123 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13978 12470 14042 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13978 12470 14042 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13978 12388 14042 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13978 12388 14042 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13978 12306 14042 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13978 12306 14042 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13978 12224 14042 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13978 12224 14042 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13978 12142 14042 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13978 12142 14042 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13978 12060 14042 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13978 12060 14042 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13978 11978 14042 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13978 11978 14042 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13978 11896 14042 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13978 11896 14042 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13978 11814 14042 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13978 11814 14042 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13978 11732 14042 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13978 11732 14042 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13978 11650 14042 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13978 11650 14042 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13897 12470 13961 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13897 12470 13961 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13897 12388 13961 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13897 12388 13961 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13897 12306 13961 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13897 12306 13961 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13897 12224 13961 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13897 12224 13961 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13897 12142 13961 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13897 12142 13961 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13897 12060 13961 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13897 12060 13961 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13897 11978 13961 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13897 11978 13961 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13897 11896 13961 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13897 11896 13961 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13897 11814 13961 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13897 11814 13961 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13897 11732 13961 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13897 11732 13961 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13897 11650 13961 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13897 11650 13961 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13816 12470 13880 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13816 12470 13880 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13816 12388 13880 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13816 12388 13880 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13816 12306 13880 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13816 12306 13880 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13816 12224 13880 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13816 12224 13880 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13816 12142 13880 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13816 12142 13880 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13816 12060 13880 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13816 12060 13880 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13816 11978 13880 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13816 11978 13880 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13816 11896 13880 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13816 11896 13880 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13816 11814 13880 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13816 11814 13880 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13816 11732 13880 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13816 11732 13880 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13816 11650 13880 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13816 11650 13880 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13735 12470 13799 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13735 12470 13799 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13735 12388 13799 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13735 12388 13799 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13735 12306 13799 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13735 12306 13799 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13735 12224 13799 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13735 12224 13799 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13735 12142 13799 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13735 12142 13799 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13735 12060 13799 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13735 12060 13799 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13735 11978 13799 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13735 11978 13799 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13735 11896 13799 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13735 11896 13799 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13735 11814 13799 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13735 11814 13799 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13735 11732 13799 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13735 11732 13799 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13735 11650 13799 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13735 11650 13799 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13654 12470 13718 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13654 12470 13718 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13654 12388 13718 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13654 12388 13718 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13654 12306 13718 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13654 12306 13718 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13654 12224 13718 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13654 12224 13718 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13654 12142 13718 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13654 12142 13718 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13654 12060 13718 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13654 12060 13718 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13654 11978 13718 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13654 11978 13718 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13654 11896 13718 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13654 11896 13718 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13654 11814 13718 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13654 11814 13718 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13654 11732 13718 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13654 11732 13718 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13654 11650 13718 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13654 11650 13718 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13573 12470 13637 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13573 12470 13637 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13573 12388 13637 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13573 12388 13637 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13573 12306 13637 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13573 12306 13637 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13573 12224 13637 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13573 12224 13637 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13573 12142 13637 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13573 12142 13637 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13573 12060 13637 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13573 12060 13637 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13573 11978 13637 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13573 11978 13637 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13573 11896 13637 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13573 11896 13637 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13573 11814 13637 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13573 11814 13637 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13573 11732 13637 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13573 11732 13637 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13573 11650 13637 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13573 11650 13637 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13492 12470 13556 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13492 12470 13556 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13492 12388 13556 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13492 12388 13556 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13492 12306 13556 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13492 12306 13556 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13492 12224 13556 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13492 12224 13556 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13492 12142 13556 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13492 12142 13556 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13492 12060 13556 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13492 12060 13556 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13492 11978 13556 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13492 11978 13556 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13492 11896 13556 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13492 11896 13556 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13492 11814 13556 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13492 11814 13556 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13492 11732 13556 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13492 11732 13556 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13492 11650 13556 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13492 11650 13556 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13411 12470 13475 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13411 12470 13475 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13411 12388 13475 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13411 12388 13475 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13411 12306 13475 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13411 12306 13475 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13411 12224 13475 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13411 12224 13475 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13411 12142 13475 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13411 12142 13475 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13411 12060 13475 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13411 12060 13475 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13411 11978 13475 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13411 11978 13475 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13411 11896 13475 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13411 11896 13475 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13411 11814 13475 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13411 11814 13475 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13411 11732 13475 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13411 11732 13475 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13411 11650 13475 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13411 11650 13475 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13330 12470 13394 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13330 12470 13394 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13330 12388 13394 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13330 12388 13394 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13330 12306 13394 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13330 12306 13394 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13330 12224 13394 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13330 12224 13394 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13330 12142 13394 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13330 12142 13394 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13330 12060 13394 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13330 12060 13394 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13330 11978 13394 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13330 11978 13394 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13330 11896 13394 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13330 11896 13394 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13330 11814 13394 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13330 11814 13394 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13330 11732 13394 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13330 11732 13394 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13330 11650 13394 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13330 11650 13394 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13249 12470 13313 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13249 12470 13313 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13249 12388 13313 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13249 12388 13313 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13249 12306 13313 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13249 12306 13313 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13249 12224 13313 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13249 12224 13313 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13249 12142 13313 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13249 12142 13313 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13249 12060 13313 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13249 12060 13313 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13249 11978 13313 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13249 11978 13313 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13249 11896 13313 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13249 11896 13313 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13249 11814 13313 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13249 11814 13313 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13249 11732 13313 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13249 11732 13313 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13249 11650 13313 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13249 11650 13313 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13168 12470 13232 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13168 12470 13232 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13168 12388 13232 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13168 12388 13232 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13168 12306 13232 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13168 12306 13232 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13168 12224 13232 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13168 12224 13232 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13168 12142 13232 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13168 12142 13232 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13168 12060 13232 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13168 12060 13232 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13168 11978 13232 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13168 11978 13232 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13168 11896 13232 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13168 11896 13232 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13168 11814 13232 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13168 11814 13232 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13168 11732 13232 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13168 11732 13232 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13168 11650 13232 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13168 11650 13232 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13087 12470 13151 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13087 12470 13151 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13087 12388 13151 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13087 12388 13151 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13087 12306 13151 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13087 12306 13151 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13087 12224 13151 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13087 12224 13151 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13087 12142 13151 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13087 12142 13151 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13087 12060 13151 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13087 12060 13151 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13087 11978 13151 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13087 11978 13151 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13087 11896 13151 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13087 11896 13151 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13087 11814 13151 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13087 11814 13151 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13087 11732 13151 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13087 11732 13151 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13087 11650 13151 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13087 11650 13151 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13006 12470 13070 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13006 12470 13070 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13006 12388 13070 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13006 12388 13070 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13006 12306 13070 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13006 12306 13070 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13006 12224 13070 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13006 12224 13070 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13006 12142 13070 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13006 12142 13070 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13006 12060 13070 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13006 12060 13070 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13006 11978 13070 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13006 11978 13070 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13006 11896 13070 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13006 11896 13070 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13006 11814 13070 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13006 11814 13070 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13006 11732 13070 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13006 11732 13070 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 13006 11650 13070 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13006 11650 13070 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12925 12470 12989 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12925 12470 12989 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12925 12388 12989 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12925 12388 12989 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12925 12306 12989 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12925 12306 12989 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12925 12224 12989 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12925 12224 12989 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12925 12142 12989 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12925 12142 12989 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12925 12060 12989 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12925 12060 12989 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12925 11978 12989 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12925 11978 12989 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12925 11896 12989 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12925 11896 12989 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12925 11814 12989 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12925 11814 12989 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12925 11732 12989 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12925 11732 12989 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12925 11650 12989 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12925 11650 12989 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12844 12470 12908 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12844 12470 12908 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12844 12388 12908 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12844 12388 12908 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12844 12306 12908 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12844 12306 12908 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12844 12224 12908 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12844 12224 12908 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12844 12142 12908 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12844 12142 12908 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12844 12060 12908 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12844 12060 12908 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12844 11978 12908 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12844 11978 12908 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12844 11896 12908 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12844 11896 12908 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12844 11814 12908 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12844 11814 12908 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12844 11732 12908 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12844 11732 12908 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12844 11650 12908 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12844 11650 12908 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12763 12470 12827 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12763 12470 12827 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12763 12388 12827 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12763 12388 12827 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12763 12306 12827 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12763 12306 12827 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12763 12224 12827 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12763 12224 12827 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12763 12142 12827 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12763 12142 12827 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12763 12060 12827 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12763 12060 12827 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12763 11978 12827 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12763 11978 12827 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12763 11896 12827 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12763 11896 12827 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12763 11814 12827 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12763 11814 12827 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12763 11732 12827 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12763 11732 12827 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12763 11650 12827 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12763 11650 12827 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12682 12470 12746 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12682 12470 12746 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12682 12388 12746 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12682 12388 12746 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12682 12306 12746 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12682 12306 12746 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12682 12224 12746 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12682 12224 12746 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12682 12142 12746 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12682 12142 12746 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12682 12060 12746 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12682 12060 12746 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12682 11978 12746 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12682 11978 12746 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12682 11896 12746 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12682 11896 12746 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12682 11814 12746 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12682 11814 12746 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12682 11732 12746 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12682 11732 12746 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12682 11650 12746 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12682 11650 12746 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12601 12470 12665 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12601 12470 12665 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12601 12388 12665 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12601 12388 12665 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12601 12306 12665 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12601 12306 12665 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12601 12224 12665 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12601 12224 12665 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12601 12142 12665 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12601 12142 12665 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12601 12060 12665 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12601 12060 12665 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12601 11978 12665 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12601 11978 12665 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12601 11896 12665 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12601 11896 12665 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12601 11814 12665 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12601 11814 12665 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12601 11732 12665 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12601 11732 12665 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12601 11650 12665 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12601 11650 12665 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12520 12470 12584 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12520 12470 12584 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12520 12388 12584 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12520 12388 12584 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12520 12306 12584 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12520 12306 12584 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12520 12224 12584 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12520 12224 12584 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12520 12142 12584 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12520 12142 12584 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12520 12060 12584 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12520 12060 12584 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12520 11978 12584 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12520 11978 12584 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12520 11896 12584 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12520 11896 12584 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12520 11814 12584 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12520 11814 12584 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12520 11732 12584 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12520 11732 12584 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12520 11650 12584 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12520 11650 12584 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12439 12470 12503 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12439 12470 12503 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12439 12388 12503 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12439 12388 12503 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12439 12306 12503 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12439 12306 12503 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12439 12224 12503 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12439 12224 12503 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12439 12142 12503 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12439 12142 12503 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12439 12060 12503 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12439 12060 12503 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12439 11978 12503 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12439 11978 12503 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12439 11896 12503 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12439 11896 12503 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12439 11814 12503 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12439 11814 12503 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12439 11732 12503 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12439 11732 12503 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12439 11650 12503 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12439 11650 12503 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12358 12470 12422 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12358 12470 12422 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12358 12388 12422 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12358 12388 12422 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12358 12306 12422 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12358 12306 12422 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12358 12224 12422 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12358 12224 12422 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12358 12142 12422 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12358 12142 12422 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12358 12060 12422 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12358 12060 12422 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12358 11978 12422 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12358 11978 12422 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12358 11896 12422 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12358 11896 12422 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12358 11814 12422 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12358 11814 12422 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12358 11732 12422 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12358 11732 12422 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12358 11650 12422 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12358 11650 12422 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12277 12470 12341 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12277 12470 12341 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12277 12388 12341 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12277 12388 12341 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12277 12306 12341 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12277 12306 12341 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12277 12224 12341 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12277 12224 12341 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12277 12142 12341 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12277 12142 12341 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12277 12060 12341 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12277 12060 12341 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12277 11978 12341 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12277 11978 12341 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12277 11896 12341 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12277 11896 12341 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12277 11814 12341 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12277 11814 12341 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12277 11732 12341 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12277 11732 12341 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12277 11650 12341 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12277 11650 12341 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12196 12470 12260 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12196 12470 12260 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12196 12388 12260 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12196 12388 12260 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12196 12306 12260 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12196 12306 12260 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12196 12224 12260 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12196 12224 12260 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12196 12142 12260 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12196 12142 12260 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12196 12060 12260 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12196 12060 12260 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12196 11978 12260 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12196 11978 12260 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12196 11896 12260 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12196 11896 12260 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12196 11814 12260 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12196 11814 12260 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12196 11732 12260 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12196 11732 12260 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12196 11650 12260 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12196 11650 12260 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12115 12470 12179 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12115 12470 12179 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12115 12388 12179 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12115 12388 12179 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12115 12306 12179 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12115 12306 12179 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12115 12224 12179 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12115 12224 12179 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12115 12142 12179 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12115 12142 12179 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12115 12060 12179 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12115 12060 12179 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12115 11978 12179 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12115 11978 12179 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12115 11896 12179 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12115 11896 12179 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12115 11814 12179 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12115 11814 12179 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12115 11732 12179 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12115 11732 12179 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12115 11650 12179 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12115 11650 12179 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12034 12470 12098 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12034 12470 12098 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12034 12388 12098 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12034 12388 12098 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12034 12306 12098 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12034 12306 12098 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12034 12224 12098 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12034 12224 12098 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12034 12142 12098 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12034 12142 12098 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12034 12060 12098 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12034 12060 12098 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12034 11978 12098 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12034 11978 12098 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12034 11896 12098 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12034 11896 12098 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12034 11814 12098 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12034 11814 12098 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12034 11732 12098 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12034 11732 12098 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 12034 11650 12098 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12034 11650 12098 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11953 12470 12017 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11953 12470 12017 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11953 12388 12017 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11953 12388 12017 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11953 12306 12017 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11953 12306 12017 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11953 12224 12017 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11953 12224 12017 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11953 12142 12017 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11953 12142 12017 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11953 12060 12017 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11953 12060 12017 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11953 11978 12017 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11953 11978 12017 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11953 11896 12017 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11953 11896 12017 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11953 11814 12017 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11953 11814 12017 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11953 11732 12017 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11953 11732 12017 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11953 11650 12017 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11953 11650 12017 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11872 12470 11936 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11872 12470 11936 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11872 12388 11936 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11872 12388 11936 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11872 12306 11936 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11872 12306 11936 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11872 12224 11936 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11872 12224 11936 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11872 12142 11936 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11872 12142 11936 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11872 12060 11936 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11872 12060 11936 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11872 11978 11936 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11872 11978 11936 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11872 11896 11936 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11872 11896 11936 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11872 11814 11936 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11872 11814 11936 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11872 11732 11936 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11872 11732 11936 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11872 11650 11936 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11872 11650 11936 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11791 12470 11855 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11791 12470 11855 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11791 12388 11855 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11791 12388 11855 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11791 12306 11855 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11791 12306 11855 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11791 12224 11855 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11791 12224 11855 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11791 12142 11855 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11791 12142 11855 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11791 12060 11855 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11791 12060 11855 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11791 11978 11855 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11791 11978 11855 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11791 11896 11855 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11791 11896 11855 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11791 11814 11855 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11791 11814 11855 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11791 11732 11855 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11791 11732 11855 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11791 11650 11855 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11791 11650 11855 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11710 12470 11774 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11710 12470 11774 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11710 12388 11774 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11710 12388 11774 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11710 12306 11774 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11710 12306 11774 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11710 12224 11774 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11710 12224 11774 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11710 12142 11774 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11710 12142 11774 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11710 12060 11774 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11710 12060 11774 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11710 11978 11774 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11710 11978 11774 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11710 11896 11774 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11710 11896 11774 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11710 11814 11774 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11710 11814 11774 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11710 11732 11774 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11710 11732 11774 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11710 11650 11774 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11710 11650 11774 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11629 12470 11693 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11629 12470 11693 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11629 12388 11693 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11629 12388 11693 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11629 12306 11693 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11629 12306 11693 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11629 12224 11693 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11629 12224 11693 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11629 12142 11693 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11629 12142 11693 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11629 12060 11693 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11629 12060 11693 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11629 11978 11693 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11629 11978 11693 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11629 11896 11693 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11629 11896 11693 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11629 11814 11693 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11629 11814 11693 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11629 11732 11693 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11629 11732 11693 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11629 11650 11693 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11629 11650 11693 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11548 12470 11612 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11548 12470 11612 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11548 12388 11612 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11548 12388 11612 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11548 12306 11612 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11548 12306 11612 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11548 12224 11612 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11548 12224 11612 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11548 12142 11612 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11548 12142 11612 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11548 12060 11612 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11548 12060 11612 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11548 11978 11612 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11548 11978 11612 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11548 11896 11612 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11548 11896 11612 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11548 11814 11612 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11548 11814 11612 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11548 11732 11612 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11548 11732 11612 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11548 11650 11612 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11548 11650 11612 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11467 12470 11531 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11467 12470 11531 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11467 12388 11531 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11467 12388 11531 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11467 12306 11531 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11467 12306 11531 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11467 12224 11531 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11467 12224 11531 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11467 12142 11531 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11467 12142 11531 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11467 12060 11531 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11467 12060 11531 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11467 11978 11531 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11467 11978 11531 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11467 11896 11531 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11467 11896 11531 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11467 11814 11531 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11467 11814 11531 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11467 11732 11531 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11467 11732 11531 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11467 11650 11531 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11467 11650 11531 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11386 12470 11450 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11386 12470 11450 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11386 12388 11450 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11386 12388 11450 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11386 12306 11450 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11386 12306 11450 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11386 12224 11450 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11386 12224 11450 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11386 12142 11450 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11386 12142 11450 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11386 12060 11450 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11386 12060 11450 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11386 11978 11450 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11386 11978 11450 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11386 11896 11450 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11386 11896 11450 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11386 11814 11450 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11386 11814 11450 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11386 11732 11450 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11386 11732 11450 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11386 11650 11450 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11386 11650 11450 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11305 12470 11369 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11305 12470 11369 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11305 12388 11369 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11305 12388 11369 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11305 12306 11369 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11305 12306 11369 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11305 12224 11369 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11305 12224 11369 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11305 12142 11369 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11305 12142 11369 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11305 12060 11369 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11305 12060 11369 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11305 11978 11369 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11305 11978 11369 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11305 11896 11369 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11305 11896 11369 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11305 11814 11369 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11305 11814 11369 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11305 11732 11369 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11305 11732 11369 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11305 11650 11369 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11305 11650 11369 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11224 12470 11288 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11224 12470 11288 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11224 12388 11288 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11224 12388 11288 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11224 12306 11288 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11224 12306 11288 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11224 12224 11288 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11224 12224 11288 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11224 12142 11288 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11224 12142 11288 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11224 12060 11288 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11224 12060 11288 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11224 11978 11288 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11224 11978 11288 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11224 11896 11288 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11224 11896 11288 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11224 11814 11288 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11224 11814 11288 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11224 11732 11288 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11224 11732 11288 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11224 11650 11288 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11224 11650 11288 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11143 12470 11207 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11143 12470 11207 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11143 12388 11207 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11143 12388 11207 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11143 12306 11207 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11143 12306 11207 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11143 12224 11207 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11143 12224 11207 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11143 12142 11207 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11143 12142 11207 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11143 12060 11207 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11143 12060 11207 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11143 11978 11207 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11143 11978 11207 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11143 11896 11207 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11143 11896 11207 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11143 11814 11207 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11143 11814 11207 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11143 11732 11207 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11143 11732 11207 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11143 11650 11207 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11143 11650 11207 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11062 12470 11126 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11062 12470 11126 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11062 12388 11126 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11062 12388 11126 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11062 12306 11126 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11062 12306 11126 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11062 12224 11126 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11062 12224 11126 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11062 12142 11126 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11062 12142 11126 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11062 12060 11126 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11062 12060 11126 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11062 11978 11126 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11062 11978 11126 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11062 11896 11126 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11062 11896 11126 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11062 11814 11126 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11062 11814 11126 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11062 11732 11126 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11062 11732 11126 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 11062 11650 11126 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11062 11650 11126 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10981 12470 11045 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10981 12470 11045 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10981 12388 11045 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10981 12388 11045 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10981 12306 11045 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10981 12306 11045 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10981 12224 11045 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10981 12224 11045 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10981 12142 11045 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10981 12142 11045 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10981 12060 11045 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10981 12060 11045 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10981 11978 11045 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10981 11978 11045 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10981 11896 11045 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10981 11896 11045 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10981 11814 11045 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10981 11814 11045 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10981 11732 11045 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10981 11732 11045 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10981 11650 11045 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10981 11650 11045 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10900 12470 10964 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10900 12470 10964 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10900 12388 10964 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10900 12388 10964 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10900 12306 10964 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10900 12306 10964 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10900 12224 10964 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10900 12224 10964 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10900 12142 10964 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10900 12142 10964 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10900 12060 10964 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10900 12060 10964 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10900 11978 10964 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10900 11978 10964 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10900 11896 10964 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10900 11896 10964 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10900 11814 10964 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10900 11814 10964 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10900 11732 10964 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10900 11732 10964 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10900 11650 10964 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10900 11650 10964 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10819 12470 10883 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10819 12470 10883 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10819 12388 10883 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10819 12388 10883 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10819 12306 10883 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10819 12306 10883 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10819 12224 10883 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10819 12224 10883 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10819 12142 10883 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10819 12142 10883 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10819 12060 10883 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10819 12060 10883 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10819 11978 10883 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10819 11978 10883 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10819 11896 10883 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10819 11896 10883 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10819 11814 10883 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10819 11814 10883 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10819 11732 10883 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10819 11732 10883 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10819 11650 10883 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10819 11650 10883 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10738 12470 10802 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10738 12470 10802 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10738 12388 10802 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10738 12388 10802 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10738 12306 10802 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10738 12306 10802 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10738 12224 10802 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10738 12224 10802 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10738 12142 10802 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10738 12142 10802 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10738 12060 10802 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10738 12060 10802 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10738 11978 10802 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10738 11978 10802 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10738 11896 10802 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10738 11896 10802 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10738 11814 10802 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10738 11814 10802 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10738 11732 10802 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10738 11732 10802 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10738 11650 10802 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10738 11650 10802 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10657 12470 10721 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10657 12470 10721 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10657 12388 10721 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10657 12388 10721 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10657 12306 10721 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10657 12306 10721 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10657 12224 10721 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10657 12224 10721 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10657 12142 10721 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10657 12142 10721 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10657 12060 10721 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10657 12060 10721 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10657 11978 10721 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10657 11978 10721 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10657 11896 10721 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10657 11896 10721 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10657 11814 10721 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10657 11814 10721 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10657 11732 10721 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10657 11732 10721 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10657 11650 10721 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10657 11650 10721 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10576 12470 10640 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10576 12470 10640 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10576 12388 10640 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10576 12388 10640 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10576 12306 10640 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10576 12306 10640 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10576 12224 10640 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10576 12224 10640 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10576 12142 10640 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10576 12142 10640 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10576 12060 10640 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10576 12060 10640 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10576 11978 10640 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10576 11978 10640 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10576 11896 10640 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10576 11896 10640 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10576 11814 10640 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10576 11814 10640 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10576 11732 10640 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10576 11732 10640 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10576 11650 10640 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10576 11650 10640 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10494 12470 10558 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10494 12470 10558 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10494 12388 10558 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10494 12388 10558 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10494 12306 10558 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10494 12306 10558 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10494 12224 10558 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10494 12224 10558 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10494 12142 10558 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10494 12142 10558 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10494 12060 10558 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10494 12060 10558 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10494 11978 10558 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10494 11978 10558 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10494 11896 10558 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10494 11896 10558 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10494 11814 10558 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10494 11814 10558 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10494 11732 10558 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10494 11732 10558 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10494 11650 10558 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10494 11650 10558 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10412 12470 10476 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10412 12470 10476 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10412 12388 10476 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10412 12388 10476 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10412 12306 10476 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10412 12306 10476 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10412 12224 10476 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10412 12224 10476 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10412 12142 10476 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10412 12142 10476 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10412 12060 10476 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10412 12060 10476 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10412 11978 10476 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10412 11978 10476 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10412 11896 10476 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10412 11896 10476 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10412 11814 10476 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10412 11814 10476 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10412 11732 10476 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10412 11732 10476 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10412 11650 10476 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10412 11650 10476 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10330 12470 10394 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10330 12470 10394 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10330 12388 10394 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10330 12388 10394 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10330 12306 10394 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10330 12306 10394 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10330 12224 10394 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10330 12224 10394 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10330 12142 10394 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10330 12142 10394 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10330 12060 10394 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10330 12060 10394 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10330 11978 10394 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10330 11978 10394 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10330 11896 10394 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10330 11896 10394 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10330 11814 10394 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10330 11814 10394 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10330 11732 10394 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10330 11732 10394 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10330 11650 10394 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10330 11650 10394 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10248 12470 10312 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10248 12470 10312 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10248 12388 10312 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10248 12388 10312 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10248 12306 10312 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10248 12306 10312 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10248 12224 10312 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10248 12224 10312 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10248 12142 10312 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10248 12142 10312 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10248 12060 10312 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10248 12060 10312 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10248 11978 10312 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10248 11978 10312 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10248 11896 10312 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10248 11896 10312 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10248 11814 10312 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10248 11814 10312 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10248 11732 10312 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10248 11732 10312 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10248 11650 10312 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10248 11650 10312 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10166 12470 10230 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10166 12470 10230 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10166 12388 10230 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10166 12388 10230 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10166 12306 10230 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10166 12306 10230 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10166 12224 10230 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10166 12224 10230 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10166 12142 10230 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10166 12142 10230 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10166 12060 10230 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10166 12060 10230 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10166 11978 10230 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10166 11978 10230 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10166 11896 10230 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10166 11896 10230 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10166 11814 10230 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10166 11814 10230 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10166 11732 10230 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10166 11732 10230 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10166 11650 10230 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10166 11650 10230 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10084 12470 10148 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10084 12470 10148 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10084 12388 10148 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10084 12388 10148 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10084 12306 10148 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10084 12306 10148 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10084 12224 10148 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10084 12224 10148 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10084 12142 10148 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10084 12142 10148 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10084 12060 10148 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10084 12060 10148 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10084 11978 10148 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10084 11978 10148 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10084 11896 10148 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10084 11896 10148 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10084 11814 10148 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10084 11814 10148 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10084 11732 10148 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10084 11732 10148 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10084 11650 10148 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10084 11650 10148 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4809 12470 4873 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4809 12470 4873 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4809 12388 4873 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4809 12388 4873 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4809 12306 4873 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4809 12306 4873 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4809 12224 4873 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4809 12224 4873 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4809 12142 4873 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4809 12142 4873 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4809 12060 4873 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4809 12060 4873 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4809 11978 4873 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4809 11978 4873 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4809 11896 4873 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4809 11896 4873 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4809 11814 4873 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4809 11814 4873 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4809 11732 4873 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4809 11732 4873 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4809 11650 4873 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4809 11650 4873 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4728 12470 4792 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4728 12470 4792 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4728 12388 4792 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4728 12388 4792 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4728 12306 4792 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4728 12306 4792 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4728 12224 4792 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4728 12224 4792 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4728 12142 4792 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4728 12142 4792 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4728 12060 4792 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4728 12060 4792 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4728 11978 4792 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4728 11978 4792 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4728 11896 4792 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4728 11896 4792 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4728 11814 4792 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4728 11814 4792 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4728 11732 4792 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4728 11732 4792 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4728 11650 4792 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4728 11650 4792 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4647 12470 4711 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4647 12470 4711 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4647 12388 4711 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4647 12388 4711 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4647 12306 4711 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4647 12306 4711 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4647 12224 4711 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4647 12224 4711 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4647 12142 4711 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4647 12142 4711 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4647 12060 4711 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4647 12060 4711 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4647 11978 4711 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4647 11978 4711 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4647 11896 4711 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4647 11896 4711 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4647 11814 4711 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4647 11814 4711 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4647 11732 4711 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4647 11732 4711 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4647 11650 4711 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4647 11650 4711 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4566 12470 4630 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4566 12470 4630 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4566 12388 4630 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4566 12388 4630 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4566 12306 4630 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4566 12306 4630 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4566 12224 4630 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4566 12224 4630 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4566 12142 4630 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4566 12142 4630 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4566 12060 4630 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4566 12060 4630 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4566 11978 4630 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4566 11978 4630 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4566 11896 4630 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4566 11896 4630 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4566 11814 4630 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4566 11814 4630 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4566 11732 4630 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4566 11732 4630 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4566 11650 4630 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4566 11650 4630 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4485 12470 4549 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4485 12470 4549 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4485 12388 4549 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4485 12388 4549 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4485 12306 4549 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4485 12306 4549 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4485 12224 4549 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4485 12224 4549 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4485 12142 4549 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4485 12142 4549 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4485 12060 4549 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4485 12060 4549 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4485 11978 4549 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4485 11978 4549 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4485 11896 4549 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4485 11896 4549 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4485 11814 4549 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4485 11814 4549 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4485 11732 4549 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4485 11732 4549 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4485 11650 4549 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4485 11650 4549 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4404 12470 4468 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4404 12470 4468 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4404 12388 4468 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4404 12388 4468 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4404 12306 4468 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4404 12306 4468 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4404 12224 4468 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4404 12224 4468 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4404 12142 4468 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4404 12142 4468 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4404 12060 4468 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4404 12060 4468 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4404 11978 4468 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4404 11978 4468 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4404 11896 4468 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4404 11896 4468 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4404 11814 4468 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4404 11814 4468 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4404 11732 4468 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4404 11732 4468 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4404 11650 4468 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4404 11650 4468 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4323 12470 4387 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4323 12470 4387 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4323 12388 4387 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4323 12388 4387 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4323 12306 4387 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4323 12306 4387 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4323 12224 4387 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4323 12224 4387 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4323 12142 4387 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4323 12142 4387 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4323 12060 4387 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4323 12060 4387 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4323 11978 4387 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4323 11978 4387 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4323 11896 4387 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4323 11896 4387 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4323 11814 4387 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4323 11814 4387 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4323 11732 4387 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4323 11732 4387 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4323 11650 4387 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4323 11650 4387 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4242 12470 4306 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4242 12470 4306 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4242 12388 4306 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4242 12388 4306 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4242 12306 4306 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4242 12306 4306 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4242 12224 4306 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4242 12224 4306 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4242 12142 4306 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4242 12142 4306 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4242 12060 4306 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4242 12060 4306 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4242 11978 4306 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4242 11978 4306 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4242 11896 4306 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4242 11896 4306 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4242 11814 4306 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4242 11814 4306 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4242 11732 4306 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4242 11732 4306 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4242 11650 4306 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4242 11650 4306 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4161 12470 4225 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4161 12470 4225 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4161 12388 4225 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4161 12388 4225 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4161 12306 4225 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4161 12306 4225 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4161 12224 4225 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4161 12224 4225 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4161 12142 4225 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4161 12142 4225 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4161 12060 4225 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4161 12060 4225 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4161 11978 4225 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4161 11978 4225 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4161 11896 4225 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4161 11896 4225 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4161 11814 4225 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4161 11814 4225 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4161 11732 4225 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4161 11732 4225 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4161 11650 4225 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4161 11650 4225 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4080 12470 4144 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4080 12470 4144 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4080 12388 4144 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4080 12388 4144 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4080 12306 4144 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4080 12306 4144 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4080 12224 4144 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4080 12224 4144 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4080 12142 4144 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4080 12142 4144 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4080 12060 4144 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4080 12060 4144 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4080 11978 4144 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4080 11978 4144 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4080 11896 4144 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4080 11896 4144 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4080 11814 4144 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4080 11814 4144 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4080 11732 4144 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4080 11732 4144 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 4080 11650 4144 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4080 11650 4144 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3999 12470 4063 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3999 12470 4063 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3999 12388 4063 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3999 12388 4063 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3999 12306 4063 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3999 12306 4063 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3999 12224 4063 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3999 12224 4063 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3999 12142 4063 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3999 12142 4063 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3999 12060 4063 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3999 12060 4063 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3999 11978 4063 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3999 11978 4063 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3999 11896 4063 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3999 11896 4063 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3999 11814 4063 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3999 11814 4063 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3999 11732 4063 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3999 11732 4063 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3999 11650 4063 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3999 11650 4063 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3918 12470 3982 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3918 12470 3982 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3918 12388 3982 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3918 12388 3982 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3918 12306 3982 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3918 12306 3982 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3918 12224 3982 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3918 12224 3982 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3918 12142 3982 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3918 12142 3982 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3918 12060 3982 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3918 12060 3982 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3918 11978 3982 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3918 11978 3982 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3918 11896 3982 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3918 11896 3982 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3918 11814 3982 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3918 11814 3982 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3918 11732 3982 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3918 11732 3982 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3918 11650 3982 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3918 11650 3982 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3837 12470 3901 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3837 12470 3901 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3837 12388 3901 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3837 12388 3901 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3837 12306 3901 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3837 12306 3901 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3837 12224 3901 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3837 12224 3901 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3837 12142 3901 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3837 12142 3901 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3837 12060 3901 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3837 12060 3901 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3837 11978 3901 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3837 11978 3901 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3837 11896 3901 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3837 11896 3901 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3837 11814 3901 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3837 11814 3901 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3837 11732 3901 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3837 11732 3901 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3837 11650 3901 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3837 11650 3901 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3756 12470 3820 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3756 12470 3820 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3756 12388 3820 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3756 12388 3820 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3756 12306 3820 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3756 12306 3820 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3756 12224 3820 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3756 12224 3820 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3756 12142 3820 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3756 12142 3820 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3756 12060 3820 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3756 12060 3820 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3756 11978 3820 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3756 11978 3820 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3756 11896 3820 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3756 11896 3820 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3756 11814 3820 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3756 11814 3820 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3756 11732 3820 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3756 11732 3820 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3756 11650 3820 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3756 11650 3820 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3675 12470 3739 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3675 12470 3739 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3675 12388 3739 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3675 12388 3739 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3675 12306 3739 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3675 12306 3739 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3675 12224 3739 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3675 12224 3739 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3675 12142 3739 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3675 12142 3739 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3675 12060 3739 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3675 12060 3739 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3675 11978 3739 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3675 11978 3739 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3675 11896 3739 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3675 11896 3739 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3675 11814 3739 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3675 11814 3739 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3675 11732 3739 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3675 11732 3739 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3675 11650 3739 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3675 11650 3739 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3594 12470 3658 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3594 12470 3658 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3594 12388 3658 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3594 12388 3658 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3594 12306 3658 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3594 12306 3658 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3594 12224 3658 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3594 12224 3658 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3594 12142 3658 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3594 12142 3658 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3594 12060 3658 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3594 12060 3658 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3594 11978 3658 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3594 11978 3658 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3594 11896 3658 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3594 11896 3658 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3594 11814 3658 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3594 11814 3658 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3594 11732 3658 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3594 11732 3658 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3594 11650 3658 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3594 11650 3658 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3513 12470 3577 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3513 12470 3577 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3513 12388 3577 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3513 12388 3577 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3513 12306 3577 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3513 12306 3577 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3513 12224 3577 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3513 12224 3577 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3513 12142 3577 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3513 12142 3577 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3513 12060 3577 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3513 12060 3577 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3513 11978 3577 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3513 11978 3577 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3513 11896 3577 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3513 11896 3577 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3513 11814 3577 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3513 11814 3577 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3513 11732 3577 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3513 11732 3577 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3513 11650 3577 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3513 11650 3577 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3432 12470 3496 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3432 12470 3496 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3432 12388 3496 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3432 12388 3496 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3432 12306 3496 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3432 12306 3496 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3432 12224 3496 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3432 12224 3496 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3432 12142 3496 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3432 12142 3496 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3432 12060 3496 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3432 12060 3496 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3432 11978 3496 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3432 11978 3496 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3432 11896 3496 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3432 11896 3496 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3432 11814 3496 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3432 11814 3496 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3432 11732 3496 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3432 11732 3496 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3432 11650 3496 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3432 11650 3496 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3351 12470 3415 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3351 12470 3415 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3351 12388 3415 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3351 12388 3415 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3351 12306 3415 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3351 12306 3415 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3351 12224 3415 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3351 12224 3415 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3351 12142 3415 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3351 12142 3415 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3351 12060 3415 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3351 12060 3415 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3351 11978 3415 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3351 11978 3415 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3351 11896 3415 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3351 11896 3415 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3351 11814 3415 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3351 11814 3415 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3351 11732 3415 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3351 11732 3415 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3351 11650 3415 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3351 11650 3415 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3270 12470 3334 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3270 12470 3334 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3270 12388 3334 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3270 12388 3334 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3270 12306 3334 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3270 12306 3334 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3270 12224 3334 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3270 12224 3334 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3270 12142 3334 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3270 12142 3334 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3270 12060 3334 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3270 12060 3334 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3270 11978 3334 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3270 11978 3334 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3270 11896 3334 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3270 11896 3334 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3270 11814 3334 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3270 11814 3334 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3270 11732 3334 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3270 11732 3334 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3270 11650 3334 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3270 11650 3334 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3189 12470 3253 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3189 12470 3253 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3189 12388 3253 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3189 12388 3253 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3189 12306 3253 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3189 12306 3253 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3189 12224 3253 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3189 12224 3253 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3189 12142 3253 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3189 12142 3253 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3189 12060 3253 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3189 12060 3253 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3189 11978 3253 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3189 11978 3253 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3189 11896 3253 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3189 11896 3253 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3189 11814 3253 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3189 11814 3253 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3189 11732 3253 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3189 11732 3253 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3189 11650 3253 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3189 11650 3253 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3108 12470 3172 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3108 12470 3172 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3108 12388 3172 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3108 12388 3172 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3108 12306 3172 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3108 12306 3172 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3108 12224 3172 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3108 12224 3172 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3108 12142 3172 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3108 12142 3172 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3108 12060 3172 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3108 12060 3172 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3108 11978 3172 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3108 11978 3172 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3108 11896 3172 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3108 11896 3172 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3108 11814 3172 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3108 11814 3172 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3108 11732 3172 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3108 11732 3172 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3108 11650 3172 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3108 11650 3172 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3027 12470 3091 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3027 12470 3091 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3027 12388 3091 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3027 12388 3091 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3027 12306 3091 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3027 12306 3091 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3027 12224 3091 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3027 12224 3091 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3027 12142 3091 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3027 12142 3091 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3027 12060 3091 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3027 12060 3091 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3027 11978 3091 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3027 11978 3091 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3027 11896 3091 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3027 11896 3091 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3027 11814 3091 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3027 11814 3091 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3027 11732 3091 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3027 11732 3091 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 3027 11650 3091 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3027 11650 3091 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2946 12470 3010 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2946 12470 3010 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2946 12388 3010 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2946 12388 3010 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2946 12306 3010 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2946 12306 3010 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2946 12224 3010 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2946 12224 3010 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2946 12142 3010 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2946 12142 3010 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2946 12060 3010 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2946 12060 3010 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2946 11978 3010 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2946 11978 3010 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2946 11896 3010 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2946 11896 3010 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2946 11814 3010 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2946 11814 3010 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2946 11732 3010 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2946 11732 3010 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2946 11650 3010 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2946 11650 3010 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2865 12470 2929 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2865 12470 2929 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2865 12388 2929 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2865 12388 2929 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2865 12306 2929 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2865 12306 2929 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2865 12224 2929 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2865 12224 2929 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2865 12142 2929 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2865 12142 2929 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2865 12060 2929 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2865 12060 2929 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2865 11978 2929 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2865 11978 2929 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2865 11896 2929 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2865 11896 2929 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2865 11814 2929 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2865 11814 2929 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2865 11732 2929 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2865 11732 2929 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2865 11650 2929 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2865 11650 2929 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2784 12470 2848 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2784 12470 2848 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2784 12388 2848 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2784 12388 2848 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2784 12306 2848 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2784 12306 2848 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2784 12224 2848 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2784 12224 2848 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2784 12142 2848 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2784 12142 2848 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2784 12060 2848 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2784 12060 2848 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2784 11978 2848 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2784 11978 2848 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2784 11896 2848 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2784 11896 2848 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2784 11814 2848 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2784 11814 2848 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2784 11732 2848 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2784 11732 2848 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2784 11650 2848 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2784 11650 2848 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2703 12470 2767 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2703 12470 2767 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2703 12388 2767 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2703 12388 2767 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2703 12306 2767 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2703 12306 2767 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2703 12224 2767 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2703 12224 2767 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2703 12142 2767 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2703 12142 2767 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2703 12060 2767 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2703 12060 2767 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2703 11978 2767 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2703 11978 2767 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2703 11896 2767 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2703 11896 2767 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2703 11814 2767 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2703 11814 2767 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2703 11732 2767 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2703 11732 2767 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2703 11650 2767 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2703 11650 2767 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2622 12470 2686 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2622 12470 2686 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2622 12388 2686 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2622 12388 2686 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2622 12306 2686 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2622 12306 2686 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2622 12224 2686 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2622 12224 2686 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2622 12142 2686 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2622 12142 2686 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2622 12060 2686 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2622 12060 2686 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2622 11978 2686 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2622 11978 2686 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2622 11896 2686 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2622 11896 2686 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2622 11814 2686 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2622 11814 2686 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2622 11732 2686 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2622 11732 2686 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2622 11650 2686 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2622 11650 2686 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2541 12470 2605 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2541 12470 2605 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2541 12388 2605 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2541 12388 2605 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2541 12306 2605 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2541 12306 2605 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2541 12224 2605 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2541 12224 2605 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2541 12142 2605 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2541 12142 2605 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2541 12060 2605 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2541 12060 2605 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2541 11978 2605 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2541 11978 2605 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2541 11896 2605 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2541 11896 2605 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2541 11814 2605 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2541 11814 2605 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2541 11732 2605 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2541 11732 2605 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2541 11650 2605 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2541 11650 2605 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2460 12470 2524 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2460 12470 2524 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2460 12388 2524 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2460 12388 2524 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2460 12306 2524 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2460 12306 2524 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2460 12224 2524 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2460 12224 2524 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2460 12142 2524 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2460 12142 2524 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2460 12060 2524 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2460 12060 2524 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2460 11978 2524 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2460 11978 2524 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2460 11896 2524 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2460 11896 2524 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2460 11814 2524 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2460 11814 2524 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2460 11732 2524 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2460 11732 2524 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2460 11650 2524 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2460 11650 2524 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2379 12470 2443 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2379 12470 2443 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2379 12388 2443 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2379 12388 2443 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2379 12306 2443 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2379 12306 2443 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2379 12224 2443 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2379 12224 2443 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2379 12142 2443 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2379 12142 2443 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2379 12060 2443 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2379 12060 2443 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2379 11978 2443 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2379 11978 2443 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2379 11896 2443 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2379 11896 2443 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2379 11814 2443 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2379 11814 2443 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2379 11732 2443 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2379 11732 2443 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2379 11650 2443 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2379 11650 2443 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2298 12470 2362 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2298 12470 2362 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2298 12388 2362 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2298 12388 2362 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2298 12306 2362 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2298 12306 2362 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2298 12224 2362 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2298 12224 2362 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2298 12142 2362 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2298 12142 2362 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2298 12060 2362 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2298 12060 2362 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2298 11978 2362 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2298 11978 2362 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2298 11896 2362 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2298 11896 2362 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2298 11814 2362 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2298 11814 2362 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2298 11732 2362 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2298 11732 2362 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2298 11650 2362 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2298 11650 2362 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2217 12470 2281 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2217 12470 2281 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2217 12388 2281 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2217 12388 2281 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2217 12306 2281 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2217 12306 2281 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2217 12224 2281 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2217 12224 2281 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2217 12142 2281 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2217 12142 2281 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2217 12060 2281 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2217 12060 2281 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2217 11978 2281 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2217 11978 2281 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2217 11896 2281 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2217 11896 2281 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2217 11814 2281 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2217 11814 2281 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2217 11732 2281 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2217 11732 2281 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2217 11650 2281 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2217 11650 2281 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2136 12470 2200 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2136 12470 2200 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2136 12388 2200 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2136 12388 2200 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2136 12306 2200 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2136 12306 2200 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2136 12224 2200 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2136 12224 2200 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2136 12142 2200 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2136 12142 2200 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2136 12060 2200 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2136 12060 2200 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2136 11978 2200 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2136 11978 2200 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2136 11896 2200 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2136 11896 2200 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2136 11814 2200 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2136 11814 2200 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2136 11732 2200 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2136 11732 2200 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2136 11650 2200 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2136 11650 2200 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2055 12470 2119 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2055 12470 2119 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2055 12388 2119 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2055 12388 2119 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2055 12306 2119 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2055 12306 2119 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2055 12224 2119 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2055 12224 2119 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2055 12142 2119 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2055 12142 2119 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2055 12060 2119 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2055 12060 2119 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2055 11978 2119 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2055 11978 2119 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2055 11896 2119 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2055 11896 2119 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2055 11814 2119 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2055 11814 2119 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2055 11732 2119 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2055 11732 2119 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 2055 11650 2119 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2055 11650 2119 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1974 12470 2038 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1974 12470 2038 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1974 12388 2038 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1974 12388 2038 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1974 12306 2038 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1974 12306 2038 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1974 12224 2038 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1974 12224 2038 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1974 12142 2038 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1974 12142 2038 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1974 12060 2038 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1974 12060 2038 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1974 11978 2038 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1974 11978 2038 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1974 11896 2038 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1974 11896 2038 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1974 11814 2038 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1974 11814 2038 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1974 11732 2038 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1974 11732 2038 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1974 11650 2038 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1974 11650 2038 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1893 12470 1957 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1893 12470 1957 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1893 12388 1957 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1893 12388 1957 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1893 12306 1957 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1893 12306 1957 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1893 12224 1957 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1893 12224 1957 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1893 12142 1957 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1893 12142 1957 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1893 12060 1957 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1893 12060 1957 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1893 11978 1957 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1893 11978 1957 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1893 11896 1957 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1893 11896 1957 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1893 11814 1957 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1893 11814 1957 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1893 11732 1957 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1893 11732 1957 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1893 11650 1957 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1893 11650 1957 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1812 12470 1876 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1812 12470 1876 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1812 12388 1876 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1812 12388 1876 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1812 12306 1876 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1812 12306 1876 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1812 12224 1876 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1812 12224 1876 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1812 12142 1876 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1812 12142 1876 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1812 12060 1876 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1812 12060 1876 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1812 11978 1876 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1812 11978 1876 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1812 11896 1876 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1812 11896 1876 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1812 11814 1876 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1812 11814 1876 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1812 11732 1876 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1812 11732 1876 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1812 11650 1876 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1812 11650 1876 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1731 12470 1795 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1731 12470 1795 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1731 12388 1795 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1731 12388 1795 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1731 12306 1795 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1731 12306 1795 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1731 12224 1795 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1731 12224 1795 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1731 12142 1795 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1731 12142 1795 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1731 12060 1795 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1731 12060 1795 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1731 11978 1795 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1731 11978 1795 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1731 11896 1795 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1731 11896 1795 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1731 11814 1795 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1731 11814 1795 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1731 11732 1795 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1731 11732 1795 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1731 11650 1795 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1731 11650 1795 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1650 12470 1714 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1650 12470 1714 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1650 12388 1714 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1650 12388 1714 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1650 12306 1714 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1650 12306 1714 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1650 12224 1714 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1650 12224 1714 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1650 12142 1714 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1650 12142 1714 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1650 12060 1714 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1650 12060 1714 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1650 11978 1714 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1650 11978 1714 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1650 11896 1714 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1650 11896 1714 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1650 11814 1714 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1650 11814 1714 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1650 11732 1714 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1650 11732 1714 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1650 11650 1714 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1650 11650 1714 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1569 12470 1633 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1569 12470 1633 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1569 12388 1633 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1569 12388 1633 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1569 12306 1633 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1569 12306 1633 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1569 12224 1633 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1569 12224 1633 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1569 12142 1633 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1569 12142 1633 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1569 12060 1633 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1569 12060 1633 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1569 11978 1633 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1569 11978 1633 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1569 11896 1633 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1569 11896 1633 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1569 11814 1633 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1569 11814 1633 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1569 11732 1633 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1569 11732 1633 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1569 11650 1633 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1569 11650 1633 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1488 12470 1552 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1488 12470 1552 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1488 12388 1552 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1488 12388 1552 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1488 12306 1552 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1488 12306 1552 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1488 12224 1552 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1488 12224 1552 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1488 12142 1552 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1488 12142 1552 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1488 12060 1552 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1488 12060 1552 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1488 11978 1552 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1488 11978 1552 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1488 11896 1552 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1488 11896 1552 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1488 11814 1552 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1488 11814 1552 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1488 11732 1552 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1488 11732 1552 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1488 11650 1552 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1488 11650 1552 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1407 12470 1471 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1407 12470 1471 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1407 12388 1471 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1407 12388 1471 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1407 12306 1471 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1407 12306 1471 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1407 12224 1471 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1407 12224 1471 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1407 12142 1471 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1407 12142 1471 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1407 12060 1471 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1407 12060 1471 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1407 11978 1471 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1407 11978 1471 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1407 11896 1471 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1407 11896 1471 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1407 11814 1471 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1407 11814 1471 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1407 11732 1471 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1407 11732 1471 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1407 11650 1471 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1407 11650 1471 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1326 12470 1390 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1326 12470 1390 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1326 12388 1390 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1326 12388 1390 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1326 12306 1390 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1326 12306 1390 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1326 12224 1390 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1326 12224 1390 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1326 12142 1390 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1326 12142 1390 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1326 12060 1390 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1326 12060 1390 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1326 11978 1390 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1326 11978 1390 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1326 11896 1390 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1326 11896 1390 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1326 11814 1390 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1326 11814 1390 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1326 11732 1390 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1326 11732 1390 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1326 11650 1390 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1326 11650 1390 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1245 12470 1309 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1245 12470 1309 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1245 12388 1309 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1245 12388 1309 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1245 12306 1309 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1245 12306 1309 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1245 12224 1309 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1245 12224 1309 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1245 12142 1309 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1245 12142 1309 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1245 12060 1309 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1245 12060 1309 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1245 11978 1309 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1245 11978 1309 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1245 11896 1309 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1245 11896 1309 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1245 11814 1309 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1245 11814 1309 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1245 11732 1309 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1245 11732 1309 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1245 11650 1309 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1245 11650 1309 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1164 12470 1228 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1164 12470 1228 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1164 12388 1228 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1164 12388 1228 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1164 12306 1228 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1164 12306 1228 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1164 12224 1228 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1164 12224 1228 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1164 12142 1228 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1164 12142 1228 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1164 12060 1228 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1164 12060 1228 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1164 11978 1228 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1164 11978 1228 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1164 11896 1228 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1164 11896 1228 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1164 11814 1228 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1164 11814 1228 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1164 11732 1228 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1164 11732 1228 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1164 11650 1228 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1164 11650 1228 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1083 12470 1147 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1083 12470 1147 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1083 12388 1147 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1083 12388 1147 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1083 12306 1147 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1083 12306 1147 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1083 12224 1147 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1083 12224 1147 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1083 12142 1147 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1083 12142 1147 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1083 12060 1147 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1083 12060 1147 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1083 11978 1147 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1083 11978 1147 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1083 11896 1147 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1083 11896 1147 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1083 11814 1147 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1083 11814 1147 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1083 11732 1147 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1083 11732 1147 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1083 11650 1147 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1083 11650 1147 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1002 12470 1066 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1002 12470 1066 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1002 12388 1066 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1002 12388 1066 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1002 12306 1066 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1002 12306 1066 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1002 12224 1066 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1002 12224 1066 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1002 12142 1066 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1002 12142 1066 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1002 12060 1066 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1002 12060 1066 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1002 11978 1066 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1002 11978 1066 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1002 11896 1066 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1002 11896 1066 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1002 11814 1066 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1002 11814 1066 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1002 11732 1066 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1002 11732 1066 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 1002 11650 1066 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1002 11650 1066 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 921 12470 985 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 921 12470 985 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 921 12388 985 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 921 12388 985 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 921 12306 985 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 921 12306 985 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 921 12224 985 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 921 12224 985 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 921 12142 985 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 921 12142 985 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 921 12060 985 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 921 12060 985 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 921 11978 985 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 921 11978 985 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 921 11896 985 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 921 11896 985 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 921 11814 985 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 921 11814 985 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 921 11732 985 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 921 11732 985 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 921 11650 985 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 921 11650 985 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 840 12470 904 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 840 12470 904 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 840 12388 904 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 840 12388 904 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 840 12306 904 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 840 12306 904 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 840 12224 904 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 840 12224 904 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 840 12142 904 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 840 12142 904 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 840 12060 904 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 840 12060 904 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 840 11978 904 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 840 11978 904 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 840 11896 904 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 840 11896 904 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 840 11814 904 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 840 11814 904 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 840 11732 904 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 840 11732 904 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 840 11650 904 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 840 11650 904 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 759 12470 823 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 759 12470 823 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 759 12388 823 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 759 12388 823 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 759 12306 823 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 759 12306 823 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 759 12224 823 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 759 12224 823 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 759 12142 823 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 759 12142 823 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 759 12060 823 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 759 12060 823 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 759 11978 823 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 759 11978 823 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 759 11896 823 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 759 11896 823 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 759 11814 823 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 759 11814 823 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 759 11732 823 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 759 11732 823 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 759 11650 823 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 759 11650 823 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 678 12470 742 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 678 12470 742 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 678 12388 742 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 678 12388 742 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 678 12306 742 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 678 12306 742 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 678 12224 742 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 678 12224 742 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 678 12142 742 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 678 12142 742 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 678 12060 742 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 678 12060 742 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 678 11978 742 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 678 11978 742 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 678 11896 742 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 678 11896 742 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 678 11814 742 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 678 11814 742 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 678 11732 742 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 678 11732 742 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 678 11650 742 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 678 11650 742 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 597 12470 661 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 597 12470 661 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 597 12388 661 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 597 12388 661 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 597 12306 661 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 597 12306 661 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 597 12224 661 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 597 12224 661 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 597 12142 661 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 597 12142 661 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 597 12060 661 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 597 12060 661 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 597 11978 661 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 597 11978 661 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 597 11896 661 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 597 11896 661 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 597 11814 661 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 597 11814 661 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 597 11732 661 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 597 11732 661 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 597 11650 661 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 597 11650 661 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 515 12470 579 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 515 12470 579 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 515 12388 579 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 515 12388 579 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 515 12306 579 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 515 12306 579 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 515 12224 579 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 515 12224 579 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 515 12142 579 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 515 12142 579 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 515 12060 579 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 515 12060 579 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 515 11978 579 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 515 11978 579 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 515 11896 579 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 515 11896 579 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 515 11814 579 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 515 11814 579 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 515 11732 579 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 515 11732 579 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 515 11650 579 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 515 11650 579 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 433 12470 497 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 433 12470 497 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 433 12388 497 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 433 12388 497 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 433 12306 497 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 433 12306 497 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 433 12224 497 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 433 12224 497 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 433 12142 497 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 433 12142 497 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 433 12060 497 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 433 12060 497 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 433 11978 497 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 433 11978 497 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 433 11896 497 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 433 11896 497 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 433 11814 497 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 433 11814 497 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 433 11732 497 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 433 11732 497 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 433 11650 497 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 433 11650 497 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 351 12470 415 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 351 12470 415 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 351 12388 415 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 351 12388 415 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 351 12306 415 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 351 12306 415 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 351 12224 415 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 351 12224 415 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 351 12142 415 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 351 12142 415 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 351 12060 415 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 351 12060 415 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 351 11978 415 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 351 11978 415 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 351 11896 415 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 351 11896 415 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 351 11814 415 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 351 11814 415 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 351 11732 415 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 351 11732 415 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 351 11650 415 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 351 11650 415 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 269 12470 333 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 269 12470 333 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 269 12388 333 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 269 12388 333 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 269 12306 333 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 269 12306 333 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 269 12224 333 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 269 12224 333 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 269 12142 333 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 269 12142 333 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 269 12060 333 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 269 12060 333 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 269 11978 333 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 269 11978 333 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 269 11896 333 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 269 11896 333 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 269 11814 333 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 269 11814 333 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 269 11732 333 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 269 11732 333 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 269 11650 333 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 269 11650 333 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 187 12470 251 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 187 12388 251 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 187 12306 251 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 187 12224 251 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 187 12142 251 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 187 12060 251 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 187 11978 251 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 187 11896 251 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 187 11814 251 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 187 11732 251 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 187 11650 251 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 105 12470 169 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 105 12388 169 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 105 12306 169 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 105 12224 169 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 105 12142 169 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 105 12060 169 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 105 11978 169 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 105 11896 169 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 105 11814 169 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 105 11732 169 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 105 11650 169 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal5 s 0 3007 193 3657 6 VDDA
port 8 nsew power bidirectional
rlabel metal5 s 14807 3007 15000 3657 6 VDDA
port 8 nsew power bidirectional
rlabel metal4 s 0 2987 193 3677 6 VDDA
port 8 nsew power bidirectional
rlabel metal4 s 14807 2987 15000 3677 6 VDDA
port 8 nsew power bidirectional
rlabel metal5 s 0 1797 254 2687 6 VCCD
port 9 nsew power bidirectional
rlabel metal5 s 14746 1797 15000 2687 6 VCCD
port 9 nsew power bidirectional
rlabel metal4 s 0 1777 254 2707 6 VCCD
port 9 nsew power bidirectional
rlabel metal4 s 14746 1777 15000 2707 6 VCCD
port 9 nsew power bidirectional
rlabel metal5 s 0 427 254 1477 6 VCCHIB
port 10 nsew power bidirectional
rlabel metal5 s 14746 427 15000 1477 6 VCCHIB
port 10 nsew power bidirectional
rlabel metal4 s 0 407 254 1497 6 VCCHIB
port 10 nsew power bidirectional
rlabel metal4 s 14746 407 15000 1497 6 VCCHIB
port 10 nsew power bidirectional
rlabel metal4 s 0 9673 15000 10269 6 AMUXBUS_B
port 11 nsew signal bidirectional
rlabel metal4 s 0 10625 15000 11221 6 AMUXBUS_A
port 12 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 15000 40000
string LEFclass PAD
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 12408642
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 11933472
<< end >>
