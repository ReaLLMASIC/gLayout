magic
tech sky130A
timestamp 1701704242
<< metal1 >>
rect 0 0 3 122
rect 157 0 160 122
<< via1 >>
rect 3 0 157 122
<< metal2 >>
rect 0 0 3 122
rect 157 0 160 122
<< properties >>
string GDS_END 85426374
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85424962
<< end >>
