magic
tech sky130A
timestamp 1701704242
<< properties >>
string GDS_END 90827054
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 90826350
<< end >>
