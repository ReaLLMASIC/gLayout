magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< dnwell >>
rect 626 9736 14336 36182
<< nwell >>
rect 517 35918 14447 36293
rect 517 10000 832 35918
rect 1593 28312 13423 28975
rect 1593 27622 2336 28312
rect 12680 27622 13423 28312
rect 1593 26878 13423 27622
rect 14072 10000 14447 35918
rect 517 9625 14447 10000
<< pwell >>
rect 219 36363 14750 36600
rect 219 9554 456 36363
rect 1093 34577 13913 34747
rect 1093 10345 1263 34577
rect 13743 10345 13913 34577
rect 1093 10175 13913 10345
rect 14513 9554 14750 36363
rect 219 9317 14750 9554
<< mvpsubdiff >>
rect 245 36497 14724 36574
rect 245 36463 455 36497
rect 489 36463 523 36497
rect 557 36463 591 36497
rect 625 36463 659 36497
rect 693 36463 727 36497
rect 761 36463 795 36497
rect 829 36463 863 36497
rect 897 36463 931 36497
rect 965 36463 999 36497
rect 1033 36463 1067 36497
rect 1101 36463 1135 36497
rect 1169 36463 1203 36497
rect 1237 36463 1271 36497
rect 1305 36463 1339 36497
rect 1373 36463 1407 36497
rect 1441 36463 1475 36497
rect 1509 36463 1543 36497
rect 1577 36463 1611 36497
rect 1645 36463 1679 36497
rect 1713 36463 1747 36497
rect 1781 36463 1815 36497
rect 1849 36463 1883 36497
rect 1917 36463 1951 36497
rect 1985 36463 2019 36497
rect 2053 36463 2087 36497
rect 2121 36463 2155 36497
rect 2189 36463 2223 36497
rect 2257 36463 2291 36497
rect 2325 36463 2359 36497
rect 2393 36463 2427 36497
rect 2461 36463 2495 36497
rect 2529 36463 2563 36497
rect 2597 36463 2631 36497
rect 2665 36463 2699 36497
rect 2733 36463 2767 36497
rect 2801 36463 2835 36497
rect 2869 36463 2903 36497
rect 2937 36463 2971 36497
rect 3005 36463 3039 36497
rect 3073 36463 3107 36497
rect 3141 36463 3175 36497
rect 3209 36463 3243 36497
rect 3277 36463 3311 36497
rect 3345 36463 3379 36497
rect 3413 36463 3447 36497
rect 3481 36463 3515 36497
rect 3549 36463 3583 36497
rect 3617 36463 3651 36497
rect 3685 36463 3719 36497
rect 3753 36463 3787 36497
rect 3821 36463 3855 36497
rect 3889 36463 3923 36497
rect 3957 36463 3991 36497
rect 4025 36463 4059 36497
rect 4093 36463 4127 36497
rect 4161 36463 4195 36497
rect 4229 36463 4263 36497
rect 4297 36463 4331 36497
rect 4365 36463 4399 36497
rect 4433 36463 4467 36497
rect 4501 36463 4535 36497
rect 4569 36463 4603 36497
rect 4637 36463 4671 36497
rect 4705 36463 4739 36497
rect 4773 36463 4807 36497
rect 4841 36463 4875 36497
rect 4909 36463 4943 36497
rect 4977 36463 5011 36497
rect 5045 36463 5079 36497
rect 5113 36463 5147 36497
rect 5181 36463 5215 36497
rect 5249 36463 5283 36497
rect 5317 36463 5351 36497
rect 5385 36463 5419 36497
rect 5453 36463 5487 36497
rect 5521 36463 5555 36497
rect 5589 36463 5623 36497
rect 5657 36463 5691 36497
rect 5725 36463 5759 36497
rect 5793 36463 5827 36497
rect 5861 36463 5895 36497
rect 5929 36463 5963 36497
rect 5997 36463 6031 36497
rect 6065 36463 6099 36497
rect 6133 36463 6167 36497
rect 6201 36463 6235 36497
rect 6269 36463 6303 36497
rect 6337 36463 6371 36497
rect 6405 36463 6439 36497
rect 6473 36463 6507 36497
rect 6541 36463 6575 36497
rect 6609 36463 6643 36497
rect 6677 36463 6711 36497
rect 6745 36463 6779 36497
rect 6813 36463 6847 36497
rect 6881 36463 6915 36497
rect 6949 36463 6983 36497
rect 7017 36463 7051 36497
rect 7085 36463 7119 36497
rect 7153 36463 7187 36497
rect 7221 36463 7255 36497
rect 7289 36463 7323 36497
rect 7357 36463 7391 36497
rect 7425 36463 7459 36497
rect 7493 36463 7527 36497
rect 7561 36463 7595 36497
rect 7629 36463 7663 36497
rect 7697 36463 7731 36497
rect 7765 36463 7799 36497
rect 7833 36463 7867 36497
rect 7901 36463 7935 36497
rect 7969 36463 8003 36497
rect 8037 36463 8071 36497
rect 8105 36463 8139 36497
rect 8173 36463 8207 36497
rect 8241 36463 8275 36497
rect 8309 36463 8343 36497
rect 8377 36463 8411 36497
rect 8445 36463 8479 36497
rect 8513 36463 8547 36497
rect 8581 36463 8615 36497
rect 8649 36463 8683 36497
rect 8717 36463 8751 36497
rect 8785 36463 8819 36497
rect 8853 36463 8887 36497
rect 8921 36463 8955 36497
rect 8989 36463 9023 36497
rect 9057 36463 9091 36497
rect 9125 36463 9159 36497
rect 9193 36463 9227 36497
rect 9261 36463 9295 36497
rect 9329 36463 9363 36497
rect 9397 36463 9431 36497
rect 9465 36463 9499 36497
rect 9533 36463 9567 36497
rect 9601 36463 9635 36497
rect 9669 36463 9703 36497
rect 9737 36463 9771 36497
rect 9805 36463 9839 36497
rect 9873 36463 9907 36497
rect 9941 36463 9975 36497
rect 10009 36463 10043 36497
rect 10077 36463 10111 36497
rect 10145 36463 10179 36497
rect 10213 36463 10247 36497
rect 10281 36463 10315 36497
rect 10349 36463 10383 36497
rect 10417 36463 10451 36497
rect 10485 36463 10519 36497
rect 10553 36463 10587 36497
rect 10621 36463 10655 36497
rect 10689 36463 10723 36497
rect 10757 36463 10791 36497
rect 10825 36463 10859 36497
rect 10893 36463 10927 36497
rect 10961 36463 10995 36497
rect 11029 36463 11063 36497
rect 11097 36463 11131 36497
rect 11165 36463 11199 36497
rect 11233 36463 11267 36497
rect 11301 36463 11335 36497
rect 11369 36463 11403 36497
rect 11437 36463 11471 36497
rect 11505 36463 11539 36497
rect 11573 36463 11607 36497
rect 11641 36463 11675 36497
rect 11709 36463 11743 36497
rect 11777 36463 11811 36497
rect 11845 36463 11879 36497
rect 11913 36463 11947 36497
rect 11981 36463 12015 36497
rect 12049 36463 12083 36497
rect 12117 36463 12151 36497
rect 12185 36463 12219 36497
rect 12253 36463 12287 36497
rect 12321 36463 12355 36497
rect 12389 36463 12423 36497
rect 12457 36463 12491 36497
rect 12525 36463 12559 36497
rect 12593 36463 12627 36497
rect 12661 36463 12695 36497
rect 12729 36463 12763 36497
rect 12797 36463 12831 36497
rect 12865 36463 12899 36497
rect 12933 36463 12967 36497
rect 13001 36463 13035 36497
rect 13069 36463 13103 36497
rect 13137 36463 13171 36497
rect 13205 36463 13239 36497
rect 13273 36463 13307 36497
rect 13341 36463 13375 36497
rect 13409 36463 13443 36497
rect 13477 36463 13511 36497
rect 13545 36463 13579 36497
rect 13613 36463 13647 36497
rect 13681 36463 13715 36497
rect 13749 36463 13783 36497
rect 13817 36463 13851 36497
rect 13885 36463 13919 36497
rect 13953 36463 13987 36497
rect 14021 36463 14055 36497
rect 14089 36463 14123 36497
rect 14157 36463 14191 36497
rect 14225 36463 14259 36497
rect 14293 36463 14327 36497
rect 14361 36463 14395 36497
rect 14429 36463 14463 36497
rect 14497 36463 14724 36497
rect 245 36389 14724 36463
rect 245 36338 430 36389
rect 245 36304 312 36338
rect 346 36304 430 36338
rect 245 36270 430 36304
rect 245 36236 312 36270
rect 346 36236 430 36270
rect 245 36202 430 36236
rect 14539 36344 14724 36389
rect 14539 36310 14607 36344
rect 14641 36310 14724 36344
rect 14539 36276 14724 36310
rect 14539 36242 14607 36276
rect 14641 36242 14724 36276
rect 245 36168 312 36202
rect 346 36168 430 36202
rect 245 36134 430 36168
rect 245 36100 312 36134
rect 346 36100 430 36134
rect 245 36066 430 36100
rect 245 36032 312 36066
rect 346 36032 430 36066
rect 245 35998 430 36032
rect 245 35964 312 35998
rect 346 35964 430 35998
rect 245 35930 430 35964
rect 245 35896 312 35930
rect 346 35896 430 35930
rect 245 35862 430 35896
rect 245 35828 312 35862
rect 346 35828 430 35862
rect 245 35794 430 35828
rect 245 35760 312 35794
rect 346 35760 430 35794
rect 245 35726 430 35760
rect 245 35692 312 35726
rect 346 35692 430 35726
rect 245 35658 430 35692
rect 245 35624 312 35658
rect 346 35624 430 35658
rect 245 35590 430 35624
rect 245 35556 312 35590
rect 346 35556 430 35590
rect 245 35522 430 35556
rect 245 35488 312 35522
rect 346 35488 430 35522
rect 245 35454 430 35488
rect 245 35420 312 35454
rect 346 35420 430 35454
rect 245 35386 430 35420
rect 245 35352 312 35386
rect 346 35352 430 35386
rect 245 35318 430 35352
rect 245 35284 312 35318
rect 346 35284 430 35318
rect 245 35250 430 35284
rect 245 35216 312 35250
rect 346 35216 430 35250
rect 245 35182 430 35216
rect 245 35148 312 35182
rect 346 35148 430 35182
rect 245 35114 430 35148
rect 245 35080 312 35114
rect 346 35080 430 35114
rect 245 35046 430 35080
rect 245 35012 312 35046
rect 346 35012 430 35046
rect 245 34978 430 35012
rect 245 34944 312 34978
rect 346 34944 430 34978
rect 245 34910 430 34944
rect 245 34876 312 34910
rect 346 34876 430 34910
rect 245 34842 430 34876
rect 245 34808 312 34842
rect 346 34808 430 34842
rect 245 34774 430 34808
rect 245 34740 312 34774
rect 346 34740 430 34774
rect 245 34706 430 34740
rect 245 34672 312 34706
rect 346 34672 430 34706
rect 245 34638 430 34672
rect 245 34604 312 34638
rect 346 34604 430 34638
rect 245 34570 430 34604
rect 245 34536 312 34570
rect 346 34536 430 34570
rect 245 34502 430 34536
rect 245 34468 312 34502
rect 346 34468 430 34502
rect 245 34434 430 34468
rect 245 34400 312 34434
rect 346 34400 430 34434
rect 245 34366 430 34400
rect 245 34332 312 34366
rect 346 34332 430 34366
rect 245 34298 430 34332
rect 245 34264 312 34298
rect 346 34264 430 34298
rect 245 34230 430 34264
rect 245 34196 312 34230
rect 346 34196 430 34230
rect 245 34162 430 34196
rect 245 34128 312 34162
rect 346 34128 430 34162
rect 245 34094 430 34128
rect 245 34060 312 34094
rect 346 34060 430 34094
rect 245 34026 430 34060
rect 245 33992 312 34026
rect 346 33992 430 34026
rect 245 33958 430 33992
rect 245 33924 312 33958
rect 346 33924 430 33958
rect 245 33890 430 33924
rect 245 33856 312 33890
rect 346 33856 430 33890
rect 245 33822 430 33856
rect 245 33788 312 33822
rect 346 33788 430 33822
rect 245 33754 430 33788
rect 245 33720 312 33754
rect 346 33720 430 33754
rect 245 33686 430 33720
rect 245 33652 312 33686
rect 346 33652 430 33686
rect 245 33618 430 33652
rect 245 33584 312 33618
rect 346 33584 430 33618
rect 245 33550 430 33584
rect 245 33516 312 33550
rect 346 33516 430 33550
rect 245 33482 430 33516
rect 245 33448 312 33482
rect 346 33448 430 33482
rect 245 33414 430 33448
rect 245 33380 312 33414
rect 346 33380 430 33414
rect 245 33346 430 33380
rect 245 33312 312 33346
rect 346 33312 430 33346
rect 245 33278 430 33312
rect 245 33244 312 33278
rect 346 33244 430 33278
rect 245 33210 430 33244
rect 245 33176 312 33210
rect 346 33176 430 33210
rect 245 33142 430 33176
rect 245 33108 312 33142
rect 346 33108 430 33142
rect 245 33074 430 33108
rect 245 33040 312 33074
rect 346 33040 430 33074
rect 245 33006 430 33040
rect 245 32972 312 33006
rect 346 32972 430 33006
rect 245 32938 430 32972
rect 245 32904 312 32938
rect 346 32904 430 32938
rect 245 32870 430 32904
rect 245 32836 312 32870
rect 346 32836 430 32870
rect 245 32802 430 32836
rect 245 32768 312 32802
rect 346 32768 430 32802
rect 245 32734 430 32768
rect 245 32700 312 32734
rect 346 32700 430 32734
rect 245 32666 430 32700
rect 245 32632 312 32666
rect 346 32632 430 32666
rect 245 32598 430 32632
rect 245 32564 312 32598
rect 346 32564 430 32598
rect 245 32530 430 32564
rect 245 32496 312 32530
rect 346 32496 430 32530
rect 245 32462 430 32496
rect 245 32428 312 32462
rect 346 32428 430 32462
rect 245 32394 430 32428
rect 245 32360 312 32394
rect 346 32360 430 32394
rect 245 32326 430 32360
rect 245 32292 312 32326
rect 346 32292 430 32326
rect 245 32258 430 32292
rect 245 32224 312 32258
rect 346 32224 430 32258
rect 245 32190 430 32224
rect 245 32156 312 32190
rect 346 32156 430 32190
rect 245 32122 430 32156
rect 245 32088 312 32122
rect 346 32088 430 32122
rect 245 32054 430 32088
rect 245 32020 312 32054
rect 346 32020 430 32054
rect 245 31986 430 32020
rect 245 31952 312 31986
rect 346 31952 430 31986
rect 245 31918 430 31952
rect 245 31884 312 31918
rect 346 31884 430 31918
rect 245 31850 430 31884
rect 245 31816 312 31850
rect 346 31816 430 31850
rect 245 31782 430 31816
rect 245 31748 312 31782
rect 346 31748 430 31782
rect 245 31714 430 31748
rect 245 31680 312 31714
rect 346 31680 430 31714
rect 245 31646 430 31680
rect 245 31612 312 31646
rect 346 31612 430 31646
rect 245 31578 430 31612
rect 245 31544 312 31578
rect 346 31544 430 31578
rect 245 31510 430 31544
rect 245 31476 312 31510
rect 346 31476 430 31510
rect 245 31442 430 31476
rect 245 31408 312 31442
rect 346 31408 430 31442
rect 245 31374 430 31408
rect 245 31340 312 31374
rect 346 31340 430 31374
rect 245 31306 430 31340
rect 245 31272 312 31306
rect 346 31272 430 31306
rect 245 31238 430 31272
rect 245 31204 312 31238
rect 346 31204 430 31238
rect 245 31170 430 31204
rect 245 31136 312 31170
rect 346 31136 430 31170
rect 245 31102 430 31136
rect 245 31068 312 31102
rect 346 31068 430 31102
rect 245 31034 430 31068
rect 245 31000 312 31034
rect 346 31000 430 31034
rect 245 30966 430 31000
rect 245 30932 312 30966
rect 346 30932 430 30966
rect 245 30898 430 30932
rect 245 30864 312 30898
rect 346 30864 430 30898
rect 245 30830 430 30864
rect 245 30796 312 30830
rect 346 30796 430 30830
rect 245 30762 430 30796
rect 245 30728 312 30762
rect 346 30728 430 30762
rect 245 30694 430 30728
rect 245 30660 312 30694
rect 346 30660 430 30694
rect 245 30626 430 30660
rect 245 30592 312 30626
rect 346 30592 430 30626
rect 245 30558 430 30592
rect 245 30524 312 30558
rect 346 30524 430 30558
rect 245 30490 430 30524
rect 245 30456 312 30490
rect 346 30456 430 30490
rect 245 30422 430 30456
rect 245 30388 312 30422
rect 346 30388 430 30422
rect 245 30354 430 30388
rect 245 30320 312 30354
rect 346 30320 430 30354
rect 245 30286 430 30320
rect 245 30252 312 30286
rect 346 30252 430 30286
rect 245 30218 430 30252
rect 245 30184 312 30218
rect 346 30184 430 30218
rect 245 30150 430 30184
rect 245 30116 312 30150
rect 346 30116 430 30150
rect 245 30082 430 30116
rect 245 30048 312 30082
rect 346 30048 430 30082
rect 245 30014 430 30048
rect 245 29980 312 30014
rect 346 29980 430 30014
rect 245 29946 430 29980
rect 245 29912 312 29946
rect 346 29912 430 29946
rect 245 29878 430 29912
rect 245 29844 312 29878
rect 346 29844 430 29878
rect 245 29810 430 29844
rect 245 29776 312 29810
rect 346 29776 430 29810
rect 245 29742 430 29776
rect 245 29708 312 29742
rect 346 29708 430 29742
rect 245 29674 430 29708
rect 245 29640 312 29674
rect 346 29640 430 29674
rect 245 29606 430 29640
rect 245 29572 312 29606
rect 346 29572 430 29606
rect 245 29538 430 29572
rect 245 29504 312 29538
rect 346 29504 430 29538
rect 245 29470 430 29504
rect 245 29436 312 29470
rect 346 29436 430 29470
rect 245 29402 430 29436
rect 245 29368 312 29402
rect 346 29368 430 29402
rect 245 29334 430 29368
rect 245 29300 312 29334
rect 346 29300 430 29334
rect 245 29266 430 29300
rect 245 29232 312 29266
rect 346 29232 430 29266
rect 245 29198 430 29232
rect 245 29164 312 29198
rect 346 29164 430 29198
rect 245 29130 430 29164
rect 245 29096 312 29130
rect 346 29096 430 29130
rect 245 29062 430 29096
rect 245 29028 312 29062
rect 346 29028 430 29062
rect 245 28994 430 29028
rect 245 28960 312 28994
rect 346 28960 430 28994
rect 245 28926 430 28960
rect 245 28892 312 28926
rect 346 28892 430 28926
rect 245 28858 430 28892
rect 245 28824 312 28858
rect 346 28824 430 28858
rect 245 28790 430 28824
rect 245 28756 312 28790
rect 346 28756 430 28790
rect 245 28722 430 28756
rect 245 28688 312 28722
rect 346 28688 430 28722
rect 245 28654 430 28688
rect 245 28620 312 28654
rect 346 28620 430 28654
rect 245 28586 430 28620
rect 245 28552 312 28586
rect 346 28552 430 28586
rect 245 28518 430 28552
rect 245 28484 312 28518
rect 346 28484 430 28518
rect 245 28450 430 28484
rect 245 28416 312 28450
rect 346 28416 430 28450
rect 245 28382 430 28416
rect 245 28348 312 28382
rect 346 28348 430 28382
rect 245 28314 430 28348
rect 245 28280 312 28314
rect 346 28280 430 28314
rect 245 28246 430 28280
rect 245 28212 312 28246
rect 346 28212 430 28246
rect 245 28178 430 28212
rect 245 28144 312 28178
rect 346 28144 430 28178
rect 245 28110 430 28144
rect 245 28076 312 28110
rect 346 28076 430 28110
rect 245 28042 430 28076
rect 245 28008 312 28042
rect 346 28008 430 28042
rect 245 27974 430 28008
rect 245 27940 312 27974
rect 346 27940 430 27974
rect 245 27906 430 27940
rect 245 27872 312 27906
rect 346 27872 430 27906
rect 245 27838 430 27872
rect 245 27804 312 27838
rect 346 27804 430 27838
rect 245 27770 430 27804
rect 245 27736 312 27770
rect 346 27736 430 27770
rect 245 27702 430 27736
rect 245 27668 312 27702
rect 346 27668 430 27702
rect 245 27634 430 27668
rect 245 27600 312 27634
rect 346 27600 430 27634
rect 245 27566 430 27600
rect 245 27532 312 27566
rect 346 27532 430 27566
rect 245 27498 430 27532
rect 245 27464 312 27498
rect 346 27464 430 27498
rect 245 27430 430 27464
rect 245 27396 312 27430
rect 346 27396 430 27430
rect 245 27362 430 27396
rect 245 27328 312 27362
rect 346 27328 430 27362
rect 245 27294 430 27328
rect 245 27260 312 27294
rect 346 27260 430 27294
rect 245 27226 430 27260
rect 245 27192 312 27226
rect 346 27192 430 27226
rect 245 27158 430 27192
rect 245 27124 312 27158
rect 346 27124 430 27158
rect 245 27090 430 27124
rect 245 27056 312 27090
rect 346 27056 430 27090
rect 245 27022 430 27056
rect 245 26988 312 27022
rect 346 26988 430 27022
rect 245 26954 430 26988
rect 245 26920 312 26954
rect 346 26920 430 26954
rect 245 26886 430 26920
rect 245 26852 312 26886
rect 346 26852 430 26886
rect 245 26818 430 26852
rect 245 26784 312 26818
rect 346 26784 430 26818
rect 245 26750 430 26784
rect 245 26716 312 26750
rect 346 26716 430 26750
rect 245 26682 430 26716
rect 245 26648 312 26682
rect 346 26648 430 26682
rect 245 26614 430 26648
rect 245 26580 312 26614
rect 346 26580 430 26614
rect 245 26546 430 26580
rect 245 26512 312 26546
rect 346 26512 430 26546
rect 245 26478 430 26512
rect 245 26444 312 26478
rect 346 26444 430 26478
rect 245 26410 430 26444
rect 245 26376 312 26410
rect 346 26376 430 26410
rect 245 26342 430 26376
rect 245 26308 312 26342
rect 346 26308 430 26342
rect 245 26274 430 26308
rect 245 26240 312 26274
rect 346 26240 430 26274
rect 245 26206 430 26240
rect 245 26172 312 26206
rect 346 26172 430 26206
rect 245 26138 430 26172
rect 245 26104 312 26138
rect 346 26104 430 26138
rect 245 26070 430 26104
rect 245 26036 312 26070
rect 346 26036 430 26070
rect 245 26002 430 26036
rect 245 25968 312 26002
rect 346 25968 430 26002
rect 245 25934 430 25968
rect 245 25900 312 25934
rect 346 25900 430 25934
rect 245 25866 430 25900
rect 245 25832 312 25866
rect 346 25832 430 25866
rect 245 25798 430 25832
rect 245 25764 312 25798
rect 346 25764 430 25798
rect 245 25730 430 25764
rect 245 25696 312 25730
rect 346 25696 430 25730
rect 245 25662 430 25696
rect 245 25628 312 25662
rect 346 25628 430 25662
rect 245 25594 430 25628
rect 245 25560 312 25594
rect 346 25560 430 25594
rect 245 25526 430 25560
rect 245 25492 312 25526
rect 346 25492 430 25526
rect 245 25458 430 25492
rect 245 25424 312 25458
rect 346 25424 430 25458
rect 245 25390 430 25424
rect 245 25356 312 25390
rect 346 25356 430 25390
rect 245 25322 430 25356
rect 245 25288 312 25322
rect 346 25288 430 25322
rect 245 25254 430 25288
rect 245 25220 312 25254
rect 346 25220 430 25254
rect 245 25186 430 25220
rect 245 25152 312 25186
rect 346 25152 430 25186
rect 245 25118 430 25152
rect 245 25084 312 25118
rect 346 25084 430 25118
rect 245 25050 430 25084
rect 245 25016 312 25050
rect 346 25016 430 25050
rect 245 24982 430 25016
rect 245 24948 312 24982
rect 346 24948 430 24982
rect 245 24914 430 24948
rect 245 24880 312 24914
rect 346 24880 430 24914
rect 245 24846 430 24880
rect 245 24812 312 24846
rect 346 24812 430 24846
rect 245 24778 430 24812
rect 245 24744 312 24778
rect 346 24744 430 24778
rect 245 24710 430 24744
rect 245 24676 312 24710
rect 346 24676 430 24710
rect 245 24642 430 24676
rect 245 24608 312 24642
rect 346 24608 430 24642
rect 245 24574 430 24608
rect 245 24540 312 24574
rect 346 24540 430 24574
rect 245 24506 430 24540
rect 245 24472 312 24506
rect 346 24472 430 24506
rect 245 24438 430 24472
rect 245 24404 312 24438
rect 346 24404 430 24438
rect 245 24370 430 24404
rect 245 24336 312 24370
rect 346 24336 430 24370
rect 245 24302 430 24336
rect 245 24268 312 24302
rect 346 24268 430 24302
rect 245 24234 430 24268
rect 245 24200 312 24234
rect 346 24200 430 24234
rect 245 24166 430 24200
rect 245 24132 312 24166
rect 346 24132 430 24166
rect 245 24098 430 24132
rect 245 24064 312 24098
rect 346 24064 430 24098
rect 245 24030 430 24064
rect 245 23996 312 24030
rect 346 23996 430 24030
rect 245 23962 430 23996
rect 245 23928 312 23962
rect 346 23928 430 23962
rect 245 23894 430 23928
rect 245 23860 312 23894
rect 346 23860 430 23894
rect 245 23826 430 23860
rect 245 23792 312 23826
rect 346 23792 430 23826
rect 245 23758 430 23792
rect 245 23724 312 23758
rect 346 23724 430 23758
rect 245 23690 430 23724
rect 245 23656 312 23690
rect 346 23656 430 23690
rect 245 23622 430 23656
rect 245 23588 312 23622
rect 346 23588 430 23622
rect 245 23554 430 23588
rect 245 23520 312 23554
rect 346 23520 430 23554
rect 245 23486 430 23520
rect 245 23452 312 23486
rect 346 23452 430 23486
rect 245 23418 430 23452
rect 245 23384 312 23418
rect 346 23384 430 23418
rect 245 23350 430 23384
rect 245 23316 312 23350
rect 346 23316 430 23350
rect 245 23282 430 23316
rect 245 23248 312 23282
rect 346 23248 430 23282
rect 245 23214 430 23248
rect 245 23180 312 23214
rect 346 23180 430 23214
rect 245 23146 430 23180
rect 245 23112 312 23146
rect 346 23112 430 23146
rect 245 23078 430 23112
rect 245 23044 312 23078
rect 346 23044 430 23078
rect 245 23010 430 23044
rect 245 22976 312 23010
rect 346 22976 430 23010
rect 245 22942 430 22976
rect 245 22908 312 22942
rect 346 22908 430 22942
rect 245 22874 430 22908
rect 245 22840 312 22874
rect 346 22840 430 22874
rect 245 22806 430 22840
rect 245 22772 312 22806
rect 346 22772 430 22806
rect 245 22738 430 22772
rect 245 22704 312 22738
rect 346 22704 430 22738
rect 245 22670 430 22704
rect 245 22636 312 22670
rect 346 22636 430 22670
rect 245 22602 430 22636
rect 245 22568 312 22602
rect 346 22568 430 22602
rect 245 22534 430 22568
rect 245 22500 312 22534
rect 346 22500 430 22534
rect 245 22466 430 22500
rect 245 22432 312 22466
rect 346 22432 430 22466
rect 245 22398 430 22432
rect 245 22364 312 22398
rect 346 22364 430 22398
rect 245 22330 430 22364
rect 245 22296 312 22330
rect 346 22296 430 22330
rect 245 22262 430 22296
rect 245 22228 312 22262
rect 346 22228 430 22262
rect 245 22194 430 22228
rect 245 22160 312 22194
rect 346 22160 430 22194
rect 245 22126 430 22160
rect 245 22092 312 22126
rect 346 22092 430 22126
rect 245 22058 430 22092
rect 245 22024 312 22058
rect 346 22024 430 22058
rect 245 21990 430 22024
rect 245 21956 312 21990
rect 346 21956 430 21990
rect 245 21922 430 21956
rect 245 21888 312 21922
rect 346 21888 430 21922
rect 245 21854 430 21888
rect 245 21820 312 21854
rect 346 21820 430 21854
rect 245 21786 430 21820
rect 245 21752 312 21786
rect 346 21752 430 21786
rect 245 21718 430 21752
rect 245 21684 312 21718
rect 346 21684 430 21718
rect 245 21650 430 21684
rect 245 21616 312 21650
rect 346 21616 430 21650
rect 245 21582 430 21616
rect 245 21548 312 21582
rect 346 21548 430 21582
rect 245 21514 430 21548
rect 245 21480 312 21514
rect 346 21480 430 21514
rect 245 21446 430 21480
rect 245 21412 312 21446
rect 346 21412 430 21446
rect 245 21378 430 21412
rect 245 21344 312 21378
rect 346 21344 430 21378
rect 245 21310 430 21344
rect 245 21276 312 21310
rect 346 21276 430 21310
rect 245 21242 430 21276
rect 245 21208 312 21242
rect 346 21208 430 21242
rect 245 21174 430 21208
rect 245 21140 312 21174
rect 346 21140 430 21174
rect 245 21106 430 21140
rect 245 21072 312 21106
rect 346 21072 430 21106
rect 245 21038 430 21072
rect 245 21004 312 21038
rect 346 21004 430 21038
rect 245 20970 430 21004
rect 245 20936 312 20970
rect 346 20936 430 20970
rect 245 20902 430 20936
rect 245 20868 312 20902
rect 346 20868 430 20902
rect 245 20834 430 20868
rect 245 20800 312 20834
rect 346 20800 430 20834
rect 245 20766 430 20800
rect 245 20732 312 20766
rect 346 20732 430 20766
rect 245 20698 430 20732
rect 245 20664 312 20698
rect 346 20664 430 20698
rect 245 20630 430 20664
rect 245 20596 312 20630
rect 346 20596 430 20630
rect 245 20562 430 20596
rect 245 20528 312 20562
rect 346 20528 430 20562
rect 245 20494 430 20528
rect 245 20460 312 20494
rect 346 20460 430 20494
rect 245 20426 430 20460
rect 245 20392 312 20426
rect 346 20392 430 20426
rect 245 20358 430 20392
rect 245 20324 312 20358
rect 346 20324 430 20358
rect 245 20290 430 20324
rect 245 20256 312 20290
rect 346 20256 430 20290
rect 245 20222 430 20256
rect 245 20188 312 20222
rect 346 20188 430 20222
rect 245 20154 430 20188
rect 245 20120 312 20154
rect 346 20120 430 20154
rect 245 20086 430 20120
rect 245 20052 312 20086
rect 346 20052 430 20086
rect 245 20018 430 20052
rect 245 19984 312 20018
rect 346 19984 430 20018
rect 245 19950 430 19984
rect 245 19916 312 19950
rect 346 19916 430 19950
rect 245 19882 430 19916
rect 245 19848 312 19882
rect 346 19848 430 19882
rect 245 19814 430 19848
rect 245 19780 312 19814
rect 346 19780 430 19814
rect 245 19746 430 19780
rect 245 19712 312 19746
rect 346 19712 430 19746
rect 245 19678 430 19712
rect 245 19644 312 19678
rect 346 19644 430 19678
rect 245 19610 430 19644
rect 245 19576 312 19610
rect 346 19576 430 19610
rect 245 19542 430 19576
rect 245 19508 312 19542
rect 346 19508 430 19542
rect 245 19474 430 19508
rect 245 19440 312 19474
rect 346 19440 430 19474
rect 245 19406 430 19440
rect 245 19372 312 19406
rect 346 19372 430 19406
rect 245 19338 430 19372
rect 245 19304 312 19338
rect 346 19304 430 19338
rect 245 19270 430 19304
rect 245 19236 312 19270
rect 346 19236 430 19270
rect 245 19202 430 19236
rect 245 19168 312 19202
rect 346 19168 430 19202
rect 245 19134 430 19168
rect 245 19100 312 19134
rect 346 19100 430 19134
rect 245 19066 430 19100
rect 245 19032 312 19066
rect 346 19032 430 19066
rect 245 18998 430 19032
rect 245 18964 312 18998
rect 346 18964 430 18998
rect 245 18930 430 18964
rect 245 18896 312 18930
rect 346 18896 430 18930
rect 245 18862 430 18896
rect 245 18828 312 18862
rect 346 18828 430 18862
rect 245 18794 430 18828
rect 245 18760 312 18794
rect 346 18760 430 18794
rect 245 18726 430 18760
rect 245 18692 312 18726
rect 346 18692 430 18726
rect 245 18658 430 18692
rect 245 18624 312 18658
rect 346 18624 430 18658
rect 245 18590 430 18624
rect 245 18556 312 18590
rect 346 18556 430 18590
rect 245 18522 430 18556
rect 245 18488 312 18522
rect 346 18488 430 18522
rect 245 18454 430 18488
rect 245 18420 312 18454
rect 346 18420 430 18454
rect 245 18386 430 18420
rect 245 18352 312 18386
rect 346 18352 430 18386
rect 245 18318 430 18352
rect 245 18284 312 18318
rect 346 18284 430 18318
rect 245 18250 430 18284
rect 245 18216 312 18250
rect 346 18216 430 18250
rect 245 18182 430 18216
rect 245 18148 312 18182
rect 346 18148 430 18182
rect 245 18114 430 18148
rect 245 18080 312 18114
rect 346 18080 430 18114
rect 245 18046 430 18080
rect 245 18012 312 18046
rect 346 18012 430 18046
rect 245 17978 430 18012
rect 245 17944 312 17978
rect 346 17944 430 17978
rect 245 17910 430 17944
rect 245 17876 312 17910
rect 346 17876 430 17910
rect 245 17842 430 17876
rect 245 17808 312 17842
rect 346 17808 430 17842
rect 245 17774 430 17808
rect 245 17740 312 17774
rect 346 17740 430 17774
rect 245 17706 430 17740
rect 245 17672 312 17706
rect 346 17672 430 17706
rect 245 17638 430 17672
rect 245 17604 312 17638
rect 346 17604 430 17638
rect 245 17570 430 17604
rect 245 17536 312 17570
rect 346 17536 430 17570
rect 245 17502 430 17536
rect 245 17468 312 17502
rect 346 17468 430 17502
rect 245 17434 430 17468
rect 245 17400 312 17434
rect 346 17400 430 17434
rect 245 17366 430 17400
rect 245 17332 312 17366
rect 346 17332 430 17366
rect 245 17298 430 17332
rect 245 17264 312 17298
rect 346 17264 430 17298
rect 245 17230 430 17264
rect 245 17196 312 17230
rect 346 17196 430 17230
rect 245 17162 430 17196
rect 245 17128 312 17162
rect 346 17128 430 17162
rect 245 17094 430 17128
rect 245 17060 312 17094
rect 346 17060 430 17094
rect 245 17026 430 17060
rect 245 16992 312 17026
rect 346 16992 430 17026
rect 245 16958 430 16992
rect 245 16924 312 16958
rect 346 16924 430 16958
rect 245 16890 430 16924
rect 245 16856 312 16890
rect 346 16856 430 16890
rect 245 16822 430 16856
rect 245 16788 312 16822
rect 346 16788 430 16822
rect 245 16754 430 16788
rect 245 16720 312 16754
rect 346 16720 430 16754
rect 245 16686 430 16720
rect 245 16652 312 16686
rect 346 16652 430 16686
rect 245 16618 430 16652
rect 245 16584 312 16618
rect 346 16584 430 16618
rect 245 16550 430 16584
rect 245 16516 312 16550
rect 346 16516 430 16550
rect 245 16482 430 16516
rect 245 16448 312 16482
rect 346 16448 430 16482
rect 245 16414 430 16448
rect 245 16380 312 16414
rect 346 16380 430 16414
rect 245 16346 430 16380
rect 245 16312 312 16346
rect 346 16312 430 16346
rect 245 16278 430 16312
rect 245 16244 312 16278
rect 346 16244 430 16278
rect 245 16210 430 16244
rect 245 16176 312 16210
rect 346 16176 430 16210
rect 245 16142 430 16176
rect 245 16108 312 16142
rect 346 16108 430 16142
rect 245 16074 430 16108
rect 245 16040 312 16074
rect 346 16040 430 16074
rect 245 16006 430 16040
rect 245 15972 312 16006
rect 346 15972 430 16006
rect 245 15938 430 15972
rect 245 15904 312 15938
rect 346 15904 430 15938
rect 245 15870 430 15904
rect 245 15836 312 15870
rect 346 15836 430 15870
rect 245 15802 430 15836
rect 245 15768 312 15802
rect 346 15768 430 15802
rect 245 15734 430 15768
rect 245 15700 312 15734
rect 346 15700 430 15734
rect 245 15666 430 15700
rect 245 15632 312 15666
rect 346 15632 430 15666
rect 245 15598 430 15632
rect 245 15564 312 15598
rect 346 15564 430 15598
rect 245 15530 430 15564
rect 245 15496 312 15530
rect 346 15496 430 15530
rect 245 15462 430 15496
rect 245 15428 312 15462
rect 346 15428 430 15462
rect 245 15394 430 15428
rect 245 15360 312 15394
rect 346 15360 430 15394
rect 245 15326 430 15360
rect 245 15292 312 15326
rect 346 15292 430 15326
rect 245 15258 430 15292
rect 245 15224 312 15258
rect 346 15224 430 15258
rect 245 15190 430 15224
rect 245 15156 312 15190
rect 346 15156 430 15190
rect 245 15122 430 15156
rect 245 15088 312 15122
rect 346 15088 430 15122
rect 245 15054 430 15088
rect 245 15020 312 15054
rect 346 15020 430 15054
rect 245 14986 430 15020
rect 245 14952 312 14986
rect 346 14952 430 14986
rect 245 14918 430 14952
rect 245 14884 312 14918
rect 346 14884 430 14918
rect 245 14850 430 14884
rect 245 14816 312 14850
rect 346 14816 430 14850
rect 245 14782 430 14816
rect 245 14748 312 14782
rect 346 14748 430 14782
rect 245 14714 430 14748
rect 245 14680 312 14714
rect 346 14680 430 14714
rect 245 14646 430 14680
rect 245 14612 312 14646
rect 346 14612 430 14646
rect 245 14578 430 14612
rect 245 14544 312 14578
rect 346 14544 430 14578
rect 245 14510 430 14544
rect 245 14476 312 14510
rect 346 14476 430 14510
rect 245 14442 430 14476
rect 245 14408 312 14442
rect 346 14408 430 14442
rect 245 14374 430 14408
rect 245 14340 312 14374
rect 346 14340 430 14374
rect 245 14306 430 14340
rect 245 14272 312 14306
rect 346 14272 430 14306
rect 245 14238 430 14272
rect 245 14204 312 14238
rect 346 14204 430 14238
rect 245 14170 430 14204
rect 245 14136 312 14170
rect 346 14136 430 14170
rect 245 14102 430 14136
rect 245 14068 312 14102
rect 346 14068 430 14102
rect 245 14034 430 14068
rect 245 14000 312 14034
rect 346 14000 430 14034
rect 245 13966 430 14000
rect 245 13932 312 13966
rect 346 13932 430 13966
rect 245 13898 430 13932
rect 245 13864 312 13898
rect 346 13864 430 13898
rect 245 13830 430 13864
rect 245 13796 312 13830
rect 346 13796 430 13830
rect 245 13762 430 13796
rect 245 13728 312 13762
rect 346 13728 430 13762
rect 245 13694 430 13728
rect 245 13660 312 13694
rect 346 13660 430 13694
rect 245 13626 430 13660
rect 245 13592 312 13626
rect 346 13592 430 13626
rect 245 13558 430 13592
rect 245 13524 312 13558
rect 346 13524 430 13558
rect 245 13490 430 13524
rect 245 13456 312 13490
rect 346 13456 430 13490
rect 245 13422 430 13456
rect 245 13388 312 13422
rect 346 13388 430 13422
rect 245 13354 430 13388
rect 245 13320 312 13354
rect 346 13320 430 13354
rect 245 13286 430 13320
rect 245 13252 312 13286
rect 346 13252 430 13286
rect 245 13218 430 13252
rect 245 13184 312 13218
rect 346 13184 430 13218
rect 245 13150 430 13184
rect 245 13116 312 13150
rect 346 13116 430 13150
rect 245 13082 430 13116
rect 245 13048 312 13082
rect 346 13048 430 13082
rect 245 13014 430 13048
rect 245 12980 312 13014
rect 346 12980 430 13014
rect 245 12946 430 12980
rect 245 12912 312 12946
rect 346 12912 430 12946
rect 245 12878 430 12912
rect 245 12844 312 12878
rect 346 12844 430 12878
rect 245 12810 430 12844
rect 245 12776 312 12810
rect 346 12776 430 12810
rect 245 12742 430 12776
rect 245 12708 312 12742
rect 346 12708 430 12742
rect 245 12674 430 12708
rect 245 12640 312 12674
rect 346 12640 430 12674
rect 245 12606 430 12640
rect 245 12572 312 12606
rect 346 12572 430 12606
rect 245 12538 430 12572
rect 245 12504 312 12538
rect 346 12504 430 12538
rect 245 12470 430 12504
rect 245 12436 312 12470
rect 346 12436 430 12470
rect 245 12402 430 12436
rect 245 12368 312 12402
rect 346 12368 430 12402
rect 245 12334 430 12368
rect 245 12300 312 12334
rect 346 12300 430 12334
rect 245 12266 430 12300
rect 245 12232 312 12266
rect 346 12232 430 12266
rect 245 12198 430 12232
rect 245 12164 312 12198
rect 346 12164 430 12198
rect 245 12130 430 12164
rect 245 12096 312 12130
rect 346 12096 430 12130
rect 245 12062 430 12096
rect 245 12028 312 12062
rect 346 12028 430 12062
rect 245 11994 430 12028
rect 245 11960 312 11994
rect 346 11960 430 11994
rect 245 11926 430 11960
rect 245 11892 312 11926
rect 346 11892 430 11926
rect 245 11858 430 11892
rect 245 11824 312 11858
rect 346 11824 430 11858
rect 245 11790 430 11824
rect 245 11756 312 11790
rect 346 11756 430 11790
rect 245 11722 430 11756
rect 245 11688 312 11722
rect 346 11688 430 11722
rect 245 11654 430 11688
rect 245 11620 312 11654
rect 346 11620 430 11654
rect 245 11586 430 11620
rect 245 11552 312 11586
rect 346 11552 430 11586
rect 245 11518 430 11552
rect 245 11484 312 11518
rect 346 11484 430 11518
rect 245 11450 430 11484
rect 245 11416 312 11450
rect 346 11416 430 11450
rect 245 11382 430 11416
rect 245 11348 312 11382
rect 346 11348 430 11382
rect 245 11314 430 11348
rect 245 11280 312 11314
rect 346 11280 430 11314
rect 245 11246 430 11280
rect 245 11212 312 11246
rect 346 11212 430 11246
rect 245 11178 430 11212
rect 245 11144 312 11178
rect 346 11144 430 11178
rect 245 11110 430 11144
rect 245 11076 312 11110
rect 346 11076 430 11110
rect 245 11042 430 11076
rect 245 11008 312 11042
rect 346 11008 430 11042
rect 245 10974 430 11008
rect 245 10940 312 10974
rect 346 10940 430 10974
rect 245 10906 430 10940
rect 245 10872 312 10906
rect 346 10872 430 10906
rect 245 10838 430 10872
rect 245 10804 312 10838
rect 346 10804 430 10838
rect 245 10770 430 10804
rect 245 10736 312 10770
rect 346 10736 430 10770
rect 245 10702 430 10736
rect 245 10668 312 10702
rect 346 10668 430 10702
rect 245 10634 430 10668
rect 245 10600 312 10634
rect 346 10600 430 10634
rect 245 10566 430 10600
rect 245 10532 312 10566
rect 346 10532 430 10566
rect 245 10498 430 10532
rect 245 10464 312 10498
rect 346 10464 430 10498
rect 245 10430 430 10464
rect 245 10396 312 10430
rect 346 10396 430 10430
rect 245 10362 430 10396
rect 245 10328 312 10362
rect 346 10328 430 10362
rect 245 10294 430 10328
rect 245 10260 312 10294
rect 346 10260 430 10294
rect 245 10226 430 10260
rect 245 10192 312 10226
rect 346 10192 430 10226
rect 245 10158 430 10192
rect 245 10124 312 10158
rect 346 10124 430 10158
rect 245 10090 430 10124
rect 245 10056 312 10090
rect 346 10056 430 10090
rect 245 10022 430 10056
rect 245 9988 312 10022
rect 346 9988 430 10022
rect 245 9954 430 9988
rect 245 9920 312 9954
rect 346 9920 430 9954
rect 245 9886 430 9920
rect 245 9852 312 9886
rect 346 9852 430 9886
rect 245 9818 430 9852
rect 245 9784 312 9818
rect 346 9784 430 9818
rect 245 9750 430 9784
rect 245 9716 312 9750
rect 346 9716 430 9750
rect 245 9682 430 9716
rect 1119 34679 13887 34721
rect 1119 34645 1305 34679
rect 1339 34645 1373 34679
rect 1407 34645 1441 34679
rect 1475 34645 1509 34679
rect 1543 34645 1577 34679
rect 1611 34645 1645 34679
rect 1679 34645 1713 34679
rect 1747 34645 1781 34679
rect 1815 34645 1849 34679
rect 1883 34645 1917 34679
rect 1951 34645 1985 34679
rect 2019 34645 2053 34679
rect 2087 34645 2121 34679
rect 2155 34645 2189 34679
rect 2223 34645 2257 34679
rect 2291 34645 2325 34679
rect 2359 34645 2393 34679
rect 2427 34645 2461 34679
rect 2495 34645 2529 34679
rect 2563 34645 2597 34679
rect 2631 34645 2665 34679
rect 2699 34645 2733 34679
rect 2767 34645 2801 34679
rect 2835 34645 2869 34679
rect 2903 34645 2937 34679
rect 2971 34645 3005 34679
rect 3039 34645 3073 34679
rect 3107 34645 3141 34679
rect 3175 34645 3209 34679
rect 3243 34645 3277 34679
rect 3311 34645 3345 34679
rect 3379 34645 3413 34679
rect 3447 34645 3481 34679
rect 3515 34645 3549 34679
rect 3583 34645 3617 34679
rect 3651 34645 3685 34679
rect 3719 34645 3753 34679
rect 3787 34645 3821 34679
rect 3855 34645 3889 34679
rect 3923 34645 3957 34679
rect 3991 34645 4025 34679
rect 4059 34645 4093 34679
rect 4127 34645 4161 34679
rect 4195 34645 4229 34679
rect 4263 34645 4297 34679
rect 4331 34645 4365 34679
rect 4399 34645 4433 34679
rect 4467 34645 4501 34679
rect 4535 34645 4569 34679
rect 4603 34645 4637 34679
rect 4671 34645 4705 34679
rect 4739 34645 4773 34679
rect 4807 34645 4841 34679
rect 4875 34645 4909 34679
rect 4943 34645 4977 34679
rect 5011 34645 5045 34679
rect 5079 34645 5113 34679
rect 5147 34645 5181 34679
rect 5215 34645 5249 34679
rect 5283 34645 5317 34679
rect 5351 34645 5385 34679
rect 5419 34645 5453 34679
rect 5487 34645 5521 34679
rect 5555 34645 5589 34679
rect 5623 34645 5657 34679
rect 5691 34645 5725 34679
rect 5759 34645 5793 34679
rect 5827 34645 5861 34679
rect 5895 34645 5929 34679
rect 5963 34645 5997 34679
rect 6031 34645 6065 34679
rect 6099 34645 6133 34679
rect 6167 34645 6201 34679
rect 6235 34645 6269 34679
rect 6303 34645 6337 34679
rect 6371 34645 6405 34679
rect 6439 34645 6473 34679
rect 6507 34645 6541 34679
rect 6575 34645 6609 34679
rect 6643 34645 6677 34679
rect 6711 34645 6745 34679
rect 6779 34645 6813 34679
rect 6847 34645 6881 34679
rect 6915 34645 6949 34679
rect 6983 34645 7017 34679
rect 7051 34645 7085 34679
rect 7119 34645 7153 34679
rect 7187 34645 7221 34679
rect 7255 34645 7289 34679
rect 7323 34645 7357 34679
rect 7391 34645 7425 34679
rect 7459 34645 7493 34679
rect 7527 34645 7561 34679
rect 7595 34645 7629 34679
rect 7663 34645 7697 34679
rect 7731 34645 7765 34679
rect 7799 34645 7833 34679
rect 7867 34645 7901 34679
rect 7935 34645 7969 34679
rect 8003 34645 8037 34679
rect 8071 34645 8105 34679
rect 8139 34645 8173 34679
rect 8207 34645 8241 34679
rect 8275 34645 8309 34679
rect 8343 34645 8377 34679
rect 8411 34645 8445 34679
rect 8479 34645 8513 34679
rect 8547 34645 8581 34679
rect 8615 34645 8649 34679
rect 8683 34645 8717 34679
rect 8751 34645 8785 34679
rect 8819 34645 8853 34679
rect 8887 34645 8921 34679
rect 8955 34645 8989 34679
rect 9023 34645 9057 34679
rect 9091 34645 9125 34679
rect 9159 34645 9193 34679
rect 9227 34645 9261 34679
rect 9295 34645 9329 34679
rect 9363 34645 9397 34679
rect 9431 34645 9465 34679
rect 9499 34645 9533 34679
rect 9567 34645 9601 34679
rect 9635 34645 9669 34679
rect 9703 34645 9737 34679
rect 9771 34645 9805 34679
rect 9839 34645 9873 34679
rect 9907 34645 9941 34679
rect 9975 34645 10009 34679
rect 10043 34645 10077 34679
rect 10111 34645 10145 34679
rect 10179 34645 10213 34679
rect 10247 34645 10281 34679
rect 10315 34645 10349 34679
rect 10383 34645 10417 34679
rect 10451 34645 10485 34679
rect 10519 34645 10553 34679
rect 10587 34645 10621 34679
rect 10655 34645 10689 34679
rect 10723 34645 10757 34679
rect 10791 34645 10825 34679
rect 10859 34645 10893 34679
rect 10927 34645 10961 34679
rect 10995 34645 11029 34679
rect 11063 34645 11097 34679
rect 11131 34645 11165 34679
rect 11199 34645 11233 34679
rect 11267 34645 11301 34679
rect 11335 34645 11369 34679
rect 11403 34645 11437 34679
rect 11471 34645 11505 34679
rect 11539 34645 11573 34679
rect 11607 34645 11641 34679
rect 11675 34645 11709 34679
rect 11743 34645 11777 34679
rect 11811 34645 11845 34679
rect 11879 34645 11913 34679
rect 11947 34645 11981 34679
rect 12015 34645 12049 34679
rect 12083 34645 12117 34679
rect 12151 34645 12185 34679
rect 12219 34645 12253 34679
rect 12287 34645 12321 34679
rect 12355 34645 12389 34679
rect 12423 34645 12457 34679
rect 12491 34645 12525 34679
rect 12559 34645 12593 34679
rect 12627 34645 12661 34679
rect 12695 34645 12729 34679
rect 12763 34645 12797 34679
rect 12831 34645 12865 34679
rect 12899 34645 12933 34679
rect 12967 34645 13001 34679
rect 13035 34645 13069 34679
rect 13103 34645 13137 34679
rect 13171 34645 13205 34679
rect 13239 34645 13273 34679
rect 13307 34645 13341 34679
rect 13375 34645 13409 34679
rect 13443 34645 13477 34679
rect 13511 34645 13545 34679
rect 13579 34645 13613 34679
rect 13647 34645 13681 34679
rect 13715 34645 13887 34679
rect 1119 34603 13887 34645
rect 1119 34478 1237 34603
rect 1119 34444 1161 34478
rect 1195 34444 1237 34478
rect 1119 34410 1237 34444
rect 1119 34376 1161 34410
rect 1195 34376 1237 34410
rect 1119 34342 1237 34376
rect 1119 34308 1161 34342
rect 1195 34308 1237 34342
rect 1119 34274 1237 34308
rect 1119 34240 1161 34274
rect 1195 34240 1237 34274
rect 1119 34206 1237 34240
rect 1119 34172 1161 34206
rect 1195 34172 1237 34206
rect 1119 34138 1237 34172
rect 1119 34104 1161 34138
rect 1195 34104 1237 34138
rect 1119 34070 1237 34104
rect 1119 34036 1161 34070
rect 1195 34036 1237 34070
rect 1119 34002 1237 34036
rect 1119 33968 1161 34002
rect 1195 33968 1237 34002
rect 1119 33934 1237 33968
rect 1119 33900 1161 33934
rect 1195 33900 1237 33934
rect 1119 33866 1237 33900
rect 1119 33832 1161 33866
rect 1195 33832 1237 33866
rect 1119 33798 1237 33832
rect 1119 33764 1161 33798
rect 1195 33764 1237 33798
rect 1119 33730 1237 33764
rect 1119 33696 1161 33730
rect 1195 33696 1237 33730
rect 1119 33662 1237 33696
rect 1119 33628 1161 33662
rect 1195 33628 1237 33662
rect 1119 33594 1237 33628
rect 1119 33560 1161 33594
rect 1195 33560 1237 33594
rect 1119 33526 1237 33560
rect 1119 33492 1161 33526
rect 1195 33492 1237 33526
rect 1119 33458 1237 33492
rect 1119 33424 1161 33458
rect 1195 33424 1237 33458
rect 1119 33390 1237 33424
rect 1119 33356 1161 33390
rect 1195 33356 1237 33390
rect 1119 33322 1237 33356
rect 1119 33288 1161 33322
rect 1195 33288 1237 33322
rect 1119 33254 1237 33288
rect 1119 33220 1161 33254
rect 1195 33220 1237 33254
rect 1119 33186 1237 33220
rect 1119 33152 1161 33186
rect 1195 33152 1237 33186
rect 1119 33118 1237 33152
rect 1119 33084 1161 33118
rect 1195 33084 1237 33118
rect 1119 33050 1237 33084
rect 1119 33016 1161 33050
rect 1195 33016 1237 33050
rect 1119 32982 1237 33016
rect 1119 32948 1161 32982
rect 1195 32948 1237 32982
rect 1119 32914 1237 32948
rect 1119 32880 1161 32914
rect 1195 32880 1237 32914
rect 1119 32846 1237 32880
rect 1119 32812 1161 32846
rect 1195 32812 1237 32846
rect 1119 32778 1237 32812
rect 1119 32744 1161 32778
rect 1195 32744 1237 32778
rect 1119 32710 1237 32744
rect 1119 32676 1161 32710
rect 1195 32676 1237 32710
rect 1119 32642 1237 32676
rect 1119 32608 1161 32642
rect 1195 32608 1237 32642
rect 1119 32574 1237 32608
rect 1119 32540 1161 32574
rect 1195 32540 1237 32574
rect 1119 32506 1237 32540
rect 1119 32472 1161 32506
rect 1195 32472 1237 32506
rect 1119 32438 1237 32472
rect 1119 32404 1161 32438
rect 1195 32404 1237 32438
rect 1119 32370 1237 32404
rect 1119 32336 1161 32370
rect 1195 32336 1237 32370
rect 1119 32302 1237 32336
rect 1119 32268 1161 32302
rect 1195 32268 1237 32302
rect 1119 32234 1237 32268
rect 1119 32200 1161 32234
rect 1195 32200 1237 32234
rect 1119 32166 1237 32200
rect 1119 32132 1161 32166
rect 1195 32132 1237 32166
rect 1119 32098 1237 32132
rect 1119 32064 1161 32098
rect 1195 32064 1237 32098
rect 1119 32030 1237 32064
rect 1119 31996 1161 32030
rect 1195 31996 1237 32030
rect 1119 31962 1237 31996
rect 1119 31928 1161 31962
rect 1195 31928 1237 31962
rect 1119 31894 1237 31928
rect 1119 31860 1161 31894
rect 1195 31860 1237 31894
rect 1119 31826 1237 31860
rect 1119 31792 1161 31826
rect 1195 31792 1237 31826
rect 1119 31758 1237 31792
rect 1119 31724 1161 31758
rect 1195 31724 1237 31758
rect 1119 31690 1237 31724
rect 1119 31656 1161 31690
rect 1195 31656 1237 31690
rect 1119 31622 1237 31656
rect 1119 31588 1161 31622
rect 1195 31588 1237 31622
rect 1119 31554 1237 31588
rect 1119 31520 1161 31554
rect 1195 31520 1237 31554
rect 1119 31486 1237 31520
rect 1119 31452 1161 31486
rect 1195 31452 1237 31486
rect 1119 31418 1237 31452
rect 1119 31384 1161 31418
rect 1195 31384 1237 31418
rect 1119 31350 1237 31384
rect 1119 31316 1161 31350
rect 1195 31316 1237 31350
rect 1119 31282 1237 31316
rect 1119 31248 1161 31282
rect 1195 31248 1237 31282
rect 1119 31214 1237 31248
rect 1119 31180 1161 31214
rect 1195 31180 1237 31214
rect 1119 31146 1237 31180
rect 1119 31112 1161 31146
rect 1195 31112 1237 31146
rect 1119 31078 1237 31112
rect 1119 31044 1161 31078
rect 1195 31044 1237 31078
rect 1119 31010 1237 31044
rect 1119 30976 1161 31010
rect 1195 30976 1237 31010
rect 1119 30942 1237 30976
rect 1119 30908 1161 30942
rect 1195 30908 1237 30942
rect 1119 30874 1237 30908
rect 1119 30840 1161 30874
rect 1195 30840 1237 30874
rect 1119 30806 1237 30840
rect 1119 30772 1161 30806
rect 1195 30772 1237 30806
rect 1119 30738 1237 30772
rect 1119 30704 1161 30738
rect 1195 30704 1237 30738
rect 1119 30670 1237 30704
rect 1119 30636 1161 30670
rect 1195 30636 1237 30670
rect 1119 30602 1237 30636
rect 1119 30568 1161 30602
rect 1195 30568 1237 30602
rect 1119 30534 1237 30568
rect 1119 30500 1161 30534
rect 1195 30500 1237 30534
rect 1119 30466 1237 30500
rect 1119 30432 1161 30466
rect 1195 30432 1237 30466
rect 1119 30398 1237 30432
rect 1119 30364 1161 30398
rect 1195 30364 1237 30398
rect 1119 30330 1237 30364
rect 1119 30296 1161 30330
rect 1195 30296 1237 30330
rect 1119 30262 1237 30296
rect 1119 30228 1161 30262
rect 1195 30228 1237 30262
rect 1119 30194 1237 30228
rect 1119 30160 1161 30194
rect 1195 30160 1237 30194
rect 1119 30126 1237 30160
rect 1119 30092 1161 30126
rect 1195 30092 1237 30126
rect 1119 30058 1237 30092
rect 1119 30024 1161 30058
rect 1195 30024 1237 30058
rect 1119 29990 1237 30024
rect 1119 29956 1161 29990
rect 1195 29956 1237 29990
rect 1119 29922 1237 29956
rect 1119 29888 1161 29922
rect 1195 29888 1237 29922
rect 1119 29854 1237 29888
rect 1119 29820 1161 29854
rect 1195 29820 1237 29854
rect 1119 29786 1237 29820
rect 1119 29752 1161 29786
rect 1195 29752 1237 29786
rect 1119 29718 1237 29752
rect 1119 29684 1161 29718
rect 1195 29684 1237 29718
rect 1119 29650 1237 29684
rect 1119 29616 1161 29650
rect 1195 29616 1237 29650
rect 1119 29582 1237 29616
rect 1119 29548 1161 29582
rect 1195 29548 1237 29582
rect 1119 29514 1237 29548
rect 1119 29480 1161 29514
rect 1195 29480 1237 29514
rect 1119 29446 1237 29480
rect 1119 29412 1161 29446
rect 1195 29412 1237 29446
rect 1119 29378 1237 29412
rect 1119 29344 1161 29378
rect 1195 29344 1237 29378
rect 1119 29310 1237 29344
rect 1119 29276 1161 29310
rect 1195 29276 1237 29310
rect 1119 29242 1237 29276
rect 1119 29208 1161 29242
rect 1195 29208 1237 29242
rect 1119 29174 1237 29208
rect 1119 29140 1161 29174
rect 1195 29140 1237 29174
rect 1119 29106 1237 29140
rect 1119 29072 1161 29106
rect 1195 29072 1237 29106
rect 1119 29038 1237 29072
rect 1119 29004 1161 29038
rect 1195 29004 1237 29038
rect 1119 28970 1237 29004
rect 1119 28936 1161 28970
rect 1195 28936 1237 28970
rect 1119 28902 1237 28936
rect 13769 34473 13887 34603
rect 13769 34439 13809 34473
rect 13843 34439 13887 34473
rect 13769 34405 13887 34439
rect 13769 34371 13809 34405
rect 13843 34371 13887 34405
rect 13769 34337 13887 34371
rect 13769 34303 13809 34337
rect 13843 34303 13887 34337
rect 13769 34269 13887 34303
rect 13769 34235 13809 34269
rect 13843 34235 13887 34269
rect 13769 34201 13887 34235
rect 13769 34167 13809 34201
rect 13843 34167 13887 34201
rect 13769 34133 13887 34167
rect 13769 34099 13809 34133
rect 13843 34099 13887 34133
rect 13769 34065 13887 34099
rect 13769 34031 13809 34065
rect 13843 34031 13887 34065
rect 13769 33997 13887 34031
rect 13769 33963 13809 33997
rect 13843 33963 13887 33997
rect 13769 33929 13887 33963
rect 13769 33895 13809 33929
rect 13843 33895 13887 33929
rect 13769 33861 13887 33895
rect 13769 33827 13809 33861
rect 13843 33827 13887 33861
rect 13769 33793 13887 33827
rect 13769 33759 13809 33793
rect 13843 33759 13887 33793
rect 13769 33725 13887 33759
rect 13769 33691 13809 33725
rect 13843 33691 13887 33725
rect 13769 33657 13887 33691
rect 13769 33623 13809 33657
rect 13843 33623 13887 33657
rect 13769 33589 13887 33623
rect 13769 33555 13809 33589
rect 13843 33555 13887 33589
rect 13769 33521 13887 33555
rect 13769 33487 13809 33521
rect 13843 33487 13887 33521
rect 13769 33453 13887 33487
rect 13769 33419 13809 33453
rect 13843 33419 13887 33453
rect 13769 33385 13887 33419
rect 13769 33351 13809 33385
rect 13843 33351 13887 33385
rect 13769 33317 13887 33351
rect 13769 33283 13809 33317
rect 13843 33283 13887 33317
rect 13769 33249 13887 33283
rect 13769 33215 13809 33249
rect 13843 33215 13887 33249
rect 13769 33181 13887 33215
rect 13769 33147 13809 33181
rect 13843 33147 13887 33181
rect 13769 33113 13887 33147
rect 13769 33079 13809 33113
rect 13843 33079 13887 33113
rect 13769 33045 13887 33079
rect 13769 33011 13809 33045
rect 13843 33011 13887 33045
rect 13769 32977 13887 33011
rect 13769 32943 13809 32977
rect 13843 32943 13887 32977
rect 13769 32909 13887 32943
rect 13769 32875 13809 32909
rect 13843 32875 13887 32909
rect 13769 32841 13887 32875
rect 13769 32807 13809 32841
rect 13843 32807 13887 32841
rect 13769 32773 13887 32807
rect 13769 32739 13809 32773
rect 13843 32739 13887 32773
rect 13769 32705 13887 32739
rect 13769 32671 13809 32705
rect 13843 32671 13887 32705
rect 13769 32637 13887 32671
rect 13769 32603 13809 32637
rect 13843 32603 13887 32637
rect 13769 32569 13887 32603
rect 13769 32535 13809 32569
rect 13843 32535 13887 32569
rect 13769 32501 13887 32535
rect 13769 32467 13809 32501
rect 13843 32467 13887 32501
rect 13769 32433 13887 32467
rect 13769 32399 13809 32433
rect 13843 32399 13887 32433
rect 13769 32365 13887 32399
rect 13769 32331 13809 32365
rect 13843 32331 13887 32365
rect 13769 32297 13887 32331
rect 13769 32263 13809 32297
rect 13843 32263 13887 32297
rect 13769 32229 13887 32263
rect 13769 32195 13809 32229
rect 13843 32195 13887 32229
rect 13769 32161 13887 32195
rect 13769 32127 13809 32161
rect 13843 32127 13887 32161
rect 13769 32093 13887 32127
rect 13769 32059 13809 32093
rect 13843 32059 13887 32093
rect 13769 32025 13887 32059
rect 13769 31991 13809 32025
rect 13843 31991 13887 32025
rect 13769 31957 13887 31991
rect 13769 31923 13809 31957
rect 13843 31923 13887 31957
rect 13769 31889 13887 31923
rect 13769 31855 13809 31889
rect 13843 31855 13887 31889
rect 13769 31821 13887 31855
rect 13769 31787 13809 31821
rect 13843 31787 13887 31821
rect 13769 31753 13887 31787
rect 13769 31719 13809 31753
rect 13843 31719 13887 31753
rect 13769 31685 13887 31719
rect 13769 31651 13809 31685
rect 13843 31651 13887 31685
rect 13769 31617 13887 31651
rect 13769 31583 13809 31617
rect 13843 31583 13887 31617
rect 13769 31549 13887 31583
rect 13769 31515 13809 31549
rect 13843 31515 13887 31549
rect 13769 31481 13887 31515
rect 13769 31447 13809 31481
rect 13843 31447 13887 31481
rect 13769 31413 13887 31447
rect 13769 31379 13809 31413
rect 13843 31379 13887 31413
rect 13769 31345 13887 31379
rect 13769 31311 13809 31345
rect 13843 31311 13887 31345
rect 13769 31277 13887 31311
rect 13769 31243 13809 31277
rect 13843 31243 13887 31277
rect 13769 31209 13887 31243
rect 13769 31175 13809 31209
rect 13843 31175 13887 31209
rect 13769 31141 13887 31175
rect 13769 31107 13809 31141
rect 13843 31107 13887 31141
rect 13769 31073 13887 31107
rect 13769 31039 13809 31073
rect 13843 31039 13887 31073
rect 13769 31005 13887 31039
rect 13769 30971 13809 31005
rect 13843 30971 13887 31005
rect 13769 30937 13887 30971
rect 13769 30903 13809 30937
rect 13843 30903 13887 30937
rect 13769 30869 13887 30903
rect 13769 30835 13809 30869
rect 13843 30835 13887 30869
rect 13769 30801 13887 30835
rect 13769 30767 13809 30801
rect 13843 30767 13887 30801
rect 13769 30733 13887 30767
rect 13769 30699 13809 30733
rect 13843 30699 13887 30733
rect 13769 30665 13887 30699
rect 13769 30631 13809 30665
rect 13843 30631 13887 30665
rect 13769 30597 13887 30631
rect 13769 30563 13809 30597
rect 13843 30563 13887 30597
rect 13769 30529 13887 30563
rect 13769 30495 13809 30529
rect 13843 30495 13887 30529
rect 13769 30461 13887 30495
rect 13769 30427 13809 30461
rect 13843 30427 13887 30461
rect 13769 30393 13887 30427
rect 13769 30359 13809 30393
rect 13843 30359 13887 30393
rect 13769 30325 13887 30359
rect 13769 30291 13809 30325
rect 13843 30291 13887 30325
rect 13769 30257 13887 30291
rect 13769 30223 13809 30257
rect 13843 30223 13887 30257
rect 13769 30189 13887 30223
rect 13769 30155 13809 30189
rect 13843 30155 13887 30189
rect 13769 30121 13887 30155
rect 13769 30087 13809 30121
rect 13843 30087 13887 30121
rect 13769 30053 13887 30087
rect 13769 30019 13809 30053
rect 13843 30019 13887 30053
rect 13769 29985 13887 30019
rect 13769 29951 13809 29985
rect 13843 29951 13887 29985
rect 13769 29917 13887 29951
rect 13769 29883 13809 29917
rect 13843 29883 13887 29917
rect 13769 29849 13887 29883
rect 13769 29815 13809 29849
rect 13843 29815 13887 29849
rect 13769 29781 13887 29815
rect 13769 29747 13809 29781
rect 13843 29747 13887 29781
rect 13769 29713 13887 29747
rect 13769 29679 13809 29713
rect 13843 29679 13887 29713
rect 13769 29645 13887 29679
rect 13769 29611 13809 29645
rect 13843 29611 13887 29645
rect 13769 29577 13887 29611
rect 13769 29543 13809 29577
rect 13843 29543 13887 29577
rect 13769 29509 13887 29543
rect 13769 29475 13809 29509
rect 13843 29475 13887 29509
rect 13769 29441 13887 29475
rect 13769 29407 13809 29441
rect 13843 29407 13887 29441
rect 13769 29373 13887 29407
rect 13769 29339 13809 29373
rect 13843 29339 13887 29373
rect 13769 29305 13887 29339
rect 13769 29271 13809 29305
rect 13843 29271 13887 29305
rect 13769 29237 13887 29271
rect 13769 29203 13809 29237
rect 13843 29203 13887 29237
rect 13769 29169 13887 29203
rect 13769 29135 13809 29169
rect 13843 29135 13887 29169
rect 13769 29101 13887 29135
rect 13769 29067 13809 29101
rect 13843 29067 13887 29101
rect 13769 29033 13887 29067
rect 13769 28999 13809 29033
rect 13843 28999 13887 29033
rect 13769 28965 13887 28999
rect 13769 28931 13809 28965
rect 13843 28931 13887 28965
rect 1119 28868 1161 28902
rect 1195 28868 1237 28902
rect 1119 28834 1237 28868
rect 1119 28800 1161 28834
rect 1195 28800 1237 28834
rect 1119 28766 1237 28800
rect 1119 28732 1161 28766
rect 1195 28732 1237 28766
rect 1119 28698 1237 28732
rect 1119 28664 1161 28698
rect 1195 28664 1237 28698
rect 1119 28630 1237 28664
rect 1119 28596 1161 28630
rect 1195 28596 1237 28630
rect 1119 28562 1237 28596
rect 1119 28528 1161 28562
rect 1195 28528 1237 28562
rect 1119 28494 1237 28528
rect 1119 28460 1161 28494
rect 1195 28460 1237 28494
rect 1119 28426 1237 28460
rect 1119 28392 1161 28426
rect 1195 28392 1237 28426
rect 1119 28358 1237 28392
rect 1119 28324 1161 28358
rect 1195 28324 1237 28358
rect 1119 28290 1237 28324
rect 1119 28256 1161 28290
rect 1195 28256 1237 28290
rect 1119 28222 1237 28256
rect 1119 28188 1161 28222
rect 1195 28188 1237 28222
rect 1119 28154 1237 28188
rect 1119 28120 1161 28154
rect 1195 28120 1237 28154
rect 1119 28086 1237 28120
rect 1119 28052 1161 28086
rect 1195 28052 1237 28086
rect 1119 28018 1237 28052
rect 1119 27984 1161 28018
rect 1195 27984 1237 28018
rect 1119 27950 1237 27984
rect 1119 27916 1161 27950
rect 1195 27916 1237 27950
rect 1119 27882 1237 27916
rect 1119 27848 1161 27882
rect 1195 27848 1237 27882
rect 1119 27814 1237 27848
rect 1119 27780 1161 27814
rect 1195 27780 1237 27814
rect 1119 27746 1237 27780
rect 1119 27712 1161 27746
rect 1195 27712 1237 27746
rect 1119 27678 1237 27712
rect 1119 27644 1161 27678
rect 1195 27644 1237 27678
rect 1119 27610 1237 27644
rect 1119 27576 1161 27610
rect 1195 27576 1237 27610
rect 1119 27542 1237 27576
rect 1119 27508 1161 27542
rect 1195 27508 1237 27542
rect 1119 27474 1237 27508
rect 1119 27440 1161 27474
rect 1195 27440 1237 27474
rect 1119 27406 1237 27440
rect 1119 27372 1161 27406
rect 1195 27372 1237 27406
rect 1119 27338 1237 27372
rect 1119 27304 1161 27338
rect 1195 27304 1237 27338
rect 1119 27270 1237 27304
rect 1119 27236 1161 27270
rect 1195 27236 1237 27270
rect 1119 27202 1237 27236
rect 1119 27168 1161 27202
rect 1195 27168 1237 27202
rect 1119 27134 1237 27168
rect 1119 27100 1161 27134
rect 1195 27100 1237 27134
rect 1119 27066 1237 27100
rect 1119 27032 1161 27066
rect 1195 27032 1237 27066
rect 1119 26998 1237 27032
rect 13769 28897 13887 28931
rect 13769 28863 13809 28897
rect 13843 28863 13887 28897
rect 13769 28829 13887 28863
rect 13769 28795 13809 28829
rect 13843 28795 13887 28829
rect 13769 28761 13887 28795
rect 13769 28727 13809 28761
rect 13843 28727 13887 28761
rect 13769 28693 13887 28727
rect 13769 28659 13809 28693
rect 13843 28659 13887 28693
rect 13769 28625 13887 28659
rect 13769 28591 13809 28625
rect 13843 28591 13887 28625
rect 13769 28557 13887 28591
rect 13769 28523 13809 28557
rect 13843 28523 13887 28557
rect 13769 28489 13887 28523
rect 13769 28455 13809 28489
rect 13843 28455 13887 28489
rect 13769 28421 13887 28455
rect 13769 28387 13809 28421
rect 13843 28387 13887 28421
rect 13769 28353 13887 28387
rect 13769 28319 13809 28353
rect 13843 28319 13887 28353
rect 13769 28285 13887 28319
rect 13769 28251 13809 28285
rect 13843 28251 13887 28285
rect 13769 28217 13887 28251
rect 13769 28183 13809 28217
rect 13843 28183 13887 28217
rect 13769 28149 13887 28183
rect 13769 28115 13809 28149
rect 13843 28115 13887 28149
rect 13769 28081 13887 28115
rect 13769 28047 13809 28081
rect 13843 28047 13887 28081
rect 13769 28013 13887 28047
rect 13769 27979 13809 28013
rect 13843 27979 13887 28013
rect 13769 27945 13887 27979
rect 13769 27911 13809 27945
rect 13843 27911 13887 27945
rect 13769 27877 13887 27911
rect 13769 27843 13809 27877
rect 13843 27843 13887 27877
rect 13769 27809 13887 27843
rect 13769 27775 13809 27809
rect 13843 27775 13887 27809
rect 13769 27741 13887 27775
rect 13769 27707 13809 27741
rect 13843 27707 13887 27741
rect 13769 27673 13887 27707
rect 13769 27639 13809 27673
rect 13843 27639 13887 27673
rect 13769 27605 13887 27639
rect 13769 27571 13809 27605
rect 13843 27571 13887 27605
rect 13769 27537 13887 27571
rect 13769 27503 13809 27537
rect 13843 27503 13887 27537
rect 13769 27469 13887 27503
rect 13769 27435 13809 27469
rect 13843 27435 13887 27469
rect 13769 27401 13887 27435
rect 13769 27367 13809 27401
rect 13843 27367 13887 27401
rect 13769 27333 13887 27367
rect 13769 27299 13809 27333
rect 13843 27299 13887 27333
rect 13769 27265 13887 27299
rect 13769 27231 13809 27265
rect 13843 27231 13887 27265
rect 13769 27197 13887 27231
rect 13769 27163 13809 27197
rect 13843 27163 13887 27197
rect 13769 27129 13887 27163
rect 13769 27095 13809 27129
rect 13843 27095 13887 27129
rect 13769 27061 13887 27095
rect 13769 27027 13809 27061
rect 13843 27027 13887 27061
rect 1119 26964 1161 26998
rect 1195 26964 1237 26998
rect 1119 26930 1237 26964
rect 1119 26896 1161 26930
rect 1195 26896 1237 26930
rect 1119 26862 1237 26896
rect 1119 26828 1161 26862
rect 1195 26828 1237 26862
rect 1119 26794 1237 26828
rect 1119 26760 1161 26794
rect 1195 26760 1237 26794
rect 1119 26726 1237 26760
rect 1119 26692 1161 26726
rect 1195 26692 1237 26726
rect 1119 26658 1237 26692
rect 1119 26624 1161 26658
rect 1195 26624 1237 26658
rect 1119 26590 1237 26624
rect 1119 26556 1161 26590
rect 1195 26556 1237 26590
rect 1119 26522 1237 26556
rect 1119 26488 1161 26522
rect 1195 26488 1237 26522
rect 1119 26454 1237 26488
rect 1119 26420 1161 26454
rect 1195 26420 1237 26454
rect 1119 26386 1237 26420
rect 1119 26352 1161 26386
rect 1195 26352 1237 26386
rect 1119 26318 1237 26352
rect 1119 26284 1161 26318
rect 1195 26284 1237 26318
rect 1119 26250 1237 26284
rect 1119 26216 1161 26250
rect 1195 26216 1237 26250
rect 1119 26182 1237 26216
rect 1119 26148 1161 26182
rect 1195 26148 1237 26182
rect 1119 26114 1237 26148
rect 1119 26080 1161 26114
rect 1195 26080 1237 26114
rect 1119 26046 1237 26080
rect 1119 26012 1161 26046
rect 1195 26012 1237 26046
rect 1119 25978 1237 26012
rect 1119 25944 1161 25978
rect 1195 25944 1237 25978
rect 1119 25910 1237 25944
rect 1119 25876 1161 25910
rect 1195 25876 1237 25910
rect 1119 25842 1237 25876
rect 1119 25808 1161 25842
rect 1195 25808 1237 25842
rect 1119 25774 1237 25808
rect 1119 25740 1161 25774
rect 1195 25740 1237 25774
rect 1119 25706 1237 25740
rect 1119 25672 1161 25706
rect 1195 25672 1237 25706
rect 1119 25638 1237 25672
rect 1119 25604 1161 25638
rect 1195 25604 1237 25638
rect 1119 25570 1237 25604
rect 1119 25536 1161 25570
rect 1195 25536 1237 25570
rect 1119 25502 1237 25536
rect 1119 25468 1161 25502
rect 1195 25468 1237 25502
rect 1119 25434 1237 25468
rect 1119 25400 1161 25434
rect 1195 25400 1237 25434
rect 1119 25366 1237 25400
rect 1119 25332 1161 25366
rect 1195 25332 1237 25366
rect 1119 25298 1237 25332
rect 1119 25264 1161 25298
rect 1195 25264 1237 25298
rect 1119 25230 1237 25264
rect 1119 25196 1161 25230
rect 1195 25196 1237 25230
rect 1119 25162 1237 25196
rect 1119 25128 1161 25162
rect 1195 25128 1237 25162
rect 1119 25094 1237 25128
rect 1119 25060 1161 25094
rect 1195 25060 1237 25094
rect 1119 25026 1237 25060
rect 1119 24992 1161 25026
rect 1195 24992 1237 25026
rect 1119 24958 1237 24992
rect 1119 24924 1161 24958
rect 1195 24924 1237 24958
rect 1119 24890 1237 24924
rect 1119 24856 1161 24890
rect 1195 24856 1237 24890
rect 1119 24822 1237 24856
rect 1119 24788 1161 24822
rect 1195 24788 1237 24822
rect 1119 24754 1237 24788
rect 1119 24720 1161 24754
rect 1195 24720 1237 24754
rect 1119 24686 1237 24720
rect 1119 24652 1161 24686
rect 1195 24652 1237 24686
rect 1119 24618 1237 24652
rect 1119 24584 1161 24618
rect 1195 24584 1237 24618
rect 1119 24550 1237 24584
rect 1119 24516 1161 24550
rect 1195 24516 1237 24550
rect 1119 24482 1237 24516
rect 1119 24448 1161 24482
rect 1195 24448 1237 24482
rect 1119 24414 1237 24448
rect 1119 24380 1161 24414
rect 1195 24380 1237 24414
rect 1119 24346 1237 24380
rect 1119 24312 1161 24346
rect 1195 24312 1237 24346
rect 1119 24278 1237 24312
rect 1119 24244 1161 24278
rect 1195 24244 1237 24278
rect 1119 24210 1237 24244
rect 1119 24176 1161 24210
rect 1195 24176 1237 24210
rect 1119 24142 1237 24176
rect 1119 24108 1161 24142
rect 1195 24108 1237 24142
rect 1119 24074 1237 24108
rect 1119 24040 1161 24074
rect 1195 24040 1237 24074
rect 1119 24006 1237 24040
rect 1119 23972 1161 24006
rect 1195 23972 1237 24006
rect 1119 23938 1237 23972
rect 1119 23904 1161 23938
rect 1195 23904 1237 23938
rect 1119 23870 1237 23904
rect 1119 23836 1161 23870
rect 1195 23836 1237 23870
rect 1119 23802 1237 23836
rect 1119 23768 1161 23802
rect 1195 23768 1237 23802
rect 1119 23734 1237 23768
rect 1119 23700 1161 23734
rect 1195 23700 1237 23734
rect 1119 23666 1237 23700
rect 1119 23632 1161 23666
rect 1195 23632 1237 23666
rect 1119 23598 1237 23632
rect 1119 23564 1161 23598
rect 1195 23564 1237 23598
rect 1119 23530 1237 23564
rect 1119 23496 1161 23530
rect 1195 23496 1237 23530
rect 1119 23462 1237 23496
rect 1119 23428 1161 23462
rect 1195 23428 1237 23462
rect 1119 23394 1237 23428
rect 1119 23360 1161 23394
rect 1195 23360 1237 23394
rect 1119 23326 1237 23360
rect 1119 23292 1161 23326
rect 1195 23292 1237 23326
rect 1119 23258 1237 23292
rect 1119 23224 1161 23258
rect 1195 23224 1237 23258
rect 1119 23190 1237 23224
rect 1119 23156 1161 23190
rect 1195 23156 1237 23190
rect 1119 23122 1237 23156
rect 1119 23088 1161 23122
rect 1195 23088 1237 23122
rect 1119 23054 1237 23088
rect 1119 23020 1161 23054
rect 1195 23020 1237 23054
rect 1119 22986 1237 23020
rect 1119 22952 1161 22986
rect 1195 22952 1237 22986
rect 1119 22918 1237 22952
rect 1119 22884 1161 22918
rect 1195 22884 1237 22918
rect 1119 22850 1237 22884
rect 1119 22816 1161 22850
rect 1195 22816 1237 22850
rect 1119 22782 1237 22816
rect 1119 22748 1161 22782
rect 1195 22748 1237 22782
rect 1119 22714 1237 22748
rect 1119 22680 1161 22714
rect 1195 22680 1237 22714
rect 1119 22646 1237 22680
rect 1119 22612 1161 22646
rect 1195 22612 1237 22646
rect 1119 22578 1237 22612
rect 1119 22544 1161 22578
rect 1195 22544 1237 22578
rect 1119 22510 1237 22544
rect 1119 22476 1161 22510
rect 1195 22476 1237 22510
rect 1119 22442 1237 22476
rect 1119 22408 1161 22442
rect 1195 22408 1237 22442
rect 1119 22374 1237 22408
rect 1119 22340 1161 22374
rect 1195 22340 1237 22374
rect 1119 22306 1237 22340
rect 1119 22272 1161 22306
rect 1195 22272 1237 22306
rect 1119 22238 1237 22272
rect 1119 22204 1161 22238
rect 1195 22204 1237 22238
rect 1119 22170 1237 22204
rect 1119 22136 1161 22170
rect 1195 22136 1237 22170
rect 1119 22102 1237 22136
rect 1119 22068 1161 22102
rect 1195 22068 1237 22102
rect 1119 22034 1237 22068
rect 1119 22000 1161 22034
rect 1195 22000 1237 22034
rect 1119 21966 1237 22000
rect 1119 21932 1161 21966
rect 1195 21932 1237 21966
rect 1119 21898 1237 21932
rect 1119 21864 1161 21898
rect 1195 21864 1237 21898
rect 1119 21830 1237 21864
rect 1119 21796 1161 21830
rect 1195 21796 1237 21830
rect 1119 21762 1237 21796
rect 1119 21728 1161 21762
rect 1195 21728 1237 21762
rect 1119 21694 1237 21728
rect 1119 21660 1161 21694
rect 1195 21660 1237 21694
rect 1119 21626 1237 21660
rect 1119 21592 1161 21626
rect 1195 21592 1237 21626
rect 1119 21558 1237 21592
rect 1119 21524 1161 21558
rect 1195 21524 1237 21558
rect 1119 21490 1237 21524
rect 1119 21456 1161 21490
rect 1195 21456 1237 21490
rect 1119 21422 1237 21456
rect 1119 21388 1161 21422
rect 1195 21388 1237 21422
rect 1119 21354 1237 21388
rect 1119 21320 1161 21354
rect 1195 21320 1237 21354
rect 1119 21286 1237 21320
rect 1119 21252 1161 21286
rect 1195 21252 1237 21286
rect 1119 21218 1237 21252
rect 1119 21184 1161 21218
rect 1195 21184 1237 21218
rect 1119 21150 1237 21184
rect 1119 21116 1161 21150
rect 1195 21116 1237 21150
rect 1119 21082 1237 21116
rect 1119 21048 1161 21082
rect 1195 21048 1237 21082
rect 1119 21014 1237 21048
rect 1119 20980 1161 21014
rect 1195 20980 1237 21014
rect 1119 20946 1237 20980
rect 1119 20912 1161 20946
rect 1195 20912 1237 20946
rect 1119 20878 1237 20912
rect 1119 20844 1161 20878
rect 1195 20844 1237 20878
rect 1119 20810 1237 20844
rect 1119 20776 1161 20810
rect 1195 20776 1237 20810
rect 1119 20742 1237 20776
rect 1119 20708 1161 20742
rect 1195 20708 1237 20742
rect 1119 20674 1237 20708
rect 1119 20640 1161 20674
rect 1195 20640 1237 20674
rect 1119 20606 1237 20640
rect 1119 20572 1161 20606
rect 1195 20572 1237 20606
rect 1119 20538 1237 20572
rect 1119 20504 1161 20538
rect 1195 20504 1237 20538
rect 1119 20470 1237 20504
rect 1119 20436 1161 20470
rect 1195 20436 1237 20470
rect 1119 20402 1237 20436
rect 1119 20368 1161 20402
rect 1195 20368 1237 20402
rect 1119 20334 1237 20368
rect 1119 20300 1161 20334
rect 1195 20300 1237 20334
rect 1119 20266 1237 20300
rect 1119 20232 1161 20266
rect 1195 20232 1237 20266
rect 1119 20198 1237 20232
rect 1119 20164 1161 20198
rect 1195 20164 1237 20198
rect 1119 20130 1237 20164
rect 1119 20096 1161 20130
rect 1195 20096 1237 20130
rect 1119 20062 1237 20096
rect 1119 20028 1161 20062
rect 1195 20028 1237 20062
rect 1119 19994 1237 20028
rect 1119 19960 1161 19994
rect 1195 19960 1237 19994
rect 1119 19926 1237 19960
rect 1119 19892 1161 19926
rect 1195 19892 1237 19926
rect 1119 19858 1237 19892
rect 1119 19824 1161 19858
rect 1195 19824 1237 19858
rect 1119 19790 1237 19824
rect 1119 19756 1161 19790
rect 1195 19756 1237 19790
rect 1119 19722 1237 19756
rect 1119 19688 1161 19722
rect 1195 19688 1237 19722
rect 1119 19654 1237 19688
rect 1119 19620 1161 19654
rect 1195 19620 1237 19654
rect 1119 19586 1237 19620
rect 1119 19552 1161 19586
rect 1195 19552 1237 19586
rect 1119 19518 1237 19552
rect 1119 19484 1161 19518
rect 1195 19484 1237 19518
rect 1119 19450 1237 19484
rect 1119 19416 1161 19450
rect 1195 19416 1237 19450
rect 1119 19382 1237 19416
rect 1119 19348 1161 19382
rect 1195 19348 1237 19382
rect 1119 19314 1237 19348
rect 1119 19280 1161 19314
rect 1195 19280 1237 19314
rect 1119 19246 1237 19280
rect 1119 19212 1161 19246
rect 1195 19212 1237 19246
rect 1119 19178 1237 19212
rect 1119 19144 1161 19178
rect 1195 19144 1237 19178
rect 1119 19110 1237 19144
rect 1119 19076 1161 19110
rect 1195 19076 1237 19110
rect 1119 19042 1237 19076
rect 1119 19008 1161 19042
rect 1195 19008 1237 19042
rect 1119 18974 1237 19008
rect 1119 18940 1161 18974
rect 1195 18940 1237 18974
rect 1119 18906 1237 18940
rect 1119 18872 1161 18906
rect 1195 18872 1237 18906
rect 1119 18838 1237 18872
rect 1119 18804 1161 18838
rect 1195 18804 1237 18838
rect 1119 18770 1237 18804
rect 1119 18736 1161 18770
rect 1195 18736 1237 18770
rect 1119 18702 1237 18736
rect 1119 18668 1161 18702
rect 1195 18668 1237 18702
rect 1119 18634 1237 18668
rect 1119 18600 1161 18634
rect 1195 18600 1237 18634
rect 1119 18566 1237 18600
rect 1119 18532 1161 18566
rect 1195 18532 1237 18566
rect 1119 18498 1237 18532
rect 1119 18464 1161 18498
rect 1195 18464 1237 18498
rect 1119 18430 1237 18464
rect 1119 18396 1161 18430
rect 1195 18396 1237 18430
rect 1119 18362 1237 18396
rect 1119 18328 1161 18362
rect 1195 18328 1237 18362
rect 1119 18294 1237 18328
rect 1119 18260 1161 18294
rect 1195 18260 1237 18294
rect 1119 18226 1237 18260
rect 1119 18192 1161 18226
rect 1195 18192 1237 18226
rect 1119 18158 1237 18192
rect 1119 18124 1161 18158
rect 1195 18124 1237 18158
rect 1119 18090 1237 18124
rect 1119 18056 1161 18090
rect 1195 18056 1237 18090
rect 1119 18022 1237 18056
rect 1119 17988 1161 18022
rect 1195 17988 1237 18022
rect 1119 17954 1237 17988
rect 1119 17920 1161 17954
rect 1195 17920 1237 17954
rect 1119 17886 1237 17920
rect 1119 17852 1161 17886
rect 1195 17852 1237 17886
rect 1119 17818 1237 17852
rect 1119 17784 1161 17818
rect 1195 17784 1237 17818
rect 1119 17750 1237 17784
rect 1119 17716 1161 17750
rect 1195 17716 1237 17750
rect 1119 17682 1237 17716
rect 1119 17648 1161 17682
rect 1195 17648 1237 17682
rect 1119 17614 1237 17648
rect 1119 17580 1161 17614
rect 1195 17580 1237 17614
rect 1119 17546 1237 17580
rect 1119 17512 1161 17546
rect 1195 17512 1237 17546
rect 1119 17478 1237 17512
rect 1119 17444 1161 17478
rect 1195 17444 1237 17478
rect 1119 17410 1237 17444
rect 1119 17376 1161 17410
rect 1195 17376 1237 17410
rect 1119 17342 1237 17376
rect 1119 17308 1161 17342
rect 1195 17308 1237 17342
rect 1119 17274 1237 17308
rect 1119 17240 1161 17274
rect 1195 17240 1237 17274
rect 1119 17206 1237 17240
rect 1119 17172 1161 17206
rect 1195 17172 1237 17206
rect 1119 17138 1237 17172
rect 1119 17104 1161 17138
rect 1195 17104 1237 17138
rect 1119 17070 1237 17104
rect 1119 17036 1161 17070
rect 1195 17036 1237 17070
rect 1119 17002 1237 17036
rect 1119 16968 1161 17002
rect 1195 16968 1237 17002
rect 1119 16934 1237 16968
rect 1119 16900 1161 16934
rect 1195 16900 1237 16934
rect 1119 16866 1237 16900
rect 1119 16832 1161 16866
rect 1195 16832 1237 16866
rect 1119 16798 1237 16832
rect 1119 16764 1161 16798
rect 1195 16764 1237 16798
rect 1119 16730 1237 16764
rect 1119 16696 1161 16730
rect 1195 16696 1237 16730
rect 1119 16662 1237 16696
rect 1119 16628 1161 16662
rect 1195 16628 1237 16662
rect 1119 16594 1237 16628
rect 1119 16560 1161 16594
rect 1195 16560 1237 16594
rect 1119 16526 1237 16560
rect 1119 16492 1161 16526
rect 1195 16492 1237 16526
rect 1119 16458 1237 16492
rect 1119 16424 1161 16458
rect 1195 16424 1237 16458
rect 1119 16390 1237 16424
rect 1119 16356 1161 16390
rect 1195 16356 1237 16390
rect 1119 16322 1237 16356
rect 1119 16288 1161 16322
rect 1195 16288 1237 16322
rect 1119 16254 1237 16288
rect 1119 16220 1161 16254
rect 1195 16220 1237 16254
rect 1119 16186 1237 16220
rect 1119 16152 1161 16186
rect 1195 16152 1237 16186
rect 1119 16118 1237 16152
rect 1119 16084 1161 16118
rect 1195 16084 1237 16118
rect 1119 16050 1237 16084
rect 1119 16016 1161 16050
rect 1195 16016 1237 16050
rect 1119 15982 1237 16016
rect 1119 15948 1161 15982
rect 1195 15948 1237 15982
rect 1119 15914 1237 15948
rect 1119 15880 1161 15914
rect 1195 15880 1237 15914
rect 1119 15846 1237 15880
rect 1119 15812 1161 15846
rect 1195 15812 1237 15846
rect 1119 15778 1237 15812
rect 1119 15744 1161 15778
rect 1195 15744 1237 15778
rect 1119 15710 1237 15744
rect 1119 15676 1161 15710
rect 1195 15676 1237 15710
rect 1119 15642 1237 15676
rect 1119 15608 1161 15642
rect 1195 15608 1237 15642
rect 1119 15574 1237 15608
rect 1119 15540 1161 15574
rect 1195 15540 1237 15574
rect 1119 15506 1237 15540
rect 1119 15472 1161 15506
rect 1195 15472 1237 15506
rect 1119 15438 1237 15472
rect 1119 15404 1161 15438
rect 1195 15404 1237 15438
rect 1119 15370 1237 15404
rect 1119 15336 1161 15370
rect 1195 15336 1237 15370
rect 1119 15302 1237 15336
rect 1119 15268 1161 15302
rect 1195 15268 1237 15302
rect 1119 15234 1237 15268
rect 1119 15200 1161 15234
rect 1195 15200 1237 15234
rect 1119 15166 1237 15200
rect 1119 15132 1161 15166
rect 1195 15132 1237 15166
rect 1119 15098 1237 15132
rect 1119 15064 1161 15098
rect 1195 15064 1237 15098
rect 1119 15030 1237 15064
rect 1119 14996 1161 15030
rect 1195 14996 1237 15030
rect 1119 14962 1237 14996
rect 1119 14928 1161 14962
rect 1195 14928 1237 14962
rect 1119 14894 1237 14928
rect 1119 14860 1161 14894
rect 1195 14860 1237 14894
rect 1119 14826 1237 14860
rect 1119 14792 1161 14826
rect 1195 14792 1237 14826
rect 1119 14758 1237 14792
rect 1119 14724 1161 14758
rect 1195 14724 1237 14758
rect 1119 14690 1237 14724
rect 1119 14656 1161 14690
rect 1195 14656 1237 14690
rect 1119 14622 1237 14656
rect 1119 14588 1161 14622
rect 1195 14588 1237 14622
rect 1119 14554 1237 14588
rect 1119 14520 1161 14554
rect 1195 14520 1237 14554
rect 1119 14486 1237 14520
rect 1119 14452 1161 14486
rect 1195 14452 1237 14486
rect 1119 14418 1237 14452
rect 1119 14384 1161 14418
rect 1195 14384 1237 14418
rect 1119 14350 1237 14384
rect 1119 14316 1161 14350
rect 1195 14316 1237 14350
rect 1119 14282 1237 14316
rect 1119 14248 1161 14282
rect 1195 14248 1237 14282
rect 1119 14214 1237 14248
rect 1119 14180 1161 14214
rect 1195 14180 1237 14214
rect 1119 14146 1237 14180
rect 1119 14112 1161 14146
rect 1195 14112 1237 14146
rect 1119 14078 1237 14112
rect 1119 14044 1161 14078
rect 1195 14044 1237 14078
rect 1119 14010 1237 14044
rect 1119 13976 1161 14010
rect 1195 13976 1237 14010
rect 1119 13942 1237 13976
rect 1119 13908 1161 13942
rect 1195 13908 1237 13942
rect 1119 13874 1237 13908
rect 1119 13840 1161 13874
rect 1195 13840 1237 13874
rect 1119 13806 1237 13840
rect 1119 13772 1161 13806
rect 1195 13772 1237 13806
rect 1119 13738 1237 13772
rect 1119 13704 1161 13738
rect 1195 13704 1237 13738
rect 1119 13670 1237 13704
rect 1119 13636 1161 13670
rect 1195 13636 1237 13670
rect 1119 13602 1237 13636
rect 1119 13568 1161 13602
rect 1195 13568 1237 13602
rect 1119 13534 1237 13568
rect 1119 13500 1161 13534
rect 1195 13500 1237 13534
rect 1119 13466 1237 13500
rect 1119 13432 1161 13466
rect 1195 13432 1237 13466
rect 1119 13398 1237 13432
rect 1119 13364 1161 13398
rect 1195 13364 1237 13398
rect 1119 13330 1237 13364
rect 1119 13296 1161 13330
rect 1195 13296 1237 13330
rect 1119 13262 1237 13296
rect 1119 13228 1161 13262
rect 1195 13228 1237 13262
rect 1119 13194 1237 13228
rect 1119 13160 1161 13194
rect 1195 13160 1237 13194
rect 1119 13126 1237 13160
rect 1119 13092 1161 13126
rect 1195 13092 1237 13126
rect 1119 13058 1237 13092
rect 1119 13024 1161 13058
rect 1195 13024 1237 13058
rect 1119 12990 1237 13024
rect 1119 12956 1161 12990
rect 1195 12956 1237 12990
rect 1119 12922 1237 12956
rect 1119 12888 1161 12922
rect 1195 12888 1237 12922
rect 1119 12854 1237 12888
rect 1119 12820 1161 12854
rect 1195 12820 1237 12854
rect 1119 12786 1237 12820
rect 1119 12752 1161 12786
rect 1195 12752 1237 12786
rect 1119 12718 1237 12752
rect 1119 12684 1161 12718
rect 1195 12684 1237 12718
rect 1119 12650 1237 12684
rect 1119 12616 1161 12650
rect 1195 12616 1237 12650
rect 1119 12582 1237 12616
rect 1119 12548 1161 12582
rect 1195 12548 1237 12582
rect 1119 12514 1237 12548
rect 1119 12480 1161 12514
rect 1195 12480 1237 12514
rect 1119 12446 1237 12480
rect 1119 12412 1161 12446
rect 1195 12412 1237 12446
rect 1119 12378 1237 12412
rect 1119 12344 1161 12378
rect 1195 12344 1237 12378
rect 1119 12310 1237 12344
rect 1119 12276 1161 12310
rect 1195 12276 1237 12310
rect 1119 12242 1237 12276
rect 1119 12208 1161 12242
rect 1195 12208 1237 12242
rect 1119 12174 1237 12208
rect 1119 12140 1161 12174
rect 1195 12140 1237 12174
rect 1119 12106 1237 12140
rect 1119 12072 1161 12106
rect 1195 12072 1237 12106
rect 1119 12038 1237 12072
rect 1119 12004 1161 12038
rect 1195 12004 1237 12038
rect 1119 11970 1237 12004
rect 1119 11936 1161 11970
rect 1195 11936 1237 11970
rect 1119 11902 1237 11936
rect 1119 11868 1161 11902
rect 1195 11868 1237 11902
rect 1119 11834 1237 11868
rect 1119 11800 1161 11834
rect 1195 11800 1237 11834
rect 1119 11766 1237 11800
rect 1119 11732 1161 11766
rect 1195 11732 1237 11766
rect 1119 11698 1237 11732
rect 1119 11664 1161 11698
rect 1195 11664 1237 11698
rect 1119 11630 1237 11664
rect 1119 11596 1161 11630
rect 1195 11596 1237 11630
rect 1119 11562 1237 11596
rect 1119 11528 1161 11562
rect 1195 11528 1237 11562
rect 1119 11494 1237 11528
rect 1119 11460 1161 11494
rect 1195 11460 1237 11494
rect 1119 11426 1237 11460
rect 1119 11392 1161 11426
rect 1195 11392 1237 11426
rect 1119 11358 1237 11392
rect 1119 11324 1161 11358
rect 1195 11324 1237 11358
rect 1119 11290 1237 11324
rect 1119 11256 1161 11290
rect 1195 11256 1237 11290
rect 1119 11222 1237 11256
rect 1119 11188 1161 11222
rect 1195 11188 1237 11222
rect 1119 11154 1237 11188
rect 1119 11120 1161 11154
rect 1195 11120 1237 11154
rect 1119 11086 1237 11120
rect 1119 11052 1161 11086
rect 1195 11052 1237 11086
rect 1119 11018 1237 11052
rect 1119 10984 1161 11018
rect 1195 10984 1237 11018
rect 1119 10950 1237 10984
rect 1119 10916 1161 10950
rect 1195 10916 1237 10950
rect 1119 10882 1237 10916
rect 1119 10848 1161 10882
rect 1195 10848 1237 10882
rect 1119 10814 1237 10848
rect 1119 10780 1161 10814
rect 1195 10780 1237 10814
rect 1119 10746 1237 10780
rect 1119 10712 1161 10746
rect 1195 10712 1237 10746
rect 1119 10678 1237 10712
rect 1119 10644 1161 10678
rect 1195 10644 1237 10678
rect 1119 10610 1237 10644
rect 1119 10576 1161 10610
rect 1195 10576 1237 10610
rect 1119 10542 1237 10576
rect 1119 10508 1161 10542
rect 1195 10508 1237 10542
rect 1119 10474 1237 10508
rect 1119 10440 1161 10474
rect 1195 10440 1237 10474
rect 1119 10406 1237 10440
rect 1119 10372 1161 10406
rect 1195 10372 1237 10406
rect 1119 10319 1237 10372
rect 13769 26993 13887 27027
rect 13769 26959 13809 26993
rect 13843 26959 13887 26993
rect 13769 26925 13887 26959
rect 13769 26891 13809 26925
rect 13843 26891 13887 26925
rect 13769 26857 13887 26891
rect 13769 26823 13809 26857
rect 13843 26823 13887 26857
rect 13769 26789 13887 26823
rect 13769 26755 13809 26789
rect 13843 26755 13887 26789
rect 13769 26721 13887 26755
rect 13769 26687 13809 26721
rect 13843 26687 13887 26721
rect 13769 26653 13887 26687
rect 13769 26619 13809 26653
rect 13843 26619 13887 26653
rect 13769 26585 13887 26619
rect 13769 26551 13809 26585
rect 13843 26551 13887 26585
rect 13769 26517 13887 26551
rect 13769 26483 13809 26517
rect 13843 26483 13887 26517
rect 13769 26449 13887 26483
rect 13769 26415 13809 26449
rect 13843 26415 13887 26449
rect 13769 26381 13887 26415
rect 13769 26347 13809 26381
rect 13843 26347 13887 26381
rect 13769 26313 13887 26347
rect 13769 26279 13809 26313
rect 13843 26279 13887 26313
rect 13769 26245 13887 26279
rect 13769 26211 13809 26245
rect 13843 26211 13887 26245
rect 13769 26177 13887 26211
rect 13769 26143 13809 26177
rect 13843 26143 13887 26177
rect 13769 26109 13887 26143
rect 13769 26075 13809 26109
rect 13843 26075 13887 26109
rect 13769 26041 13887 26075
rect 13769 26007 13809 26041
rect 13843 26007 13887 26041
rect 13769 25973 13887 26007
rect 13769 25939 13809 25973
rect 13843 25939 13887 25973
rect 13769 25905 13887 25939
rect 13769 25871 13809 25905
rect 13843 25871 13887 25905
rect 13769 25837 13887 25871
rect 13769 25803 13809 25837
rect 13843 25803 13887 25837
rect 13769 25769 13887 25803
rect 13769 25735 13809 25769
rect 13843 25735 13887 25769
rect 13769 25701 13887 25735
rect 13769 25667 13809 25701
rect 13843 25667 13887 25701
rect 13769 25633 13887 25667
rect 13769 25599 13809 25633
rect 13843 25599 13887 25633
rect 13769 25565 13887 25599
rect 13769 25531 13809 25565
rect 13843 25531 13887 25565
rect 13769 25497 13887 25531
rect 13769 25463 13809 25497
rect 13843 25463 13887 25497
rect 13769 25429 13887 25463
rect 13769 25395 13809 25429
rect 13843 25395 13887 25429
rect 13769 25361 13887 25395
rect 13769 25327 13809 25361
rect 13843 25327 13887 25361
rect 13769 25293 13887 25327
rect 13769 25259 13809 25293
rect 13843 25259 13887 25293
rect 13769 25225 13887 25259
rect 13769 25191 13809 25225
rect 13843 25191 13887 25225
rect 13769 25157 13887 25191
rect 13769 25123 13809 25157
rect 13843 25123 13887 25157
rect 13769 25089 13887 25123
rect 13769 25055 13809 25089
rect 13843 25055 13887 25089
rect 13769 25021 13887 25055
rect 13769 24987 13809 25021
rect 13843 24987 13887 25021
rect 13769 24953 13887 24987
rect 13769 24919 13809 24953
rect 13843 24919 13887 24953
rect 13769 24885 13887 24919
rect 13769 24851 13809 24885
rect 13843 24851 13887 24885
rect 13769 24817 13887 24851
rect 13769 24783 13809 24817
rect 13843 24783 13887 24817
rect 13769 24749 13887 24783
rect 13769 24715 13809 24749
rect 13843 24715 13887 24749
rect 13769 24681 13887 24715
rect 13769 24647 13809 24681
rect 13843 24647 13887 24681
rect 13769 24613 13887 24647
rect 13769 24579 13809 24613
rect 13843 24579 13887 24613
rect 13769 24545 13887 24579
rect 13769 24511 13809 24545
rect 13843 24511 13887 24545
rect 13769 24477 13887 24511
rect 13769 24443 13809 24477
rect 13843 24443 13887 24477
rect 13769 24409 13887 24443
rect 13769 24375 13809 24409
rect 13843 24375 13887 24409
rect 13769 24341 13887 24375
rect 13769 24307 13809 24341
rect 13843 24307 13887 24341
rect 13769 24273 13887 24307
rect 13769 24239 13809 24273
rect 13843 24239 13887 24273
rect 13769 24205 13887 24239
rect 13769 24171 13809 24205
rect 13843 24171 13887 24205
rect 13769 24137 13887 24171
rect 13769 24103 13809 24137
rect 13843 24103 13887 24137
rect 13769 24069 13887 24103
rect 13769 24035 13809 24069
rect 13843 24035 13887 24069
rect 13769 24001 13887 24035
rect 13769 23967 13809 24001
rect 13843 23967 13887 24001
rect 13769 23933 13887 23967
rect 13769 23899 13809 23933
rect 13843 23899 13887 23933
rect 13769 23865 13887 23899
rect 13769 23831 13809 23865
rect 13843 23831 13887 23865
rect 13769 23797 13887 23831
rect 13769 23763 13809 23797
rect 13843 23763 13887 23797
rect 13769 23729 13887 23763
rect 13769 23695 13809 23729
rect 13843 23695 13887 23729
rect 13769 23661 13887 23695
rect 13769 23627 13809 23661
rect 13843 23627 13887 23661
rect 13769 23593 13887 23627
rect 13769 23559 13809 23593
rect 13843 23559 13887 23593
rect 13769 23525 13887 23559
rect 13769 23491 13809 23525
rect 13843 23491 13887 23525
rect 13769 23457 13887 23491
rect 13769 23423 13809 23457
rect 13843 23423 13887 23457
rect 13769 23389 13887 23423
rect 13769 23355 13809 23389
rect 13843 23355 13887 23389
rect 13769 23321 13887 23355
rect 13769 23287 13809 23321
rect 13843 23287 13887 23321
rect 13769 23253 13887 23287
rect 13769 23219 13809 23253
rect 13843 23219 13887 23253
rect 13769 23185 13887 23219
rect 13769 23151 13809 23185
rect 13843 23151 13887 23185
rect 13769 23117 13887 23151
rect 13769 23083 13809 23117
rect 13843 23083 13887 23117
rect 13769 23049 13887 23083
rect 13769 23015 13809 23049
rect 13843 23015 13887 23049
rect 13769 22981 13887 23015
rect 13769 22947 13809 22981
rect 13843 22947 13887 22981
rect 13769 22913 13887 22947
rect 13769 22879 13809 22913
rect 13843 22879 13887 22913
rect 13769 22845 13887 22879
rect 13769 22811 13809 22845
rect 13843 22811 13887 22845
rect 13769 22777 13887 22811
rect 13769 22743 13809 22777
rect 13843 22743 13887 22777
rect 13769 22709 13887 22743
rect 13769 22675 13809 22709
rect 13843 22675 13887 22709
rect 13769 22641 13887 22675
rect 13769 22607 13809 22641
rect 13843 22607 13887 22641
rect 13769 22573 13887 22607
rect 13769 22539 13809 22573
rect 13843 22539 13887 22573
rect 13769 22505 13887 22539
rect 13769 22471 13809 22505
rect 13843 22471 13887 22505
rect 13769 22437 13887 22471
rect 13769 22403 13809 22437
rect 13843 22403 13887 22437
rect 13769 22369 13887 22403
rect 13769 22335 13809 22369
rect 13843 22335 13887 22369
rect 13769 22301 13887 22335
rect 13769 22267 13809 22301
rect 13843 22267 13887 22301
rect 13769 22233 13887 22267
rect 13769 22199 13809 22233
rect 13843 22199 13887 22233
rect 13769 22165 13887 22199
rect 13769 22131 13809 22165
rect 13843 22131 13887 22165
rect 13769 22097 13887 22131
rect 13769 22063 13809 22097
rect 13843 22063 13887 22097
rect 13769 22029 13887 22063
rect 13769 21995 13809 22029
rect 13843 21995 13887 22029
rect 13769 21961 13887 21995
rect 13769 21927 13809 21961
rect 13843 21927 13887 21961
rect 13769 21893 13887 21927
rect 13769 21859 13809 21893
rect 13843 21859 13887 21893
rect 13769 21825 13887 21859
rect 13769 21791 13809 21825
rect 13843 21791 13887 21825
rect 13769 21757 13887 21791
rect 13769 21723 13809 21757
rect 13843 21723 13887 21757
rect 13769 21689 13887 21723
rect 13769 21655 13809 21689
rect 13843 21655 13887 21689
rect 13769 21621 13887 21655
rect 13769 21587 13809 21621
rect 13843 21587 13887 21621
rect 13769 21553 13887 21587
rect 13769 21519 13809 21553
rect 13843 21519 13887 21553
rect 13769 21485 13887 21519
rect 13769 21451 13809 21485
rect 13843 21451 13887 21485
rect 13769 21417 13887 21451
rect 13769 21383 13809 21417
rect 13843 21383 13887 21417
rect 13769 21349 13887 21383
rect 13769 21315 13809 21349
rect 13843 21315 13887 21349
rect 13769 21281 13887 21315
rect 13769 21247 13809 21281
rect 13843 21247 13887 21281
rect 13769 21213 13887 21247
rect 13769 21179 13809 21213
rect 13843 21179 13887 21213
rect 13769 21145 13887 21179
rect 13769 21111 13809 21145
rect 13843 21111 13887 21145
rect 13769 21077 13887 21111
rect 13769 21043 13809 21077
rect 13843 21043 13887 21077
rect 13769 21009 13887 21043
rect 13769 20975 13809 21009
rect 13843 20975 13887 21009
rect 13769 20941 13887 20975
rect 13769 20907 13809 20941
rect 13843 20907 13887 20941
rect 13769 20873 13887 20907
rect 13769 20839 13809 20873
rect 13843 20839 13887 20873
rect 13769 20805 13887 20839
rect 13769 20771 13809 20805
rect 13843 20771 13887 20805
rect 13769 20737 13887 20771
rect 13769 20703 13809 20737
rect 13843 20703 13887 20737
rect 13769 20669 13887 20703
rect 13769 20635 13809 20669
rect 13843 20635 13887 20669
rect 13769 20601 13887 20635
rect 13769 20567 13809 20601
rect 13843 20567 13887 20601
rect 13769 20533 13887 20567
rect 13769 20499 13809 20533
rect 13843 20499 13887 20533
rect 13769 20465 13887 20499
rect 13769 20431 13809 20465
rect 13843 20431 13887 20465
rect 13769 20397 13887 20431
rect 13769 20363 13809 20397
rect 13843 20363 13887 20397
rect 13769 20329 13887 20363
rect 13769 20295 13809 20329
rect 13843 20295 13887 20329
rect 13769 20261 13887 20295
rect 13769 20227 13809 20261
rect 13843 20227 13887 20261
rect 13769 20193 13887 20227
rect 13769 20159 13809 20193
rect 13843 20159 13887 20193
rect 13769 20125 13887 20159
rect 13769 20091 13809 20125
rect 13843 20091 13887 20125
rect 13769 20057 13887 20091
rect 13769 20023 13809 20057
rect 13843 20023 13887 20057
rect 13769 19989 13887 20023
rect 13769 19955 13809 19989
rect 13843 19955 13887 19989
rect 13769 19921 13887 19955
rect 13769 19887 13809 19921
rect 13843 19887 13887 19921
rect 13769 19853 13887 19887
rect 13769 19819 13809 19853
rect 13843 19819 13887 19853
rect 13769 19785 13887 19819
rect 13769 19751 13809 19785
rect 13843 19751 13887 19785
rect 13769 19717 13887 19751
rect 13769 19683 13809 19717
rect 13843 19683 13887 19717
rect 13769 19649 13887 19683
rect 13769 19615 13809 19649
rect 13843 19615 13887 19649
rect 13769 19581 13887 19615
rect 13769 19547 13809 19581
rect 13843 19547 13887 19581
rect 13769 19513 13887 19547
rect 13769 19479 13809 19513
rect 13843 19479 13887 19513
rect 13769 19445 13887 19479
rect 13769 19411 13809 19445
rect 13843 19411 13887 19445
rect 13769 19377 13887 19411
rect 13769 19343 13809 19377
rect 13843 19343 13887 19377
rect 13769 19309 13887 19343
rect 13769 19275 13809 19309
rect 13843 19275 13887 19309
rect 13769 19241 13887 19275
rect 13769 19207 13809 19241
rect 13843 19207 13887 19241
rect 13769 19173 13887 19207
rect 13769 19139 13809 19173
rect 13843 19139 13887 19173
rect 13769 19105 13887 19139
rect 13769 19071 13809 19105
rect 13843 19071 13887 19105
rect 13769 19037 13887 19071
rect 13769 19003 13809 19037
rect 13843 19003 13887 19037
rect 13769 18969 13887 19003
rect 13769 18935 13809 18969
rect 13843 18935 13887 18969
rect 13769 18901 13887 18935
rect 13769 18867 13809 18901
rect 13843 18867 13887 18901
rect 13769 18833 13887 18867
rect 13769 18799 13809 18833
rect 13843 18799 13887 18833
rect 13769 18765 13887 18799
rect 13769 18731 13809 18765
rect 13843 18731 13887 18765
rect 13769 18697 13887 18731
rect 13769 18663 13809 18697
rect 13843 18663 13887 18697
rect 13769 18629 13887 18663
rect 13769 18595 13809 18629
rect 13843 18595 13887 18629
rect 13769 18561 13887 18595
rect 13769 18527 13809 18561
rect 13843 18527 13887 18561
rect 13769 18493 13887 18527
rect 13769 18459 13809 18493
rect 13843 18459 13887 18493
rect 13769 18425 13887 18459
rect 13769 18391 13809 18425
rect 13843 18391 13887 18425
rect 13769 18357 13887 18391
rect 13769 18323 13809 18357
rect 13843 18323 13887 18357
rect 13769 18289 13887 18323
rect 13769 18255 13809 18289
rect 13843 18255 13887 18289
rect 13769 18221 13887 18255
rect 13769 18187 13809 18221
rect 13843 18187 13887 18221
rect 13769 18153 13887 18187
rect 13769 18119 13809 18153
rect 13843 18119 13887 18153
rect 13769 18085 13887 18119
rect 13769 18051 13809 18085
rect 13843 18051 13887 18085
rect 13769 18017 13887 18051
rect 13769 17983 13809 18017
rect 13843 17983 13887 18017
rect 13769 17949 13887 17983
rect 13769 17915 13809 17949
rect 13843 17915 13887 17949
rect 13769 17881 13887 17915
rect 13769 17847 13809 17881
rect 13843 17847 13887 17881
rect 13769 17813 13887 17847
rect 13769 17779 13809 17813
rect 13843 17779 13887 17813
rect 13769 17745 13887 17779
rect 13769 17711 13809 17745
rect 13843 17711 13887 17745
rect 13769 17677 13887 17711
rect 13769 17643 13809 17677
rect 13843 17643 13887 17677
rect 13769 17609 13887 17643
rect 13769 17575 13809 17609
rect 13843 17575 13887 17609
rect 13769 17541 13887 17575
rect 13769 17507 13809 17541
rect 13843 17507 13887 17541
rect 13769 17473 13887 17507
rect 13769 17439 13809 17473
rect 13843 17439 13887 17473
rect 13769 17405 13887 17439
rect 13769 17371 13809 17405
rect 13843 17371 13887 17405
rect 13769 17337 13887 17371
rect 13769 17303 13809 17337
rect 13843 17303 13887 17337
rect 13769 17269 13887 17303
rect 13769 17235 13809 17269
rect 13843 17235 13887 17269
rect 13769 17201 13887 17235
rect 13769 17167 13809 17201
rect 13843 17167 13887 17201
rect 13769 17133 13887 17167
rect 13769 17099 13809 17133
rect 13843 17099 13887 17133
rect 13769 17065 13887 17099
rect 13769 17031 13809 17065
rect 13843 17031 13887 17065
rect 13769 16997 13887 17031
rect 13769 16963 13809 16997
rect 13843 16963 13887 16997
rect 13769 16929 13887 16963
rect 13769 16895 13809 16929
rect 13843 16895 13887 16929
rect 13769 16861 13887 16895
rect 13769 16827 13809 16861
rect 13843 16827 13887 16861
rect 13769 16793 13887 16827
rect 13769 16759 13809 16793
rect 13843 16759 13887 16793
rect 13769 16725 13887 16759
rect 13769 16691 13809 16725
rect 13843 16691 13887 16725
rect 13769 16657 13887 16691
rect 13769 16623 13809 16657
rect 13843 16623 13887 16657
rect 13769 16589 13887 16623
rect 13769 16555 13809 16589
rect 13843 16555 13887 16589
rect 13769 16521 13887 16555
rect 13769 16487 13809 16521
rect 13843 16487 13887 16521
rect 13769 16453 13887 16487
rect 13769 16419 13809 16453
rect 13843 16419 13887 16453
rect 13769 16385 13887 16419
rect 13769 16351 13809 16385
rect 13843 16351 13887 16385
rect 13769 16317 13887 16351
rect 13769 16283 13809 16317
rect 13843 16283 13887 16317
rect 13769 16249 13887 16283
rect 13769 16215 13809 16249
rect 13843 16215 13887 16249
rect 13769 16181 13887 16215
rect 13769 16147 13809 16181
rect 13843 16147 13887 16181
rect 13769 16113 13887 16147
rect 13769 16079 13809 16113
rect 13843 16079 13887 16113
rect 13769 16045 13887 16079
rect 13769 16011 13809 16045
rect 13843 16011 13887 16045
rect 13769 15977 13887 16011
rect 13769 15943 13809 15977
rect 13843 15943 13887 15977
rect 13769 15909 13887 15943
rect 13769 15875 13809 15909
rect 13843 15875 13887 15909
rect 13769 15841 13887 15875
rect 13769 15807 13809 15841
rect 13843 15807 13887 15841
rect 13769 15773 13887 15807
rect 13769 15739 13809 15773
rect 13843 15739 13887 15773
rect 13769 15705 13887 15739
rect 13769 15671 13809 15705
rect 13843 15671 13887 15705
rect 13769 15637 13887 15671
rect 13769 15603 13809 15637
rect 13843 15603 13887 15637
rect 13769 15569 13887 15603
rect 13769 15535 13809 15569
rect 13843 15535 13887 15569
rect 13769 15501 13887 15535
rect 13769 15467 13809 15501
rect 13843 15467 13887 15501
rect 13769 15433 13887 15467
rect 13769 15399 13809 15433
rect 13843 15399 13887 15433
rect 13769 15365 13887 15399
rect 13769 15331 13809 15365
rect 13843 15331 13887 15365
rect 13769 15297 13887 15331
rect 13769 15263 13809 15297
rect 13843 15263 13887 15297
rect 13769 15229 13887 15263
rect 13769 15195 13809 15229
rect 13843 15195 13887 15229
rect 13769 15161 13887 15195
rect 13769 15127 13809 15161
rect 13843 15127 13887 15161
rect 13769 15093 13887 15127
rect 13769 15059 13809 15093
rect 13843 15059 13887 15093
rect 13769 15025 13887 15059
rect 13769 14991 13809 15025
rect 13843 14991 13887 15025
rect 13769 14957 13887 14991
rect 13769 14923 13809 14957
rect 13843 14923 13887 14957
rect 13769 14889 13887 14923
rect 13769 14855 13809 14889
rect 13843 14855 13887 14889
rect 13769 14821 13887 14855
rect 13769 14787 13809 14821
rect 13843 14787 13887 14821
rect 13769 14753 13887 14787
rect 13769 14719 13809 14753
rect 13843 14719 13887 14753
rect 13769 14685 13887 14719
rect 13769 14651 13809 14685
rect 13843 14651 13887 14685
rect 13769 14617 13887 14651
rect 13769 14583 13809 14617
rect 13843 14583 13887 14617
rect 13769 14549 13887 14583
rect 13769 14515 13809 14549
rect 13843 14515 13887 14549
rect 13769 14481 13887 14515
rect 13769 14447 13809 14481
rect 13843 14447 13887 14481
rect 13769 14413 13887 14447
rect 13769 14379 13809 14413
rect 13843 14379 13887 14413
rect 13769 14345 13887 14379
rect 13769 14311 13809 14345
rect 13843 14311 13887 14345
rect 13769 14277 13887 14311
rect 13769 14243 13809 14277
rect 13843 14243 13887 14277
rect 13769 14209 13887 14243
rect 13769 14175 13809 14209
rect 13843 14175 13887 14209
rect 13769 14141 13887 14175
rect 13769 14107 13809 14141
rect 13843 14107 13887 14141
rect 13769 14073 13887 14107
rect 13769 14039 13809 14073
rect 13843 14039 13887 14073
rect 13769 14005 13887 14039
rect 13769 13971 13809 14005
rect 13843 13971 13887 14005
rect 13769 13937 13887 13971
rect 13769 13903 13809 13937
rect 13843 13903 13887 13937
rect 13769 13869 13887 13903
rect 13769 13835 13809 13869
rect 13843 13835 13887 13869
rect 13769 13801 13887 13835
rect 13769 13767 13809 13801
rect 13843 13767 13887 13801
rect 13769 13733 13887 13767
rect 13769 13699 13809 13733
rect 13843 13699 13887 13733
rect 13769 13665 13887 13699
rect 13769 13631 13809 13665
rect 13843 13631 13887 13665
rect 13769 13597 13887 13631
rect 13769 13563 13809 13597
rect 13843 13563 13887 13597
rect 13769 13529 13887 13563
rect 13769 13495 13809 13529
rect 13843 13495 13887 13529
rect 13769 13461 13887 13495
rect 13769 13427 13809 13461
rect 13843 13427 13887 13461
rect 13769 13393 13887 13427
rect 13769 13359 13809 13393
rect 13843 13359 13887 13393
rect 13769 13325 13887 13359
rect 13769 13291 13809 13325
rect 13843 13291 13887 13325
rect 13769 13257 13887 13291
rect 13769 13223 13809 13257
rect 13843 13223 13887 13257
rect 13769 13189 13887 13223
rect 13769 13155 13809 13189
rect 13843 13155 13887 13189
rect 13769 13121 13887 13155
rect 13769 13087 13809 13121
rect 13843 13087 13887 13121
rect 13769 13053 13887 13087
rect 13769 13019 13809 13053
rect 13843 13019 13887 13053
rect 13769 12985 13887 13019
rect 13769 12951 13809 12985
rect 13843 12951 13887 12985
rect 13769 12917 13887 12951
rect 13769 12883 13809 12917
rect 13843 12883 13887 12917
rect 13769 12849 13887 12883
rect 13769 12815 13809 12849
rect 13843 12815 13887 12849
rect 13769 12781 13887 12815
rect 13769 12747 13809 12781
rect 13843 12747 13887 12781
rect 13769 12713 13887 12747
rect 13769 12679 13809 12713
rect 13843 12679 13887 12713
rect 13769 12645 13887 12679
rect 13769 12611 13809 12645
rect 13843 12611 13887 12645
rect 13769 12577 13887 12611
rect 13769 12543 13809 12577
rect 13843 12543 13887 12577
rect 13769 12509 13887 12543
rect 13769 12475 13809 12509
rect 13843 12475 13887 12509
rect 13769 12441 13887 12475
rect 13769 12407 13809 12441
rect 13843 12407 13887 12441
rect 13769 12373 13887 12407
rect 13769 12339 13809 12373
rect 13843 12339 13887 12373
rect 13769 12305 13887 12339
rect 13769 12271 13809 12305
rect 13843 12271 13887 12305
rect 13769 12237 13887 12271
rect 13769 12203 13809 12237
rect 13843 12203 13887 12237
rect 13769 12169 13887 12203
rect 13769 12135 13809 12169
rect 13843 12135 13887 12169
rect 13769 12101 13887 12135
rect 13769 12067 13809 12101
rect 13843 12067 13887 12101
rect 13769 12033 13887 12067
rect 13769 11999 13809 12033
rect 13843 11999 13887 12033
rect 13769 11965 13887 11999
rect 13769 11931 13809 11965
rect 13843 11931 13887 11965
rect 13769 11897 13887 11931
rect 13769 11863 13809 11897
rect 13843 11863 13887 11897
rect 13769 11829 13887 11863
rect 13769 11795 13809 11829
rect 13843 11795 13887 11829
rect 13769 11761 13887 11795
rect 13769 11727 13809 11761
rect 13843 11727 13887 11761
rect 13769 11693 13887 11727
rect 13769 11659 13809 11693
rect 13843 11659 13887 11693
rect 13769 11625 13887 11659
rect 13769 11591 13809 11625
rect 13843 11591 13887 11625
rect 13769 11557 13887 11591
rect 13769 11523 13809 11557
rect 13843 11523 13887 11557
rect 13769 11489 13887 11523
rect 13769 11455 13809 11489
rect 13843 11455 13887 11489
rect 13769 11421 13887 11455
rect 13769 11387 13809 11421
rect 13843 11387 13887 11421
rect 13769 11353 13887 11387
rect 13769 11319 13809 11353
rect 13843 11319 13887 11353
rect 13769 11285 13887 11319
rect 13769 11251 13809 11285
rect 13843 11251 13887 11285
rect 13769 11217 13887 11251
rect 13769 11183 13809 11217
rect 13843 11183 13887 11217
rect 13769 11149 13887 11183
rect 13769 11115 13809 11149
rect 13843 11115 13887 11149
rect 13769 11081 13887 11115
rect 13769 11047 13809 11081
rect 13843 11047 13887 11081
rect 13769 11013 13887 11047
rect 13769 10979 13809 11013
rect 13843 10979 13887 11013
rect 13769 10945 13887 10979
rect 13769 10911 13809 10945
rect 13843 10911 13887 10945
rect 13769 10877 13887 10911
rect 13769 10843 13809 10877
rect 13843 10843 13887 10877
rect 13769 10809 13887 10843
rect 13769 10775 13809 10809
rect 13843 10775 13887 10809
rect 13769 10741 13887 10775
rect 13769 10707 13809 10741
rect 13843 10707 13887 10741
rect 13769 10673 13887 10707
rect 13769 10639 13809 10673
rect 13843 10639 13887 10673
rect 13769 10605 13887 10639
rect 13769 10571 13809 10605
rect 13843 10571 13887 10605
rect 13769 10537 13887 10571
rect 13769 10503 13809 10537
rect 13843 10503 13887 10537
rect 13769 10469 13887 10503
rect 13769 10435 13809 10469
rect 13843 10435 13887 10469
rect 13769 10401 13887 10435
rect 13769 10367 13809 10401
rect 13843 10367 13887 10401
rect 13769 10319 13887 10367
rect 1119 10278 13887 10319
rect 1119 10244 1302 10278
rect 1336 10244 1370 10278
rect 1404 10244 1438 10278
rect 1472 10244 1506 10278
rect 1540 10244 1574 10278
rect 1608 10244 1642 10278
rect 1676 10244 1710 10278
rect 1744 10244 1778 10278
rect 1812 10244 1846 10278
rect 1880 10244 1914 10278
rect 1948 10244 1982 10278
rect 2016 10244 2050 10278
rect 2084 10244 2118 10278
rect 2152 10244 2186 10278
rect 2220 10244 2254 10278
rect 2288 10244 2322 10278
rect 2356 10244 2390 10278
rect 2424 10244 2458 10278
rect 2492 10244 2526 10278
rect 2560 10244 2594 10278
rect 2628 10244 2662 10278
rect 2696 10244 2730 10278
rect 2764 10244 2798 10278
rect 2832 10244 2866 10278
rect 2900 10244 2934 10278
rect 2968 10244 3002 10278
rect 3036 10244 3070 10278
rect 3104 10244 3138 10278
rect 3172 10244 3206 10278
rect 3240 10244 3274 10278
rect 3308 10244 3342 10278
rect 3376 10244 3410 10278
rect 3444 10244 3478 10278
rect 3512 10244 3546 10278
rect 3580 10244 3614 10278
rect 3648 10244 3682 10278
rect 3716 10244 3750 10278
rect 3784 10244 3818 10278
rect 3852 10244 3886 10278
rect 3920 10244 3954 10278
rect 3988 10244 4022 10278
rect 4056 10244 4090 10278
rect 4124 10244 4158 10278
rect 4192 10244 4226 10278
rect 4260 10244 4294 10278
rect 4328 10244 4362 10278
rect 4396 10244 4430 10278
rect 4464 10244 4498 10278
rect 4532 10244 4566 10278
rect 4600 10244 4634 10278
rect 4668 10244 4702 10278
rect 4736 10244 4770 10278
rect 4804 10244 4838 10278
rect 4872 10244 4906 10278
rect 4940 10244 4974 10278
rect 5008 10244 5042 10278
rect 5076 10244 5110 10278
rect 5144 10244 5178 10278
rect 5212 10244 5246 10278
rect 5280 10244 5314 10278
rect 5348 10244 5382 10278
rect 5416 10244 5450 10278
rect 5484 10244 5518 10278
rect 5552 10244 5586 10278
rect 5620 10244 5654 10278
rect 5688 10244 5722 10278
rect 5756 10244 5790 10278
rect 5824 10244 5858 10278
rect 5892 10244 5926 10278
rect 5960 10244 5994 10278
rect 6028 10244 6062 10278
rect 6096 10244 6130 10278
rect 6164 10244 6198 10278
rect 6232 10244 6266 10278
rect 6300 10244 6334 10278
rect 6368 10244 6402 10278
rect 6436 10244 6470 10278
rect 6504 10244 6538 10278
rect 6572 10244 6606 10278
rect 6640 10244 6674 10278
rect 6708 10244 6742 10278
rect 6776 10244 6810 10278
rect 6844 10244 6878 10278
rect 6912 10244 6946 10278
rect 6980 10244 7014 10278
rect 7048 10244 7082 10278
rect 7116 10244 7150 10278
rect 7184 10244 7218 10278
rect 7252 10244 7286 10278
rect 7320 10244 7354 10278
rect 7388 10244 7422 10278
rect 7456 10244 7490 10278
rect 7524 10244 7558 10278
rect 7592 10244 7626 10278
rect 7660 10244 7694 10278
rect 7728 10244 7762 10278
rect 7796 10244 7830 10278
rect 7864 10244 7898 10278
rect 7932 10244 7966 10278
rect 8000 10244 8034 10278
rect 8068 10244 8102 10278
rect 8136 10244 8170 10278
rect 8204 10244 8238 10278
rect 8272 10244 8306 10278
rect 8340 10244 8374 10278
rect 8408 10244 8442 10278
rect 8476 10244 8510 10278
rect 8544 10244 8578 10278
rect 8612 10244 8646 10278
rect 8680 10244 8714 10278
rect 8748 10244 8782 10278
rect 8816 10244 8850 10278
rect 8884 10244 8918 10278
rect 8952 10244 8986 10278
rect 9020 10244 9054 10278
rect 9088 10244 9122 10278
rect 9156 10244 9190 10278
rect 9224 10244 9258 10278
rect 9292 10244 9326 10278
rect 9360 10244 9394 10278
rect 9428 10244 9462 10278
rect 9496 10244 9530 10278
rect 9564 10244 9598 10278
rect 9632 10244 9666 10278
rect 9700 10244 9734 10278
rect 9768 10244 9802 10278
rect 9836 10244 9870 10278
rect 9904 10244 9938 10278
rect 9972 10244 10006 10278
rect 10040 10244 10074 10278
rect 10108 10244 10142 10278
rect 10176 10244 10210 10278
rect 10244 10244 10278 10278
rect 10312 10244 10346 10278
rect 10380 10244 10414 10278
rect 10448 10244 10482 10278
rect 10516 10244 10550 10278
rect 10584 10244 10618 10278
rect 10652 10244 10686 10278
rect 10720 10244 10754 10278
rect 10788 10244 10822 10278
rect 10856 10244 10890 10278
rect 10924 10244 10958 10278
rect 10992 10244 11026 10278
rect 11060 10244 11094 10278
rect 11128 10244 11162 10278
rect 11196 10244 11230 10278
rect 11264 10244 11298 10278
rect 11332 10244 11366 10278
rect 11400 10244 11434 10278
rect 11468 10244 11502 10278
rect 11536 10244 11570 10278
rect 11604 10244 11638 10278
rect 11672 10244 11706 10278
rect 11740 10244 11774 10278
rect 11808 10244 11842 10278
rect 11876 10244 11910 10278
rect 11944 10244 11978 10278
rect 12012 10244 12046 10278
rect 12080 10244 12114 10278
rect 12148 10244 12182 10278
rect 12216 10244 12250 10278
rect 12284 10244 12318 10278
rect 12352 10244 12386 10278
rect 12420 10244 12454 10278
rect 12488 10244 12522 10278
rect 12556 10244 12590 10278
rect 12624 10244 12658 10278
rect 12692 10244 12726 10278
rect 12760 10244 12794 10278
rect 12828 10244 12862 10278
rect 12896 10244 12930 10278
rect 12964 10244 12998 10278
rect 13032 10244 13066 10278
rect 13100 10244 13134 10278
rect 13168 10244 13202 10278
rect 13236 10244 13270 10278
rect 13304 10244 13338 10278
rect 13372 10244 13406 10278
rect 13440 10244 13474 10278
rect 13508 10244 13542 10278
rect 13576 10244 13610 10278
rect 13644 10244 13678 10278
rect 13712 10244 13887 10278
rect 1119 10201 13887 10244
rect 14539 36208 14724 36242
rect 14539 36174 14607 36208
rect 14641 36174 14724 36208
rect 14539 36140 14724 36174
rect 14539 36106 14607 36140
rect 14641 36106 14724 36140
rect 14539 36072 14724 36106
rect 14539 36038 14607 36072
rect 14641 36038 14724 36072
rect 14539 36004 14724 36038
rect 14539 35970 14607 36004
rect 14641 35970 14724 36004
rect 14539 35936 14724 35970
rect 14539 35902 14607 35936
rect 14641 35902 14724 35936
rect 14539 35868 14724 35902
rect 14539 35834 14607 35868
rect 14641 35834 14724 35868
rect 14539 35800 14724 35834
rect 14539 35766 14607 35800
rect 14641 35766 14724 35800
rect 14539 35732 14724 35766
rect 14539 35698 14607 35732
rect 14641 35698 14724 35732
rect 14539 35664 14724 35698
rect 14539 35630 14607 35664
rect 14641 35630 14724 35664
rect 14539 35596 14724 35630
rect 14539 35562 14607 35596
rect 14641 35562 14724 35596
rect 14539 35528 14724 35562
rect 14539 35494 14607 35528
rect 14641 35494 14724 35528
rect 14539 35460 14724 35494
rect 14539 35426 14607 35460
rect 14641 35426 14724 35460
rect 14539 35392 14724 35426
rect 14539 35358 14607 35392
rect 14641 35358 14724 35392
rect 14539 35324 14724 35358
rect 14539 35290 14607 35324
rect 14641 35290 14724 35324
rect 14539 35256 14724 35290
rect 14539 35222 14607 35256
rect 14641 35222 14724 35256
rect 14539 35188 14724 35222
rect 14539 35154 14607 35188
rect 14641 35154 14724 35188
rect 14539 35120 14724 35154
rect 14539 35086 14607 35120
rect 14641 35086 14724 35120
rect 14539 35052 14724 35086
rect 14539 35018 14607 35052
rect 14641 35018 14724 35052
rect 14539 34984 14724 35018
rect 14539 34950 14607 34984
rect 14641 34950 14724 34984
rect 14539 34916 14724 34950
rect 14539 34882 14607 34916
rect 14641 34882 14724 34916
rect 14539 34848 14724 34882
rect 14539 34814 14607 34848
rect 14641 34814 14724 34848
rect 14539 34780 14724 34814
rect 14539 34746 14607 34780
rect 14641 34746 14724 34780
rect 14539 34712 14724 34746
rect 14539 34678 14607 34712
rect 14641 34678 14724 34712
rect 14539 34644 14724 34678
rect 14539 34610 14607 34644
rect 14641 34610 14724 34644
rect 14539 34576 14724 34610
rect 14539 34542 14607 34576
rect 14641 34542 14724 34576
rect 14539 34508 14724 34542
rect 14539 34474 14607 34508
rect 14641 34474 14724 34508
rect 14539 34440 14724 34474
rect 14539 34406 14607 34440
rect 14641 34406 14724 34440
rect 14539 34372 14724 34406
rect 14539 34338 14607 34372
rect 14641 34338 14724 34372
rect 14539 34304 14724 34338
rect 14539 34270 14607 34304
rect 14641 34270 14724 34304
rect 14539 34236 14724 34270
rect 14539 34202 14607 34236
rect 14641 34202 14724 34236
rect 14539 34168 14724 34202
rect 14539 34134 14607 34168
rect 14641 34134 14724 34168
rect 14539 34100 14724 34134
rect 14539 34066 14607 34100
rect 14641 34066 14724 34100
rect 14539 34032 14724 34066
rect 14539 33998 14607 34032
rect 14641 33998 14724 34032
rect 14539 33964 14724 33998
rect 14539 33930 14607 33964
rect 14641 33930 14724 33964
rect 14539 33896 14724 33930
rect 14539 33862 14607 33896
rect 14641 33862 14724 33896
rect 14539 33828 14724 33862
rect 14539 33794 14607 33828
rect 14641 33794 14724 33828
rect 14539 33760 14724 33794
rect 14539 33726 14607 33760
rect 14641 33726 14724 33760
rect 14539 33692 14724 33726
rect 14539 33658 14607 33692
rect 14641 33658 14724 33692
rect 14539 33624 14724 33658
rect 14539 33590 14607 33624
rect 14641 33590 14724 33624
rect 14539 33556 14724 33590
rect 14539 33522 14607 33556
rect 14641 33522 14724 33556
rect 14539 33488 14724 33522
rect 14539 33454 14607 33488
rect 14641 33454 14724 33488
rect 14539 33420 14724 33454
rect 14539 33386 14607 33420
rect 14641 33386 14724 33420
rect 14539 33352 14724 33386
rect 14539 33318 14607 33352
rect 14641 33318 14724 33352
rect 14539 33284 14724 33318
rect 14539 33250 14607 33284
rect 14641 33250 14724 33284
rect 14539 33216 14724 33250
rect 14539 33182 14607 33216
rect 14641 33182 14724 33216
rect 14539 33148 14724 33182
rect 14539 33114 14607 33148
rect 14641 33114 14724 33148
rect 14539 33080 14724 33114
rect 14539 33046 14607 33080
rect 14641 33046 14724 33080
rect 14539 33012 14724 33046
rect 14539 32978 14607 33012
rect 14641 32978 14724 33012
rect 14539 32944 14724 32978
rect 14539 32910 14607 32944
rect 14641 32910 14724 32944
rect 14539 32876 14724 32910
rect 14539 32842 14607 32876
rect 14641 32842 14724 32876
rect 14539 32808 14724 32842
rect 14539 32774 14607 32808
rect 14641 32774 14724 32808
rect 14539 32740 14724 32774
rect 14539 32706 14607 32740
rect 14641 32706 14724 32740
rect 14539 32672 14724 32706
rect 14539 32638 14607 32672
rect 14641 32638 14724 32672
rect 14539 32604 14724 32638
rect 14539 32570 14607 32604
rect 14641 32570 14724 32604
rect 14539 32536 14724 32570
rect 14539 32502 14607 32536
rect 14641 32502 14724 32536
rect 14539 32468 14724 32502
rect 14539 32434 14607 32468
rect 14641 32434 14724 32468
rect 14539 32400 14724 32434
rect 14539 32366 14607 32400
rect 14641 32366 14724 32400
rect 14539 32332 14724 32366
rect 14539 32298 14607 32332
rect 14641 32298 14724 32332
rect 14539 32264 14724 32298
rect 14539 32230 14607 32264
rect 14641 32230 14724 32264
rect 14539 32196 14724 32230
rect 14539 32162 14607 32196
rect 14641 32162 14724 32196
rect 14539 32128 14724 32162
rect 14539 32094 14607 32128
rect 14641 32094 14724 32128
rect 14539 32060 14724 32094
rect 14539 32026 14607 32060
rect 14641 32026 14724 32060
rect 14539 31992 14724 32026
rect 14539 31958 14607 31992
rect 14641 31958 14724 31992
rect 14539 31924 14724 31958
rect 14539 31890 14607 31924
rect 14641 31890 14724 31924
rect 14539 31856 14724 31890
rect 14539 31822 14607 31856
rect 14641 31822 14724 31856
rect 14539 31788 14724 31822
rect 14539 31754 14607 31788
rect 14641 31754 14724 31788
rect 14539 31720 14724 31754
rect 14539 31686 14607 31720
rect 14641 31686 14724 31720
rect 14539 31652 14724 31686
rect 14539 31618 14607 31652
rect 14641 31618 14724 31652
rect 14539 31584 14724 31618
rect 14539 31550 14607 31584
rect 14641 31550 14724 31584
rect 14539 31516 14724 31550
rect 14539 31482 14607 31516
rect 14641 31482 14724 31516
rect 14539 31448 14724 31482
rect 14539 31414 14607 31448
rect 14641 31414 14724 31448
rect 14539 31380 14724 31414
rect 14539 31346 14607 31380
rect 14641 31346 14724 31380
rect 14539 31312 14724 31346
rect 14539 31278 14607 31312
rect 14641 31278 14724 31312
rect 14539 31244 14724 31278
rect 14539 31210 14607 31244
rect 14641 31210 14724 31244
rect 14539 31176 14724 31210
rect 14539 31142 14607 31176
rect 14641 31142 14724 31176
rect 14539 31108 14724 31142
rect 14539 31074 14607 31108
rect 14641 31074 14724 31108
rect 14539 31040 14724 31074
rect 14539 31006 14607 31040
rect 14641 31006 14724 31040
rect 14539 30972 14724 31006
rect 14539 30938 14607 30972
rect 14641 30938 14724 30972
rect 14539 30904 14724 30938
rect 14539 30870 14607 30904
rect 14641 30870 14724 30904
rect 14539 30836 14724 30870
rect 14539 30802 14607 30836
rect 14641 30802 14724 30836
rect 14539 30768 14724 30802
rect 14539 30734 14607 30768
rect 14641 30734 14724 30768
rect 14539 30700 14724 30734
rect 14539 30666 14607 30700
rect 14641 30666 14724 30700
rect 14539 30632 14724 30666
rect 14539 30598 14607 30632
rect 14641 30598 14724 30632
rect 14539 30564 14724 30598
rect 14539 30530 14607 30564
rect 14641 30530 14724 30564
rect 14539 30496 14724 30530
rect 14539 30462 14607 30496
rect 14641 30462 14724 30496
rect 14539 30428 14724 30462
rect 14539 30394 14607 30428
rect 14641 30394 14724 30428
rect 14539 30360 14724 30394
rect 14539 30326 14607 30360
rect 14641 30326 14724 30360
rect 14539 30292 14724 30326
rect 14539 30258 14607 30292
rect 14641 30258 14724 30292
rect 14539 30224 14724 30258
rect 14539 30190 14607 30224
rect 14641 30190 14724 30224
rect 14539 30156 14724 30190
rect 14539 30122 14607 30156
rect 14641 30122 14724 30156
rect 14539 30088 14724 30122
rect 14539 30054 14607 30088
rect 14641 30054 14724 30088
rect 14539 30020 14724 30054
rect 14539 29986 14607 30020
rect 14641 29986 14724 30020
rect 14539 29952 14724 29986
rect 14539 29918 14607 29952
rect 14641 29918 14724 29952
rect 14539 29884 14724 29918
rect 14539 29850 14607 29884
rect 14641 29850 14724 29884
rect 14539 29816 14724 29850
rect 14539 29782 14607 29816
rect 14641 29782 14724 29816
rect 14539 29748 14724 29782
rect 14539 29714 14607 29748
rect 14641 29714 14724 29748
rect 14539 29680 14724 29714
rect 14539 29646 14607 29680
rect 14641 29646 14724 29680
rect 14539 29612 14724 29646
rect 14539 29578 14607 29612
rect 14641 29578 14724 29612
rect 14539 29544 14724 29578
rect 14539 29510 14607 29544
rect 14641 29510 14724 29544
rect 14539 29476 14724 29510
rect 14539 29442 14607 29476
rect 14641 29442 14724 29476
rect 14539 29408 14724 29442
rect 14539 29374 14607 29408
rect 14641 29374 14724 29408
rect 14539 29340 14724 29374
rect 14539 29306 14607 29340
rect 14641 29306 14724 29340
rect 14539 29272 14724 29306
rect 14539 29238 14607 29272
rect 14641 29238 14724 29272
rect 14539 29204 14724 29238
rect 14539 29170 14607 29204
rect 14641 29170 14724 29204
rect 14539 29136 14724 29170
rect 14539 29102 14607 29136
rect 14641 29102 14724 29136
rect 14539 29068 14724 29102
rect 14539 29034 14607 29068
rect 14641 29034 14724 29068
rect 14539 29000 14724 29034
rect 14539 28966 14607 29000
rect 14641 28966 14724 29000
rect 14539 28932 14724 28966
rect 14539 28898 14607 28932
rect 14641 28898 14724 28932
rect 14539 28864 14724 28898
rect 14539 28830 14607 28864
rect 14641 28830 14724 28864
rect 14539 28796 14724 28830
rect 14539 28762 14607 28796
rect 14641 28762 14724 28796
rect 14539 28728 14724 28762
rect 14539 28694 14607 28728
rect 14641 28694 14724 28728
rect 14539 28660 14724 28694
rect 14539 28626 14607 28660
rect 14641 28626 14724 28660
rect 14539 28592 14724 28626
rect 14539 28558 14607 28592
rect 14641 28558 14724 28592
rect 14539 28524 14724 28558
rect 14539 28490 14607 28524
rect 14641 28490 14724 28524
rect 14539 28456 14724 28490
rect 14539 28422 14607 28456
rect 14641 28422 14724 28456
rect 14539 28388 14724 28422
rect 14539 28354 14607 28388
rect 14641 28354 14724 28388
rect 14539 28320 14724 28354
rect 14539 28286 14607 28320
rect 14641 28286 14724 28320
rect 14539 28252 14724 28286
rect 14539 28218 14607 28252
rect 14641 28218 14724 28252
rect 14539 28184 14724 28218
rect 14539 28150 14607 28184
rect 14641 28150 14724 28184
rect 14539 28116 14724 28150
rect 14539 28082 14607 28116
rect 14641 28082 14724 28116
rect 14539 28048 14724 28082
rect 14539 28014 14607 28048
rect 14641 28014 14724 28048
rect 14539 27980 14724 28014
rect 14539 27946 14607 27980
rect 14641 27946 14724 27980
rect 14539 27912 14724 27946
rect 14539 27878 14607 27912
rect 14641 27878 14724 27912
rect 14539 27844 14724 27878
rect 14539 27810 14607 27844
rect 14641 27810 14724 27844
rect 14539 27776 14724 27810
rect 14539 27742 14607 27776
rect 14641 27742 14724 27776
rect 14539 27708 14724 27742
rect 14539 27674 14607 27708
rect 14641 27674 14724 27708
rect 14539 27640 14724 27674
rect 14539 27606 14607 27640
rect 14641 27606 14724 27640
rect 14539 27572 14724 27606
rect 14539 27538 14607 27572
rect 14641 27538 14724 27572
rect 14539 27504 14724 27538
rect 14539 27470 14607 27504
rect 14641 27470 14724 27504
rect 14539 27436 14724 27470
rect 14539 27402 14607 27436
rect 14641 27402 14724 27436
rect 14539 27368 14724 27402
rect 14539 27334 14607 27368
rect 14641 27334 14724 27368
rect 14539 27300 14724 27334
rect 14539 27266 14607 27300
rect 14641 27266 14724 27300
rect 14539 27232 14724 27266
rect 14539 27198 14607 27232
rect 14641 27198 14724 27232
rect 14539 27164 14724 27198
rect 14539 27130 14607 27164
rect 14641 27130 14724 27164
rect 14539 27096 14724 27130
rect 14539 27062 14607 27096
rect 14641 27062 14724 27096
rect 14539 27028 14724 27062
rect 14539 26994 14607 27028
rect 14641 26994 14724 27028
rect 14539 26960 14724 26994
rect 14539 26926 14607 26960
rect 14641 26926 14724 26960
rect 14539 26892 14724 26926
rect 14539 26858 14607 26892
rect 14641 26858 14724 26892
rect 14539 26824 14724 26858
rect 14539 26790 14607 26824
rect 14641 26790 14724 26824
rect 14539 26756 14724 26790
rect 14539 26722 14607 26756
rect 14641 26722 14724 26756
rect 14539 26688 14724 26722
rect 14539 26654 14607 26688
rect 14641 26654 14724 26688
rect 14539 26620 14724 26654
rect 14539 26586 14607 26620
rect 14641 26586 14724 26620
rect 14539 26552 14724 26586
rect 14539 26518 14607 26552
rect 14641 26518 14724 26552
rect 14539 26484 14724 26518
rect 14539 26450 14607 26484
rect 14641 26450 14724 26484
rect 14539 26416 14724 26450
rect 14539 26382 14607 26416
rect 14641 26382 14724 26416
rect 14539 26348 14724 26382
rect 14539 26314 14607 26348
rect 14641 26314 14724 26348
rect 14539 26280 14724 26314
rect 14539 26246 14607 26280
rect 14641 26246 14724 26280
rect 14539 26212 14724 26246
rect 14539 26178 14607 26212
rect 14641 26178 14724 26212
rect 14539 26144 14724 26178
rect 14539 26110 14607 26144
rect 14641 26110 14724 26144
rect 14539 26076 14724 26110
rect 14539 26042 14607 26076
rect 14641 26042 14724 26076
rect 14539 26008 14724 26042
rect 14539 25974 14607 26008
rect 14641 25974 14724 26008
rect 14539 25940 14724 25974
rect 14539 25906 14607 25940
rect 14641 25906 14724 25940
rect 14539 25872 14724 25906
rect 14539 25838 14607 25872
rect 14641 25838 14724 25872
rect 14539 25804 14724 25838
rect 14539 25770 14607 25804
rect 14641 25770 14724 25804
rect 14539 25736 14724 25770
rect 14539 25702 14607 25736
rect 14641 25702 14724 25736
rect 14539 25668 14724 25702
rect 14539 25634 14607 25668
rect 14641 25634 14724 25668
rect 14539 25600 14724 25634
rect 14539 25566 14607 25600
rect 14641 25566 14724 25600
rect 14539 25532 14724 25566
rect 14539 25498 14607 25532
rect 14641 25498 14724 25532
rect 14539 25464 14724 25498
rect 14539 25430 14607 25464
rect 14641 25430 14724 25464
rect 14539 25396 14724 25430
rect 14539 25362 14607 25396
rect 14641 25362 14724 25396
rect 14539 25328 14724 25362
rect 14539 25294 14607 25328
rect 14641 25294 14724 25328
rect 14539 25260 14724 25294
rect 14539 25226 14607 25260
rect 14641 25226 14724 25260
rect 14539 25192 14724 25226
rect 14539 25158 14607 25192
rect 14641 25158 14724 25192
rect 14539 25124 14724 25158
rect 14539 25090 14607 25124
rect 14641 25090 14724 25124
rect 14539 25056 14724 25090
rect 14539 25022 14607 25056
rect 14641 25022 14724 25056
rect 14539 24988 14724 25022
rect 14539 24954 14607 24988
rect 14641 24954 14724 24988
rect 14539 24920 14724 24954
rect 14539 24886 14607 24920
rect 14641 24886 14724 24920
rect 14539 24852 14724 24886
rect 14539 24818 14607 24852
rect 14641 24818 14724 24852
rect 14539 24784 14724 24818
rect 14539 24750 14607 24784
rect 14641 24750 14724 24784
rect 14539 24716 14724 24750
rect 14539 24682 14607 24716
rect 14641 24682 14724 24716
rect 14539 24648 14724 24682
rect 14539 24614 14607 24648
rect 14641 24614 14724 24648
rect 14539 24580 14724 24614
rect 14539 24546 14607 24580
rect 14641 24546 14724 24580
rect 14539 24512 14724 24546
rect 14539 24478 14607 24512
rect 14641 24478 14724 24512
rect 14539 24444 14724 24478
rect 14539 24410 14607 24444
rect 14641 24410 14724 24444
rect 14539 24376 14724 24410
rect 14539 24342 14607 24376
rect 14641 24342 14724 24376
rect 14539 24308 14724 24342
rect 14539 24274 14607 24308
rect 14641 24274 14724 24308
rect 14539 24240 14724 24274
rect 14539 24206 14607 24240
rect 14641 24206 14724 24240
rect 14539 24172 14724 24206
rect 14539 24138 14607 24172
rect 14641 24138 14724 24172
rect 14539 24104 14724 24138
rect 14539 24070 14607 24104
rect 14641 24070 14724 24104
rect 14539 24036 14724 24070
rect 14539 24002 14607 24036
rect 14641 24002 14724 24036
rect 14539 23968 14724 24002
rect 14539 23934 14607 23968
rect 14641 23934 14724 23968
rect 14539 23900 14724 23934
rect 14539 23866 14607 23900
rect 14641 23866 14724 23900
rect 14539 23832 14724 23866
rect 14539 23798 14607 23832
rect 14641 23798 14724 23832
rect 14539 23764 14724 23798
rect 14539 23730 14607 23764
rect 14641 23730 14724 23764
rect 14539 23696 14724 23730
rect 14539 23662 14607 23696
rect 14641 23662 14724 23696
rect 14539 23628 14724 23662
rect 14539 23594 14607 23628
rect 14641 23594 14724 23628
rect 14539 23560 14724 23594
rect 14539 23526 14607 23560
rect 14641 23526 14724 23560
rect 14539 23492 14724 23526
rect 14539 23458 14607 23492
rect 14641 23458 14724 23492
rect 14539 23424 14724 23458
rect 14539 23390 14607 23424
rect 14641 23390 14724 23424
rect 14539 23356 14724 23390
rect 14539 23322 14607 23356
rect 14641 23322 14724 23356
rect 14539 23288 14724 23322
rect 14539 23254 14607 23288
rect 14641 23254 14724 23288
rect 14539 23220 14724 23254
rect 14539 23186 14607 23220
rect 14641 23186 14724 23220
rect 14539 23152 14724 23186
rect 14539 23118 14607 23152
rect 14641 23118 14724 23152
rect 14539 23084 14724 23118
rect 14539 23050 14607 23084
rect 14641 23050 14724 23084
rect 14539 23016 14724 23050
rect 14539 22982 14607 23016
rect 14641 22982 14724 23016
rect 14539 22948 14724 22982
rect 14539 22914 14607 22948
rect 14641 22914 14724 22948
rect 14539 22880 14724 22914
rect 14539 22846 14607 22880
rect 14641 22846 14724 22880
rect 14539 22812 14724 22846
rect 14539 22778 14607 22812
rect 14641 22778 14724 22812
rect 14539 22744 14724 22778
rect 14539 22710 14607 22744
rect 14641 22710 14724 22744
rect 14539 22676 14724 22710
rect 14539 22642 14607 22676
rect 14641 22642 14724 22676
rect 14539 22608 14724 22642
rect 14539 22574 14607 22608
rect 14641 22574 14724 22608
rect 14539 22540 14724 22574
rect 14539 22506 14607 22540
rect 14641 22506 14724 22540
rect 14539 22472 14724 22506
rect 14539 22438 14607 22472
rect 14641 22438 14724 22472
rect 14539 22404 14724 22438
rect 14539 22370 14607 22404
rect 14641 22370 14724 22404
rect 14539 22336 14724 22370
rect 14539 22302 14607 22336
rect 14641 22302 14724 22336
rect 14539 22268 14724 22302
rect 14539 22234 14607 22268
rect 14641 22234 14724 22268
rect 14539 22200 14724 22234
rect 14539 22166 14607 22200
rect 14641 22166 14724 22200
rect 14539 22132 14724 22166
rect 14539 22098 14607 22132
rect 14641 22098 14724 22132
rect 14539 22064 14724 22098
rect 14539 22030 14607 22064
rect 14641 22030 14724 22064
rect 14539 21996 14724 22030
rect 14539 21962 14607 21996
rect 14641 21962 14724 21996
rect 14539 21928 14724 21962
rect 14539 21894 14607 21928
rect 14641 21894 14724 21928
rect 14539 21860 14724 21894
rect 14539 21826 14607 21860
rect 14641 21826 14724 21860
rect 14539 21792 14724 21826
rect 14539 21758 14607 21792
rect 14641 21758 14724 21792
rect 14539 21724 14724 21758
rect 14539 21690 14607 21724
rect 14641 21690 14724 21724
rect 14539 21656 14724 21690
rect 14539 21622 14607 21656
rect 14641 21622 14724 21656
rect 14539 21588 14724 21622
rect 14539 21554 14607 21588
rect 14641 21554 14724 21588
rect 14539 21520 14724 21554
rect 14539 21486 14607 21520
rect 14641 21486 14724 21520
rect 14539 21452 14724 21486
rect 14539 21418 14607 21452
rect 14641 21418 14724 21452
rect 14539 21384 14724 21418
rect 14539 21350 14607 21384
rect 14641 21350 14724 21384
rect 14539 21316 14724 21350
rect 14539 21282 14607 21316
rect 14641 21282 14724 21316
rect 14539 21248 14724 21282
rect 14539 21214 14607 21248
rect 14641 21214 14724 21248
rect 14539 21180 14724 21214
rect 14539 21146 14607 21180
rect 14641 21146 14724 21180
rect 14539 21112 14724 21146
rect 14539 21078 14607 21112
rect 14641 21078 14724 21112
rect 14539 21044 14724 21078
rect 14539 21010 14607 21044
rect 14641 21010 14724 21044
rect 14539 20976 14724 21010
rect 14539 20942 14607 20976
rect 14641 20942 14724 20976
rect 14539 20908 14724 20942
rect 14539 20874 14607 20908
rect 14641 20874 14724 20908
rect 14539 20840 14724 20874
rect 14539 20806 14607 20840
rect 14641 20806 14724 20840
rect 14539 20772 14724 20806
rect 14539 20738 14607 20772
rect 14641 20738 14724 20772
rect 14539 20704 14724 20738
rect 14539 20670 14607 20704
rect 14641 20670 14724 20704
rect 14539 20636 14724 20670
rect 14539 20602 14607 20636
rect 14641 20602 14724 20636
rect 14539 20568 14724 20602
rect 14539 20534 14607 20568
rect 14641 20534 14724 20568
rect 14539 20500 14724 20534
rect 14539 20466 14607 20500
rect 14641 20466 14724 20500
rect 14539 20432 14724 20466
rect 14539 20398 14607 20432
rect 14641 20398 14724 20432
rect 14539 20364 14724 20398
rect 14539 20330 14607 20364
rect 14641 20330 14724 20364
rect 14539 20296 14724 20330
rect 14539 20262 14607 20296
rect 14641 20262 14724 20296
rect 14539 20228 14724 20262
rect 14539 20194 14607 20228
rect 14641 20194 14724 20228
rect 14539 20160 14724 20194
rect 14539 20126 14607 20160
rect 14641 20126 14724 20160
rect 14539 20092 14724 20126
rect 14539 20058 14607 20092
rect 14641 20058 14724 20092
rect 14539 20024 14724 20058
rect 14539 19990 14607 20024
rect 14641 19990 14724 20024
rect 14539 19956 14724 19990
rect 14539 19922 14607 19956
rect 14641 19922 14724 19956
rect 14539 19888 14724 19922
rect 14539 19854 14607 19888
rect 14641 19854 14724 19888
rect 14539 19820 14724 19854
rect 14539 19786 14607 19820
rect 14641 19786 14724 19820
rect 14539 19752 14724 19786
rect 14539 19718 14607 19752
rect 14641 19718 14724 19752
rect 14539 19684 14724 19718
rect 14539 19650 14607 19684
rect 14641 19650 14724 19684
rect 14539 19616 14724 19650
rect 14539 19582 14607 19616
rect 14641 19582 14724 19616
rect 14539 19548 14724 19582
rect 14539 19514 14607 19548
rect 14641 19514 14724 19548
rect 14539 19480 14724 19514
rect 14539 19446 14607 19480
rect 14641 19446 14724 19480
rect 14539 19412 14724 19446
rect 14539 19378 14607 19412
rect 14641 19378 14724 19412
rect 14539 19344 14724 19378
rect 14539 19310 14607 19344
rect 14641 19310 14724 19344
rect 14539 19276 14724 19310
rect 14539 19242 14607 19276
rect 14641 19242 14724 19276
rect 14539 19208 14724 19242
rect 14539 19174 14607 19208
rect 14641 19174 14724 19208
rect 14539 19140 14724 19174
rect 14539 19106 14607 19140
rect 14641 19106 14724 19140
rect 14539 19072 14724 19106
rect 14539 19038 14607 19072
rect 14641 19038 14724 19072
rect 14539 19004 14724 19038
rect 14539 18970 14607 19004
rect 14641 18970 14724 19004
rect 14539 18936 14724 18970
rect 14539 18902 14607 18936
rect 14641 18902 14724 18936
rect 14539 18868 14724 18902
rect 14539 18834 14607 18868
rect 14641 18834 14724 18868
rect 14539 18800 14724 18834
rect 14539 18766 14607 18800
rect 14641 18766 14724 18800
rect 14539 18732 14724 18766
rect 14539 18698 14607 18732
rect 14641 18698 14724 18732
rect 14539 18664 14724 18698
rect 14539 18630 14607 18664
rect 14641 18630 14724 18664
rect 14539 18596 14724 18630
rect 14539 18562 14607 18596
rect 14641 18562 14724 18596
rect 14539 18528 14724 18562
rect 14539 18494 14607 18528
rect 14641 18494 14724 18528
rect 14539 18460 14724 18494
rect 14539 18426 14607 18460
rect 14641 18426 14724 18460
rect 14539 18392 14724 18426
rect 14539 18358 14607 18392
rect 14641 18358 14724 18392
rect 14539 18324 14724 18358
rect 14539 18290 14607 18324
rect 14641 18290 14724 18324
rect 14539 18256 14724 18290
rect 14539 18222 14607 18256
rect 14641 18222 14724 18256
rect 14539 18188 14724 18222
rect 14539 18154 14607 18188
rect 14641 18154 14724 18188
rect 14539 18120 14724 18154
rect 14539 18086 14607 18120
rect 14641 18086 14724 18120
rect 14539 18052 14724 18086
rect 14539 18018 14607 18052
rect 14641 18018 14724 18052
rect 14539 17984 14724 18018
rect 14539 17950 14607 17984
rect 14641 17950 14724 17984
rect 14539 17916 14724 17950
rect 14539 17882 14607 17916
rect 14641 17882 14724 17916
rect 14539 17848 14724 17882
rect 14539 17814 14607 17848
rect 14641 17814 14724 17848
rect 14539 17780 14724 17814
rect 14539 17746 14607 17780
rect 14641 17746 14724 17780
rect 14539 17712 14724 17746
rect 14539 17678 14607 17712
rect 14641 17678 14724 17712
rect 14539 17644 14724 17678
rect 14539 17610 14607 17644
rect 14641 17610 14724 17644
rect 14539 17576 14724 17610
rect 14539 17542 14607 17576
rect 14641 17542 14724 17576
rect 14539 17508 14724 17542
rect 14539 17474 14607 17508
rect 14641 17474 14724 17508
rect 14539 17440 14724 17474
rect 14539 17406 14607 17440
rect 14641 17406 14724 17440
rect 14539 17372 14724 17406
rect 14539 17338 14607 17372
rect 14641 17338 14724 17372
rect 14539 17304 14724 17338
rect 14539 17270 14607 17304
rect 14641 17270 14724 17304
rect 14539 17236 14724 17270
rect 14539 17202 14607 17236
rect 14641 17202 14724 17236
rect 14539 17168 14724 17202
rect 14539 17134 14607 17168
rect 14641 17134 14724 17168
rect 14539 17100 14724 17134
rect 14539 17066 14607 17100
rect 14641 17066 14724 17100
rect 14539 17032 14724 17066
rect 14539 16998 14607 17032
rect 14641 16998 14724 17032
rect 14539 16964 14724 16998
rect 14539 16930 14607 16964
rect 14641 16930 14724 16964
rect 14539 16896 14724 16930
rect 14539 16862 14607 16896
rect 14641 16862 14724 16896
rect 14539 16828 14724 16862
rect 14539 16794 14607 16828
rect 14641 16794 14724 16828
rect 14539 16760 14724 16794
rect 14539 16726 14607 16760
rect 14641 16726 14724 16760
rect 14539 16692 14724 16726
rect 14539 16658 14607 16692
rect 14641 16658 14724 16692
rect 14539 16624 14724 16658
rect 14539 16590 14607 16624
rect 14641 16590 14724 16624
rect 14539 16556 14724 16590
rect 14539 16522 14607 16556
rect 14641 16522 14724 16556
rect 14539 16488 14724 16522
rect 14539 16454 14607 16488
rect 14641 16454 14724 16488
rect 14539 16420 14724 16454
rect 14539 16386 14607 16420
rect 14641 16386 14724 16420
rect 14539 16352 14724 16386
rect 14539 16318 14607 16352
rect 14641 16318 14724 16352
rect 14539 16284 14724 16318
rect 14539 16250 14607 16284
rect 14641 16250 14724 16284
rect 14539 16216 14724 16250
rect 14539 16182 14607 16216
rect 14641 16182 14724 16216
rect 14539 16148 14724 16182
rect 14539 16114 14607 16148
rect 14641 16114 14724 16148
rect 14539 16080 14724 16114
rect 14539 16046 14607 16080
rect 14641 16046 14724 16080
rect 14539 16012 14724 16046
rect 14539 15978 14607 16012
rect 14641 15978 14724 16012
rect 14539 15944 14724 15978
rect 14539 15910 14607 15944
rect 14641 15910 14724 15944
rect 14539 15876 14724 15910
rect 14539 15842 14607 15876
rect 14641 15842 14724 15876
rect 14539 15808 14724 15842
rect 14539 15774 14607 15808
rect 14641 15774 14724 15808
rect 14539 15740 14724 15774
rect 14539 15706 14607 15740
rect 14641 15706 14724 15740
rect 14539 15672 14724 15706
rect 14539 15638 14607 15672
rect 14641 15638 14724 15672
rect 14539 15604 14724 15638
rect 14539 15570 14607 15604
rect 14641 15570 14724 15604
rect 14539 15536 14724 15570
rect 14539 15502 14607 15536
rect 14641 15502 14724 15536
rect 14539 15468 14724 15502
rect 14539 15434 14607 15468
rect 14641 15434 14724 15468
rect 14539 15400 14724 15434
rect 14539 15366 14607 15400
rect 14641 15366 14724 15400
rect 14539 15332 14724 15366
rect 14539 15298 14607 15332
rect 14641 15298 14724 15332
rect 14539 15264 14724 15298
rect 14539 15230 14607 15264
rect 14641 15230 14724 15264
rect 14539 15196 14724 15230
rect 14539 15162 14607 15196
rect 14641 15162 14724 15196
rect 14539 15128 14724 15162
rect 14539 15094 14607 15128
rect 14641 15094 14724 15128
rect 14539 15060 14724 15094
rect 14539 15026 14607 15060
rect 14641 15026 14724 15060
rect 14539 14992 14724 15026
rect 14539 14958 14607 14992
rect 14641 14958 14724 14992
rect 14539 14924 14724 14958
rect 14539 14890 14607 14924
rect 14641 14890 14724 14924
rect 14539 14856 14724 14890
rect 14539 14822 14607 14856
rect 14641 14822 14724 14856
rect 14539 14788 14724 14822
rect 14539 14754 14607 14788
rect 14641 14754 14724 14788
rect 14539 14720 14724 14754
rect 14539 14686 14607 14720
rect 14641 14686 14724 14720
rect 14539 14652 14724 14686
rect 14539 14618 14607 14652
rect 14641 14618 14724 14652
rect 14539 14584 14724 14618
rect 14539 14550 14607 14584
rect 14641 14550 14724 14584
rect 14539 14516 14724 14550
rect 14539 14482 14607 14516
rect 14641 14482 14724 14516
rect 14539 14448 14724 14482
rect 14539 14414 14607 14448
rect 14641 14414 14724 14448
rect 14539 14380 14724 14414
rect 14539 14346 14607 14380
rect 14641 14346 14724 14380
rect 14539 14312 14724 14346
rect 14539 14278 14607 14312
rect 14641 14278 14724 14312
rect 14539 14244 14724 14278
rect 14539 14210 14607 14244
rect 14641 14210 14724 14244
rect 14539 14176 14724 14210
rect 14539 14142 14607 14176
rect 14641 14142 14724 14176
rect 14539 14108 14724 14142
rect 14539 14074 14607 14108
rect 14641 14074 14724 14108
rect 14539 14040 14724 14074
rect 14539 14006 14607 14040
rect 14641 14006 14724 14040
rect 14539 13972 14724 14006
rect 14539 13938 14607 13972
rect 14641 13938 14724 13972
rect 14539 13904 14724 13938
rect 14539 13870 14607 13904
rect 14641 13870 14724 13904
rect 14539 13836 14724 13870
rect 14539 13802 14607 13836
rect 14641 13802 14724 13836
rect 14539 13768 14724 13802
rect 14539 13734 14607 13768
rect 14641 13734 14724 13768
rect 14539 13700 14724 13734
rect 14539 13666 14607 13700
rect 14641 13666 14724 13700
rect 14539 13632 14724 13666
rect 14539 13598 14607 13632
rect 14641 13598 14724 13632
rect 14539 13564 14724 13598
rect 14539 13530 14607 13564
rect 14641 13530 14724 13564
rect 14539 13496 14724 13530
rect 14539 13462 14607 13496
rect 14641 13462 14724 13496
rect 14539 13428 14724 13462
rect 14539 13394 14607 13428
rect 14641 13394 14724 13428
rect 14539 13360 14724 13394
rect 14539 13326 14607 13360
rect 14641 13326 14724 13360
rect 14539 13292 14724 13326
rect 14539 13258 14607 13292
rect 14641 13258 14724 13292
rect 14539 13224 14724 13258
rect 14539 13190 14607 13224
rect 14641 13190 14724 13224
rect 14539 13156 14724 13190
rect 14539 13122 14607 13156
rect 14641 13122 14724 13156
rect 14539 13088 14724 13122
rect 14539 13054 14607 13088
rect 14641 13054 14724 13088
rect 14539 13020 14724 13054
rect 14539 12986 14607 13020
rect 14641 12986 14724 13020
rect 14539 12952 14724 12986
rect 14539 12918 14607 12952
rect 14641 12918 14724 12952
rect 14539 12884 14724 12918
rect 14539 12850 14607 12884
rect 14641 12850 14724 12884
rect 14539 12816 14724 12850
rect 14539 12782 14607 12816
rect 14641 12782 14724 12816
rect 14539 12748 14724 12782
rect 14539 12714 14607 12748
rect 14641 12714 14724 12748
rect 14539 12680 14724 12714
rect 14539 12646 14607 12680
rect 14641 12646 14724 12680
rect 14539 12612 14724 12646
rect 14539 12578 14607 12612
rect 14641 12578 14724 12612
rect 14539 12544 14724 12578
rect 14539 12510 14607 12544
rect 14641 12510 14724 12544
rect 14539 12476 14724 12510
rect 14539 12442 14607 12476
rect 14641 12442 14724 12476
rect 14539 12408 14724 12442
rect 14539 12374 14607 12408
rect 14641 12374 14724 12408
rect 14539 12340 14724 12374
rect 14539 12306 14607 12340
rect 14641 12306 14724 12340
rect 14539 12272 14724 12306
rect 14539 12238 14607 12272
rect 14641 12238 14724 12272
rect 14539 12204 14724 12238
rect 14539 12170 14607 12204
rect 14641 12170 14724 12204
rect 14539 12136 14724 12170
rect 14539 12102 14607 12136
rect 14641 12102 14724 12136
rect 14539 12068 14724 12102
rect 14539 12034 14607 12068
rect 14641 12034 14724 12068
rect 14539 12000 14724 12034
rect 14539 11966 14607 12000
rect 14641 11966 14724 12000
rect 14539 11932 14724 11966
rect 14539 11898 14607 11932
rect 14641 11898 14724 11932
rect 14539 11864 14724 11898
rect 14539 11830 14607 11864
rect 14641 11830 14724 11864
rect 14539 11796 14724 11830
rect 14539 11762 14607 11796
rect 14641 11762 14724 11796
rect 14539 11728 14724 11762
rect 14539 11694 14607 11728
rect 14641 11694 14724 11728
rect 14539 11660 14724 11694
rect 14539 11626 14607 11660
rect 14641 11626 14724 11660
rect 14539 11592 14724 11626
rect 14539 11558 14607 11592
rect 14641 11558 14724 11592
rect 14539 11524 14724 11558
rect 14539 11490 14607 11524
rect 14641 11490 14724 11524
rect 14539 11456 14724 11490
rect 14539 11422 14607 11456
rect 14641 11422 14724 11456
rect 14539 11388 14724 11422
rect 14539 11354 14607 11388
rect 14641 11354 14724 11388
rect 14539 11320 14724 11354
rect 14539 11286 14607 11320
rect 14641 11286 14724 11320
rect 14539 11252 14724 11286
rect 14539 11218 14607 11252
rect 14641 11218 14724 11252
rect 14539 11184 14724 11218
rect 14539 11150 14607 11184
rect 14641 11150 14724 11184
rect 14539 11116 14724 11150
rect 14539 11082 14607 11116
rect 14641 11082 14724 11116
rect 14539 11048 14724 11082
rect 14539 11014 14607 11048
rect 14641 11014 14724 11048
rect 14539 10980 14724 11014
rect 14539 10946 14607 10980
rect 14641 10946 14724 10980
rect 14539 10912 14724 10946
rect 14539 10878 14607 10912
rect 14641 10878 14724 10912
rect 14539 10844 14724 10878
rect 14539 10810 14607 10844
rect 14641 10810 14724 10844
rect 14539 10776 14724 10810
rect 14539 10742 14607 10776
rect 14641 10742 14724 10776
rect 14539 10708 14724 10742
rect 14539 10674 14607 10708
rect 14641 10674 14724 10708
rect 14539 10640 14724 10674
rect 14539 10606 14607 10640
rect 14641 10606 14724 10640
rect 14539 10572 14724 10606
rect 14539 10538 14607 10572
rect 14641 10538 14724 10572
rect 14539 10504 14724 10538
rect 14539 10470 14607 10504
rect 14641 10470 14724 10504
rect 14539 10436 14724 10470
rect 14539 10402 14607 10436
rect 14641 10402 14724 10436
rect 14539 10368 14724 10402
rect 14539 10334 14607 10368
rect 14641 10334 14724 10368
rect 14539 10300 14724 10334
rect 14539 10266 14607 10300
rect 14641 10266 14724 10300
rect 14539 10232 14724 10266
rect 14539 10198 14607 10232
rect 14641 10198 14724 10232
rect 14539 10164 14724 10198
rect 14539 10130 14607 10164
rect 14641 10130 14724 10164
rect 14539 10096 14724 10130
rect 14539 10062 14607 10096
rect 14641 10062 14724 10096
rect 14539 10028 14724 10062
rect 14539 9994 14607 10028
rect 14641 9994 14724 10028
rect 14539 9960 14724 9994
rect 14539 9926 14607 9960
rect 14641 9926 14724 9960
rect 14539 9892 14724 9926
rect 14539 9858 14607 9892
rect 14641 9858 14724 9892
rect 14539 9824 14724 9858
rect 14539 9790 14607 9824
rect 14641 9790 14724 9824
rect 14539 9756 14724 9790
rect 14539 9722 14607 9756
rect 14641 9722 14724 9756
rect 245 9648 312 9682
rect 346 9648 430 9682
rect 245 9614 430 9648
rect 245 9580 312 9614
rect 346 9580 430 9614
rect 245 9528 430 9580
rect 14539 9688 14724 9722
rect 14539 9654 14607 9688
rect 14641 9654 14724 9688
rect 14539 9620 14724 9654
rect 14539 9586 14607 9620
rect 14641 9586 14724 9620
rect 14539 9528 14724 9586
rect 245 9451 14724 9528
rect 245 9417 476 9451
rect 510 9417 544 9451
rect 578 9417 612 9451
rect 646 9417 680 9451
rect 714 9417 748 9451
rect 782 9417 816 9451
rect 850 9417 884 9451
rect 918 9417 952 9451
rect 986 9417 1020 9451
rect 1054 9417 1088 9451
rect 1122 9417 1156 9451
rect 1190 9417 1224 9451
rect 1258 9417 1292 9451
rect 1326 9417 1360 9451
rect 1394 9417 1428 9451
rect 1462 9417 1496 9451
rect 1530 9417 1564 9451
rect 1598 9417 1632 9451
rect 1666 9417 1700 9451
rect 1734 9417 1768 9451
rect 1802 9417 1836 9451
rect 1870 9417 1904 9451
rect 1938 9417 1972 9451
rect 2006 9417 2040 9451
rect 2074 9417 2108 9451
rect 2142 9417 2176 9451
rect 2210 9417 2244 9451
rect 2278 9417 2312 9451
rect 2346 9417 2380 9451
rect 2414 9417 2448 9451
rect 2482 9417 2516 9451
rect 2550 9417 2584 9451
rect 2618 9417 2652 9451
rect 2686 9417 2720 9451
rect 2754 9417 2788 9451
rect 2822 9417 2856 9451
rect 2890 9417 2924 9451
rect 2958 9417 2992 9451
rect 3026 9417 3060 9451
rect 3094 9417 3128 9451
rect 3162 9417 3196 9451
rect 3230 9417 3264 9451
rect 3298 9417 3332 9451
rect 3366 9417 3400 9451
rect 3434 9417 3468 9451
rect 3502 9417 3536 9451
rect 3570 9417 3604 9451
rect 3638 9417 3672 9451
rect 3706 9417 3740 9451
rect 3774 9417 3808 9451
rect 3842 9417 3876 9451
rect 3910 9417 3944 9451
rect 3978 9417 4012 9451
rect 4046 9417 4080 9451
rect 4114 9417 4148 9451
rect 4182 9417 4216 9451
rect 4250 9417 4284 9451
rect 4318 9417 4352 9451
rect 4386 9417 4420 9451
rect 4454 9417 4488 9451
rect 4522 9417 4556 9451
rect 4590 9417 4624 9451
rect 4658 9417 4692 9451
rect 4726 9417 4760 9451
rect 4794 9417 4828 9451
rect 4862 9417 4896 9451
rect 4930 9417 4964 9451
rect 4998 9417 5032 9451
rect 5066 9417 5100 9451
rect 5134 9417 5168 9451
rect 5202 9417 5236 9451
rect 5270 9417 5304 9451
rect 5338 9417 5372 9451
rect 5406 9417 5440 9451
rect 5474 9417 5508 9451
rect 5542 9417 5576 9451
rect 5610 9417 5644 9451
rect 5678 9417 5712 9451
rect 5746 9417 5780 9451
rect 5814 9417 5848 9451
rect 5882 9417 5916 9451
rect 5950 9417 5984 9451
rect 6018 9417 6052 9451
rect 6086 9417 6120 9451
rect 6154 9417 6188 9451
rect 6222 9417 6256 9451
rect 6290 9417 6324 9451
rect 6358 9417 6392 9451
rect 6426 9417 6460 9451
rect 6494 9417 6528 9451
rect 6562 9417 6596 9451
rect 6630 9417 6664 9451
rect 6698 9417 6732 9451
rect 6766 9417 6800 9451
rect 6834 9417 6868 9451
rect 6902 9417 6936 9451
rect 6970 9417 7004 9451
rect 7038 9417 7072 9451
rect 7106 9417 7140 9451
rect 7174 9417 7208 9451
rect 7242 9417 7276 9451
rect 7310 9417 7344 9451
rect 7378 9417 7412 9451
rect 7446 9417 7480 9451
rect 7514 9417 7548 9451
rect 7582 9417 7616 9451
rect 7650 9417 7684 9451
rect 7718 9417 7752 9451
rect 7786 9417 7820 9451
rect 7854 9417 7888 9451
rect 7922 9417 7956 9451
rect 7990 9417 8024 9451
rect 8058 9417 8092 9451
rect 8126 9417 8160 9451
rect 8194 9417 8228 9451
rect 8262 9417 8296 9451
rect 8330 9417 8364 9451
rect 8398 9417 8432 9451
rect 8466 9417 8500 9451
rect 8534 9417 8568 9451
rect 8602 9417 8636 9451
rect 8670 9417 8704 9451
rect 8738 9417 8772 9451
rect 8806 9417 8840 9451
rect 8874 9417 8908 9451
rect 8942 9417 8976 9451
rect 9010 9417 9044 9451
rect 9078 9417 9112 9451
rect 9146 9417 9180 9451
rect 9214 9417 9248 9451
rect 9282 9417 9316 9451
rect 9350 9417 9384 9451
rect 9418 9417 9452 9451
rect 9486 9417 9520 9451
rect 9554 9417 9588 9451
rect 9622 9417 9656 9451
rect 9690 9417 9724 9451
rect 9758 9417 9792 9451
rect 9826 9417 9860 9451
rect 9894 9417 9928 9451
rect 9962 9417 9996 9451
rect 10030 9417 10064 9451
rect 10098 9417 10132 9451
rect 10166 9417 10200 9451
rect 10234 9417 10268 9451
rect 10302 9417 10336 9451
rect 10370 9417 10404 9451
rect 10438 9417 10472 9451
rect 10506 9417 10540 9451
rect 10574 9417 10608 9451
rect 10642 9417 10676 9451
rect 10710 9417 10744 9451
rect 10778 9417 10812 9451
rect 10846 9417 10880 9451
rect 10914 9417 10948 9451
rect 10982 9417 11016 9451
rect 11050 9417 11084 9451
rect 11118 9417 11152 9451
rect 11186 9417 11220 9451
rect 11254 9417 11288 9451
rect 11322 9417 11356 9451
rect 11390 9417 11424 9451
rect 11458 9417 11492 9451
rect 11526 9417 11560 9451
rect 11594 9417 11628 9451
rect 11662 9417 11696 9451
rect 11730 9417 11764 9451
rect 11798 9417 11832 9451
rect 11866 9417 11900 9451
rect 11934 9417 11968 9451
rect 12002 9417 12036 9451
rect 12070 9417 12104 9451
rect 12138 9417 12172 9451
rect 12206 9417 12240 9451
rect 12274 9417 12308 9451
rect 12342 9417 12376 9451
rect 12410 9417 12444 9451
rect 12478 9417 12512 9451
rect 12546 9417 12580 9451
rect 12614 9417 12648 9451
rect 12682 9417 12716 9451
rect 12750 9417 12784 9451
rect 12818 9417 12852 9451
rect 12886 9417 12920 9451
rect 12954 9417 12988 9451
rect 13022 9417 13056 9451
rect 13090 9417 13124 9451
rect 13158 9417 13192 9451
rect 13226 9417 13260 9451
rect 13294 9417 13328 9451
rect 13362 9417 13396 9451
rect 13430 9417 13464 9451
rect 13498 9417 13532 9451
rect 13566 9417 13600 9451
rect 13634 9417 13668 9451
rect 13702 9417 13736 9451
rect 13770 9417 13804 9451
rect 13838 9417 13872 9451
rect 13906 9417 13940 9451
rect 13974 9417 14008 9451
rect 14042 9417 14076 9451
rect 14110 9417 14144 9451
rect 14178 9417 14212 9451
rect 14246 9417 14280 9451
rect 14314 9417 14348 9451
rect 14382 9417 14416 9451
rect 14450 9417 14484 9451
rect 14518 9417 14724 9451
rect 245 9343 14724 9417
<< mvnsubdiff >>
rect 583 36177 14381 36227
rect 583 36143 766 36177
rect 800 36143 834 36177
rect 868 36143 902 36177
rect 936 36143 970 36177
rect 1004 36143 1038 36177
rect 1072 36143 1106 36177
rect 1140 36143 1174 36177
rect 1208 36143 1242 36177
rect 1276 36143 1310 36177
rect 1344 36143 1378 36177
rect 1412 36143 1446 36177
rect 1480 36143 1514 36177
rect 1548 36143 1582 36177
rect 1616 36143 1650 36177
rect 1684 36143 1718 36177
rect 1752 36143 1786 36177
rect 1820 36143 1854 36177
rect 1888 36143 1922 36177
rect 1956 36143 1990 36177
rect 2024 36143 2058 36177
rect 2092 36143 2126 36177
rect 2160 36143 2194 36177
rect 2228 36143 2262 36177
rect 2296 36143 2330 36177
rect 2364 36143 2398 36177
rect 2432 36143 2466 36177
rect 2500 36143 2534 36177
rect 2568 36143 2602 36177
rect 2636 36143 2670 36177
rect 2704 36143 2738 36177
rect 2772 36143 2806 36177
rect 2840 36143 2874 36177
rect 2908 36143 2942 36177
rect 2976 36143 3010 36177
rect 3044 36143 3078 36177
rect 3112 36143 3146 36177
rect 3180 36143 3214 36177
rect 3248 36143 3282 36177
rect 3316 36143 3350 36177
rect 3384 36143 3418 36177
rect 3452 36143 3486 36177
rect 3520 36143 3554 36177
rect 3588 36143 3622 36177
rect 3656 36143 3690 36177
rect 3724 36143 3758 36177
rect 3792 36143 3826 36177
rect 3860 36143 3894 36177
rect 3928 36143 3962 36177
rect 3996 36143 4030 36177
rect 4064 36143 4098 36177
rect 4132 36143 4166 36177
rect 4200 36143 4234 36177
rect 4268 36143 4302 36177
rect 4336 36143 4370 36177
rect 4404 36143 4438 36177
rect 4472 36143 4506 36177
rect 4540 36143 4574 36177
rect 4608 36143 4642 36177
rect 4676 36143 4710 36177
rect 4744 36143 4778 36177
rect 4812 36143 4846 36177
rect 4880 36143 4914 36177
rect 4948 36143 4982 36177
rect 5016 36143 5050 36177
rect 5084 36143 5118 36177
rect 5152 36143 5186 36177
rect 5220 36143 5254 36177
rect 5288 36143 5322 36177
rect 5356 36143 5390 36177
rect 5424 36143 5458 36177
rect 5492 36143 5526 36177
rect 5560 36143 5594 36177
rect 5628 36143 5662 36177
rect 5696 36143 5730 36177
rect 5764 36143 5798 36177
rect 5832 36143 5866 36177
rect 5900 36143 5934 36177
rect 5968 36143 6002 36177
rect 6036 36143 6070 36177
rect 6104 36143 6138 36177
rect 6172 36143 6206 36177
rect 6240 36143 6274 36177
rect 6308 36143 6342 36177
rect 6376 36143 6410 36177
rect 6444 36143 6478 36177
rect 6512 36143 6546 36177
rect 6580 36143 6614 36177
rect 6648 36143 6682 36177
rect 6716 36143 6750 36177
rect 6784 36143 6818 36177
rect 6852 36143 6886 36177
rect 6920 36143 6954 36177
rect 6988 36143 7022 36177
rect 7056 36143 7090 36177
rect 7124 36143 7158 36177
rect 7192 36143 7226 36177
rect 7260 36143 7294 36177
rect 7328 36143 7362 36177
rect 7396 36143 7430 36177
rect 7464 36143 7498 36177
rect 7532 36143 7566 36177
rect 7600 36143 7634 36177
rect 7668 36143 7702 36177
rect 7736 36143 7770 36177
rect 7804 36143 7838 36177
rect 7872 36143 7906 36177
rect 7940 36143 7974 36177
rect 8008 36143 8042 36177
rect 8076 36143 8110 36177
rect 8144 36143 8178 36177
rect 8212 36143 8246 36177
rect 8280 36143 8314 36177
rect 8348 36143 8382 36177
rect 8416 36143 8450 36177
rect 8484 36143 8518 36177
rect 8552 36143 8586 36177
rect 8620 36143 8654 36177
rect 8688 36143 8722 36177
rect 8756 36143 8790 36177
rect 8824 36143 8858 36177
rect 8892 36143 8926 36177
rect 8960 36143 8994 36177
rect 9028 36143 9062 36177
rect 9096 36143 9130 36177
rect 9164 36143 9198 36177
rect 9232 36143 9266 36177
rect 9300 36143 9334 36177
rect 9368 36143 9402 36177
rect 9436 36143 9470 36177
rect 9504 36143 9538 36177
rect 9572 36143 9606 36177
rect 9640 36143 9674 36177
rect 9708 36143 9742 36177
rect 9776 36143 9810 36177
rect 9844 36143 9878 36177
rect 9912 36143 9946 36177
rect 9980 36143 10014 36177
rect 10048 36143 10082 36177
rect 10116 36143 10150 36177
rect 10184 36143 10218 36177
rect 10252 36143 10286 36177
rect 10320 36143 10354 36177
rect 10388 36143 10422 36177
rect 10456 36143 10490 36177
rect 10524 36143 10558 36177
rect 10592 36143 10626 36177
rect 10660 36143 10694 36177
rect 10728 36143 10762 36177
rect 10796 36143 10830 36177
rect 10864 36143 10898 36177
rect 10932 36143 10966 36177
rect 11000 36143 11034 36177
rect 11068 36143 11102 36177
rect 11136 36143 11170 36177
rect 11204 36143 11238 36177
rect 11272 36143 11306 36177
rect 11340 36143 11374 36177
rect 11408 36143 11442 36177
rect 11476 36143 11510 36177
rect 11544 36143 11578 36177
rect 11612 36143 11646 36177
rect 11680 36143 11714 36177
rect 11748 36143 11782 36177
rect 11816 36143 11850 36177
rect 11884 36143 11918 36177
rect 11952 36143 11986 36177
rect 12020 36143 12054 36177
rect 12088 36143 12122 36177
rect 12156 36143 12190 36177
rect 12224 36143 12258 36177
rect 12292 36143 12326 36177
rect 12360 36143 12394 36177
rect 12428 36143 12462 36177
rect 12496 36143 12530 36177
rect 12564 36143 12598 36177
rect 12632 36143 12666 36177
rect 12700 36143 12734 36177
rect 12768 36143 12802 36177
rect 12836 36143 12870 36177
rect 12904 36143 12938 36177
rect 12972 36143 13006 36177
rect 13040 36143 13074 36177
rect 13108 36143 13142 36177
rect 13176 36143 13210 36177
rect 13244 36143 13278 36177
rect 13312 36143 13346 36177
rect 13380 36143 13414 36177
rect 13448 36143 13482 36177
rect 13516 36143 13550 36177
rect 13584 36143 13618 36177
rect 13652 36143 13686 36177
rect 13720 36143 13754 36177
rect 13788 36143 13822 36177
rect 13856 36143 13890 36177
rect 13924 36143 13958 36177
rect 13992 36143 14026 36177
rect 14060 36143 14094 36177
rect 14128 36143 14162 36177
rect 14196 36143 14381 36177
rect 583 36093 14381 36143
rect 583 36032 715 36093
rect 583 35998 632 36032
rect 666 35998 715 36032
rect 583 35964 715 35998
rect 583 35930 632 35964
rect 666 35930 715 35964
rect 583 35896 715 35930
rect 583 35862 632 35896
rect 666 35862 715 35896
rect 583 35828 715 35862
rect 583 35794 632 35828
rect 666 35794 715 35828
rect 583 35760 715 35794
rect 583 35726 632 35760
rect 666 35726 715 35760
rect 583 35692 715 35726
rect 583 35658 632 35692
rect 666 35658 715 35692
rect 583 35624 715 35658
rect 583 35590 632 35624
rect 666 35590 715 35624
rect 583 35556 715 35590
rect 583 35522 632 35556
rect 666 35522 715 35556
rect 583 35488 715 35522
rect 583 35454 632 35488
rect 666 35454 715 35488
rect 583 35420 715 35454
rect 583 35386 632 35420
rect 666 35386 715 35420
rect 583 35352 715 35386
rect 583 35318 632 35352
rect 666 35318 715 35352
rect 583 35284 715 35318
rect 583 35250 632 35284
rect 666 35250 715 35284
rect 583 35216 715 35250
rect 583 35182 632 35216
rect 666 35182 715 35216
rect 583 35148 715 35182
rect 583 35114 632 35148
rect 666 35114 715 35148
rect 583 35080 715 35114
rect 583 35046 632 35080
rect 666 35046 715 35080
rect 583 35012 715 35046
rect 583 34978 632 35012
rect 666 34978 715 35012
rect 583 34944 715 34978
rect 583 34910 632 34944
rect 666 34910 715 34944
rect 583 34876 715 34910
rect 583 34842 632 34876
rect 666 34842 715 34876
rect 583 34808 715 34842
rect 583 34774 632 34808
rect 666 34774 715 34808
rect 583 34740 715 34774
rect 583 34706 632 34740
rect 666 34706 715 34740
rect 14247 36032 14381 36093
rect 14247 35998 14297 36032
rect 14331 35998 14381 36032
rect 14247 35964 14381 35998
rect 14247 35930 14297 35964
rect 14331 35930 14381 35964
rect 14247 35896 14381 35930
rect 14247 35862 14297 35896
rect 14331 35862 14381 35896
rect 14247 35828 14381 35862
rect 14247 35794 14297 35828
rect 14331 35794 14381 35828
rect 14247 35760 14381 35794
rect 14247 35726 14297 35760
rect 14331 35726 14381 35760
rect 14247 35692 14381 35726
rect 14247 35658 14297 35692
rect 14331 35658 14381 35692
rect 14247 35624 14381 35658
rect 14247 35590 14297 35624
rect 14331 35590 14381 35624
rect 14247 35556 14381 35590
rect 14247 35522 14297 35556
rect 14331 35522 14381 35556
rect 14247 35488 14381 35522
rect 14247 35454 14297 35488
rect 14331 35454 14381 35488
rect 14247 35420 14381 35454
rect 14247 35386 14297 35420
rect 14331 35386 14381 35420
rect 14247 35352 14381 35386
rect 14247 35318 14297 35352
rect 14331 35318 14381 35352
rect 14247 35284 14381 35318
rect 14247 35250 14297 35284
rect 14331 35250 14381 35284
rect 14247 35216 14381 35250
rect 14247 35182 14297 35216
rect 14331 35182 14381 35216
rect 14247 35148 14381 35182
rect 14247 35114 14297 35148
rect 14331 35114 14381 35148
rect 14247 35080 14381 35114
rect 14247 35046 14297 35080
rect 14331 35046 14381 35080
rect 14247 35012 14381 35046
rect 14247 34978 14297 35012
rect 14331 34978 14381 35012
rect 14247 34944 14381 34978
rect 14247 34910 14297 34944
rect 14331 34910 14381 34944
rect 14247 34876 14381 34910
rect 14247 34842 14297 34876
rect 14331 34842 14381 34876
rect 14247 34808 14381 34842
rect 14247 34774 14297 34808
rect 14331 34774 14381 34808
rect 14247 34740 14381 34774
rect 583 34672 715 34706
rect 583 34638 632 34672
rect 666 34638 715 34672
rect 583 34604 715 34638
rect 583 34570 632 34604
rect 666 34570 715 34604
rect 583 34536 715 34570
rect 583 34502 632 34536
rect 666 34502 715 34536
rect 583 34468 715 34502
rect 583 34434 632 34468
rect 666 34434 715 34468
rect 583 34400 715 34434
rect 583 34366 632 34400
rect 666 34366 715 34400
rect 583 34332 715 34366
rect 583 34298 632 34332
rect 666 34298 715 34332
rect 583 34264 715 34298
rect 583 34230 632 34264
rect 666 34230 715 34264
rect 583 34196 715 34230
rect 583 34162 632 34196
rect 666 34162 715 34196
rect 583 34128 715 34162
rect 583 34094 632 34128
rect 666 34094 715 34128
rect 583 34060 715 34094
rect 583 34026 632 34060
rect 666 34026 715 34060
rect 583 33992 715 34026
rect 583 33958 632 33992
rect 666 33958 715 33992
rect 583 33924 715 33958
rect 583 33890 632 33924
rect 666 33890 715 33924
rect 583 33856 715 33890
rect 583 33822 632 33856
rect 666 33822 715 33856
rect 583 33788 715 33822
rect 583 33754 632 33788
rect 666 33754 715 33788
rect 583 33720 715 33754
rect 583 33686 632 33720
rect 666 33686 715 33720
rect 583 33652 715 33686
rect 583 33618 632 33652
rect 666 33618 715 33652
rect 583 33584 715 33618
rect 583 33550 632 33584
rect 666 33550 715 33584
rect 583 33516 715 33550
rect 583 33482 632 33516
rect 666 33482 715 33516
rect 583 33448 715 33482
rect 583 33414 632 33448
rect 666 33414 715 33448
rect 583 33380 715 33414
rect 583 33346 632 33380
rect 666 33346 715 33380
rect 583 33312 715 33346
rect 583 33278 632 33312
rect 666 33278 715 33312
rect 583 33244 715 33278
rect 583 33210 632 33244
rect 666 33210 715 33244
rect 583 33176 715 33210
rect 583 33142 632 33176
rect 666 33142 715 33176
rect 583 33108 715 33142
rect 583 33074 632 33108
rect 666 33074 715 33108
rect 583 33040 715 33074
rect 583 33006 632 33040
rect 666 33006 715 33040
rect 583 32972 715 33006
rect 583 32938 632 32972
rect 666 32938 715 32972
rect 583 32904 715 32938
rect 583 32870 632 32904
rect 666 32870 715 32904
rect 583 32836 715 32870
rect 583 32802 632 32836
rect 666 32802 715 32836
rect 583 32768 715 32802
rect 583 32734 632 32768
rect 666 32734 715 32768
rect 583 32700 715 32734
rect 583 32666 632 32700
rect 666 32666 715 32700
rect 583 32632 715 32666
rect 583 32598 632 32632
rect 666 32598 715 32632
rect 583 32564 715 32598
rect 583 32530 632 32564
rect 666 32530 715 32564
rect 583 32496 715 32530
rect 583 32462 632 32496
rect 666 32462 715 32496
rect 583 32428 715 32462
rect 583 32394 632 32428
rect 666 32394 715 32428
rect 583 32360 715 32394
rect 583 32326 632 32360
rect 666 32326 715 32360
rect 583 32292 715 32326
rect 583 32258 632 32292
rect 666 32258 715 32292
rect 583 32224 715 32258
rect 583 32190 632 32224
rect 666 32190 715 32224
rect 583 32156 715 32190
rect 583 32122 632 32156
rect 666 32122 715 32156
rect 583 32088 715 32122
rect 583 32054 632 32088
rect 666 32054 715 32088
rect 583 32020 715 32054
rect 583 31986 632 32020
rect 666 31986 715 32020
rect 583 31952 715 31986
rect 583 31918 632 31952
rect 666 31918 715 31952
rect 583 31884 715 31918
rect 583 31850 632 31884
rect 666 31850 715 31884
rect 583 31816 715 31850
rect 583 31782 632 31816
rect 666 31782 715 31816
rect 583 31748 715 31782
rect 583 31714 632 31748
rect 666 31714 715 31748
rect 583 31680 715 31714
rect 583 31646 632 31680
rect 666 31646 715 31680
rect 583 31612 715 31646
rect 583 31578 632 31612
rect 666 31578 715 31612
rect 583 31544 715 31578
rect 583 31510 632 31544
rect 666 31510 715 31544
rect 583 31476 715 31510
rect 583 31442 632 31476
rect 666 31442 715 31476
rect 583 31408 715 31442
rect 583 31374 632 31408
rect 666 31374 715 31408
rect 583 31340 715 31374
rect 583 31306 632 31340
rect 666 31306 715 31340
rect 583 31272 715 31306
rect 583 31238 632 31272
rect 666 31238 715 31272
rect 583 31204 715 31238
rect 583 31170 632 31204
rect 666 31170 715 31204
rect 583 31136 715 31170
rect 583 31102 632 31136
rect 666 31102 715 31136
rect 583 31068 715 31102
rect 583 31034 632 31068
rect 666 31034 715 31068
rect 583 31000 715 31034
rect 583 30966 632 31000
rect 666 30966 715 31000
rect 583 30932 715 30966
rect 583 30898 632 30932
rect 666 30898 715 30932
rect 583 30864 715 30898
rect 583 30830 632 30864
rect 666 30830 715 30864
rect 583 30796 715 30830
rect 583 30762 632 30796
rect 666 30762 715 30796
rect 583 30728 715 30762
rect 583 30694 632 30728
rect 666 30694 715 30728
rect 583 30660 715 30694
rect 583 30626 632 30660
rect 666 30626 715 30660
rect 583 30592 715 30626
rect 583 30558 632 30592
rect 666 30558 715 30592
rect 583 30524 715 30558
rect 583 30490 632 30524
rect 666 30490 715 30524
rect 583 30456 715 30490
rect 583 30422 632 30456
rect 666 30422 715 30456
rect 583 30388 715 30422
rect 583 30354 632 30388
rect 666 30354 715 30388
rect 583 30320 715 30354
rect 583 30286 632 30320
rect 666 30286 715 30320
rect 583 30252 715 30286
rect 583 30218 632 30252
rect 666 30218 715 30252
rect 583 30184 715 30218
rect 583 30150 632 30184
rect 666 30150 715 30184
rect 583 30116 715 30150
rect 583 30082 632 30116
rect 666 30082 715 30116
rect 583 30048 715 30082
rect 583 30014 632 30048
rect 666 30014 715 30048
rect 583 29980 715 30014
rect 583 29946 632 29980
rect 666 29946 715 29980
rect 583 29912 715 29946
rect 583 29878 632 29912
rect 666 29878 715 29912
rect 583 29844 715 29878
rect 583 29810 632 29844
rect 666 29810 715 29844
rect 583 29776 715 29810
rect 583 29742 632 29776
rect 666 29742 715 29776
rect 583 29708 715 29742
rect 583 29674 632 29708
rect 666 29674 715 29708
rect 583 29640 715 29674
rect 583 29606 632 29640
rect 666 29606 715 29640
rect 583 29572 715 29606
rect 583 29538 632 29572
rect 666 29538 715 29572
rect 583 29504 715 29538
rect 583 29470 632 29504
rect 666 29470 715 29504
rect 583 29436 715 29470
rect 583 29402 632 29436
rect 666 29402 715 29436
rect 583 29368 715 29402
rect 583 29334 632 29368
rect 666 29334 715 29368
rect 583 29300 715 29334
rect 583 29266 632 29300
rect 666 29266 715 29300
rect 583 29232 715 29266
rect 583 29198 632 29232
rect 666 29198 715 29232
rect 583 29164 715 29198
rect 583 29130 632 29164
rect 666 29130 715 29164
rect 583 29096 715 29130
rect 583 29062 632 29096
rect 666 29062 715 29096
rect 583 29028 715 29062
rect 583 28994 632 29028
rect 666 28994 715 29028
rect 583 28960 715 28994
rect 583 28926 632 28960
rect 666 28926 715 28960
rect 583 28892 715 28926
rect 583 28858 632 28892
rect 666 28858 715 28892
rect 583 28824 715 28858
rect 583 28790 632 28824
rect 666 28790 715 28824
rect 583 28756 715 28790
rect 583 28722 632 28756
rect 666 28722 715 28756
rect 583 28688 715 28722
rect 583 28654 632 28688
rect 666 28654 715 28688
rect 583 28620 715 28654
rect 583 28586 632 28620
rect 666 28586 715 28620
rect 583 28552 715 28586
rect 583 28518 632 28552
rect 666 28518 715 28552
rect 583 28484 715 28518
rect 583 28450 632 28484
rect 666 28450 715 28484
rect 583 28416 715 28450
rect 583 28382 632 28416
rect 666 28382 715 28416
rect 583 28348 715 28382
rect 583 28314 632 28348
rect 666 28314 715 28348
rect 583 28280 715 28314
rect 583 28246 632 28280
rect 666 28246 715 28280
rect 583 28212 715 28246
rect 583 28178 632 28212
rect 666 28178 715 28212
rect 583 28144 715 28178
rect 583 28110 632 28144
rect 666 28110 715 28144
rect 583 28076 715 28110
rect 583 28042 632 28076
rect 666 28042 715 28076
rect 583 28008 715 28042
rect 583 27974 632 28008
rect 666 27974 715 28008
rect 583 27940 715 27974
rect 583 27906 632 27940
rect 666 27906 715 27940
rect 583 27872 715 27906
rect 583 27838 632 27872
rect 666 27838 715 27872
rect 583 27804 715 27838
rect 583 27770 632 27804
rect 666 27770 715 27804
rect 583 27736 715 27770
rect 583 27702 632 27736
rect 666 27702 715 27736
rect 583 27668 715 27702
rect 583 27634 632 27668
rect 666 27634 715 27668
rect 583 27600 715 27634
rect 583 27566 632 27600
rect 666 27566 715 27600
rect 583 27532 715 27566
rect 583 27498 632 27532
rect 666 27498 715 27532
rect 583 27464 715 27498
rect 583 27430 632 27464
rect 666 27430 715 27464
rect 583 27396 715 27430
rect 583 27362 632 27396
rect 666 27362 715 27396
rect 583 27328 715 27362
rect 583 27294 632 27328
rect 666 27294 715 27328
rect 583 27260 715 27294
rect 583 27226 632 27260
rect 666 27226 715 27260
rect 583 27192 715 27226
rect 583 27158 632 27192
rect 666 27158 715 27192
rect 583 27124 715 27158
rect 583 27090 632 27124
rect 666 27090 715 27124
rect 583 27056 715 27090
rect 583 27022 632 27056
rect 666 27022 715 27056
rect 583 26988 715 27022
rect 583 26954 632 26988
rect 666 26954 715 26988
rect 583 26920 715 26954
rect 583 26886 632 26920
rect 666 26886 715 26920
rect 583 26852 715 26886
rect 583 26818 632 26852
rect 666 26818 715 26852
rect 583 26784 715 26818
rect 583 26750 632 26784
rect 666 26750 715 26784
rect 583 26716 715 26750
rect 583 26682 632 26716
rect 666 26682 715 26716
rect 583 26648 715 26682
rect 583 26614 632 26648
rect 666 26614 715 26648
rect 583 26580 715 26614
rect 583 26546 632 26580
rect 666 26546 715 26580
rect 583 26512 715 26546
rect 583 26478 632 26512
rect 666 26478 715 26512
rect 583 26444 715 26478
rect 583 26410 632 26444
rect 666 26410 715 26444
rect 583 26376 715 26410
rect 583 26342 632 26376
rect 666 26342 715 26376
rect 583 26308 715 26342
rect 583 26274 632 26308
rect 666 26274 715 26308
rect 583 26240 715 26274
rect 583 26206 632 26240
rect 666 26206 715 26240
rect 583 26172 715 26206
rect 583 26138 632 26172
rect 666 26138 715 26172
rect 583 26104 715 26138
rect 583 26070 632 26104
rect 666 26070 715 26104
rect 583 26036 715 26070
rect 583 26002 632 26036
rect 666 26002 715 26036
rect 583 25968 715 26002
rect 583 25934 632 25968
rect 666 25934 715 25968
rect 583 25900 715 25934
rect 583 25866 632 25900
rect 666 25866 715 25900
rect 583 25832 715 25866
rect 583 25798 632 25832
rect 666 25798 715 25832
rect 583 25764 715 25798
rect 583 25730 632 25764
rect 666 25730 715 25764
rect 583 25696 715 25730
rect 583 25662 632 25696
rect 666 25662 715 25696
rect 583 25628 715 25662
rect 583 25594 632 25628
rect 666 25594 715 25628
rect 583 25560 715 25594
rect 583 25526 632 25560
rect 666 25526 715 25560
rect 583 25492 715 25526
rect 583 25458 632 25492
rect 666 25458 715 25492
rect 583 25424 715 25458
rect 583 25390 632 25424
rect 666 25390 715 25424
rect 583 25356 715 25390
rect 583 25322 632 25356
rect 666 25322 715 25356
rect 583 25288 715 25322
rect 583 25254 632 25288
rect 666 25254 715 25288
rect 583 25220 715 25254
rect 583 25186 632 25220
rect 666 25186 715 25220
rect 583 25152 715 25186
rect 583 25118 632 25152
rect 666 25118 715 25152
rect 583 25084 715 25118
rect 583 25050 632 25084
rect 666 25050 715 25084
rect 583 25016 715 25050
rect 583 24982 632 25016
rect 666 24982 715 25016
rect 583 24948 715 24982
rect 583 24914 632 24948
rect 666 24914 715 24948
rect 583 24880 715 24914
rect 583 24846 632 24880
rect 666 24846 715 24880
rect 583 24812 715 24846
rect 583 24778 632 24812
rect 666 24778 715 24812
rect 583 24744 715 24778
rect 583 24710 632 24744
rect 666 24710 715 24744
rect 583 24676 715 24710
rect 583 24642 632 24676
rect 666 24642 715 24676
rect 583 24608 715 24642
rect 583 24574 632 24608
rect 666 24574 715 24608
rect 583 24540 715 24574
rect 583 24506 632 24540
rect 666 24506 715 24540
rect 583 24472 715 24506
rect 583 24438 632 24472
rect 666 24438 715 24472
rect 583 24404 715 24438
rect 583 24370 632 24404
rect 666 24370 715 24404
rect 583 24336 715 24370
rect 583 24302 632 24336
rect 666 24302 715 24336
rect 583 24268 715 24302
rect 583 24234 632 24268
rect 666 24234 715 24268
rect 583 24200 715 24234
rect 583 24166 632 24200
rect 666 24166 715 24200
rect 583 24132 715 24166
rect 583 24098 632 24132
rect 666 24098 715 24132
rect 583 24064 715 24098
rect 583 24030 632 24064
rect 666 24030 715 24064
rect 583 23996 715 24030
rect 583 23962 632 23996
rect 666 23962 715 23996
rect 583 23928 715 23962
rect 583 23894 632 23928
rect 666 23894 715 23928
rect 583 23860 715 23894
rect 583 23826 632 23860
rect 666 23826 715 23860
rect 583 23792 715 23826
rect 583 23758 632 23792
rect 666 23758 715 23792
rect 583 23724 715 23758
rect 583 23690 632 23724
rect 666 23690 715 23724
rect 583 23656 715 23690
rect 583 23622 632 23656
rect 666 23622 715 23656
rect 583 23588 715 23622
rect 583 23554 632 23588
rect 666 23554 715 23588
rect 583 23520 715 23554
rect 583 23486 632 23520
rect 666 23486 715 23520
rect 583 23452 715 23486
rect 583 23418 632 23452
rect 666 23418 715 23452
rect 583 23384 715 23418
rect 583 23350 632 23384
rect 666 23350 715 23384
rect 583 23316 715 23350
rect 583 23282 632 23316
rect 666 23282 715 23316
rect 583 23248 715 23282
rect 583 23214 632 23248
rect 666 23214 715 23248
rect 583 23180 715 23214
rect 583 23146 632 23180
rect 666 23146 715 23180
rect 583 23112 715 23146
rect 583 23078 632 23112
rect 666 23078 715 23112
rect 583 23044 715 23078
rect 583 23010 632 23044
rect 666 23010 715 23044
rect 583 22976 715 23010
rect 583 22942 632 22976
rect 666 22942 715 22976
rect 583 22908 715 22942
rect 583 22874 632 22908
rect 666 22874 715 22908
rect 583 22840 715 22874
rect 583 22806 632 22840
rect 666 22806 715 22840
rect 583 22772 715 22806
rect 583 22738 632 22772
rect 666 22738 715 22772
rect 583 22704 715 22738
rect 583 22670 632 22704
rect 666 22670 715 22704
rect 583 22636 715 22670
rect 583 22602 632 22636
rect 666 22602 715 22636
rect 583 22568 715 22602
rect 583 22534 632 22568
rect 666 22534 715 22568
rect 583 22500 715 22534
rect 583 22466 632 22500
rect 666 22466 715 22500
rect 583 22432 715 22466
rect 583 22398 632 22432
rect 666 22398 715 22432
rect 583 22364 715 22398
rect 583 22330 632 22364
rect 666 22330 715 22364
rect 583 22296 715 22330
rect 583 22262 632 22296
rect 666 22262 715 22296
rect 583 22228 715 22262
rect 583 22194 632 22228
rect 666 22194 715 22228
rect 583 22160 715 22194
rect 583 22126 632 22160
rect 666 22126 715 22160
rect 583 22092 715 22126
rect 583 22058 632 22092
rect 666 22058 715 22092
rect 583 22024 715 22058
rect 583 21990 632 22024
rect 666 21990 715 22024
rect 583 21956 715 21990
rect 583 21922 632 21956
rect 666 21922 715 21956
rect 583 21888 715 21922
rect 583 21854 632 21888
rect 666 21854 715 21888
rect 583 21820 715 21854
rect 583 21786 632 21820
rect 666 21786 715 21820
rect 583 21752 715 21786
rect 583 21718 632 21752
rect 666 21718 715 21752
rect 583 21684 715 21718
rect 583 21650 632 21684
rect 666 21650 715 21684
rect 583 21616 715 21650
rect 583 21582 632 21616
rect 666 21582 715 21616
rect 583 21548 715 21582
rect 583 21514 632 21548
rect 666 21514 715 21548
rect 583 21480 715 21514
rect 583 21446 632 21480
rect 666 21446 715 21480
rect 583 21412 715 21446
rect 583 21378 632 21412
rect 666 21378 715 21412
rect 583 21344 715 21378
rect 583 21310 632 21344
rect 666 21310 715 21344
rect 583 21276 715 21310
rect 583 21242 632 21276
rect 666 21242 715 21276
rect 583 21208 715 21242
rect 583 21174 632 21208
rect 666 21174 715 21208
rect 583 21140 715 21174
rect 583 21106 632 21140
rect 666 21106 715 21140
rect 583 21072 715 21106
rect 583 21038 632 21072
rect 666 21038 715 21072
rect 583 21004 715 21038
rect 583 20970 632 21004
rect 666 20970 715 21004
rect 583 20936 715 20970
rect 583 20902 632 20936
rect 666 20902 715 20936
rect 583 20868 715 20902
rect 583 20834 632 20868
rect 666 20834 715 20868
rect 583 20800 715 20834
rect 583 20766 632 20800
rect 666 20766 715 20800
rect 583 20732 715 20766
rect 583 20698 632 20732
rect 666 20698 715 20732
rect 583 20664 715 20698
rect 583 20630 632 20664
rect 666 20630 715 20664
rect 583 20596 715 20630
rect 583 20562 632 20596
rect 666 20562 715 20596
rect 583 20528 715 20562
rect 583 20494 632 20528
rect 666 20494 715 20528
rect 583 20460 715 20494
rect 583 20426 632 20460
rect 666 20426 715 20460
rect 583 20392 715 20426
rect 583 20358 632 20392
rect 666 20358 715 20392
rect 583 20324 715 20358
rect 583 20290 632 20324
rect 666 20290 715 20324
rect 583 20256 715 20290
rect 583 20222 632 20256
rect 666 20222 715 20256
rect 583 20188 715 20222
rect 583 20154 632 20188
rect 666 20154 715 20188
rect 583 20120 715 20154
rect 583 20086 632 20120
rect 666 20086 715 20120
rect 583 20052 715 20086
rect 583 20018 632 20052
rect 666 20018 715 20052
rect 583 19984 715 20018
rect 583 19950 632 19984
rect 666 19950 715 19984
rect 583 19916 715 19950
rect 583 19882 632 19916
rect 666 19882 715 19916
rect 583 19848 715 19882
rect 583 19814 632 19848
rect 666 19814 715 19848
rect 583 19780 715 19814
rect 583 19746 632 19780
rect 666 19746 715 19780
rect 583 19712 715 19746
rect 583 19678 632 19712
rect 666 19678 715 19712
rect 583 19644 715 19678
rect 583 19610 632 19644
rect 666 19610 715 19644
rect 583 19576 715 19610
rect 583 19542 632 19576
rect 666 19542 715 19576
rect 583 19508 715 19542
rect 583 19474 632 19508
rect 666 19474 715 19508
rect 583 19440 715 19474
rect 583 19406 632 19440
rect 666 19406 715 19440
rect 583 19372 715 19406
rect 583 19338 632 19372
rect 666 19338 715 19372
rect 583 19304 715 19338
rect 583 19270 632 19304
rect 666 19270 715 19304
rect 583 19236 715 19270
rect 583 19202 632 19236
rect 666 19202 715 19236
rect 583 19168 715 19202
rect 583 19134 632 19168
rect 666 19134 715 19168
rect 583 19100 715 19134
rect 583 19066 632 19100
rect 666 19066 715 19100
rect 583 19032 715 19066
rect 583 18998 632 19032
rect 666 18998 715 19032
rect 583 18964 715 18998
rect 583 18930 632 18964
rect 666 18930 715 18964
rect 583 18896 715 18930
rect 583 18862 632 18896
rect 666 18862 715 18896
rect 583 18828 715 18862
rect 583 18794 632 18828
rect 666 18794 715 18828
rect 583 18760 715 18794
rect 583 18726 632 18760
rect 666 18726 715 18760
rect 583 18692 715 18726
rect 583 18658 632 18692
rect 666 18658 715 18692
rect 583 18624 715 18658
rect 583 18590 632 18624
rect 666 18590 715 18624
rect 583 18556 715 18590
rect 583 18522 632 18556
rect 666 18522 715 18556
rect 583 18488 715 18522
rect 583 18454 632 18488
rect 666 18454 715 18488
rect 583 18420 715 18454
rect 583 18386 632 18420
rect 666 18386 715 18420
rect 583 18352 715 18386
rect 583 18318 632 18352
rect 666 18318 715 18352
rect 583 18284 715 18318
rect 583 18250 632 18284
rect 666 18250 715 18284
rect 583 18216 715 18250
rect 583 18182 632 18216
rect 666 18182 715 18216
rect 583 18148 715 18182
rect 583 18114 632 18148
rect 666 18114 715 18148
rect 583 18080 715 18114
rect 583 18046 632 18080
rect 666 18046 715 18080
rect 583 18012 715 18046
rect 583 17978 632 18012
rect 666 17978 715 18012
rect 583 17944 715 17978
rect 583 17910 632 17944
rect 666 17910 715 17944
rect 583 17876 715 17910
rect 583 17842 632 17876
rect 666 17842 715 17876
rect 583 17808 715 17842
rect 583 17774 632 17808
rect 666 17774 715 17808
rect 583 17740 715 17774
rect 583 17706 632 17740
rect 666 17706 715 17740
rect 583 17672 715 17706
rect 583 17638 632 17672
rect 666 17638 715 17672
rect 583 17604 715 17638
rect 583 17570 632 17604
rect 666 17570 715 17604
rect 583 17536 715 17570
rect 583 17502 632 17536
rect 666 17502 715 17536
rect 583 17468 715 17502
rect 583 17434 632 17468
rect 666 17434 715 17468
rect 583 17400 715 17434
rect 583 17366 632 17400
rect 666 17366 715 17400
rect 583 17332 715 17366
rect 583 17298 632 17332
rect 666 17298 715 17332
rect 583 17264 715 17298
rect 583 17230 632 17264
rect 666 17230 715 17264
rect 583 17196 715 17230
rect 583 17162 632 17196
rect 666 17162 715 17196
rect 583 17128 715 17162
rect 583 17094 632 17128
rect 666 17094 715 17128
rect 583 17060 715 17094
rect 583 17026 632 17060
rect 666 17026 715 17060
rect 583 16992 715 17026
rect 583 16958 632 16992
rect 666 16958 715 16992
rect 583 16924 715 16958
rect 583 16890 632 16924
rect 666 16890 715 16924
rect 583 16856 715 16890
rect 583 16822 632 16856
rect 666 16822 715 16856
rect 583 16788 715 16822
rect 583 16754 632 16788
rect 666 16754 715 16788
rect 583 16720 715 16754
rect 583 16686 632 16720
rect 666 16686 715 16720
rect 583 16652 715 16686
rect 583 16618 632 16652
rect 666 16618 715 16652
rect 583 16584 715 16618
rect 583 16550 632 16584
rect 666 16550 715 16584
rect 583 16516 715 16550
rect 583 16482 632 16516
rect 666 16482 715 16516
rect 583 16448 715 16482
rect 583 16414 632 16448
rect 666 16414 715 16448
rect 583 16380 715 16414
rect 583 16346 632 16380
rect 666 16346 715 16380
rect 583 16312 715 16346
rect 583 16278 632 16312
rect 666 16278 715 16312
rect 583 16244 715 16278
rect 583 16210 632 16244
rect 666 16210 715 16244
rect 583 16176 715 16210
rect 583 16142 632 16176
rect 666 16142 715 16176
rect 583 16108 715 16142
rect 583 16074 632 16108
rect 666 16074 715 16108
rect 583 16040 715 16074
rect 583 16006 632 16040
rect 666 16006 715 16040
rect 583 15972 715 16006
rect 583 15938 632 15972
rect 666 15938 715 15972
rect 583 15904 715 15938
rect 583 15870 632 15904
rect 666 15870 715 15904
rect 583 15836 715 15870
rect 583 15802 632 15836
rect 666 15802 715 15836
rect 583 15768 715 15802
rect 583 15734 632 15768
rect 666 15734 715 15768
rect 583 15700 715 15734
rect 583 15666 632 15700
rect 666 15666 715 15700
rect 583 15632 715 15666
rect 583 15598 632 15632
rect 666 15598 715 15632
rect 583 15564 715 15598
rect 583 15530 632 15564
rect 666 15530 715 15564
rect 583 15496 715 15530
rect 583 15462 632 15496
rect 666 15462 715 15496
rect 583 15428 715 15462
rect 583 15394 632 15428
rect 666 15394 715 15428
rect 583 15360 715 15394
rect 583 15326 632 15360
rect 666 15326 715 15360
rect 583 15292 715 15326
rect 583 15258 632 15292
rect 666 15258 715 15292
rect 583 15224 715 15258
rect 583 15190 632 15224
rect 666 15190 715 15224
rect 583 15156 715 15190
rect 583 15122 632 15156
rect 666 15122 715 15156
rect 583 15088 715 15122
rect 583 15054 632 15088
rect 666 15054 715 15088
rect 583 15020 715 15054
rect 583 14986 632 15020
rect 666 14986 715 15020
rect 583 14952 715 14986
rect 583 14918 632 14952
rect 666 14918 715 14952
rect 583 14884 715 14918
rect 583 14850 632 14884
rect 666 14850 715 14884
rect 583 14816 715 14850
rect 583 14782 632 14816
rect 666 14782 715 14816
rect 583 14748 715 14782
rect 583 14714 632 14748
rect 666 14714 715 14748
rect 583 14680 715 14714
rect 583 14646 632 14680
rect 666 14646 715 14680
rect 583 14612 715 14646
rect 583 14578 632 14612
rect 666 14578 715 14612
rect 583 14544 715 14578
rect 583 14510 632 14544
rect 666 14510 715 14544
rect 583 14476 715 14510
rect 583 14442 632 14476
rect 666 14442 715 14476
rect 583 14408 715 14442
rect 583 14374 632 14408
rect 666 14374 715 14408
rect 583 14340 715 14374
rect 583 14306 632 14340
rect 666 14306 715 14340
rect 583 14272 715 14306
rect 583 14238 632 14272
rect 666 14238 715 14272
rect 583 14204 715 14238
rect 583 14170 632 14204
rect 666 14170 715 14204
rect 583 14136 715 14170
rect 583 14102 632 14136
rect 666 14102 715 14136
rect 583 14068 715 14102
rect 583 14034 632 14068
rect 666 14034 715 14068
rect 583 14000 715 14034
rect 583 13966 632 14000
rect 666 13966 715 14000
rect 583 13932 715 13966
rect 583 13898 632 13932
rect 666 13898 715 13932
rect 583 13864 715 13898
rect 583 13830 632 13864
rect 666 13830 715 13864
rect 583 13796 715 13830
rect 583 13762 632 13796
rect 666 13762 715 13796
rect 583 13728 715 13762
rect 583 13694 632 13728
rect 666 13694 715 13728
rect 583 13660 715 13694
rect 583 13626 632 13660
rect 666 13626 715 13660
rect 583 13592 715 13626
rect 583 13558 632 13592
rect 666 13558 715 13592
rect 583 13524 715 13558
rect 583 13490 632 13524
rect 666 13490 715 13524
rect 583 13456 715 13490
rect 583 13422 632 13456
rect 666 13422 715 13456
rect 583 13388 715 13422
rect 583 13354 632 13388
rect 666 13354 715 13388
rect 583 13320 715 13354
rect 583 13286 632 13320
rect 666 13286 715 13320
rect 583 13252 715 13286
rect 583 13218 632 13252
rect 666 13218 715 13252
rect 583 13184 715 13218
rect 583 13150 632 13184
rect 666 13150 715 13184
rect 583 13116 715 13150
rect 583 13082 632 13116
rect 666 13082 715 13116
rect 583 13048 715 13082
rect 583 13014 632 13048
rect 666 13014 715 13048
rect 583 12980 715 13014
rect 583 12946 632 12980
rect 666 12946 715 12980
rect 583 12912 715 12946
rect 583 12878 632 12912
rect 666 12878 715 12912
rect 583 12844 715 12878
rect 583 12810 632 12844
rect 666 12810 715 12844
rect 583 12776 715 12810
rect 583 12742 632 12776
rect 666 12742 715 12776
rect 583 12708 715 12742
rect 583 12674 632 12708
rect 666 12674 715 12708
rect 583 12640 715 12674
rect 583 12606 632 12640
rect 666 12606 715 12640
rect 583 12572 715 12606
rect 583 12538 632 12572
rect 666 12538 715 12572
rect 583 12504 715 12538
rect 583 12470 632 12504
rect 666 12470 715 12504
rect 583 12436 715 12470
rect 583 12402 632 12436
rect 666 12402 715 12436
rect 583 12368 715 12402
rect 583 12334 632 12368
rect 666 12334 715 12368
rect 583 12300 715 12334
rect 583 12266 632 12300
rect 666 12266 715 12300
rect 583 12232 715 12266
rect 583 12198 632 12232
rect 666 12198 715 12232
rect 583 12164 715 12198
rect 583 12130 632 12164
rect 666 12130 715 12164
rect 583 12096 715 12130
rect 583 12062 632 12096
rect 666 12062 715 12096
rect 583 12028 715 12062
rect 583 11994 632 12028
rect 666 11994 715 12028
rect 583 11960 715 11994
rect 583 11926 632 11960
rect 666 11926 715 11960
rect 583 11892 715 11926
rect 583 11858 632 11892
rect 666 11858 715 11892
rect 583 11824 715 11858
rect 583 11790 632 11824
rect 666 11790 715 11824
rect 583 11756 715 11790
rect 583 11722 632 11756
rect 666 11722 715 11756
rect 583 11688 715 11722
rect 583 11654 632 11688
rect 666 11654 715 11688
rect 583 11620 715 11654
rect 583 11586 632 11620
rect 666 11586 715 11620
rect 583 11552 715 11586
rect 583 11518 632 11552
rect 666 11518 715 11552
rect 583 11484 715 11518
rect 583 11450 632 11484
rect 666 11450 715 11484
rect 583 11416 715 11450
rect 583 11382 632 11416
rect 666 11382 715 11416
rect 583 11348 715 11382
rect 583 11314 632 11348
rect 666 11314 715 11348
rect 583 11280 715 11314
rect 583 11246 632 11280
rect 666 11246 715 11280
rect 583 11212 715 11246
rect 583 11178 632 11212
rect 666 11178 715 11212
rect 583 11144 715 11178
rect 583 11110 632 11144
rect 666 11110 715 11144
rect 583 11076 715 11110
rect 583 11042 632 11076
rect 666 11042 715 11076
rect 583 11008 715 11042
rect 583 10974 632 11008
rect 666 10974 715 11008
rect 583 10940 715 10974
rect 583 10906 632 10940
rect 666 10906 715 10940
rect 583 10872 715 10906
rect 583 10838 632 10872
rect 666 10838 715 10872
rect 583 10804 715 10838
rect 583 10770 632 10804
rect 666 10770 715 10804
rect 583 10736 715 10770
rect 583 10702 632 10736
rect 666 10702 715 10736
rect 583 10668 715 10702
rect 583 10634 632 10668
rect 666 10634 715 10668
rect 583 10600 715 10634
rect 583 10566 632 10600
rect 666 10566 715 10600
rect 583 10532 715 10566
rect 583 10498 632 10532
rect 666 10498 715 10532
rect 583 10464 715 10498
rect 583 10430 632 10464
rect 666 10430 715 10464
rect 583 10396 715 10430
rect 583 10362 632 10396
rect 666 10362 715 10396
rect 583 10328 715 10362
rect 583 10294 632 10328
rect 666 10294 715 10328
rect 583 10260 715 10294
rect 583 10226 632 10260
rect 666 10226 715 10260
rect 583 10192 715 10226
rect 1659 28879 13357 28909
rect 1659 28505 2119 28879
rect 12897 28505 13357 28879
rect 1659 28475 13357 28505
rect 1659 28422 2093 28475
rect 1659 27504 1689 28422
rect 2063 27504 2093 28422
rect 1659 27451 2093 27504
rect 12923 28422 13357 28475
rect 12923 27504 12953 28422
rect 13327 27504 13357 28422
rect 12923 27451 13357 27504
rect 1659 27421 13357 27451
rect 1659 27047 2119 27421
rect 12897 27047 13357 27421
rect 1659 27017 13357 27047
rect 14247 34706 14297 34740
rect 14331 34706 14381 34740
rect 14247 34672 14381 34706
rect 14247 34638 14297 34672
rect 14331 34638 14381 34672
rect 14247 34604 14381 34638
rect 14247 34570 14297 34604
rect 14331 34570 14381 34604
rect 14247 34536 14381 34570
rect 14247 34502 14297 34536
rect 14331 34502 14381 34536
rect 14247 34468 14381 34502
rect 14247 34434 14297 34468
rect 14331 34434 14381 34468
rect 14247 34400 14381 34434
rect 14247 34366 14297 34400
rect 14331 34366 14381 34400
rect 14247 34332 14381 34366
rect 14247 34298 14297 34332
rect 14331 34298 14381 34332
rect 14247 34264 14381 34298
rect 14247 34230 14297 34264
rect 14331 34230 14381 34264
rect 14247 34196 14381 34230
rect 14247 34162 14297 34196
rect 14331 34162 14381 34196
rect 14247 34128 14381 34162
rect 14247 34094 14297 34128
rect 14331 34094 14381 34128
rect 14247 34060 14381 34094
rect 14247 34026 14297 34060
rect 14331 34026 14381 34060
rect 14247 33992 14381 34026
rect 14247 33958 14297 33992
rect 14331 33958 14381 33992
rect 14247 33924 14381 33958
rect 14247 33890 14297 33924
rect 14331 33890 14381 33924
rect 14247 33856 14381 33890
rect 14247 33822 14297 33856
rect 14331 33822 14381 33856
rect 14247 33788 14381 33822
rect 14247 33754 14297 33788
rect 14331 33754 14381 33788
rect 14247 33720 14381 33754
rect 14247 33686 14297 33720
rect 14331 33686 14381 33720
rect 14247 33652 14381 33686
rect 14247 33618 14297 33652
rect 14331 33618 14381 33652
rect 14247 33584 14381 33618
rect 14247 33550 14297 33584
rect 14331 33550 14381 33584
rect 14247 33516 14381 33550
rect 14247 33482 14297 33516
rect 14331 33482 14381 33516
rect 14247 33448 14381 33482
rect 14247 33414 14297 33448
rect 14331 33414 14381 33448
rect 14247 33380 14381 33414
rect 14247 33346 14297 33380
rect 14331 33346 14381 33380
rect 14247 33312 14381 33346
rect 14247 33278 14297 33312
rect 14331 33278 14381 33312
rect 14247 33244 14381 33278
rect 14247 33210 14297 33244
rect 14331 33210 14381 33244
rect 14247 33176 14381 33210
rect 14247 33142 14297 33176
rect 14331 33142 14381 33176
rect 14247 33108 14381 33142
rect 14247 33074 14297 33108
rect 14331 33074 14381 33108
rect 14247 33040 14381 33074
rect 14247 33006 14297 33040
rect 14331 33006 14381 33040
rect 14247 32972 14381 33006
rect 14247 32938 14297 32972
rect 14331 32938 14381 32972
rect 14247 32904 14381 32938
rect 14247 32870 14297 32904
rect 14331 32870 14381 32904
rect 14247 32836 14381 32870
rect 14247 32802 14297 32836
rect 14331 32802 14381 32836
rect 14247 32768 14381 32802
rect 14247 32734 14297 32768
rect 14331 32734 14381 32768
rect 14247 32700 14381 32734
rect 14247 32666 14297 32700
rect 14331 32666 14381 32700
rect 14247 32632 14381 32666
rect 14247 32598 14297 32632
rect 14331 32598 14381 32632
rect 14247 32564 14381 32598
rect 14247 32530 14297 32564
rect 14331 32530 14381 32564
rect 14247 32496 14381 32530
rect 14247 32462 14297 32496
rect 14331 32462 14381 32496
rect 14247 32428 14381 32462
rect 14247 32394 14297 32428
rect 14331 32394 14381 32428
rect 14247 32360 14381 32394
rect 14247 32326 14297 32360
rect 14331 32326 14381 32360
rect 14247 32292 14381 32326
rect 14247 32258 14297 32292
rect 14331 32258 14381 32292
rect 14247 32224 14381 32258
rect 14247 32190 14297 32224
rect 14331 32190 14381 32224
rect 14247 32156 14381 32190
rect 14247 32122 14297 32156
rect 14331 32122 14381 32156
rect 14247 32088 14381 32122
rect 14247 32054 14297 32088
rect 14331 32054 14381 32088
rect 14247 32020 14381 32054
rect 14247 31986 14297 32020
rect 14331 31986 14381 32020
rect 14247 31952 14381 31986
rect 14247 31918 14297 31952
rect 14331 31918 14381 31952
rect 14247 31884 14381 31918
rect 14247 31850 14297 31884
rect 14331 31850 14381 31884
rect 14247 31816 14381 31850
rect 14247 31782 14297 31816
rect 14331 31782 14381 31816
rect 14247 31748 14381 31782
rect 14247 31714 14297 31748
rect 14331 31714 14381 31748
rect 14247 31680 14381 31714
rect 14247 31646 14297 31680
rect 14331 31646 14381 31680
rect 14247 31612 14381 31646
rect 14247 31578 14297 31612
rect 14331 31578 14381 31612
rect 14247 31544 14381 31578
rect 14247 31510 14297 31544
rect 14331 31510 14381 31544
rect 14247 31476 14381 31510
rect 14247 31442 14297 31476
rect 14331 31442 14381 31476
rect 14247 31408 14381 31442
rect 14247 31374 14297 31408
rect 14331 31374 14381 31408
rect 14247 31340 14381 31374
rect 14247 31306 14297 31340
rect 14331 31306 14381 31340
rect 14247 31272 14381 31306
rect 14247 31238 14297 31272
rect 14331 31238 14381 31272
rect 14247 31204 14381 31238
rect 14247 31170 14297 31204
rect 14331 31170 14381 31204
rect 14247 31136 14381 31170
rect 14247 31102 14297 31136
rect 14331 31102 14381 31136
rect 14247 31068 14381 31102
rect 14247 31034 14297 31068
rect 14331 31034 14381 31068
rect 14247 31000 14381 31034
rect 14247 30966 14297 31000
rect 14331 30966 14381 31000
rect 14247 30932 14381 30966
rect 14247 30898 14297 30932
rect 14331 30898 14381 30932
rect 14247 30864 14381 30898
rect 14247 30830 14297 30864
rect 14331 30830 14381 30864
rect 14247 30796 14381 30830
rect 14247 30762 14297 30796
rect 14331 30762 14381 30796
rect 14247 30728 14381 30762
rect 14247 30694 14297 30728
rect 14331 30694 14381 30728
rect 14247 30660 14381 30694
rect 14247 30626 14297 30660
rect 14331 30626 14381 30660
rect 14247 30592 14381 30626
rect 14247 30558 14297 30592
rect 14331 30558 14381 30592
rect 14247 30524 14381 30558
rect 14247 30490 14297 30524
rect 14331 30490 14381 30524
rect 14247 30456 14381 30490
rect 14247 30422 14297 30456
rect 14331 30422 14381 30456
rect 14247 30388 14381 30422
rect 14247 30354 14297 30388
rect 14331 30354 14381 30388
rect 14247 30320 14381 30354
rect 14247 30286 14297 30320
rect 14331 30286 14381 30320
rect 14247 30252 14381 30286
rect 14247 30218 14297 30252
rect 14331 30218 14381 30252
rect 14247 30184 14381 30218
rect 14247 30150 14297 30184
rect 14331 30150 14381 30184
rect 14247 30116 14381 30150
rect 14247 30082 14297 30116
rect 14331 30082 14381 30116
rect 14247 30048 14381 30082
rect 14247 30014 14297 30048
rect 14331 30014 14381 30048
rect 14247 29980 14381 30014
rect 14247 29946 14297 29980
rect 14331 29946 14381 29980
rect 14247 29912 14381 29946
rect 14247 29878 14297 29912
rect 14331 29878 14381 29912
rect 14247 29844 14381 29878
rect 14247 29810 14297 29844
rect 14331 29810 14381 29844
rect 14247 29776 14381 29810
rect 14247 29742 14297 29776
rect 14331 29742 14381 29776
rect 14247 29708 14381 29742
rect 14247 29674 14297 29708
rect 14331 29674 14381 29708
rect 14247 29640 14381 29674
rect 14247 29606 14297 29640
rect 14331 29606 14381 29640
rect 14247 29572 14381 29606
rect 14247 29538 14297 29572
rect 14331 29538 14381 29572
rect 14247 29504 14381 29538
rect 14247 29470 14297 29504
rect 14331 29470 14381 29504
rect 14247 29436 14381 29470
rect 14247 29402 14297 29436
rect 14331 29402 14381 29436
rect 14247 29368 14381 29402
rect 14247 29334 14297 29368
rect 14331 29334 14381 29368
rect 14247 29300 14381 29334
rect 14247 29266 14297 29300
rect 14331 29266 14381 29300
rect 14247 29232 14381 29266
rect 14247 29198 14297 29232
rect 14331 29198 14381 29232
rect 14247 29164 14381 29198
rect 14247 29130 14297 29164
rect 14331 29130 14381 29164
rect 14247 29096 14381 29130
rect 14247 29062 14297 29096
rect 14331 29062 14381 29096
rect 14247 29028 14381 29062
rect 14247 28994 14297 29028
rect 14331 28994 14381 29028
rect 14247 28960 14381 28994
rect 14247 28926 14297 28960
rect 14331 28926 14381 28960
rect 14247 28892 14381 28926
rect 14247 28858 14297 28892
rect 14331 28858 14381 28892
rect 14247 28824 14381 28858
rect 14247 28790 14297 28824
rect 14331 28790 14381 28824
rect 14247 28756 14381 28790
rect 14247 28722 14297 28756
rect 14331 28722 14381 28756
rect 14247 28688 14381 28722
rect 14247 28654 14297 28688
rect 14331 28654 14381 28688
rect 14247 28620 14381 28654
rect 14247 28586 14297 28620
rect 14331 28586 14381 28620
rect 14247 28552 14381 28586
rect 14247 28518 14297 28552
rect 14331 28518 14381 28552
rect 14247 28484 14381 28518
rect 14247 28450 14297 28484
rect 14331 28450 14381 28484
rect 14247 28416 14381 28450
rect 14247 28382 14297 28416
rect 14331 28382 14381 28416
rect 14247 28348 14381 28382
rect 14247 28314 14297 28348
rect 14331 28314 14381 28348
rect 14247 28280 14381 28314
rect 14247 28246 14297 28280
rect 14331 28246 14381 28280
rect 14247 28212 14381 28246
rect 14247 28178 14297 28212
rect 14331 28178 14381 28212
rect 14247 28144 14381 28178
rect 14247 28110 14297 28144
rect 14331 28110 14381 28144
rect 14247 28076 14381 28110
rect 14247 28042 14297 28076
rect 14331 28042 14381 28076
rect 14247 28008 14381 28042
rect 14247 27974 14297 28008
rect 14331 27974 14381 28008
rect 14247 27940 14381 27974
rect 14247 27906 14297 27940
rect 14331 27906 14381 27940
rect 14247 27872 14381 27906
rect 14247 27838 14297 27872
rect 14331 27838 14381 27872
rect 14247 27804 14381 27838
rect 14247 27770 14297 27804
rect 14331 27770 14381 27804
rect 14247 27736 14381 27770
rect 14247 27702 14297 27736
rect 14331 27702 14381 27736
rect 14247 27668 14381 27702
rect 14247 27634 14297 27668
rect 14331 27634 14381 27668
rect 14247 27600 14381 27634
rect 14247 27566 14297 27600
rect 14331 27566 14381 27600
rect 14247 27532 14381 27566
rect 14247 27498 14297 27532
rect 14331 27498 14381 27532
rect 14247 27464 14381 27498
rect 14247 27430 14297 27464
rect 14331 27430 14381 27464
rect 14247 27396 14381 27430
rect 14247 27362 14297 27396
rect 14331 27362 14381 27396
rect 14247 27328 14381 27362
rect 14247 27294 14297 27328
rect 14331 27294 14381 27328
rect 14247 27260 14381 27294
rect 14247 27226 14297 27260
rect 14331 27226 14381 27260
rect 14247 27192 14381 27226
rect 14247 27158 14297 27192
rect 14331 27158 14381 27192
rect 14247 27124 14381 27158
rect 14247 27090 14297 27124
rect 14331 27090 14381 27124
rect 14247 27056 14381 27090
rect 14247 27022 14297 27056
rect 14331 27022 14381 27056
rect 14247 26988 14381 27022
rect 14247 26954 14297 26988
rect 14331 26954 14381 26988
rect 14247 26920 14381 26954
rect 14247 26886 14297 26920
rect 14331 26886 14381 26920
rect 14247 26852 14381 26886
rect 14247 26818 14297 26852
rect 14331 26818 14381 26852
rect 14247 26784 14381 26818
rect 14247 26750 14297 26784
rect 14331 26750 14381 26784
rect 14247 26716 14381 26750
rect 14247 26682 14297 26716
rect 14331 26682 14381 26716
rect 14247 26648 14381 26682
rect 14247 26614 14297 26648
rect 14331 26614 14381 26648
rect 14247 26580 14381 26614
rect 14247 26546 14297 26580
rect 14331 26546 14381 26580
rect 14247 26512 14381 26546
rect 14247 26478 14297 26512
rect 14331 26478 14381 26512
rect 14247 26444 14381 26478
rect 14247 26410 14297 26444
rect 14331 26410 14381 26444
rect 14247 26376 14381 26410
rect 14247 26342 14297 26376
rect 14331 26342 14381 26376
rect 14247 26308 14381 26342
rect 14247 26274 14297 26308
rect 14331 26274 14381 26308
rect 14247 26240 14381 26274
rect 14247 26206 14297 26240
rect 14331 26206 14381 26240
rect 14247 26172 14381 26206
rect 14247 26138 14297 26172
rect 14331 26138 14381 26172
rect 14247 26104 14381 26138
rect 14247 26070 14297 26104
rect 14331 26070 14381 26104
rect 14247 26036 14381 26070
rect 14247 26002 14297 26036
rect 14331 26002 14381 26036
rect 14247 25968 14381 26002
rect 14247 25934 14297 25968
rect 14331 25934 14381 25968
rect 14247 25900 14381 25934
rect 14247 25866 14297 25900
rect 14331 25866 14381 25900
rect 14247 25832 14381 25866
rect 14247 25798 14297 25832
rect 14331 25798 14381 25832
rect 14247 25764 14381 25798
rect 14247 25730 14297 25764
rect 14331 25730 14381 25764
rect 14247 25696 14381 25730
rect 14247 25662 14297 25696
rect 14331 25662 14381 25696
rect 14247 25628 14381 25662
rect 14247 25594 14297 25628
rect 14331 25594 14381 25628
rect 14247 25560 14381 25594
rect 14247 25526 14297 25560
rect 14331 25526 14381 25560
rect 14247 25492 14381 25526
rect 14247 25458 14297 25492
rect 14331 25458 14381 25492
rect 14247 25424 14381 25458
rect 14247 25390 14297 25424
rect 14331 25390 14381 25424
rect 14247 25356 14381 25390
rect 14247 25322 14297 25356
rect 14331 25322 14381 25356
rect 14247 25288 14381 25322
rect 14247 25254 14297 25288
rect 14331 25254 14381 25288
rect 14247 25220 14381 25254
rect 14247 25186 14297 25220
rect 14331 25186 14381 25220
rect 14247 25152 14381 25186
rect 14247 25118 14297 25152
rect 14331 25118 14381 25152
rect 14247 25084 14381 25118
rect 14247 25050 14297 25084
rect 14331 25050 14381 25084
rect 14247 25016 14381 25050
rect 14247 24982 14297 25016
rect 14331 24982 14381 25016
rect 14247 24948 14381 24982
rect 14247 24914 14297 24948
rect 14331 24914 14381 24948
rect 14247 24880 14381 24914
rect 14247 24846 14297 24880
rect 14331 24846 14381 24880
rect 14247 24812 14381 24846
rect 14247 24778 14297 24812
rect 14331 24778 14381 24812
rect 14247 24744 14381 24778
rect 14247 24710 14297 24744
rect 14331 24710 14381 24744
rect 14247 24676 14381 24710
rect 14247 24642 14297 24676
rect 14331 24642 14381 24676
rect 14247 24608 14381 24642
rect 14247 24574 14297 24608
rect 14331 24574 14381 24608
rect 14247 24540 14381 24574
rect 14247 24506 14297 24540
rect 14331 24506 14381 24540
rect 14247 24472 14381 24506
rect 14247 24438 14297 24472
rect 14331 24438 14381 24472
rect 14247 24404 14381 24438
rect 14247 24370 14297 24404
rect 14331 24370 14381 24404
rect 14247 24336 14381 24370
rect 14247 24302 14297 24336
rect 14331 24302 14381 24336
rect 14247 24268 14381 24302
rect 14247 24234 14297 24268
rect 14331 24234 14381 24268
rect 14247 24200 14381 24234
rect 14247 24166 14297 24200
rect 14331 24166 14381 24200
rect 14247 24132 14381 24166
rect 14247 24098 14297 24132
rect 14331 24098 14381 24132
rect 14247 24064 14381 24098
rect 14247 24030 14297 24064
rect 14331 24030 14381 24064
rect 14247 23996 14381 24030
rect 14247 23962 14297 23996
rect 14331 23962 14381 23996
rect 14247 23928 14381 23962
rect 14247 23894 14297 23928
rect 14331 23894 14381 23928
rect 14247 23860 14381 23894
rect 14247 23826 14297 23860
rect 14331 23826 14381 23860
rect 14247 23792 14381 23826
rect 14247 23758 14297 23792
rect 14331 23758 14381 23792
rect 14247 23724 14381 23758
rect 14247 23690 14297 23724
rect 14331 23690 14381 23724
rect 14247 23656 14381 23690
rect 14247 23622 14297 23656
rect 14331 23622 14381 23656
rect 14247 23588 14381 23622
rect 14247 23554 14297 23588
rect 14331 23554 14381 23588
rect 14247 23520 14381 23554
rect 14247 23486 14297 23520
rect 14331 23486 14381 23520
rect 14247 23452 14381 23486
rect 14247 23418 14297 23452
rect 14331 23418 14381 23452
rect 14247 23384 14381 23418
rect 14247 23350 14297 23384
rect 14331 23350 14381 23384
rect 14247 23316 14381 23350
rect 14247 23282 14297 23316
rect 14331 23282 14381 23316
rect 14247 23248 14381 23282
rect 14247 23214 14297 23248
rect 14331 23214 14381 23248
rect 14247 23180 14381 23214
rect 14247 23146 14297 23180
rect 14331 23146 14381 23180
rect 14247 23112 14381 23146
rect 14247 23078 14297 23112
rect 14331 23078 14381 23112
rect 14247 23044 14381 23078
rect 14247 23010 14297 23044
rect 14331 23010 14381 23044
rect 14247 22976 14381 23010
rect 14247 22942 14297 22976
rect 14331 22942 14381 22976
rect 14247 22908 14381 22942
rect 14247 22874 14297 22908
rect 14331 22874 14381 22908
rect 14247 22840 14381 22874
rect 14247 22806 14297 22840
rect 14331 22806 14381 22840
rect 14247 22772 14381 22806
rect 14247 22738 14297 22772
rect 14331 22738 14381 22772
rect 14247 22704 14381 22738
rect 14247 22670 14297 22704
rect 14331 22670 14381 22704
rect 14247 22636 14381 22670
rect 14247 22602 14297 22636
rect 14331 22602 14381 22636
rect 14247 22568 14381 22602
rect 14247 22534 14297 22568
rect 14331 22534 14381 22568
rect 14247 22500 14381 22534
rect 14247 22466 14297 22500
rect 14331 22466 14381 22500
rect 14247 22432 14381 22466
rect 14247 22398 14297 22432
rect 14331 22398 14381 22432
rect 14247 22364 14381 22398
rect 14247 22330 14297 22364
rect 14331 22330 14381 22364
rect 14247 22296 14381 22330
rect 14247 22262 14297 22296
rect 14331 22262 14381 22296
rect 14247 22228 14381 22262
rect 14247 22194 14297 22228
rect 14331 22194 14381 22228
rect 14247 22160 14381 22194
rect 14247 22126 14297 22160
rect 14331 22126 14381 22160
rect 14247 22092 14381 22126
rect 14247 22058 14297 22092
rect 14331 22058 14381 22092
rect 14247 22024 14381 22058
rect 14247 21990 14297 22024
rect 14331 21990 14381 22024
rect 14247 21956 14381 21990
rect 14247 21922 14297 21956
rect 14331 21922 14381 21956
rect 14247 21888 14381 21922
rect 14247 21854 14297 21888
rect 14331 21854 14381 21888
rect 14247 21820 14381 21854
rect 14247 21786 14297 21820
rect 14331 21786 14381 21820
rect 14247 21752 14381 21786
rect 14247 21718 14297 21752
rect 14331 21718 14381 21752
rect 14247 21684 14381 21718
rect 14247 21650 14297 21684
rect 14331 21650 14381 21684
rect 14247 21616 14381 21650
rect 14247 21582 14297 21616
rect 14331 21582 14381 21616
rect 14247 21548 14381 21582
rect 14247 21514 14297 21548
rect 14331 21514 14381 21548
rect 14247 21480 14381 21514
rect 14247 21446 14297 21480
rect 14331 21446 14381 21480
rect 14247 21412 14381 21446
rect 14247 21378 14297 21412
rect 14331 21378 14381 21412
rect 14247 21344 14381 21378
rect 14247 21310 14297 21344
rect 14331 21310 14381 21344
rect 14247 21276 14381 21310
rect 14247 21242 14297 21276
rect 14331 21242 14381 21276
rect 14247 21208 14381 21242
rect 14247 21174 14297 21208
rect 14331 21174 14381 21208
rect 14247 21140 14381 21174
rect 14247 21106 14297 21140
rect 14331 21106 14381 21140
rect 14247 21072 14381 21106
rect 14247 21038 14297 21072
rect 14331 21038 14381 21072
rect 14247 21004 14381 21038
rect 14247 20970 14297 21004
rect 14331 20970 14381 21004
rect 14247 20936 14381 20970
rect 14247 20902 14297 20936
rect 14331 20902 14381 20936
rect 14247 20868 14381 20902
rect 14247 20834 14297 20868
rect 14331 20834 14381 20868
rect 14247 20800 14381 20834
rect 14247 20766 14297 20800
rect 14331 20766 14381 20800
rect 14247 20732 14381 20766
rect 14247 20698 14297 20732
rect 14331 20698 14381 20732
rect 14247 20664 14381 20698
rect 14247 20630 14297 20664
rect 14331 20630 14381 20664
rect 14247 20596 14381 20630
rect 14247 20562 14297 20596
rect 14331 20562 14381 20596
rect 14247 20528 14381 20562
rect 14247 20494 14297 20528
rect 14331 20494 14381 20528
rect 14247 20460 14381 20494
rect 14247 20426 14297 20460
rect 14331 20426 14381 20460
rect 14247 20392 14381 20426
rect 14247 20358 14297 20392
rect 14331 20358 14381 20392
rect 14247 20324 14381 20358
rect 14247 20290 14297 20324
rect 14331 20290 14381 20324
rect 14247 20256 14381 20290
rect 14247 20222 14297 20256
rect 14331 20222 14381 20256
rect 14247 20188 14381 20222
rect 14247 20154 14297 20188
rect 14331 20154 14381 20188
rect 14247 20120 14381 20154
rect 14247 20086 14297 20120
rect 14331 20086 14381 20120
rect 14247 20052 14381 20086
rect 14247 20018 14297 20052
rect 14331 20018 14381 20052
rect 14247 19984 14381 20018
rect 14247 19950 14297 19984
rect 14331 19950 14381 19984
rect 14247 19916 14381 19950
rect 14247 19882 14297 19916
rect 14331 19882 14381 19916
rect 14247 19848 14381 19882
rect 14247 19814 14297 19848
rect 14331 19814 14381 19848
rect 14247 19780 14381 19814
rect 14247 19746 14297 19780
rect 14331 19746 14381 19780
rect 14247 19712 14381 19746
rect 14247 19678 14297 19712
rect 14331 19678 14381 19712
rect 14247 19644 14381 19678
rect 14247 19610 14297 19644
rect 14331 19610 14381 19644
rect 14247 19576 14381 19610
rect 14247 19542 14297 19576
rect 14331 19542 14381 19576
rect 14247 19508 14381 19542
rect 14247 19474 14297 19508
rect 14331 19474 14381 19508
rect 14247 19440 14381 19474
rect 14247 19406 14297 19440
rect 14331 19406 14381 19440
rect 14247 19372 14381 19406
rect 14247 19338 14297 19372
rect 14331 19338 14381 19372
rect 14247 19304 14381 19338
rect 14247 19270 14297 19304
rect 14331 19270 14381 19304
rect 14247 19236 14381 19270
rect 14247 19202 14297 19236
rect 14331 19202 14381 19236
rect 14247 19168 14381 19202
rect 14247 19134 14297 19168
rect 14331 19134 14381 19168
rect 14247 19100 14381 19134
rect 14247 19066 14297 19100
rect 14331 19066 14381 19100
rect 14247 19032 14381 19066
rect 14247 18998 14297 19032
rect 14331 18998 14381 19032
rect 14247 18964 14381 18998
rect 14247 18930 14297 18964
rect 14331 18930 14381 18964
rect 14247 18896 14381 18930
rect 14247 18862 14297 18896
rect 14331 18862 14381 18896
rect 14247 18828 14381 18862
rect 14247 18794 14297 18828
rect 14331 18794 14381 18828
rect 14247 18760 14381 18794
rect 14247 18726 14297 18760
rect 14331 18726 14381 18760
rect 14247 18692 14381 18726
rect 14247 18658 14297 18692
rect 14331 18658 14381 18692
rect 14247 18624 14381 18658
rect 14247 18590 14297 18624
rect 14331 18590 14381 18624
rect 14247 18556 14381 18590
rect 14247 18522 14297 18556
rect 14331 18522 14381 18556
rect 14247 18488 14381 18522
rect 14247 18454 14297 18488
rect 14331 18454 14381 18488
rect 14247 18420 14381 18454
rect 14247 18386 14297 18420
rect 14331 18386 14381 18420
rect 14247 18352 14381 18386
rect 14247 18318 14297 18352
rect 14331 18318 14381 18352
rect 14247 18284 14381 18318
rect 14247 18250 14297 18284
rect 14331 18250 14381 18284
rect 14247 18216 14381 18250
rect 14247 18182 14297 18216
rect 14331 18182 14381 18216
rect 14247 18148 14381 18182
rect 14247 18114 14297 18148
rect 14331 18114 14381 18148
rect 14247 18080 14381 18114
rect 14247 18046 14297 18080
rect 14331 18046 14381 18080
rect 14247 18012 14381 18046
rect 14247 17978 14297 18012
rect 14331 17978 14381 18012
rect 14247 17944 14381 17978
rect 14247 17910 14297 17944
rect 14331 17910 14381 17944
rect 14247 17876 14381 17910
rect 14247 17842 14297 17876
rect 14331 17842 14381 17876
rect 14247 17808 14381 17842
rect 14247 17774 14297 17808
rect 14331 17774 14381 17808
rect 14247 17740 14381 17774
rect 14247 17706 14297 17740
rect 14331 17706 14381 17740
rect 14247 17672 14381 17706
rect 14247 17638 14297 17672
rect 14331 17638 14381 17672
rect 14247 17604 14381 17638
rect 14247 17570 14297 17604
rect 14331 17570 14381 17604
rect 14247 17536 14381 17570
rect 14247 17502 14297 17536
rect 14331 17502 14381 17536
rect 14247 17468 14381 17502
rect 14247 17434 14297 17468
rect 14331 17434 14381 17468
rect 14247 17400 14381 17434
rect 14247 17366 14297 17400
rect 14331 17366 14381 17400
rect 14247 17332 14381 17366
rect 14247 17298 14297 17332
rect 14331 17298 14381 17332
rect 14247 17264 14381 17298
rect 14247 17230 14297 17264
rect 14331 17230 14381 17264
rect 14247 17196 14381 17230
rect 14247 17162 14297 17196
rect 14331 17162 14381 17196
rect 14247 17128 14381 17162
rect 14247 17094 14297 17128
rect 14331 17094 14381 17128
rect 14247 17060 14381 17094
rect 14247 17026 14297 17060
rect 14331 17026 14381 17060
rect 14247 16992 14381 17026
rect 14247 16958 14297 16992
rect 14331 16958 14381 16992
rect 14247 16924 14381 16958
rect 14247 16890 14297 16924
rect 14331 16890 14381 16924
rect 14247 16856 14381 16890
rect 14247 16822 14297 16856
rect 14331 16822 14381 16856
rect 14247 16788 14381 16822
rect 14247 16754 14297 16788
rect 14331 16754 14381 16788
rect 14247 16720 14381 16754
rect 14247 16686 14297 16720
rect 14331 16686 14381 16720
rect 14247 16652 14381 16686
rect 14247 16618 14297 16652
rect 14331 16618 14381 16652
rect 14247 16584 14381 16618
rect 14247 16550 14297 16584
rect 14331 16550 14381 16584
rect 14247 16516 14381 16550
rect 14247 16482 14297 16516
rect 14331 16482 14381 16516
rect 14247 16448 14381 16482
rect 14247 16414 14297 16448
rect 14331 16414 14381 16448
rect 14247 16380 14381 16414
rect 14247 16346 14297 16380
rect 14331 16346 14381 16380
rect 14247 16312 14381 16346
rect 14247 16278 14297 16312
rect 14331 16278 14381 16312
rect 14247 16244 14381 16278
rect 14247 16210 14297 16244
rect 14331 16210 14381 16244
rect 14247 16176 14381 16210
rect 14247 16142 14297 16176
rect 14331 16142 14381 16176
rect 14247 16108 14381 16142
rect 14247 16074 14297 16108
rect 14331 16074 14381 16108
rect 14247 16040 14381 16074
rect 14247 16006 14297 16040
rect 14331 16006 14381 16040
rect 14247 15972 14381 16006
rect 14247 15938 14297 15972
rect 14331 15938 14381 15972
rect 14247 15904 14381 15938
rect 14247 15870 14297 15904
rect 14331 15870 14381 15904
rect 14247 15836 14381 15870
rect 14247 15802 14297 15836
rect 14331 15802 14381 15836
rect 14247 15768 14381 15802
rect 14247 15734 14297 15768
rect 14331 15734 14381 15768
rect 14247 15700 14381 15734
rect 14247 15666 14297 15700
rect 14331 15666 14381 15700
rect 14247 15632 14381 15666
rect 14247 15598 14297 15632
rect 14331 15598 14381 15632
rect 14247 15564 14381 15598
rect 14247 15530 14297 15564
rect 14331 15530 14381 15564
rect 14247 15496 14381 15530
rect 14247 15462 14297 15496
rect 14331 15462 14381 15496
rect 14247 15428 14381 15462
rect 14247 15394 14297 15428
rect 14331 15394 14381 15428
rect 14247 15360 14381 15394
rect 14247 15326 14297 15360
rect 14331 15326 14381 15360
rect 14247 15292 14381 15326
rect 14247 15258 14297 15292
rect 14331 15258 14381 15292
rect 14247 15224 14381 15258
rect 14247 15190 14297 15224
rect 14331 15190 14381 15224
rect 14247 15156 14381 15190
rect 14247 15122 14297 15156
rect 14331 15122 14381 15156
rect 14247 15088 14381 15122
rect 14247 15054 14297 15088
rect 14331 15054 14381 15088
rect 14247 15020 14381 15054
rect 14247 14986 14297 15020
rect 14331 14986 14381 15020
rect 14247 14952 14381 14986
rect 14247 14918 14297 14952
rect 14331 14918 14381 14952
rect 14247 14884 14381 14918
rect 14247 14850 14297 14884
rect 14331 14850 14381 14884
rect 14247 14816 14381 14850
rect 14247 14782 14297 14816
rect 14331 14782 14381 14816
rect 14247 14748 14381 14782
rect 14247 14714 14297 14748
rect 14331 14714 14381 14748
rect 14247 14680 14381 14714
rect 14247 14646 14297 14680
rect 14331 14646 14381 14680
rect 14247 14612 14381 14646
rect 14247 14578 14297 14612
rect 14331 14578 14381 14612
rect 14247 14544 14381 14578
rect 14247 14510 14297 14544
rect 14331 14510 14381 14544
rect 14247 14476 14381 14510
rect 14247 14442 14297 14476
rect 14331 14442 14381 14476
rect 14247 14408 14381 14442
rect 14247 14374 14297 14408
rect 14331 14374 14381 14408
rect 14247 14340 14381 14374
rect 14247 14306 14297 14340
rect 14331 14306 14381 14340
rect 14247 14272 14381 14306
rect 14247 14238 14297 14272
rect 14331 14238 14381 14272
rect 14247 14204 14381 14238
rect 14247 14170 14297 14204
rect 14331 14170 14381 14204
rect 14247 14136 14381 14170
rect 14247 14102 14297 14136
rect 14331 14102 14381 14136
rect 14247 14068 14381 14102
rect 14247 14034 14297 14068
rect 14331 14034 14381 14068
rect 14247 14000 14381 14034
rect 14247 13966 14297 14000
rect 14331 13966 14381 14000
rect 14247 13932 14381 13966
rect 14247 13898 14297 13932
rect 14331 13898 14381 13932
rect 14247 13864 14381 13898
rect 14247 13830 14297 13864
rect 14331 13830 14381 13864
rect 14247 13796 14381 13830
rect 14247 13762 14297 13796
rect 14331 13762 14381 13796
rect 14247 13728 14381 13762
rect 14247 13694 14297 13728
rect 14331 13694 14381 13728
rect 14247 13660 14381 13694
rect 14247 13626 14297 13660
rect 14331 13626 14381 13660
rect 14247 13592 14381 13626
rect 14247 13558 14297 13592
rect 14331 13558 14381 13592
rect 14247 13524 14381 13558
rect 14247 13490 14297 13524
rect 14331 13490 14381 13524
rect 14247 13456 14381 13490
rect 14247 13422 14297 13456
rect 14331 13422 14381 13456
rect 14247 13388 14381 13422
rect 14247 13354 14297 13388
rect 14331 13354 14381 13388
rect 14247 13320 14381 13354
rect 14247 13286 14297 13320
rect 14331 13286 14381 13320
rect 14247 13252 14381 13286
rect 14247 13218 14297 13252
rect 14331 13218 14381 13252
rect 14247 13184 14381 13218
rect 14247 13150 14297 13184
rect 14331 13150 14381 13184
rect 14247 13116 14381 13150
rect 14247 13082 14297 13116
rect 14331 13082 14381 13116
rect 14247 13048 14381 13082
rect 14247 13014 14297 13048
rect 14331 13014 14381 13048
rect 14247 12980 14381 13014
rect 14247 12946 14297 12980
rect 14331 12946 14381 12980
rect 14247 12912 14381 12946
rect 14247 12878 14297 12912
rect 14331 12878 14381 12912
rect 14247 12844 14381 12878
rect 14247 12810 14297 12844
rect 14331 12810 14381 12844
rect 14247 12776 14381 12810
rect 14247 12742 14297 12776
rect 14331 12742 14381 12776
rect 14247 12708 14381 12742
rect 14247 12674 14297 12708
rect 14331 12674 14381 12708
rect 14247 12640 14381 12674
rect 14247 12606 14297 12640
rect 14331 12606 14381 12640
rect 14247 12572 14381 12606
rect 14247 12538 14297 12572
rect 14331 12538 14381 12572
rect 14247 12504 14381 12538
rect 14247 12470 14297 12504
rect 14331 12470 14381 12504
rect 14247 12436 14381 12470
rect 14247 12402 14297 12436
rect 14331 12402 14381 12436
rect 14247 12368 14381 12402
rect 14247 12334 14297 12368
rect 14331 12334 14381 12368
rect 14247 12300 14381 12334
rect 14247 12266 14297 12300
rect 14331 12266 14381 12300
rect 14247 12232 14381 12266
rect 14247 12198 14297 12232
rect 14331 12198 14381 12232
rect 14247 12164 14381 12198
rect 14247 12130 14297 12164
rect 14331 12130 14381 12164
rect 14247 12096 14381 12130
rect 14247 12062 14297 12096
rect 14331 12062 14381 12096
rect 14247 12028 14381 12062
rect 14247 11994 14297 12028
rect 14331 11994 14381 12028
rect 14247 11960 14381 11994
rect 14247 11926 14297 11960
rect 14331 11926 14381 11960
rect 14247 11892 14381 11926
rect 14247 11858 14297 11892
rect 14331 11858 14381 11892
rect 14247 11824 14381 11858
rect 14247 11790 14297 11824
rect 14331 11790 14381 11824
rect 14247 11756 14381 11790
rect 14247 11722 14297 11756
rect 14331 11722 14381 11756
rect 14247 11688 14381 11722
rect 14247 11654 14297 11688
rect 14331 11654 14381 11688
rect 14247 11620 14381 11654
rect 14247 11586 14297 11620
rect 14331 11586 14381 11620
rect 14247 11552 14381 11586
rect 14247 11518 14297 11552
rect 14331 11518 14381 11552
rect 14247 11484 14381 11518
rect 14247 11450 14297 11484
rect 14331 11450 14381 11484
rect 14247 11416 14381 11450
rect 14247 11382 14297 11416
rect 14331 11382 14381 11416
rect 14247 11348 14381 11382
rect 14247 11314 14297 11348
rect 14331 11314 14381 11348
rect 14247 11280 14381 11314
rect 14247 11246 14297 11280
rect 14331 11246 14381 11280
rect 14247 11212 14381 11246
rect 14247 11178 14297 11212
rect 14331 11178 14381 11212
rect 14247 11144 14381 11178
rect 14247 11110 14297 11144
rect 14331 11110 14381 11144
rect 14247 11076 14381 11110
rect 14247 11042 14297 11076
rect 14331 11042 14381 11076
rect 14247 11008 14381 11042
rect 14247 10974 14297 11008
rect 14331 10974 14381 11008
rect 14247 10940 14381 10974
rect 14247 10906 14297 10940
rect 14331 10906 14381 10940
rect 14247 10872 14381 10906
rect 14247 10838 14297 10872
rect 14331 10838 14381 10872
rect 14247 10804 14381 10838
rect 14247 10770 14297 10804
rect 14331 10770 14381 10804
rect 14247 10736 14381 10770
rect 14247 10702 14297 10736
rect 14331 10702 14381 10736
rect 14247 10668 14381 10702
rect 14247 10634 14297 10668
rect 14331 10634 14381 10668
rect 14247 10600 14381 10634
rect 14247 10566 14297 10600
rect 14331 10566 14381 10600
rect 14247 10532 14381 10566
rect 14247 10498 14297 10532
rect 14331 10498 14381 10532
rect 14247 10464 14381 10498
rect 14247 10430 14297 10464
rect 14331 10430 14381 10464
rect 14247 10396 14381 10430
rect 14247 10362 14297 10396
rect 14331 10362 14381 10396
rect 14247 10328 14381 10362
rect 14247 10294 14297 10328
rect 14331 10294 14381 10328
rect 14247 10260 14381 10294
rect 14247 10226 14297 10260
rect 14331 10226 14381 10260
rect 583 10158 632 10192
rect 666 10158 715 10192
rect 583 10124 715 10158
rect 583 10090 632 10124
rect 666 10090 715 10124
rect 583 10056 715 10090
rect 583 10022 632 10056
rect 666 10022 715 10056
rect 583 9988 715 10022
rect 583 9954 632 9988
rect 666 9954 715 9988
rect 583 9920 715 9954
rect 583 9886 632 9920
rect 666 9886 715 9920
rect 583 9825 715 9886
rect 14247 10192 14381 10226
rect 14247 10158 14297 10192
rect 14331 10158 14381 10192
rect 14247 10124 14381 10158
rect 14247 10090 14297 10124
rect 14331 10090 14381 10124
rect 14247 10056 14381 10090
rect 14247 10022 14297 10056
rect 14331 10022 14381 10056
rect 14247 9988 14381 10022
rect 14247 9954 14297 9988
rect 14331 9954 14381 9988
rect 14247 9920 14381 9954
rect 14247 9886 14297 9920
rect 14331 9886 14381 9920
rect 14247 9825 14381 9886
rect 583 9775 14381 9825
rect 583 9741 766 9775
rect 800 9741 834 9775
rect 868 9741 902 9775
rect 936 9741 970 9775
rect 1004 9741 1038 9775
rect 1072 9741 1106 9775
rect 1140 9741 1174 9775
rect 1208 9741 1242 9775
rect 1276 9741 1310 9775
rect 1344 9741 1378 9775
rect 1412 9741 1446 9775
rect 1480 9741 1514 9775
rect 1548 9741 1582 9775
rect 1616 9741 1650 9775
rect 1684 9741 1718 9775
rect 1752 9741 1786 9775
rect 1820 9741 1854 9775
rect 1888 9741 1922 9775
rect 1956 9741 1990 9775
rect 2024 9741 2058 9775
rect 2092 9741 2126 9775
rect 2160 9741 2194 9775
rect 2228 9741 2262 9775
rect 2296 9741 2330 9775
rect 2364 9741 2398 9775
rect 2432 9741 2466 9775
rect 2500 9741 2534 9775
rect 2568 9741 2602 9775
rect 2636 9741 2670 9775
rect 2704 9741 2738 9775
rect 2772 9741 2806 9775
rect 2840 9741 2874 9775
rect 2908 9741 2942 9775
rect 2976 9741 3010 9775
rect 3044 9741 3078 9775
rect 3112 9741 3146 9775
rect 3180 9741 3214 9775
rect 3248 9741 3282 9775
rect 3316 9741 3350 9775
rect 3384 9741 3418 9775
rect 3452 9741 3486 9775
rect 3520 9741 3554 9775
rect 3588 9741 3622 9775
rect 3656 9741 3690 9775
rect 3724 9741 3758 9775
rect 3792 9741 3826 9775
rect 3860 9741 3894 9775
rect 3928 9741 3962 9775
rect 3996 9741 4030 9775
rect 4064 9741 4098 9775
rect 4132 9741 4166 9775
rect 4200 9741 4234 9775
rect 4268 9741 4302 9775
rect 4336 9741 4370 9775
rect 4404 9741 4438 9775
rect 4472 9741 4506 9775
rect 4540 9741 4574 9775
rect 4608 9741 4642 9775
rect 4676 9741 4710 9775
rect 4744 9741 4778 9775
rect 4812 9741 4846 9775
rect 4880 9741 4914 9775
rect 4948 9741 4982 9775
rect 5016 9741 5050 9775
rect 5084 9741 5118 9775
rect 5152 9741 5186 9775
rect 5220 9741 5254 9775
rect 5288 9741 5322 9775
rect 5356 9741 5390 9775
rect 5424 9741 5458 9775
rect 5492 9741 5526 9775
rect 5560 9741 5594 9775
rect 5628 9741 5662 9775
rect 5696 9741 5730 9775
rect 5764 9741 5798 9775
rect 5832 9741 5866 9775
rect 5900 9741 5934 9775
rect 5968 9741 6002 9775
rect 6036 9741 6070 9775
rect 6104 9741 6138 9775
rect 6172 9741 6206 9775
rect 6240 9741 6274 9775
rect 6308 9741 6342 9775
rect 6376 9741 6410 9775
rect 6444 9741 6478 9775
rect 6512 9741 6546 9775
rect 6580 9741 6614 9775
rect 6648 9741 6682 9775
rect 6716 9741 6750 9775
rect 6784 9741 6818 9775
rect 6852 9741 6886 9775
rect 6920 9741 6954 9775
rect 6988 9741 7022 9775
rect 7056 9741 7090 9775
rect 7124 9741 7158 9775
rect 7192 9741 7226 9775
rect 7260 9741 7294 9775
rect 7328 9741 7362 9775
rect 7396 9741 7430 9775
rect 7464 9741 7498 9775
rect 7532 9741 7566 9775
rect 7600 9741 7634 9775
rect 7668 9741 7702 9775
rect 7736 9741 7770 9775
rect 7804 9741 7838 9775
rect 7872 9741 7906 9775
rect 7940 9741 7974 9775
rect 8008 9741 8042 9775
rect 8076 9741 8110 9775
rect 8144 9741 8178 9775
rect 8212 9741 8246 9775
rect 8280 9741 8314 9775
rect 8348 9741 8382 9775
rect 8416 9741 8450 9775
rect 8484 9741 8518 9775
rect 8552 9741 8586 9775
rect 8620 9741 8654 9775
rect 8688 9741 8722 9775
rect 8756 9741 8790 9775
rect 8824 9741 8858 9775
rect 8892 9741 8926 9775
rect 8960 9741 8994 9775
rect 9028 9741 9062 9775
rect 9096 9741 9130 9775
rect 9164 9741 9198 9775
rect 9232 9741 9266 9775
rect 9300 9741 9334 9775
rect 9368 9741 9402 9775
rect 9436 9741 9470 9775
rect 9504 9741 9538 9775
rect 9572 9741 9606 9775
rect 9640 9741 9674 9775
rect 9708 9741 9742 9775
rect 9776 9741 9810 9775
rect 9844 9741 9878 9775
rect 9912 9741 9946 9775
rect 9980 9741 10014 9775
rect 10048 9741 10082 9775
rect 10116 9741 10150 9775
rect 10184 9741 10218 9775
rect 10252 9741 10286 9775
rect 10320 9741 10354 9775
rect 10388 9741 10422 9775
rect 10456 9741 10490 9775
rect 10524 9741 10558 9775
rect 10592 9741 10626 9775
rect 10660 9741 10694 9775
rect 10728 9741 10762 9775
rect 10796 9741 10830 9775
rect 10864 9741 10898 9775
rect 10932 9741 10966 9775
rect 11000 9741 11034 9775
rect 11068 9741 11102 9775
rect 11136 9741 11170 9775
rect 11204 9741 11238 9775
rect 11272 9741 11306 9775
rect 11340 9741 11374 9775
rect 11408 9741 11442 9775
rect 11476 9741 11510 9775
rect 11544 9741 11578 9775
rect 11612 9741 11646 9775
rect 11680 9741 11714 9775
rect 11748 9741 11782 9775
rect 11816 9741 11850 9775
rect 11884 9741 11918 9775
rect 11952 9741 11986 9775
rect 12020 9741 12054 9775
rect 12088 9741 12122 9775
rect 12156 9741 12190 9775
rect 12224 9741 12258 9775
rect 12292 9741 12326 9775
rect 12360 9741 12394 9775
rect 12428 9741 12462 9775
rect 12496 9741 12530 9775
rect 12564 9741 12598 9775
rect 12632 9741 12666 9775
rect 12700 9741 12734 9775
rect 12768 9741 12802 9775
rect 12836 9741 12870 9775
rect 12904 9741 12938 9775
rect 12972 9741 13006 9775
rect 13040 9741 13074 9775
rect 13108 9741 13142 9775
rect 13176 9741 13210 9775
rect 13244 9741 13278 9775
rect 13312 9741 13346 9775
rect 13380 9741 13414 9775
rect 13448 9741 13482 9775
rect 13516 9741 13550 9775
rect 13584 9741 13618 9775
rect 13652 9741 13686 9775
rect 13720 9741 13754 9775
rect 13788 9741 13822 9775
rect 13856 9741 13890 9775
rect 13924 9741 13958 9775
rect 13992 9741 14026 9775
rect 14060 9741 14094 9775
rect 14128 9741 14162 9775
rect 14196 9741 14381 9775
rect 583 9691 14381 9741
<< mvpsubdiffcont >>
rect 455 36463 489 36497
rect 523 36463 557 36497
rect 591 36463 625 36497
rect 659 36463 693 36497
rect 727 36463 761 36497
rect 795 36463 829 36497
rect 863 36463 897 36497
rect 931 36463 965 36497
rect 999 36463 1033 36497
rect 1067 36463 1101 36497
rect 1135 36463 1169 36497
rect 1203 36463 1237 36497
rect 1271 36463 1305 36497
rect 1339 36463 1373 36497
rect 1407 36463 1441 36497
rect 1475 36463 1509 36497
rect 1543 36463 1577 36497
rect 1611 36463 1645 36497
rect 1679 36463 1713 36497
rect 1747 36463 1781 36497
rect 1815 36463 1849 36497
rect 1883 36463 1917 36497
rect 1951 36463 1985 36497
rect 2019 36463 2053 36497
rect 2087 36463 2121 36497
rect 2155 36463 2189 36497
rect 2223 36463 2257 36497
rect 2291 36463 2325 36497
rect 2359 36463 2393 36497
rect 2427 36463 2461 36497
rect 2495 36463 2529 36497
rect 2563 36463 2597 36497
rect 2631 36463 2665 36497
rect 2699 36463 2733 36497
rect 2767 36463 2801 36497
rect 2835 36463 2869 36497
rect 2903 36463 2937 36497
rect 2971 36463 3005 36497
rect 3039 36463 3073 36497
rect 3107 36463 3141 36497
rect 3175 36463 3209 36497
rect 3243 36463 3277 36497
rect 3311 36463 3345 36497
rect 3379 36463 3413 36497
rect 3447 36463 3481 36497
rect 3515 36463 3549 36497
rect 3583 36463 3617 36497
rect 3651 36463 3685 36497
rect 3719 36463 3753 36497
rect 3787 36463 3821 36497
rect 3855 36463 3889 36497
rect 3923 36463 3957 36497
rect 3991 36463 4025 36497
rect 4059 36463 4093 36497
rect 4127 36463 4161 36497
rect 4195 36463 4229 36497
rect 4263 36463 4297 36497
rect 4331 36463 4365 36497
rect 4399 36463 4433 36497
rect 4467 36463 4501 36497
rect 4535 36463 4569 36497
rect 4603 36463 4637 36497
rect 4671 36463 4705 36497
rect 4739 36463 4773 36497
rect 4807 36463 4841 36497
rect 4875 36463 4909 36497
rect 4943 36463 4977 36497
rect 5011 36463 5045 36497
rect 5079 36463 5113 36497
rect 5147 36463 5181 36497
rect 5215 36463 5249 36497
rect 5283 36463 5317 36497
rect 5351 36463 5385 36497
rect 5419 36463 5453 36497
rect 5487 36463 5521 36497
rect 5555 36463 5589 36497
rect 5623 36463 5657 36497
rect 5691 36463 5725 36497
rect 5759 36463 5793 36497
rect 5827 36463 5861 36497
rect 5895 36463 5929 36497
rect 5963 36463 5997 36497
rect 6031 36463 6065 36497
rect 6099 36463 6133 36497
rect 6167 36463 6201 36497
rect 6235 36463 6269 36497
rect 6303 36463 6337 36497
rect 6371 36463 6405 36497
rect 6439 36463 6473 36497
rect 6507 36463 6541 36497
rect 6575 36463 6609 36497
rect 6643 36463 6677 36497
rect 6711 36463 6745 36497
rect 6779 36463 6813 36497
rect 6847 36463 6881 36497
rect 6915 36463 6949 36497
rect 6983 36463 7017 36497
rect 7051 36463 7085 36497
rect 7119 36463 7153 36497
rect 7187 36463 7221 36497
rect 7255 36463 7289 36497
rect 7323 36463 7357 36497
rect 7391 36463 7425 36497
rect 7459 36463 7493 36497
rect 7527 36463 7561 36497
rect 7595 36463 7629 36497
rect 7663 36463 7697 36497
rect 7731 36463 7765 36497
rect 7799 36463 7833 36497
rect 7867 36463 7901 36497
rect 7935 36463 7969 36497
rect 8003 36463 8037 36497
rect 8071 36463 8105 36497
rect 8139 36463 8173 36497
rect 8207 36463 8241 36497
rect 8275 36463 8309 36497
rect 8343 36463 8377 36497
rect 8411 36463 8445 36497
rect 8479 36463 8513 36497
rect 8547 36463 8581 36497
rect 8615 36463 8649 36497
rect 8683 36463 8717 36497
rect 8751 36463 8785 36497
rect 8819 36463 8853 36497
rect 8887 36463 8921 36497
rect 8955 36463 8989 36497
rect 9023 36463 9057 36497
rect 9091 36463 9125 36497
rect 9159 36463 9193 36497
rect 9227 36463 9261 36497
rect 9295 36463 9329 36497
rect 9363 36463 9397 36497
rect 9431 36463 9465 36497
rect 9499 36463 9533 36497
rect 9567 36463 9601 36497
rect 9635 36463 9669 36497
rect 9703 36463 9737 36497
rect 9771 36463 9805 36497
rect 9839 36463 9873 36497
rect 9907 36463 9941 36497
rect 9975 36463 10009 36497
rect 10043 36463 10077 36497
rect 10111 36463 10145 36497
rect 10179 36463 10213 36497
rect 10247 36463 10281 36497
rect 10315 36463 10349 36497
rect 10383 36463 10417 36497
rect 10451 36463 10485 36497
rect 10519 36463 10553 36497
rect 10587 36463 10621 36497
rect 10655 36463 10689 36497
rect 10723 36463 10757 36497
rect 10791 36463 10825 36497
rect 10859 36463 10893 36497
rect 10927 36463 10961 36497
rect 10995 36463 11029 36497
rect 11063 36463 11097 36497
rect 11131 36463 11165 36497
rect 11199 36463 11233 36497
rect 11267 36463 11301 36497
rect 11335 36463 11369 36497
rect 11403 36463 11437 36497
rect 11471 36463 11505 36497
rect 11539 36463 11573 36497
rect 11607 36463 11641 36497
rect 11675 36463 11709 36497
rect 11743 36463 11777 36497
rect 11811 36463 11845 36497
rect 11879 36463 11913 36497
rect 11947 36463 11981 36497
rect 12015 36463 12049 36497
rect 12083 36463 12117 36497
rect 12151 36463 12185 36497
rect 12219 36463 12253 36497
rect 12287 36463 12321 36497
rect 12355 36463 12389 36497
rect 12423 36463 12457 36497
rect 12491 36463 12525 36497
rect 12559 36463 12593 36497
rect 12627 36463 12661 36497
rect 12695 36463 12729 36497
rect 12763 36463 12797 36497
rect 12831 36463 12865 36497
rect 12899 36463 12933 36497
rect 12967 36463 13001 36497
rect 13035 36463 13069 36497
rect 13103 36463 13137 36497
rect 13171 36463 13205 36497
rect 13239 36463 13273 36497
rect 13307 36463 13341 36497
rect 13375 36463 13409 36497
rect 13443 36463 13477 36497
rect 13511 36463 13545 36497
rect 13579 36463 13613 36497
rect 13647 36463 13681 36497
rect 13715 36463 13749 36497
rect 13783 36463 13817 36497
rect 13851 36463 13885 36497
rect 13919 36463 13953 36497
rect 13987 36463 14021 36497
rect 14055 36463 14089 36497
rect 14123 36463 14157 36497
rect 14191 36463 14225 36497
rect 14259 36463 14293 36497
rect 14327 36463 14361 36497
rect 14395 36463 14429 36497
rect 14463 36463 14497 36497
rect 312 36304 346 36338
rect 312 36236 346 36270
rect 14607 36310 14641 36344
rect 14607 36242 14641 36276
rect 312 36168 346 36202
rect 312 36100 346 36134
rect 312 36032 346 36066
rect 312 35964 346 35998
rect 312 35896 346 35930
rect 312 35828 346 35862
rect 312 35760 346 35794
rect 312 35692 346 35726
rect 312 35624 346 35658
rect 312 35556 346 35590
rect 312 35488 346 35522
rect 312 35420 346 35454
rect 312 35352 346 35386
rect 312 35284 346 35318
rect 312 35216 346 35250
rect 312 35148 346 35182
rect 312 35080 346 35114
rect 312 35012 346 35046
rect 312 34944 346 34978
rect 312 34876 346 34910
rect 312 34808 346 34842
rect 312 34740 346 34774
rect 312 34672 346 34706
rect 312 34604 346 34638
rect 312 34536 346 34570
rect 312 34468 346 34502
rect 312 34400 346 34434
rect 312 34332 346 34366
rect 312 34264 346 34298
rect 312 34196 346 34230
rect 312 34128 346 34162
rect 312 34060 346 34094
rect 312 33992 346 34026
rect 312 33924 346 33958
rect 312 33856 346 33890
rect 312 33788 346 33822
rect 312 33720 346 33754
rect 312 33652 346 33686
rect 312 33584 346 33618
rect 312 33516 346 33550
rect 312 33448 346 33482
rect 312 33380 346 33414
rect 312 33312 346 33346
rect 312 33244 346 33278
rect 312 33176 346 33210
rect 312 33108 346 33142
rect 312 33040 346 33074
rect 312 32972 346 33006
rect 312 32904 346 32938
rect 312 32836 346 32870
rect 312 32768 346 32802
rect 312 32700 346 32734
rect 312 32632 346 32666
rect 312 32564 346 32598
rect 312 32496 346 32530
rect 312 32428 346 32462
rect 312 32360 346 32394
rect 312 32292 346 32326
rect 312 32224 346 32258
rect 312 32156 346 32190
rect 312 32088 346 32122
rect 312 32020 346 32054
rect 312 31952 346 31986
rect 312 31884 346 31918
rect 312 31816 346 31850
rect 312 31748 346 31782
rect 312 31680 346 31714
rect 312 31612 346 31646
rect 312 31544 346 31578
rect 312 31476 346 31510
rect 312 31408 346 31442
rect 312 31340 346 31374
rect 312 31272 346 31306
rect 312 31204 346 31238
rect 312 31136 346 31170
rect 312 31068 346 31102
rect 312 31000 346 31034
rect 312 30932 346 30966
rect 312 30864 346 30898
rect 312 30796 346 30830
rect 312 30728 346 30762
rect 312 30660 346 30694
rect 312 30592 346 30626
rect 312 30524 346 30558
rect 312 30456 346 30490
rect 312 30388 346 30422
rect 312 30320 346 30354
rect 312 30252 346 30286
rect 312 30184 346 30218
rect 312 30116 346 30150
rect 312 30048 346 30082
rect 312 29980 346 30014
rect 312 29912 346 29946
rect 312 29844 346 29878
rect 312 29776 346 29810
rect 312 29708 346 29742
rect 312 29640 346 29674
rect 312 29572 346 29606
rect 312 29504 346 29538
rect 312 29436 346 29470
rect 312 29368 346 29402
rect 312 29300 346 29334
rect 312 29232 346 29266
rect 312 29164 346 29198
rect 312 29096 346 29130
rect 312 29028 346 29062
rect 312 28960 346 28994
rect 312 28892 346 28926
rect 312 28824 346 28858
rect 312 28756 346 28790
rect 312 28688 346 28722
rect 312 28620 346 28654
rect 312 28552 346 28586
rect 312 28484 346 28518
rect 312 28416 346 28450
rect 312 28348 346 28382
rect 312 28280 346 28314
rect 312 28212 346 28246
rect 312 28144 346 28178
rect 312 28076 346 28110
rect 312 28008 346 28042
rect 312 27940 346 27974
rect 312 27872 346 27906
rect 312 27804 346 27838
rect 312 27736 346 27770
rect 312 27668 346 27702
rect 312 27600 346 27634
rect 312 27532 346 27566
rect 312 27464 346 27498
rect 312 27396 346 27430
rect 312 27328 346 27362
rect 312 27260 346 27294
rect 312 27192 346 27226
rect 312 27124 346 27158
rect 312 27056 346 27090
rect 312 26988 346 27022
rect 312 26920 346 26954
rect 312 26852 346 26886
rect 312 26784 346 26818
rect 312 26716 346 26750
rect 312 26648 346 26682
rect 312 26580 346 26614
rect 312 26512 346 26546
rect 312 26444 346 26478
rect 312 26376 346 26410
rect 312 26308 346 26342
rect 312 26240 346 26274
rect 312 26172 346 26206
rect 312 26104 346 26138
rect 312 26036 346 26070
rect 312 25968 346 26002
rect 312 25900 346 25934
rect 312 25832 346 25866
rect 312 25764 346 25798
rect 312 25696 346 25730
rect 312 25628 346 25662
rect 312 25560 346 25594
rect 312 25492 346 25526
rect 312 25424 346 25458
rect 312 25356 346 25390
rect 312 25288 346 25322
rect 312 25220 346 25254
rect 312 25152 346 25186
rect 312 25084 346 25118
rect 312 25016 346 25050
rect 312 24948 346 24982
rect 312 24880 346 24914
rect 312 24812 346 24846
rect 312 24744 346 24778
rect 312 24676 346 24710
rect 312 24608 346 24642
rect 312 24540 346 24574
rect 312 24472 346 24506
rect 312 24404 346 24438
rect 312 24336 346 24370
rect 312 24268 346 24302
rect 312 24200 346 24234
rect 312 24132 346 24166
rect 312 24064 346 24098
rect 312 23996 346 24030
rect 312 23928 346 23962
rect 312 23860 346 23894
rect 312 23792 346 23826
rect 312 23724 346 23758
rect 312 23656 346 23690
rect 312 23588 346 23622
rect 312 23520 346 23554
rect 312 23452 346 23486
rect 312 23384 346 23418
rect 312 23316 346 23350
rect 312 23248 346 23282
rect 312 23180 346 23214
rect 312 23112 346 23146
rect 312 23044 346 23078
rect 312 22976 346 23010
rect 312 22908 346 22942
rect 312 22840 346 22874
rect 312 22772 346 22806
rect 312 22704 346 22738
rect 312 22636 346 22670
rect 312 22568 346 22602
rect 312 22500 346 22534
rect 312 22432 346 22466
rect 312 22364 346 22398
rect 312 22296 346 22330
rect 312 22228 346 22262
rect 312 22160 346 22194
rect 312 22092 346 22126
rect 312 22024 346 22058
rect 312 21956 346 21990
rect 312 21888 346 21922
rect 312 21820 346 21854
rect 312 21752 346 21786
rect 312 21684 346 21718
rect 312 21616 346 21650
rect 312 21548 346 21582
rect 312 21480 346 21514
rect 312 21412 346 21446
rect 312 21344 346 21378
rect 312 21276 346 21310
rect 312 21208 346 21242
rect 312 21140 346 21174
rect 312 21072 346 21106
rect 312 21004 346 21038
rect 312 20936 346 20970
rect 312 20868 346 20902
rect 312 20800 346 20834
rect 312 20732 346 20766
rect 312 20664 346 20698
rect 312 20596 346 20630
rect 312 20528 346 20562
rect 312 20460 346 20494
rect 312 20392 346 20426
rect 312 20324 346 20358
rect 312 20256 346 20290
rect 312 20188 346 20222
rect 312 20120 346 20154
rect 312 20052 346 20086
rect 312 19984 346 20018
rect 312 19916 346 19950
rect 312 19848 346 19882
rect 312 19780 346 19814
rect 312 19712 346 19746
rect 312 19644 346 19678
rect 312 19576 346 19610
rect 312 19508 346 19542
rect 312 19440 346 19474
rect 312 19372 346 19406
rect 312 19304 346 19338
rect 312 19236 346 19270
rect 312 19168 346 19202
rect 312 19100 346 19134
rect 312 19032 346 19066
rect 312 18964 346 18998
rect 312 18896 346 18930
rect 312 18828 346 18862
rect 312 18760 346 18794
rect 312 18692 346 18726
rect 312 18624 346 18658
rect 312 18556 346 18590
rect 312 18488 346 18522
rect 312 18420 346 18454
rect 312 18352 346 18386
rect 312 18284 346 18318
rect 312 18216 346 18250
rect 312 18148 346 18182
rect 312 18080 346 18114
rect 312 18012 346 18046
rect 312 17944 346 17978
rect 312 17876 346 17910
rect 312 17808 346 17842
rect 312 17740 346 17774
rect 312 17672 346 17706
rect 312 17604 346 17638
rect 312 17536 346 17570
rect 312 17468 346 17502
rect 312 17400 346 17434
rect 312 17332 346 17366
rect 312 17264 346 17298
rect 312 17196 346 17230
rect 312 17128 346 17162
rect 312 17060 346 17094
rect 312 16992 346 17026
rect 312 16924 346 16958
rect 312 16856 346 16890
rect 312 16788 346 16822
rect 312 16720 346 16754
rect 312 16652 346 16686
rect 312 16584 346 16618
rect 312 16516 346 16550
rect 312 16448 346 16482
rect 312 16380 346 16414
rect 312 16312 346 16346
rect 312 16244 346 16278
rect 312 16176 346 16210
rect 312 16108 346 16142
rect 312 16040 346 16074
rect 312 15972 346 16006
rect 312 15904 346 15938
rect 312 15836 346 15870
rect 312 15768 346 15802
rect 312 15700 346 15734
rect 312 15632 346 15666
rect 312 15564 346 15598
rect 312 15496 346 15530
rect 312 15428 346 15462
rect 312 15360 346 15394
rect 312 15292 346 15326
rect 312 15224 346 15258
rect 312 15156 346 15190
rect 312 15088 346 15122
rect 312 15020 346 15054
rect 312 14952 346 14986
rect 312 14884 346 14918
rect 312 14816 346 14850
rect 312 14748 346 14782
rect 312 14680 346 14714
rect 312 14612 346 14646
rect 312 14544 346 14578
rect 312 14476 346 14510
rect 312 14408 346 14442
rect 312 14340 346 14374
rect 312 14272 346 14306
rect 312 14204 346 14238
rect 312 14136 346 14170
rect 312 14068 346 14102
rect 312 14000 346 14034
rect 312 13932 346 13966
rect 312 13864 346 13898
rect 312 13796 346 13830
rect 312 13728 346 13762
rect 312 13660 346 13694
rect 312 13592 346 13626
rect 312 13524 346 13558
rect 312 13456 346 13490
rect 312 13388 346 13422
rect 312 13320 346 13354
rect 312 13252 346 13286
rect 312 13184 346 13218
rect 312 13116 346 13150
rect 312 13048 346 13082
rect 312 12980 346 13014
rect 312 12912 346 12946
rect 312 12844 346 12878
rect 312 12776 346 12810
rect 312 12708 346 12742
rect 312 12640 346 12674
rect 312 12572 346 12606
rect 312 12504 346 12538
rect 312 12436 346 12470
rect 312 12368 346 12402
rect 312 12300 346 12334
rect 312 12232 346 12266
rect 312 12164 346 12198
rect 312 12096 346 12130
rect 312 12028 346 12062
rect 312 11960 346 11994
rect 312 11892 346 11926
rect 312 11824 346 11858
rect 312 11756 346 11790
rect 312 11688 346 11722
rect 312 11620 346 11654
rect 312 11552 346 11586
rect 312 11484 346 11518
rect 312 11416 346 11450
rect 312 11348 346 11382
rect 312 11280 346 11314
rect 312 11212 346 11246
rect 312 11144 346 11178
rect 312 11076 346 11110
rect 312 11008 346 11042
rect 312 10940 346 10974
rect 312 10872 346 10906
rect 312 10804 346 10838
rect 312 10736 346 10770
rect 312 10668 346 10702
rect 312 10600 346 10634
rect 312 10532 346 10566
rect 312 10464 346 10498
rect 312 10396 346 10430
rect 312 10328 346 10362
rect 312 10260 346 10294
rect 312 10192 346 10226
rect 312 10124 346 10158
rect 312 10056 346 10090
rect 312 9988 346 10022
rect 312 9920 346 9954
rect 312 9852 346 9886
rect 312 9784 346 9818
rect 312 9716 346 9750
rect 1305 34645 1339 34679
rect 1373 34645 1407 34679
rect 1441 34645 1475 34679
rect 1509 34645 1543 34679
rect 1577 34645 1611 34679
rect 1645 34645 1679 34679
rect 1713 34645 1747 34679
rect 1781 34645 1815 34679
rect 1849 34645 1883 34679
rect 1917 34645 1951 34679
rect 1985 34645 2019 34679
rect 2053 34645 2087 34679
rect 2121 34645 2155 34679
rect 2189 34645 2223 34679
rect 2257 34645 2291 34679
rect 2325 34645 2359 34679
rect 2393 34645 2427 34679
rect 2461 34645 2495 34679
rect 2529 34645 2563 34679
rect 2597 34645 2631 34679
rect 2665 34645 2699 34679
rect 2733 34645 2767 34679
rect 2801 34645 2835 34679
rect 2869 34645 2903 34679
rect 2937 34645 2971 34679
rect 3005 34645 3039 34679
rect 3073 34645 3107 34679
rect 3141 34645 3175 34679
rect 3209 34645 3243 34679
rect 3277 34645 3311 34679
rect 3345 34645 3379 34679
rect 3413 34645 3447 34679
rect 3481 34645 3515 34679
rect 3549 34645 3583 34679
rect 3617 34645 3651 34679
rect 3685 34645 3719 34679
rect 3753 34645 3787 34679
rect 3821 34645 3855 34679
rect 3889 34645 3923 34679
rect 3957 34645 3991 34679
rect 4025 34645 4059 34679
rect 4093 34645 4127 34679
rect 4161 34645 4195 34679
rect 4229 34645 4263 34679
rect 4297 34645 4331 34679
rect 4365 34645 4399 34679
rect 4433 34645 4467 34679
rect 4501 34645 4535 34679
rect 4569 34645 4603 34679
rect 4637 34645 4671 34679
rect 4705 34645 4739 34679
rect 4773 34645 4807 34679
rect 4841 34645 4875 34679
rect 4909 34645 4943 34679
rect 4977 34645 5011 34679
rect 5045 34645 5079 34679
rect 5113 34645 5147 34679
rect 5181 34645 5215 34679
rect 5249 34645 5283 34679
rect 5317 34645 5351 34679
rect 5385 34645 5419 34679
rect 5453 34645 5487 34679
rect 5521 34645 5555 34679
rect 5589 34645 5623 34679
rect 5657 34645 5691 34679
rect 5725 34645 5759 34679
rect 5793 34645 5827 34679
rect 5861 34645 5895 34679
rect 5929 34645 5963 34679
rect 5997 34645 6031 34679
rect 6065 34645 6099 34679
rect 6133 34645 6167 34679
rect 6201 34645 6235 34679
rect 6269 34645 6303 34679
rect 6337 34645 6371 34679
rect 6405 34645 6439 34679
rect 6473 34645 6507 34679
rect 6541 34645 6575 34679
rect 6609 34645 6643 34679
rect 6677 34645 6711 34679
rect 6745 34645 6779 34679
rect 6813 34645 6847 34679
rect 6881 34645 6915 34679
rect 6949 34645 6983 34679
rect 7017 34645 7051 34679
rect 7085 34645 7119 34679
rect 7153 34645 7187 34679
rect 7221 34645 7255 34679
rect 7289 34645 7323 34679
rect 7357 34645 7391 34679
rect 7425 34645 7459 34679
rect 7493 34645 7527 34679
rect 7561 34645 7595 34679
rect 7629 34645 7663 34679
rect 7697 34645 7731 34679
rect 7765 34645 7799 34679
rect 7833 34645 7867 34679
rect 7901 34645 7935 34679
rect 7969 34645 8003 34679
rect 8037 34645 8071 34679
rect 8105 34645 8139 34679
rect 8173 34645 8207 34679
rect 8241 34645 8275 34679
rect 8309 34645 8343 34679
rect 8377 34645 8411 34679
rect 8445 34645 8479 34679
rect 8513 34645 8547 34679
rect 8581 34645 8615 34679
rect 8649 34645 8683 34679
rect 8717 34645 8751 34679
rect 8785 34645 8819 34679
rect 8853 34645 8887 34679
rect 8921 34645 8955 34679
rect 8989 34645 9023 34679
rect 9057 34645 9091 34679
rect 9125 34645 9159 34679
rect 9193 34645 9227 34679
rect 9261 34645 9295 34679
rect 9329 34645 9363 34679
rect 9397 34645 9431 34679
rect 9465 34645 9499 34679
rect 9533 34645 9567 34679
rect 9601 34645 9635 34679
rect 9669 34645 9703 34679
rect 9737 34645 9771 34679
rect 9805 34645 9839 34679
rect 9873 34645 9907 34679
rect 9941 34645 9975 34679
rect 10009 34645 10043 34679
rect 10077 34645 10111 34679
rect 10145 34645 10179 34679
rect 10213 34645 10247 34679
rect 10281 34645 10315 34679
rect 10349 34645 10383 34679
rect 10417 34645 10451 34679
rect 10485 34645 10519 34679
rect 10553 34645 10587 34679
rect 10621 34645 10655 34679
rect 10689 34645 10723 34679
rect 10757 34645 10791 34679
rect 10825 34645 10859 34679
rect 10893 34645 10927 34679
rect 10961 34645 10995 34679
rect 11029 34645 11063 34679
rect 11097 34645 11131 34679
rect 11165 34645 11199 34679
rect 11233 34645 11267 34679
rect 11301 34645 11335 34679
rect 11369 34645 11403 34679
rect 11437 34645 11471 34679
rect 11505 34645 11539 34679
rect 11573 34645 11607 34679
rect 11641 34645 11675 34679
rect 11709 34645 11743 34679
rect 11777 34645 11811 34679
rect 11845 34645 11879 34679
rect 11913 34645 11947 34679
rect 11981 34645 12015 34679
rect 12049 34645 12083 34679
rect 12117 34645 12151 34679
rect 12185 34645 12219 34679
rect 12253 34645 12287 34679
rect 12321 34645 12355 34679
rect 12389 34645 12423 34679
rect 12457 34645 12491 34679
rect 12525 34645 12559 34679
rect 12593 34645 12627 34679
rect 12661 34645 12695 34679
rect 12729 34645 12763 34679
rect 12797 34645 12831 34679
rect 12865 34645 12899 34679
rect 12933 34645 12967 34679
rect 13001 34645 13035 34679
rect 13069 34645 13103 34679
rect 13137 34645 13171 34679
rect 13205 34645 13239 34679
rect 13273 34645 13307 34679
rect 13341 34645 13375 34679
rect 13409 34645 13443 34679
rect 13477 34645 13511 34679
rect 13545 34645 13579 34679
rect 13613 34645 13647 34679
rect 13681 34645 13715 34679
rect 1161 34444 1195 34478
rect 1161 34376 1195 34410
rect 1161 34308 1195 34342
rect 1161 34240 1195 34274
rect 1161 34172 1195 34206
rect 1161 34104 1195 34138
rect 1161 34036 1195 34070
rect 1161 33968 1195 34002
rect 1161 33900 1195 33934
rect 1161 33832 1195 33866
rect 1161 33764 1195 33798
rect 1161 33696 1195 33730
rect 1161 33628 1195 33662
rect 1161 33560 1195 33594
rect 1161 33492 1195 33526
rect 1161 33424 1195 33458
rect 1161 33356 1195 33390
rect 1161 33288 1195 33322
rect 1161 33220 1195 33254
rect 1161 33152 1195 33186
rect 1161 33084 1195 33118
rect 1161 33016 1195 33050
rect 1161 32948 1195 32982
rect 1161 32880 1195 32914
rect 1161 32812 1195 32846
rect 1161 32744 1195 32778
rect 1161 32676 1195 32710
rect 1161 32608 1195 32642
rect 1161 32540 1195 32574
rect 1161 32472 1195 32506
rect 1161 32404 1195 32438
rect 1161 32336 1195 32370
rect 1161 32268 1195 32302
rect 1161 32200 1195 32234
rect 1161 32132 1195 32166
rect 1161 32064 1195 32098
rect 1161 31996 1195 32030
rect 1161 31928 1195 31962
rect 1161 31860 1195 31894
rect 1161 31792 1195 31826
rect 1161 31724 1195 31758
rect 1161 31656 1195 31690
rect 1161 31588 1195 31622
rect 1161 31520 1195 31554
rect 1161 31452 1195 31486
rect 1161 31384 1195 31418
rect 1161 31316 1195 31350
rect 1161 31248 1195 31282
rect 1161 31180 1195 31214
rect 1161 31112 1195 31146
rect 1161 31044 1195 31078
rect 1161 30976 1195 31010
rect 1161 30908 1195 30942
rect 1161 30840 1195 30874
rect 1161 30772 1195 30806
rect 1161 30704 1195 30738
rect 1161 30636 1195 30670
rect 1161 30568 1195 30602
rect 1161 30500 1195 30534
rect 1161 30432 1195 30466
rect 1161 30364 1195 30398
rect 1161 30296 1195 30330
rect 1161 30228 1195 30262
rect 1161 30160 1195 30194
rect 1161 30092 1195 30126
rect 1161 30024 1195 30058
rect 1161 29956 1195 29990
rect 1161 29888 1195 29922
rect 1161 29820 1195 29854
rect 1161 29752 1195 29786
rect 1161 29684 1195 29718
rect 1161 29616 1195 29650
rect 1161 29548 1195 29582
rect 1161 29480 1195 29514
rect 1161 29412 1195 29446
rect 1161 29344 1195 29378
rect 1161 29276 1195 29310
rect 1161 29208 1195 29242
rect 1161 29140 1195 29174
rect 1161 29072 1195 29106
rect 1161 29004 1195 29038
rect 1161 28936 1195 28970
rect 13809 34439 13843 34473
rect 13809 34371 13843 34405
rect 13809 34303 13843 34337
rect 13809 34235 13843 34269
rect 13809 34167 13843 34201
rect 13809 34099 13843 34133
rect 13809 34031 13843 34065
rect 13809 33963 13843 33997
rect 13809 33895 13843 33929
rect 13809 33827 13843 33861
rect 13809 33759 13843 33793
rect 13809 33691 13843 33725
rect 13809 33623 13843 33657
rect 13809 33555 13843 33589
rect 13809 33487 13843 33521
rect 13809 33419 13843 33453
rect 13809 33351 13843 33385
rect 13809 33283 13843 33317
rect 13809 33215 13843 33249
rect 13809 33147 13843 33181
rect 13809 33079 13843 33113
rect 13809 33011 13843 33045
rect 13809 32943 13843 32977
rect 13809 32875 13843 32909
rect 13809 32807 13843 32841
rect 13809 32739 13843 32773
rect 13809 32671 13843 32705
rect 13809 32603 13843 32637
rect 13809 32535 13843 32569
rect 13809 32467 13843 32501
rect 13809 32399 13843 32433
rect 13809 32331 13843 32365
rect 13809 32263 13843 32297
rect 13809 32195 13843 32229
rect 13809 32127 13843 32161
rect 13809 32059 13843 32093
rect 13809 31991 13843 32025
rect 13809 31923 13843 31957
rect 13809 31855 13843 31889
rect 13809 31787 13843 31821
rect 13809 31719 13843 31753
rect 13809 31651 13843 31685
rect 13809 31583 13843 31617
rect 13809 31515 13843 31549
rect 13809 31447 13843 31481
rect 13809 31379 13843 31413
rect 13809 31311 13843 31345
rect 13809 31243 13843 31277
rect 13809 31175 13843 31209
rect 13809 31107 13843 31141
rect 13809 31039 13843 31073
rect 13809 30971 13843 31005
rect 13809 30903 13843 30937
rect 13809 30835 13843 30869
rect 13809 30767 13843 30801
rect 13809 30699 13843 30733
rect 13809 30631 13843 30665
rect 13809 30563 13843 30597
rect 13809 30495 13843 30529
rect 13809 30427 13843 30461
rect 13809 30359 13843 30393
rect 13809 30291 13843 30325
rect 13809 30223 13843 30257
rect 13809 30155 13843 30189
rect 13809 30087 13843 30121
rect 13809 30019 13843 30053
rect 13809 29951 13843 29985
rect 13809 29883 13843 29917
rect 13809 29815 13843 29849
rect 13809 29747 13843 29781
rect 13809 29679 13843 29713
rect 13809 29611 13843 29645
rect 13809 29543 13843 29577
rect 13809 29475 13843 29509
rect 13809 29407 13843 29441
rect 13809 29339 13843 29373
rect 13809 29271 13843 29305
rect 13809 29203 13843 29237
rect 13809 29135 13843 29169
rect 13809 29067 13843 29101
rect 13809 28999 13843 29033
rect 13809 28931 13843 28965
rect 1161 28868 1195 28902
rect 1161 28800 1195 28834
rect 1161 28732 1195 28766
rect 1161 28664 1195 28698
rect 1161 28596 1195 28630
rect 1161 28528 1195 28562
rect 1161 28460 1195 28494
rect 1161 28392 1195 28426
rect 1161 28324 1195 28358
rect 1161 28256 1195 28290
rect 1161 28188 1195 28222
rect 1161 28120 1195 28154
rect 1161 28052 1195 28086
rect 1161 27984 1195 28018
rect 1161 27916 1195 27950
rect 1161 27848 1195 27882
rect 1161 27780 1195 27814
rect 1161 27712 1195 27746
rect 1161 27644 1195 27678
rect 1161 27576 1195 27610
rect 1161 27508 1195 27542
rect 1161 27440 1195 27474
rect 1161 27372 1195 27406
rect 1161 27304 1195 27338
rect 1161 27236 1195 27270
rect 1161 27168 1195 27202
rect 1161 27100 1195 27134
rect 1161 27032 1195 27066
rect 13809 28863 13843 28897
rect 13809 28795 13843 28829
rect 13809 28727 13843 28761
rect 13809 28659 13843 28693
rect 13809 28591 13843 28625
rect 13809 28523 13843 28557
rect 13809 28455 13843 28489
rect 13809 28387 13843 28421
rect 13809 28319 13843 28353
rect 13809 28251 13843 28285
rect 13809 28183 13843 28217
rect 13809 28115 13843 28149
rect 13809 28047 13843 28081
rect 13809 27979 13843 28013
rect 13809 27911 13843 27945
rect 13809 27843 13843 27877
rect 13809 27775 13843 27809
rect 13809 27707 13843 27741
rect 13809 27639 13843 27673
rect 13809 27571 13843 27605
rect 13809 27503 13843 27537
rect 13809 27435 13843 27469
rect 13809 27367 13843 27401
rect 13809 27299 13843 27333
rect 13809 27231 13843 27265
rect 13809 27163 13843 27197
rect 13809 27095 13843 27129
rect 13809 27027 13843 27061
rect 1161 26964 1195 26998
rect 1161 26896 1195 26930
rect 1161 26828 1195 26862
rect 1161 26760 1195 26794
rect 1161 26692 1195 26726
rect 1161 26624 1195 26658
rect 1161 26556 1195 26590
rect 1161 26488 1195 26522
rect 1161 26420 1195 26454
rect 1161 26352 1195 26386
rect 1161 26284 1195 26318
rect 1161 26216 1195 26250
rect 1161 26148 1195 26182
rect 1161 26080 1195 26114
rect 1161 26012 1195 26046
rect 1161 25944 1195 25978
rect 1161 25876 1195 25910
rect 1161 25808 1195 25842
rect 1161 25740 1195 25774
rect 1161 25672 1195 25706
rect 1161 25604 1195 25638
rect 1161 25536 1195 25570
rect 1161 25468 1195 25502
rect 1161 25400 1195 25434
rect 1161 25332 1195 25366
rect 1161 25264 1195 25298
rect 1161 25196 1195 25230
rect 1161 25128 1195 25162
rect 1161 25060 1195 25094
rect 1161 24992 1195 25026
rect 1161 24924 1195 24958
rect 1161 24856 1195 24890
rect 1161 24788 1195 24822
rect 1161 24720 1195 24754
rect 1161 24652 1195 24686
rect 1161 24584 1195 24618
rect 1161 24516 1195 24550
rect 1161 24448 1195 24482
rect 1161 24380 1195 24414
rect 1161 24312 1195 24346
rect 1161 24244 1195 24278
rect 1161 24176 1195 24210
rect 1161 24108 1195 24142
rect 1161 24040 1195 24074
rect 1161 23972 1195 24006
rect 1161 23904 1195 23938
rect 1161 23836 1195 23870
rect 1161 23768 1195 23802
rect 1161 23700 1195 23734
rect 1161 23632 1195 23666
rect 1161 23564 1195 23598
rect 1161 23496 1195 23530
rect 1161 23428 1195 23462
rect 1161 23360 1195 23394
rect 1161 23292 1195 23326
rect 1161 23224 1195 23258
rect 1161 23156 1195 23190
rect 1161 23088 1195 23122
rect 1161 23020 1195 23054
rect 1161 22952 1195 22986
rect 1161 22884 1195 22918
rect 1161 22816 1195 22850
rect 1161 22748 1195 22782
rect 1161 22680 1195 22714
rect 1161 22612 1195 22646
rect 1161 22544 1195 22578
rect 1161 22476 1195 22510
rect 1161 22408 1195 22442
rect 1161 22340 1195 22374
rect 1161 22272 1195 22306
rect 1161 22204 1195 22238
rect 1161 22136 1195 22170
rect 1161 22068 1195 22102
rect 1161 22000 1195 22034
rect 1161 21932 1195 21966
rect 1161 21864 1195 21898
rect 1161 21796 1195 21830
rect 1161 21728 1195 21762
rect 1161 21660 1195 21694
rect 1161 21592 1195 21626
rect 1161 21524 1195 21558
rect 1161 21456 1195 21490
rect 1161 21388 1195 21422
rect 1161 21320 1195 21354
rect 1161 21252 1195 21286
rect 1161 21184 1195 21218
rect 1161 21116 1195 21150
rect 1161 21048 1195 21082
rect 1161 20980 1195 21014
rect 1161 20912 1195 20946
rect 1161 20844 1195 20878
rect 1161 20776 1195 20810
rect 1161 20708 1195 20742
rect 1161 20640 1195 20674
rect 1161 20572 1195 20606
rect 1161 20504 1195 20538
rect 1161 20436 1195 20470
rect 1161 20368 1195 20402
rect 1161 20300 1195 20334
rect 1161 20232 1195 20266
rect 1161 20164 1195 20198
rect 1161 20096 1195 20130
rect 1161 20028 1195 20062
rect 1161 19960 1195 19994
rect 1161 19892 1195 19926
rect 1161 19824 1195 19858
rect 1161 19756 1195 19790
rect 1161 19688 1195 19722
rect 1161 19620 1195 19654
rect 1161 19552 1195 19586
rect 1161 19484 1195 19518
rect 1161 19416 1195 19450
rect 1161 19348 1195 19382
rect 1161 19280 1195 19314
rect 1161 19212 1195 19246
rect 1161 19144 1195 19178
rect 1161 19076 1195 19110
rect 1161 19008 1195 19042
rect 1161 18940 1195 18974
rect 1161 18872 1195 18906
rect 1161 18804 1195 18838
rect 1161 18736 1195 18770
rect 1161 18668 1195 18702
rect 1161 18600 1195 18634
rect 1161 18532 1195 18566
rect 1161 18464 1195 18498
rect 1161 18396 1195 18430
rect 1161 18328 1195 18362
rect 1161 18260 1195 18294
rect 1161 18192 1195 18226
rect 1161 18124 1195 18158
rect 1161 18056 1195 18090
rect 1161 17988 1195 18022
rect 1161 17920 1195 17954
rect 1161 17852 1195 17886
rect 1161 17784 1195 17818
rect 1161 17716 1195 17750
rect 1161 17648 1195 17682
rect 1161 17580 1195 17614
rect 1161 17512 1195 17546
rect 1161 17444 1195 17478
rect 1161 17376 1195 17410
rect 1161 17308 1195 17342
rect 1161 17240 1195 17274
rect 1161 17172 1195 17206
rect 1161 17104 1195 17138
rect 1161 17036 1195 17070
rect 1161 16968 1195 17002
rect 1161 16900 1195 16934
rect 1161 16832 1195 16866
rect 1161 16764 1195 16798
rect 1161 16696 1195 16730
rect 1161 16628 1195 16662
rect 1161 16560 1195 16594
rect 1161 16492 1195 16526
rect 1161 16424 1195 16458
rect 1161 16356 1195 16390
rect 1161 16288 1195 16322
rect 1161 16220 1195 16254
rect 1161 16152 1195 16186
rect 1161 16084 1195 16118
rect 1161 16016 1195 16050
rect 1161 15948 1195 15982
rect 1161 15880 1195 15914
rect 1161 15812 1195 15846
rect 1161 15744 1195 15778
rect 1161 15676 1195 15710
rect 1161 15608 1195 15642
rect 1161 15540 1195 15574
rect 1161 15472 1195 15506
rect 1161 15404 1195 15438
rect 1161 15336 1195 15370
rect 1161 15268 1195 15302
rect 1161 15200 1195 15234
rect 1161 15132 1195 15166
rect 1161 15064 1195 15098
rect 1161 14996 1195 15030
rect 1161 14928 1195 14962
rect 1161 14860 1195 14894
rect 1161 14792 1195 14826
rect 1161 14724 1195 14758
rect 1161 14656 1195 14690
rect 1161 14588 1195 14622
rect 1161 14520 1195 14554
rect 1161 14452 1195 14486
rect 1161 14384 1195 14418
rect 1161 14316 1195 14350
rect 1161 14248 1195 14282
rect 1161 14180 1195 14214
rect 1161 14112 1195 14146
rect 1161 14044 1195 14078
rect 1161 13976 1195 14010
rect 1161 13908 1195 13942
rect 1161 13840 1195 13874
rect 1161 13772 1195 13806
rect 1161 13704 1195 13738
rect 1161 13636 1195 13670
rect 1161 13568 1195 13602
rect 1161 13500 1195 13534
rect 1161 13432 1195 13466
rect 1161 13364 1195 13398
rect 1161 13296 1195 13330
rect 1161 13228 1195 13262
rect 1161 13160 1195 13194
rect 1161 13092 1195 13126
rect 1161 13024 1195 13058
rect 1161 12956 1195 12990
rect 1161 12888 1195 12922
rect 1161 12820 1195 12854
rect 1161 12752 1195 12786
rect 1161 12684 1195 12718
rect 1161 12616 1195 12650
rect 1161 12548 1195 12582
rect 1161 12480 1195 12514
rect 1161 12412 1195 12446
rect 1161 12344 1195 12378
rect 1161 12276 1195 12310
rect 1161 12208 1195 12242
rect 1161 12140 1195 12174
rect 1161 12072 1195 12106
rect 1161 12004 1195 12038
rect 1161 11936 1195 11970
rect 1161 11868 1195 11902
rect 1161 11800 1195 11834
rect 1161 11732 1195 11766
rect 1161 11664 1195 11698
rect 1161 11596 1195 11630
rect 1161 11528 1195 11562
rect 1161 11460 1195 11494
rect 1161 11392 1195 11426
rect 1161 11324 1195 11358
rect 1161 11256 1195 11290
rect 1161 11188 1195 11222
rect 1161 11120 1195 11154
rect 1161 11052 1195 11086
rect 1161 10984 1195 11018
rect 1161 10916 1195 10950
rect 1161 10848 1195 10882
rect 1161 10780 1195 10814
rect 1161 10712 1195 10746
rect 1161 10644 1195 10678
rect 1161 10576 1195 10610
rect 1161 10508 1195 10542
rect 1161 10440 1195 10474
rect 1161 10372 1195 10406
rect 13809 26959 13843 26993
rect 13809 26891 13843 26925
rect 13809 26823 13843 26857
rect 13809 26755 13843 26789
rect 13809 26687 13843 26721
rect 13809 26619 13843 26653
rect 13809 26551 13843 26585
rect 13809 26483 13843 26517
rect 13809 26415 13843 26449
rect 13809 26347 13843 26381
rect 13809 26279 13843 26313
rect 13809 26211 13843 26245
rect 13809 26143 13843 26177
rect 13809 26075 13843 26109
rect 13809 26007 13843 26041
rect 13809 25939 13843 25973
rect 13809 25871 13843 25905
rect 13809 25803 13843 25837
rect 13809 25735 13843 25769
rect 13809 25667 13843 25701
rect 13809 25599 13843 25633
rect 13809 25531 13843 25565
rect 13809 25463 13843 25497
rect 13809 25395 13843 25429
rect 13809 25327 13843 25361
rect 13809 25259 13843 25293
rect 13809 25191 13843 25225
rect 13809 25123 13843 25157
rect 13809 25055 13843 25089
rect 13809 24987 13843 25021
rect 13809 24919 13843 24953
rect 13809 24851 13843 24885
rect 13809 24783 13843 24817
rect 13809 24715 13843 24749
rect 13809 24647 13843 24681
rect 13809 24579 13843 24613
rect 13809 24511 13843 24545
rect 13809 24443 13843 24477
rect 13809 24375 13843 24409
rect 13809 24307 13843 24341
rect 13809 24239 13843 24273
rect 13809 24171 13843 24205
rect 13809 24103 13843 24137
rect 13809 24035 13843 24069
rect 13809 23967 13843 24001
rect 13809 23899 13843 23933
rect 13809 23831 13843 23865
rect 13809 23763 13843 23797
rect 13809 23695 13843 23729
rect 13809 23627 13843 23661
rect 13809 23559 13843 23593
rect 13809 23491 13843 23525
rect 13809 23423 13843 23457
rect 13809 23355 13843 23389
rect 13809 23287 13843 23321
rect 13809 23219 13843 23253
rect 13809 23151 13843 23185
rect 13809 23083 13843 23117
rect 13809 23015 13843 23049
rect 13809 22947 13843 22981
rect 13809 22879 13843 22913
rect 13809 22811 13843 22845
rect 13809 22743 13843 22777
rect 13809 22675 13843 22709
rect 13809 22607 13843 22641
rect 13809 22539 13843 22573
rect 13809 22471 13843 22505
rect 13809 22403 13843 22437
rect 13809 22335 13843 22369
rect 13809 22267 13843 22301
rect 13809 22199 13843 22233
rect 13809 22131 13843 22165
rect 13809 22063 13843 22097
rect 13809 21995 13843 22029
rect 13809 21927 13843 21961
rect 13809 21859 13843 21893
rect 13809 21791 13843 21825
rect 13809 21723 13843 21757
rect 13809 21655 13843 21689
rect 13809 21587 13843 21621
rect 13809 21519 13843 21553
rect 13809 21451 13843 21485
rect 13809 21383 13843 21417
rect 13809 21315 13843 21349
rect 13809 21247 13843 21281
rect 13809 21179 13843 21213
rect 13809 21111 13843 21145
rect 13809 21043 13843 21077
rect 13809 20975 13843 21009
rect 13809 20907 13843 20941
rect 13809 20839 13843 20873
rect 13809 20771 13843 20805
rect 13809 20703 13843 20737
rect 13809 20635 13843 20669
rect 13809 20567 13843 20601
rect 13809 20499 13843 20533
rect 13809 20431 13843 20465
rect 13809 20363 13843 20397
rect 13809 20295 13843 20329
rect 13809 20227 13843 20261
rect 13809 20159 13843 20193
rect 13809 20091 13843 20125
rect 13809 20023 13843 20057
rect 13809 19955 13843 19989
rect 13809 19887 13843 19921
rect 13809 19819 13843 19853
rect 13809 19751 13843 19785
rect 13809 19683 13843 19717
rect 13809 19615 13843 19649
rect 13809 19547 13843 19581
rect 13809 19479 13843 19513
rect 13809 19411 13843 19445
rect 13809 19343 13843 19377
rect 13809 19275 13843 19309
rect 13809 19207 13843 19241
rect 13809 19139 13843 19173
rect 13809 19071 13843 19105
rect 13809 19003 13843 19037
rect 13809 18935 13843 18969
rect 13809 18867 13843 18901
rect 13809 18799 13843 18833
rect 13809 18731 13843 18765
rect 13809 18663 13843 18697
rect 13809 18595 13843 18629
rect 13809 18527 13843 18561
rect 13809 18459 13843 18493
rect 13809 18391 13843 18425
rect 13809 18323 13843 18357
rect 13809 18255 13843 18289
rect 13809 18187 13843 18221
rect 13809 18119 13843 18153
rect 13809 18051 13843 18085
rect 13809 17983 13843 18017
rect 13809 17915 13843 17949
rect 13809 17847 13843 17881
rect 13809 17779 13843 17813
rect 13809 17711 13843 17745
rect 13809 17643 13843 17677
rect 13809 17575 13843 17609
rect 13809 17507 13843 17541
rect 13809 17439 13843 17473
rect 13809 17371 13843 17405
rect 13809 17303 13843 17337
rect 13809 17235 13843 17269
rect 13809 17167 13843 17201
rect 13809 17099 13843 17133
rect 13809 17031 13843 17065
rect 13809 16963 13843 16997
rect 13809 16895 13843 16929
rect 13809 16827 13843 16861
rect 13809 16759 13843 16793
rect 13809 16691 13843 16725
rect 13809 16623 13843 16657
rect 13809 16555 13843 16589
rect 13809 16487 13843 16521
rect 13809 16419 13843 16453
rect 13809 16351 13843 16385
rect 13809 16283 13843 16317
rect 13809 16215 13843 16249
rect 13809 16147 13843 16181
rect 13809 16079 13843 16113
rect 13809 16011 13843 16045
rect 13809 15943 13843 15977
rect 13809 15875 13843 15909
rect 13809 15807 13843 15841
rect 13809 15739 13843 15773
rect 13809 15671 13843 15705
rect 13809 15603 13843 15637
rect 13809 15535 13843 15569
rect 13809 15467 13843 15501
rect 13809 15399 13843 15433
rect 13809 15331 13843 15365
rect 13809 15263 13843 15297
rect 13809 15195 13843 15229
rect 13809 15127 13843 15161
rect 13809 15059 13843 15093
rect 13809 14991 13843 15025
rect 13809 14923 13843 14957
rect 13809 14855 13843 14889
rect 13809 14787 13843 14821
rect 13809 14719 13843 14753
rect 13809 14651 13843 14685
rect 13809 14583 13843 14617
rect 13809 14515 13843 14549
rect 13809 14447 13843 14481
rect 13809 14379 13843 14413
rect 13809 14311 13843 14345
rect 13809 14243 13843 14277
rect 13809 14175 13843 14209
rect 13809 14107 13843 14141
rect 13809 14039 13843 14073
rect 13809 13971 13843 14005
rect 13809 13903 13843 13937
rect 13809 13835 13843 13869
rect 13809 13767 13843 13801
rect 13809 13699 13843 13733
rect 13809 13631 13843 13665
rect 13809 13563 13843 13597
rect 13809 13495 13843 13529
rect 13809 13427 13843 13461
rect 13809 13359 13843 13393
rect 13809 13291 13843 13325
rect 13809 13223 13843 13257
rect 13809 13155 13843 13189
rect 13809 13087 13843 13121
rect 13809 13019 13843 13053
rect 13809 12951 13843 12985
rect 13809 12883 13843 12917
rect 13809 12815 13843 12849
rect 13809 12747 13843 12781
rect 13809 12679 13843 12713
rect 13809 12611 13843 12645
rect 13809 12543 13843 12577
rect 13809 12475 13843 12509
rect 13809 12407 13843 12441
rect 13809 12339 13843 12373
rect 13809 12271 13843 12305
rect 13809 12203 13843 12237
rect 13809 12135 13843 12169
rect 13809 12067 13843 12101
rect 13809 11999 13843 12033
rect 13809 11931 13843 11965
rect 13809 11863 13843 11897
rect 13809 11795 13843 11829
rect 13809 11727 13843 11761
rect 13809 11659 13843 11693
rect 13809 11591 13843 11625
rect 13809 11523 13843 11557
rect 13809 11455 13843 11489
rect 13809 11387 13843 11421
rect 13809 11319 13843 11353
rect 13809 11251 13843 11285
rect 13809 11183 13843 11217
rect 13809 11115 13843 11149
rect 13809 11047 13843 11081
rect 13809 10979 13843 11013
rect 13809 10911 13843 10945
rect 13809 10843 13843 10877
rect 13809 10775 13843 10809
rect 13809 10707 13843 10741
rect 13809 10639 13843 10673
rect 13809 10571 13843 10605
rect 13809 10503 13843 10537
rect 13809 10435 13843 10469
rect 13809 10367 13843 10401
rect 1302 10244 1336 10278
rect 1370 10244 1404 10278
rect 1438 10244 1472 10278
rect 1506 10244 1540 10278
rect 1574 10244 1608 10278
rect 1642 10244 1676 10278
rect 1710 10244 1744 10278
rect 1778 10244 1812 10278
rect 1846 10244 1880 10278
rect 1914 10244 1948 10278
rect 1982 10244 2016 10278
rect 2050 10244 2084 10278
rect 2118 10244 2152 10278
rect 2186 10244 2220 10278
rect 2254 10244 2288 10278
rect 2322 10244 2356 10278
rect 2390 10244 2424 10278
rect 2458 10244 2492 10278
rect 2526 10244 2560 10278
rect 2594 10244 2628 10278
rect 2662 10244 2696 10278
rect 2730 10244 2764 10278
rect 2798 10244 2832 10278
rect 2866 10244 2900 10278
rect 2934 10244 2968 10278
rect 3002 10244 3036 10278
rect 3070 10244 3104 10278
rect 3138 10244 3172 10278
rect 3206 10244 3240 10278
rect 3274 10244 3308 10278
rect 3342 10244 3376 10278
rect 3410 10244 3444 10278
rect 3478 10244 3512 10278
rect 3546 10244 3580 10278
rect 3614 10244 3648 10278
rect 3682 10244 3716 10278
rect 3750 10244 3784 10278
rect 3818 10244 3852 10278
rect 3886 10244 3920 10278
rect 3954 10244 3988 10278
rect 4022 10244 4056 10278
rect 4090 10244 4124 10278
rect 4158 10244 4192 10278
rect 4226 10244 4260 10278
rect 4294 10244 4328 10278
rect 4362 10244 4396 10278
rect 4430 10244 4464 10278
rect 4498 10244 4532 10278
rect 4566 10244 4600 10278
rect 4634 10244 4668 10278
rect 4702 10244 4736 10278
rect 4770 10244 4804 10278
rect 4838 10244 4872 10278
rect 4906 10244 4940 10278
rect 4974 10244 5008 10278
rect 5042 10244 5076 10278
rect 5110 10244 5144 10278
rect 5178 10244 5212 10278
rect 5246 10244 5280 10278
rect 5314 10244 5348 10278
rect 5382 10244 5416 10278
rect 5450 10244 5484 10278
rect 5518 10244 5552 10278
rect 5586 10244 5620 10278
rect 5654 10244 5688 10278
rect 5722 10244 5756 10278
rect 5790 10244 5824 10278
rect 5858 10244 5892 10278
rect 5926 10244 5960 10278
rect 5994 10244 6028 10278
rect 6062 10244 6096 10278
rect 6130 10244 6164 10278
rect 6198 10244 6232 10278
rect 6266 10244 6300 10278
rect 6334 10244 6368 10278
rect 6402 10244 6436 10278
rect 6470 10244 6504 10278
rect 6538 10244 6572 10278
rect 6606 10244 6640 10278
rect 6674 10244 6708 10278
rect 6742 10244 6776 10278
rect 6810 10244 6844 10278
rect 6878 10244 6912 10278
rect 6946 10244 6980 10278
rect 7014 10244 7048 10278
rect 7082 10244 7116 10278
rect 7150 10244 7184 10278
rect 7218 10244 7252 10278
rect 7286 10244 7320 10278
rect 7354 10244 7388 10278
rect 7422 10244 7456 10278
rect 7490 10244 7524 10278
rect 7558 10244 7592 10278
rect 7626 10244 7660 10278
rect 7694 10244 7728 10278
rect 7762 10244 7796 10278
rect 7830 10244 7864 10278
rect 7898 10244 7932 10278
rect 7966 10244 8000 10278
rect 8034 10244 8068 10278
rect 8102 10244 8136 10278
rect 8170 10244 8204 10278
rect 8238 10244 8272 10278
rect 8306 10244 8340 10278
rect 8374 10244 8408 10278
rect 8442 10244 8476 10278
rect 8510 10244 8544 10278
rect 8578 10244 8612 10278
rect 8646 10244 8680 10278
rect 8714 10244 8748 10278
rect 8782 10244 8816 10278
rect 8850 10244 8884 10278
rect 8918 10244 8952 10278
rect 8986 10244 9020 10278
rect 9054 10244 9088 10278
rect 9122 10244 9156 10278
rect 9190 10244 9224 10278
rect 9258 10244 9292 10278
rect 9326 10244 9360 10278
rect 9394 10244 9428 10278
rect 9462 10244 9496 10278
rect 9530 10244 9564 10278
rect 9598 10244 9632 10278
rect 9666 10244 9700 10278
rect 9734 10244 9768 10278
rect 9802 10244 9836 10278
rect 9870 10244 9904 10278
rect 9938 10244 9972 10278
rect 10006 10244 10040 10278
rect 10074 10244 10108 10278
rect 10142 10244 10176 10278
rect 10210 10244 10244 10278
rect 10278 10244 10312 10278
rect 10346 10244 10380 10278
rect 10414 10244 10448 10278
rect 10482 10244 10516 10278
rect 10550 10244 10584 10278
rect 10618 10244 10652 10278
rect 10686 10244 10720 10278
rect 10754 10244 10788 10278
rect 10822 10244 10856 10278
rect 10890 10244 10924 10278
rect 10958 10244 10992 10278
rect 11026 10244 11060 10278
rect 11094 10244 11128 10278
rect 11162 10244 11196 10278
rect 11230 10244 11264 10278
rect 11298 10244 11332 10278
rect 11366 10244 11400 10278
rect 11434 10244 11468 10278
rect 11502 10244 11536 10278
rect 11570 10244 11604 10278
rect 11638 10244 11672 10278
rect 11706 10244 11740 10278
rect 11774 10244 11808 10278
rect 11842 10244 11876 10278
rect 11910 10244 11944 10278
rect 11978 10244 12012 10278
rect 12046 10244 12080 10278
rect 12114 10244 12148 10278
rect 12182 10244 12216 10278
rect 12250 10244 12284 10278
rect 12318 10244 12352 10278
rect 12386 10244 12420 10278
rect 12454 10244 12488 10278
rect 12522 10244 12556 10278
rect 12590 10244 12624 10278
rect 12658 10244 12692 10278
rect 12726 10244 12760 10278
rect 12794 10244 12828 10278
rect 12862 10244 12896 10278
rect 12930 10244 12964 10278
rect 12998 10244 13032 10278
rect 13066 10244 13100 10278
rect 13134 10244 13168 10278
rect 13202 10244 13236 10278
rect 13270 10244 13304 10278
rect 13338 10244 13372 10278
rect 13406 10244 13440 10278
rect 13474 10244 13508 10278
rect 13542 10244 13576 10278
rect 13610 10244 13644 10278
rect 13678 10244 13712 10278
rect 14607 36174 14641 36208
rect 14607 36106 14641 36140
rect 14607 36038 14641 36072
rect 14607 35970 14641 36004
rect 14607 35902 14641 35936
rect 14607 35834 14641 35868
rect 14607 35766 14641 35800
rect 14607 35698 14641 35732
rect 14607 35630 14641 35664
rect 14607 35562 14641 35596
rect 14607 35494 14641 35528
rect 14607 35426 14641 35460
rect 14607 35358 14641 35392
rect 14607 35290 14641 35324
rect 14607 35222 14641 35256
rect 14607 35154 14641 35188
rect 14607 35086 14641 35120
rect 14607 35018 14641 35052
rect 14607 34950 14641 34984
rect 14607 34882 14641 34916
rect 14607 34814 14641 34848
rect 14607 34746 14641 34780
rect 14607 34678 14641 34712
rect 14607 34610 14641 34644
rect 14607 34542 14641 34576
rect 14607 34474 14641 34508
rect 14607 34406 14641 34440
rect 14607 34338 14641 34372
rect 14607 34270 14641 34304
rect 14607 34202 14641 34236
rect 14607 34134 14641 34168
rect 14607 34066 14641 34100
rect 14607 33998 14641 34032
rect 14607 33930 14641 33964
rect 14607 33862 14641 33896
rect 14607 33794 14641 33828
rect 14607 33726 14641 33760
rect 14607 33658 14641 33692
rect 14607 33590 14641 33624
rect 14607 33522 14641 33556
rect 14607 33454 14641 33488
rect 14607 33386 14641 33420
rect 14607 33318 14641 33352
rect 14607 33250 14641 33284
rect 14607 33182 14641 33216
rect 14607 33114 14641 33148
rect 14607 33046 14641 33080
rect 14607 32978 14641 33012
rect 14607 32910 14641 32944
rect 14607 32842 14641 32876
rect 14607 32774 14641 32808
rect 14607 32706 14641 32740
rect 14607 32638 14641 32672
rect 14607 32570 14641 32604
rect 14607 32502 14641 32536
rect 14607 32434 14641 32468
rect 14607 32366 14641 32400
rect 14607 32298 14641 32332
rect 14607 32230 14641 32264
rect 14607 32162 14641 32196
rect 14607 32094 14641 32128
rect 14607 32026 14641 32060
rect 14607 31958 14641 31992
rect 14607 31890 14641 31924
rect 14607 31822 14641 31856
rect 14607 31754 14641 31788
rect 14607 31686 14641 31720
rect 14607 31618 14641 31652
rect 14607 31550 14641 31584
rect 14607 31482 14641 31516
rect 14607 31414 14641 31448
rect 14607 31346 14641 31380
rect 14607 31278 14641 31312
rect 14607 31210 14641 31244
rect 14607 31142 14641 31176
rect 14607 31074 14641 31108
rect 14607 31006 14641 31040
rect 14607 30938 14641 30972
rect 14607 30870 14641 30904
rect 14607 30802 14641 30836
rect 14607 30734 14641 30768
rect 14607 30666 14641 30700
rect 14607 30598 14641 30632
rect 14607 30530 14641 30564
rect 14607 30462 14641 30496
rect 14607 30394 14641 30428
rect 14607 30326 14641 30360
rect 14607 30258 14641 30292
rect 14607 30190 14641 30224
rect 14607 30122 14641 30156
rect 14607 30054 14641 30088
rect 14607 29986 14641 30020
rect 14607 29918 14641 29952
rect 14607 29850 14641 29884
rect 14607 29782 14641 29816
rect 14607 29714 14641 29748
rect 14607 29646 14641 29680
rect 14607 29578 14641 29612
rect 14607 29510 14641 29544
rect 14607 29442 14641 29476
rect 14607 29374 14641 29408
rect 14607 29306 14641 29340
rect 14607 29238 14641 29272
rect 14607 29170 14641 29204
rect 14607 29102 14641 29136
rect 14607 29034 14641 29068
rect 14607 28966 14641 29000
rect 14607 28898 14641 28932
rect 14607 28830 14641 28864
rect 14607 28762 14641 28796
rect 14607 28694 14641 28728
rect 14607 28626 14641 28660
rect 14607 28558 14641 28592
rect 14607 28490 14641 28524
rect 14607 28422 14641 28456
rect 14607 28354 14641 28388
rect 14607 28286 14641 28320
rect 14607 28218 14641 28252
rect 14607 28150 14641 28184
rect 14607 28082 14641 28116
rect 14607 28014 14641 28048
rect 14607 27946 14641 27980
rect 14607 27878 14641 27912
rect 14607 27810 14641 27844
rect 14607 27742 14641 27776
rect 14607 27674 14641 27708
rect 14607 27606 14641 27640
rect 14607 27538 14641 27572
rect 14607 27470 14641 27504
rect 14607 27402 14641 27436
rect 14607 27334 14641 27368
rect 14607 27266 14641 27300
rect 14607 27198 14641 27232
rect 14607 27130 14641 27164
rect 14607 27062 14641 27096
rect 14607 26994 14641 27028
rect 14607 26926 14641 26960
rect 14607 26858 14641 26892
rect 14607 26790 14641 26824
rect 14607 26722 14641 26756
rect 14607 26654 14641 26688
rect 14607 26586 14641 26620
rect 14607 26518 14641 26552
rect 14607 26450 14641 26484
rect 14607 26382 14641 26416
rect 14607 26314 14641 26348
rect 14607 26246 14641 26280
rect 14607 26178 14641 26212
rect 14607 26110 14641 26144
rect 14607 26042 14641 26076
rect 14607 25974 14641 26008
rect 14607 25906 14641 25940
rect 14607 25838 14641 25872
rect 14607 25770 14641 25804
rect 14607 25702 14641 25736
rect 14607 25634 14641 25668
rect 14607 25566 14641 25600
rect 14607 25498 14641 25532
rect 14607 25430 14641 25464
rect 14607 25362 14641 25396
rect 14607 25294 14641 25328
rect 14607 25226 14641 25260
rect 14607 25158 14641 25192
rect 14607 25090 14641 25124
rect 14607 25022 14641 25056
rect 14607 24954 14641 24988
rect 14607 24886 14641 24920
rect 14607 24818 14641 24852
rect 14607 24750 14641 24784
rect 14607 24682 14641 24716
rect 14607 24614 14641 24648
rect 14607 24546 14641 24580
rect 14607 24478 14641 24512
rect 14607 24410 14641 24444
rect 14607 24342 14641 24376
rect 14607 24274 14641 24308
rect 14607 24206 14641 24240
rect 14607 24138 14641 24172
rect 14607 24070 14641 24104
rect 14607 24002 14641 24036
rect 14607 23934 14641 23968
rect 14607 23866 14641 23900
rect 14607 23798 14641 23832
rect 14607 23730 14641 23764
rect 14607 23662 14641 23696
rect 14607 23594 14641 23628
rect 14607 23526 14641 23560
rect 14607 23458 14641 23492
rect 14607 23390 14641 23424
rect 14607 23322 14641 23356
rect 14607 23254 14641 23288
rect 14607 23186 14641 23220
rect 14607 23118 14641 23152
rect 14607 23050 14641 23084
rect 14607 22982 14641 23016
rect 14607 22914 14641 22948
rect 14607 22846 14641 22880
rect 14607 22778 14641 22812
rect 14607 22710 14641 22744
rect 14607 22642 14641 22676
rect 14607 22574 14641 22608
rect 14607 22506 14641 22540
rect 14607 22438 14641 22472
rect 14607 22370 14641 22404
rect 14607 22302 14641 22336
rect 14607 22234 14641 22268
rect 14607 22166 14641 22200
rect 14607 22098 14641 22132
rect 14607 22030 14641 22064
rect 14607 21962 14641 21996
rect 14607 21894 14641 21928
rect 14607 21826 14641 21860
rect 14607 21758 14641 21792
rect 14607 21690 14641 21724
rect 14607 21622 14641 21656
rect 14607 21554 14641 21588
rect 14607 21486 14641 21520
rect 14607 21418 14641 21452
rect 14607 21350 14641 21384
rect 14607 21282 14641 21316
rect 14607 21214 14641 21248
rect 14607 21146 14641 21180
rect 14607 21078 14641 21112
rect 14607 21010 14641 21044
rect 14607 20942 14641 20976
rect 14607 20874 14641 20908
rect 14607 20806 14641 20840
rect 14607 20738 14641 20772
rect 14607 20670 14641 20704
rect 14607 20602 14641 20636
rect 14607 20534 14641 20568
rect 14607 20466 14641 20500
rect 14607 20398 14641 20432
rect 14607 20330 14641 20364
rect 14607 20262 14641 20296
rect 14607 20194 14641 20228
rect 14607 20126 14641 20160
rect 14607 20058 14641 20092
rect 14607 19990 14641 20024
rect 14607 19922 14641 19956
rect 14607 19854 14641 19888
rect 14607 19786 14641 19820
rect 14607 19718 14641 19752
rect 14607 19650 14641 19684
rect 14607 19582 14641 19616
rect 14607 19514 14641 19548
rect 14607 19446 14641 19480
rect 14607 19378 14641 19412
rect 14607 19310 14641 19344
rect 14607 19242 14641 19276
rect 14607 19174 14641 19208
rect 14607 19106 14641 19140
rect 14607 19038 14641 19072
rect 14607 18970 14641 19004
rect 14607 18902 14641 18936
rect 14607 18834 14641 18868
rect 14607 18766 14641 18800
rect 14607 18698 14641 18732
rect 14607 18630 14641 18664
rect 14607 18562 14641 18596
rect 14607 18494 14641 18528
rect 14607 18426 14641 18460
rect 14607 18358 14641 18392
rect 14607 18290 14641 18324
rect 14607 18222 14641 18256
rect 14607 18154 14641 18188
rect 14607 18086 14641 18120
rect 14607 18018 14641 18052
rect 14607 17950 14641 17984
rect 14607 17882 14641 17916
rect 14607 17814 14641 17848
rect 14607 17746 14641 17780
rect 14607 17678 14641 17712
rect 14607 17610 14641 17644
rect 14607 17542 14641 17576
rect 14607 17474 14641 17508
rect 14607 17406 14641 17440
rect 14607 17338 14641 17372
rect 14607 17270 14641 17304
rect 14607 17202 14641 17236
rect 14607 17134 14641 17168
rect 14607 17066 14641 17100
rect 14607 16998 14641 17032
rect 14607 16930 14641 16964
rect 14607 16862 14641 16896
rect 14607 16794 14641 16828
rect 14607 16726 14641 16760
rect 14607 16658 14641 16692
rect 14607 16590 14641 16624
rect 14607 16522 14641 16556
rect 14607 16454 14641 16488
rect 14607 16386 14641 16420
rect 14607 16318 14641 16352
rect 14607 16250 14641 16284
rect 14607 16182 14641 16216
rect 14607 16114 14641 16148
rect 14607 16046 14641 16080
rect 14607 15978 14641 16012
rect 14607 15910 14641 15944
rect 14607 15842 14641 15876
rect 14607 15774 14641 15808
rect 14607 15706 14641 15740
rect 14607 15638 14641 15672
rect 14607 15570 14641 15604
rect 14607 15502 14641 15536
rect 14607 15434 14641 15468
rect 14607 15366 14641 15400
rect 14607 15298 14641 15332
rect 14607 15230 14641 15264
rect 14607 15162 14641 15196
rect 14607 15094 14641 15128
rect 14607 15026 14641 15060
rect 14607 14958 14641 14992
rect 14607 14890 14641 14924
rect 14607 14822 14641 14856
rect 14607 14754 14641 14788
rect 14607 14686 14641 14720
rect 14607 14618 14641 14652
rect 14607 14550 14641 14584
rect 14607 14482 14641 14516
rect 14607 14414 14641 14448
rect 14607 14346 14641 14380
rect 14607 14278 14641 14312
rect 14607 14210 14641 14244
rect 14607 14142 14641 14176
rect 14607 14074 14641 14108
rect 14607 14006 14641 14040
rect 14607 13938 14641 13972
rect 14607 13870 14641 13904
rect 14607 13802 14641 13836
rect 14607 13734 14641 13768
rect 14607 13666 14641 13700
rect 14607 13598 14641 13632
rect 14607 13530 14641 13564
rect 14607 13462 14641 13496
rect 14607 13394 14641 13428
rect 14607 13326 14641 13360
rect 14607 13258 14641 13292
rect 14607 13190 14641 13224
rect 14607 13122 14641 13156
rect 14607 13054 14641 13088
rect 14607 12986 14641 13020
rect 14607 12918 14641 12952
rect 14607 12850 14641 12884
rect 14607 12782 14641 12816
rect 14607 12714 14641 12748
rect 14607 12646 14641 12680
rect 14607 12578 14641 12612
rect 14607 12510 14641 12544
rect 14607 12442 14641 12476
rect 14607 12374 14641 12408
rect 14607 12306 14641 12340
rect 14607 12238 14641 12272
rect 14607 12170 14641 12204
rect 14607 12102 14641 12136
rect 14607 12034 14641 12068
rect 14607 11966 14641 12000
rect 14607 11898 14641 11932
rect 14607 11830 14641 11864
rect 14607 11762 14641 11796
rect 14607 11694 14641 11728
rect 14607 11626 14641 11660
rect 14607 11558 14641 11592
rect 14607 11490 14641 11524
rect 14607 11422 14641 11456
rect 14607 11354 14641 11388
rect 14607 11286 14641 11320
rect 14607 11218 14641 11252
rect 14607 11150 14641 11184
rect 14607 11082 14641 11116
rect 14607 11014 14641 11048
rect 14607 10946 14641 10980
rect 14607 10878 14641 10912
rect 14607 10810 14641 10844
rect 14607 10742 14641 10776
rect 14607 10674 14641 10708
rect 14607 10606 14641 10640
rect 14607 10538 14641 10572
rect 14607 10470 14641 10504
rect 14607 10402 14641 10436
rect 14607 10334 14641 10368
rect 14607 10266 14641 10300
rect 14607 10198 14641 10232
rect 14607 10130 14641 10164
rect 14607 10062 14641 10096
rect 14607 9994 14641 10028
rect 14607 9926 14641 9960
rect 14607 9858 14641 9892
rect 14607 9790 14641 9824
rect 14607 9722 14641 9756
rect 312 9648 346 9682
rect 312 9580 346 9614
rect 14607 9654 14641 9688
rect 14607 9586 14641 9620
rect 476 9417 510 9451
rect 544 9417 578 9451
rect 612 9417 646 9451
rect 680 9417 714 9451
rect 748 9417 782 9451
rect 816 9417 850 9451
rect 884 9417 918 9451
rect 952 9417 986 9451
rect 1020 9417 1054 9451
rect 1088 9417 1122 9451
rect 1156 9417 1190 9451
rect 1224 9417 1258 9451
rect 1292 9417 1326 9451
rect 1360 9417 1394 9451
rect 1428 9417 1462 9451
rect 1496 9417 1530 9451
rect 1564 9417 1598 9451
rect 1632 9417 1666 9451
rect 1700 9417 1734 9451
rect 1768 9417 1802 9451
rect 1836 9417 1870 9451
rect 1904 9417 1938 9451
rect 1972 9417 2006 9451
rect 2040 9417 2074 9451
rect 2108 9417 2142 9451
rect 2176 9417 2210 9451
rect 2244 9417 2278 9451
rect 2312 9417 2346 9451
rect 2380 9417 2414 9451
rect 2448 9417 2482 9451
rect 2516 9417 2550 9451
rect 2584 9417 2618 9451
rect 2652 9417 2686 9451
rect 2720 9417 2754 9451
rect 2788 9417 2822 9451
rect 2856 9417 2890 9451
rect 2924 9417 2958 9451
rect 2992 9417 3026 9451
rect 3060 9417 3094 9451
rect 3128 9417 3162 9451
rect 3196 9417 3230 9451
rect 3264 9417 3298 9451
rect 3332 9417 3366 9451
rect 3400 9417 3434 9451
rect 3468 9417 3502 9451
rect 3536 9417 3570 9451
rect 3604 9417 3638 9451
rect 3672 9417 3706 9451
rect 3740 9417 3774 9451
rect 3808 9417 3842 9451
rect 3876 9417 3910 9451
rect 3944 9417 3978 9451
rect 4012 9417 4046 9451
rect 4080 9417 4114 9451
rect 4148 9417 4182 9451
rect 4216 9417 4250 9451
rect 4284 9417 4318 9451
rect 4352 9417 4386 9451
rect 4420 9417 4454 9451
rect 4488 9417 4522 9451
rect 4556 9417 4590 9451
rect 4624 9417 4658 9451
rect 4692 9417 4726 9451
rect 4760 9417 4794 9451
rect 4828 9417 4862 9451
rect 4896 9417 4930 9451
rect 4964 9417 4998 9451
rect 5032 9417 5066 9451
rect 5100 9417 5134 9451
rect 5168 9417 5202 9451
rect 5236 9417 5270 9451
rect 5304 9417 5338 9451
rect 5372 9417 5406 9451
rect 5440 9417 5474 9451
rect 5508 9417 5542 9451
rect 5576 9417 5610 9451
rect 5644 9417 5678 9451
rect 5712 9417 5746 9451
rect 5780 9417 5814 9451
rect 5848 9417 5882 9451
rect 5916 9417 5950 9451
rect 5984 9417 6018 9451
rect 6052 9417 6086 9451
rect 6120 9417 6154 9451
rect 6188 9417 6222 9451
rect 6256 9417 6290 9451
rect 6324 9417 6358 9451
rect 6392 9417 6426 9451
rect 6460 9417 6494 9451
rect 6528 9417 6562 9451
rect 6596 9417 6630 9451
rect 6664 9417 6698 9451
rect 6732 9417 6766 9451
rect 6800 9417 6834 9451
rect 6868 9417 6902 9451
rect 6936 9417 6970 9451
rect 7004 9417 7038 9451
rect 7072 9417 7106 9451
rect 7140 9417 7174 9451
rect 7208 9417 7242 9451
rect 7276 9417 7310 9451
rect 7344 9417 7378 9451
rect 7412 9417 7446 9451
rect 7480 9417 7514 9451
rect 7548 9417 7582 9451
rect 7616 9417 7650 9451
rect 7684 9417 7718 9451
rect 7752 9417 7786 9451
rect 7820 9417 7854 9451
rect 7888 9417 7922 9451
rect 7956 9417 7990 9451
rect 8024 9417 8058 9451
rect 8092 9417 8126 9451
rect 8160 9417 8194 9451
rect 8228 9417 8262 9451
rect 8296 9417 8330 9451
rect 8364 9417 8398 9451
rect 8432 9417 8466 9451
rect 8500 9417 8534 9451
rect 8568 9417 8602 9451
rect 8636 9417 8670 9451
rect 8704 9417 8738 9451
rect 8772 9417 8806 9451
rect 8840 9417 8874 9451
rect 8908 9417 8942 9451
rect 8976 9417 9010 9451
rect 9044 9417 9078 9451
rect 9112 9417 9146 9451
rect 9180 9417 9214 9451
rect 9248 9417 9282 9451
rect 9316 9417 9350 9451
rect 9384 9417 9418 9451
rect 9452 9417 9486 9451
rect 9520 9417 9554 9451
rect 9588 9417 9622 9451
rect 9656 9417 9690 9451
rect 9724 9417 9758 9451
rect 9792 9417 9826 9451
rect 9860 9417 9894 9451
rect 9928 9417 9962 9451
rect 9996 9417 10030 9451
rect 10064 9417 10098 9451
rect 10132 9417 10166 9451
rect 10200 9417 10234 9451
rect 10268 9417 10302 9451
rect 10336 9417 10370 9451
rect 10404 9417 10438 9451
rect 10472 9417 10506 9451
rect 10540 9417 10574 9451
rect 10608 9417 10642 9451
rect 10676 9417 10710 9451
rect 10744 9417 10778 9451
rect 10812 9417 10846 9451
rect 10880 9417 10914 9451
rect 10948 9417 10982 9451
rect 11016 9417 11050 9451
rect 11084 9417 11118 9451
rect 11152 9417 11186 9451
rect 11220 9417 11254 9451
rect 11288 9417 11322 9451
rect 11356 9417 11390 9451
rect 11424 9417 11458 9451
rect 11492 9417 11526 9451
rect 11560 9417 11594 9451
rect 11628 9417 11662 9451
rect 11696 9417 11730 9451
rect 11764 9417 11798 9451
rect 11832 9417 11866 9451
rect 11900 9417 11934 9451
rect 11968 9417 12002 9451
rect 12036 9417 12070 9451
rect 12104 9417 12138 9451
rect 12172 9417 12206 9451
rect 12240 9417 12274 9451
rect 12308 9417 12342 9451
rect 12376 9417 12410 9451
rect 12444 9417 12478 9451
rect 12512 9417 12546 9451
rect 12580 9417 12614 9451
rect 12648 9417 12682 9451
rect 12716 9417 12750 9451
rect 12784 9417 12818 9451
rect 12852 9417 12886 9451
rect 12920 9417 12954 9451
rect 12988 9417 13022 9451
rect 13056 9417 13090 9451
rect 13124 9417 13158 9451
rect 13192 9417 13226 9451
rect 13260 9417 13294 9451
rect 13328 9417 13362 9451
rect 13396 9417 13430 9451
rect 13464 9417 13498 9451
rect 13532 9417 13566 9451
rect 13600 9417 13634 9451
rect 13668 9417 13702 9451
rect 13736 9417 13770 9451
rect 13804 9417 13838 9451
rect 13872 9417 13906 9451
rect 13940 9417 13974 9451
rect 14008 9417 14042 9451
rect 14076 9417 14110 9451
rect 14144 9417 14178 9451
rect 14212 9417 14246 9451
rect 14280 9417 14314 9451
rect 14348 9417 14382 9451
rect 14416 9417 14450 9451
rect 14484 9417 14518 9451
<< mvnsubdiffcont >>
rect 766 36143 800 36177
rect 834 36143 868 36177
rect 902 36143 936 36177
rect 970 36143 1004 36177
rect 1038 36143 1072 36177
rect 1106 36143 1140 36177
rect 1174 36143 1208 36177
rect 1242 36143 1276 36177
rect 1310 36143 1344 36177
rect 1378 36143 1412 36177
rect 1446 36143 1480 36177
rect 1514 36143 1548 36177
rect 1582 36143 1616 36177
rect 1650 36143 1684 36177
rect 1718 36143 1752 36177
rect 1786 36143 1820 36177
rect 1854 36143 1888 36177
rect 1922 36143 1956 36177
rect 1990 36143 2024 36177
rect 2058 36143 2092 36177
rect 2126 36143 2160 36177
rect 2194 36143 2228 36177
rect 2262 36143 2296 36177
rect 2330 36143 2364 36177
rect 2398 36143 2432 36177
rect 2466 36143 2500 36177
rect 2534 36143 2568 36177
rect 2602 36143 2636 36177
rect 2670 36143 2704 36177
rect 2738 36143 2772 36177
rect 2806 36143 2840 36177
rect 2874 36143 2908 36177
rect 2942 36143 2976 36177
rect 3010 36143 3044 36177
rect 3078 36143 3112 36177
rect 3146 36143 3180 36177
rect 3214 36143 3248 36177
rect 3282 36143 3316 36177
rect 3350 36143 3384 36177
rect 3418 36143 3452 36177
rect 3486 36143 3520 36177
rect 3554 36143 3588 36177
rect 3622 36143 3656 36177
rect 3690 36143 3724 36177
rect 3758 36143 3792 36177
rect 3826 36143 3860 36177
rect 3894 36143 3928 36177
rect 3962 36143 3996 36177
rect 4030 36143 4064 36177
rect 4098 36143 4132 36177
rect 4166 36143 4200 36177
rect 4234 36143 4268 36177
rect 4302 36143 4336 36177
rect 4370 36143 4404 36177
rect 4438 36143 4472 36177
rect 4506 36143 4540 36177
rect 4574 36143 4608 36177
rect 4642 36143 4676 36177
rect 4710 36143 4744 36177
rect 4778 36143 4812 36177
rect 4846 36143 4880 36177
rect 4914 36143 4948 36177
rect 4982 36143 5016 36177
rect 5050 36143 5084 36177
rect 5118 36143 5152 36177
rect 5186 36143 5220 36177
rect 5254 36143 5288 36177
rect 5322 36143 5356 36177
rect 5390 36143 5424 36177
rect 5458 36143 5492 36177
rect 5526 36143 5560 36177
rect 5594 36143 5628 36177
rect 5662 36143 5696 36177
rect 5730 36143 5764 36177
rect 5798 36143 5832 36177
rect 5866 36143 5900 36177
rect 5934 36143 5968 36177
rect 6002 36143 6036 36177
rect 6070 36143 6104 36177
rect 6138 36143 6172 36177
rect 6206 36143 6240 36177
rect 6274 36143 6308 36177
rect 6342 36143 6376 36177
rect 6410 36143 6444 36177
rect 6478 36143 6512 36177
rect 6546 36143 6580 36177
rect 6614 36143 6648 36177
rect 6682 36143 6716 36177
rect 6750 36143 6784 36177
rect 6818 36143 6852 36177
rect 6886 36143 6920 36177
rect 6954 36143 6988 36177
rect 7022 36143 7056 36177
rect 7090 36143 7124 36177
rect 7158 36143 7192 36177
rect 7226 36143 7260 36177
rect 7294 36143 7328 36177
rect 7362 36143 7396 36177
rect 7430 36143 7464 36177
rect 7498 36143 7532 36177
rect 7566 36143 7600 36177
rect 7634 36143 7668 36177
rect 7702 36143 7736 36177
rect 7770 36143 7804 36177
rect 7838 36143 7872 36177
rect 7906 36143 7940 36177
rect 7974 36143 8008 36177
rect 8042 36143 8076 36177
rect 8110 36143 8144 36177
rect 8178 36143 8212 36177
rect 8246 36143 8280 36177
rect 8314 36143 8348 36177
rect 8382 36143 8416 36177
rect 8450 36143 8484 36177
rect 8518 36143 8552 36177
rect 8586 36143 8620 36177
rect 8654 36143 8688 36177
rect 8722 36143 8756 36177
rect 8790 36143 8824 36177
rect 8858 36143 8892 36177
rect 8926 36143 8960 36177
rect 8994 36143 9028 36177
rect 9062 36143 9096 36177
rect 9130 36143 9164 36177
rect 9198 36143 9232 36177
rect 9266 36143 9300 36177
rect 9334 36143 9368 36177
rect 9402 36143 9436 36177
rect 9470 36143 9504 36177
rect 9538 36143 9572 36177
rect 9606 36143 9640 36177
rect 9674 36143 9708 36177
rect 9742 36143 9776 36177
rect 9810 36143 9844 36177
rect 9878 36143 9912 36177
rect 9946 36143 9980 36177
rect 10014 36143 10048 36177
rect 10082 36143 10116 36177
rect 10150 36143 10184 36177
rect 10218 36143 10252 36177
rect 10286 36143 10320 36177
rect 10354 36143 10388 36177
rect 10422 36143 10456 36177
rect 10490 36143 10524 36177
rect 10558 36143 10592 36177
rect 10626 36143 10660 36177
rect 10694 36143 10728 36177
rect 10762 36143 10796 36177
rect 10830 36143 10864 36177
rect 10898 36143 10932 36177
rect 10966 36143 11000 36177
rect 11034 36143 11068 36177
rect 11102 36143 11136 36177
rect 11170 36143 11204 36177
rect 11238 36143 11272 36177
rect 11306 36143 11340 36177
rect 11374 36143 11408 36177
rect 11442 36143 11476 36177
rect 11510 36143 11544 36177
rect 11578 36143 11612 36177
rect 11646 36143 11680 36177
rect 11714 36143 11748 36177
rect 11782 36143 11816 36177
rect 11850 36143 11884 36177
rect 11918 36143 11952 36177
rect 11986 36143 12020 36177
rect 12054 36143 12088 36177
rect 12122 36143 12156 36177
rect 12190 36143 12224 36177
rect 12258 36143 12292 36177
rect 12326 36143 12360 36177
rect 12394 36143 12428 36177
rect 12462 36143 12496 36177
rect 12530 36143 12564 36177
rect 12598 36143 12632 36177
rect 12666 36143 12700 36177
rect 12734 36143 12768 36177
rect 12802 36143 12836 36177
rect 12870 36143 12904 36177
rect 12938 36143 12972 36177
rect 13006 36143 13040 36177
rect 13074 36143 13108 36177
rect 13142 36143 13176 36177
rect 13210 36143 13244 36177
rect 13278 36143 13312 36177
rect 13346 36143 13380 36177
rect 13414 36143 13448 36177
rect 13482 36143 13516 36177
rect 13550 36143 13584 36177
rect 13618 36143 13652 36177
rect 13686 36143 13720 36177
rect 13754 36143 13788 36177
rect 13822 36143 13856 36177
rect 13890 36143 13924 36177
rect 13958 36143 13992 36177
rect 14026 36143 14060 36177
rect 14094 36143 14128 36177
rect 14162 36143 14196 36177
rect 632 35998 666 36032
rect 632 35930 666 35964
rect 632 35862 666 35896
rect 632 35794 666 35828
rect 632 35726 666 35760
rect 632 35658 666 35692
rect 632 35590 666 35624
rect 632 35522 666 35556
rect 632 35454 666 35488
rect 632 35386 666 35420
rect 632 35318 666 35352
rect 632 35250 666 35284
rect 632 35182 666 35216
rect 632 35114 666 35148
rect 632 35046 666 35080
rect 632 34978 666 35012
rect 632 34910 666 34944
rect 632 34842 666 34876
rect 632 34774 666 34808
rect 632 34706 666 34740
rect 14297 35998 14331 36032
rect 14297 35930 14331 35964
rect 14297 35862 14331 35896
rect 14297 35794 14331 35828
rect 14297 35726 14331 35760
rect 14297 35658 14331 35692
rect 14297 35590 14331 35624
rect 14297 35522 14331 35556
rect 14297 35454 14331 35488
rect 14297 35386 14331 35420
rect 14297 35318 14331 35352
rect 14297 35250 14331 35284
rect 14297 35182 14331 35216
rect 14297 35114 14331 35148
rect 14297 35046 14331 35080
rect 14297 34978 14331 35012
rect 14297 34910 14331 34944
rect 14297 34842 14331 34876
rect 14297 34774 14331 34808
rect 632 34638 666 34672
rect 632 34570 666 34604
rect 632 34502 666 34536
rect 632 34434 666 34468
rect 632 34366 666 34400
rect 632 34298 666 34332
rect 632 34230 666 34264
rect 632 34162 666 34196
rect 632 34094 666 34128
rect 632 34026 666 34060
rect 632 33958 666 33992
rect 632 33890 666 33924
rect 632 33822 666 33856
rect 632 33754 666 33788
rect 632 33686 666 33720
rect 632 33618 666 33652
rect 632 33550 666 33584
rect 632 33482 666 33516
rect 632 33414 666 33448
rect 632 33346 666 33380
rect 632 33278 666 33312
rect 632 33210 666 33244
rect 632 33142 666 33176
rect 632 33074 666 33108
rect 632 33006 666 33040
rect 632 32938 666 32972
rect 632 32870 666 32904
rect 632 32802 666 32836
rect 632 32734 666 32768
rect 632 32666 666 32700
rect 632 32598 666 32632
rect 632 32530 666 32564
rect 632 32462 666 32496
rect 632 32394 666 32428
rect 632 32326 666 32360
rect 632 32258 666 32292
rect 632 32190 666 32224
rect 632 32122 666 32156
rect 632 32054 666 32088
rect 632 31986 666 32020
rect 632 31918 666 31952
rect 632 31850 666 31884
rect 632 31782 666 31816
rect 632 31714 666 31748
rect 632 31646 666 31680
rect 632 31578 666 31612
rect 632 31510 666 31544
rect 632 31442 666 31476
rect 632 31374 666 31408
rect 632 31306 666 31340
rect 632 31238 666 31272
rect 632 31170 666 31204
rect 632 31102 666 31136
rect 632 31034 666 31068
rect 632 30966 666 31000
rect 632 30898 666 30932
rect 632 30830 666 30864
rect 632 30762 666 30796
rect 632 30694 666 30728
rect 632 30626 666 30660
rect 632 30558 666 30592
rect 632 30490 666 30524
rect 632 30422 666 30456
rect 632 30354 666 30388
rect 632 30286 666 30320
rect 632 30218 666 30252
rect 632 30150 666 30184
rect 632 30082 666 30116
rect 632 30014 666 30048
rect 632 29946 666 29980
rect 632 29878 666 29912
rect 632 29810 666 29844
rect 632 29742 666 29776
rect 632 29674 666 29708
rect 632 29606 666 29640
rect 632 29538 666 29572
rect 632 29470 666 29504
rect 632 29402 666 29436
rect 632 29334 666 29368
rect 632 29266 666 29300
rect 632 29198 666 29232
rect 632 29130 666 29164
rect 632 29062 666 29096
rect 632 28994 666 29028
rect 632 28926 666 28960
rect 632 28858 666 28892
rect 632 28790 666 28824
rect 632 28722 666 28756
rect 632 28654 666 28688
rect 632 28586 666 28620
rect 632 28518 666 28552
rect 632 28450 666 28484
rect 632 28382 666 28416
rect 632 28314 666 28348
rect 632 28246 666 28280
rect 632 28178 666 28212
rect 632 28110 666 28144
rect 632 28042 666 28076
rect 632 27974 666 28008
rect 632 27906 666 27940
rect 632 27838 666 27872
rect 632 27770 666 27804
rect 632 27702 666 27736
rect 632 27634 666 27668
rect 632 27566 666 27600
rect 632 27498 666 27532
rect 632 27430 666 27464
rect 632 27362 666 27396
rect 632 27294 666 27328
rect 632 27226 666 27260
rect 632 27158 666 27192
rect 632 27090 666 27124
rect 632 27022 666 27056
rect 632 26954 666 26988
rect 632 26886 666 26920
rect 632 26818 666 26852
rect 632 26750 666 26784
rect 632 26682 666 26716
rect 632 26614 666 26648
rect 632 26546 666 26580
rect 632 26478 666 26512
rect 632 26410 666 26444
rect 632 26342 666 26376
rect 632 26274 666 26308
rect 632 26206 666 26240
rect 632 26138 666 26172
rect 632 26070 666 26104
rect 632 26002 666 26036
rect 632 25934 666 25968
rect 632 25866 666 25900
rect 632 25798 666 25832
rect 632 25730 666 25764
rect 632 25662 666 25696
rect 632 25594 666 25628
rect 632 25526 666 25560
rect 632 25458 666 25492
rect 632 25390 666 25424
rect 632 25322 666 25356
rect 632 25254 666 25288
rect 632 25186 666 25220
rect 632 25118 666 25152
rect 632 25050 666 25084
rect 632 24982 666 25016
rect 632 24914 666 24948
rect 632 24846 666 24880
rect 632 24778 666 24812
rect 632 24710 666 24744
rect 632 24642 666 24676
rect 632 24574 666 24608
rect 632 24506 666 24540
rect 632 24438 666 24472
rect 632 24370 666 24404
rect 632 24302 666 24336
rect 632 24234 666 24268
rect 632 24166 666 24200
rect 632 24098 666 24132
rect 632 24030 666 24064
rect 632 23962 666 23996
rect 632 23894 666 23928
rect 632 23826 666 23860
rect 632 23758 666 23792
rect 632 23690 666 23724
rect 632 23622 666 23656
rect 632 23554 666 23588
rect 632 23486 666 23520
rect 632 23418 666 23452
rect 632 23350 666 23384
rect 632 23282 666 23316
rect 632 23214 666 23248
rect 632 23146 666 23180
rect 632 23078 666 23112
rect 632 23010 666 23044
rect 632 22942 666 22976
rect 632 22874 666 22908
rect 632 22806 666 22840
rect 632 22738 666 22772
rect 632 22670 666 22704
rect 632 22602 666 22636
rect 632 22534 666 22568
rect 632 22466 666 22500
rect 632 22398 666 22432
rect 632 22330 666 22364
rect 632 22262 666 22296
rect 632 22194 666 22228
rect 632 22126 666 22160
rect 632 22058 666 22092
rect 632 21990 666 22024
rect 632 21922 666 21956
rect 632 21854 666 21888
rect 632 21786 666 21820
rect 632 21718 666 21752
rect 632 21650 666 21684
rect 632 21582 666 21616
rect 632 21514 666 21548
rect 632 21446 666 21480
rect 632 21378 666 21412
rect 632 21310 666 21344
rect 632 21242 666 21276
rect 632 21174 666 21208
rect 632 21106 666 21140
rect 632 21038 666 21072
rect 632 20970 666 21004
rect 632 20902 666 20936
rect 632 20834 666 20868
rect 632 20766 666 20800
rect 632 20698 666 20732
rect 632 20630 666 20664
rect 632 20562 666 20596
rect 632 20494 666 20528
rect 632 20426 666 20460
rect 632 20358 666 20392
rect 632 20290 666 20324
rect 632 20222 666 20256
rect 632 20154 666 20188
rect 632 20086 666 20120
rect 632 20018 666 20052
rect 632 19950 666 19984
rect 632 19882 666 19916
rect 632 19814 666 19848
rect 632 19746 666 19780
rect 632 19678 666 19712
rect 632 19610 666 19644
rect 632 19542 666 19576
rect 632 19474 666 19508
rect 632 19406 666 19440
rect 632 19338 666 19372
rect 632 19270 666 19304
rect 632 19202 666 19236
rect 632 19134 666 19168
rect 632 19066 666 19100
rect 632 18998 666 19032
rect 632 18930 666 18964
rect 632 18862 666 18896
rect 632 18794 666 18828
rect 632 18726 666 18760
rect 632 18658 666 18692
rect 632 18590 666 18624
rect 632 18522 666 18556
rect 632 18454 666 18488
rect 632 18386 666 18420
rect 632 18318 666 18352
rect 632 18250 666 18284
rect 632 18182 666 18216
rect 632 18114 666 18148
rect 632 18046 666 18080
rect 632 17978 666 18012
rect 632 17910 666 17944
rect 632 17842 666 17876
rect 632 17774 666 17808
rect 632 17706 666 17740
rect 632 17638 666 17672
rect 632 17570 666 17604
rect 632 17502 666 17536
rect 632 17434 666 17468
rect 632 17366 666 17400
rect 632 17298 666 17332
rect 632 17230 666 17264
rect 632 17162 666 17196
rect 632 17094 666 17128
rect 632 17026 666 17060
rect 632 16958 666 16992
rect 632 16890 666 16924
rect 632 16822 666 16856
rect 632 16754 666 16788
rect 632 16686 666 16720
rect 632 16618 666 16652
rect 632 16550 666 16584
rect 632 16482 666 16516
rect 632 16414 666 16448
rect 632 16346 666 16380
rect 632 16278 666 16312
rect 632 16210 666 16244
rect 632 16142 666 16176
rect 632 16074 666 16108
rect 632 16006 666 16040
rect 632 15938 666 15972
rect 632 15870 666 15904
rect 632 15802 666 15836
rect 632 15734 666 15768
rect 632 15666 666 15700
rect 632 15598 666 15632
rect 632 15530 666 15564
rect 632 15462 666 15496
rect 632 15394 666 15428
rect 632 15326 666 15360
rect 632 15258 666 15292
rect 632 15190 666 15224
rect 632 15122 666 15156
rect 632 15054 666 15088
rect 632 14986 666 15020
rect 632 14918 666 14952
rect 632 14850 666 14884
rect 632 14782 666 14816
rect 632 14714 666 14748
rect 632 14646 666 14680
rect 632 14578 666 14612
rect 632 14510 666 14544
rect 632 14442 666 14476
rect 632 14374 666 14408
rect 632 14306 666 14340
rect 632 14238 666 14272
rect 632 14170 666 14204
rect 632 14102 666 14136
rect 632 14034 666 14068
rect 632 13966 666 14000
rect 632 13898 666 13932
rect 632 13830 666 13864
rect 632 13762 666 13796
rect 632 13694 666 13728
rect 632 13626 666 13660
rect 632 13558 666 13592
rect 632 13490 666 13524
rect 632 13422 666 13456
rect 632 13354 666 13388
rect 632 13286 666 13320
rect 632 13218 666 13252
rect 632 13150 666 13184
rect 632 13082 666 13116
rect 632 13014 666 13048
rect 632 12946 666 12980
rect 632 12878 666 12912
rect 632 12810 666 12844
rect 632 12742 666 12776
rect 632 12674 666 12708
rect 632 12606 666 12640
rect 632 12538 666 12572
rect 632 12470 666 12504
rect 632 12402 666 12436
rect 632 12334 666 12368
rect 632 12266 666 12300
rect 632 12198 666 12232
rect 632 12130 666 12164
rect 632 12062 666 12096
rect 632 11994 666 12028
rect 632 11926 666 11960
rect 632 11858 666 11892
rect 632 11790 666 11824
rect 632 11722 666 11756
rect 632 11654 666 11688
rect 632 11586 666 11620
rect 632 11518 666 11552
rect 632 11450 666 11484
rect 632 11382 666 11416
rect 632 11314 666 11348
rect 632 11246 666 11280
rect 632 11178 666 11212
rect 632 11110 666 11144
rect 632 11042 666 11076
rect 632 10974 666 11008
rect 632 10906 666 10940
rect 632 10838 666 10872
rect 632 10770 666 10804
rect 632 10702 666 10736
rect 632 10634 666 10668
rect 632 10566 666 10600
rect 632 10498 666 10532
rect 632 10430 666 10464
rect 632 10362 666 10396
rect 632 10294 666 10328
rect 632 10226 666 10260
rect 2119 28505 12897 28879
rect 1689 27504 2063 28422
rect 12953 27504 13327 28422
rect 2119 27047 12897 27421
rect 14297 34706 14331 34740
rect 14297 34638 14331 34672
rect 14297 34570 14331 34604
rect 14297 34502 14331 34536
rect 14297 34434 14331 34468
rect 14297 34366 14331 34400
rect 14297 34298 14331 34332
rect 14297 34230 14331 34264
rect 14297 34162 14331 34196
rect 14297 34094 14331 34128
rect 14297 34026 14331 34060
rect 14297 33958 14331 33992
rect 14297 33890 14331 33924
rect 14297 33822 14331 33856
rect 14297 33754 14331 33788
rect 14297 33686 14331 33720
rect 14297 33618 14331 33652
rect 14297 33550 14331 33584
rect 14297 33482 14331 33516
rect 14297 33414 14331 33448
rect 14297 33346 14331 33380
rect 14297 33278 14331 33312
rect 14297 33210 14331 33244
rect 14297 33142 14331 33176
rect 14297 33074 14331 33108
rect 14297 33006 14331 33040
rect 14297 32938 14331 32972
rect 14297 32870 14331 32904
rect 14297 32802 14331 32836
rect 14297 32734 14331 32768
rect 14297 32666 14331 32700
rect 14297 32598 14331 32632
rect 14297 32530 14331 32564
rect 14297 32462 14331 32496
rect 14297 32394 14331 32428
rect 14297 32326 14331 32360
rect 14297 32258 14331 32292
rect 14297 32190 14331 32224
rect 14297 32122 14331 32156
rect 14297 32054 14331 32088
rect 14297 31986 14331 32020
rect 14297 31918 14331 31952
rect 14297 31850 14331 31884
rect 14297 31782 14331 31816
rect 14297 31714 14331 31748
rect 14297 31646 14331 31680
rect 14297 31578 14331 31612
rect 14297 31510 14331 31544
rect 14297 31442 14331 31476
rect 14297 31374 14331 31408
rect 14297 31306 14331 31340
rect 14297 31238 14331 31272
rect 14297 31170 14331 31204
rect 14297 31102 14331 31136
rect 14297 31034 14331 31068
rect 14297 30966 14331 31000
rect 14297 30898 14331 30932
rect 14297 30830 14331 30864
rect 14297 30762 14331 30796
rect 14297 30694 14331 30728
rect 14297 30626 14331 30660
rect 14297 30558 14331 30592
rect 14297 30490 14331 30524
rect 14297 30422 14331 30456
rect 14297 30354 14331 30388
rect 14297 30286 14331 30320
rect 14297 30218 14331 30252
rect 14297 30150 14331 30184
rect 14297 30082 14331 30116
rect 14297 30014 14331 30048
rect 14297 29946 14331 29980
rect 14297 29878 14331 29912
rect 14297 29810 14331 29844
rect 14297 29742 14331 29776
rect 14297 29674 14331 29708
rect 14297 29606 14331 29640
rect 14297 29538 14331 29572
rect 14297 29470 14331 29504
rect 14297 29402 14331 29436
rect 14297 29334 14331 29368
rect 14297 29266 14331 29300
rect 14297 29198 14331 29232
rect 14297 29130 14331 29164
rect 14297 29062 14331 29096
rect 14297 28994 14331 29028
rect 14297 28926 14331 28960
rect 14297 28858 14331 28892
rect 14297 28790 14331 28824
rect 14297 28722 14331 28756
rect 14297 28654 14331 28688
rect 14297 28586 14331 28620
rect 14297 28518 14331 28552
rect 14297 28450 14331 28484
rect 14297 28382 14331 28416
rect 14297 28314 14331 28348
rect 14297 28246 14331 28280
rect 14297 28178 14331 28212
rect 14297 28110 14331 28144
rect 14297 28042 14331 28076
rect 14297 27974 14331 28008
rect 14297 27906 14331 27940
rect 14297 27838 14331 27872
rect 14297 27770 14331 27804
rect 14297 27702 14331 27736
rect 14297 27634 14331 27668
rect 14297 27566 14331 27600
rect 14297 27498 14331 27532
rect 14297 27430 14331 27464
rect 14297 27362 14331 27396
rect 14297 27294 14331 27328
rect 14297 27226 14331 27260
rect 14297 27158 14331 27192
rect 14297 27090 14331 27124
rect 14297 27022 14331 27056
rect 14297 26954 14331 26988
rect 14297 26886 14331 26920
rect 14297 26818 14331 26852
rect 14297 26750 14331 26784
rect 14297 26682 14331 26716
rect 14297 26614 14331 26648
rect 14297 26546 14331 26580
rect 14297 26478 14331 26512
rect 14297 26410 14331 26444
rect 14297 26342 14331 26376
rect 14297 26274 14331 26308
rect 14297 26206 14331 26240
rect 14297 26138 14331 26172
rect 14297 26070 14331 26104
rect 14297 26002 14331 26036
rect 14297 25934 14331 25968
rect 14297 25866 14331 25900
rect 14297 25798 14331 25832
rect 14297 25730 14331 25764
rect 14297 25662 14331 25696
rect 14297 25594 14331 25628
rect 14297 25526 14331 25560
rect 14297 25458 14331 25492
rect 14297 25390 14331 25424
rect 14297 25322 14331 25356
rect 14297 25254 14331 25288
rect 14297 25186 14331 25220
rect 14297 25118 14331 25152
rect 14297 25050 14331 25084
rect 14297 24982 14331 25016
rect 14297 24914 14331 24948
rect 14297 24846 14331 24880
rect 14297 24778 14331 24812
rect 14297 24710 14331 24744
rect 14297 24642 14331 24676
rect 14297 24574 14331 24608
rect 14297 24506 14331 24540
rect 14297 24438 14331 24472
rect 14297 24370 14331 24404
rect 14297 24302 14331 24336
rect 14297 24234 14331 24268
rect 14297 24166 14331 24200
rect 14297 24098 14331 24132
rect 14297 24030 14331 24064
rect 14297 23962 14331 23996
rect 14297 23894 14331 23928
rect 14297 23826 14331 23860
rect 14297 23758 14331 23792
rect 14297 23690 14331 23724
rect 14297 23622 14331 23656
rect 14297 23554 14331 23588
rect 14297 23486 14331 23520
rect 14297 23418 14331 23452
rect 14297 23350 14331 23384
rect 14297 23282 14331 23316
rect 14297 23214 14331 23248
rect 14297 23146 14331 23180
rect 14297 23078 14331 23112
rect 14297 23010 14331 23044
rect 14297 22942 14331 22976
rect 14297 22874 14331 22908
rect 14297 22806 14331 22840
rect 14297 22738 14331 22772
rect 14297 22670 14331 22704
rect 14297 22602 14331 22636
rect 14297 22534 14331 22568
rect 14297 22466 14331 22500
rect 14297 22398 14331 22432
rect 14297 22330 14331 22364
rect 14297 22262 14331 22296
rect 14297 22194 14331 22228
rect 14297 22126 14331 22160
rect 14297 22058 14331 22092
rect 14297 21990 14331 22024
rect 14297 21922 14331 21956
rect 14297 21854 14331 21888
rect 14297 21786 14331 21820
rect 14297 21718 14331 21752
rect 14297 21650 14331 21684
rect 14297 21582 14331 21616
rect 14297 21514 14331 21548
rect 14297 21446 14331 21480
rect 14297 21378 14331 21412
rect 14297 21310 14331 21344
rect 14297 21242 14331 21276
rect 14297 21174 14331 21208
rect 14297 21106 14331 21140
rect 14297 21038 14331 21072
rect 14297 20970 14331 21004
rect 14297 20902 14331 20936
rect 14297 20834 14331 20868
rect 14297 20766 14331 20800
rect 14297 20698 14331 20732
rect 14297 20630 14331 20664
rect 14297 20562 14331 20596
rect 14297 20494 14331 20528
rect 14297 20426 14331 20460
rect 14297 20358 14331 20392
rect 14297 20290 14331 20324
rect 14297 20222 14331 20256
rect 14297 20154 14331 20188
rect 14297 20086 14331 20120
rect 14297 20018 14331 20052
rect 14297 19950 14331 19984
rect 14297 19882 14331 19916
rect 14297 19814 14331 19848
rect 14297 19746 14331 19780
rect 14297 19678 14331 19712
rect 14297 19610 14331 19644
rect 14297 19542 14331 19576
rect 14297 19474 14331 19508
rect 14297 19406 14331 19440
rect 14297 19338 14331 19372
rect 14297 19270 14331 19304
rect 14297 19202 14331 19236
rect 14297 19134 14331 19168
rect 14297 19066 14331 19100
rect 14297 18998 14331 19032
rect 14297 18930 14331 18964
rect 14297 18862 14331 18896
rect 14297 18794 14331 18828
rect 14297 18726 14331 18760
rect 14297 18658 14331 18692
rect 14297 18590 14331 18624
rect 14297 18522 14331 18556
rect 14297 18454 14331 18488
rect 14297 18386 14331 18420
rect 14297 18318 14331 18352
rect 14297 18250 14331 18284
rect 14297 18182 14331 18216
rect 14297 18114 14331 18148
rect 14297 18046 14331 18080
rect 14297 17978 14331 18012
rect 14297 17910 14331 17944
rect 14297 17842 14331 17876
rect 14297 17774 14331 17808
rect 14297 17706 14331 17740
rect 14297 17638 14331 17672
rect 14297 17570 14331 17604
rect 14297 17502 14331 17536
rect 14297 17434 14331 17468
rect 14297 17366 14331 17400
rect 14297 17298 14331 17332
rect 14297 17230 14331 17264
rect 14297 17162 14331 17196
rect 14297 17094 14331 17128
rect 14297 17026 14331 17060
rect 14297 16958 14331 16992
rect 14297 16890 14331 16924
rect 14297 16822 14331 16856
rect 14297 16754 14331 16788
rect 14297 16686 14331 16720
rect 14297 16618 14331 16652
rect 14297 16550 14331 16584
rect 14297 16482 14331 16516
rect 14297 16414 14331 16448
rect 14297 16346 14331 16380
rect 14297 16278 14331 16312
rect 14297 16210 14331 16244
rect 14297 16142 14331 16176
rect 14297 16074 14331 16108
rect 14297 16006 14331 16040
rect 14297 15938 14331 15972
rect 14297 15870 14331 15904
rect 14297 15802 14331 15836
rect 14297 15734 14331 15768
rect 14297 15666 14331 15700
rect 14297 15598 14331 15632
rect 14297 15530 14331 15564
rect 14297 15462 14331 15496
rect 14297 15394 14331 15428
rect 14297 15326 14331 15360
rect 14297 15258 14331 15292
rect 14297 15190 14331 15224
rect 14297 15122 14331 15156
rect 14297 15054 14331 15088
rect 14297 14986 14331 15020
rect 14297 14918 14331 14952
rect 14297 14850 14331 14884
rect 14297 14782 14331 14816
rect 14297 14714 14331 14748
rect 14297 14646 14331 14680
rect 14297 14578 14331 14612
rect 14297 14510 14331 14544
rect 14297 14442 14331 14476
rect 14297 14374 14331 14408
rect 14297 14306 14331 14340
rect 14297 14238 14331 14272
rect 14297 14170 14331 14204
rect 14297 14102 14331 14136
rect 14297 14034 14331 14068
rect 14297 13966 14331 14000
rect 14297 13898 14331 13932
rect 14297 13830 14331 13864
rect 14297 13762 14331 13796
rect 14297 13694 14331 13728
rect 14297 13626 14331 13660
rect 14297 13558 14331 13592
rect 14297 13490 14331 13524
rect 14297 13422 14331 13456
rect 14297 13354 14331 13388
rect 14297 13286 14331 13320
rect 14297 13218 14331 13252
rect 14297 13150 14331 13184
rect 14297 13082 14331 13116
rect 14297 13014 14331 13048
rect 14297 12946 14331 12980
rect 14297 12878 14331 12912
rect 14297 12810 14331 12844
rect 14297 12742 14331 12776
rect 14297 12674 14331 12708
rect 14297 12606 14331 12640
rect 14297 12538 14331 12572
rect 14297 12470 14331 12504
rect 14297 12402 14331 12436
rect 14297 12334 14331 12368
rect 14297 12266 14331 12300
rect 14297 12198 14331 12232
rect 14297 12130 14331 12164
rect 14297 12062 14331 12096
rect 14297 11994 14331 12028
rect 14297 11926 14331 11960
rect 14297 11858 14331 11892
rect 14297 11790 14331 11824
rect 14297 11722 14331 11756
rect 14297 11654 14331 11688
rect 14297 11586 14331 11620
rect 14297 11518 14331 11552
rect 14297 11450 14331 11484
rect 14297 11382 14331 11416
rect 14297 11314 14331 11348
rect 14297 11246 14331 11280
rect 14297 11178 14331 11212
rect 14297 11110 14331 11144
rect 14297 11042 14331 11076
rect 14297 10974 14331 11008
rect 14297 10906 14331 10940
rect 14297 10838 14331 10872
rect 14297 10770 14331 10804
rect 14297 10702 14331 10736
rect 14297 10634 14331 10668
rect 14297 10566 14331 10600
rect 14297 10498 14331 10532
rect 14297 10430 14331 10464
rect 14297 10362 14331 10396
rect 14297 10294 14331 10328
rect 14297 10226 14331 10260
rect 632 10158 666 10192
rect 632 10090 666 10124
rect 632 10022 666 10056
rect 632 9954 666 9988
rect 632 9886 666 9920
rect 14297 10158 14331 10192
rect 14297 10090 14331 10124
rect 14297 10022 14331 10056
rect 14297 9954 14331 9988
rect 14297 9886 14331 9920
rect 766 9741 800 9775
rect 834 9741 868 9775
rect 902 9741 936 9775
rect 970 9741 1004 9775
rect 1038 9741 1072 9775
rect 1106 9741 1140 9775
rect 1174 9741 1208 9775
rect 1242 9741 1276 9775
rect 1310 9741 1344 9775
rect 1378 9741 1412 9775
rect 1446 9741 1480 9775
rect 1514 9741 1548 9775
rect 1582 9741 1616 9775
rect 1650 9741 1684 9775
rect 1718 9741 1752 9775
rect 1786 9741 1820 9775
rect 1854 9741 1888 9775
rect 1922 9741 1956 9775
rect 1990 9741 2024 9775
rect 2058 9741 2092 9775
rect 2126 9741 2160 9775
rect 2194 9741 2228 9775
rect 2262 9741 2296 9775
rect 2330 9741 2364 9775
rect 2398 9741 2432 9775
rect 2466 9741 2500 9775
rect 2534 9741 2568 9775
rect 2602 9741 2636 9775
rect 2670 9741 2704 9775
rect 2738 9741 2772 9775
rect 2806 9741 2840 9775
rect 2874 9741 2908 9775
rect 2942 9741 2976 9775
rect 3010 9741 3044 9775
rect 3078 9741 3112 9775
rect 3146 9741 3180 9775
rect 3214 9741 3248 9775
rect 3282 9741 3316 9775
rect 3350 9741 3384 9775
rect 3418 9741 3452 9775
rect 3486 9741 3520 9775
rect 3554 9741 3588 9775
rect 3622 9741 3656 9775
rect 3690 9741 3724 9775
rect 3758 9741 3792 9775
rect 3826 9741 3860 9775
rect 3894 9741 3928 9775
rect 3962 9741 3996 9775
rect 4030 9741 4064 9775
rect 4098 9741 4132 9775
rect 4166 9741 4200 9775
rect 4234 9741 4268 9775
rect 4302 9741 4336 9775
rect 4370 9741 4404 9775
rect 4438 9741 4472 9775
rect 4506 9741 4540 9775
rect 4574 9741 4608 9775
rect 4642 9741 4676 9775
rect 4710 9741 4744 9775
rect 4778 9741 4812 9775
rect 4846 9741 4880 9775
rect 4914 9741 4948 9775
rect 4982 9741 5016 9775
rect 5050 9741 5084 9775
rect 5118 9741 5152 9775
rect 5186 9741 5220 9775
rect 5254 9741 5288 9775
rect 5322 9741 5356 9775
rect 5390 9741 5424 9775
rect 5458 9741 5492 9775
rect 5526 9741 5560 9775
rect 5594 9741 5628 9775
rect 5662 9741 5696 9775
rect 5730 9741 5764 9775
rect 5798 9741 5832 9775
rect 5866 9741 5900 9775
rect 5934 9741 5968 9775
rect 6002 9741 6036 9775
rect 6070 9741 6104 9775
rect 6138 9741 6172 9775
rect 6206 9741 6240 9775
rect 6274 9741 6308 9775
rect 6342 9741 6376 9775
rect 6410 9741 6444 9775
rect 6478 9741 6512 9775
rect 6546 9741 6580 9775
rect 6614 9741 6648 9775
rect 6682 9741 6716 9775
rect 6750 9741 6784 9775
rect 6818 9741 6852 9775
rect 6886 9741 6920 9775
rect 6954 9741 6988 9775
rect 7022 9741 7056 9775
rect 7090 9741 7124 9775
rect 7158 9741 7192 9775
rect 7226 9741 7260 9775
rect 7294 9741 7328 9775
rect 7362 9741 7396 9775
rect 7430 9741 7464 9775
rect 7498 9741 7532 9775
rect 7566 9741 7600 9775
rect 7634 9741 7668 9775
rect 7702 9741 7736 9775
rect 7770 9741 7804 9775
rect 7838 9741 7872 9775
rect 7906 9741 7940 9775
rect 7974 9741 8008 9775
rect 8042 9741 8076 9775
rect 8110 9741 8144 9775
rect 8178 9741 8212 9775
rect 8246 9741 8280 9775
rect 8314 9741 8348 9775
rect 8382 9741 8416 9775
rect 8450 9741 8484 9775
rect 8518 9741 8552 9775
rect 8586 9741 8620 9775
rect 8654 9741 8688 9775
rect 8722 9741 8756 9775
rect 8790 9741 8824 9775
rect 8858 9741 8892 9775
rect 8926 9741 8960 9775
rect 8994 9741 9028 9775
rect 9062 9741 9096 9775
rect 9130 9741 9164 9775
rect 9198 9741 9232 9775
rect 9266 9741 9300 9775
rect 9334 9741 9368 9775
rect 9402 9741 9436 9775
rect 9470 9741 9504 9775
rect 9538 9741 9572 9775
rect 9606 9741 9640 9775
rect 9674 9741 9708 9775
rect 9742 9741 9776 9775
rect 9810 9741 9844 9775
rect 9878 9741 9912 9775
rect 9946 9741 9980 9775
rect 10014 9741 10048 9775
rect 10082 9741 10116 9775
rect 10150 9741 10184 9775
rect 10218 9741 10252 9775
rect 10286 9741 10320 9775
rect 10354 9741 10388 9775
rect 10422 9741 10456 9775
rect 10490 9741 10524 9775
rect 10558 9741 10592 9775
rect 10626 9741 10660 9775
rect 10694 9741 10728 9775
rect 10762 9741 10796 9775
rect 10830 9741 10864 9775
rect 10898 9741 10932 9775
rect 10966 9741 11000 9775
rect 11034 9741 11068 9775
rect 11102 9741 11136 9775
rect 11170 9741 11204 9775
rect 11238 9741 11272 9775
rect 11306 9741 11340 9775
rect 11374 9741 11408 9775
rect 11442 9741 11476 9775
rect 11510 9741 11544 9775
rect 11578 9741 11612 9775
rect 11646 9741 11680 9775
rect 11714 9741 11748 9775
rect 11782 9741 11816 9775
rect 11850 9741 11884 9775
rect 11918 9741 11952 9775
rect 11986 9741 12020 9775
rect 12054 9741 12088 9775
rect 12122 9741 12156 9775
rect 12190 9741 12224 9775
rect 12258 9741 12292 9775
rect 12326 9741 12360 9775
rect 12394 9741 12428 9775
rect 12462 9741 12496 9775
rect 12530 9741 12564 9775
rect 12598 9741 12632 9775
rect 12666 9741 12700 9775
rect 12734 9741 12768 9775
rect 12802 9741 12836 9775
rect 12870 9741 12904 9775
rect 12938 9741 12972 9775
rect 13006 9741 13040 9775
rect 13074 9741 13108 9775
rect 13142 9741 13176 9775
rect 13210 9741 13244 9775
rect 13278 9741 13312 9775
rect 13346 9741 13380 9775
rect 13414 9741 13448 9775
rect 13482 9741 13516 9775
rect 13550 9741 13584 9775
rect 13618 9741 13652 9775
rect 13686 9741 13720 9775
rect 13754 9741 13788 9775
rect 13822 9741 13856 9775
rect 13890 9741 13924 9775
rect 13958 9741 13992 9775
rect 14026 9741 14060 9775
rect 14094 9741 14128 9775
rect 14162 9741 14196 9775
<< locali >>
rect 245 36534 14724 36574
rect 245 36500 320 36534
rect 354 36533 14724 36534
rect 354 36500 14614 36533
rect 245 36499 14614 36500
rect 14648 36499 14724 36533
rect 245 36498 14724 36499
rect 245 36497 556 36498
rect 590 36497 628 36498
rect 662 36497 700 36498
rect 734 36497 772 36498
rect 806 36497 844 36498
rect 878 36497 916 36498
rect 950 36497 988 36498
rect 1022 36497 1060 36498
rect 1094 36497 1132 36498
rect 1166 36497 1204 36498
rect 1238 36497 1276 36498
rect 1310 36497 1348 36498
rect 1382 36497 1420 36498
rect 1454 36497 1492 36498
rect 1526 36497 1564 36498
rect 1598 36497 1636 36498
rect 1670 36497 1708 36498
rect 1742 36497 1780 36498
rect 1814 36497 1852 36498
rect 1886 36497 1924 36498
rect 1958 36497 1996 36498
rect 2030 36497 2068 36498
rect 2102 36497 2140 36498
rect 2174 36497 2212 36498
rect 2246 36497 2284 36498
rect 2318 36497 2356 36498
rect 2390 36497 2428 36498
rect 2462 36497 2500 36498
rect 2534 36497 2572 36498
rect 2606 36497 2644 36498
rect 2678 36497 2716 36498
rect 2750 36497 2788 36498
rect 2822 36497 2860 36498
rect 2894 36497 2932 36498
rect 2966 36497 3004 36498
rect 3038 36497 3076 36498
rect 3110 36497 3148 36498
rect 3182 36497 3220 36498
rect 3254 36497 3292 36498
rect 3326 36497 3364 36498
rect 3398 36497 3436 36498
rect 3470 36497 3508 36498
rect 3542 36497 3580 36498
rect 3614 36497 3652 36498
rect 3686 36497 3724 36498
rect 3758 36497 3796 36498
rect 3830 36497 3868 36498
rect 3902 36497 3940 36498
rect 3974 36497 4012 36498
rect 4046 36497 4084 36498
rect 4118 36497 4156 36498
rect 4190 36497 4228 36498
rect 4262 36497 4300 36498
rect 4334 36497 4372 36498
rect 4406 36497 4444 36498
rect 4478 36497 4516 36498
rect 4550 36497 4588 36498
rect 4622 36497 4660 36498
rect 4694 36497 4732 36498
rect 4766 36497 4804 36498
rect 4838 36497 4876 36498
rect 4910 36497 4948 36498
rect 4982 36497 5020 36498
rect 5054 36497 5092 36498
rect 5126 36497 5164 36498
rect 5198 36497 5236 36498
rect 5270 36497 5308 36498
rect 5342 36497 5380 36498
rect 5414 36497 5452 36498
rect 5486 36497 5524 36498
rect 5558 36497 5596 36498
rect 5630 36497 5668 36498
rect 5702 36497 5740 36498
rect 5774 36497 5812 36498
rect 5846 36497 5884 36498
rect 5918 36497 5956 36498
rect 5990 36497 6028 36498
rect 6062 36497 6100 36498
rect 6134 36497 6172 36498
rect 6206 36497 6244 36498
rect 6278 36497 6316 36498
rect 6350 36497 6388 36498
rect 6422 36497 6460 36498
rect 6494 36497 6532 36498
rect 6566 36497 6604 36498
rect 6638 36497 6676 36498
rect 6710 36497 6748 36498
rect 6782 36497 6820 36498
rect 6854 36497 6892 36498
rect 6926 36497 6964 36498
rect 6998 36497 7036 36498
rect 7070 36497 7108 36498
rect 7142 36497 7180 36498
rect 7214 36497 7252 36498
rect 7286 36497 7324 36498
rect 7358 36497 7396 36498
rect 7430 36497 7468 36498
rect 7502 36497 7540 36498
rect 7574 36497 7612 36498
rect 7646 36497 7684 36498
rect 7718 36497 7756 36498
rect 7790 36497 7828 36498
rect 7862 36497 7900 36498
rect 7934 36497 7972 36498
rect 8006 36497 8044 36498
rect 8078 36497 8116 36498
rect 8150 36497 8188 36498
rect 8222 36497 8260 36498
rect 8294 36497 8332 36498
rect 8366 36497 8404 36498
rect 8438 36497 8476 36498
rect 8510 36497 8548 36498
rect 8582 36497 8620 36498
rect 8654 36497 8692 36498
rect 8726 36497 8764 36498
rect 8798 36497 8836 36498
rect 8870 36497 8908 36498
rect 8942 36497 8980 36498
rect 9014 36497 9052 36498
rect 9086 36497 9124 36498
rect 9158 36497 9196 36498
rect 9230 36497 9268 36498
rect 9302 36497 9340 36498
rect 9374 36497 9412 36498
rect 9446 36497 9484 36498
rect 9518 36497 9556 36498
rect 9590 36497 9628 36498
rect 9662 36497 9700 36498
rect 9734 36497 9772 36498
rect 9806 36497 9844 36498
rect 9878 36497 9916 36498
rect 9950 36497 9988 36498
rect 10022 36497 10060 36498
rect 10094 36497 10132 36498
rect 10166 36497 10204 36498
rect 10238 36497 10276 36498
rect 10310 36497 10348 36498
rect 10382 36497 10420 36498
rect 10454 36497 10492 36498
rect 10526 36497 10564 36498
rect 10598 36497 10636 36498
rect 10670 36497 10708 36498
rect 10742 36497 10780 36498
rect 10814 36497 10852 36498
rect 10886 36497 10924 36498
rect 10958 36497 10996 36498
rect 11030 36497 11068 36498
rect 11102 36497 11140 36498
rect 11174 36497 11212 36498
rect 11246 36497 11284 36498
rect 11318 36497 11356 36498
rect 11390 36497 11428 36498
rect 11462 36497 11500 36498
rect 11534 36497 11572 36498
rect 11606 36497 11644 36498
rect 11678 36497 11716 36498
rect 11750 36497 11788 36498
rect 11822 36497 11860 36498
rect 11894 36497 11932 36498
rect 11966 36497 12004 36498
rect 12038 36497 12076 36498
rect 12110 36497 12148 36498
rect 12182 36497 12220 36498
rect 12254 36497 12292 36498
rect 12326 36497 12364 36498
rect 12398 36497 12436 36498
rect 12470 36497 12508 36498
rect 12542 36497 12580 36498
rect 12614 36497 12652 36498
rect 12686 36497 12724 36498
rect 12758 36497 12796 36498
rect 12830 36497 12868 36498
rect 12902 36497 12940 36498
rect 12974 36497 13012 36498
rect 13046 36497 13084 36498
rect 13118 36497 13156 36498
rect 13190 36497 13228 36498
rect 13262 36497 13300 36498
rect 13334 36497 13372 36498
rect 13406 36497 13444 36498
rect 13478 36497 13516 36498
rect 13550 36497 13588 36498
rect 13622 36497 13660 36498
rect 13694 36497 13732 36498
rect 13766 36497 13804 36498
rect 13838 36497 13876 36498
rect 13910 36497 13948 36498
rect 13982 36497 14020 36498
rect 14054 36497 14092 36498
rect 14126 36497 14164 36498
rect 14198 36497 14236 36498
rect 14270 36497 14308 36498
rect 14342 36497 14380 36498
rect 14414 36497 14724 36498
rect 245 36463 455 36497
rect 489 36463 523 36497
rect 590 36464 591 36497
rect 557 36463 591 36464
rect 625 36464 628 36497
rect 693 36464 700 36497
rect 761 36464 772 36497
rect 829 36464 844 36497
rect 897 36464 916 36497
rect 965 36464 988 36497
rect 1033 36464 1060 36497
rect 1101 36464 1132 36497
rect 625 36463 659 36464
rect 693 36463 727 36464
rect 761 36463 795 36464
rect 829 36463 863 36464
rect 897 36463 931 36464
rect 965 36463 999 36464
rect 1033 36463 1067 36464
rect 1101 36463 1135 36464
rect 1169 36463 1203 36497
rect 1238 36464 1271 36497
rect 1310 36464 1339 36497
rect 1382 36464 1407 36497
rect 1454 36464 1475 36497
rect 1526 36464 1543 36497
rect 1598 36464 1611 36497
rect 1670 36464 1679 36497
rect 1742 36464 1747 36497
rect 1814 36464 1815 36497
rect 1237 36463 1271 36464
rect 1305 36463 1339 36464
rect 1373 36463 1407 36464
rect 1441 36463 1475 36464
rect 1509 36463 1543 36464
rect 1577 36463 1611 36464
rect 1645 36463 1679 36464
rect 1713 36463 1747 36464
rect 1781 36463 1815 36464
rect 1849 36464 1852 36497
rect 1917 36464 1924 36497
rect 1985 36464 1996 36497
rect 2053 36464 2068 36497
rect 2121 36464 2140 36497
rect 2189 36464 2212 36497
rect 2257 36464 2284 36497
rect 2325 36464 2356 36497
rect 1849 36463 1883 36464
rect 1917 36463 1951 36464
rect 1985 36463 2019 36464
rect 2053 36463 2087 36464
rect 2121 36463 2155 36464
rect 2189 36463 2223 36464
rect 2257 36463 2291 36464
rect 2325 36463 2359 36464
rect 2393 36463 2427 36497
rect 2462 36464 2495 36497
rect 2534 36464 2563 36497
rect 2606 36464 2631 36497
rect 2678 36464 2699 36497
rect 2750 36464 2767 36497
rect 2822 36464 2835 36497
rect 2894 36464 2903 36497
rect 2966 36464 2971 36497
rect 3038 36464 3039 36497
rect 2461 36463 2495 36464
rect 2529 36463 2563 36464
rect 2597 36463 2631 36464
rect 2665 36463 2699 36464
rect 2733 36463 2767 36464
rect 2801 36463 2835 36464
rect 2869 36463 2903 36464
rect 2937 36463 2971 36464
rect 3005 36463 3039 36464
rect 3073 36464 3076 36497
rect 3141 36464 3148 36497
rect 3209 36464 3220 36497
rect 3277 36464 3292 36497
rect 3345 36464 3364 36497
rect 3413 36464 3436 36497
rect 3481 36464 3508 36497
rect 3549 36464 3580 36497
rect 3073 36463 3107 36464
rect 3141 36463 3175 36464
rect 3209 36463 3243 36464
rect 3277 36463 3311 36464
rect 3345 36463 3379 36464
rect 3413 36463 3447 36464
rect 3481 36463 3515 36464
rect 3549 36463 3583 36464
rect 3617 36463 3651 36497
rect 3686 36464 3719 36497
rect 3758 36464 3787 36497
rect 3830 36464 3855 36497
rect 3902 36464 3923 36497
rect 3974 36464 3991 36497
rect 4046 36464 4059 36497
rect 4118 36464 4127 36497
rect 4190 36464 4195 36497
rect 4262 36464 4263 36497
rect 3685 36463 3719 36464
rect 3753 36463 3787 36464
rect 3821 36463 3855 36464
rect 3889 36463 3923 36464
rect 3957 36463 3991 36464
rect 4025 36463 4059 36464
rect 4093 36463 4127 36464
rect 4161 36463 4195 36464
rect 4229 36463 4263 36464
rect 4297 36464 4300 36497
rect 4365 36464 4372 36497
rect 4433 36464 4444 36497
rect 4501 36464 4516 36497
rect 4569 36464 4588 36497
rect 4637 36464 4660 36497
rect 4705 36464 4732 36497
rect 4773 36464 4804 36497
rect 4297 36463 4331 36464
rect 4365 36463 4399 36464
rect 4433 36463 4467 36464
rect 4501 36463 4535 36464
rect 4569 36463 4603 36464
rect 4637 36463 4671 36464
rect 4705 36463 4739 36464
rect 4773 36463 4807 36464
rect 4841 36463 4875 36497
rect 4910 36464 4943 36497
rect 4982 36464 5011 36497
rect 5054 36464 5079 36497
rect 5126 36464 5147 36497
rect 5198 36464 5215 36497
rect 5270 36464 5283 36497
rect 5342 36464 5351 36497
rect 5414 36464 5419 36497
rect 5486 36464 5487 36497
rect 4909 36463 4943 36464
rect 4977 36463 5011 36464
rect 5045 36463 5079 36464
rect 5113 36463 5147 36464
rect 5181 36463 5215 36464
rect 5249 36463 5283 36464
rect 5317 36463 5351 36464
rect 5385 36463 5419 36464
rect 5453 36463 5487 36464
rect 5521 36464 5524 36497
rect 5589 36464 5596 36497
rect 5657 36464 5668 36497
rect 5725 36464 5740 36497
rect 5793 36464 5812 36497
rect 5861 36464 5884 36497
rect 5929 36464 5956 36497
rect 5997 36464 6028 36497
rect 5521 36463 5555 36464
rect 5589 36463 5623 36464
rect 5657 36463 5691 36464
rect 5725 36463 5759 36464
rect 5793 36463 5827 36464
rect 5861 36463 5895 36464
rect 5929 36463 5963 36464
rect 5997 36463 6031 36464
rect 6065 36463 6099 36497
rect 6134 36464 6167 36497
rect 6206 36464 6235 36497
rect 6278 36464 6303 36497
rect 6350 36464 6371 36497
rect 6422 36464 6439 36497
rect 6494 36464 6507 36497
rect 6566 36464 6575 36497
rect 6638 36464 6643 36497
rect 6710 36464 6711 36497
rect 6133 36463 6167 36464
rect 6201 36463 6235 36464
rect 6269 36463 6303 36464
rect 6337 36463 6371 36464
rect 6405 36463 6439 36464
rect 6473 36463 6507 36464
rect 6541 36463 6575 36464
rect 6609 36463 6643 36464
rect 6677 36463 6711 36464
rect 6745 36464 6748 36497
rect 6813 36464 6820 36497
rect 6881 36464 6892 36497
rect 6949 36464 6964 36497
rect 7017 36464 7036 36497
rect 7085 36464 7108 36497
rect 7153 36464 7180 36497
rect 7221 36464 7252 36497
rect 6745 36463 6779 36464
rect 6813 36463 6847 36464
rect 6881 36463 6915 36464
rect 6949 36463 6983 36464
rect 7017 36463 7051 36464
rect 7085 36463 7119 36464
rect 7153 36463 7187 36464
rect 7221 36463 7255 36464
rect 7289 36463 7323 36497
rect 7358 36464 7391 36497
rect 7430 36464 7459 36497
rect 7502 36464 7527 36497
rect 7574 36464 7595 36497
rect 7646 36464 7663 36497
rect 7718 36464 7731 36497
rect 7790 36464 7799 36497
rect 7862 36464 7867 36497
rect 7934 36464 7935 36497
rect 7357 36463 7391 36464
rect 7425 36463 7459 36464
rect 7493 36463 7527 36464
rect 7561 36463 7595 36464
rect 7629 36463 7663 36464
rect 7697 36463 7731 36464
rect 7765 36463 7799 36464
rect 7833 36463 7867 36464
rect 7901 36463 7935 36464
rect 7969 36464 7972 36497
rect 8037 36464 8044 36497
rect 8105 36464 8116 36497
rect 8173 36464 8188 36497
rect 8241 36464 8260 36497
rect 8309 36464 8332 36497
rect 8377 36464 8404 36497
rect 8445 36464 8476 36497
rect 7969 36463 8003 36464
rect 8037 36463 8071 36464
rect 8105 36463 8139 36464
rect 8173 36463 8207 36464
rect 8241 36463 8275 36464
rect 8309 36463 8343 36464
rect 8377 36463 8411 36464
rect 8445 36463 8479 36464
rect 8513 36463 8547 36497
rect 8582 36464 8615 36497
rect 8654 36464 8683 36497
rect 8726 36464 8751 36497
rect 8798 36464 8819 36497
rect 8870 36464 8887 36497
rect 8942 36464 8955 36497
rect 9014 36464 9023 36497
rect 9086 36464 9091 36497
rect 9158 36464 9159 36497
rect 8581 36463 8615 36464
rect 8649 36463 8683 36464
rect 8717 36463 8751 36464
rect 8785 36463 8819 36464
rect 8853 36463 8887 36464
rect 8921 36463 8955 36464
rect 8989 36463 9023 36464
rect 9057 36463 9091 36464
rect 9125 36463 9159 36464
rect 9193 36464 9196 36497
rect 9261 36464 9268 36497
rect 9329 36464 9340 36497
rect 9397 36464 9412 36497
rect 9465 36464 9484 36497
rect 9533 36464 9556 36497
rect 9601 36464 9628 36497
rect 9669 36464 9700 36497
rect 9193 36463 9227 36464
rect 9261 36463 9295 36464
rect 9329 36463 9363 36464
rect 9397 36463 9431 36464
rect 9465 36463 9499 36464
rect 9533 36463 9567 36464
rect 9601 36463 9635 36464
rect 9669 36463 9703 36464
rect 9737 36463 9771 36497
rect 9806 36464 9839 36497
rect 9878 36464 9907 36497
rect 9950 36464 9975 36497
rect 10022 36464 10043 36497
rect 10094 36464 10111 36497
rect 10166 36464 10179 36497
rect 10238 36464 10247 36497
rect 10310 36464 10315 36497
rect 10382 36464 10383 36497
rect 9805 36463 9839 36464
rect 9873 36463 9907 36464
rect 9941 36463 9975 36464
rect 10009 36463 10043 36464
rect 10077 36463 10111 36464
rect 10145 36463 10179 36464
rect 10213 36463 10247 36464
rect 10281 36463 10315 36464
rect 10349 36463 10383 36464
rect 10417 36464 10420 36497
rect 10485 36464 10492 36497
rect 10553 36464 10564 36497
rect 10621 36464 10636 36497
rect 10689 36464 10708 36497
rect 10757 36464 10780 36497
rect 10825 36464 10852 36497
rect 10893 36464 10924 36497
rect 10417 36463 10451 36464
rect 10485 36463 10519 36464
rect 10553 36463 10587 36464
rect 10621 36463 10655 36464
rect 10689 36463 10723 36464
rect 10757 36463 10791 36464
rect 10825 36463 10859 36464
rect 10893 36463 10927 36464
rect 10961 36463 10995 36497
rect 11030 36464 11063 36497
rect 11102 36464 11131 36497
rect 11174 36464 11199 36497
rect 11246 36464 11267 36497
rect 11318 36464 11335 36497
rect 11390 36464 11403 36497
rect 11462 36464 11471 36497
rect 11534 36464 11539 36497
rect 11606 36464 11607 36497
rect 11029 36463 11063 36464
rect 11097 36463 11131 36464
rect 11165 36463 11199 36464
rect 11233 36463 11267 36464
rect 11301 36463 11335 36464
rect 11369 36463 11403 36464
rect 11437 36463 11471 36464
rect 11505 36463 11539 36464
rect 11573 36463 11607 36464
rect 11641 36464 11644 36497
rect 11709 36464 11716 36497
rect 11777 36464 11788 36497
rect 11845 36464 11860 36497
rect 11913 36464 11932 36497
rect 11981 36464 12004 36497
rect 12049 36464 12076 36497
rect 12117 36464 12148 36497
rect 11641 36463 11675 36464
rect 11709 36463 11743 36464
rect 11777 36463 11811 36464
rect 11845 36463 11879 36464
rect 11913 36463 11947 36464
rect 11981 36463 12015 36464
rect 12049 36463 12083 36464
rect 12117 36463 12151 36464
rect 12185 36463 12219 36497
rect 12254 36464 12287 36497
rect 12326 36464 12355 36497
rect 12398 36464 12423 36497
rect 12470 36464 12491 36497
rect 12542 36464 12559 36497
rect 12614 36464 12627 36497
rect 12686 36464 12695 36497
rect 12758 36464 12763 36497
rect 12830 36464 12831 36497
rect 12253 36463 12287 36464
rect 12321 36463 12355 36464
rect 12389 36463 12423 36464
rect 12457 36463 12491 36464
rect 12525 36463 12559 36464
rect 12593 36463 12627 36464
rect 12661 36463 12695 36464
rect 12729 36463 12763 36464
rect 12797 36463 12831 36464
rect 12865 36464 12868 36497
rect 12933 36464 12940 36497
rect 13001 36464 13012 36497
rect 13069 36464 13084 36497
rect 13137 36464 13156 36497
rect 13205 36464 13228 36497
rect 13273 36464 13300 36497
rect 13341 36464 13372 36497
rect 12865 36463 12899 36464
rect 12933 36463 12967 36464
rect 13001 36463 13035 36464
rect 13069 36463 13103 36464
rect 13137 36463 13171 36464
rect 13205 36463 13239 36464
rect 13273 36463 13307 36464
rect 13341 36463 13375 36464
rect 13409 36463 13443 36497
rect 13478 36464 13511 36497
rect 13550 36464 13579 36497
rect 13622 36464 13647 36497
rect 13694 36464 13715 36497
rect 13766 36464 13783 36497
rect 13838 36464 13851 36497
rect 13910 36464 13919 36497
rect 13982 36464 13987 36497
rect 14054 36464 14055 36497
rect 13477 36463 13511 36464
rect 13545 36463 13579 36464
rect 13613 36463 13647 36464
rect 13681 36463 13715 36464
rect 13749 36463 13783 36464
rect 13817 36463 13851 36464
rect 13885 36463 13919 36464
rect 13953 36463 13987 36464
rect 14021 36463 14055 36464
rect 14089 36464 14092 36497
rect 14157 36464 14164 36497
rect 14225 36464 14236 36497
rect 14293 36464 14308 36497
rect 14361 36464 14380 36497
rect 14089 36463 14123 36464
rect 14157 36463 14191 36464
rect 14225 36463 14259 36464
rect 14293 36463 14327 36464
rect 14361 36463 14395 36464
rect 14429 36463 14463 36497
rect 14497 36463 14724 36497
rect 245 36462 14724 36463
rect 245 36428 320 36462
rect 354 36461 14724 36462
rect 354 36428 14614 36461
rect 245 36427 14614 36428
rect 14648 36427 14724 36461
rect 245 36389 14724 36427
rect 245 36338 430 36389
rect 245 36304 312 36338
rect 346 36304 430 36338
rect 245 36270 430 36304
rect 245 36236 312 36270
rect 346 36265 430 36270
rect 245 36231 320 36236
rect 354 36231 430 36265
rect 245 36202 430 36231
rect 14539 36344 14724 36389
rect 14539 36310 14607 36344
rect 14641 36310 14724 36344
rect 14539 36276 14724 36310
rect 14539 36242 14607 36276
rect 14641 36262 14724 36276
rect 14539 36228 14614 36242
rect 14648 36228 14724 36262
rect 14539 36208 14724 36228
rect 245 36168 312 36202
rect 346 36193 430 36202
rect 245 36159 320 36168
rect 354 36159 430 36193
rect 245 36134 430 36159
rect 245 36100 312 36134
rect 346 36121 430 36134
rect 245 36087 320 36100
rect 354 36087 430 36121
rect 245 36066 430 36087
rect 245 36032 312 36066
rect 346 36049 430 36066
rect 245 36015 320 36032
rect 354 36015 430 36049
rect 245 35998 430 36015
rect 245 35964 312 35998
rect 346 35977 430 35998
rect 245 35943 320 35964
rect 354 35943 430 35977
rect 245 35930 430 35943
rect 245 35896 312 35930
rect 346 35905 430 35930
rect 245 35871 320 35896
rect 354 35871 430 35905
rect 245 35862 430 35871
rect 245 35828 312 35862
rect 346 35833 430 35862
rect 245 35799 320 35828
rect 354 35799 430 35833
rect 245 35794 430 35799
rect 245 35760 312 35794
rect 346 35761 430 35794
rect 245 35727 320 35760
rect 354 35727 430 35761
rect 245 35726 430 35727
rect 245 35692 312 35726
rect 346 35692 430 35726
rect 245 35689 430 35692
rect 245 35658 320 35689
rect 245 35624 312 35658
rect 354 35655 430 35689
rect 346 35624 430 35655
rect 245 35617 430 35624
rect 245 35590 320 35617
rect 245 35556 312 35590
rect 354 35583 430 35617
rect 346 35556 430 35583
rect 245 35545 430 35556
rect 245 35522 320 35545
rect 245 35488 312 35522
rect 354 35511 430 35545
rect 346 35488 430 35511
rect 245 35473 430 35488
rect 245 35454 320 35473
rect 245 35420 312 35454
rect 354 35439 430 35473
rect 346 35420 430 35439
rect 245 35401 430 35420
rect 245 35386 320 35401
rect 245 35352 312 35386
rect 354 35367 430 35401
rect 346 35352 430 35367
rect 245 35329 430 35352
rect 245 35318 320 35329
rect 245 35284 312 35318
rect 354 35295 430 35329
rect 346 35284 430 35295
rect 245 35257 430 35284
rect 245 35250 320 35257
rect 245 35216 312 35250
rect 354 35223 430 35257
rect 346 35216 430 35223
rect 245 35185 430 35216
rect 245 35182 320 35185
rect 245 35148 312 35182
rect 354 35151 430 35185
rect 346 35148 430 35151
rect 245 35114 430 35148
rect 245 35080 312 35114
rect 346 35113 430 35114
rect 245 35079 320 35080
rect 354 35079 430 35113
rect 245 35046 430 35079
rect 245 35012 312 35046
rect 346 35041 430 35046
rect 245 35007 320 35012
rect 354 35007 430 35041
rect 245 34978 430 35007
rect 245 34944 312 34978
rect 346 34969 430 34978
rect 245 34935 320 34944
rect 354 34935 430 34969
rect 245 34910 430 34935
rect 245 34876 312 34910
rect 346 34897 430 34910
rect 245 34863 320 34876
rect 354 34863 430 34897
rect 245 34842 430 34863
rect 245 34808 312 34842
rect 346 34825 430 34842
rect 245 34791 320 34808
rect 354 34791 430 34825
rect 245 34774 430 34791
rect 245 34740 312 34774
rect 346 34753 430 34774
rect 245 34719 320 34740
rect 354 34719 430 34753
rect 245 34706 430 34719
rect 245 34672 312 34706
rect 346 34681 430 34706
rect 245 34647 320 34672
rect 354 34647 430 34681
rect 245 34638 430 34647
rect 245 34604 312 34638
rect 346 34609 430 34638
rect 245 34575 320 34604
rect 354 34575 430 34609
rect 245 34570 430 34575
rect 245 34536 312 34570
rect 346 34537 430 34570
rect 245 34503 320 34536
rect 354 34503 430 34537
rect 245 34502 430 34503
rect 245 34468 312 34502
rect 346 34468 430 34502
rect 245 34465 430 34468
rect 245 34434 320 34465
rect 245 34400 312 34434
rect 354 34431 430 34465
rect 346 34400 430 34431
rect 245 34393 430 34400
rect 245 34366 320 34393
rect 245 34332 312 34366
rect 354 34359 430 34393
rect 346 34332 430 34359
rect 245 34321 430 34332
rect 245 34298 320 34321
rect 245 34264 312 34298
rect 354 34287 430 34321
rect 346 34264 430 34287
rect 245 34249 430 34264
rect 245 34230 320 34249
rect 245 34196 312 34230
rect 354 34215 430 34249
rect 346 34196 430 34215
rect 245 34177 430 34196
rect 245 34162 320 34177
rect 245 34128 312 34162
rect 354 34143 430 34177
rect 346 34128 430 34143
rect 245 34105 430 34128
rect 245 34094 320 34105
rect 245 34060 312 34094
rect 354 34071 430 34105
rect 346 34060 430 34071
rect 245 34033 430 34060
rect 245 34026 320 34033
rect 245 33992 312 34026
rect 354 33999 430 34033
rect 346 33992 430 33999
rect 245 33961 430 33992
rect 245 33958 320 33961
rect 245 33924 312 33958
rect 354 33927 430 33961
rect 346 33924 430 33927
rect 245 33890 430 33924
rect 245 33856 312 33890
rect 346 33889 430 33890
rect 245 33855 320 33856
rect 354 33855 430 33889
rect 245 33822 430 33855
rect 245 33788 312 33822
rect 346 33817 430 33822
rect 245 33783 320 33788
rect 354 33783 430 33817
rect 245 33754 430 33783
rect 245 33720 312 33754
rect 346 33745 430 33754
rect 245 33711 320 33720
rect 354 33711 430 33745
rect 245 33686 430 33711
rect 245 33652 312 33686
rect 346 33673 430 33686
rect 245 33639 320 33652
rect 354 33639 430 33673
rect 245 33618 430 33639
rect 245 33584 312 33618
rect 346 33601 430 33618
rect 245 33567 320 33584
rect 354 33567 430 33601
rect 245 33550 430 33567
rect 245 33516 312 33550
rect 346 33529 430 33550
rect 245 33495 320 33516
rect 354 33495 430 33529
rect 245 33482 430 33495
rect 245 33448 312 33482
rect 346 33457 430 33482
rect 245 33423 320 33448
rect 354 33423 430 33457
rect 245 33414 430 33423
rect 245 33380 312 33414
rect 346 33385 430 33414
rect 245 33351 320 33380
rect 354 33351 430 33385
rect 245 33346 430 33351
rect 245 33312 312 33346
rect 346 33313 430 33346
rect 245 33279 320 33312
rect 354 33279 430 33313
rect 245 33278 430 33279
rect 245 33244 312 33278
rect 346 33244 430 33278
rect 245 33241 430 33244
rect 245 33210 320 33241
rect 245 33176 312 33210
rect 354 33207 430 33241
rect 346 33176 430 33207
rect 245 33169 430 33176
rect 245 33142 320 33169
rect 245 33108 312 33142
rect 354 33135 430 33169
rect 346 33108 430 33135
rect 245 33097 430 33108
rect 245 33074 320 33097
rect 245 33040 312 33074
rect 354 33063 430 33097
rect 346 33040 430 33063
rect 245 33025 430 33040
rect 245 33006 320 33025
rect 245 32972 312 33006
rect 354 32991 430 33025
rect 346 32972 430 32991
rect 245 32953 430 32972
rect 245 32938 320 32953
rect 245 32904 312 32938
rect 354 32919 430 32953
rect 346 32904 430 32919
rect 245 32881 430 32904
rect 245 32870 320 32881
rect 245 32836 312 32870
rect 354 32847 430 32881
rect 346 32836 430 32847
rect 245 32809 430 32836
rect 245 32802 320 32809
rect 245 32768 312 32802
rect 354 32775 430 32809
rect 346 32768 430 32775
rect 245 32737 430 32768
rect 245 32734 320 32737
rect 245 32700 312 32734
rect 354 32703 430 32737
rect 346 32700 430 32703
rect 245 32666 430 32700
rect 245 32632 312 32666
rect 346 32665 430 32666
rect 245 32631 320 32632
rect 354 32631 430 32665
rect 245 32598 430 32631
rect 245 32564 312 32598
rect 346 32593 430 32598
rect 245 32559 320 32564
rect 354 32559 430 32593
rect 245 32530 430 32559
rect 245 32496 312 32530
rect 346 32521 430 32530
rect 245 32487 320 32496
rect 354 32487 430 32521
rect 245 32462 430 32487
rect 245 32428 312 32462
rect 346 32449 430 32462
rect 245 32415 320 32428
rect 354 32415 430 32449
rect 245 32394 430 32415
rect 245 32360 312 32394
rect 346 32377 430 32394
rect 245 32343 320 32360
rect 354 32343 430 32377
rect 245 32326 430 32343
rect 245 32292 312 32326
rect 346 32305 430 32326
rect 245 32271 320 32292
rect 354 32271 430 32305
rect 245 32258 430 32271
rect 245 32224 312 32258
rect 346 32233 430 32258
rect 245 32199 320 32224
rect 354 32199 430 32233
rect 245 32190 430 32199
rect 245 32156 312 32190
rect 346 32161 430 32190
rect 245 32127 320 32156
rect 354 32127 430 32161
rect 245 32122 430 32127
rect 245 32088 312 32122
rect 346 32089 430 32122
rect 245 32055 320 32088
rect 354 32055 430 32089
rect 245 32054 430 32055
rect 245 32020 312 32054
rect 346 32020 430 32054
rect 245 32017 430 32020
rect 245 31986 320 32017
rect 245 31952 312 31986
rect 354 31983 430 32017
rect 346 31952 430 31983
rect 245 31945 430 31952
rect 245 31918 320 31945
rect 245 31884 312 31918
rect 354 31911 430 31945
rect 346 31884 430 31911
rect 245 31873 430 31884
rect 245 31850 320 31873
rect 245 31816 312 31850
rect 354 31839 430 31873
rect 346 31816 430 31839
rect 245 31801 430 31816
rect 245 31782 320 31801
rect 245 31748 312 31782
rect 354 31767 430 31801
rect 346 31748 430 31767
rect 245 31729 430 31748
rect 245 31714 320 31729
rect 245 31680 312 31714
rect 354 31695 430 31729
rect 346 31680 430 31695
rect 245 31657 430 31680
rect 245 31646 320 31657
rect 245 31612 312 31646
rect 354 31623 430 31657
rect 346 31612 430 31623
rect 245 31585 430 31612
rect 245 31578 320 31585
rect 245 31544 312 31578
rect 354 31551 430 31585
rect 346 31544 430 31551
rect 245 31513 430 31544
rect 245 31510 320 31513
rect 245 31476 312 31510
rect 354 31479 430 31513
rect 346 31476 430 31479
rect 245 31442 430 31476
rect 245 31408 312 31442
rect 346 31441 430 31442
rect 245 31407 320 31408
rect 354 31407 430 31441
rect 245 31374 430 31407
rect 245 31340 312 31374
rect 346 31369 430 31374
rect 245 31335 320 31340
rect 354 31335 430 31369
rect 245 31306 430 31335
rect 245 31272 312 31306
rect 346 31297 430 31306
rect 245 31263 320 31272
rect 354 31263 430 31297
rect 245 31238 430 31263
rect 245 31204 312 31238
rect 346 31225 430 31238
rect 245 31191 320 31204
rect 354 31191 430 31225
rect 245 31170 430 31191
rect 245 31136 312 31170
rect 346 31153 430 31170
rect 245 31119 320 31136
rect 354 31119 430 31153
rect 245 31102 430 31119
rect 245 31068 312 31102
rect 346 31081 430 31102
rect 245 31047 320 31068
rect 354 31047 430 31081
rect 245 31034 430 31047
rect 245 31000 312 31034
rect 346 31009 430 31034
rect 245 30975 320 31000
rect 354 30975 430 31009
rect 245 30966 430 30975
rect 245 30932 312 30966
rect 346 30937 430 30966
rect 245 30903 320 30932
rect 354 30903 430 30937
rect 245 30898 430 30903
rect 245 30864 312 30898
rect 346 30865 430 30898
rect 245 30831 320 30864
rect 354 30831 430 30865
rect 245 30830 430 30831
rect 245 30796 312 30830
rect 346 30796 430 30830
rect 245 30793 430 30796
rect 245 30762 320 30793
rect 245 30728 312 30762
rect 354 30759 430 30793
rect 346 30728 430 30759
rect 245 30721 430 30728
rect 245 30694 320 30721
rect 245 30660 312 30694
rect 354 30687 430 30721
rect 346 30660 430 30687
rect 245 30649 430 30660
rect 245 30626 320 30649
rect 245 30592 312 30626
rect 354 30615 430 30649
rect 346 30592 430 30615
rect 245 30577 430 30592
rect 245 30558 320 30577
rect 245 30524 312 30558
rect 354 30543 430 30577
rect 346 30524 430 30543
rect 245 30505 430 30524
rect 245 30490 320 30505
rect 245 30456 312 30490
rect 354 30471 430 30505
rect 346 30456 430 30471
rect 245 30433 430 30456
rect 245 30422 320 30433
rect 245 30388 312 30422
rect 354 30399 430 30433
rect 346 30388 430 30399
rect 245 30361 430 30388
rect 245 30354 320 30361
rect 245 30320 312 30354
rect 354 30327 430 30361
rect 346 30320 430 30327
rect 245 30289 430 30320
rect 245 30286 320 30289
rect 245 30252 312 30286
rect 354 30255 430 30289
rect 346 30252 430 30255
rect 245 30218 430 30252
rect 245 30184 312 30218
rect 346 30217 430 30218
rect 245 30183 320 30184
rect 354 30183 430 30217
rect 245 30150 430 30183
rect 245 30116 312 30150
rect 346 30145 430 30150
rect 245 30111 320 30116
rect 354 30111 430 30145
rect 245 30082 430 30111
rect 245 30048 312 30082
rect 346 30073 430 30082
rect 245 30039 320 30048
rect 354 30039 430 30073
rect 245 30014 430 30039
rect 245 29980 312 30014
rect 346 30001 430 30014
rect 245 29967 320 29980
rect 354 29967 430 30001
rect 245 29946 430 29967
rect 245 29912 312 29946
rect 346 29929 430 29946
rect 245 29895 320 29912
rect 354 29895 430 29929
rect 245 29878 430 29895
rect 245 29844 312 29878
rect 346 29857 430 29878
rect 245 29823 320 29844
rect 354 29823 430 29857
rect 245 29810 430 29823
rect 245 29776 312 29810
rect 346 29785 430 29810
rect 245 29751 320 29776
rect 354 29751 430 29785
rect 245 29742 430 29751
rect 245 29708 312 29742
rect 346 29713 430 29742
rect 245 29679 320 29708
rect 354 29679 430 29713
rect 245 29674 430 29679
rect 245 29640 312 29674
rect 346 29641 430 29674
rect 245 29607 320 29640
rect 354 29607 430 29641
rect 245 29606 430 29607
rect 245 29572 312 29606
rect 346 29572 430 29606
rect 245 29569 430 29572
rect 245 29538 320 29569
rect 245 29504 312 29538
rect 354 29535 430 29569
rect 346 29504 430 29535
rect 245 29497 430 29504
rect 245 29470 320 29497
rect 245 29436 312 29470
rect 354 29463 430 29497
rect 346 29436 430 29463
rect 245 29425 430 29436
rect 245 29402 320 29425
rect 245 29368 312 29402
rect 354 29391 430 29425
rect 346 29368 430 29391
rect 245 29353 430 29368
rect 245 29334 320 29353
rect 245 29300 312 29334
rect 354 29319 430 29353
rect 346 29300 430 29319
rect 245 29281 430 29300
rect 245 29266 320 29281
rect 245 29232 312 29266
rect 354 29247 430 29281
rect 346 29232 430 29247
rect 245 29209 430 29232
rect 245 29198 320 29209
rect 245 29164 312 29198
rect 354 29175 430 29209
rect 346 29164 430 29175
rect 245 29137 430 29164
rect 245 29130 320 29137
rect 245 29096 312 29130
rect 354 29103 430 29137
rect 346 29096 430 29103
rect 245 29065 430 29096
rect 245 29062 320 29065
rect 245 29028 312 29062
rect 354 29031 430 29065
rect 346 29028 430 29031
rect 245 28994 430 29028
rect 245 28960 312 28994
rect 346 28993 430 28994
rect 245 28959 320 28960
rect 354 28959 430 28993
rect 245 28926 430 28959
rect 245 28892 312 28926
rect 346 28921 430 28926
rect 245 28887 320 28892
rect 354 28887 430 28921
rect 245 28858 430 28887
rect 245 28824 312 28858
rect 346 28849 430 28858
rect 245 28815 320 28824
rect 354 28815 430 28849
rect 245 28790 430 28815
rect 245 28756 312 28790
rect 346 28777 430 28790
rect 245 28743 320 28756
rect 354 28743 430 28777
rect 245 28722 430 28743
rect 245 28688 312 28722
rect 346 28705 430 28722
rect 245 28671 320 28688
rect 354 28671 430 28705
rect 245 28654 430 28671
rect 245 28620 312 28654
rect 346 28633 430 28654
rect 245 28599 320 28620
rect 354 28599 430 28633
rect 245 28586 430 28599
rect 245 28552 312 28586
rect 346 28561 430 28586
rect 245 28527 320 28552
rect 354 28527 430 28561
rect 245 28518 430 28527
rect 245 28484 312 28518
rect 346 28489 430 28518
rect 245 28455 320 28484
rect 354 28455 430 28489
rect 245 28450 430 28455
rect 245 28416 312 28450
rect 346 28417 430 28450
rect 245 28383 320 28416
rect 354 28383 430 28417
rect 245 28382 430 28383
rect 245 28348 312 28382
rect 346 28348 430 28382
rect 245 28345 430 28348
rect 245 28314 320 28345
rect 245 28280 312 28314
rect 354 28311 430 28345
rect 346 28280 430 28311
rect 245 28273 430 28280
rect 245 28246 320 28273
rect 245 28212 312 28246
rect 354 28239 430 28273
rect 346 28212 430 28239
rect 245 28201 430 28212
rect 245 28178 320 28201
rect 245 28144 312 28178
rect 354 28167 430 28201
rect 346 28144 430 28167
rect 245 28129 430 28144
rect 245 28110 320 28129
rect 245 28076 312 28110
rect 354 28095 430 28129
rect 346 28076 430 28095
rect 245 28057 430 28076
rect 245 28042 320 28057
rect 245 28008 312 28042
rect 354 28023 430 28057
rect 346 28008 430 28023
rect 245 27985 430 28008
rect 245 27974 320 27985
rect 245 27940 312 27974
rect 354 27951 430 27985
rect 346 27940 430 27951
rect 245 27913 430 27940
rect 245 27906 320 27913
rect 245 27872 312 27906
rect 354 27879 430 27913
rect 346 27872 430 27879
rect 245 27841 430 27872
rect 245 27838 320 27841
rect 245 27804 312 27838
rect 354 27807 430 27841
rect 346 27804 430 27807
rect 245 27770 430 27804
rect 245 27736 312 27770
rect 346 27769 430 27770
rect 245 27735 320 27736
rect 354 27735 430 27769
rect 245 27702 430 27735
rect 245 27668 312 27702
rect 346 27697 430 27702
rect 245 27663 320 27668
rect 354 27663 430 27697
rect 245 27634 430 27663
rect 245 27600 312 27634
rect 346 27625 430 27634
rect 245 27591 320 27600
rect 354 27591 430 27625
rect 245 27566 430 27591
rect 245 27532 312 27566
rect 346 27553 430 27566
rect 245 27519 320 27532
rect 354 27519 430 27553
rect 245 27498 430 27519
rect 245 27464 312 27498
rect 346 27481 430 27498
rect 245 27447 320 27464
rect 354 27447 430 27481
rect 245 27430 430 27447
rect 245 27396 312 27430
rect 346 27409 430 27430
rect 245 27375 320 27396
rect 354 27375 430 27409
rect 245 27362 430 27375
rect 245 27328 312 27362
rect 346 27337 430 27362
rect 245 27303 320 27328
rect 354 27303 430 27337
rect 245 27294 430 27303
rect 245 27260 312 27294
rect 346 27265 430 27294
rect 245 27231 320 27260
rect 354 27231 430 27265
rect 245 27226 430 27231
rect 245 27192 312 27226
rect 346 27193 430 27226
rect 245 27159 320 27192
rect 354 27159 430 27193
rect 245 27158 430 27159
rect 245 27124 312 27158
rect 346 27124 430 27158
rect 245 27121 430 27124
rect 245 27090 320 27121
rect 245 27056 312 27090
rect 354 27087 430 27121
rect 346 27056 430 27087
rect 245 27049 430 27056
rect 245 27022 320 27049
rect 245 26988 312 27022
rect 354 27015 430 27049
rect 346 26988 430 27015
rect 245 26977 430 26988
rect 245 26954 320 26977
rect 245 26920 312 26954
rect 354 26943 430 26977
rect 346 26920 430 26943
rect 245 26905 430 26920
rect 245 26886 320 26905
rect 245 26852 312 26886
rect 354 26871 430 26905
rect 346 26852 430 26871
rect 245 26833 430 26852
rect 245 26818 320 26833
rect 245 26784 312 26818
rect 354 26799 430 26833
rect 346 26784 430 26799
rect 245 26761 430 26784
rect 245 26750 320 26761
rect 245 26716 312 26750
rect 354 26727 430 26761
rect 346 26716 430 26727
rect 245 26689 430 26716
rect 245 26682 320 26689
rect 245 26648 312 26682
rect 354 26655 430 26689
rect 346 26648 430 26655
rect 245 26617 430 26648
rect 245 26614 320 26617
rect 245 26580 312 26614
rect 354 26583 430 26617
rect 346 26580 430 26583
rect 245 26546 430 26580
rect 245 26512 312 26546
rect 346 26545 430 26546
rect 245 26511 320 26512
rect 354 26511 430 26545
rect 245 26478 430 26511
rect 245 26444 312 26478
rect 346 26473 430 26478
rect 245 26439 320 26444
rect 354 26439 430 26473
rect 245 26410 430 26439
rect 245 26376 312 26410
rect 346 26401 430 26410
rect 245 26367 320 26376
rect 354 26367 430 26401
rect 245 26342 430 26367
rect 245 26308 312 26342
rect 346 26329 430 26342
rect 245 26295 320 26308
rect 354 26295 430 26329
rect 245 26274 430 26295
rect 245 26240 312 26274
rect 346 26257 430 26274
rect 245 26223 320 26240
rect 354 26223 430 26257
rect 245 26206 430 26223
rect 245 26172 312 26206
rect 346 26185 430 26206
rect 245 26151 320 26172
rect 354 26151 430 26185
rect 245 26138 430 26151
rect 245 26104 312 26138
rect 346 26113 430 26138
rect 245 26079 320 26104
rect 354 26079 430 26113
rect 245 26070 430 26079
rect 245 26036 312 26070
rect 346 26041 430 26070
rect 245 26007 320 26036
rect 354 26007 430 26041
rect 245 26002 430 26007
rect 245 25968 312 26002
rect 346 25969 430 26002
rect 245 25935 320 25968
rect 354 25935 430 25969
rect 245 25934 430 25935
rect 245 25900 312 25934
rect 346 25900 430 25934
rect 245 25897 430 25900
rect 245 25866 320 25897
rect 245 25832 312 25866
rect 354 25863 430 25897
rect 346 25832 430 25863
rect 245 25825 430 25832
rect 245 25798 320 25825
rect 245 25764 312 25798
rect 354 25791 430 25825
rect 346 25764 430 25791
rect 245 25753 430 25764
rect 245 25730 320 25753
rect 245 25696 312 25730
rect 354 25719 430 25753
rect 346 25696 430 25719
rect 245 25681 430 25696
rect 245 25662 320 25681
rect 245 25628 312 25662
rect 354 25647 430 25681
rect 346 25628 430 25647
rect 245 25609 430 25628
rect 245 25594 320 25609
rect 245 25560 312 25594
rect 354 25575 430 25609
rect 346 25560 430 25575
rect 245 25537 430 25560
rect 245 25526 320 25537
rect 245 25492 312 25526
rect 354 25503 430 25537
rect 346 25492 430 25503
rect 245 25465 430 25492
rect 245 25458 320 25465
rect 245 25424 312 25458
rect 354 25431 430 25465
rect 346 25424 430 25431
rect 245 25393 430 25424
rect 245 25390 320 25393
rect 245 25356 312 25390
rect 354 25359 430 25393
rect 346 25356 430 25359
rect 245 25322 430 25356
rect 245 25288 312 25322
rect 346 25321 430 25322
rect 245 25287 320 25288
rect 354 25287 430 25321
rect 245 25254 430 25287
rect 245 25220 312 25254
rect 346 25249 430 25254
rect 245 25215 320 25220
rect 354 25215 430 25249
rect 245 25186 430 25215
rect 245 25152 312 25186
rect 346 25177 430 25186
rect 245 25143 320 25152
rect 354 25143 430 25177
rect 245 25118 430 25143
rect 245 25084 312 25118
rect 346 25105 430 25118
rect 245 25071 320 25084
rect 354 25071 430 25105
rect 245 25050 430 25071
rect 245 25016 312 25050
rect 346 25033 430 25050
rect 245 24999 320 25016
rect 354 24999 430 25033
rect 245 24982 430 24999
rect 245 24948 312 24982
rect 346 24961 430 24982
rect 245 24927 320 24948
rect 354 24927 430 24961
rect 245 24914 430 24927
rect 245 24880 312 24914
rect 346 24889 430 24914
rect 245 24855 320 24880
rect 354 24855 430 24889
rect 245 24846 430 24855
rect 245 24812 312 24846
rect 346 24817 430 24846
rect 245 24783 320 24812
rect 354 24783 430 24817
rect 245 24778 430 24783
rect 245 24744 312 24778
rect 346 24745 430 24778
rect 245 24711 320 24744
rect 354 24711 430 24745
rect 245 24710 430 24711
rect 245 24676 312 24710
rect 346 24676 430 24710
rect 245 24673 430 24676
rect 245 24642 320 24673
rect 245 24608 312 24642
rect 354 24639 430 24673
rect 346 24608 430 24639
rect 245 24601 430 24608
rect 245 24574 320 24601
rect 245 24540 312 24574
rect 354 24567 430 24601
rect 346 24540 430 24567
rect 245 24529 430 24540
rect 245 24506 320 24529
rect 245 24472 312 24506
rect 354 24495 430 24529
rect 346 24472 430 24495
rect 245 24457 430 24472
rect 245 24438 320 24457
rect 245 24404 312 24438
rect 354 24423 430 24457
rect 346 24404 430 24423
rect 245 24385 430 24404
rect 245 24370 320 24385
rect 245 24336 312 24370
rect 354 24351 430 24385
rect 346 24336 430 24351
rect 245 24313 430 24336
rect 245 24302 320 24313
rect 245 24268 312 24302
rect 354 24279 430 24313
rect 346 24268 430 24279
rect 245 24241 430 24268
rect 245 24234 320 24241
rect 245 24200 312 24234
rect 354 24207 430 24241
rect 346 24200 430 24207
rect 245 24169 430 24200
rect 245 24166 320 24169
rect 245 24132 312 24166
rect 354 24135 430 24169
rect 346 24132 430 24135
rect 245 24098 430 24132
rect 245 24064 312 24098
rect 346 24097 430 24098
rect 245 24063 320 24064
rect 354 24063 430 24097
rect 245 24030 430 24063
rect 245 23996 312 24030
rect 346 24025 430 24030
rect 245 23991 320 23996
rect 354 23991 430 24025
rect 245 23962 430 23991
rect 245 23928 312 23962
rect 346 23953 430 23962
rect 245 23919 320 23928
rect 354 23919 430 23953
rect 245 23894 430 23919
rect 245 23860 312 23894
rect 346 23881 430 23894
rect 245 23847 320 23860
rect 354 23847 430 23881
rect 245 23826 430 23847
rect 245 23792 312 23826
rect 346 23809 430 23826
rect 245 23775 320 23792
rect 354 23775 430 23809
rect 245 23758 430 23775
rect 245 23724 312 23758
rect 346 23737 430 23758
rect 245 23703 320 23724
rect 354 23703 430 23737
rect 245 23690 430 23703
rect 245 23656 312 23690
rect 346 23665 430 23690
rect 245 23631 320 23656
rect 354 23631 430 23665
rect 245 23622 430 23631
rect 245 23588 312 23622
rect 346 23593 430 23622
rect 245 23559 320 23588
rect 354 23559 430 23593
rect 245 23554 430 23559
rect 245 23520 312 23554
rect 346 23521 430 23554
rect 245 23487 320 23520
rect 354 23487 430 23521
rect 245 23486 430 23487
rect 245 23452 312 23486
rect 346 23452 430 23486
rect 245 23449 430 23452
rect 245 23418 320 23449
rect 245 23384 312 23418
rect 354 23415 430 23449
rect 346 23384 430 23415
rect 245 23377 430 23384
rect 245 23350 320 23377
rect 245 23316 312 23350
rect 354 23343 430 23377
rect 346 23316 430 23343
rect 245 23305 430 23316
rect 245 23282 320 23305
rect 245 23248 312 23282
rect 354 23271 430 23305
rect 346 23248 430 23271
rect 245 23233 430 23248
rect 245 23214 320 23233
rect 245 23180 312 23214
rect 354 23199 430 23233
rect 346 23180 430 23199
rect 245 23161 430 23180
rect 245 23146 320 23161
rect 245 23112 312 23146
rect 354 23127 430 23161
rect 346 23112 430 23127
rect 245 23089 430 23112
rect 245 23078 320 23089
rect 245 23044 312 23078
rect 354 23055 430 23089
rect 346 23044 430 23055
rect 245 23017 430 23044
rect 245 23010 320 23017
rect 245 22976 312 23010
rect 354 22983 430 23017
rect 346 22976 430 22983
rect 245 22945 430 22976
rect 245 22942 320 22945
rect 245 22908 312 22942
rect 354 22911 430 22945
rect 346 22908 430 22911
rect 245 22874 430 22908
rect 245 22840 312 22874
rect 346 22873 430 22874
rect 245 22839 320 22840
rect 354 22839 430 22873
rect 245 22806 430 22839
rect 245 22772 312 22806
rect 346 22801 430 22806
rect 245 22767 320 22772
rect 354 22767 430 22801
rect 245 22738 430 22767
rect 245 22704 312 22738
rect 346 22729 430 22738
rect 245 22695 320 22704
rect 354 22695 430 22729
rect 245 22670 430 22695
rect 245 22636 312 22670
rect 346 22657 430 22670
rect 245 22623 320 22636
rect 354 22623 430 22657
rect 245 22602 430 22623
rect 245 22568 312 22602
rect 346 22585 430 22602
rect 245 22551 320 22568
rect 354 22551 430 22585
rect 245 22534 430 22551
rect 245 22500 312 22534
rect 346 22513 430 22534
rect 245 22479 320 22500
rect 354 22479 430 22513
rect 245 22466 430 22479
rect 245 22432 312 22466
rect 346 22441 430 22466
rect 245 22407 320 22432
rect 354 22407 430 22441
rect 245 22398 430 22407
rect 245 22364 312 22398
rect 346 22369 430 22398
rect 245 22335 320 22364
rect 354 22335 430 22369
rect 245 22330 430 22335
rect 245 22296 312 22330
rect 346 22297 430 22330
rect 245 22263 320 22296
rect 354 22263 430 22297
rect 245 22262 430 22263
rect 245 22228 312 22262
rect 346 22228 430 22262
rect 245 22225 430 22228
rect 245 22194 320 22225
rect 245 22160 312 22194
rect 354 22191 430 22225
rect 346 22160 430 22191
rect 245 22153 430 22160
rect 245 22126 320 22153
rect 245 22092 312 22126
rect 354 22119 430 22153
rect 346 22092 430 22119
rect 245 22081 430 22092
rect 245 22058 320 22081
rect 245 22024 312 22058
rect 354 22047 430 22081
rect 346 22024 430 22047
rect 245 22009 430 22024
rect 245 21990 320 22009
rect 245 21956 312 21990
rect 354 21975 430 22009
rect 346 21956 430 21975
rect 245 21937 430 21956
rect 245 21922 320 21937
rect 245 21888 312 21922
rect 354 21903 430 21937
rect 346 21888 430 21903
rect 245 21865 430 21888
rect 245 21854 320 21865
rect 245 21820 312 21854
rect 354 21831 430 21865
rect 346 21820 430 21831
rect 245 21793 430 21820
rect 245 21786 320 21793
rect 245 21752 312 21786
rect 354 21759 430 21793
rect 346 21752 430 21759
rect 245 21721 430 21752
rect 245 21718 320 21721
rect 245 21684 312 21718
rect 354 21687 430 21721
rect 346 21684 430 21687
rect 245 21650 430 21684
rect 245 21616 312 21650
rect 346 21649 430 21650
rect 245 21615 320 21616
rect 354 21615 430 21649
rect 245 21582 430 21615
rect 245 21548 312 21582
rect 346 21577 430 21582
rect 245 21543 320 21548
rect 354 21543 430 21577
rect 245 21514 430 21543
rect 245 21480 312 21514
rect 346 21505 430 21514
rect 245 21471 320 21480
rect 354 21471 430 21505
rect 245 21446 430 21471
rect 245 21412 312 21446
rect 346 21433 430 21446
rect 245 21399 320 21412
rect 354 21399 430 21433
rect 245 21378 430 21399
rect 245 21344 312 21378
rect 346 21361 430 21378
rect 245 21327 320 21344
rect 354 21327 430 21361
rect 245 21310 430 21327
rect 245 21276 312 21310
rect 346 21289 430 21310
rect 245 21255 320 21276
rect 354 21255 430 21289
rect 245 21242 430 21255
rect 245 21208 312 21242
rect 346 21217 430 21242
rect 245 21183 320 21208
rect 354 21183 430 21217
rect 245 21174 430 21183
rect 245 21140 312 21174
rect 346 21145 430 21174
rect 245 21111 320 21140
rect 354 21111 430 21145
rect 245 21106 430 21111
rect 245 21072 312 21106
rect 346 21073 430 21106
rect 245 21039 320 21072
rect 354 21039 430 21073
rect 245 21038 430 21039
rect 245 21004 312 21038
rect 346 21004 430 21038
rect 245 21001 430 21004
rect 245 20970 320 21001
rect 245 20936 312 20970
rect 354 20967 430 21001
rect 346 20936 430 20967
rect 245 20929 430 20936
rect 245 20902 320 20929
rect 245 20868 312 20902
rect 354 20895 430 20929
rect 346 20868 430 20895
rect 245 20857 430 20868
rect 245 20834 320 20857
rect 245 20800 312 20834
rect 354 20823 430 20857
rect 346 20800 430 20823
rect 245 20785 430 20800
rect 245 20766 320 20785
rect 245 20732 312 20766
rect 354 20751 430 20785
rect 346 20732 430 20751
rect 245 20713 430 20732
rect 245 20698 320 20713
rect 245 20664 312 20698
rect 354 20679 430 20713
rect 346 20664 430 20679
rect 245 20641 430 20664
rect 245 20630 320 20641
rect 245 20596 312 20630
rect 354 20607 430 20641
rect 346 20596 430 20607
rect 245 20569 430 20596
rect 245 20562 320 20569
rect 245 20528 312 20562
rect 354 20535 430 20569
rect 346 20528 430 20535
rect 245 20497 430 20528
rect 245 20494 320 20497
rect 245 20460 312 20494
rect 354 20463 430 20497
rect 346 20460 430 20463
rect 245 20426 430 20460
rect 245 20392 312 20426
rect 346 20425 430 20426
rect 245 20391 320 20392
rect 354 20391 430 20425
rect 245 20358 430 20391
rect 245 20324 312 20358
rect 346 20353 430 20358
rect 245 20319 320 20324
rect 354 20319 430 20353
rect 245 20290 430 20319
rect 245 20256 312 20290
rect 346 20281 430 20290
rect 245 20247 320 20256
rect 354 20247 430 20281
rect 245 20222 430 20247
rect 245 20188 312 20222
rect 346 20209 430 20222
rect 245 20175 320 20188
rect 354 20175 430 20209
rect 245 20154 430 20175
rect 245 20120 312 20154
rect 346 20137 430 20154
rect 245 20103 320 20120
rect 354 20103 430 20137
rect 245 20086 430 20103
rect 245 20052 312 20086
rect 346 20065 430 20086
rect 245 20031 320 20052
rect 354 20031 430 20065
rect 245 20018 430 20031
rect 245 19984 312 20018
rect 346 19993 430 20018
rect 245 19959 320 19984
rect 354 19959 430 19993
rect 245 19950 430 19959
rect 245 19916 312 19950
rect 346 19921 430 19950
rect 245 19887 320 19916
rect 354 19887 430 19921
rect 245 19882 430 19887
rect 245 19848 312 19882
rect 346 19849 430 19882
rect 245 19815 320 19848
rect 354 19815 430 19849
rect 245 19814 430 19815
rect 245 19780 312 19814
rect 346 19780 430 19814
rect 245 19777 430 19780
rect 245 19746 320 19777
rect 245 19712 312 19746
rect 354 19743 430 19777
rect 346 19712 430 19743
rect 245 19705 430 19712
rect 245 19678 320 19705
rect 245 19644 312 19678
rect 354 19671 430 19705
rect 346 19644 430 19671
rect 245 19633 430 19644
rect 245 19610 320 19633
rect 245 19576 312 19610
rect 354 19599 430 19633
rect 346 19576 430 19599
rect 245 19561 430 19576
rect 245 19542 320 19561
rect 245 19508 312 19542
rect 354 19527 430 19561
rect 346 19508 430 19527
rect 245 19489 430 19508
rect 245 19474 320 19489
rect 245 19440 312 19474
rect 354 19455 430 19489
rect 346 19440 430 19455
rect 245 19417 430 19440
rect 245 19406 320 19417
rect 245 19372 312 19406
rect 354 19383 430 19417
rect 346 19372 430 19383
rect 245 19345 430 19372
rect 245 19338 320 19345
rect 245 19304 312 19338
rect 354 19311 430 19345
rect 346 19304 430 19311
rect 245 19273 430 19304
rect 245 19270 320 19273
rect 245 19236 312 19270
rect 354 19239 430 19273
rect 346 19236 430 19239
rect 245 19202 430 19236
rect 245 19168 312 19202
rect 346 19201 430 19202
rect 245 19167 320 19168
rect 354 19167 430 19201
rect 245 19134 430 19167
rect 245 19100 312 19134
rect 346 19129 430 19134
rect 245 19095 320 19100
rect 354 19095 430 19129
rect 245 19066 430 19095
rect 245 19032 312 19066
rect 346 19057 430 19066
rect 245 19023 320 19032
rect 354 19023 430 19057
rect 245 18998 430 19023
rect 245 18964 312 18998
rect 346 18985 430 18998
rect 245 18951 320 18964
rect 354 18951 430 18985
rect 245 18930 430 18951
rect 245 18896 312 18930
rect 346 18913 430 18930
rect 245 18879 320 18896
rect 354 18879 430 18913
rect 245 18862 430 18879
rect 245 18828 312 18862
rect 346 18841 430 18862
rect 245 18807 320 18828
rect 354 18807 430 18841
rect 245 18794 430 18807
rect 245 18760 312 18794
rect 346 18769 430 18794
rect 245 18735 320 18760
rect 354 18735 430 18769
rect 245 18726 430 18735
rect 245 18692 312 18726
rect 346 18697 430 18726
rect 245 18663 320 18692
rect 354 18663 430 18697
rect 245 18658 430 18663
rect 245 18624 312 18658
rect 346 18625 430 18658
rect 245 18591 320 18624
rect 354 18591 430 18625
rect 245 18590 430 18591
rect 245 18556 312 18590
rect 346 18556 430 18590
rect 245 18553 430 18556
rect 245 18522 320 18553
rect 245 18488 312 18522
rect 354 18519 430 18553
rect 346 18488 430 18519
rect 245 18481 430 18488
rect 245 18454 320 18481
rect 245 18420 312 18454
rect 354 18447 430 18481
rect 346 18420 430 18447
rect 245 18409 430 18420
rect 245 18386 320 18409
rect 245 18352 312 18386
rect 354 18375 430 18409
rect 346 18352 430 18375
rect 245 18337 430 18352
rect 245 18318 320 18337
rect 245 18284 312 18318
rect 354 18303 430 18337
rect 346 18284 430 18303
rect 245 18265 430 18284
rect 245 18250 320 18265
rect 245 18216 312 18250
rect 354 18231 430 18265
rect 346 18216 430 18231
rect 245 18193 430 18216
rect 245 18182 320 18193
rect 245 18148 312 18182
rect 354 18159 430 18193
rect 346 18148 430 18159
rect 245 18121 430 18148
rect 245 18114 320 18121
rect 245 18080 312 18114
rect 354 18087 430 18121
rect 346 18080 430 18087
rect 245 18049 430 18080
rect 245 18046 320 18049
rect 245 18012 312 18046
rect 354 18015 430 18049
rect 346 18012 430 18015
rect 245 17978 430 18012
rect 245 17944 312 17978
rect 346 17977 430 17978
rect 245 17943 320 17944
rect 354 17943 430 17977
rect 245 17910 430 17943
rect 245 17876 312 17910
rect 346 17905 430 17910
rect 245 17871 320 17876
rect 354 17871 430 17905
rect 245 17842 430 17871
rect 245 17808 312 17842
rect 346 17833 430 17842
rect 245 17799 320 17808
rect 354 17799 430 17833
rect 245 17774 430 17799
rect 245 17740 312 17774
rect 346 17761 430 17774
rect 245 17727 320 17740
rect 354 17727 430 17761
rect 245 17706 430 17727
rect 245 17672 312 17706
rect 346 17689 430 17706
rect 245 17655 320 17672
rect 354 17655 430 17689
rect 245 17638 430 17655
rect 245 17604 312 17638
rect 346 17617 430 17638
rect 245 17583 320 17604
rect 354 17583 430 17617
rect 245 17570 430 17583
rect 245 17536 312 17570
rect 346 17545 430 17570
rect 245 17511 320 17536
rect 354 17511 430 17545
rect 245 17502 430 17511
rect 245 17468 312 17502
rect 346 17473 430 17502
rect 245 17439 320 17468
rect 354 17439 430 17473
rect 245 17434 430 17439
rect 245 17400 312 17434
rect 346 17401 430 17434
rect 245 17367 320 17400
rect 354 17367 430 17401
rect 245 17366 430 17367
rect 245 17332 312 17366
rect 346 17332 430 17366
rect 245 17329 430 17332
rect 245 17298 320 17329
rect 245 17264 312 17298
rect 354 17295 430 17329
rect 346 17264 430 17295
rect 245 17257 430 17264
rect 245 17230 320 17257
rect 245 17196 312 17230
rect 354 17223 430 17257
rect 346 17196 430 17223
rect 245 17185 430 17196
rect 245 17162 320 17185
rect 245 17128 312 17162
rect 354 17151 430 17185
rect 346 17128 430 17151
rect 245 17113 430 17128
rect 245 17094 320 17113
rect 245 17060 312 17094
rect 354 17079 430 17113
rect 346 17060 430 17079
rect 245 17041 430 17060
rect 245 17026 320 17041
rect 245 16992 312 17026
rect 354 17007 430 17041
rect 346 16992 430 17007
rect 245 16969 430 16992
rect 245 16958 320 16969
rect 245 16924 312 16958
rect 354 16935 430 16969
rect 346 16924 430 16935
rect 245 16897 430 16924
rect 245 16890 320 16897
rect 245 16856 312 16890
rect 354 16863 430 16897
rect 346 16856 430 16863
rect 245 16825 430 16856
rect 245 16822 320 16825
rect 245 16788 312 16822
rect 354 16791 430 16825
rect 346 16788 430 16791
rect 245 16754 430 16788
rect 245 16720 312 16754
rect 346 16753 430 16754
rect 245 16719 320 16720
rect 354 16719 430 16753
rect 245 16686 430 16719
rect 245 16652 312 16686
rect 346 16681 430 16686
rect 245 16647 320 16652
rect 354 16647 430 16681
rect 245 16618 430 16647
rect 245 16584 312 16618
rect 346 16609 430 16618
rect 245 16575 320 16584
rect 354 16575 430 16609
rect 245 16550 430 16575
rect 245 16516 312 16550
rect 346 16537 430 16550
rect 245 16503 320 16516
rect 354 16503 430 16537
rect 245 16482 430 16503
rect 245 16448 312 16482
rect 346 16465 430 16482
rect 245 16431 320 16448
rect 354 16431 430 16465
rect 245 16414 430 16431
rect 245 16380 312 16414
rect 346 16393 430 16414
rect 245 16359 320 16380
rect 354 16359 430 16393
rect 245 16346 430 16359
rect 245 16312 312 16346
rect 346 16321 430 16346
rect 245 16287 320 16312
rect 354 16287 430 16321
rect 245 16278 430 16287
rect 245 16244 312 16278
rect 346 16249 430 16278
rect 245 16215 320 16244
rect 354 16215 430 16249
rect 245 16210 430 16215
rect 245 16176 312 16210
rect 346 16177 430 16210
rect 245 16143 320 16176
rect 354 16143 430 16177
rect 245 16142 430 16143
rect 245 16108 312 16142
rect 346 16108 430 16142
rect 245 16105 430 16108
rect 245 16074 320 16105
rect 245 16040 312 16074
rect 354 16071 430 16105
rect 346 16040 430 16071
rect 245 16033 430 16040
rect 245 16006 320 16033
rect 245 15972 312 16006
rect 354 15999 430 16033
rect 346 15972 430 15999
rect 245 15961 430 15972
rect 245 15938 320 15961
rect 245 15904 312 15938
rect 354 15927 430 15961
rect 346 15904 430 15927
rect 245 15889 430 15904
rect 245 15870 320 15889
rect 245 15836 312 15870
rect 354 15855 430 15889
rect 346 15836 430 15855
rect 245 15817 430 15836
rect 245 15802 320 15817
rect 245 15768 312 15802
rect 354 15783 430 15817
rect 346 15768 430 15783
rect 245 15745 430 15768
rect 245 15734 320 15745
rect 245 15700 312 15734
rect 354 15711 430 15745
rect 346 15700 430 15711
rect 245 15673 430 15700
rect 245 15666 320 15673
rect 245 15632 312 15666
rect 354 15639 430 15673
rect 346 15632 430 15639
rect 245 15601 430 15632
rect 245 15598 320 15601
rect 245 15564 312 15598
rect 354 15567 430 15601
rect 346 15564 430 15567
rect 245 15530 430 15564
rect 245 15496 312 15530
rect 346 15529 430 15530
rect 245 15495 320 15496
rect 354 15495 430 15529
rect 245 15462 430 15495
rect 245 15428 312 15462
rect 346 15457 430 15462
rect 245 15423 320 15428
rect 354 15423 430 15457
rect 245 15394 430 15423
rect 245 15360 312 15394
rect 346 15385 430 15394
rect 245 15351 320 15360
rect 354 15351 430 15385
rect 245 15326 430 15351
rect 245 15292 312 15326
rect 346 15313 430 15326
rect 245 15279 320 15292
rect 354 15279 430 15313
rect 245 15258 430 15279
rect 245 15224 312 15258
rect 346 15241 430 15258
rect 245 15207 320 15224
rect 354 15207 430 15241
rect 245 15190 430 15207
rect 245 15156 312 15190
rect 346 15169 430 15190
rect 245 15135 320 15156
rect 354 15135 430 15169
rect 245 15122 430 15135
rect 245 15088 312 15122
rect 346 15097 430 15122
rect 245 15063 320 15088
rect 354 15063 430 15097
rect 245 15054 430 15063
rect 245 15020 312 15054
rect 346 15025 430 15054
rect 245 14991 320 15020
rect 354 14991 430 15025
rect 245 14986 430 14991
rect 245 14952 312 14986
rect 346 14953 430 14986
rect 245 14919 320 14952
rect 354 14919 430 14953
rect 245 14918 430 14919
rect 245 14884 312 14918
rect 346 14884 430 14918
rect 245 14881 430 14884
rect 245 14850 320 14881
rect 245 14816 312 14850
rect 354 14847 430 14881
rect 346 14816 430 14847
rect 245 14809 430 14816
rect 245 14782 320 14809
rect 245 14748 312 14782
rect 354 14775 430 14809
rect 346 14748 430 14775
rect 245 14737 430 14748
rect 245 14714 320 14737
rect 245 14680 312 14714
rect 354 14703 430 14737
rect 346 14680 430 14703
rect 245 14665 430 14680
rect 245 14646 320 14665
rect 245 14612 312 14646
rect 354 14631 430 14665
rect 346 14612 430 14631
rect 245 14593 430 14612
rect 245 14578 320 14593
rect 245 14544 312 14578
rect 354 14559 430 14593
rect 346 14544 430 14559
rect 245 14521 430 14544
rect 245 14510 320 14521
rect 245 14476 312 14510
rect 354 14487 430 14521
rect 346 14476 430 14487
rect 245 14449 430 14476
rect 245 14442 320 14449
rect 245 14408 312 14442
rect 354 14415 430 14449
rect 346 14408 430 14415
rect 245 14377 430 14408
rect 245 14374 320 14377
rect 245 14340 312 14374
rect 354 14343 430 14377
rect 346 14340 430 14343
rect 245 14306 430 14340
rect 245 14272 312 14306
rect 346 14305 430 14306
rect 245 14271 320 14272
rect 354 14271 430 14305
rect 245 14238 430 14271
rect 245 14204 312 14238
rect 346 14233 430 14238
rect 245 14199 320 14204
rect 354 14199 430 14233
rect 245 14170 430 14199
rect 245 14136 312 14170
rect 346 14161 430 14170
rect 245 14127 320 14136
rect 354 14127 430 14161
rect 245 14102 430 14127
rect 245 14068 312 14102
rect 346 14089 430 14102
rect 245 14055 320 14068
rect 354 14055 430 14089
rect 245 14034 430 14055
rect 245 14000 312 14034
rect 346 14017 430 14034
rect 245 13983 320 14000
rect 354 13983 430 14017
rect 245 13966 430 13983
rect 245 13932 312 13966
rect 346 13945 430 13966
rect 245 13911 320 13932
rect 354 13911 430 13945
rect 245 13898 430 13911
rect 245 13864 312 13898
rect 346 13873 430 13898
rect 245 13839 320 13864
rect 354 13839 430 13873
rect 245 13830 430 13839
rect 245 13796 312 13830
rect 346 13801 430 13830
rect 245 13767 320 13796
rect 354 13767 430 13801
rect 245 13762 430 13767
rect 245 13728 312 13762
rect 346 13729 430 13762
rect 245 13695 320 13728
rect 354 13695 430 13729
rect 245 13694 430 13695
rect 245 13660 312 13694
rect 346 13660 430 13694
rect 245 13657 430 13660
rect 245 13626 320 13657
rect 245 13592 312 13626
rect 354 13623 430 13657
rect 346 13592 430 13623
rect 245 13585 430 13592
rect 245 13558 320 13585
rect 245 13524 312 13558
rect 354 13551 430 13585
rect 346 13524 430 13551
rect 245 13513 430 13524
rect 245 13490 320 13513
rect 245 13456 312 13490
rect 354 13479 430 13513
rect 346 13456 430 13479
rect 245 13441 430 13456
rect 245 13422 320 13441
rect 245 13388 312 13422
rect 354 13407 430 13441
rect 346 13388 430 13407
rect 245 13369 430 13388
rect 245 13354 320 13369
rect 245 13320 312 13354
rect 354 13335 430 13369
rect 346 13320 430 13335
rect 245 13297 430 13320
rect 245 13286 320 13297
rect 245 13252 312 13286
rect 354 13263 430 13297
rect 346 13252 430 13263
rect 245 13225 430 13252
rect 245 13218 320 13225
rect 245 13184 312 13218
rect 354 13191 430 13225
rect 346 13184 430 13191
rect 245 13153 430 13184
rect 245 13150 320 13153
rect 245 13116 312 13150
rect 354 13119 430 13153
rect 346 13116 430 13119
rect 245 13082 430 13116
rect 245 13048 312 13082
rect 346 13081 430 13082
rect 245 13047 320 13048
rect 354 13047 430 13081
rect 245 13014 430 13047
rect 245 12980 312 13014
rect 346 13009 430 13014
rect 245 12975 320 12980
rect 354 12975 430 13009
rect 245 12946 430 12975
rect 245 12912 312 12946
rect 346 12937 430 12946
rect 245 12903 320 12912
rect 354 12903 430 12937
rect 245 12878 430 12903
rect 245 12844 312 12878
rect 346 12865 430 12878
rect 245 12831 320 12844
rect 354 12831 430 12865
rect 245 12810 430 12831
rect 245 12776 312 12810
rect 346 12793 430 12810
rect 245 12759 320 12776
rect 354 12759 430 12793
rect 245 12742 430 12759
rect 245 12708 312 12742
rect 346 12721 430 12742
rect 245 12687 320 12708
rect 354 12687 430 12721
rect 245 12674 430 12687
rect 245 12640 312 12674
rect 346 12649 430 12674
rect 245 12615 320 12640
rect 354 12615 430 12649
rect 245 12606 430 12615
rect 245 12572 312 12606
rect 346 12577 430 12606
rect 245 12543 320 12572
rect 354 12543 430 12577
rect 245 12538 430 12543
rect 245 12504 312 12538
rect 346 12505 430 12538
rect 245 12471 320 12504
rect 354 12471 430 12505
rect 245 12470 430 12471
rect 245 12436 312 12470
rect 346 12436 430 12470
rect 245 12433 430 12436
rect 245 12402 320 12433
rect 245 12368 312 12402
rect 354 12399 430 12433
rect 346 12368 430 12399
rect 245 12361 430 12368
rect 245 12334 320 12361
rect 245 12300 312 12334
rect 354 12327 430 12361
rect 346 12300 430 12327
rect 245 12289 430 12300
rect 245 12266 320 12289
rect 245 12232 312 12266
rect 354 12255 430 12289
rect 346 12232 430 12255
rect 245 12217 430 12232
rect 245 12198 320 12217
rect 245 12164 312 12198
rect 354 12183 430 12217
rect 346 12164 430 12183
rect 245 12145 430 12164
rect 245 12130 320 12145
rect 245 12096 312 12130
rect 354 12111 430 12145
rect 346 12096 430 12111
rect 245 12073 430 12096
rect 245 12062 320 12073
rect 245 12028 312 12062
rect 354 12039 430 12073
rect 346 12028 430 12039
rect 245 12001 430 12028
rect 245 11994 320 12001
rect 245 11960 312 11994
rect 354 11967 430 12001
rect 346 11960 430 11967
rect 245 11929 430 11960
rect 245 11926 320 11929
rect 245 11892 312 11926
rect 354 11895 430 11929
rect 346 11892 430 11895
rect 245 11858 430 11892
rect 245 11824 312 11858
rect 346 11857 430 11858
rect 245 11823 320 11824
rect 354 11823 430 11857
rect 245 11790 430 11823
rect 245 11756 312 11790
rect 346 11785 430 11790
rect 245 11751 320 11756
rect 354 11751 430 11785
rect 245 11722 430 11751
rect 245 11688 312 11722
rect 346 11713 430 11722
rect 245 11679 320 11688
rect 354 11679 430 11713
rect 245 11654 430 11679
rect 245 11620 312 11654
rect 346 11641 430 11654
rect 245 11607 320 11620
rect 354 11607 430 11641
rect 245 11586 430 11607
rect 245 11552 312 11586
rect 346 11569 430 11586
rect 245 11535 320 11552
rect 354 11535 430 11569
rect 245 11518 430 11535
rect 245 11484 312 11518
rect 346 11497 430 11518
rect 245 11463 320 11484
rect 354 11463 430 11497
rect 245 11450 430 11463
rect 245 11416 312 11450
rect 346 11425 430 11450
rect 245 11391 320 11416
rect 354 11391 430 11425
rect 245 11382 430 11391
rect 245 11348 312 11382
rect 346 11353 430 11382
rect 245 11319 320 11348
rect 354 11319 430 11353
rect 245 11314 430 11319
rect 245 11280 312 11314
rect 346 11281 430 11314
rect 245 11247 320 11280
rect 354 11247 430 11281
rect 245 11246 430 11247
rect 245 11212 312 11246
rect 346 11212 430 11246
rect 245 11209 430 11212
rect 245 11178 320 11209
rect 245 11144 312 11178
rect 354 11175 430 11209
rect 346 11144 430 11175
rect 245 11137 430 11144
rect 245 11110 320 11137
rect 245 11076 312 11110
rect 354 11103 430 11137
rect 346 11076 430 11103
rect 245 11065 430 11076
rect 245 11042 320 11065
rect 245 11008 312 11042
rect 354 11031 430 11065
rect 346 11008 430 11031
rect 245 10993 430 11008
rect 245 10974 320 10993
rect 245 10940 312 10974
rect 354 10959 430 10993
rect 346 10940 430 10959
rect 245 10921 430 10940
rect 245 10906 320 10921
rect 245 10872 312 10906
rect 354 10887 430 10921
rect 346 10872 430 10887
rect 245 10849 430 10872
rect 245 10838 320 10849
rect 245 10804 312 10838
rect 354 10815 430 10849
rect 346 10804 430 10815
rect 245 10777 430 10804
rect 245 10770 320 10777
rect 245 10736 312 10770
rect 354 10743 430 10777
rect 346 10736 430 10743
rect 245 10705 430 10736
rect 245 10702 320 10705
rect 245 10668 312 10702
rect 354 10671 430 10705
rect 346 10668 430 10671
rect 245 10634 430 10668
rect 245 10600 312 10634
rect 346 10633 430 10634
rect 245 10599 320 10600
rect 354 10599 430 10633
rect 245 10566 430 10599
rect 245 10532 312 10566
rect 346 10561 430 10566
rect 245 10527 320 10532
rect 354 10527 430 10561
rect 245 10498 430 10527
rect 245 10464 312 10498
rect 346 10489 430 10498
rect 245 10455 320 10464
rect 354 10455 430 10489
rect 245 10430 430 10455
rect 245 10396 312 10430
rect 346 10417 430 10430
rect 245 10383 320 10396
rect 354 10383 430 10417
rect 245 10362 430 10383
rect 245 10328 312 10362
rect 346 10345 430 10362
rect 245 10311 320 10328
rect 354 10311 430 10345
rect 245 10294 430 10311
rect 245 10260 312 10294
rect 346 10273 430 10294
rect 245 10239 320 10260
rect 354 10239 430 10273
rect 245 10226 430 10239
rect 245 10192 312 10226
rect 346 10201 430 10226
rect 245 10167 320 10192
rect 354 10167 430 10201
rect 245 10158 430 10167
rect 245 10124 312 10158
rect 346 10129 430 10158
rect 245 10095 320 10124
rect 354 10095 430 10129
rect 245 10090 430 10095
rect 245 10056 312 10090
rect 346 10057 430 10090
rect 245 10023 320 10056
rect 354 10023 430 10057
rect 245 10022 430 10023
rect 245 9988 312 10022
rect 346 9988 430 10022
rect 245 9985 430 9988
rect 245 9954 320 9985
rect 245 9920 312 9954
rect 354 9951 430 9985
rect 346 9920 430 9951
rect 245 9913 430 9920
rect 245 9886 320 9913
rect 245 9852 312 9886
rect 354 9879 430 9913
rect 346 9852 430 9879
rect 245 9841 430 9852
rect 245 9818 320 9841
rect 245 9784 312 9818
rect 354 9807 430 9841
rect 346 9784 430 9807
rect 245 9769 430 9784
rect 245 9750 320 9769
rect 245 9716 312 9750
rect 354 9735 430 9769
rect 346 9716 430 9735
rect 245 9697 430 9716
rect 603 36177 14361 36207
rect 603 36143 766 36177
rect 800 36143 834 36177
rect 868 36143 902 36177
rect 936 36143 970 36177
rect 1004 36143 1038 36177
rect 1072 36143 1106 36177
rect 1140 36143 1174 36177
rect 1208 36143 1242 36177
rect 1276 36143 1310 36177
rect 1344 36143 1378 36177
rect 1412 36143 1446 36177
rect 1480 36143 1514 36177
rect 1548 36143 1582 36177
rect 1616 36143 1650 36177
rect 1684 36143 1718 36177
rect 1752 36143 1786 36177
rect 1820 36143 1854 36177
rect 1888 36143 1922 36177
rect 1956 36143 1990 36177
rect 2024 36143 2058 36177
rect 2092 36143 2126 36177
rect 2160 36143 2194 36177
rect 2228 36143 2262 36177
rect 2296 36143 2330 36177
rect 2364 36143 2398 36177
rect 2432 36143 2466 36177
rect 2500 36143 2534 36177
rect 2568 36143 2602 36177
rect 2636 36143 2670 36177
rect 2704 36143 2738 36177
rect 2772 36143 2806 36177
rect 2840 36143 2874 36177
rect 2908 36143 2942 36177
rect 2976 36143 3010 36177
rect 3044 36143 3078 36177
rect 3112 36143 3146 36177
rect 3180 36143 3214 36177
rect 3248 36143 3282 36177
rect 3316 36143 3350 36177
rect 3384 36143 3418 36177
rect 3452 36143 3486 36177
rect 3520 36143 3554 36177
rect 3588 36143 3622 36177
rect 3656 36143 3690 36177
rect 3724 36143 3758 36177
rect 3792 36143 3826 36177
rect 3860 36143 3894 36177
rect 3928 36143 3962 36177
rect 3996 36143 4030 36177
rect 4064 36143 4098 36177
rect 4132 36143 4166 36177
rect 4200 36143 4234 36177
rect 4268 36143 4302 36177
rect 4336 36143 4370 36177
rect 4404 36143 4438 36177
rect 4472 36143 4506 36177
rect 4540 36143 4574 36177
rect 4608 36143 4642 36177
rect 4676 36143 4710 36177
rect 4744 36143 4778 36177
rect 4812 36143 4846 36177
rect 4880 36143 4914 36177
rect 4948 36143 4982 36177
rect 5016 36143 5050 36177
rect 5084 36143 5118 36177
rect 5152 36143 5186 36177
rect 5220 36143 5254 36177
rect 5288 36143 5322 36177
rect 5356 36143 5390 36177
rect 5424 36143 5458 36177
rect 5492 36143 5526 36177
rect 5560 36143 5594 36177
rect 5628 36143 5662 36177
rect 5696 36143 5730 36177
rect 5764 36143 5798 36177
rect 5832 36143 5866 36177
rect 5900 36143 5934 36177
rect 5968 36143 6002 36177
rect 6036 36143 6070 36177
rect 6104 36143 6138 36177
rect 6172 36143 6206 36177
rect 6240 36143 6274 36177
rect 6308 36143 6342 36177
rect 6376 36143 6410 36177
rect 6444 36143 6478 36177
rect 6512 36143 6546 36177
rect 6580 36143 6614 36177
rect 6648 36143 6682 36177
rect 6716 36143 6750 36177
rect 6784 36143 6818 36177
rect 6852 36143 6886 36177
rect 6920 36143 6954 36177
rect 6988 36143 7022 36177
rect 7056 36143 7090 36177
rect 7124 36143 7158 36177
rect 7192 36143 7226 36177
rect 7260 36143 7294 36177
rect 7328 36143 7362 36177
rect 7396 36143 7430 36177
rect 7464 36143 7498 36177
rect 7532 36143 7566 36177
rect 7600 36143 7634 36177
rect 7668 36143 7702 36177
rect 7736 36143 7770 36177
rect 7804 36143 7838 36177
rect 7872 36143 7906 36177
rect 7940 36143 7974 36177
rect 8008 36143 8042 36177
rect 8076 36143 8110 36177
rect 8144 36143 8178 36177
rect 8212 36143 8246 36177
rect 8280 36143 8314 36177
rect 8348 36143 8382 36177
rect 8416 36143 8450 36177
rect 8484 36143 8518 36177
rect 8552 36143 8586 36177
rect 8620 36143 8654 36177
rect 8688 36143 8722 36177
rect 8756 36143 8790 36177
rect 8824 36143 8858 36177
rect 8892 36143 8926 36177
rect 8960 36143 8994 36177
rect 9028 36143 9062 36177
rect 9096 36143 9130 36177
rect 9164 36143 9198 36177
rect 9232 36143 9266 36177
rect 9300 36143 9334 36177
rect 9368 36143 9402 36177
rect 9436 36143 9470 36177
rect 9504 36143 9538 36177
rect 9572 36143 9606 36177
rect 9640 36143 9674 36177
rect 9708 36143 9742 36177
rect 9776 36143 9810 36177
rect 9844 36143 9878 36177
rect 9912 36143 9946 36177
rect 9980 36143 10014 36177
rect 10048 36143 10082 36177
rect 10116 36143 10150 36177
rect 10184 36143 10218 36177
rect 10252 36143 10286 36177
rect 10320 36143 10354 36177
rect 10388 36143 10422 36177
rect 10456 36143 10490 36177
rect 10524 36143 10558 36177
rect 10592 36143 10626 36177
rect 10660 36143 10694 36177
rect 10728 36143 10762 36177
rect 10796 36143 10830 36177
rect 10864 36143 10898 36177
rect 10932 36143 10966 36177
rect 11000 36143 11034 36177
rect 11068 36143 11102 36177
rect 11136 36143 11170 36177
rect 11204 36143 11238 36177
rect 11272 36143 11306 36177
rect 11340 36143 11374 36177
rect 11408 36143 11442 36177
rect 11476 36143 11510 36177
rect 11544 36143 11578 36177
rect 11612 36143 11646 36177
rect 11680 36143 11714 36177
rect 11748 36143 11782 36177
rect 11816 36143 11850 36177
rect 11884 36143 11918 36177
rect 11952 36143 11986 36177
rect 12020 36143 12054 36177
rect 12088 36143 12122 36177
rect 12156 36143 12190 36177
rect 12224 36143 12258 36177
rect 12292 36143 12326 36177
rect 12360 36143 12394 36177
rect 12428 36143 12462 36177
rect 12496 36143 12530 36177
rect 12564 36143 12598 36177
rect 12632 36143 12666 36177
rect 12700 36143 12734 36177
rect 12768 36143 12802 36177
rect 12836 36143 12870 36177
rect 12904 36143 12938 36177
rect 12972 36143 13006 36177
rect 13040 36143 13074 36177
rect 13108 36143 13142 36177
rect 13176 36143 13210 36177
rect 13244 36143 13278 36177
rect 13312 36143 13346 36177
rect 13380 36143 13414 36177
rect 13448 36143 13482 36177
rect 13516 36143 13550 36177
rect 13584 36143 13618 36177
rect 13652 36143 13686 36177
rect 13720 36143 13754 36177
rect 13788 36143 13822 36177
rect 13856 36143 13890 36177
rect 13924 36143 13958 36177
rect 13992 36143 14026 36177
rect 14060 36143 14094 36177
rect 14128 36143 14162 36177
rect 14196 36143 14361 36177
rect 603 36032 14361 36143
rect 603 35998 632 36032
rect 666 36003 14297 36032
rect 666 35998 1009 36003
rect 603 35969 1009 35998
rect 1043 35969 1081 36003
rect 1115 35969 1153 36003
rect 1187 35969 1225 36003
rect 1259 35969 1297 36003
rect 1331 35969 1369 36003
rect 1403 35969 1441 36003
rect 1475 35969 1513 36003
rect 1547 35969 1585 36003
rect 1619 35969 1657 36003
rect 1691 35969 1729 36003
rect 1763 35969 1801 36003
rect 1835 35969 1873 36003
rect 1907 35969 1945 36003
rect 1979 35969 2017 36003
rect 2051 35969 2089 36003
rect 2123 35969 2161 36003
rect 2195 35969 2233 36003
rect 2267 35969 2305 36003
rect 2339 35969 2377 36003
rect 2411 35969 2449 36003
rect 2483 35969 2521 36003
rect 2555 35969 2593 36003
rect 2627 35969 2665 36003
rect 2699 35969 2737 36003
rect 2771 35969 2809 36003
rect 2843 35969 2881 36003
rect 2915 35969 2953 36003
rect 2987 35969 3025 36003
rect 3059 35969 3097 36003
rect 3131 35969 3169 36003
rect 3203 35969 3241 36003
rect 3275 35969 3313 36003
rect 3347 35969 3385 36003
rect 3419 35969 3457 36003
rect 3491 35969 3529 36003
rect 3563 35969 3601 36003
rect 3635 35969 3673 36003
rect 3707 35969 3745 36003
rect 3779 35969 3817 36003
rect 3851 35969 3889 36003
rect 3923 35969 3961 36003
rect 3995 35969 4033 36003
rect 4067 35969 4105 36003
rect 4139 35969 4177 36003
rect 4211 35969 4249 36003
rect 4283 35969 4321 36003
rect 4355 35969 4393 36003
rect 4427 35969 4465 36003
rect 4499 35969 4537 36003
rect 4571 35969 4609 36003
rect 4643 35969 4681 36003
rect 4715 35969 4753 36003
rect 4787 35969 4825 36003
rect 4859 35969 4897 36003
rect 4931 35969 4969 36003
rect 5003 35969 5041 36003
rect 5075 35969 5113 36003
rect 5147 35969 5185 36003
rect 5219 35969 5257 36003
rect 5291 35969 5329 36003
rect 5363 35969 5401 36003
rect 5435 35969 5473 36003
rect 5507 35969 5545 36003
rect 5579 35969 5617 36003
rect 5651 35969 5689 36003
rect 5723 35969 5761 36003
rect 5795 35969 5833 36003
rect 5867 35969 5905 36003
rect 5939 35969 5977 36003
rect 6011 35969 6049 36003
rect 6083 35969 6121 36003
rect 6155 35969 6193 36003
rect 6227 35969 6265 36003
rect 6299 35969 6337 36003
rect 6371 35969 6409 36003
rect 6443 35969 6481 36003
rect 6515 35969 6553 36003
rect 6587 35969 6625 36003
rect 6659 35969 6697 36003
rect 6731 35969 6769 36003
rect 6803 35969 6841 36003
rect 6875 35969 6913 36003
rect 6947 35969 6985 36003
rect 7019 35969 7057 36003
rect 7091 35969 7129 36003
rect 7163 35969 7201 36003
rect 7235 35969 7273 36003
rect 7307 35969 7345 36003
rect 7379 35969 7417 36003
rect 7451 35969 7489 36003
rect 7523 35969 7561 36003
rect 7595 35969 7633 36003
rect 7667 35969 7705 36003
rect 7739 35969 7777 36003
rect 7811 35969 7849 36003
rect 7883 35969 7921 36003
rect 7955 35969 7993 36003
rect 8027 35969 8065 36003
rect 8099 35969 8137 36003
rect 8171 35969 8209 36003
rect 8243 35969 8281 36003
rect 8315 35969 8353 36003
rect 8387 35969 8425 36003
rect 8459 35969 8497 36003
rect 8531 35969 8569 36003
rect 8603 35969 8641 36003
rect 8675 35969 8713 36003
rect 8747 35969 8785 36003
rect 8819 35969 8857 36003
rect 8891 35969 8929 36003
rect 8963 35969 9001 36003
rect 9035 35969 9073 36003
rect 9107 35969 9145 36003
rect 9179 35969 9217 36003
rect 9251 35969 9289 36003
rect 9323 35969 9361 36003
rect 9395 35969 9433 36003
rect 9467 35969 9505 36003
rect 9539 35969 9577 36003
rect 9611 35969 9649 36003
rect 9683 35969 9721 36003
rect 9755 35969 9793 36003
rect 9827 35969 9865 36003
rect 9899 35969 9937 36003
rect 9971 35969 10009 36003
rect 10043 35969 10081 36003
rect 10115 35969 10153 36003
rect 10187 35969 10225 36003
rect 10259 35969 10297 36003
rect 10331 35969 10369 36003
rect 10403 35969 10441 36003
rect 10475 35969 10513 36003
rect 10547 35969 10585 36003
rect 10619 35969 10657 36003
rect 10691 35969 10729 36003
rect 10763 35969 10801 36003
rect 10835 35969 10873 36003
rect 10907 35969 10945 36003
rect 10979 35969 11017 36003
rect 11051 35969 11089 36003
rect 11123 35969 11161 36003
rect 11195 35969 11233 36003
rect 11267 35969 11305 36003
rect 11339 35969 11377 36003
rect 11411 35969 11449 36003
rect 11483 35969 11521 36003
rect 11555 35969 11593 36003
rect 11627 35969 11665 36003
rect 11699 35969 11737 36003
rect 11771 35969 11809 36003
rect 11843 35969 11881 36003
rect 11915 35969 11953 36003
rect 11987 35969 12025 36003
rect 12059 35969 12097 36003
rect 12131 35969 12169 36003
rect 12203 35969 12241 36003
rect 12275 35969 12313 36003
rect 12347 35969 12385 36003
rect 12419 35969 12457 36003
rect 12491 35969 12529 36003
rect 12563 35969 12601 36003
rect 12635 35969 12673 36003
rect 12707 35969 12745 36003
rect 12779 35969 12817 36003
rect 12851 35969 12889 36003
rect 12923 35969 12961 36003
rect 12995 35969 13033 36003
rect 13067 35969 13105 36003
rect 13139 35969 13177 36003
rect 13211 35969 13249 36003
rect 13283 35969 13321 36003
rect 13355 35969 13393 36003
rect 13427 35969 13465 36003
rect 13499 35969 13537 36003
rect 13571 35969 13609 36003
rect 13643 35969 13681 36003
rect 13715 35969 13753 36003
rect 13787 35969 13825 36003
rect 13859 35969 13897 36003
rect 13931 35969 13969 36003
rect 14003 35998 14297 36003
rect 14331 35998 14361 36032
rect 14003 35969 14361 35998
rect 603 35964 14361 35969
rect 603 35930 632 35964
rect 666 35930 14297 35964
rect 14331 35930 14361 35964
rect 603 35896 14361 35930
rect 603 35862 632 35896
rect 666 35884 14297 35896
rect 666 35862 807 35884
rect 603 35850 807 35862
rect 841 35862 14297 35884
rect 14331 35862 14361 35896
rect 841 35850 14361 35862
rect 603 35828 14361 35850
rect 603 35794 632 35828
rect 666 35812 14297 35828
rect 666 35794 807 35812
rect 603 35778 807 35794
rect 841 35805 14297 35812
rect 841 35778 14122 35805
rect 603 35771 14122 35778
rect 14156 35794 14297 35805
rect 14331 35794 14361 35828
rect 14156 35771 14361 35794
rect 603 35760 14361 35771
rect 603 35726 632 35760
rect 666 35740 14297 35760
rect 666 35726 807 35740
rect 603 35706 807 35726
rect 841 35733 14297 35740
rect 841 35706 14122 35733
rect 603 35699 14122 35706
rect 14156 35726 14297 35733
rect 14331 35726 14361 35760
rect 14156 35699 14361 35726
rect 603 35692 14361 35699
rect 603 35658 632 35692
rect 666 35668 14297 35692
rect 666 35658 807 35668
rect 603 35634 807 35658
rect 841 35661 14297 35668
rect 841 35634 14122 35661
rect 603 35627 14122 35634
rect 14156 35658 14297 35661
rect 14331 35658 14361 35692
rect 14156 35627 14361 35658
rect 603 35624 14361 35627
rect 603 35590 632 35624
rect 666 35596 14297 35624
rect 666 35590 807 35596
rect 603 35562 807 35590
rect 841 35590 14297 35596
rect 14331 35590 14361 35624
rect 841 35589 14361 35590
rect 841 35562 14122 35589
rect 603 35556 14122 35562
rect 603 35522 632 35556
rect 666 35555 14122 35556
rect 14156 35556 14361 35589
rect 14156 35555 14297 35556
rect 666 35524 14297 35555
rect 666 35522 807 35524
rect 603 35490 807 35522
rect 841 35522 14297 35524
rect 14331 35522 14361 35556
rect 841 35517 14361 35522
rect 841 35490 14122 35517
rect 603 35488 14122 35490
rect 603 35454 632 35488
rect 666 35483 14122 35488
rect 14156 35488 14361 35517
rect 14156 35483 14297 35488
rect 666 35454 14297 35483
rect 14331 35454 14361 35488
rect 603 35452 14361 35454
rect 603 35420 807 35452
rect 603 35386 632 35420
rect 666 35418 807 35420
rect 841 35445 14361 35452
rect 841 35418 14122 35445
rect 666 35411 14122 35418
rect 14156 35420 14361 35445
rect 14156 35411 14297 35420
rect 666 35386 14297 35411
rect 14331 35386 14361 35420
rect 603 35380 14361 35386
rect 603 35352 807 35380
rect 603 35318 632 35352
rect 666 35346 807 35352
rect 841 35373 14361 35380
rect 841 35346 14122 35373
rect 666 35339 14122 35346
rect 14156 35352 14361 35373
rect 14156 35339 14297 35352
rect 666 35318 14297 35339
rect 14331 35318 14361 35352
rect 603 35308 14361 35318
rect 603 35284 807 35308
rect 603 35250 632 35284
rect 666 35274 807 35284
rect 841 35301 14361 35308
rect 841 35274 14122 35301
rect 666 35267 14122 35274
rect 14156 35284 14361 35301
rect 14156 35267 14297 35284
rect 666 35250 14297 35267
rect 14331 35250 14361 35284
rect 603 35236 14361 35250
rect 603 35216 807 35236
rect 603 35182 632 35216
rect 666 35202 807 35216
rect 841 35229 14361 35236
rect 841 35202 14122 35229
rect 666 35195 14122 35202
rect 14156 35216 14361 35229
rect 14156 35195 14297 35216
rect 666 35182 14297 35195
rect 14331 35182 14361 35216
rect 603 35164 14361 35182
rect 603 35148 807 35164
rect 603 35114 632 35148
rect 666 35130 807 35148
rect 841 35157 14361 35164
rect 841 35130 14122 35157
rect 666 35123 14122 35130
rect 14156 35148 14361 35157
rect 14156 35123 14297 35148
rect 666 35114 14297 35123
rect 14331 35114 14361 35148
rect 603 35092 14361 35114
rect 603 35080 807 35092
rect 603 35046 632 35080
rect 666 35058 807 35080
rect 841 35085 14361 35092
rect 841 35058 14122 35085
rect 666 35051 14122 35058
rect 14156 35080 14361 35085
rect 14156 35051 14297 35080
rect 666 35046 14297 35051
rect 14331 35046 14361 35080
rect 603 35020 14361 35046
rect 603 35012 807 35020
rect 603 34978 632 35012
rect 666 34986 807 35012
rect 841 35013 14361 35020
rect 841 34986 14122 35013
rect 666 34979 14122 34986
rect 14156 35012 14361 35013
rect 14156 34979 14297 35012
rect 666 34978 14297 34979
rect 14331 34978 14361 35012
rect 603 34948 14361 34978
rect 603 34944 807 34948
rect 603 34910 632 34944
rect 666 34914 807 34944
rect 841 34944 14361 34948
rect 841 34941 14297 34944
rect 841 34914 14122 34941
rect 666 34910 14122 34914
rect 603 34907 14122 34910
rect 14156 34910 14297 34941
rect 14331 34910 14361 34944
rect 14156 34907 14361 34910
rect 603 34876 14361 34907
rect 603 34842 632 34876
rect 666 34842 807 34876
rect 841 34869 14297 34876
rect 841 34842 14122 34869
rect 603 34835 14122 34842
rect 14156 34842 14297 34869
rect 14331 34842 14361 34876
rect 14156 34835 14361 34842
rect 603 34831 14361 34835
rect 603 34808 1026 34831
rect 603 34774 632 34808
rect 666 34804 1026 34808
rect 666 34774 807 34804
rect 603 34770 807 34774
rect 841 34770 1026 34804
rect 603 34740 1026 34770
rect 603 34706 632 34740
rect 666 34732 1026 34740
rect 666 34706 807 34732
rect 603 34698 807 34706
rect 841 34698 1026 34732
rect 13968 34808 14361 34831
rect 13968 34797 14297 34808
rect 13968 34763 14122 34797
rect 14156 34774 14297 34797
rect 14331 34774 14361 34808
rect 14156 34763 14361 34774
rect 13968 34740 14361 34763
rect 13968 34725 14297 34740
rect 603 34672 1026 34698
rect 603 34638 632 34672
rect 666 34660 1026 34672
rect 666 34638 807 34660
rect 603 34626 807 34638
rect 841 34626 1026 34660
rect 603 34604 1026 34626
rect 603 34570 632 34604
rect 666 34588 1026 34604
rect 666 34570 807 34588
rect 603 34554 807 34570
rect 841 34554 1026 34588
rect 603 34536 1026 34554
rect 603 34502 632 34536
rect 666 34516 1026 34536
rect 666 34502 807 34516
rect 603 34482 807 34502
rect 841 34482 1026 34516
rect 603 34468 1026 34482
rect 603 34434 632 34468
rect 666 34444 1026 34468
rect 666 34434 807 34444
rect 603 34410 807 34434
rect 841 34410 1026 34444
rect 603 34400 1026 34410
rect 603 34366 632 34400
rect 666 34372 1026 34400
rect 666 34366 807 34372
rect 603 34338 807 34366
rect 841 34338 1026 34372
rect 603 34332 1026 34338
rect 603 34298 632 34332
rect 666 34300 1026 34332
rect 666 34298 807 34300
rect 603 34266 807 34298
rect 841 34266 1026 34300
rect 603 34264 1026 34266
rect 603 34230 632 34264
rect 666 34230 1026 34264
rect 603 34228 1026 34230
rect 603 34196 807 34228
rect 603 34162 632 34196
rect 666 34194 807 34196
rect 841 34194 1026 34228
rect 666 34162 1026 34194
rect 603 34156 1026 34162
rect 603 34128 807 34156
rect 603 34094 632 34128
rect 666 34122 807 34128
rect 841 34122 1026 34156
rect 666 34094 1026 34122
rect 603 34084 1026 34094
rect 603 34060 807 34084
rect 603 34026 632 34060
rect 666 34050 807 34060
rect 841 34050 1026 34084
rect 666 34026 1026 34050
rect 603 34012 1026 34026
rect 603 33992 807 34012
rect 603 33958 632 33992
rect 666 33978 807 33992
rect 841 33978 1026 34012
rect 666 33958 1026 33978
rect 603 33940 1026 33958
rect 603 33924 807 33940
rect 603 33890 632 33924
rect 666 33906 807 33924
rect 841 33906 1026 33940
rect 666 33890 1026 33906
rect 603 33868 1026 33890
rect 603 33856 807 33868
rect 603 33822 632 33856
rect 666 33834 807 33856
rect 841 33834 1026 33868
rect 666 33822 1026 33834
rect 603 33796 1026 33822
rect 603 33788 807 33796
rect 603 33754 632 33788
rect 666 33762 807 33788
rect 841 33762 1026 33796
rect 666 33754 1026 33762
rect 603 33724 1026 33754
rect 603 33720 807 33724
rect 603 33686 632 33720
rect 666 33690 807 33720
rect 841 33690 1026 33724
rect 666 33686 1026 33690
rect 603 33652 1026 33686
rect 603 33618 632 33652
rect 666 33618 807 33652
rect 841 33618 1026 33652
rect 603 33584 1026 33618
rect 603 33550 632 33584
rect 666 33580 1026 33584
rect 666 33550 807 33580
rect 603 33546 807 33550
rect 841 33546 1026 33580
rect 603 33516 1026 33546
rect 603 33482 632 33516
rect 666 33508 1026 33516
rect 666 33482 807 33508
rect 603 33474 807 33482
rect 841 33474 1026 33508
rect 603 33448 1026 33474
rect 603 33414 632 33448
rect 666 33436 1026 33448
rect 666 33414 807 33436
rect 603 33402 807 33414
rect 841 33402 1026 33436
rect 603 33380 1026 33402
rect 603 33346 632 33380
rect 666 33364 1026 33380
rect 666 33346 807 33364
rect 603 33330 807 33346
rect 841 33330 1026 33364
rect 603 33312 1026 33330
rect 603 33278 632 33312
rect 666 33292 1026 33312
rect 666 33278 807 33292
rect 603 33258 807 33278
rect 841 33258 1026 33292
rect 603 33244 1026 33258
rect 603 33210 632 33244
rect 666 33220 1026 33244
rect 666 33210 807 33220
rect 603 33186 807 33210
rect 841 33186 1026 33220
rect 603 33176 1026 33186
rect 603 33142 632 33176
rect 666 33148 1026 33176
rect 666 33142 807 33148
rect 603 33114 807 33142
rect 841 33114 1026 33148
rect 603 33108 1026 33114
rect 603 33074 632 33108
rect 666 33076 1026 33108
rect 666 33074 807 33076
rect 603 33042 807 33074
rect 841 33042 1026 33076
rect 603 33040 1026 33042
rect 603 33006 632 33040
rect 666 33006 1026 33040
rect 603 33004 1026 33006
rect 603 32972 807 33004
rect 603 32938 632 32972
rect 666 32970 807 32972
rect 841 32970 1026 33004
rect 666 32938 1026 32970
rect 603 32932 1026 32938
rect 603 32904 807 32932
rect 603 32870 632 32904
rect 666 32898 807 32904
rect 841 32898 1026 32932
rect 666 32870 1026 32898
rect 603 32860 1026 32870
rect 603 32836 807 32860
rect 603 32802 632 32836
rect 666 32826 807 32836
rect 841 32826 1026 32860
rect 666 32802 1026 32826
rect 603 32788 1026 32802
rect 603 32768 807 32788
rect 603 32734 632 32768
rect 666 32754 807 32768
rect 841 32754 1026 32788
rect 666 32734 1026 32754
rect 603 32716 1026 32734
rect 603 32700 807 32716
rect 603 32666 632 32700
rect 666 32682 807 32700
rect 841 32682 1026 32716
rect 666 32666 1026 32682
rect 603 32644 1026 32666
rect 603 32632 807 32644
rect 603 32598 632 32632
rect 666 32610 807 32632
rect 841 32610 1026 32644
rect 666 32598 1026 32610
rect 603 32572 1026 32598
rect 603 32564 807 32572
rect 603 32530 632 32564
rect 666 32538 807 32564
rect 841 32538 1026 32572
rect 666 32530 1026 32538
rect 603 32500 1026 32530
rect 603 32496 807 32500
rect 603 32462 632 32496
rect 666 32466 807 32496
rect 841 32466 1026 32500
rect 666 32462 1026 32466
rect 603 32428 1026 32462
rect 603 32394 632 32428
rect 666 32394 807 32428
rect 841 32394 1026 32428
rect 603 32360 1026 32394
rect 603 32326 632 32360
rect 666 32356 1026 32360
rect 666 32326 807 32356
rect 603 32322 807 32326
rect 841 32322 1026 32356
rect 603 32292 1026 32322
rect 603 32258 632 32292
rect 666 32284 1026 32292
rect 666 32258 807 32284
rect 603 32250 807 32258
rect 841 32250 1026 32284
rect 603 32224 1026 32250
rect 603 32190 632 32224
rect 666 32212 1026 32224
rect 666 32190 807 32212
rect 603 32178 807 32190
rect 841 32178 1026 32212
rect 603 32156 1026 32178
rect 603 32122 632 32156
rect 666 32140 1026 32156
rect 666 32122 807 32140
rect 603 32106 807 32122
rect 841 32106 1026 32140
rect 603 32088 1026 32106
rect 603 32054 632 32088
rect 666 32068 1026 32088
rect 666 32054 807 32068
rect 603 32034 807 32054
rect 841 32034 1026 32068
rect 603 32020 1026 32034
rect 603 31986 632 32020
rect 666 31996 1026 32020
rect 666 31986 807 31996
rect 603 31962 807 31986
rect 841 31962 1026 31996
rect 603 31952 1026 31962
rect 603 31918 632 31952
rect 666 31924 1026 31952
rect 666 31918 807 31924
rect 603 31890 807 31918
rect 841 31890 1026 31924
rect 603 31884 1026 31890
rect 603 31850 632 31884
rect 666 31852 1026 31884
rect 666 31850 807 31852
rect 603 31818 807 31850
rect 841 31818 1026 31852
rect 603 31816 1026 31818
rect 603 31782 632 31816
rect 666 31782 1026 31816
rect 603 31780 1026 31782
rect 603 31748 807 31780
rect 603 31714 632 31748
rect 666 31746 807 31748
rect 841 31746 1026 31780
rect 666 31714 1026 31746
rect 603 31708 1026 31714
rect 603 31680 807 31708
rect 603 31646 632 31680
rect 666 31674 807 31680
rect 841 31674 1026 31708
rect 666 31646 1026 31674
rect 603 31636 1026 31646
rect 603 31612 807 31636
rect 603 31578 632 31612
rect 666 31602 807 31612
rect 841 31602 1026 31636
rect 666 31578 1026 31602
rect 603 31564 1026 31578
rect 603 31544 807 31564
rect 603 31510 632 31544
rect 666 31530 807 31544
rect 841 31530 1026 31564
rect 666 31510 1026 31530
rect 603 31492 1026 31510
rect 603 31476 807 31492
rect 603 31442 632 31476
rect 666 31458 807 31476
rect 841 31458 1026 31492
rect 666 31442 1026 31458
rect 603 31420 1026 31442
rect 603 31408 807 31420
rect 603 31374 632 31408
rect 666 31386 807 31408
rect 841 31386 1026 31420
rect 666 31374 1026 31386
rect 603 31348 1026 31374
rect 603 31340 807 31348
rect 603 31306 632 31340
rect 666 31314 807 31340
rect 841 31314 1026 31348
rect 666 31306 1026 31314
rect 603 31276 1026 31306
rect 603 31272 807 31276
rect 603 31238 632 31272
rect 666 31242 807 31272
rect 841 31242 1026 31276
rect 666 31238 1026 31242
rect 603 31204 1026 31238
rect 603 31170 632 31204
rect 666 31170 807 31204
rect 841 31170 1026 31204
rect 603 31136 1026 31170
rect 603 31102 632 31136
rect 666 31132 1026 31136
rect 666 31102 807 31132
rect 603 31098 807 31102
rect 841 31098 1026 31132
rect 603 31068 1026 31098
rect 603 31034 632 31068
rect 666 31060 1026 31068
rect 666 31034 807 31060
rect 603 31026 807 31034
rect 841 31026 1026 31060
rect 603 31000 1026 31026
rect 603 30966 632 31000
rect 666 30988 1026 31000
rect 666 30966 807 30988
rect 603 30954 807 30966
rect 841 30954 1026 30988
rect 603 30932 1026 30954
rect 603 30898 632 30932
rect 666 30916 1026 30932
rect 666 30898 807 30916
rect 603 30882 807 30898
rect 841 30882 1026 30916
rect 603 30864 1026 30882
rect 603 30830 632 30864
rect 666 30844 1026 30864
rect 666 30830 807 30844
rect 603 30810 807 30830
rect 841 30810 1026 30844
rect 603 30796 1026 30810
rect 603 30762 632 30796
rect 666 30772 1026 30796
rect 666 30762 807 30772
rect 603 30738 807 30762
rect 841 30738 1026 30772
rect 603 30728 1026 30738
rect 603 30694 632 30728
rect 666 30700 1026 30728
rect 666 30694 807 30700
rect 603 30666 807 30694
rect 841 30666 1026 30700
rect 603 30660 1026 30666
rect 603 30626 632 30660
rect 666 30628 1026 30660
rect 666 30626 807 30628
rect 603 30594 807 30626
rect 841 30594 1026 30628
rect 603 30592 1026 30594
rect 603 30558 632 30592
rect 666 30558 1026 30592
rect 603 30556 1026 30558
rect 603 30524 807 30556
rect 603 30490 632 30524
rect 666 30522 807 30524
rect 841 30522 1026 30556
rect 666 30490 1026 30522
rect 603 30484 1026 30490
rect 603 30456 807 30484
rect 603 30422 632 30456
rect 666 30450 807 30456
rect 841 30450 1026 30484
rect 666 30422 1026 30450
rect 603 30412 1026 30422
rect 603 30388 807 30412
rect 603 30354 632 30388
rect 666 30378 807 30388
rect 841 30378 1026 30412
rect 666 30354 1026 30378
rect 603 30340 1026 30354
rect 603 30320 807 30340
rect 603 30286 632 30320
rect 666 30306 807 30320
rect 841 30306 1026 30340
rect 666 30286 1026 30306
rect 603 30268 1026 30286
rect 603 30252 807 30268
rect 603 30218 632 30252
rect 666 30234 807 30252
rect 841 30234 1026 30268
rect 666 30218 1026 30234
rect 603 30196 1026 30218
rect 603 30184 807 30196
rect 603 30150 632 30184
rect 666 30162 807 30184
rect 841 30162 1026 30196
rect 666 30150 1026 30162
rect 603 30124 1026 30150
rect 603 30116 807 30124
rect 603 30082 632 30116
rect 666 30090 807 30116
rect 841 30090 1026 30124
rect 666 30082 1026 30090
rect 603 30052 1026 30082
rect 603 30048 807 30052
rect 603 30014 632 30048
rect 666 30018 807 30048
rect 841 30018 1026 30052
rect 666 30014 1026 30018
rect 603 29980 1026 30014
rect 603 29946 632 29980
rect 666 29946 807 29980
rect 841 29946 1026 29980
rect 603 29912 1026 29946
rect 603 29878 632 29912
rect 666 29908 1026 29912
rect 666 29878 807 29908
rect 603 29874 807 29878
rect 841 29874 1026 29908
rect 603 29844 1026 29874
rect 603 29810 632 29844
rect 666 29836 1026 29844
rect 666 29810 807 29836
rect 603 29802 807 29810
rect 841 29802 1026 29836
rect 603 29776 1026 29802
rect 603 29742 632 29776
rect 666 29764 1026 29776
rect 666 29742 807 29764
rect 603 29730 807 29742
rect 841 29730 1026 29764
rect 603 29708 1026 29730
rect 603 29674 632 29708
rect 666 29692 1026 29708
rect 666 29674 807 29692
rect 603 29658 807 29674
rect 841 29658 1026 29692
rect 603 29640 1026 29658
rect 603 29606 632 29640
rect 666 29620 1026 29640
rect 666 29606 807 29620
rect 603 29586 807 29606
rect 841 29586 1026 29620
rect 603 29572 1026 29586
rect 603 29538 632 29572
rect 666 29548 1026 29572
rect 666 29538 807 29548
rect 603 29514 807 29538
rect 841 29514 1026 29548
rect 603 29504 1026 29514
rect 603 29470 632 29504
rect 666 29476 1026 29504
rect 666 29470 807 29476
rect 603 29442 807 29470
rect 841 29442 1026 29476
rect 603 29436 1026 29442
rect 603 29402 632 29436
rect 666 29404 1026 29436
rect 666 29402 807 29404
rect 603 29370 807 29402
rect 841 29370 1026 29404
rect 603 29368 1026 29370
rect 603 29334 632 29368
rect 666 29334 1026 29368
rect 603 29332 1026 29334
rect 603 29300 807 29332
rect 603 29266 632 29300
rect 666 29298 807 29300
rect 841 29298 1026 29332
rect 666 29266 1026 29298
rect 603 29260 1026 29266
rect 603 29232 807 29260
rect 603 29198 632 29232
rect 666 29226 807 29232
rect 841 29226 1026 29260
rect 666 29198 1026 29226
rect 603 29188 1026 29198
rect 603 29164 807 29188
rect 603 29130 632 29164
rect 666 29154 807 29164
rect 841 29154 1026 29188
rect 666 29130 1026 29154
rect 603 29116 1026 29130
rect 603 29096 807 29116
rect 603 29062 632 29096
rect 666 29082 807 29096
rect 841 29082 1026 29116
rect 666 29062 1026 29082
rect 603 29044 1026 29062
rect 603 29028 807 29044
rect 603 28994 632 29028
rect 666 29010 807 29028
rect 841 29010 1026 29044
rect 666 28994 1026 29010
rect 603 28972 1026 28994
rect 603 28960 807 28972
rect 603 28926 632 28960
rect 666 28938 807 28960
rect 841 28938 1026 28972
rect 666 28926 1026 28938
rect 603 28900 1026 28926
rect 603 28892 807 28900
rect 603 28858 632 28892
rect 666 28866 807 28892
rect 841 28866 1026 28900
rect 666 28858 1026 28866
rect 603 28828 1026 28858
rect 603 28824 807 28828
rect 603 28790 632 28824
rect 666 28794 807 28824
rect 841 28794 1026 28828
rect 666 28790 1026 28794
rect 603 28756 1026 28790
rect 603 28722 632 28756
rect 666 28722 807 28756
rect 841 28722 1026 28756
rect 603 28688 1026 28722
rect 603 28654 632 28688
rect 666 28684 1026 28688
rect 666 28654 807 28684
rect 603 28650 807 28654
rect 841 28650 1026 28684
rect 603 28620 1026 28650
rect 603 28586 632 28620
rect 666 28612 1026 28620
rect 666 28586 807 28612
rect 603 28578 807 28586
rect 841 28578 1026 28612
rect 603 28552 1026 28578
rect 603 28518 632 28552
rect 666 28540 1026 28552
rect 666 28518 807 28540
rect 603 28506 807 28518
rect 841 28506 1026 28540
rect 603 28484 1026 28506
rect 603 28450 632 28484
rect 666 28468 1026 28484
rect 666 28450 807 28468
rect 603 28434 807 28450
rect 841 28434 1026 28468
rect 603 28416 1026 28434
rect 603 28382 632 28416
rect 666 28396 1026 28416
rect 666 28382 807 28396
rect 603 28362 807 28382
rect 841 28362 1026 28396
rect 603 28348 1026 28362
rect 603 28314 632 28348
rect 666 28324 1026 28348
rect 666 28314 807 28324
rect 603 28290 807 28314
rect 841 28290 1026 28324
rect 603 28280 1026 28290
rect 603 28246 632 28280
rect 666 28252 1026 28280
rect 666 28246 807 28252
rect 603 28218 807 28246
rect 841 28218 1026 28252
rect 603 28212 1026 28218
rect 603 28178 632 28212
rect 666 28180 1026 28212
rect 666 28178 807 28180
rect 603 28146 807 28178
rect 841 28146 1026 28180
rect 603 28144 1026 28146
rect 603 28110 632 28144
rect 666 28110 1026 28144
rect 603 28108 1026 28110
rect 603 28076 807 28108
rect 603 28042 632 28076
rect 666 28074 807 28076
rect 841 28074 1026 28108
rect 666 28042 1026 28074
rect 603 28036 1026 28042
rect 603 28008 807 28036
rect 603 27974 632 28008
rect 666 28002 807 28008
rect 841 28002 1026 28036
rect 666 27974 1026 28002
rect 603 27964 1026 27974
rect 603 27940 807 27964
rect 603 27906 632 27940
rect 666 27930 807 27940
rect 841 27930 1026 27964
rect 666 27906 1026 27930
rect 603 27892 1026 27906
rect 603 27872 807 27892
rect 603 27838 632 27872
rect 666 27858 807 27872
rect 841 27858 1026 27892
rect 666 27838 1026 27858
rect 603 27820 1026 27838
rect 603 27804 807 27820
rect 603 27770 632 27804
rect 666 27786 807 27804
rect 841 27786 1026 27820
rect 666 27770 1026 27786
rect 603 27748 1026 27770
rect 603 27736 807 27748
rect 603 27702 632 27736
rect 666 27714 807 27736
rect 841 27714 1026 27748
rect 666 27702 1026 27714
rect 603 27676 1026 27702
rect 603 27668 807 27676
rect 603 27634 632 27668
rect 666 27642 807 27668
rect 841 27642 1026 27676
rect 666 27634 1026 27642
rect 603 27604 1026 27634
rect 603 27600 807 27604
rect 603 27566 632 27600
rect 666 27570 807 27600
rect 841 27570 1026 27604
rect 666 27566 1026 27570
rect 603 27532 1026 27566
rect 603 27498 632 27532
rect 666 27498 807 27532
rect 841 27498 1026 27532
rect 603 27464 1026 27498
rect 603 27430 632 27464
rect 666 27460 1026 27464
rect 666 27430 807 27460
rect 603 27426 807 27430
rect 841 27426 1026 27460
rect 603 27396 1026 27426
rect 603 27362 632 27396
rect 666 27388 1026 27396
rect 666 27362 807 27388
rect 603 27354 807 27362
rect 841 27354 1026 27388
rect 603 27328 1026 27354
rect 603 27294 632 27328
rect 666 27316 1026 27328
rect 666 27294 807 27316
rect 603 27282 807 27294
rect 841 27282 1026 27316
rect 603 27260 1026 27282
rect 603 27226 632 27260
rect 666 27244 1026 27260
rect 666 27226 807 27244
rect 603 27210 807 27226
rect 841 27210 1026 27244
rect 603 27192 1026 27210
rect 603 27158 632 27192
rect 666 27172 1026 27192
rect 666 27158 807 27172
rect 603 27138 807 27158
rect 841 27138 1026 27172
rect 603 27124 1026 27138
rect 603 27090 632 27124
rect 666 27100 1026 27124
rect 666 27090 807 27100
rect 603 27066 807 27090
rect 841 27066 1026 27100
rect 603 27056 1026 27066
rect 603 27022 632 27056
rect 666 27028 1026 27056
rect 666 27022 807 27028
rect 603 26994 807 27022
rect 841 26994 1026 27028
rect 603 26988 1026 26994
rect 603 26954 632 26988
rect 666 26956 1026 26988
rect 666 26954 807 26956
rect 603 26922 807 26954
rect 841 26922 1026 26956
rect 603 26920 1026 26922
rect 603 26886 632 26920
rect 666 26886 1026 26920
rect 603 26884 1026 26886
rect 603 26852 807 26884
rect 603 26818 632 26852
rect 666 26850 807 26852
rect 841 26850 1026 26884
rect 666 26818 1026 26850
rect 603 26812 1026 26818
rect 603 26784 807 26812
rect 603 26750 632 26784
rect 666 26778 807 26784
rect 841 26778 1026 26812
rect 666 26750 1026 26778
rect 603 26740 1026 26750
rect 603 26716 807 26740
rect 603 26682 632 26716
rect 666 26706 807 26716
rect 841 26706 1026 26740
rect 666 26682 1026 26706
rect 603 26668 1026 26682
rect 603 26648 807 26668
rect 603 26614 632 26648
rect 666 26634 807 26648
rect 841 26634 1026 26668
rect 666 26614 1026 26634
rect 603 26596 1026 26614
rect 603 26580 807 26596
rect 603 26546 632 26580
rect 666 26562 807 26580
rect 841 26562 1026 26596
rect 666 26546 1026 26562
rect 603 26524 1026 26546
rect 603 26512 807 26524
rect 603 26478 632 26512
rect 666 26490 807 26512
rect 841 26490 1026 26524
rect 666 26478 1026 26490
rect 603 26452 1026 26478
rect 603 26444 807 26452
rect 603 26410 632 26444
rect 666 26418 807 26444
rect 841 26418 1026 26452
rect 666 26410 1026 26418
rect 603 26380 1026 26410
rect 603 26376 807 26380
rect 603 26342 632 26376
rect 666 26346 807 26376
rect 841 26346 1026 26380
rect 666 26342 1026 26346
rect 603 26308 1026 26342
rect 603 26274 632 26308
rect 666 26274 807 26308
rect 841 26274 1026 26308
rect 603 26240 1026 26274
rect 603 26206 632 26240
rect 666 26236 1026 26240
rect 666 26206 807 26236
rect 603 26202 807 26206
rect 841 26202 1026 26236
rect 603 26172 1026 26202
rect 603 26138 632 26172
rect 666 26164 1026 26172
rect 666 26138 807 26164
rect 603 26130 807 26138
rect 841 26130 1026 26164
rect 603 26104 1026 26130
rect 603 26070 632 26104
rect 666 26092 1026 26104
rect 666 26070 807 26092
rect 603 26058 807 26070
rect 841 26058 1026 26092
rect 603 26036 1026 26058
rect 603 26002 632 26036
rect 666 26020 1026 26036
rect 666 26002 807 26020
rect 603 25986 807 26002
rect 841 25986 1026 26020
rect 603 25968 1026 25986
rect 603 25934 632 25968
rect 666 25948 1026 25968
rect 666 25934 807 25948
rect 603 25914 807 25934
rect 841 25914 1026 25948
rect 603 25900 1026 25914
rect 603 25866 632 25900
rect 666 25876 1026 25900
rect 666 25866 807 25876
rect 603 25842 807 25866
rect 841 25842 1026 25876
rect 603 25832 1026 25842
rect 603 25798 632 25832
rect 666 25804 1026 25832
rect 666 25798 807 25804
rect 603 25770 807 25798
rect 841 25770 1026 25804
rect 603 25764 1026 25770
rect 603 25730 632 25764
rect 666 25732 1026 25764
rect 666 25730 807 25732
rect 603 25698 807 25730
rect 841 25698 1026 25732
rect 603 25696 1026 25698
rect 603 25662 632 25696
rect 666 25662 1026 25696
rect 603 25660 1026 25662
rect 603 25628 807 25660
rect 603 25594 632 25628
rect 666 25626 807 25628
rect 841 25626 1026 25660
rect 666 25594 1026 25626
rect 603 25588 1026 25594
rect 603 25560 807 25588
rect 603 25526 632 25560
rect 666 25554 807 25560
rect 841 25554 1026 25588
rect 666 25526 1026 25554
rect 603 25516 1026 25526
rect 603 25492 807 25516
rect 603 25458 632 25492
rect 666 25482 807 25492
rect 841 25482 1026 25516
rect 666 25458 1026 25482
rect 603 25444 1026 25458
rect 603 25424 807 25444
rect 603 25390 632 25424
rect 666 25410 807 25424
rect 841 25410 1026 25444
rect 666 25390 1026 25410
rect 603 25372 1026 25390
rect 603 25356 807 25372
rect 603 25322 632 25356
rect 666 25338 807 25356
rect 841 25338 1026 25372
rect 666 25322 1026 25338
rect 603 25300 1026 25322
rect 603 25288 807 25300
rect 603 25254 632 25288
rect 666 25266 807 25288
rect 841 25266 1026 25300
rect 666 25254 1026 25266
rect 603 25228 1026 25254
rect 603 25220 807 25228
rect 603 25186 632 25220
rect 666 25194 807 25220
rect 841 25194 1026 25228
rect 666 25186 1026 25194
rect 603 25156 1026 25186
rect 603 25152 807 25156
rect 603 25118 632 25152
rect 666 25122 807 25152
rect 841 25122 1026 25156
rect 666 25118 1026 25122
rect 603 25084 1026 25118
rect 603 25050 632 25084
rect 666 25050 807 25084
rect 841 25050 1026 25084
rect 603 25016 1026 25050
rect 603 24982 632 25016
rect 666 25012 1026 25016
rect 666 24982 807 25012
rect 603 24978 807 24982
rect 841 24978 1026 25012
rect 603 24948 1026 24978
rect 603 24914 632 24948
rect 666 24940 1026 24948
rect 666 24914 807 24940
rect 603 24906 807 24914
rect 841 24906 1026 24940
rect 603 24880 1026 24906
rect 603 24846 632 24880
rect 666 24868 1026 24880
rect 666 24846 807 24868
rect 603 24834 807 24846
rect 841 24834 1026 24868
rect 603 24812 1026 24834
rect 603 24778 632 24812
rect 666 24796 1026 24812
rect 666 24778 807 24796
rect 603 24762 807 24778
rect 841 24762 1026 24796
rect 603 24744 1026 24762
rect 603 24710 632 24744
rect 666 24724 1026 24744
rect 666 24710 807 24724
rect 603 24690 807 24710
rect 841 24690 1026 24724
rect 603 24676 1026 24690
rect 603 24642 632 24676
rect 666 24652 1026 24676
rect 666 24642 807 24652
rect 603 24618 807 24642
rect 841 24618 1026 24652
rect 603 24608 1026 24618
rect 603 24574 632 24608
rect 666 24580 1026 24608
rect 666 24574 807 24580
rect 603 24546 807 24574
rect 841 24546 1026 24580
rect 603 24540 1026 24546
rect 603 24506 632 24540
rect 666 24508 1026 24540
rect 666 24506 807 24508
rect 603 24474 807 24506
rect 841 24474 1026 24508
rect 603 24472 1026 24474
rect 603 24438 632 24472
rect 666 24438 1026 24472
rect 603 24436 1026 24438
rect 603 24404 807 24436
rect 603 24370 632 24404
rect 666 24402 807 24404
rect 841 24402 1026 24436
rect 666 24370 1026 24402
rect 603 24364 1026 24370
rect 603 24336 807 24364
rect 603 24302 632 24336
rect 666 24330 807 24336
rect 841 24330 1026 24364
rect 666 24302 1026 24330
rect 603 24292 1026 24302
rect 603 24268 807 24292
rect 603 24234 632 24268
rect 666 24258 807 24268
rect 841 24258 1026 24292
rect 666 24234 1026 24258
rect 603 24220 1026 24234
rect 603 24200 807 24220
rect 603 24166 632 24200
rect 666 24186 807 24200
rect 841 24186 1026 24220
rect 666 24166 1026 24186
rect 603 24148 1026 24166
rect 603 24132 807 24148
rect 603 24098 632 24132
rect 666 24114 807 24132
rect 841 24114 1026 24148
rect 666 24098 1026 24114
rect 603 24076 1026 24098
rect 603 24064 807 24076
rect 603 24030 632 24064
rect 666 24042 807 24064
rect 841 24042 1026 24076
rect 666 24030 1026 24042
rect 603 24004 1026 24030
rect 603 23996 807 24004
rect 603 23962 632 23996
rect 666 23970 807 23996
rect 841 23970 1026 24004
rect 666 23962 1026 23970
rect 603 23932 1026 23962
rect 603 23928 807 23932
rect 603 23894 632 23928
rect 666 23898 807 23928
rect 841 23898 1026 23932
rect 666 23894 1026 23898
rect 603 23860 1026 23894
rect 603 23826 632 23860
rect 666 23826 807 23860
rect 841 23826 1026 23860
rect 603 23792 1026 23826
rect 603 23758 632 23792
rect 666 23788 1026 23792
rect 666 23758 807 23788
rect 603 23754 807 23758
rect 841 23754 1026 23788
rect 603 23724 1026 23754
rect 603 23690 632 23724
rect 666 23716 1026 23724
rect 666 23690 807 23716
rect 603 23682 807 23690
rect 841 23682 1026 23716
rect 603 23656 1026 23682
rect 603 23622 632 23656
rect 666 23644 1026 23656
rect 666 23622 807 23644
rect 603 23610 807 23622
rect 841 23610 1026 23644
rect 603 23588 1026 23610
rect 603 23554 632 23588
rect 666 23572 1026 23588
rect 666 23554 807 23572
rect 603 23538 807 23554
rect 841 23538 1026 23572
rect 603 23520 1026 23538
rect 603 23486 632 23520
rect 666 23500 1026 23520
rect 666 23486 807 23500
rect 603 23466 807 23486
rect 841 23466 1026 23500
rect 603 23452 1026 23466
rect 603 23418 632 23452
rect 666 23428 1026 23452
rect 666 23418 807 23428
rect 603 23394 807 23418
rect 841 23394 1026 23428
rect 603 23384 1026 23394
rect 603 23350 632 23384
rect 666 23356 1026 23384
rect 666 23350 807 23356
rect 603 23322 807 23350
rect 841 23322 1026 23356
rect 603 23316 1026 23322
rect 603 23282 632 23316
rect 666 23284 1026 23316
rect 666 23282 807 23284
rect 603 23250 807 23282
rect 841 23250 1026 23284
rect 603 23248 1026 23250
rect 603 23214 632 23248
rect 666 23214 1026 23248
rect 603 23212 1026 23214
rect 603 23180 807 23212
rect 603 23146 632 23180
rect 666 23178 807 23180
rect 841 23178 1026 23212
rect 666 23146 1026 23178
rect 603 23140 1026 23146
rect 603 23112 807 23140
rect 603 23078 632 23112
rect 666 23106 807 23112
rect 841 23106 1026 23140
rect 666 23078 1026 23106
rect 603 23068 1026 23078
rect 603 23044 807 23068
rect 603 23010 632 23044
rect 666 23034 807 23044
rect 841 23034 1026 23068
rect 666 23010 1026 23034
rect 603 22996 1026 23010
rect 603 22976 807 22996
rect 603 22942 632 22976
rect 666 22962 807 22976
rect 841 22962 1026 22996
rect 666 22942 1026 22962
rect 603 22924 1026 22942
rect 603 22908 807 22924
rect 603 22874 632 22908
rect 666 22890 807 22908
rect 841 22890 1026 22924
rect 666 22874 1026 22890
rect 603 22852 1026 22874
rect 603 22840 807 22852
rect 603 22806 632 22840
rect 666 22818 807 22840
rect 841 22818 1026 22852
rect 666 22806 1026 22818
rect 603 22780 1026 22806
rect 603 22772 807 22780
rect 603 22738 632 22772
rect 666 22746 807 22772
rect 841 22746 1026 22780
rect 666 22738 1026 22746
rect 603 22708 1026 22738
rect 603 22704 807 22708
rect 603 22670 632 22704
rect 666 22674 807 22704
rect 841 22674 1026 22708
rect 666 22670 1026 22674
rect 603 22636 1026 22670
rect 603 22602 632 22636
rect 666 22602 807 22636
rect 841 22602 1026 22636
rect 603 22568 1026 22602
rect 603 22534 632 22568
rect 666 22564 1026 22568
rect 666 22534 807 22564
rect 603 22530 807 22534
rect 841 22530 1026 22564
rect 603 22500 1026 22530
rect 603 22466 632 22500
rect 666 22492 1026 22500
rect 666 22466 807 22492
rect 603 22458 807 22466
rect 841 22458 1026 22492
rect 603 22432 1026 22458
rect 603 22398 632 22432
rect 666 22420 1026 22432
rect 666 22398 807 22420
rect 603 22386 807 22398
rect 841 22386 1026 22420
rect 603 22364 1026 22386
rect 603 22330 632 22364
rect 666 22348 1026 22364
rect 666 22330 807 22348
rect 603 22314 807 22330
rect 841 22314 1026 22348
rect 603 22296 1026 22314
rect 603 22262 632 22296
rect 666 22276 1026 22296
rect 666 22262 807 22276
rect 603 22242 807 22262
rect 841 22242 1026 22276
rect 603 22228 1026 22242
rect 603 22194 632 22228
rect 666 22204 1026 22228
rect 666 22194 807 22204
rect 603 22170 807 22194
rect 841 22170 1026 22204
rect 603 22160 1026 22170
rect 603 22126 632 22160
rect 666 22132 1026 22160
rect 666 22126 807 22132
rect 603 22098 807 22126
rect 841 22098 1026 22132
rect 603 22092 1026 22098
rect 603 22058 632 22092
rect 666 22060 1026 22092
rect 666 22058 807 22060
rect 603 22026 807 22058
rect 841 22026 1026 22060
rect 603 22024 1026 22026
rect 603 21990 632 22024
rect 666 21990 1026 22024
rect 603 21988 1026 21990
rect 603 21956 807 21988
rect 603 21922 632 21956
rect 666 21954 807 21956
rect 841 21954 1026 21988
rect 666 21922 1026 21954
rect 603 21916 1026 21922
rect 603 21888 807 21916
rect 603 21854 632 21888
rect 666 21882 807 21888
rect 841 21882 1026 21916
rect 666 21854 1026 21882
rect 603 21844 1026 21854
rect 603 21820 807 21844
rect 603 21786 632 21820
rect 666 21810 807 21820
rect 841 21810 1026 21844
rect 666 21786 1026 21810
rect 603 21772 1026 21786
rect 603 21752 807 21772
rect 603 21718 632 21752
rect 666 21738 807 21752
rect 841 21738 1026 21772
rect 666 21718 1026 21738
rect 603 21700 1026 21718
rect 603 21684 807 21700
rect 603 21650 632 21684
rect 666 21666 807 21684
rect 841 21666 1026 21700
rect 666 21650 1026 21666
rect 603 21628 1026 21650
rect 603 21616 807 21628
rect 603 21582 632 21616
rect 666 21594 807 21616
rect 841 21594 1026 21628
rect 666 21582 1026 21594
rect 603 21556 1026 21582
rect 603 21548 807 21556
rect 603 21514 632 21548
rect 666 21522 807 21548
rect 841 21522 1026 21556
rect 666 21514 1026 21522
rect 603 21484 1026 21514
rect 603 21480 807 21484
rect 603 21446 632 21480
rect 666 21450 807 21480
rect 841 21450 1026 21484
rect 666 21446 1026 21450
rect 603 21412 1026 21446
rect 603 21378 632 21412
rect 666 21378 807 21412
rect 841 21378 1026 21412
rect 603 21344 1026 21378
rect 603 21310 632 21344
rect 666 21340 1026 21344
rect 666 21310 807 21340
rect 603 21306 807 21310
rect 841 21306 1026 21340
rect 603 21276 1026 21306
rect 603 21242 632 21276
rect 666 21268 1026 21276
rect 666 21242 807 21268
rect 603 21234 807 21242
rect 841 21234 1026 21268
rect 603 21208 1026 21234
rect 603 21174 632 21208
rect 666 21196 1026 21208
rect 666 21174 807 21196
rect 603 21162 807 21174
rect 841 21162 1026 21196
rect 603 21140 1026 21162
rect 603 21106 632 21140
rect 666 21124 1026 21140
rect 666 21106 807 21124
rect 603 21090 807 21106
rect 841 21090 1026 21124
rect 603 21072 1026 21090
rect 603 21038 632 21072
rect 666 21052 1026 21072
rect 666 21038 807 21052
rect 603 21018 807 21038
rect 841 21018 1026 21052
rect 603 21004 1026 21018
rect 603 20970 632 21004
rect 666 20980 1026 21004
rect 666 20970 807 20980
rect 603 20946 807 20970
rect 841 20946 1026 20980
rect 603 20936 1026 20946
rect 603 20902 632 20936
rect 666 20908 1026 20936
rect 666 20902 807 20908
rect 603 20874 807 20902
rect 841 20874 1026 20908
rect 603 20868 1026 20874
rect 603 20834 632 20868
rect 666 20836 1026 20868
rect 666 20834 807 20836
rect 603 20802 807 20834
rect 841 20802 1026 20836
rect 603 20800 1026 20802
rect 603 20766 632 20800
rect 666 20766 1026 20800
rect 603 20764 1026 20766
rect 603 20732 807 20764
rect 603 20698 632 20732
rect 666 20730 807 20732
rect 841 20730 1026 20764
rect 666 20698 1026 20730
rect 603 20692 1026 20698
rect 603 20664 807 20692
rect 603 20630 632 20664
rect 666 20658 807 20664
rect 841 20658 1026 20692
rect 666 20630 1026 20658
rect 603 20620 1026 20630
rect 603 20596 807 20620
rect 603 20562 632 20596
rect 666 20586 807 20596
rect 841 20586 1026 20620
rect 666 20562 1026 20586
rect 603 20548 1026 20562
rect 603 20528 807 20548
rect 603 20494 632 20528
rect 666 20514 807 20528
rect 841 20514 1026 20548
rect 666 20494 1026 20514
rect 603 20476 1026 20494
rect 603 20460 807 20476
rect 603 20426 632 20460
rect 666 20442 807 20460
rect 841 20442 1026 20476
rect 666 20426 1026 20442
rect 603 20404 1026 20426
rect 603 20392 807 20404
rect 603 20358 632 20392
rect 666 20370 807 20392
rect 841 20370 1026 20404
rect 666 20358 1026 20370
rect 603 20332 1026 20358
rect 603 20324 807 20332
rect 603 20290 632 20324
rect 666 20298 807 20324
rect 841 20298 1026 20332
rect 666 20290 1026 20298
rect 603 20260 1026 20290
rect 603 20256 807 20260
rect 603 20222 632 20256
rect 666 20226 807 20256
rect 841 20226 1026 20260
rect 666 20222 1026 20226
rect 603 20188 1026 20222
rect 603 20154 632 20188
rect 666 20154 807 20188
rect 841 20154 1026 20188
rect 603 20120 1026 20154
rect 603 20086 632 20120
rect 666 20116 1026 20120
rect 666 20086 807 20116
rect 603 20082 807 20086
rect 841 20082 1026 20116
rect 603 20052 1026 20082
rect 603 20018 632 20052
rect 666 20044 1026 20052
rect 666 20018 807 20044
rect 603 20010 807 20018
rect 841 20010 1026 20044
rect 603 19984 1026 20010
rect 603 19950 632 19984
rect 666 19972 1026 19984
rect 666 19950 807 19972
rect 603 19938 807 19950
rect 841 19938 1026 19972
rect 603 19916 1026 19938
rect 603 19882 632 19916
rect 666 19900 1026 19916
rect 666 19882 807 19900
rect 603 19866 807 19882
rect 841 19866 1026 19900
rect 603 19848 1026 19866
rect 603 19814 632 19848
rect 666 19828 1026 19848
rect 666 19814 807 19828
rect 603 19794 807 19814
rect 841 19794 1026 19828
rect 603 19780 1026 19794
rect 603 19746 632 19780
rect 666 19756 1026 19780
rect 666 19746 807 19756
rect 603 19722 807 19746
rect 841 19722 1026 19756
rect 603 19712 1026 19722
rect 603 19678 632 19712
rect 666 19684 1026 19712
rect 666 19678 807 19684
rect 603 19650 807 19678
rect 841 19650 1026 19684
rect 603 19644 1026 19650
rect 603 19610 632 19644
rect 666 19612 1026 19644
rect 666 19610 807 19612
rect 603 19578 807 19610
rect 841 19578 1026 19612
rect 603 19576 1026 19578
rect 603 19542 632 19576
rect 666 19542 1026 19576
rect 603 19540 1026 19542
rect 603 19508 807 19540
rect 603 19474 632 19508
rect 666 19506 807 19508
rect 841 19506 1026 19540
rect 666 19474 1026 19506
rect 603 19468 1026 19474
rect 603 19440 807 19468
rect 603 19406 632 19440
rect 666 19434 807 19440
rect 841 19434 1026 19468
rect 666 19406 1026 19434
rect 603 19396 1026 19406
rect 603 19372 807 19396
rect 603 19338 632 19372
rect 666 19362 807 19372
rect 841 19362 1026 19396
rect 666 19338 1026 19362
rect 603 19324 1026 19338
rect 603 19304 807 19324
rect 603 19270 632 19304
rect 666 19290 807 19304
rect 841 19290 1026 19324
rect 666 19270 1026 19290
rect 603 19252 1026 19270
rect 603 19236 807 19252
rect 603 19202 632 19236
rect 666 19218 807 19236
rect 841 19218 1026 19252
rect 666 19202 1026 19218
rect 603 19180 1026 19202
rect 603 19168 807 19180
rect 603 19134 632 19168
rect 666 19146 807 19168
rect 841 19146 1026 19180
rect 666 19134 1026 19146
rect 603 19108 1026 19134
rect 603 19100 807 19108
rect 603 19066 632 19100
rect 666 19074 807 19100
rect 841 19074 1026 19108
rect 666 19066 1026 19074
rect 603 19036 1026 19066
rect 603 19032 807 19036
rect 603 18998 632 19032
rect 666 19002 807 19032
rect 841 19002 1026 19036
rect 666 18998 1026 19002
rect 603 18964 1026 18998
rect 603 18930 632 18964
rect 666 18930 807 18964
rect 841 18930 1026 18964
rect 603 18896 1026 18930
rect 603 18862 632 18896
rect 666 18892 1026 18896
rect 666 18862 807 18892
rect 603 18858 807 18862
rect 841 18858 1026 18892
rect 603 18828 1026 18858
rect 603 18794 632 18828
rect 666 18820 1026 18828
rect 666 18794 807 18820
rect 603 18786 807 18794
rect 841 18786 1026 18820
rect 603 18760 1026 18786
rect 603 18726 632 18760
rect 666 18748 1026 18760
rect 666 18726 807 18748
rect 603 18714 807 18726
rect 841 18714 1026 18748
rect 603 18692 1026 18714
rect 603 18658 632 18692
rect 666 18676 1026 18692
rect 666 18658 807 18676
rect 603 18642 807 18658
rect 841 18642 1026 18676
rect 603 18624 1026 18642
rect 603 18590 632 18624
rect 666 18604 1026 18624
rect 666 18590 807 18604
rect 603 18570 807 18590
rect 841 18570 1026 18604
rect 603 18556 1026 18570
rect 603 18522 632 18556
rect 666 18532 1026 18556
rect 666 18522 807 18532
rect 603 18498 807 18522
rect 841 18498 1026 18532
rect 603 18488 1026 18498
rect 603 18454 632 18488
rect 666 18460 1026 18488
rect 666 18454 807 18460
rect 603 18426 807 18454
rect 841 18426 1026 18460
rect 603 18420 1026 18426
rect 603 18386 632 18420
rect 666 18388 1026 18420
rect 666 18386 807 18388
rect 603 18354 807 18386
rect 841 18354 1026 18388
rect 603 18352 1026 18354
rect 603 18318 632 18352
rect 666 18318 1026 18352
rect 603 18316 1026 18318
rect 603 18284 807 18316
rect 603 18250 632 18284
rect 666 18282 807 18284
rect 841 18282 1026 18316
rect 666 18250 1026 18282
rect 603 18244 1026 18250
rect 603 18216 807 18244
rect 603 18182 632 18216
rect 666 18210 807 18216
rect 841 18210 1026 18244
rect 666 18182 1026 18210
rect 603 18172 1026 18182
rect 603 18148 807 18172
rect 603 18114 632 18148
rect 666 18138 807 18148
rect 841 18138 1026 18172
rect 666 18114 1026 18138
rect 603 18100 1026 18114
rect 603 18080 807 18100
rect 603 18046 632 18080
rect 666 18066 807 18080
rect 841 18066 1026 18100
rect 666 18046 1026 18066
rect 603 18028 1026 18046
rect 603 18012 807 18028
rect 603 17978 632 18012
rect 666 17994 807 18012
rect 841 17994 1026 18028
rect 666 17978 1026 17994
rect 603 17956 1026 17978
rect 603 17944 807 17956
rect 603 17910 632 17944
rect 666 17922 807 17944
rect 841 17922 1026 17956
rect 666 17910 1026 17922
rect 603 17884 1026 17910
rect 603 17876 807 17884
rect 603 17842 632 17876
rect 666 17850 807 17876
rect 841 17850 1026 17884
rect 666 17842 1026 17850
rect 603 17812 1026 17842
rect 603 17808 807 17812
rect 603 17774 632 17808
rect 666 17778 807 17808
rect 841 17778 1026 17812
rect 666 17774 1026 17778
rect 603 17740 1026 17774
rect 603 17706 632 17740
rect 666 17706 807 17740
rect 841 17706 1026 17740
rect 603 17672 1026 17706
rect 603 17638 632 17672
rect 666 17668 1026 17672
rect 666 17638 807 17668
rect 603 17634 807 17638
rect 841 17634 1026 17668
rect 603 17604 1026 17634
rect 603 17570 632 17604
rect 666 17596 1026 17604
rect 666 17570 807 17596
rect 603 17562 807 17570
rect 841 17562 1026 17596
rect 603 17536 1026 17562
rect 603 17502 632 17536
rect 666 17524 1026 17536
rect 666 17502 807 17524
rect 603 17490 807 17502
rect 841 17490 1026 17524
rect 603 17468 1026 17490
rect 603 17434 632 17468
rect 666 17452 1026 17468
rect 666 17434 807 17452
rect 603 17418 807 17434
rect 841 17418 1026 17452
rect 603 17400 1026 17418
rect 603 17366 632 17400
rect 666 17380 1026 17400
rect 666 17366 807 17380
rect 603 17346 807 17366
rect 841 17346 1026 17380
rect 603 17332 1026 17346
rect 603 17298 632 17332
rect 666 17308 1026 17332
rect 666 17298 807 17308
rect 603 17274 807 17298
rect 841 17274 1026 17308
rect 603 17264 1026 17274
rect 603 17230 632 17264
rect 666 17236 1026 17264
rect 666 17230 807 17236
rect 603 17202 807 17230
rect 841 17202 1026 17236
rect 603 17196 1026 17202
rect 603 17162 632 17196
rect 666 17164 1026 17196
rect 666 17162 807 17164
rect 603 17130 807 17162
rect 841 17130 1026 17164
rect 603 17128 1026 17130
rect 603 17094 632 17128
rect 666 17094 1026 17128
rect 603 17092 1026 17094
rect 603 17060 807 17092
rect 603 17026 632 17060
rect 666 17058 807 17060
rect 841 17058 1026 17092
rect 666 17026 1026 17058
rect 603 17020 1026 17026
rect 603 16992 807 17020
rect 603 16958 632 16992
rect 666 16986 807 16992
rect 841 16986 1026 17020
rect 666 16958 1026 16986
rect 603 16948 1026 16958
rect 603 16924 807 16948
rect 603 16890 632 16924
rect 666 16914 807 16924
rect 841 16914 1026 16948
rect 666 16890 1026 16914
rect 603 16876 1026 16890
rect 603 16856 807 16876
rect 603 16822 632 16856
rect 666 16842 807 16856
rect 841 16842 1026 16876
rect 666 16822 1026 16842
rect 603 16804 1026 16822
rect 603 16788 807 16804
rect 603 16754 632 16788
rect 666 16770 807 16788
rect 841 16770 1026 16804
rect 666 16754 1026 16770
rect 603 16732 1026 16754
rect 603 16720 807 16732
rect 603 16686 632 16720
rect 666 16698 807 16720
rect 841 16698 1026 16732
rect 666 16686 1026 16698
rect 603 16660 1026 16686
rect 603 16652 807 16660
rect 603 16618 632 16652
rect 666 16626 807 16652
rect 841 16626 1026 16660
rect 666 16618 1026 16626
rect 603 16588 1026 16618
rect 603 16584 807 16588
rect 603 16550 632 16584
rect 666 16554 807 16584
rect 841 16554 1026 16588
rect 666 16550 1026 16554
rect 603 16516 1026 16550
rect 603 16482 632 16516
rect 666 16482 807 16516
rect 841 16482 1026 16516
rect 603 16448 1026 16482
rect 603 16414 632 16448
rect 666 16444 1026 16448
rect 666 16414 807 16444
rect 603 16410 807 16414
rect 841 16410 1026 16444
rect 603 16380 1026 16410
rect 603 16346 632 16380
rect 666 16372 1026 16380
rect 666 16346 807 16372
rect 603 16338 807 16346
rect 841 16338 1026 16372
rect 603 16312 1026 16338
rect 603 16278 632 16312
rect 666 16300 1026 16312
rect 666 16278 807 16300
rect 603 16266 807 16278
rect 841 16266 1026 16300
rect 603 16244 1026 16266
rect 603 16210 632 16244
rect 666 16228 1026 16244
rect 666 16210 807 16228
rect 603 16194 807 16210
rect 841 16194 1026 16228
rect 603 16176 1026 16194
rect 603 16142 632 16176
rect 666 16156 1026 16176
rect 666 16142 807 16156
rect 603 16122 807 16142
rect 841 16122 1026 16156
rect 603 16108 1026 16122
rect 603 16074 632 16108
rect 666 16084 1026 16108
rect 666 16074 807 16084
rect 603 16050 807 16074
rect 841 16050 1026 16084
rect 603 16040 1026 16050
rect 603 16006 632 16040
rect 666 16012 1026 16040
rect 666 16006 807 16012
rect 603 15978 807 16006
rect 841 15978 1026 16012
rect 603 15972 1026 15978
rect 603 15938 632 15972
rect 666 15940 1026 15972
rect 666 15938 807 15940
rect 603 15906 807 15938
rect 841 15906 1026 15940
rect 603 15904 1026 15906
rect 603 15870 632 15904
rect 666 15870 1026 15904
rect 603 15868 1026 15870
rect 603 15836 807 15868
rect 603 15802 632 15836
rect 666 15834 807 15836
rect 841 15834 1026 15868
rect 666 15802 1026 15834
rect 603 15796 1026 15802
rect 603 15768 807 15796
rect 603 15734 632 15768
rect 666 15762 807 15768
rect 841 15762 1026 15796
rect 666 15734 1026 15762
rect 603 15724 1026 15734
rect 603 15700 807 15724
rect 603 15666 632 15700
rect 666 15690 807 15700
rect 841 15690 1026 15724
rect 666 15666 1026 15690
rect 603 15652 1026 15666
rect 603 15632 807 15652
rect 603 15598 632 15632
rect 666 15618 807 15632
rect 841 15618 1026 15652
rect 666 15598 1026 15618
rect 603 15580 1026 15598
rect 603 15564 807 15580
rect 603 15530 632 15564
rect 666 15546 807 15564
rect 841 15546 1026 15580
rect 666 15530 1026 15546
rect 603 15508 1026 15530
rect 603 15496 807 15508
rect 603 15462 632 15496
rect 666 15474 807 15496
rect 841 15474 1026 15508
rect 666 15462 1026 15474
rect 603 15436 1026 15462
rect 603 15428 807 15436
rect 603 15394 632 15428
rect 666 15402 807 15428
rect 841 15402 1026 15436
rect 666 15394 1026 15402
rect 603 15364 1026 15394
rect 603 15360 807 15364
rect 603 15326 632 15360
rect 666 15330 807 15360
rect 841 15330 1026 15364
rect 666 15326 1026 15330
rect 603 15292 1026 15326
rect 603 15258 632 15292
rect 666 15258 807 15292
rect 841 15258 1026 15292
rect 603 15224 1026 15258
rect 603 15190 632 15224
rect 666 15220 1026 15224
rect 666 15190 807 15220
rect 603 15186 807 15190
rect 841 15186 1026 15220
rect 603 15156 1026 15186
rect 603 15122 632 15156
rect 666 15148 1026 15156
rect 666 15122 807 15148
rect 603 15114 807 15122
rect 841 15114 1026 15148
rect 603 15088 1026 15114
rect 603 15054 632 15088
rect 666 15076 1026 15088
rect 666 15054 807 15076
rect 603 15042 807 15054
rect 841 15042 1026 15076
rect 603 15020 1026 15042
rect 603 14986 632 15020
rect 666 15004 1026 15020
rect 666 14986 807 15004
rect 603 14970 807 14986
rect 841 14970 1026 15004
rect 603 14952 1026 14970
rect 603 14918 632 14952
rect 666 14932 1026 14952
rect 666 14918 807 14932
rect 603 14898 807 14918
rect 841 14898 1026 14932
rect 603 14884 1026 14898
rect 603 14850 632 14884
rect 666 14860 1026 14884
rect 666 14850 807 14860
rect 603 14826 807 14850
rect 841 14826 1026 14860
rect 603 14816 1026 14826
rect 603 14782 632 14816
rect 666 14788 1026 14816
rect 666 14782 807 14788
rect 603 14754 807 14782
rect 841 14754 1026 14788
rect 603 14748 1026 14754
rect 603 14714 632 14748
rect 666 14716 1026 14748
rect 666 14714 807 14716
rect 603 14682 807 14714
rect 841 14682 1026 14716
rect 603 14680 1026 14682
rect 603 14646 632 14680
rect 666 14646 1026 14680
rect 603 14644 1026 14646
rect 603 14612 807 14644
rect 603 14578 632 14612
rect 666 14610 807 14612
rect 841 14610 1026 14644
rect 666 14578 1026 14610
rect 603 14572 1026 14578
rect 603 14544 807 14572
rect 603 14510 632 14544
rect 666 14538 807 14544
rect 841 14538 1026 14572
rect 666 14510 1026 14538
rect 603 14500 1026 14510
rect 603 14476 807 14500
rect 603 14442 632 14476
rect 666 14466 807 14476
rect 841 14466 1026 14500
rect 666 14442 1026 14466
rect 603 14428 1026 14442
rect 603 14408 807 14428
rect 603 14374 632 14408
rect 666 14394 807 14408
rect 841 14394 1026 14428
rect 666 14374 1026 14394
rect 603 14356 1026 14374
rect 603 14340 807 14356
rect 603 14306 632 14340
rect 666 14322 807 14340
rect 841 14322 1026 14356
rect 666 14306 1026 14322
rect 603 14284 1026 14306
rect 603 14272 807 14284
rect 603 14238 632 14272
rect 666 14250 807 14272
rect 841 14250 1026 14284
rect 666 14238 1026 14250
rect 603 14212 1026 14238
rect 603 14204 807 14212
rect 603 14170 632 14204
rect 666 14178 807 14204
rect 841 14178 1026 14212
rect 666 14170 1026 14178
rect 603 14140 1026 14170
rect 603 14136 807 14140
rect 603 14102 632 14136
rect 666 14106 807 14136
rect 841 14106 1026 14140
rect 666 14102 1026 14106
rect 603 14068 1026 14102
rect 603 14034 632 14068
rect 666 14034 807 14068
rect 841 14034 1026 14068
rect 603 14000 1026 14034
rect 603 13966 632 14000
rect 666 13996 1026 14000
rect 666 13966 807 13996
rect 603 13962 807 13966
rect 841 13962 1026 13996
rect 603 13932 1026 13962
rect 603 13898 632 13932
rect 666 13924 1026 13932
rect 666 13898 807 13924
rect 603 13890 807 13898
rect 841 13890 1026 13924
rect 603 13864 1026 13890
rect 603 13830 632 13864
rect 666 13852 1026 13864
rect 666 13830 807 13852
rect 603 13818 807 13830
rect 841 13818 1026 13852
rect 603 13796 1026 13818
rect 603 13762 632 13796
rect 666 13780 1026 13796
rect 666 13762 807 13780
rect 603 13746 807 13762
rect 841 13746 1026 13780
rect 603 13728 1026 13746
rect 603 13694 632 13728
rect 666 13708 1026 13728
rect 666 13694 807 13708
rect 603 13674 807 13694
rect 841 13674 1026 13708
rect 603 13660 1026 13674
rect 603 13626 632 13660
rect 666 13636 1026 13660
rect 666 13626 807 13636
rect 603 13602 807 13626
rect 841 13602 1026 13636
rect 603 13592 1026 13602
rect 603 13558 632 13592
rect 666 13564 1026 13592
rect 666 13558 807 13564
rect 603 13530 807 13558
rect 841 13530 1026 13564
rect 603 13524 1026 13530
rect 603 13490 632 13524
rect 666 13492 1026 13524
rect 666 13490 807 13492
rect 603 13458 807 13490
rect 841 13458 1026 13492
rect 603 13456 1026 13458
rect 603 13422 632 13456
rect 666 13422 1026 13456
rect 603 13420 1026 13422
rect 603 13388 807 13420
rect 603 13354 632 13388
rect 666 13386 807 13388
rect 841 13386 1026 13420
rect 666 13354 1026 13386
rect 603 13348 1026 13354
rect 603 13320 807 13348
rect 603 13286 632 13320
rect 666 13314 807 13320
rect 841 13314 1026 13348
rect 666 13286 1026 13314
rect 603 13276 1026 13286
rect 603 13252 807 13276
rect 603 13218 632 13252
rect 666 13242 807 13252
rect 841 13242 1026 13276
rect 666 13218 1026 13242
rect 603 13204 1026 13218
rect 603 13184 807 13204
rect 603 13150 632 13184
rect 666 13170 807 13184
rect 841 13170 1026 13204
rect 666 13150 1026 13170
rect 603 13132 1026 13150
rect 603 13116 807 13132
rect 603 13082 632 13116
rect 666 13098 807 13116
rect 841 13098 1026 13132
rect 666 13082 1026 13098
rect 603 13060 1026 13082
rect 603 13048 807 13060
rect 603 13014 632 13048
rect 666 13026 807 13048
rect 841 13026 1026 13060
rect 666 13014 1026 13026
rect 603 12988 1026 13014
rect 603 12980 807 12988
rect 603 12946 632 12980
rect 666 12954 807 12980
rect 841 12954 1026 12988
rect 666 12946 1026 12954
rect 603 12916 1026 12946
rect 603 12912 807 12916
rect 603 12878 632 12912
rect 666 12882 807 12912
rect 841 12882 1026 12916
rect 666 12878 1026 12882
rect 603 12844 1026 12878
rect 603 12810 632 12844
rect 666 12810 807 12844
rect 841 12810 1026 12844
rect 603 12776 1026 12810
rect 603 12742 632 12776
rect 666 12772 1026 12776
rect 666 12742 807 12772
rect 603 12738 807 12742
rect 841 12738 1026 12772
rect 603 12708 1026 12738
rect 603 12674 632 12708
rect 666 12700 1026 12708
rect 666 12674 807 12700
rect 603 12666 807 12674
rect 841 12666 1026 12700
rect 603 12640 1026 12666
rect 603 12606 632 12640
rect 666 12628 1026 12640
rect 666 12606 807 12628
rect 603 12594 807 12606
rect 841 12594 1026 12628
rect 603 12572 1026 12594
rect 603 12538 632 12572
rect 666 12556 1026 12572
rect 666 12538 807 12556
rect 603 12522 807 12538
rect 841 12522 1026 12556
rect 603 12504 1026 12522
rect 603 12470 632 12504
rect 666 12484 1026 12504
rect 666 12470 807 12484
rect 603 12450 807 12470
rect 841 12450 1026 12484
rect 603 12436 1026 12450
rect 603 12402 632 12436
rect 666 12412 1026 12436
rect 666 12402 807 12412
rect 603 12378 807 12402
rect 841 12378 1026 12412
rect 603 12368 1026 12378
rect 603 12334 632 12368
rect 666 12340 1026 12368
rect 666 12334 807 12340
rect 603 12306 807 12334
rect 841 12306 1026 12340
rect 603 12300 1026 12306
rect 603 12266 632 12300
rect 666 12268 1026 12300
rect 666 12266 807 12268
rect 603 12234 807 12266
rect 841 12234 1026 12268
rect 603 12232 1026 12234
rect 603 12198 632 12232
rect 666 12198 1026 12232
rect 603 12196 1026 12198
rect 603 12164 807 12196
rect 603 12130 632 12164
rect 666 12162 807 12164
rect 841 12162 1026 12196
rect 666 12130 1026 12162
rect 603 12124 1026 12130
rect 603 12096 807 12124
rect 603 12062 632 12096
rect 666 12090 807 12096
rect 841 12090 1026 12124
rect 666 12062 1026 12090
rect 603 12052 1026 12062
rect 603 12028 807 12052
rect 603 11994 632 12028
rect 666 12018 807 12028
rect 841 12018 1026 12052
rect 666 11994 1026 12018
rect 603 11980 1026 11994
rect 603 11960 807 11980
rect 603 11926 632 11960
rect 666 11946 807 11960
rect 841 11946 1026 11980
rect 666 11926 1026 11946
rect 603 11908 1026 11926
rect 603 11892 807 11908
rect 603 11858 632 11892
rect 666 11874 807 11892
rect 841 11874 1026 11908
rect 666 11858 1026 11874
rect 603 11836 1026 11858
rect 603 11824 807 11836
rect 603 11790 632 11824
rect 666 11802 807 11824
rect 841 11802 1026 11836
rect 666 11790 1026 11802
rect 603 11764 1026 11790
rect 603 11756 807 11764
rect 603 11722 632 11756
rect 666 11730 807 11756
rect 841 11730 1026 11764
rect 666 11722 1026 11730
rect 603 11692 1026 11722
rect 603 11688 807 11692
rect 603 11654 632 11688
rect 666 11658 807 11688
rect 841 11658 1026 11692
rect 666 11654 1026 11658
rect 603 11620 1026 11654
rect 603 11586 632 11620
rect 666 11586 807 11620
rect 841 11586 1026 11620
rect 603 11552 1026 11586
rect 603 11518 632 11552
rect 666 11548 1026 11552
rect 666 11518 807 11548
rect 603 11514 807 11518
rect 841 11514 1026 11548
rect 603 11484 1026 11514
rect 603 11450 632 11484
rect 666 11476 1026 11484
rect 666 11450 807 11476
rect 603 11442 807 11450
rect 841 11442 1026 11476
rect 603 11416 1026 11442
rect 603 11382 632 11416
rect 666 11404 1026 11416
rect 666 11382 807 11404
rect 603 11370 807 11382
rect 841 11370 1026 11404
rect 603 11348 1026 11370
rect 603 11314 632 11348
rect 666 11332 1026 11348
rect 666 11314 807 11332
rect 603 11298 807 11314
rect 841 11298 1026 11332
rect 603 11280 1026 11298
rect 603 11246 632 11280
rect 666 11260 1026 11280
rect 666 11246 807 11260
rect 603 11226 807 11246
rect 841 11226 1026 11260
rect 603 11212 1026 11226
rect 603 11178 632 11212
rect 666 11188 1026 11212
rect 666 11178 807 11188
rect 603 11154 807 11178
rect 841 11154 1026 11188
rect 603 11144 1026 11154
rect 603 11110 632 11144
rect 666 11116 1026 11144
rect 666 11110 807 11116
rect 603 11082 807 11110
rect 841 11082 1026 11116
rect 603 11076 1026 11082
rect 603 11042 632 11076
rect 666 11044 1026 11076
rect 666 11042 807 11044
rect 603 11010 807 11042
rect 841 11010 1026 11044
rect 603 11008 1026 11010
rect 603 10974 632 11008
rect 666 10974 1026 11008
rect 603 10972 1026 10974
rect 603 10940 807 10972
rect 603 10906 632 10940
rect 666 10938 807 10940
rect 841 10938 1026 10972
rect 666 10906 1026 10938
rect 603 10900 1026 10906
rect 603 10872 807 10900
rect 603 10838 632 10872
rect 666 10866 807 10872
rect 841 10866 1026 10900
rect 666 10838 1026 10866
rect 603 10828 1026 10838
rect 603 10804 807 10828
rect 603 10770 632 10804
rect 666 10794 807 10804
rect 841 10794 1026 10828
rect 666 10770 1026 10794
rect 603 10756 1026 10770
rect 603 10736 807 10756
rect 603 10702 632 10736
rect 666 10722 807 10736
rect 841 10722 1026 10756
rect 666 10702 1026 10722
rect 603 10684 1026 10702
rect 603 10668 807 10684
rect 603 10634 632 10668
rect 666 10650 807 10668
rect 841 10650 1026 10684
rect 666 10634 1026 10650
rect 603 10612 1026 10634
rect 603 10600 807 10612
rect 603 10566 632 10600
rect 666 10578 807 10600
rect 841 10578 1026 10612
rect 666 10566 1026 10578
rect 603 10540 1026 10566
rect 603 10532 807 10540
rect 603 10498 632 10532
rect 666 10506 807 10532
rect 841 10506 1026 10540
rect 666 10498 1026 10506
rect 603 10468 1026 10498
rect 603 10464 807 10468
rect 603 10430 632 10464
rect 666 10434 807 10464
rect 841 10434 1026 10468
rect 666 10430 1026 10434
rect 603 10396 1026 10430
rect 603 10362 632 10396
rect 666 10362 807 10396
rect 841 10362 1026 10396
rect 603 10328 1026 10362
rect 603 10294 632 10328
rect 666 10324 1026 10328
rect 666 10294 807 10324
rect 603 10290 807 10294
rect 841 10290 1026 10324
rect 603 10260 1026 10290
rect 603 10226 632 10260
rect 666 10252 1026 10260
rect 666 10226 807 10252
rect 603 10218 807 10226
rect 841 10218 1026 10252
rect 603 10192 1026 10218
rect 1119 34679 13887 34721
rect 1119 34645 1301 34679
rect 1339 34645 1373 34679
rect 1407 34645 1441 34679
rect 1479 34645 1509 34679
rect 1551 34645 1577 34679
rect 1623 34645 1645 34679
rect 1695 34645 1713 34679
rect 1767 34645 1781 34679
rect 1839 34645 1849 34679
rect 1911 34645 1917 34679
rect 1983 34645 1985 34679
rect 2019 34645 2021 34679
rect 2087 34645 2093 34679
rect 2155 34645 2165 34679
rect 2223 34645 2237 34679
rect 2291 34645 2309 34679
rect 2359 34645 2381 34679
rect 2427 34645 2453 34679
rect 2495 34645 2525 34679
rect 2563 34645 2597 34679
rect 2631 34645 2665 34679
rect 2703 34645 2733 34679
rect 2775 34645 2801 34679
rect 2847 34645 2869 34679
rect 2919 34645 2937 34679
rect 2991 34645 3005 34679
rect 3063 34645 3073 34679
rect 3135 34645 3141 34679
rect 3207 34645 3209 34679
rect 3243 34645 3245 34679
rect 3311 34645 3317 34679
rect 3379 34645 3389 34679
rect 3447 34645 3461 34679
rect 3515 34645 3533 34679
rect 3583 34645 3605 34679
rect 3651 34645 3677 34679
rect 3719 34645 3749 34679
rect 3787 34645 3821 34679
rect 3855 34645 3889 34679
rect 3927 34645 3957 34679
rect 3999 34645 4025 34679
rect 4071 34645 4093 34679
rect 4143 34645 4161 34679
rect 4215 34645 4229 34679
rect 4287 34645 4297 34679
rect 4359 34645 4365 34679
rect 4431 34645 4433 34679
rect 4467 34645 4469 34679
rect 4535 34645 4541 34679
rect 4603 34645 4613 34679
rect 4671 34645 4685 34679
rect 4739 34645 4757 34679
rect 4807 34645 4829 34679
rect 4875 34645 4901 34679
rect 4943 34645 4973 34679
rect 5011 34645 5045 34679
rect 5079 34645 5113 34679
rect 5151 34645 5181 34679
rect 5223 34645 5249 34679
rect 5295 34645 5317 34679
rect 5367 34645 5385 34679
rect 5439 34645 5453 34679
rect 5511 34645 5521 34679
rect 5583 34645 5589 34679
rect 5655 34645 5657 34679
rect 5691 34645 5693 34679
rect 5759 34645 5765 34679
rect 5827 34645 5837 34679
rect 5895 34645 5909 34679
rect 5963 34645 5981 34679
rect 6031 34645 6053 34679
rect 6099 34645 6125 34679
rect 6167 34645 6197 34679
rect 6235 34645 6269 34679
rect 6303 34645 6337 34679
rect 6375 34645 6405 34679
rect 6447 34645 6473 34679
rect 6519 34645 6541 34679
rect 6591 34645 6609 34679
rect 6663 34645 6677 34679
rect 6735 34645 6745 34679
rect 6807 34645 6813 34679
rect 6879 34645 6881 34679
rect 6915 34645 6917 34679
rect 6983 34645 6989 34679
rect 7051 34645 7061 34679
rect 7119 34645 7133 34679
rect 7187 34645 7205 34679
rect 7255 34645 7277 34679
rect 7323 34645 7349 34679
rect 7391 34645 7421 34679
rect 7459 34645 7493 34679
rect 7527 34645 7561 34679
rect 7599 34645 7629 34679
rect 7671 34645 7697 34679
rect 7743 34645 7765 34679
rect 7815 34645 7833 34679
rect 7887 34645 7901 34679
rect 7959 34645 7969 34679
rect 8031 34645 8037 34679
rect 8103 34645 8105 34679
rect 8139 34645 8141 34679
rect 8207 34645 8213 34679
rect 8275 34645 8285 34679
rect 8343 34645 8357 34679
rect 8411 34645 8429 34679
rect 8479 34645 8501 34679
rect 8547 34645 8573 34679
rect 8615 34645 8645 34679
rect 8683 34645 8717 34679
rect 8751 34645 8785 34679
rect 8823 34645 8853 34679
rect 8895 34645 8921 34679
rect 8967 34645 8989 34679
rect 9039 34645 9057 34679
rect 9111 34645 9125 34679
rect 9183 34645 9193 34679
rect 9255 34645 9261 34679
rect 9327 34645 9329 34679
rect 9363 34645 9365 34679
rect 9431 34645 9437 34679
rect 9499 34645 9509 34679
rect 9567 34645 9581 34679
rect 9635 34645 9653 34679
rect 9703 34645 9725 34679
rect 9771 34645 9797 34679
rect 9839 34645 9869 34679
rect 9907 34645 9941 34679
rect 9975 34645 10009 34679
rect 10047 34645 10077 34679
rect 10119 34645 10145 34679
rect 10191 34645 10213 34679
rect 10263 34645 10281 34679
rect 10335 34645 10349 34679
rect 10407 34645 10417 34679
rect 10479 34645 10485 34679
rect 10551 34645 10553 34679
rect 10587 34645 10589 34679
rect 10655 34645 10661 34679
rect 10723 34645 10733 34679
rect 10791 34645 10805 34679
rect 10859 34645 10877 34679
rect 10927 34645 10949 34679
rect 10995 34645 11021 34679
rect 11063 34645 11093 34679
rect 11131 34645 11165 34679
rect 11199 34645 11233 34679
rect 11271 34645 11301 34679
rect 11343 34645 11369 34679
rect 11415 34645 11437 34679
rect 11487 34645 11505 34679
rect 11559 34645 11573 34679
rect 11631 34645 11641 34679
rect 11703 34645 11709 34679
rect 11775 34645 11777 34679
rect 11811 34645 11813 34679
rect 11879 34645 11885 34679
rect 11947 34645 11957 34679
rect 12015 34645 12029 34679
rect 12083 34645 12101 34679
rect 12151 34645 12173 34679
rect 12219 34645 12245 34679
rect 12287 34645 12317 34679
rect 12355 34645 12389 34679
rect 12423 34645 12457 34679
rect 12495 34645 12525 34679
rect 12567 34645 12593 34679
rect 12639 34645 12661 34679
rect 12711 34645 12729 34679
rect 12783 34645 12797 34679
rect 12855 34645 12865 34679
rect 12927 34645 12933 34679
rect 12999 34645 13001 34679
rect 13035 34645 13037 34679
rect 13103 34645 13109 34679
rect 13171 34645 13181 34679
rect 13239 34645 13253 34679
rect 13307 34645 13325 34679
rect 13375 34645 13397 34679
rect 13443 34645 13469 34679
rect 13511 34645 13541 34679
rect 13579 34645 13613 34679
rect 13647 34645 13681 34679
rect 13719 34645 13887 34679
rect 1119 34603 13887 34645
rect 1119 34478 1237 34603
rect 1119 34432 1161 34478
rect 1195 34432 1237 34478
rect 1119 34410 1237 34432
rect 1119 34360 1161 34410
rect 1195 34360 1237 34410
rect 1119 34342 1237 34360
rect 1119 34288 1161 34342
rect 1195 34288 1237 34342
rect 1119 34274 1237 34288
rect 1119 34216 1161 34274
rect 1195 34216 1237 34274
rect 1119 34206 1237 34216
rect 1119 34144 1161 34206
rect 1195 34144 1237 34206
rect 1119 34138 1237 34144
rect 1119 34072 1161 34138
rect 1195 34072 1237 34138
rect 1119 34070 1237 34072
rect 1119 34036 1161 34070
rect 1195 34036 1237 34070
rect 1119 34034 1237 34036
rect 1119 33968 1161 34034
rect 1195 33968 1237 34034
rect 1119 33962 1237 33968
rect 1119 33900 1161 33962
rect 1195 33900 1237 33962
rect 1119 33890 1237 33900
rect 1119 33832 1161 33890
rect 1195 33832 1237 33890
rect 1119 33818 1237 33832
rect 1119 33764 1161 33818
rect 1195 33764 1237 33818
rect 1119 33746 1237 33764
rect 1119 33696 1161 33746
rect 1195 33696 1237 33746
rect 1119 33674 1237 33696
rect 1119 33628 1161 33674
rect 1195 33628 1237 33674
rect 1119 33602 1237 33628
rect 1119 33560 1161 33602
rect 1195 33560 1237 33602
rect 1119 33530 1237 33560
rect 1119 33492 1161 33530
rect 1195 33492 1237 33530
rect 1119 33458 1237 33492
rect 1119 33424 1161 33458
rect 1195 33424 1237 33458
rect 1119 33390 1237 33424
rect 1119 33352 1161 33390
rect 1195 33352 1237 33390
rect 1119 33322 1237 33352
rect 1119 33280 1161 33322
rect 1195 33280 1237 33322
rect 1119 33254 1237 33280
rect 1119 33208 1161 33254
rect 1195 33208 1237 33254
rect 1119 33186 1237 33208
rect 1119 33136 1161 33186
rect 1195 33136 1237 33186
rect 1119 33118 1237 33136
rect 1119 33064 1161 33118
rect 1195 33064 1237 33118
rect 1119 33050 1237 33064
rect 1119 32992 1161 33050
rect 1195 32992 1237 33050
rect 1119 32982 1237 32992
rect 1119 32920 1161 32982
rect 1195 32920 1237 32982
rect 1119 32914 1237 32920
rect 1119 32848 1161 32914
rect 1195 32848 1237 32914
rect 1119 32846 1237 32848
rect 1119 32812 1161 32846
rect 1195 32812 1237 32846
rect 1119 32810 1237 32812
rect 1119 32744 1161 32810
rect 1195 32744 1237 32810
rect 1119 32738 1237 32744
rect 1119 32676 1161 32738
rect 1195 32676 1237 32738
rect 1119 32666 1237 32676
rect 1119 32608 1161 32666
rect 1195 32608 1237 32666
rect 1119 32594 1237 32608
rect 1119 32540 1161 32594
rect 1195 32540 1237 32594
rect 1119 32522 1237 32540
rect 1119 32472 1161 32522
rect 1195 32472 1237 32522
rect 1119 32450 1237 32472
rect 1119 32404 1161 32450
rect 1195 32404 1237 32450
rect 1119 32378 1237 32404
rect 1119 32336 1161 32378
rect 1195 32336 1237 32378
rect 1119 32306 1237 32336
rect 1119 32268 1161 32306
rect 1195 32268 1237 32306
rect 1119 32234 1237 32268
rect 1119 32200 1161 32234
rect 1195 32200 1237 32234
rect 1119 32166 1237 32200
rect 1119 32128 1161 32166
rect 1195 32128 1237 32166
rect 1119 32098 1237 32128
rect 1119 32056 1161 32098
rect 1195 32056 1237 32098
rect 1119 32030 1237 32056
rect 1119 31984 1161 32030
rect 1195 31984 1237 32030
rect 1119 31962 1237 31984
rect 1119 31912 1161 31962
rect 1195 31912 1237 31962
rect 1119 31894 1237 31912
rect 1119 31840 1161 31894
rect 1195 31840 1237 31894
rect 1119 31826 1237 31840
rect 1119 31768 1161 31826
rect 1195 31768 1237 31826
rect 1119 31758 1237 31768
rect 1119 31696 1161 31758
rect 1195 31696 1237 31758
rect 1119 31690 1237 31696
rect 1119 31624 1161 31690
rect 1195 31624 1237 31690
rect 1119 31622 1237 31624
rect 1119 31588 1161 31622
rect 1195 31588 1237 31622
rect 1119 31586 1237 31588
rect 1119 31520 1161 31586
rect 1195 31520 1237 31586
rect 1119 31514 1237 31520
rect 1119 31452 1161 31514
rect 1195 31452 1237 31514
rect 1119 31442 1237 31452
rect 1119 31384 1161 31442
rect 1195 31384 1237 31442
rect 1119 31370 1237 31384
rect 1119 31316 1161 31370
rect 1195 31316 1237 31370
rect 1119 31298 1237 31316
rect 1119 31248 1161 31298
rect 1195 31248 1237 31298
rect 1119 31226 1237 31248
rect 1119 31180 1161 31226
rect 1195 31180 1237 31226
rect 1119 31154 1237 31180
rect 1119 31112 1161 31154
rect 1195 31112 1237 31154
rect 1119 31082 1237 31112
rect 1119 31044 1161 31082
rect 1195 31044 1237 31082
rect 1119 31010 1237 31044
rect 1119 30976 1161 31010
rect 1195 30976 1237 31010
rect 1119 30942 1237 30976
rect 1119 30904 1161 30942
rect 1195 30904 1237 30942
rect 1119 30874 1237 30904
rect 1119 30832 1161 30874
rect 1195 30832 1237 30874
rect 1119 30806 1237 30832
rect 1119 30760 1161 30806
rect 1195 30760 1237 30806
rect 1119 30738 1237 30760
rect 1119 30688 1161 30738
rect 1195 30688 1237 30738
rect 1119 30670 1237 30688
rect 1119 30616 1161 30670
rect 1195 30616 1237 30670
rect 1119 30602 1237 30616
rect 1119 30544 1161 30602
rect 1195 30544 1237 30602
rect 1119 30534 1237 30544
rect 1119 30472 1161 30534
rect 1195 30472 1237 30534
rect 1119 30466 1237 30472
rect 1119 30400 1161 30466
rect 1195 30400 1237 30466
rect 1119 30398 1237 30400
rect 1119 30364 1161 30398
rect 1195 30364 1237 30398
rect 1119 30362 1237 30364
rect 1119 30296 1161 30362
rect 1195 30296 1237 30362
rect 1119 30290 1237 30296
rect 1119 30228 1161 30290
rect 1195 30228 1237 30290
rect 1119 30218 1237 30228
rect 1119 30160 1161 30218
rect 1195 30160 1237 30218
rect 1119 30146 1237 30160
rect 1119 30092 1161 30146
rect 1195 30092 1237 30146
rect 1119 30074 1237 30092
rect 1119 30024 1161 30074
rect 1195 30024 1237 30074
rect 1119 30002 1237 30024
rect 1119 29956 1161 30002
rect 1195 29956 1237 30002
rect 1119 29930 1237 29956
rect 1119 29888 1161 29930
rect 1195 29888 1237 29930
rect 1119 29858 1237 29888
rect 1119 29820 1161 29858
rect 1195 29820 1237 29858
rect 1119 29786 1237 29820
rect 1119 29752 1161 29786
rect 1195 29752 1237 29786
rect 1119 29718 1237 29752
rect 1119 29680 1161 29718
rect 1195 29680 1237 29718
rect 1119 29650 1237 29680
rect 1119 29608 1161 29650
rect 1195 29608 1237 29650
rect 1119 29582 1237 29608
rect 1119 29536 1161 29582
rect 1195 29536 1237 29582
rect 1119 29514 1237 29536
rect 1119 29464 1161 29514
rect 1195 29464 1237 29514
rect 1119 29446 1237 29464
rect 1119 29392 1161 29446
rect 1195 29392 1237 29446
rect 1119 29378 1237 29392
rect 1119 29320 1161 29378
rect 1195 29320 1237 29378
rect 1119 29310 1237 29320
rect 1119 29248 1161 29310
rect 1195 29248 1237 29310
rect 1119 29242 1237 29248
rect 1119 29176 1161 29242
rect 1195 29176 1237 29242
rect 1119 29174 1237 29176
rect 1119 29140 1161 29174
rect 1195 29140 1237 29174
rect 1119 29138 1237 29140
rect 1119 29072 1161 29138
rect 1195 29072 1237 29138
rect 1119 29066 1237 29072
rect 1119 29004 1161 29066
rect 1195 29004 1237 29066
rect 1119 28994 1237 29004
rect 1119 28936 1161 28994
rect 1195 28936 1237 28994
rect 1119 28922 1237 28936
rect 1119 28868 1161 28922
rect 1195 28868 1237 28922
rect 13769 34474 13887 34603
rect 13769 34439 13809 34474
rect 13843 34439 13887 34474
rect 13769 34405 13887 34439
rect 13769 34368 13809 34405
rect 13843 34368 13887 34405
rect 13769 34337 13887 34368
rect 13769 34296 13809 34337
rect 13843 34296 13887 34337
rect 13769 34269 13887 34296
rect 13769 34224 13809 34269
rect 13843 34224 13887 34269
rect 13769 34201 13887 34224
rect 13769 34152 13809 34201
rect 13843 34152 13887 34201
rect 13769 34133 13887 34152
rect 13769 34080 13809 34133
rect 13843 34080 13887 34133
rect 13769 34065 13887 34080
rect 13769 34008 13809 34065
rect 13843 34008 13887 34065
rect 13769 33997 13887 34008
rect 13769 33936 13809 33997
rect 13843 33936 13887 33997
rect 13769 33929 13887 33936
rect 13769 33864 13809 33929
rect 13843 33864 13887 33929
rect 13769 33861 13887 33864
rect 13769 33827 13809 33861
rect 13843 33827 13887 33861
rect 13769 33826 13887 33827
rect 13769 33759 13809 33826
rect 13843 33759 13887 33826
rect 13769 33754 13887 33759
rect 13769 33691 13809 33754
rect 13843 33691 13887 33754
rect 13769 33682 13887 33691
rect 13769 33623 13809 33682
rect 13843 33623 13887 33682
rect 13769 33610 13887 33623
rect 13769 33555 13809 33610
rect 13843 33555 13887 33610
rect 13769 33538 13887 33555
rect 13769 33487 13809 33538
rect 13843 33487 13887 33538
rect 13769 33466 13887 33487
rect 13769 33419 13809 33466
rect 13843 33419 13887 33466
rect 13769 33394 13887 33419
rect 13769 33351 13809 33394
rect 13843 33351 13887 33394
rect 13769 33322 13887 33351
rect 13769 33283 13809 33322
rect 13843 33283 13887 33322
rect 13769 33250 13887 33283
rect 13769 33215 13809 33250
rect 13843 33215 13887 33250
rect 13769 33181 13887 33215
rect 13769 33144 13809 33181
rect 13843 33144 13887 33181
rect 13769 33113 13887 33144
rect 13769 33072 13809 33113
rect 13843 33072 13887 33113
rect 13769 33045 13887 33072
rect 13769 33000 13809 33045
rect 13843 33000 13887 33045
rect 13769 32977 13887 33000
rect 13769 32928 13809 32977
rect 13843 32928 13887 32977
rect 13769 32909 13887 32928
rect 13769 32856 13809 32909
rect 13843 32856 13887 32909
rect 13769 32841 13887 32856
rect 13769 32784 13809 32841
rect 13843 32784 13887 32841
rect 13769 32773 13887 32784
rect 13769 32712 13809 32773
rect 13843 32712 13887 32773
rect 13769 32705 13887 32712
rect 13769 32640 13809 32705
rect 13843 32640 13887 32705
rect 13769 32637 13887 32640
rect 13769 32603 13809 32637
rect 13843 32603 13887 32637
rect 13769 32602 13887 32603
rect 13769 32535 13809 32602
rect 13843 32535 13887 32602
rect 13769 32530 13887 32535
rect 13769 32467 13809 32530
rect 13843 32467 13887 32530
rect 13769 32458 13887 32467
rect 13769 32399 13809 32458
rect 13843 32399 13887 32458
rect 13769 32386 13887 32399
rect 13769 32331 13809 32386
rect 13843 32331 13887 32386
rect 13769 32314 13887 32331
rect 13769 32263 13809 32314
rect 13843 32263 13887 32314
rect 13769 32242 13887 32263
rect 13769 32195 13809 32242
rect 13843 32195 13887 32242
rect 13769 32170 13887 32195
rect 13769 32127 13809 32170
rect 13843 32127 13887 32170
rect 13769 32098 13887 32127
rect 13769 32059 13809 32098
rect 13843 32059 13887 32098
rect 13769 32026 13887 32059
rect 13769 31991 13809 32026
rect 13843 31991 13887 32026
rect 13769 31957 13887 31991
rect 13769 31920 13809 31957
rect 13843 31920 13887 31957
rect 13769 31889 13887 31920
rect 13769 31848 13809 31889
rect 13843 31848 13887 31889
rect 13769 31821 13887 31848
rect 13769 31776 13809 31821
rect 13843 31776 13887 31821
rect 13769 31753 13887 31776
rect 13769 31704 13809 31753
rect 13843 31704 13887 31753
rect 13769 31685 13887 31704
rect 13769 31632 13809 31685
rect 13843 31632 13887 31685
rect 13769 31617 13887 31632
rect 13769 31560 13809 31617
rect 13843 31560 13887 31617
rect 13769 31549 13887 31560
rect 13769 31488 13809 31549
rect 13843 31488 13887 31549
rect 13769 31481 13887 31488
rect 13769 31416 13809 31481
rect 13843 31416 13887 31481
rect 13769 31413 13887 31416
rect 13769 31379 13809 31413
rect 13843 31379 13887 31413
rect 13769 31378 13887 31379
rect 13769 31311 13809 31378
rect 13843 31311 13887 31378
rect 13769 31306 13887 31311
rect 13769 31243 13809 31306
rect 13843 31243 13887 31306
rect 13769 31234 13887 31243
rect 13769 31175 13809 31234
rect 13843 31175 13887 31234
rect 13769 31162 13887 31175
rect 13769 31107 13809 31162
rect 13843 31107 13887 31162
rect 13769 31090 13887 31107
rect 13769 31039 13809 31090
rect 13843 31039 13887 31090
rect 13769 31018 13887 31039
rect 13769 30971 13809 31018
rect 13843 30971 13887 31018
rect 13769 30946 13887 30971
rect 13769 30903 13809 30946
rect 13843 30903 13887 30946
rect 13769 30874 13887 30903
rect 13769 30835 13809 30874
rect 13843 30835 13887 30874
rect 13769 30802 13887 30835
rect 13769 30767 13809 30802
rect 13843 30767 13887 30802
rect 13769 30733 13887 30767
rect 13769 30696 13809 30733
rect 13843 30696 13887 30733
rect 13769 30665 13887 30696
rect 13769 30624 13809 30665
rect 13843 30624 13887 30665
rect 13769 30597 13887 30624
rect 13769 30552 13809 30597
rect 13843 30552 13887 30597
rect 13769 30529 13887 30552
rect 13769 30480 13809 30529
rect 13843 30480 13887 30529
rect 13769 30461 13887 30480
rect 13769 30408 13809 30461
rect 13843 30408 13887 30461
rect 13769 30393 13887 30408
rect 13769 30336 13809 30393
rect 13843 30336 13887 30393
rect 13769 30325 13887 30336
rect 13769 30264 13809 30325
rect 13843 30264 13887 30325
rect 13769 30257 13887 30264
rect 13769 30192 13809 30257
rect 13843 30192 13887 30257
rect 13769 30189 13887 30192
rect 13769 30155 13809 30189
rect 13843 30155 13887 30189
rect 13769 30154 13887 30155
rect 13769 30087 13809 30154
rect 13843 30087 13887 30154
rect 13769 30082 13887 30087
rect 13769 30019 13809 30082
rect 13843 30019 13887 30082
rect 13769 30010 13887 30019
rect 13769 29951 13809 30010
rect 13843 29951 13887 30010
rect 13769 29938 13887 29951
rect 13769 29883 13809 29938
rect 13843 29883 13887 29938
rect 13769 29866 13887 29883
rect 13769 29815 13809 29866
rect 13843 29815 13887 29866
rect 13769 29794 13887 29815
rect 13769 29747 13809 29794
rect 13843 29747 13887 29794
rect 13769 29722 13887 29747
rect 13769 29679 13809 29722
rect 13843 29679 13887 29722
rect 13769 29650 13887 29679
rect 13769 29611 13809 29650
rect 13843 29611 13887 29650
rect 13769 29578 13887 29611
rect 13769 29543 13809 29578
rect 13843 29543 13887 29578
rect 13769 29509 13887 29543
rect 13769 29472 13809 29509
rect 13843 29472 13887 29509
rect 13769 29441 13887 29472
rect 13769 29400 13809 29441
rect 13843 29400 13887 29441
rect 13769 29373 13887 29400
rect 13769 29328 13809 29373
rect 13843 29328 13887 29373
rect 13769 29305 13887 29328
rect 13769 29256 13809 29305
rect 13843 29256 13887 29305
rect 13769 29237 13887 29256
rect 13769 29184 13809 29237
rect 13843 29184 13887 29237
rect 13769 29169 13887 29184
rect 13769 29112 13809 29169
rect 13843 29112 13887 29169
rect 13769 29101 13887 29112
rect 13769 29040 13809 29101
rect 13843 29040 13887 29101
rect 13769 29033 13887 29040
rect 13769 28968 13809 29033
rect 13843 28968 13887 29033
rect 13769 28965 13887 28968
rect 13769 28931 13809 28965
rect 13843 28931 13887 28965
rect 13769 28930 13887 28931
rect 1119 28850 1237 28868
rect 1119 28800 1161 28850
rect 1195 28800 1237 28850
rect 1119 28778 1237 28800
rect 1119 28732 1161 28778
rect 1195 28732 1237 28778
rect 1119 28706 1237 28732
rect 1119 28664 1161 28706
rect 1195 28664 1237 28706
rect 1119 28634 1237 28664
rect 1119 28596 1161 28634
rect 1195 28596 1237 28634
rect 1119 28562 1237 28596
rect 1119 28528 1161 28562
rect 1195 28528 1237 28562
rect 1119 28494 1237 28528
rect 1119 28456 1161 28494
rect 1195 28456 1237 28494
rect 1119 28426 1237 28456
rect 1119 28384 1161 28426
rect 1195 28384 1237 28426
rect 1119 28358 1237 28384
rect 1119 28312 1161 28358
rect 1195 28312 1237 28358
rect 1119 28290 1237 28312
rect 1119 28240 1161 28290
rect 1195 28240 1237 28290
rect 1119 28222 1237 28240
rect 1119 28168 1161 28222
rect 1195 28168 1237 28222
rect 1119 28154 1237 28168
rect 1119 28096 1161 28154
rect 1195 28096 1237 28154
rect 1119 28086 1237 28096
rect 1119 28024 1161 28086
rect 1195 28024 1237 28086
rect 1119 28018 1237 28024
rect 1119 27952 1161 28018
rect 1195 27952 1237 28018
rect 1119 27950 1237 27952
rect 1119 27916 1161 27950
rect 1195 27916 1237 27950
rect 1119 27914 1237 27916
rect 1119 27848 1161 27914
rect 1195 27848 1237 27914
rect 1119 27842 1237 27848
rect 1119 27780 1161 27842
rect 1195 27780 1237 27842
rect 1119 27770 1237 27780
rect 1119 27712 1161 27770
rect 1195 27712 1237 27770
rect 1119 27698 1237 27712
rect 1119 27644 1161 27698
rect 1195 27644 1237 27698
rect 1119 27626 1237 27644
rect 1119 27576 1161 27626
rect 1195 27576 1237 27626
rect 1119 27554 1237 27576
rect 1119 27508 1161 27554
rect 1195 27508 1237 27554
rect 1119 27482 1237 27508
rect 1119 27440 1161 27482
rect 1195 27440 1237 27482
rect 1119 27410 1237 27440
rect 1119 27372 1161 27410
rect 1195 27372 1237 27410
rect 1119 27338 1237 27372
rect 1119 27304 1161 27338
rect 1195 27304 1237 27338
rect 1119 27270 1237 27304
rect 1119 27232 1161 27270
rect 1195 27232 1237 27270
rect 1119 27202 1237 27232
rect 1119 27160 1161 27202
rect 1195 27160 1237 27202
rect 1119 27134 1237 27160
rect 1119 27088 1161 27134
rect 1195 27088 1237 27134
rect 1119 27066 1237 27088
rect 1119 27016 1161 27066
rect 1195 27016 1237 27066
rect 1659 28879 13357 28909
rect 1659 28875 2119 28879
rect 12897 28875 13357 28879
rect 1659 28553 1982 28875
rect 13032 28553 13357 28875
rect 1659 28505 2119 28553
rect 12897 28505 13357 28553
rect 1659 28489 13357 28505
rect 1659 28422 1726 28489
rect 1976 28482 13357 28489
rect 1976 28475 13031 28482
rect 1976 28422 2093 28475
rect 1659 27504 1689 28422
rect 2063 27504 2093 28422
rect 12923 28422 13031 28475
rect 13281 28422 13357 28482
rect 2156 28172 12840 28368
rect 2156 27758 2382 28172
rect 12614 27758 12840 28172
rect 2156 27556 12840 27758
rect 1659 27447 1726 27504
rect 1976 27451 2093 27504
rect 12923 27504 12953 28422
rect 13327 27504 13357 28422
rect 12923 27451 13031 27504
rect 1976 27447 13031 27451
rect 1659 27440 13031 27447
rect 13281 27440 13357 27504
rect 1659 27421 13357 27440
rect 1659 27334 2119 27421
rect 12897 27334 13357 27421
rect 1659 27084 1985 27334
rect 13035 27084 13357 27334
rect 1659 27047 2119 27084
rect 12897 27047 13357 27084
rect 1659 27017 13357 27047
rect 13769 28863 13809 28930
rect 13843 28863 13887 28930
rect 13769 28858 13887 28863
rect 13769 28795 13809 28858
rect 13843 28795 13887 28858
rect 13769 28786 13887 28795
rect 13769 28727 13809 28786
rect 13843 28727 13887 28786
rect 13769 28693 13887 28727
rect 13769 28659 13809 28693
rect 13843 28659 13887 28693
rect 13769 28625 13887 28659
rect 13769 28591 13809 28625
rect 13843 28591 13887 28625
rect 13769 28557 13887 28591
rect 13769 28523 13809 28557
rect 13843 28523 13887 28557
rect 13769 28489 13887 28523
rect 13769 28455 13809 28489
rect 13843 28455 13887 28489
rect 13769 28421 13887 28455
rect 13769 28387 13809 28421
rect 13843 28387 13887 28421
rect 13769 28353 13887 28387
rect 13769 28319 13809 28353
rect 13843 28319 13887 28353
rect 13769 28285 13887 28319
rect 13769 28251 13809 28285
rect 13843 28251 13887 28285
rect 13769 28217 13887 28251
rect 13769 28183 13809 28217
rect 13843 28183 13887 28217
rect 13769 28149 13887 28183
rect 13769 28115 13809 28149
rect 13843 28115 13887 28149
rect 13769 28081 13887 28115
rect 13769 28047 13809 28081
rect 13843 28047 13887 28081
rect 13769 28013 13887 28047
rect 13769 27979 13809 28013
rect 13843 27979 13887 28013
rect 13769 27945 13887 27979
rect 13769 27911 13809 27945
rect 13843 27911 13887 27945
rect 13769 27877 13887 27911
rect 13769 27843 13809 27877
rect 13843 27843 13887 27877
rect 13769 27809 13887 27843
rect 13769 27775 13809 27809
rect 13843 27775 13887 27809
rect 13769 27741 13887 27775
rect 13769 27707 13809 27741
rect 13843 27707 13887 27741
rect 13769 27673 13887 27707
rect 13769 27639 13809 27673
rect 13843 27639 13887 27673
rect 13769 27605 13887 27639
rect 13769 27571 13809 27605
rect 13843 27571 13887 27605
rect 13769 27537 13887 27571
rect 13769 27503 13809 27537
rect 13843 27503 13887 27537
rect 13769 27469 13887 27503
rect 13769 27435 13809 27469
rect 13843 27435 13887 27469
rect 13769 27401 13887 27435
rect 13769 27367 13809 27401
rect 13843 27367 13887 27401
rect 13769 27333 13887 27367
rect 13769 27299 13809 27333
rect 13843 27299 13887 27333
rect 13769 27265 13887 27299
rect 13769 27231 13809 27265
rect 13843 27231 13887 27265
rect 13769 27197 13887 27231
rect 13769 27163 13809 27197
rect 13843 27163 13887 27197
rect 13769 27129 13887 27163
rect 13769 27095 13809 27129
rect 13843 27095 13887 27129
rect 13769 27061 13887 27095
rect 13769 27027 13809 27061
rect 13843 27027 13887 27061
rect 1119 26998 1237 27016
rect 1119 26944 1161 26998
rect 1195 26944 1237 26998
rect 1119 26930 1237 26944
rect 1119 26872 1161 26930
rect 1195 26872 1237 26930
rect 1119 26862 1237 26872
rect 1119 26800 1161 26862
rect 1195 26800 1237 26862
rect 1119 26794 1237 26800
rect 1119 26728 1161 26794
rect 1195 26728 1237 26794
rect 1119 26726 1237 26728
rect 1119 26692 1161 26726
rect 1195 26692 1237 26726
rect 1119 26690 1237 26692
rect 1119 26624 1161 26690
rect 1195 26624 1237 26690
rect 1119 26618 1237 26624
rect 1119 26556 1161 26618
rect 1195 26556 1237 26618
rect 13769 26993 13887 27027
rect 13769 26959 13809 26993
rect 13843 26959 13887 26993
rect 13769 26925 13887 26959
rect 13769 26891 13809 26925
rect 13843 26891 13887 26925
rect 13769 26857 13887 26891
rect 13769 26823 13809 26857
rect 13843 26823 13887 26857
rect 13769 26789 13887 26823
rect 13769 26755 13809 26789
rect 13843 26755 13887 26789
rect 13769 26721 13887 26755
rect 13769 26687 13809 26721
rect 13843 26687 13887 26721
rect 13769 26653 13887 26687
rect 13769 26619 13809 26653
rect 13843 26619 13887 26653
rect 13769 26613 13887 26619
rect 1119 26546 1237 26556
rect 1119 26488 1161 26546
rect 1195 26488 1237 26546
rect 1119 26474 1237 26488
rect 1119 26420 1161 26474
rect 1195 26420 1237 26474
rect 1119 26402 1237 26420
rect 1119 26352 1161 26402
rect 1195 26352 1237 26402
rect 1119 26330 1237 26352
rect 1119 26284 1161 26330
rect 1195 26284 1237 26330
rect 1119 26258 1237 26284
rect 1119 26216 1161 26258
rect 1195 26216 1237 26258
rect 1119 26186 1237 26216
rect 1119 26148 1161 26186
rect 1195 26148 1237 26186
rect 1119 26114 1237 26148
rect 1119 26080 1161 26114
rect 1195 26080 1237 26114
rect 1119 26046 1237 26080
rect 1119 26008 1161 26046
rect 1195 26008 1237 26046
rect 1119 25978 1237 26008
rect 1119 25936 1161 25978
rect 1195 25936 1237 25978
rect 1119 25910 1237 25936
rect 1119 25864 1161 25910
rect 1195 25864 1237 25910
rect 1119 25842 1237 25864
rect 1119 25792 1161 25842
rect 1195 25792 1237 25842
rect 1119 25774 1237 25792
rect 1119 25720 1161 25774
rect 1195 25720 1237 25774
rect 1119 25706 1237 25720
rect 1119 25648 1161 25706
rect 1195 25648 1237 25706
rect 1119 25638 1237 25648
rect 1119 25576 1161 25638
rect 1195 25576 1237 25638
rect 1119 25570 1237 25576
rect 1119 25504 1161 25570
rect 1195 25504 1237 25570
rect 1119 25502 1237 25504
rect 1119 25468 1161 25502
rect 1195 25468 1237 25502
rect 1119 25466 1237 25468
rect 1119 25400 1161 25466
rect 1195 25400 1237 25466
rect 1119 25394 1237 25400
rect 1119 25332 1161 25394
rect 1195 25332 1237 25394
rect 1119 25322 1237 25332
rect 1119 25264 1161 25322
rect 1195 25264 1237 25322
rect 1119 25250 1237 25264
rect 1119 25196 1161 25250
rect 1195 25196 1237 25250
rect 1119 25178 1237 25196
rect 1119 25128 1161 25178
rect 1195 25128 1237 25178
rect 1119 25106 1237 25128
rect 1119 25060 1161 25106
rect 1195 25060 1237 25106
rect 1119 25034 1237 25060
rect 1119 24992 1161 25034
rect 1195 24992 1237 25034
rect 1119 24962 1237 24992
rect 1119 24924 1161 24962
rect 1195 24924 1237 24962
rect 1119 24890 1237 24924
rect 1119 24856 1161 24890
rect 1195 24856 1237 24890
rect 1119 24822 1237 24856
rect 1119 24784 1161 24822
rect 1195 24784 1237 24822
rect 1119 24754 1237 24784
rect 1698 26585 13887 26613
rect 1698 26551 13809 26585
rect 13843 26551 13887 26585
rect 1698 26517 13887 26551
rect 1698 26483 13809 26517
rect 13843 26483 13887 26517
rect 1698 26449 13887 26483
rect 1698 26415 13809 26449
rect 13843 26415 13887 26449
rect 1698 26381 13887 26415
rect 1698 26347 13809 26381
rect 13843 26347 13887 26381
rect 1698 26313 13887 26347
rect 1698 26279 13809 26313
rect 13843 26279 13887 26313
rect 1698 26245 13887 26279
rect 1698 26211 13809 26245
rect 13843 26211 13887 26245
rect 1698 26177 13887 26211
rect 1698 26143 13809 26177
rect 13843 26143 13887 26177
rect 1698 26109 13887 26143
rect 1698 26080 13809 26109
rect 1698 25313 2270 26080
rect 12712 26075 13809 26080
rect 13843 26075 13887 26109
rect 12712 26041 13887 26075
rect 12712 26007 13809 26041
rect 13843 26007 13887 26041
rect 12712 25973 13887 26007
rect 12712 25939 13809 25973
rect 13843 25939 13887 25973
rect 12712 25905 13887 25939
rect 12712 25871 13809 25905
rect 13843 25871 13887 25905
rect 12712 25837 13887 25871
rect 12712 25803 13809 25837
rect 13843 25803 13887 25837
rect 12712 25769 13887 25803
rect 12712 25735 13809 25769
rect 13843 25735 13887 25769
rect 12712 25701 13887 25735
rect 12712 25667 13809 25701
rect 13843 25667 13887 25701
rect 12712 25633 13887 25667
rect 12712 25599 13809 25633
rect 13843 25599 13887 25633
rect 12712 25565 13887 25599
rect 12712 25531 13809 25565
rect 13843 25531 13887 25565
rect 12712 25497 13887 25531
rect 12712 25463 13809 25497
rect 13843 25463 13887 25497
rect 12712 25429 13887 25463
rect 12712 25395 13809 25429
rect 13843 25395 13887 25429
rect 12712 25361 13887 25395
rect 12712 25327 13809 25361
rect 13843 25327 13887 25361
rect 12712 25313 13887 25327
rect 1698 25293 13887 25313
rect 1698 25259 13809 25293
rect 13843 25259 13887 25293
rect 1698 25225 13887 25259
rect 1698 25191 13809 25225
rect 13843 25191 13887 25225
rect 1698 25157 13887 25191
rect 1698 25123 13809 25157
rect 13843 25123 13887 25157
rect 1698 25089 13887 25123
rect 1698 25055 13809 25089
rect 13843 25055 13887 25089
rect 1698 25021 13887 25055
rect 1698 24987 13809 25021
rect 13843 24987 13887 25021
rect 1698 24953 13887 24987
rect 1698 24919 13809 24953
rect 13843 24919 13887 24953
rect 1698 24885 13887 24919
rect 1698 24851 13809 24885
rect 13843 24851 13887 24885
rect 1698 24817 13887 24851
rect 1698 24783 13809 24817
rect 13843 24783 13887 24817
rect 1698 24780 13887 24783
rect 1119 24712 1161 24754
rect 1195 24712 1237 24754
rect 1119 24686 1237 24712
rect 1119 24640 1161 24686
rect 1195 24640 1237 24686
rect 1119 24618 1237 24640
rect 1119 24568 1161 24618
rect 1195 24568 1237 24618
rect 1119 24550 1237 24568
rect 1119 24496 1161 24550
rect 1195 24496 1237 24550
rect 1119 24482 1237 24496
rect 1119 24424 1161 24482
rect 1195 24424 1237 24482
rect 1119 24414 1237 24424
rect 1119 24352 1161 24414
rect 1195 24352 1237 24414
rect 1119 24346 1237 24352
rect 1119 24280 1161 24346
rect 1195 24280 1237 24346
rect 1119 24278 1237 24280
rect 1119 24244 1161 24278
rect 1195 24244 1237 24278
rect 1119 24242 1237 24244
rect 1119 24176 1161 24242
rect 1195 24176 1237 24242
rect 1119 24170 1237 24176
rect 1119 24108 1161 24170
rect 1195 24108 1237 24170
rect 1119 24098 1237 24108
rect 1119 24040 1161 24098
rect 1195 24040 1237 24098
rect 1119 24026 1237 24040
rect 1119 23972 1161 24026
rect 1195 23972 1237 24026
rect 1119 23954 1237 23972
rect 1119 23904 1161 23954
rect 1195 23904 1237 23954
rect 1119 23882 1237 23904
rect 1119 23836 1161 23882
rect 1195 23836 1237 23882
rect 1119 23810 1237 23836
rect 1119 23768 1161 23810
rect 1195 23768 1237 23810
rect 1119 23738 1237 23768
rect 1119 23700 1161 23738
rect 1195 23700 1237 23738
rect 1119 23666 1237 23700
rect 1119 23632 1161 23666
rect 1195 23632 1237 23666
rect 1119 23598 1237 23632
rect 1119 23560 1161 23598
rect 1195 23560 1237 23598
rect 1119 23530 1237 23560
rect 1119 23488 1161 23530
rect 1195 23488 1237 23530
rect 1119 23462 1237 23488
rect 1119 23416 1161 23462
rect 1195 23416 1237 23462
rect 1119 23394 1237 23416
rect 1119 23344 1161 23394
rect 1195 23344 1237 23394
rect 1119 23326 1237 23344
rect 1119 23272 1161 23326
rect 1195 23272 1237 23326
rect 1119 23258 1237 23272
rect 1119 23200 1161 23258
rect 1195 23200 1237 23258
rect 1119 23190 1237 23200
rect 1119 23128 1161 23190
rect 1195 23128 1237 23190
rect 1119 23122 1237 23128
rect 1119 23056 1161 23122
rect 1195 23056 1237 23122
rect 1119 23054 1237 23056
rect 1119 23020 1161 23054
rect 1195 23020 1237 23054
rect 1119 23018 1237 23020
rect 1119 22952 1161 23018
rect 1195 22952 1237 23018
rect 1119 22946 1237 22952
rect 1119 22884 1161 22946
rect 1195 22884 1237 22946
rect 1119 22874 1237 22884
rect 1119 22816 1161 22874
rect 1195 22816 1237 22874
rect 1119 22802 1237 22816
rect 1119 22748 1161 22802
rect 1195 22748 1237 22802
rect 1119 22730 1237 22748
rect 1119 22680 1161 22730
rect 1195 22680 1237 22730
rect 1119 22658 1237 22680
rect 1119 22612 1161 22658
rect 1195 22612 1237 22658
rect 1119 22586 1237 22612
rect 1119 22544 1161 22586
rect 1195 22544 1237 22586
rect 1119 22514 1237 22544
rect 1119 22476 1161 22514
rect 1195 22476 1237 22514
rect 1119 22442 1237 22476
rect 1119 22408 1161 22442
rect 1195 22408 1237 22442
rect 1119 22374 1237 22408
rect 1119 22336 1161 22374
rect 1195 22336 1237 22374
rect 1119 22306 1237 22336
rect 1119 22264 1161 22306
rect 1195 22264 1237 22306
rect 1119 22238 1237 22264
rect 1119 22192 1161 22238
rect 1195 22192 1237 22238
rect 1119 22170 1237 22192
rect 1119 22120 1161 22170
rect 1195 22120 1237 22170
rect 1119 22102 1237 22120
rect 1119 22048 1161 22102
rect 1195 22048 1237 22102
rect 1119 22034 1237 22048
rect 1119 21976 1161 22034
rect 1195 21976 1237 22034
rect 1119 21966 1237 21976
rect 1119 21904 1161 21966
rect 1195 21904 1237 21966
rect 1119 21898 1237 21904
rect 1119 21832 1161 21898
rect 1195 21832 1237 21898
rect 1119 21830 1237 21832
rect 1119 21796 1161 21830
rect 1195 21796 1237 21830
rect 1119 21794 1237 21796
rect 1119 21728 1161 21794
rect 1195 21728 1237 21794
rect 1119 21722 1237 21728
rect 1119 21660 1161 21722
rect 1195 21660 1237 21722
rect 1119 21650 1237 21660
rect 1119 21592 1161 21650
rect 1195 21592 1237 21650
rect 1119 21578 1237 21592
rect 1119 21524 1161 21578
rect 1195 21524 1237 21578
rect 1119 21506 1237 21524
rect 1119 21456 1161 21506
rect 1195 21456 1237 21506
rect 1119 21434 1237 21456
rect 1119 21388 1161 21434
rect 1195 21388 1237 21434
rect 1119 21362 1237 21388
rect 1119 21320 1161 21362
rect 1195 21320 1237 21362
rect 1119 21290 1237 21320
rect 1119 21252 1161 21290
rect 1195 21252 1237 21290
rect 1119 21218 1237 21252
rect 1119 21184 1161 21218
rect 1195 21184 1237 21218
rect 1119 21150 1237 21184
rect 1119 21112 1161 21150
rect 1195 21112 1237 21150
rect 1119 21082 1237 21112
rect 1119 21040 1161 21082
rect 1195 21040 1237 21082
rect 1119 21014 1237 21040
rect 1119 20968 1161 21014
rect 1195 20968 1237 21014
rect 1119 20946 1237 20968
rect 1119 20896 1161 20946
rect 1195 20896 1237 20946
rect 1119 20878 1237 20896
rect 1119 20824 1161 20878
rect 1195 20824 1237 20878
rect 1119 20810 1237 20824
rect 1119 20752 1161 20810
rect 1195 20752 1237 20810
rect 1119 20742 1237 20752
rect 1119 20680 1161 20742
rect 1195 20680 1237 20742
rect 1119 20674 1237 20680
rect 1119 20608 1161 20674
rect 1195 20608 1237 20674
rect 1119 20606 1237 20608
rect 1119 20572 1161 20606
rect 1195 20572 1237 20606
rect 1119 20570 1237 20572
rect 1119 20504 1161 20570
rect 1195 20504 1237 20570
rect 1119 20498 1237 20504
rect 1119 20436 1161 20498
rect 1195 20436 1237 20498
rect 1119 20426 1237 20436
rect 1119 20368 1161 20426
rect 1195 20368 1237 20426
rect 1119 20354 1237 20368
rect 1119 20300 1161 20354
rect 1195 20300 1237 20354
rect 1119 20282 1237 20300
rect 1119 20232 1161 20282
rect 1195 20232 1237 20282
rect 1119 20210 1237 20232
rect 1119 20164 1161 20210
rect 1195 20164 1237 20210
rect 1119 20138 1237 20164
rect 1119 20096 1161 20138
rect 1195 20096 1237 20138
rect 1119 20066 1237 20096
rect 1119 20028 1161 20066
rect 1195 20028 1237 20066
rect 1119 19994 1237 20028
rect 1119 19960 1161 19994
rect 1195 19960 1237 19994
rect 1119 19926 1237 19960
rect 1119 19888 1161 19926
rect 1195 19888 1237 19926
rect 1119 19858 1237 19888
rect 1119 19816 1161 19858
rect 1195 19816 1237 19858
rect 1119 19790 1237 19816
rect 1119 19744 1161 19790
rect 1195 19744 1237 19790
rect 1119 19722 1237 19744
rect 1119 19672 1161 19722
rect 1195 19672 1237 19722
rect 1119 19654 1237 19672
rect 1119 19600 1161 19654
rect 1195 19600 1237 19654
rect 1119 19586 1237 19600
rect 1119 19528 1161 19586
rect 1195 19528 1237 19586
rect 1119 19518 1237 19528
rect 1119 19456 1161 19518
rect 1195 19456 1237 19518
rect 1119 19450 1237 19456
rect 1119 19384 1161 19450
rect 1195 19384 1237 19450
rect 1119 19382 1237 19384
rect 1119 19348 1161 19382
rect 1195 19348 1237 19382
rect 1119 19346 1237 19348
rect 1119 19280 1161 19346
rect 1195 19280 1237 19346
rect 1119 19274 1237 19280
rect 1119 19212 1161 19274
rect 1195 19212 1237 19274
rect 1119 19202 1237 19212
rect 1119 19144 1161 19202
rect 1195 19144 1237 19202
rect 1119 19130 1237 19144
rect 1119 19076 1161 19130
rect 1195 19076 1237 19130
rect 1119 19058 1237 19076
rect 1119 19008 1161 19058
rect 1195 19008 1237 19058
rect 1119 18986 1237 19008
rect 1119 18940 1161 18986
rect 1195 18940 1237 18986
rect 1119 18914 1237 18940
rect 1119 18872 1161 18914
rect 1195 18872 1237 18914
rect 1119 18842 1237 18872
rect 1119 18804 1161 18842
rect 1195 18804 1237 18842
rect 1119 18770 1237 18804
rect 1119 18736 1161 18770
rect 1195 18736 1237 18770
rect 1119 18702 1237 18736
rect 1119 18664 1161 18702
rect 1195 18664 1237 18702
rect 1119 18634 1237 18664
rect 1119 18592 1161 18634
rect 1195 18592 1237 18634
rect 1119 18566 1237 18592
rect 1119 18520 1161 18566
rect 1195 18520 1237 18566
rect 1119 18498 1237 18520
rect 1119 18448 1161 18498
rect 1195 18448 1237 18498
rect 1119 18430 1237 18448
rect 1119 18376 1161 18430
rect 1195 18376 1237 18430
rect 1119 18362 1237 18376
rect 1119 18304 1161 18362
rect 1195 18304 1237 18362
rect 1119 18294 1237 18304
rect 1119 18232 1161 18294
rect 1195 18232 1237 18294
rect 1119 18226 1237 18232
rect 1119 18160 1161 18226
rect 1195 18160 1237 18226
rect 1119 18158 1237 18160
rect 1119 18124 1161 18158
rect 1195 18124 1237 18158
rect 1119 18122 1237 18124
rect 1119 18056 1161 18122
rect 1195 18056 1237 18122
rect 1119 18050 1237 18056
rect 1119 17988 1161 18050
rect 1195 17988 1237 18050
rect 1119 17978 1237 17988
rect 1119 17920 1161 17978
rect 1195 17920 1237 17978
rect 1119 17906 1237 17920
rect 1119 17852 1161 17906
rect 1195 17852 1237 17906
rect 1119 17834 1237 17852
rect 1119 17784 1161 17834
rect 1195 17784 1237 17834
rect 1119 17762 1237 17784
rect 1119 17716 1161 17762
rect 1195 17716 1237 17762
rect 1119 17690 1237 17716
rect 1119 17648 1161 17690
rect 1195 17648 1237 17690
rect 1119 17618 1237 17648
rect 1119 17580 1161 17618
rect 1195 17580 1237 17618
rect 1119 17546 1237 17580
rect 1119 17512 1161 17546
rect 1195 17512 1237 17546
rect 1119 17478 1237 17512
rect 1119 17440 1161 17478
rect 1195 17440 1237 17478
rect 1119 17410 1237 17440
rect 1119 17368 1161 17410
rect 1195 17368 1237 17410
rect 1119 17342 1237 17368
rect 1119 17296 1161 17342
rect 1195 17296 1237 17342
rect 1119 17274 1237 17296
rect 1119 17224 1161 17274
rect 1195 17224 1237 17274
rect 1119 17206 1237 17224
rect 1119 17152 1161 17206
rect 1195 17152 1237 17206
rect 1119 17138 1237 17152
rect 1119 17080 1161 17138
rect 1195 17080 1237 17138
rect 1119 17070 1237 17080
rect 1119 17008 1161 17070
rect 1195 17008 1237 17070
rect 1119 17002 1237 17008
rect 1119 16936 1161 17002
rect 1195 16936 1237 17002
rect 1119 16934 1237 16936
rect 1119 16900 1161 16934
rect 1195 16900 1237 16934
rect 1119 16898 1237 16900
rect 1119 16832 1161 16898
rect 1195 16832 1237 16898
rect 1119 16826 1237 16832
rect 1119 16764 1161 16826
rect 1195 16764 1237 16826
rect 1119 16754 1237 16764
rect 1119 16696 1161 16754
rect 1195 16696 1237 16754
rect 1119 16682 1237 16696
rect 1119 16628 1161 16682
rect 1195 16628 1237 16682
rect 1119 16610 1237 16628
rect 1119 16560 1161 16610
rect 1195 16560 1237 16610
rect 1119 16538 1237 16560
rect 1119 16492 1161 16538
rect 1195 16492 1237 16538
rect 1119 16466 1237 16492
rect 1119 16424 1161 16466
rect 1195 16424 1237 16466
rect 1119 16394 1237 16424
rect 1119 16356 1161 16394
rect 1195 16356 1237 16394
rect 1119 16322 1237 16356
rect 1119 16288 1161 16322
rect 1195 16288 1237 16322
rect 1119 16254 1237 16288
rect 1119 16216 1161 16254
rect 1195 16216 1237 16254
rect 1119 16186 1237 16216
rect 1119 16144 1161 16186
rect 1195 16144 1237 16186
rect 1119 16118 1237 16144
rect 1119 16072 1161 16118
rect 1195 16072 1237 16118
rect 1119 16050 1237 16072
rect 1119 16000 1161 16050
rect 1195 16000 1237 16050
rect 1119 15982 1237 16000
rect 1119 15928 1161 15982
rect 1195 15928 1237 15982
rect 1119 15914 1237 15928
rect 1119 15856 1161 15914
rect 1195 15856 1237 15914
rect 1119 15846 1237 15856
rect 1119 15784 1161 15846
rect 1195 15784 1237 15846
rect 1119 15778 1237 15784
rect 1119 15712 1161 15778
rect 1195 15712 1237 15778
rect 1119 15710 1237 15712
rect 1119 15676 1161 15710
rect 1195 15676 1237 15710
rect 1119 15674 1237 15676
rect 1119 15608 1161 15674
rect 1195 15608 1237 15674
rect 1119 15602 1237 15608
rect 1119 15540 1161 15602
rect 1195 15540 1237 15602
rect 1119 15530 1237 15540
rect 1119 15472 1161 15530
rect 1195 15472 1237 15530
rect 1119 15458 1237 15472
rect 1119 15404 1161 15458
rect 1195 15404 1237 15458
rect 1119 15386 1237 15404
rect 1119 15336 1161 15386
rect 1195 15336 1237 15386
rect 1119 15314 1237 15336
rect 1119 15268 1161 15314
rect 1195 15268 1237 15314
rect 1119 15242 1237 15268
rect 1119 15200 1161 15242
rect 1195 15200 1237 15242
rect 1119 15170 1237 15200
rect 1119 15132 1161 15170
rect 1195 15132 1237 15170
rect 1119 15098 1237 15132
rect 1119 15064 1161 15098
rect 1195 15064 1237 15098
rect 1119 15030 1237 15064
rect 1119 14992 1161 15030
rect 1195 14992 1237 15030
rect 1119 14962 1237 14992
rect 1119 14920 1161 14962
rect 1195 14920 1237 14962
rect 1119 14894 1237 14920
rect 1119 14848 1161 14894
rect 1195 14848 1237 14894
rect 1119 14826 1237 14848
rect 1119 14776 1161 14826
rect 1195 14776 1237 14826
rect 1119 14758 1237 14776
rect 1119 14704 1161 14758
rect 1195 14704 1237 14758
rect 1119 14690 1237 14704
rect 1119 14632 1161 14690
rect 1195 14632 1237 14690
rect 1119 14622 1237 14632
rect 1119 14560 1161 14622
rect 1195 14560 1237 14622
rect 1119 14554 1237 14560
rect 1119 14488 1161 14554
rect 1195 14488 1237 14554
rect 1119 14486 1237 14488
rect 1119 14452 1161 14486
rect 1195 14452 1237 14486
rect 1119 14450 1237 14452
rect 1119 14384 1161 14450
rect 1195 14384 1237 14450
rect 1119 14378 1237 14384
rect 1119 14316 1161 14378
rect 1195 14316 1237 14378
rect 1119 14306 1237 14316
rect 1119 14248 1161 14306
rect 1195 14248 1237 14306
rect 1119 14234 1237 14248
rect 1119 14180 1161 14234
rect 1195 14180 1237 14234
rect 1119 14162 1237 14180
rect 1119 14112 1161 14162
rect 1195 14112 1237 14162
rect 1119 14090 1237 14112
rect 1119 14044 1161 14090
rect 1195 14044 1237 14090
rect 1119 14018 1237 14044
rect 1119 13976 1161 14018
rect 1195 13976 1237 14018
rect 1119 13946 1237 13976
rect 1119 13908 1161 13946
rect 1195 13908 1237 13946
rect 1119 13874 1237 13908
rect 1119 13840 1161 13874
rect 1195 13840 1237 13874
rect 1119 13806 1237 13840
rect 1119 13768 1161 13806
rect 1195 13768 1237 13806
rect 1119 13738 1237 13768
rect 1119 13696 1161 13738
rect 1195 13696 1237 13738
rect 1119 13670 1237 13696
rect 1119 13624 1161 13670
rect 1195 13624 1237 13670
rect 1119 13602 1237 13624
rect 1119 13552 1161 13602
rect 1195 13552 1237 13602
rect 1119 13534 1237 13552
rect 1119 13480 1161 13534
rect 1195 13480 1237 13534
rect 1119 13466 1237 13480
rect 1119 13408 1161 13466
rect 1195 13408 1237 13466
rect 1119 13398 1237 13408
rect 1119 13336 1161 13398
rect 1195 13336 1237 13398
rect 1119 13330 1237 13336
rect 1119 13264 1161 13330
rect 1195 13264 1237 13330
rect 1119 13262 1237 13264
rect 1119 13228 1161 13262
rect 1195 13228 1237 13262
rect 1119 13226 1237 13228
rect 1119 13160 1161 13226
rect 1195 13160 1237 13226
rect 1119 13154 1237 13160
rect 1119 13092 1161 13154
rect 1195 13092 1237 13154
rect 1119 13082 1237 13092
rect 1119 13024 1161 13082
rect 1195 13024 1237 13082
rect 1119 13010 1237 13024
rect 1119 12956 1161 13010
rect 1195 12956 1237 13010
rect 1119 12938 1237 12956
rect 1119 12888 1161 12938
rect 1195 12888 1237 12938
rect 1119 12866 1237 12888
rect 1119 12820 1161 12866
rect 1195 12820 1237 12866
rect 1119 12794 1237 12820
rect 1119 12752 1161 12794
rect 1195 12752 1237 12794
rect 1119 12722 1237 12752
rect 1119 12684 1161 12722
rect 1195 12684 1237 12722
rect 1119 12650 1237 12684
rect 1119 12616 1161 12650
rect 1195 12616 1237 12650
rect 1119 12582 1237 12616
rect 1119 12544 1161 12582
rect 1195 12544 1237 12582
rect 1119 12514 1237 12544
rect 1119 12472 1161 12514
rect 1195 12472 1237 12514
rect 1119 12446 1237 12472
rect 1119 12400 1161 12446
rect 1195 12400 1237 12446
rect 1119 12378 1237 12400
rect 1119 12328 1161 12378
rect 1195 12328 1237 12378
rect 1119 12310 1237 12328
rect 1119 12256 1161 12310
rect 1195 12256 1237 12310
rect 1119 12242 1237 12256
rect 1119 12184 1161 12242
rect 1195 12184 1237 12242
rect 1119 12174 1237 12184
rect 1119 12112 1161 12174
rect 1195 12112 1237 12174
rect 1119 12106 1237 12112
rect 1119 12040 1161 12106
rect 1195 12040 1237 12106
rect 1119 12038 1237 12040
rect 1119 12004 1161 12038
rect 1195 12004 1237 12038
rect 1119 12002 1237 12004
rect 1119 11936 1161 12002
rect 1195 11936 1237 12002
rect 1119 11930 1237 11936
rect 1119 11868 1161 11930
rect 1195 11868 1237 11930
rect 1119 11858 1237 11868
rect 1119 11800 1161 11858
rect 1195 11800 1237 11858
rect 1119 11786 1237 11800
rect 1119 11732 1161 11786
rect 1195 11732 1237 11786
rect 1119 11714 1237 11732
rect 1119 11664 1161 11714
rect 1195 11664 1237 11714
rect 1119 11642 1237 11664
rect 1119 11596 1161 11642
rect 1195 11596 1237 11642
rect 1119 11570 1237 11596
rect 1119 11528 1161 11570
rect 1195 11528 1237 11570
rect 1119 11498 1237 11528
rect 1119 11460 1161 11498
rect 1195 11460 1237 11498
rect 1119 11426 1237 11460
rect 1119 11392 1161 11426
rect 1195 11392 1237 11426
rect 1119 11358 1237 11392
rect 1119 11320 1161 11358
rect 1195 11320 1237 11358
rect 1119 11290 1237 11320
rect 1119 11248 1161 11290
rect 1195 11248 1237 11290
rect 1119 11222 1237 11248
rect 1119 11176 1161 11222
rect 1195 11176 1237 11222
rect 1119 11154 1237 11176
rect 1119 11104 1161 11154
rect 1195 11104 1237 11154
rect 1119 11086 1237 11104
rect 1119 11032 1161 11086
rect 1195 11032 1237 11086
rect 1119 11018 1237 11032
rect 1119 10960 1161 11018
rect 1195 10960 1237 11018
rect 1119 10950 1237 10960
rect 1119 10888 1161 10950
rect 1195 10888 1237 10950
rect 1119 10882 1237 10888
rect 1119 10816 1161 10882
rect 1195 10816 1237 10882
rect 1119 10814 1237 10816
rect 1119 10780 1161 10814
rect 1195 10780 1237 10814
rect 1119 10778 1237 10780
rect 1119 10712 1161 10778
rect 1195 10712 1237 10778
rect 1119 10706 1237 10712
rect 1119 10644 1161 10706
rect 1195 10644 1237 10706
rect 1119 10634 1237 10644
rect 1119 10576 1161 10634
rect 1195 10576 1237 10634
rect 1119 10562 1237 10576
rect 1119 10508 1161 10562
rect 1195 10508 1237 10562
rect 1119 10490 1237 10508
rect 1119 10440 1161 10490
rect 1195 10440 1237 10490
rect 1119 10418 1237 10440
rect 1119 10372 1161 10418
rect 1195 10372 1237 10418
rect 1119 10319 1237 10372
rect 13769 24749 13887 24780
rect 13769 24715 13809 24749
rect 13843 24715 13887 24749
rect 13769 24681 13887 24715
rect 13769 24647 13809 24681
rect 13843 24647 13887 24681
rect 13769 24613 13887 24647
rect 13769 24579 13809 24613
rect 13843 24579 13887 24613
rect 13769 24545 13887 24579
rect 13769 24511 13809 24545
rect 13843 24511 13887 24545
rect 13769 24477 13887 24511
rect 13769 24443 13809 24477
rect 13843 24443 13887 24477
rect 13769 24409 13887 24443
rect 13769 24375 13809 24409
rect 13843 24375 13887 24409
rect 13769 24341 13887 24375
rect 13769 24307 13809 24341
rect 13843 24307 13887 24341
rect 13769 24273 13887 24307
rect 13769 24239 13809 24273
rect 13843 24239 13887 24273
rect 13769 24205 13887 24239
rect 13769 24171 13809 24205
rect 13843 24171 13887 24205
rect 13769 24137 13887 24171
rect 13769 24103 13809 24137
rect 13843 24103 13887 24137
rect 13769 24069 13887 24103
rect 13769 24035 13809 24069
rect 13843 24035 13887 24069
rect 13769 24001 13887 24035
rect 13769 23967 13809 24001
rect 13843 23967 13887 24001
rect 13769 23933 13887 23967
rect 13769 23899 13809 23933
rect 13843 23899 13887 23933
rect 13769 23865 13887 23899
rect 13769 23831 13809 23865
rect 13843 23831 13887 23865
rect 13769 23797 13887 23831
rect 13769 23763 13809 23797
rect 13843 23763 13887 23797
rect 13769 23729 13887 23763
rect 13769 23695 13809 23729
rect 13843 23695 13887 23729
rect 13769 23661 13887 23695
rect 13769 23627 13809 23661
rect 13843 23627 13887 23661
rect 13769 23593 13887 23627
rect 13769 23559 13809 23593
rect 13843 23559 13887 23593
rect 13769 23525 13887 23559
rect 13769 23491 13809 23525
rect 13843 23491 13887 23525
rect 13769 23457 13887 23491
rect 13769 23423 13809 23457
rect 13843 23423 13887 23457
rect 13769 23389 13887 23423
rect 13769 23347 13809 23389
rect 13843 23347 13887 23389
rect 13769 23321 13887 23347
rect 13769 23275 13809 23321
rect 13843 23275 13887 23321
rect 13769 23253 13887 23275
rect 13769 23203 13809 23253
rect 13843 23203 13887 23253
rect 13769 23185 13887 23203
rect 13769 23131 13809 23185
rect 13843 23131 13887 23185
rect 13769 23117 13887 23131
rect 13769 23059 13809 23117
rect 13843 23059 13887 23117
rect 13769 23049 13887 23059
rect 13769 22987 13809 23049
rect 13843 22987 13887 23049
rect 13769 22981 13887 22987
rect 13769 22915 13809 22981
rect 13843 22915 13887 22981
rect 13769 22913 13887 22915
rect 13769 22879 13809 22913
rect 13843 22879 13887 22913
rect 13769 22877 13887 22879
rect 13769 22811 13809 22877
rect 13843 22811 13887 22877
rect 13769 22805 13887 22811
rect 13769 22743 13809 22805
rect 13843 22743 13887 22805
rect 13769 22733 13887 22743
rect 13769 22675 13809 22733
rect 13843 22675 13887 22733
rect 13769 22661 13887 22675
rect 13769 22607 13809 22661
rect 13843 22607 13887 22661
rect 13769 22589 13887 22607
rect 13769 22539 13809 22589
rect 13843 22539 13887 22589
rect 13769 22517 13887 22539
rect 13769 22471 13809 22517
rect 13843 22471 13887 22517
rect 13769 22445 13887 22471
rect 13769 22403 13809 22445
rect 13843 22403 13887 22445
rect 13769 22373 13887 22403
rect 13769 22335 13809 22373
rect 13843 22335 13887 22373
rect 13769 22301 13887 22335
rect 13769 22267 13809 22301
rect 13843 22267 13887 22301
rect 13769 22233 13887 22267
rect 13769 22195 13809 22233
rect 13843 22195 13887 22233
rect 13769 22165 13887 22195
rect 13769 22123 13809 22165
rect 13843 22123 13887 22165
rect 13769 22097 13887 22123
rect 13769 22051 13809 22097
rect 13843 22051 13887 22097
rect 13769 22029 13887 22051
rect 13769 21979 13809 22029
rect 13843 21979 13887 22029
rect 13769 21961 13887 21979
rect 13769 21907 13809 21961
rect 13843 21907 13887 21961
rect 13769 21893 13887 21907
rect 13769 21835 13809 21893
rect 13843 21835 13887 21893
rect 13769 21825 13887 21835
rect 13769 21763 13809 21825
rect 13843 21763 13887 21825
rect 13769 21757 13887 21763
rect 13769 21691 13809 21757
rect 13843 21691 13887 21757
rect 13769 21689 13887 21691
rect 13769 21655 13809 21689
rect 13843 21655 13887 21689
rect 13769 21653 13887 21655
rect 13769 21587 13809 21653
rect 13843 21587 13887 21653
rect 13769 21581 13887 21587
rect 13769 21519 13809 21581
rect 13843 21519 13887 21581
rect 13769 21509 13887 21519
rect 13769 21451 13809 21509
rect 13843 21451 13887 21509
rect 13769 21437 13887 21451
rect 13769 21383 13809 21437
rect 13843 21383 13887 21437
rect 13769 21365 13887 21383
rect 13769 21315 13809 21365
rect 13843 21315 13887 21365
rect 13769 21293 13887 21315
rect 13769 21247 13809 21293
rect 13843 21247 13887 21293
rect 13769 21221 13887 21247
rect 13769 21179 13809 21221
rect 13843 21179 13887 21221
rect 13769 21149 13887 21179
rect 13769 21111 13809 21149
rect 13843 21111 13887 21149
rect 13769 21077 13887 21111
rect 13769 21043 13809 21077
rect 13843 21043 13887 21077
rect 13769 21009 13887 21043
rect 13769 20971 13809 21009
rect 13843 20971 13887 21009
rect 13769 20941 13887 20971
rect 13769 20899 13809 20941
rect 13843 20899 13887 20941
rect 13769 20873 13887 20899
rect 13769 20827 13809 20873
rect 13843 20827 13887 20873
rect 13769 20805 13887 20827
rect 13769 20755 13809 20805
rect 13843 20755 13887 20805
rect 13769 20737 13887 20755
rect 13769 20683 13809 20737
rect 13843 20683 13887 20737
rect 13769 20669 13887 20683
rect 13769 20611 13809 20669
rect 13843 20611 13887 20669
rect 13769 20601 13887 20611
rect 13769 20539 13809 20601
rect 13843 20539 13887 20601
rect 13769 20533 13887 20539
rect 13769 20467 13809 20533
rect 13843 20467 13887 20533
rect 13769 20465 13887 20467
rect 13769 20431 13809 20465
rect 13843 20431 13887 20465
rect 13769 20429 13887 20431
rect 13769 20363 13809 20429
rect 13843 20363 13887 20429
rect 13769 20357 13887 20363
rect 13769 20295 13809 20357
rect 13843 20295 13887 20357
rect 13769 20285 13887 20295
rect 13769 20227 13809 20285
rect 13843 20227 13887 20285
rect 13769 20213 13887 20227
rect 13769 20159 13809 20213
rect 13843 20159 13887 20213
rect 13769 20141 13887 20159
rect 13769 20091 13809 20141
rect 13843 20091 13887 20141
rect 13769 20069 13887 20091
rect 13769 20023 13809 20069
rect 13843 20023 13887 20069
rect 13769 19997 13887 20023
rect 13769 19955 13809 19997
rect 13843 19955 13887 19997
rect 13769 19925 13887 19955
rect 13769 19887 13809 19925
rect 13843 19887 13887 19925
rect 13769 19853 13887 19887
rect 13769 19819 13809 19853
rect 13843 19819 13887 19853
rect 13769 19785 13887 19819
rect 13769 19747 13809 19785
rect 13843 19747 13887 19785
rect 13769 19717 13887 19747
rect 13769 19675 13809 19717
rect 13843 19675 13887 19717
rect 13769 19649 13887 19675
rect 13769 19603 13809 19649
rect 13843 19603 13887 19649
rect 13769 19581 13887 19603
rect 13769 19531 13809 19581
rect 13843 19531 13887 19581
rect 13769 19513 13887 19531
rect 13769 19459 13809 19513
rect 13843 19459 13887 19513
rect 13769 19445 13887 19459
rect 13769 19387 13809 19445
rect 13843 19387 13887 19445
rect 13769 19377 13887 19387
rect 13769 19315 13809 19377
rect 13843 19315 13887 19377
rect 13769 19309 13887 19315
rect 13769 19243 13809 19309
rect 13843 19243 13887 19309
rect 13769 19241 13887 19243
rect 13769 19207 13809 19241
rect 13843 19207 13887 19241
rect 13769 19205 13887 19207
rect 13769 19139 13809 19205
rect 13843 19139 13887 19205
rect 13769 19133 13887 19139
rect 13769 19071 13809 19133
rect 13843 19071 13887 19133
rect 13769 19061 13887 19071
rect 13769 19003 13809 19061
rect 13843 19003 13887 19061
rect 13769 18989 13887 19003
rect 13769 18935 13809 18989
rect 13843 18935 13887 18989
rect 13769 18917 13887 18935
rect 13769 18867 13809 18917
rect 13843 18867 13887 18917
rect 13769 18845 13887 18867
rect 13769 18799 13809 18845
rect 13843 18799 13887 18845
rect 13769 18773 13887 18799
rect 13769 18731 13809 18773
rect 13843 18731 13887 18773
rect 13769 18701 13887 18731
rect 13769 18663 13809 18701
rect 13843 18663 13887 18701
rect 13769 18629 13887 18663
rect 13769 18595 13809 18629
rect 13843 18595 13887 18629
rect 13769 18561 13887 18595
rect 13769 18523 13809 18561
rect 13843 18523 13887 18561
rect 13769 18493 13887 18523
rect 13769 18451 13809 18493
rect 13843 18451 13887 18493
rect 13769 18425 13887 18451
rect 13769 18379 13809 18425
rect 13843 18379 13887 18425
rect 13769 18357 13887 18379
rect 13769 18307 13809 18357
rect 13843 18307 13887 18357
rect 13769 18289 13887 18307
rect 13769 18235 13809 18289
rect 13843 18235 13887 18289
rect 13769 18221 13887 18235
rect 13769 18163 13809 18221
rect 13843 18163 13887 18221
rect 13769 18153 13887 18163
rect 13769 18091 13809 18153
rect 13843 18091 13887 18153
rect 13769 18085 13887 18091
rect 13769 18019 13809 18085
rect 13843 18019 13887 18085
rect 13769 18017 13887 18019
rect 13769 17983 13809 18017
rect 13843 17983 13887 18017
rect 13769 17981 13887 17983
rect 13769 17915 13809 17981
rect 13843 17915 13887 17981
rect 13769 17909 13887 17915
rect 13769 17847 13809 17909
rect 13843 17847 13887 17909
rect 13769 17837 13887 17847
rect 13769 17779 13809 17837
rect 13843 17779 13887 17837
rect 13769 17765 13887 17779
rect 13769 17711 13809 17765
rect 13843 17711 13887 17765
rect 13769 17693 13887 17711
rect 13769 17643 13809 17693
rect 13843 17643 13887 17693
rect 13769 17621 13887 17643
rect 13769 17575 13809 17621
rect 13843 17575 13887 17621
rect 13769 17549 13887 17575
rect 13769 17507 13809 17549
rect 13843 17507 13887 17549
rect 13769 17477 13887 17507
rect 13769 17439 13809 17477
rect 13843 17439 13887 17477
rect 13769 17405 13887 17439
rect 13769 17371 13809 17405
rect 13843 17371 13887 17405
rect 13769 17337 13887 17371
rect 13769 17299 13809 17337
rect 13843 17299 13887 17337
rect 13769 17269 13887 17299
rect 13769 17227 13809 17269
rect 13843 17227 13887 17269
rect 13769 17201 13887 17227
rect 13769 17155 13809 17201
rect 13843 17155 13887 17201
rect 13769 17133 13887 17155
rect 13769 17083 13809 17133
rect 13843 17083 13887 17133
rect 13769 17065 13887 17083
rect 13769 17011 13809 17065
rect 13843 17011 13887 17065
rect 13769 16997 13887 17011
rect 13769 16939 13809 16997
rect 13843 16939 13887 16997
rect 13769 16929 13887 16939
rect 13769 16867 13809 16929
rect 13843 16867 13887 16929
rect 13769 16861 13887 16867
rect 13769 16795 13809 16861
rect 13843 16795 13887 16861
rect 13769 16793 13887 16795
rect 13769 16759 13809 16793
rect 13843 16759 13887 16793
rect 13769 16757 13887 16759
rect 13769 16691 13809 16757
rect 13843 16691 13887 16757
rect 13769 16685 13887 16691
rect 13769 16623 13809 16685
rect 13843 16623 13887 16685
rect 13769 16613 13887 16623
rect 13769 16555 13809 16613
rect 13843 16555 13887 16613
rect 13769 16541 13887 16555
rect 13769 16487 13809 16541
rect 13843 16487 13887 16541
rect 13769 16469 13887 16487
rect 13769 16419 13809 16469
rect 13843 16419 13887 16469
rect 13769 16397 13887 16419
rect 13769 16351 13809 16397
rect 13843 16351 13887 16397
rect 13769 16325 13887 16351
rect 13769 16283 13809 16325
rect 13843 16283 13887 16325
rect 13769 16253 13887 16283
rect 13769 16215 13809 16253
rect 13843 16215 13887 16253
rect 13769 16181 13887 16215
rect 13769 16147 13809 16181
rect 13843 16147 13887 16181
rect 13769 16113 13887 16147
rect 13769 16075 13809 16113
rect 13843 16075 13887 16113
rect 13769 16045 13887 16075
rect 13769 16003 13809 16045
rect 13843 16003 13887 16045
rect 13769 15977 13887 16003
rect 13769 15931 13809 15977
rect 13843 15931 13887 15977
rect 13769 15909 13887 15931
rect 13769 15859 13809 15909
rect 13843 15859 13887 15909
rect 13769 15841 13887 15859
rect 13769 15787 13809 15841
rect 13843 15787 13887 15841
rect 13769 15773 13887 15787
rect 13769 15715 13809 15773
rect 13843 15715 13887 15773
rect 13769 15705 13887 15715
rect 13769 15643 13809 15705
rect 13843 15643 13887 15705
rect 13769 15637 13887 15643
rect 13769 15571 13809 15637
rect 13843 15571 13887 15637
rect 13769 15569 13887 15571
rect 13769 15535 13809 15569
rect 13843 15535 13887 15569
rect 13769 15533 13887 15535
rect 13769 15467 13809 15533
rect 13843 15467 13887 15533
rect 13769 15461 13887 15467
rect 13769 15399 13809 15461
rect 13843 15399 13887 15461
rect 13769 15389 13887 15399
rect 13769 15331 13809 15389
rect 13843 15331 13887 15389
rect 13769 15317 13887 15331
rect 13769 15263 13809 15317
rect 13843 15263 13887 15317
rect 13769 15245 13887 15263
rect 13769 15195 13809 15245
rect 13843 15195 13887 15245
rect 13769 15173 13887 15195
rect 13769 15127 13809 15173
rect 13843 15127 13887 15173
rect 13769 15101 13887 15127
rect 13769 15059 13809 15101
rect 13843 15059 13887 15101
rect 13769 15029 13887 15059
rect 13769 14991 13809 15029
rect 13843 14991 13887 15029
rect 13769 14957 13887 14991
rect 13769 14923 13809 14957
rect 13843 14923 13887 14957
rect 13769 14889 13887 14923
rect 13769 14851 13809 14889
rect 13843 14851 13887 14889
rect 13769 14821 13887 14851
rect 13769 14779 13809 14821
rect 13843 14779 13887 14821
rect 13769 14753 13887 14779
rect 13769 14707 13809 14753
rect 13843 14707 13887 14753
rect 13769 14685 13887 14707
rect 13769 14635 13809 14685
rect 13843 14635 13887 14685
rect 13769 14617 13887 14635
rect 13769 14563 13809 14617
rect 13843 14563 13887 14617
rect 13769 14549 13887 14563
rect 13769 14491 13809 14549
rect 13843 14491 13887 14549
rect 13769 14481 13887 14491
rect 13769 14419 13809 14481
rect 13843 14419 13887 14481
rect 13769 14413 13887 14419
rect 13769 14347 13809 14413
rect 13843 14347 13887 14413
rect 13769 14345 13887 14347
rect 13769 14311 13809 14345
rect 13843 14311 13887 14345
rect 13769 14309 13887 14311
rect 13769 14243 13809 14309
rect 13843 14243 13887 14309
rect 13769 14237 13887 14243
rect 13769 14175 13809 14237
rect 13843 14175 13887 14237
rect 13769 14165 13887 14175
rect 13769 14107 13809 14165
rect 13843 14107 13887 14165
rect 13769 14093 13887 14107
rect 13769 14039 13809 14093
rect 13843 14039 13887 14093
rect 13769 14021 13887 14039
rect 13769 13971 13809 14021
rect 13843 13971 13887 14021
rect 13769 13949 13887 13971
rect 13769 13903 13809 13949
rect 13843 13903 13887 13949
rect 13769 13877 13887 13903
rect 13769 13835 13809 13877
rect 13843 13835 13887 13877
rect 13769 13805 13887 13835
rect 13769 13767 13809 13805
rect 13843 13767 13887 13805
rect 13769 13733 13887 13767
rect 13769 13699 13809 13733
rect 13843 13699 13887 13733
rect 13769 13665 13887 13699
rect 13769 13627 13809 13665
rect 13843 13627 13887 13665
rect 13769 13597 13887 13627
rect 13769 13555 13809 13597
rect 13843 13555 13887 13597
rect 13769 13529 13887 13555
rect 13769 13483 13809 13529
rect 13843 13483 13887 13529
rect 13769 13461 13887 13483
rect 13769 13411 13809 13461
rect 13843 13411 13887 13461
rect 13769 13393 13887 13411
rect 13769 13339 13809 13393
rect 13843 13339 13887 13393
rect 13769 13325 13887 13339
rect 13769 13267 13809 13325
rect 13843 13267 13887 13325
rect 13769 13257 13887 13267
rect 13769 13195 13809 13257
rect 13843 13195 13887 13257
rect 13769 13189 13887 13195
rect 13769 13123 13809 13189
rect 13843 13123 13887 13189
rect 13769 13121 13887 13123
rect 13769 13087 13809 13121
rect 13843 13087 13887 13121
rect 13769 13085 13887 13087
rect 13769 13019 13809 13085
rect 13843 13019 13887 13085
rect 13769 13013 13887 13019
rect 13769 12951 13809 13013
rect 13843 12951 13887 13013
rect 13769 12941 13887 12951
rect 13769 12883 13809 12941
rect 13843 12883 13887 12941
rect 13769 12869 13887 12883
rect 13769 12815 13809 12869
rect 13843 12815 13887 12869
rect 13769 12797 13887 12815
rect 13769 12747 13809 12797
rect 13843 12747 13887 12797
rect 13769 12725 13887 12747
rect 13769 12679 13809 12725
rect 13843 12679 13887 12725
rect 13769 12653 13887 12679
rect 13769 12611 13809 12653
rect 13843 12611 13887 12653
rect 13769 12581 13887 12611
rect 13769 12543 13809 12581
rect 13843 12543 13887 12581
rect 13769 12509 13887 12543
rect 13769 12475 13809 12509
rect 13843 12475 13887 12509
rect 13769 12441 13887 12475
rect 13769 12403 13809 12441
rect 13843 12403 13887 12441
rect 13769 12373 13887 12403
rect 13769 12331 13809 12373
rect 13843 12331 13887 12373
rect 13769 12305 13887 12331
rect 13769 12259 13809 12305
rect 13843 12259 13887 12305
rect 13769 12237 13887 12259
rect 13769 12187 13809 12237
rect 13843 12187 13887 12237
rect 13769 12169 13887 12187
rect 13769 12115 13809 12169
rect 13843 12115 13887 12169
rect 13769 12101 13887 12115
rect 13769 12043 13809 12101
rect 13843 12043 13887 12101
rect 13769 12033 13887 12043
rect 13769 11971 13809 12033
rect 13843 11971 13887 12033
rect 13769 11965 13887 11971
rect 13769 11899 13809 11965
rect 13843 11899 13887 11965
rect 13769 11897 13887 11899
rect 13769 11863 13809 11897
rect 13843 11863 13887 11897
rect 13769 11861 13887 11863
rect 13769 11795 13809 11861
rect 13843 11795 13887 11861
rect 13769 11789 13887 11795
rect 13769 11727 13809 11789
rect 13843 11727 13887 11789
rect 13769 11717 13887 11727
rect 13769 11659 13809 11717
rect 13843 11659 13887 11717
rect 13769 11645 13887 11659
rect 13769 11591 13809 11645
rect 13843 11591 13887 11645
rect 13769 11573 13887 11591
rect 13769 11523 13809 11573
rect 13843 11523 13887 11573
rect 13769 11501 13887 11523
rect 13769 11455 13809 11501
rect 13843 11455 13887 11501
rect 13769 11429 13887 11455
rect 13769 11387 13809 11429
rect 13843 11387 13887 11429
rect 13769 11357 13887 11387
rect 13769 11319 13809 11357
rect 13843 11319 13887 11357
rect 13769 11285 13887 11319
rect 13769 11251 13809 11285
rect 13843 11251 13887 11285
rect 13769 11217 13887 11251
rect 13769 11179 13809 11217
rect 13843 11179 13887 11217
rect 13769 11149 13887 11179
rect 13769 11107 13809 11149
rect 13843 11107 13887 11149
rect 13769 11081 13887 11107
rect 13769 11035 13809 11081
rect 13843 11035 13887 11081
rect 13769 11013 13887 11035
rect 13769 10963 13809 11013
rect 13843 10963 13887 11013
rect 13769 10945 13887 10963
rect 13769 10891 13809 10945
rect 13843 10891 13887 10945
rect 13769 10877 13887 10891
rect 13769 10819 13809 10877
rect 13843 10819 13887 10877
rect 13769 10809 13887 10819
rect 13769 10747 13809 10809
rect 13843 10747 13887 10809
rect 13769 10741 13887 10747
rect 13769 10675 13809 10741
rect 13843 10675 13887 10741
rect 13769 10673 13887 10675
rect 13769 10639 13809 10673
rect 13843 10639 13887 10673
rect 13769 10637 13887 10639
rect 13769 10571 13809 10637
rect 13843 10571 13887 10637
rect 13769 10565 13887 10571
rect 13769 10503 13809 10565
rect 13843 10503 13887 10565
rect 13769 10493 13887 10503
rect 13769 10435 13809 10493
rect 13843 10435 13887 10493
rect 13769 10421 13887 10435
rect 13769 10367 13809 10421
rect 13843 10367 13887 10421
rect 13769 10319 13887 10367
rect 1119 10278 13887 10319
rect 1119 10244 1298 10278
rect 1336 10244 1370 10278
rect 1404 10244 1438 10278
rect 1476 10244 1506 10278
rect 1548 10244 1574 10278
rect 1620 10244 1642 10278
rect 1692 10244 1710 10278
rect 1764 10244 1778 10278
rect 1836 10244 1846 10278
rect 1908 10244 1914 10278
rect 1980 10244 1982 10278
rect 2016 10244 2018 10278
rect 2084 10244 2090 10278
rect 2152 10244 2162 10278
rect 2220 10244 2234 10278
rect 2288 10244 2306 10278
rect 2356 10244 2378 10278
rect 2424 10244 2450 10278
rect 2492 10244 2522 10278
rect 2560 10244 2594 10278
rect 2628 10244 2662 10278
rect 2700 10244 2730 10278
rect 2772 10244 2798 10278
rect 2844 10244 2866 10278
rect 2916 10244 2934 10278
rect 2988 10244 3002 10278
rect 3060 10244 3070 10278
rect 3132 10244 3138 10278
rect 3204 10244 3206 10278
rect 3240 10244 3242 10278
rect 3308 10244 3314 10278
rect 3376 10244 3386 10278
rect 3444 10244 3458 10278
rect 3512 10244 3530 10278
rect 3580 10244 3602 10278
rect 3648 10244 3674 10278
rect 3716 10244 3746 10278
rect 3784 10244 3818 10278
rect 3852 10244 3886 10278
rect 3924 10244 3954 10278
rect 3996 10244 4022 10278
rect 4068 10244 4090 10278
rect 4140 10244 4158 10278
rect 4212 10244 4226 10278
rect 4284 10244 4294 10278
rect 4356 10244 4362 10278
rect 4428 10244 4430 10278
rect 4464 10244 4466 10278
rect 4532 10244 4538 10278
rect 4600 10244 4610 10278
rect 4668 10244 4682 10278
rect 4736 10244 4754 10278
rect 4804 10244 4826 10278
rect 4872 10244 4898 10278
rect 4940 10244 4970 10278
rect 5008 10244 5042 10278
rect 5076 10244 5110 10278
rect 5148 10244 5178 10278
rect 5220 10244 5246 10278
rect 5292 10244 5314 10278
rect 5364 10244 5382 10278
rect 5436 10244 5450 10278
rect 5508 10244 5518 10278
rect 5580 10244 5586 10278
rect 5652 10244 5654 10278
rect 5688 10244 5690 10278
rect 5756 10244 5762 10278
rect 5824 10244 5834 10278
rect 5892 10244 5906 10278
rect 5960 10244 5978 10278
rect 6028 10244 6050 10278
rect 6096 10244 6122 10278
rect 6164 10244 6194 10278
rect 6232 10244 6266 10278
rect 6300 10244 6334 10278
rect 6372 10244 6402 10278
rect 6444 10244 6470 10278
rect 6516 10244 6538 10278
rect 6588 10244 6606 10278
rect 6660 10244 6674 10278
rect 6732 10244 6742 10278
rect 6804 10244 6810 10278
rect 6876 10244 6878 10278
rect 6912 10244 6914 10278
rect 6980 10244 6986 10278
rect 7048 10244 7058 10278
rect 7116 10244 7130 10278
rect 7184 10244 7202 10278
rect 7252 10244 7274 10278
rect 7320 10244 7346 10278
rect 7388 10244 7418 10278
rect 7456 10244 7490 10278
rect 7524 10244 7558 10278
rect 7596 10244 7626 10278
rect 7668 10244 7694 10278
rect 7740 10244 7762 10278
rect 7812 10244 7830 10278
rect 7884 10244 7898 10278
rect 7956 10244 7966 10278
rect 8028 10244 8034 10278
rect 8100 10244 8102 10278
rect 8136 10244 8138 10278
rect 8204 10244 8210 10278
rect 8272 10244 8282 10278
rect 8340 10244 8354 10278
rect 8408 10244 8426 10278
rect 8476 10244 8498 10278
rect 8544 10244 8570 10278
rect 8612 10244 8642 10278
rect 8680 10244 8714 10278
rect 8748 10244 8782 10278
rect 8820 10244 8850 10278
rect 8892 10244 8918 10278
rect 8964 10244 8986 10278
rect 9036 10244 9054 10278
rect 9108 10244 9122 10278
rect 9180 10244 9190 10278
rect 9252 10244 9258 10278
rect 9324 10244 9326 10278
rect 9360 10244 9362 10278
rect 9428 10244 9434 10278
rect 9496 10244 9506 10278
rect 9564 10244 9578 10278
rect 9632 10244 9650 10278
rect 9700 10244 9722 10278
rect 9768 10244 9794 10278
rect 9836 10244 9866 10278
rect 9904 10244 9938 10278
rect 9972 10244 10006 10278
rect 10044 10244 10074 10278
rect 10116 10244 10142 10278
rect 10188 10244 10210 10278
rect 10260 10244 10278 10278
rect 10332 10244 10346 10278
rect 10404 10244 10414 10278
rect 10476 10244 10482 10278
rect 10548 10244 10550 10278
rect 10584 10244 10586 10278
rect 10652 10244 10658 10278
rect 10720 10244 10730 10278
rect 10788 10244 10802 10278
rect 10856 10244 10874 10278
rect 10924 10244 10946 10278
rect 10992 10244 11018 10278
rect 11060 10244 11090 10278
rect 11128 10244 11162 10278
rect 11196 10244 11230 10278
rect 11268 10244 11298 10278
rect 11340 10244 11366 10278
rect 11412 10244 11434 10278
rect 11484 10244 11502 10278
rect 11556 10244 11570 10278
rect 11628 10244 11638 10278
rect 11700 10244 11706 10278
rect 11772 10244 11774 10278
rect 11808 10244 11810 10278
rect 11876 10244 11882 10278
rect 11944 10244 11954 10278
rect 12012 10244 12026 10278
rect 12080 10244 12098 10278
rect 12148 10244 12170 10278
rect 12216 10244 12242 10278
rect 12284 10244 12314 10278
rect 12352 10244 12386 10278
rect 12420 10244 12454 10278
rect 12492 10244 12522 10278
rect 12564 10244 12590 10278
rect 12636 10244 12658 10278
rect 12708 10244 12726 10278
rect 12780 10244 12794 10278
rect 12852 10244 12862 10278
rect 12924 10244 12930 10278
rect 12996 10244 12998 10278
rect 13032 10244 13034 10278
rect 13100 10244 13106 10278
rect 13168 10244 13178 10278
rect 13236 10244 13250 10278
rect 13304 10244 13322 10278
rect 13372 10244 13394 10278
rect 13440 10244 13466 10278
rect 13508 10244 13538 10278
rect 13576 10244 13610 10278
rect 13644 10244 13678 10278
rect 13716 10244 13887 10278
rect 1119 10201 13887 10244
rect 13968 34691 14122 34725
rect 14156 34706 14297 34725
rect 14331 34706 14361 34740
rect 14156 34691 14361 34706
rect 13968 34672 14361 34691
rect 13968 34653 14297 34672
rect 13968 34619 14122 34653
rect 14156 34638 14297 34653
rect 14331 34638 14361 34672
rect 14156 34619 14361 34638
rect 13968 34604 14361 34619
rect 13968 34581 14297 34604
rect 13968 34547 14122 34581
rect 14156 34570 14297 34581
rect 14331 34570 14361 34604
rect 14156 34547 14361 34570
rect 13968 34536 14361 34547
rect 13968 34509 14297 34536
rect 13968 34475 14122 34509
rect 14156 34502 14297 34509
rect 14331 34502 14361 34536
rect 14156 34475 14361 34502
rect 13968 34468 14361 34475
rect 13968 34437 14297 34468
rect 13968 34403 14122 34437
rect 14156 34434 14297 34437
rect 14331 34434 14361 34468
rect 14156 34403 14361 34434
rect 13968 34400 14361 34403
rect 13968 34366 14297 34400
rect 14331 34366 14361 34400
rect 13968 34365 14361 34366
rect 13968 34331 14122 34365
rect 14156 34332 14361 34365
rect 14156 34331 14297 34332
rect 13968 34298 14297 34331
rect 14331 34298 14361 34332
rect 13968 34293 14361 34298
rect 13968 34259 14122 34293
rect 14156 34264 14361 34293
rect 14156 34259 14297 34264
rect 13968 34230 14297 34259
rect 14331 34230 14361 34264
rect 13968 34221 14361 34230
rect 13968 34187 14122 34221
rect 14156 34196 14361 34221
rect 14156 34187 14297 34196
rect 13968 34162 14297 34187
rect 14331 34162 14361 34196
rect 13968 34149 14361 34162
rect 13968 34115 14122 34149
rect 14156 34128 14361 34149
rect 14156 34115 14297 34128
rect 13968 34094 14297 34115
rect 14331 34094 14361 34128
rect 13968 34077 14361 34094
rect 13968 34043 14122 34077
rect 14156 34060 14361 34077
rect 14156 34043 14297 34060
rect 13968 34026 14297 34043
rect 14331 34026 14361 34060
rect 13968 34005 14361 34026
rect 13968 33971 14122 34005
rect 14156 33992 14361 34005
rect 14156 33971 14297 33992
rect 13968 33958 14297 33971
rect 14331 33958 14361 33992
rect 13968 33933 14361 33958
rect 13968 33899 14122 33933
rect 14156 33924 14361 33933
rect 14156 33899 14297 33924
rect 13968 33890 14297 33899
rect 14331 33890 14361 33924
rect 13968 33861 14361 33890
rect 13968 33827 14122 33861
rect 14156 33856 14361 33861
rect 14156 33827 14297 33856
rect 13968 33822 14297 33827
rect 14331 33822 14361 33856
rect 13968 33789 14361 33822
rect 13968 33755 14122 33789
rect 14156 33788 14361 33789
rect 14156 33755 14297 33788
rect 13968 33754 14297 33755
rect 14331 33754 14361 33788
rect 13968 33720 14361 33754
rect 13968 33717 14297 33720
rect 13968 33683 14122 33717
rect 14156 33686 14297 33717
rect 14331 33686 14361 33720
rect 14156 33683 14361 33686
rect 13968 33652 14361 33683
rect 13968 33645 14297 33652
rect 13968 33611 14122 33645
rect 14156 33618 14297 33645
rect 14331 33618 14361 33652
rect 14156 33611 14361 33618
rect 13968 33584 14361 33611
rect 13968 33573 14297 33584
rect 13968 33539 14122 33573
rect 14156 33550 14297 33573
rect 14331 33550 14361 33584
rect 14156 33539 14361 33550
rect 13968 33516 14361 33539
rect 13968 33501 14297 33516
rect 13968 33467 14122 33501
rect 14156 33482 14297 33501
rect 14331 33482 14361 33516
rect 14156 33467 14361 33482
rect 13968 33448 14361 33467
rect 13968 33429 14297 33448
rect 13968 33395 14122 33429
rect 14156 33414 14297 33429
rect 14331 33414 14361 33448
rect 14156 33395 14361 33414
rect 13968 33380 14361 33395
rect 13968 33357 14297 33380
rect 13968 33323 14122 33357
rect 14156 33346 14297 33357
rect 14331 33346 14361 33380
rect 14156 33323 14361 33346
rect 13968 33312 14361 33323
rect 13968 33285 14297 33312
rect 13968 33251 14122 33285
rect 14156 33278 14297 33285
rect 14331 33278 14361 33312
rect 14156 33251 14361 33278
rect 13968 33244 14361 33251
rect 13968 33213 14297 33244
rect 13968 33179 14122 33213
rect 14156 33210 14297 33213
rect 14331 33210 14361 33244
rect 14156 33179 14361 33210
rect 13968 33176 14361 33179
rect 13968 33142 14297 33176
rect 14331 33142 14361 33176
rect 13968 33141 14361 33142
rect 13968 33107 14122 33141
rect 14156 33108 14361 33141
rect 14156 33107 14297 33108
rect 13968 33074 14297 33107
rect 14331 33074 14361 33108
rect 13968 33069 14361 33074
rect 13968 33035 14122 33069
rect 14156 33040 14361 33069
rect 14156 33035 14297 33040
rect 13968 33006 14297 33035
rect 14331 33006 14361 33040
rect 13968 32997 14361 33006
rect 13968 32963 14122 32997
rect 14156 32972 14361 32997
rect 14156 32963 14297 32972
rect 13968 32938 14297 32963
rect 14331 32938 14361 32972
rect 13968 32925 14361 32938
rect 13968 32891 14122 32925
rect 14156 32904 14361 32925
rect 14156 32891 14297 32904
rect 13968 32870 14297 32891
rect 14331 32870 14361 32904
rect 13968 32853 14361 32870
rect 13968 32819 14122 32853
rect 14156 32836 14361 32853
rect 14156 32819 14297 32836
rect 13968 32802 14297 32819
rect 14331 32802 14361 32836
rect 13968 32781 14361 32802
rect 13968 32747 14122 32781
rect 14156 32768 14361 32781
rect 14156 32747 14297 32768
rect 13968 32734 14297 32747
rect 14331 32734 14361 32768
rect 13968 32709 14361 32734
rect 13968 32675 14122 32709
rect 14156 32700 14361 32709
rect 14156 32675 14297 32700
rect 13968 32666 14297 32675
rect 14331 32666 14361 32700
rect 13968 32637 14361 32666
rect 13968 32603 14122 32637
rect 14156 32632 14361 32637
rect 14156 32603 14297 32632
rect 13968 32598 14297 32603
rect 14331 32598 14361 32632
rect 13968 32565 14361 32598
rect 13968 32531 14122 32565
rect 14156 32564 14361 32565
rect 14156 32531 14297 32564
rect 13968 32530 14297 32531
rect 14331 32530 14361 32564
rect 13968 32496 14361 32530
rect 13968 32493 14297 32496
rect 13968 32459 14122 32493
rect 14156 32462 14297 32493
rect 14331 32462 14361 32496
rect 14156 32459 14361 32462
rect 13968 32428 14361 32459
rect 13968 32421 14297 32428
rect 13968 32387 14122 32421
rect 14156 32394 14297 32421
rect 14331 32394 14361 32428
rect 14156 32387 14361 32394
rect 13968 32360 14361 32387
rect 13968 32349 14297 32360
rect 13968 32315 14122 32349
rect 14156 32326 14297 32349
rect 14331 32326 14361 32360
rect 14156 32315 14361 32326
rect 13968 32292 14361 32315
rect 13968 32277 14297 32292
rect 13968 32243 14122 32277
rect 14156 32258 14297 32277
rect 14331 32258 14361 32292
rect 14156 32243 14361 32258
rect 13968 32224 14361 32243
rect 13968 32205 14297 32224
rect 13968 32171 14122 32205
rect 14156 32190 14297 32205
rect 14331 32190 14361 32224
rect 14156 32171 14361 32190
rect 13968 32156 14361 32171
rect 13968 32133 14297 32156
rect 13968 32099 14122 32133
rect 14156 32122 14297 32133
rect 14331 32122 14361 32156
rect 14156 32099 14361 32122
rect 13968 32088 14361 32099
rect 13968 32061 14297 32088
rect 13968 32027 14122 32061
rect 14156 32054 14297 32061
rect 14331 32054 14361 32088
rect 14156 32027 14361 32054
rect 13968 32020 14361 32027
rect 13968 31989 14297 32020
rect 13968 31955 14122 31989
rect 14156 31986 14297 31989
rect 14331 31986 14361 32020
rect 14156 31955 14361 31986
rect 13968 31952 14361 31955
rect 13968 31918 14297 31952
rect 14331 31918 14361 31952
rect 13968 31917 14361 31918
rect 13968 31883 14122 31917
rect 14156 31884 14361 31917
rect 14156 31883 14297 31884
rect 13968 31850 14297 31883
rect 14331 31850 14361 31884
rect 13968 31845 14361 31850
rect 13968 31811 14122 31845
rect 14156 31816 14361 31845
rect 14156 31811 14297 31816
rect 13968 31782 14297 31811
rect 14331 31782 14361 31816
rect 13968 31773 14361 31782
rect 13968 31739 14122 31773
rect 14156 31748 14361 31773
rect 14156 31739 14297 31748
rect 13968 31714 14297 31739
rect 14331 31714 14361 31748
rect 13968 31701 14361 31714
rect 13968 31667 14122 31701
rect 14156 31680 14361 31701
rect 14156 31667 14297 31680
rect 13968 31646 14297 31667
rect 14331 31646 14361 31680
rect 13968 31629 14361 31646
rect 13968 31595 14122 31629
rect 14156 31612 14361 31629
rect 14156 31595 14297 31612
rect 13968 31578 14297 31595
rect 14331 31578 14361 31612
rect 13968 31557 14361 31578
rect 13968 31523 14122 31557
rect 14156 31544 14361 31557
rect 14156 31523 14297 31544
rect 13968 31510 14297 31523
rect 14331 31510 14361 31544
rect 13968 31485 14361 31510
rect 13968 31451 14122 31485
rect 14156 31476 14361 31485
rect 14156 31451 14297 31476
rect 13968 31442 14297 31451
rect 14331 31442 14361 31476
rect 13968 31413 14361 31442
rect 13968 31379 14122 31413
rect 14156 31408 14361 31413
rect 14156 31379 14297 31408
rect 13968 31374 14297 31379
rect 14331 31374 14361 31408
rect 13968 31341 14361 31374
rect 13968 31307 14122 31341
rect 14156 31340 14361 31341
rect 14156 31307 14297 31340
rect 13968 31306 14297 31307
rect 14331 31306 14361 31340
rect 13968 31272 14361 31306
rect 13968 31269 14297 31272
rect 13968 31235 14122 31269
rect 14156 31238 14297 31269
rect 14331 31238 14361 31272
rect 14156 31235 14361 31238
rect 13968 31204 14361 31235
rect 13968 31197 14297 31204
rect 13968 31163 14122 31197
rect 14156 31170 14297 31197
rect 14331 31170 14361 31204
rect 14156 31163 14361 31170
rect 13968 31136 14361 31163
rect 13968 31125 14297 31136
rect 13968 31091 14122 31125
rect 14156 31102 14297 31125
rect 14331 31102 14361 31136
rect 14156 31091 14361 31102
rect 13968 31068 14361 31091
rect 13968 31053 14297 31068
rect 13968 31019 14122 31053
rect 14156 31034 14297 31053
rect 14331 31034 14361 31068
rect 14156 31019 14361 31034
rect 13968 31000 14361 31019
rect 13968 30981 14297 31000
rect 13968 30947 14122 30981
rect 14156 30966 14297 30981
rect 14331 30966 14361 31000
rect 14156 30947 14361 30966
rect 13968 30932 14361 30947
rect 13968 30909 14297 30932
rect 13968 30875 14122 30909
rect 14156 30898 14297 30909
rect 14331 30898 14361 30932
rect 14156 30875 14361 30898
rect 13968 30864 14361 30875
rect 13968 30837 14297 30864
rect 13968 30803 14122 30837
rect 14156 30830 14297 30837
rect 14331 30830 14361 30864
rect 14156 30803 14361 30830
rect 13968 30796 14361 30803
rect 13968 30765 14297 30796
rect 13968 30731 14122 30765
rect 14156 30762 14297 30765
rect 14331 30762 14361 30796
rect 14156 30731 14361 30762
rect 13968 30728 14361 30731
rect 13968 30694 14297 30728
rect 14331 30694 14361 30728
rect 13968 30693 14361 30694
rect 13968 30659 14122 30693
rect 14156 30660 14361 30693
rect 14156 30659 14297 30660
rect 13968 30626 14297 30659
rect 14331 30626 14361 30660
rect 13968 30621 14361 30626
rect 13968 30587 14122 30621
rect 14156 30592 14361 30621
rect 14156 30587 14297 30592
rect 13968 30558 14297 30587
rect 14331 30558 14361 30592
rect 13968 30549 14361 30558
rect 13968 30515 14122 30549
rect 14156 30524 14361 30549
rect 14156 30515 14297 30524
rect 13968 30490 14297 30515
rect 14331 30490 14361 30524
rect 13968 30477 14361 30490
rect 13968 30443 14122 30477
rect 14156 30456 14361 30477
rect 14156 30443 14297 30456
rect 13968 30422 14297 30443
rect 14331 30422 14361 30456
rect 13968 30405 14361 30422
rect 13968 30371 14122 30405
rect 14156 30388 14361 30405
rect 14156 30371 14297 30388
rect 13968 30354 14297 30371
rect 14331 30354 14361 30388
rect 13968 30333 14361 30354
rect 13968 30299 14122 30333
rect 14156 30320 14361 30333
rect 14156 30299 14297 30320
rect 13968 30286 14297 30299
rect 14331 30286 14361 30320
rect 13968 30261 14361 30286
rect 13968 30227 14122 30261
rect 14156 30252 14361 30261
rect 14156 30227 14297 30252
rect 13968 30218 14297 30227
rect 14331 30218 14361 30252
rect 13968 30189 14361 30218
rect 13968 30155 14122 30189
rect 14156 30184 14361 30189
rect 14156 30155 14297 30184
rect 13968 30150 14297 30155
rect 14331 30150 14361 30184
rect 13968 30117 14361 30150
rect 13968 30083 14122 30117
rect 14156 30116 14361 30117
rect 14156 30083 14297 30116
rect 13968 30082 14297 30083
rect 14331 30082 14361 30116
rect 13968 30048 14361 30082
rect 13968 30045 14297 30048
rect 13968 30011 14122 30045
rect 14156 30014 14297 30045
rect 14331 30014 14361 30048
rect 14156 30011 14361 30014
rect 13968 29980 14361 30011
rect 13968 29973 14297 29980
rect 13968 29939 14122 29973
rect 14156 29946 14297 29973
rect 14331 29946 14361 29980
rect 14156 29939 14361 29946
rect 13968 29912 14361 29939
rect 13968 29901 14297 29912
rect 13968 29867 14122 29901
rect 14156 29878 14297 29901
rect 14331 29878 14361 29912
rect 14156 29867 14361 29878
rect 13968 29844 14361 29867
rect 13968 29829 14297 29844
rect 13968 29795 14122 29829
rect 14156 29810 14297 29829
rect 14331 29810 14361 29844
rect 14156 29795 14361 29810
rect 13968 29776 14361 29795
rect 13968 29757 14297 29776
rect 13968 29723 14122 29757
rect 14156 29742 14297 29757
rect 14331 29742 14361 29776
rect 14156 29723 14361 29742
rect 13968 29708 14361 29723
rect 13968 29685 14297 29708
rect 13968 29651 14122 29685
rect 14156 29674 14297 29685
rect 14331 29674 14361 29708
rect 14156 29651 14361 29674
rect 13968 29640 14361 29651
rect 13968 29613 14297 29640
rect 13968 29579 14122 29613
rect 14156 29606 14297 29613
rect 14331 29606 14361 29640
rect 14156 29579 14361 29606
rect 13968 29572 14361 29579
rect 13968 29541 14297 29572
rect 13968 29507 14122 29541
rect 14156 29538 14297 29541
rect 14331 29538 14361 29572
rect 14156 29507 14361 29538
rect 13968 29504 14361 29507
rect 13968 29470 14297 29504
rect 14331 29470 14361 29504
rect 13968 29469 14361 29470
rect 13968 29435 14122 29469
rect 14156 29436 14361 29469
rect 14156 29435 14297 29436
rect 13968 29402 14297 29435
rect 14331 29402 14361 29436
rect 13968 29397 14361 29402
rect 13968 29363 14122 29397
rect 14156 29368 14361 29397
rect 14156 29363 14297 29368
rect 13968 29334 14297 29363
rect 14331 29334 14361 29368
rect 13968 29325 14361 29334
rect 13968 29291 14122 29325
rect 14156 29300 14361 29325
rect 14156 29291 14297 29300
rect 13968 29266 14297 29291
rect 14331 29266 14361 29300
rect 13968 29253 14361 29266
rect 13968 29219 14122 29253
rect 14156 29232 14361 29253
rect 14156 29219 14297 29232
rect 13968 29198 14297 29219
rect 14331 29198 14361 29232
rect 13968 29181 14361 29198
rect 13968 29147 14122 29181
rect 14156 29164 14361 29181
rect 14156 29147 14297 29164
rect 13968 29130 14297 29147
rect 14331 29130 14361 29164
rect 13968 29109 14361 29130
rect 13968 29075 14122 29109
rect 14156 29096 14361 29109
rect 14156 29075 14297 29096
rect 13968 29062 14297 29075
rect 14331 29062 14361 29096
rect 13968 29037 14361 29062
rect 13968 29003 14122 29037
rect 14156 29028 14361 29037
rect 14156 29003 14297 29028
rect 13968 28994 14297 29003
rect 14331 28994 14361 29028
rect 13968 28965 14361 28994
rect 13968 28931 14122 28965
rect 14156 28960 14361 28965
rect 14156 28931 14297 28960
rect 13968 28926 14297 28931
rect 14331 28926 14361 28960
rect 13968 28893 14361 28926
rect 13968 28859 14122 28893
rect 14156 28892 14361 28893
rect 14156 28859 14297 28892
rect 13968 28858 14297 28859
rect 14331 28858 14361 28892
rect 13968 28824 14361 28858
rect 13968 28821 14297 28824
rect 13968 28787 14122 28821
rect 14156 28790 14297 28821
rect 14331 28790 14361 28824
rect 14156 28787 14361 28790
rect 13968 28756 14361 28787
rect 13968 28749 14297 28756
rect 13968 28715 14122 28749
rect 14156 28722 14297 28749
rect 14331 28722 14361 28756
rect 14156 28715 14361 28722
rect 13968 28688 14361 28715
rect 13968 28677 14297 28688
rect 13968 28643 14122 28677
rect 14156 28654 14297 28677
rect 14331 28654 14361 28688
rect 14156 28643 14361 28654
rect 13968 28620 14361 28643
rect 13968 28605 14297 28620
rect 13968 28571 14122 28605
rect 14156 28586 14297 28605
rect 14331 28586 14361 28620
rect 14156 28571 14361 28586
rect 13968 28552 14361 28571
rect 13968 28533 14297 28552
rect 13968 28499 14122 28533
rect 14156 28518 14297 28533
rect 14331 28518 14361 28552
rect 14156 28499 14361 28518
rect 13968 28484 14361 28499
rect 13968 28461 14297 28484
rect 13968 28427 14122 28461
rect 14156 28450 14297 28461
rect 14331 28450 14361 28484
rect 14156 28427 14361 28450
rect 13968 28416 14361 28427
rect 13968 28389 14297 28416
rect 13968 28355 14122 28389
rect 14156 28382 14297 28389
rect 14331 28382 14361 28416
rect 14156 28355 14361 28382
rect 13968 28348 14361 28355
rect 13968 28317 14297 28348
rect 13968 28283 14122 28317
rect 14156 28314 14297 28317
rect 14331 28314 14361 28348
rect 14156 28283 14361 28314
rect 13968 28280 14361 28283
rect 13968 28246 14297 28280
rect 14331 28246 14361 28280
rect 13968 28245 14361 28246
rect 13968 28211 14122 28245
rect 14156 28212 14361 28245
rect 14156 28211 14297 28212
rect 13968 28178 14297 28211
rect 14331 28178 14361 28212
rect 13968 28173 14361 28178
rect 13968 28139 14122 28173
rect 14156 28144 14361 28173
rect 14156 28139 14297 28144
rect 13968 28110 14297 28139
rect 14331 28110 14361 28144
rect 13968 28101 14361 28110
rect 13968 28067 14122 28101
rect 14156 28076 14361 28101
rect 14156 28067 14297 28076
rect 13968 28042 14297 28067
rect 14331 28042 14361 28076
rect 13968 28029 14361 28042
rect 13968 27995 14122 28029
rect 14156 28008 14361 28029
rect 14156 27995 14297 28008
rect 13968 27974 14297 27995
rect 14331 27974 14361 28008
rect 13968 27957 14361 27974
rect 13968 27923 14122 27957
rect 14156 27940 14361 27957
rect 14156 27923 14297 27940
rect 13968 27906 14297 27923
rect 14331 27906 14361 27940
rect 13968 27885 14361 27906
rect 13968 27851 14122 27885
rect 14156 27872 14361 27885
rect 14156 27851 14297 27872
rect 13968 27838 14297 27851
rect 14331 27838 14361 27872
rect 13968 27813 14361 27838
rect 13968 27779 14122 27813
rect 14156 27804 14361 27813
rect 14156 27779 14297 27804
rect 13968 27770 14297 27779
rect 14331 27770 14361 27804
rect 13968 27741 14361 27770
rect 13968 27707 14122 27741
rect 14156 27736 14361 27741
rect 14156 27707 14297 27736
rect 13968 27702 14297 27707
rect 14331 27702 14361 27736
rect 13968 27669 14361 27702
rect 13968 27635 14122 27669
rect 14156 27668 14361 27669
rect 14156 27635 14297 27668
rect 13968 27634 14297 27635
rect 14331 27634 14361 27668
rect 13968 27600 14361 27634
rect 13968 27597 14297 27600
rect 13968 27563 14122 27597
rect 14156 27566 14297 27597
rect 14331 27566 14361 27600
rect 14156 27563 14361 27566
rect 13968 27532 14361 27563
rect 13968 27525 14297 27532
rect 13968 27491 14122 27525
rect 14156 27498 14297 27525
rect 14331 27498 14361 27532
rect 14156 27491 14361 27498
rect 13968 27464 14361 27491
rect 13968 27453 14297 27464
rect 13968 27419 14122 27453
rect 14156 27430 14297 27453
rect 14331 27430 14361 27464
rect 14156 27419 14361 27430
rect 13968 27396 14361 27419
rect 13968 27381 14297 27396
rect 13968 27347 14122 27381
rect 14156 27362 14297 27381
rect 14331 27362 14361 27396
rect 14156 27347 14361 27362
rect 13968 27328 14361 27347
rect 13968 27309 14297 27328
rect 13968 27275 14122 27309
rect 14156 27294 14297 27309
rect 14331 27294 14361 27328
rect 14156 27275 14361 27294
rect 13968 27260 14361 27275
rect 13968 27237 14297 27260
rect 13968 27203 14122 27237
rect 14156 27226 14297 27237
rect 14331 27226 14361 27260
rect 14156 27203 14361 27226
rect 13968 27192 14361 27203
rect 13968 27165 14297 27192
rect 13968 27131 14122 27165
rect 14156 27158 14297 27165
rect 14331 27158 14361 27192
rect 14156 27131 14361 27158
rect 13968 27124 14361 27131
rect 13968 27093 14297 27124
rect 13968 27059 14122 27093
rect 14156 27090 14297 27093
rect 14331 27090 14361 27124
rect 14156 27059 14361 27090
rect 13968 27056 14361 27059
rect 13968 27022 14297 27056
rect 14331 27022 14361 27056
rect 13968 27021 14361 27022
rect 13968 26987 14122 27021
rect 14156 26988 14361 27021
rect 14156 26987 14297 26988
rect 13968 26954 14297 26987
rect 14331 26954 14361 26988
rect 13968 26949 14361 26954
rect 13968 26915 14122 26949
rect 14156 26920 14361 26949
rect 14156 26915 14297 26920
rect 13968 26886 14297 26915
rect 14331 26886 14361 26920
rect 13968 26877 14361 26886
rect 13968 26843 14122 26877
rect 14156 26852 14361 26877
rect 14156 26843 14297 26852
rect 13968 26818 14297 26843
rect 14331 26818 14361 26852
rect 13968 26805 14361 26818
rect 13968 26771 14122 26805
rect 14156 26784 14361 26805
rect 14156 26771 14297 26784
rect 13968 26750 14297 26771
rect 14331 26750 14361 26784
rect 13968 26733 14361 26750
rect 13968 26699 14122 26733
rect 14156 26716 14361 26733
rect 14156 26699 14297 26716
rect 13968 26682 14297 26699
rect 14331 26682 14361 26716
rect 13968 26661 14361 26682
rect 13968 26627 14122 26661
rect 14156 26648 14361 26661
rect 14156 26627 14297 26648
rect 13968 26614 14297 26627
rect 14331 26614 14361 26648
rect 13968 26589 14361 26614
rect 13968 26555 14122 26589
rect 14156 26580 14361 26589
rect 14156 26555 14297 26580
rect 13968 26546 14297 26555
rect 14331 26546 14361 26580
rect 13968 26517 14361 26546
rect 13968 26483 14122 26517
rect 14156 26512 14361 26517
rect 14156 26483 14297 26512
rect 13968 26478 14297 26483
rect 14331 26478 14361 26512
rect 13968 26445 14361 26478
rect 13968 26411 14122 26445
rect 14156 26444 14361 26445
rect 14156 26411 14297 26444
rect 13968 26410 14297 26411
rect 14331 26410 14361 26444
rect 13968 26376 14361 26410
rect 13968 26373 14297 26376
rect 13968 26339 14122 26373
rect 14156 26342 14297 26373
rect 14331 26342 14361 26376
rect 14156 26339 14361 26342
rect 13968 26308 14361 26339
rect 13968 26301 14297 26308
rect 13968 26267 14122 26301
rect 14156 26274 14297 26301
rect 14331 26274 14361 26308
rect 14156 26267 14361 26274
rect 13968 26240 14361 26267
rect 13968 26229 14297 26240
rect 13968 26195 14122 26229
rect 14156 26206 14297 26229
rect 14331 26206 14361 26240
rect 14156 26195 14361 26206
rect 13968 26172 14361 26195
rect 13968 26157 14297 26172
rect 13968 26123 14122 26157
rect 14156 26138 14297 26157
rect 14331 26138 14361 26172
rect 14156 26123 14361 26138
rect 13968 26104 14361 26123
rect 13968 26085 14297 26104
rect 13968 26051 14122 26085
rect 14156 26070 14297 26085
rect 14331 26070 14361 26104
rect 14156 26051 14361 26070
rect 13968 26036 14361 26051
rect 13968 26013 14297 26036
rect 13968 25979 14122 26013
rect 14156 26002 14297 26013
rect 14331 26002 14361 26036
rect 14156 25979 14361 26002
rect 13968 25968 14361 25979
rect 13968 25941 14297 25968
rect 13968 25907 14122 25941
rect 14156 25934 14297 25941
rect 14331 25934 14361 25968
rect 14156 25907 14361 25934
rect 13968 25900 14361 25907
rect 13968 25869 14297 25900
rect 13968 25835 14122 25869
rect 14156 25866 14297 25869
rect 14331 25866 14361 25900
rect 14156 25835 14361 25866
rect 13968 25832 14361 25835
rect 13968 25798 14297 25832
rect 14331 25798 14361 25832
rect 13968 25797 14361 25798
rect 13968 25763 14122 25797
rect 14156 25764 14361 25797
rect 14156 25763 14297 25764
rect 13968 25730 14297 25763
rect 14331 25730 14361 25764
rect 13968 25725 14361 25730
rect 13968 25691 14122 25725
rect 14156 25696 14361 25725
rect 14156 25691 14297 25696
rect 13968 25662 14297 25691
rect 14331 25662 14361 25696
rect 13968 25653 14361 25662
rect 13968 25619 14122 25653
rect 14156 25628 14361 25653
rect 14156 25619 14297 25628
rect 13968 25594 14297 25619
rect 14331 25594 14361 25628
rect 13968 25581 14361 25594
rect 13968 25547 14122 25581
rect 14156 25560 14361 25581
rect 14156 25547 14297 25560
rect 13968 25526 14297 25547
rect 14331 25526 14361 25560
rect 13968 25509 14361 25526
rect 13968 25475 14122 25509
rect 14156 25492 14361 25509
rect 14156 25475 14297 25492
rect 13968 25458 14297 25475
rect 14331 25458 14361 25492
rect 13968 25437 14361 25458
rect 13968 25403 14122 25437
rect 14156 25424 14361 25437
rect 14156 25403 14297 25424
rect 13968 25390 14297 25403
rect 14331 25390 14361 25424
rect 13968 25365 14361 25390
rect 13968 25331 14122 25365
rect 14156 25356 14361 25365
rect 14156 25331 14297 25356
rect 13968 25322 14297 25331
rect 14331 25322 14361 25356
rect 13968 25293 14361 25322
rect 13968 25259 14122 25293
rect 14156 25288 14361 25293
rect 14156 25259 14297 25288
rect 13968 25254 14297 25259
rect 14331 25254 14361 25288
rect 13968 25221 14361 25254
rect 13968 25187 14122 25221
rect 14156 25220 14361 25221
rect 14156 25187 14297 25220
rect 13968 25186 14297 25187
rect 14331 25186 14361 25220
rect 13968 25152 14361 25186
rect 13968 25149 14297 25152
rect 13968 25115 14122 25149
rect 14156 25118 14297 25149
rect 14331 25118 14361 25152
rect 14156 25115 14361 25118
rect 13968 25084 14361 25115
rect 13968 25077 14297 25084
rect 13968 25043 14122 25077
rect 14156 25050 14297 25077
rect 14331 25050 14361 25084
rect 14156 25043 14361 25050
rect 13968 25016 14361 25043
rect 13968 25005 14297 25016
rect 13968 24971 14122 25005
rect 14156 24982 14297 25005
rect 14331 24982 14361 25016
rect 14156 24971 14361 24982
rect 13968 24948 14361 24971
rect 13968 24933 14297 24948
rect 13968 24899 14122 24933
rect 14156 24914 14297 24933
rect 14331 24914 14361 24948
rect 14156 24899 14361 24914
rect 13968 24880 14361 24899
rect 13968 24861 14297 24880
rect 13968 24827 14122 24861
rect 14156 24846 14297 24861
rect 14331 24846 14361 24880
rect 14156 24827 14361 24846
rect 13968 24812 14361 24827
rect 13968 24789 14297 24812
rect 13968 24755 14122 24789
rect 14156 24778 14297 24789
rect 14331 24778 14361 24812
rect 14156 24755 14361 24778
rect 13968 24744 14361 24755
rect 13968 24717 14297 24744
rect 13968 24683 14122 24717
rect 14156 24710 14297 24717
rect 14331 24710 14361 24744
rect 14156 24683 14361 24710
rect 13968 24676 14361 24683
rect 13968 24645 14297 24676
rect 13968 24611 14122 24645
rect 14156 24642 14297 24645
rect 14331 24642 14361 24676
rect 14156 24611 14361 24642
rect 13968 24608 14361 24611
rect 13968 24574 14297 24608
rect 14331 24574 14361 24608
rect 13968 24573 14361 24574
rect 13968 24539 14122 24573
rect 14156 24540 14361 24573
rect 14156 24539 14297 24540
rect 13968 24506 14297 24539
rect 14331 24506 14361 24540
rect 13968 24501 14361 24506
rect 13968 24467 14122 24501
rect 14156 24472 14361 24501
rect 14156 24467 14297 24472
rect 13968 24438 14297 24467
rect 14331 24438 14361 24472
rect 13968 24429 14361 24438
rect 13968 24395 14122 24429
rect 14156 24404 14361 24429
rect 14156 24395 14297 24404
rect 13968 24370 14297 24395
rect 14331 24370 14361 24404
rect 13968 24357 14361 24370
rect 13968 24323 14122 24357
rect 14156 24336 14361 24357
rect 14156 24323 14297 24336
rect 13968 24302 14297 24323
rect 14331 24302 14361 24336
rect 13968 24285 14361 24302
rect 13968 24251 14122 24285
rect 14156 24268 14361 24285
rect 14156 24251 14297 24268
rect 13968 24234 14297 24251
rect 14331 24234 14361 24268
rect 13968 24213 14361 24234
rect 13968 24179 14122 24213
rect 14156 24200 14361 24213
rect 14156 24179 14297 24200
rect 13968 24166 14297 24179
rect 14331 24166 14361 24200
rect 13968 24141 14361 24166
rect 13968 24107 14122 24141
rect 14156 24132 14361 24141
rect 14156 24107 14297 24132
rect 13968 24098 14297 24107
rect 14331 24098 14361 24132
rect 13968 24069 14361 24098
rect 13968 24035 14122 24069
rect 14156 24064 14361 24069
rect 14156 24035 14297 24064
rect 13968 24030 14297 24035
rect 14331 24030 14361 24064
rect 13968 23997 14361 24030
rect 13968 23963 14122 23997
rect 14156 23996 14361 23997
rect 14156 23963 14297 23996
rect 13968 23962 14297 23963
rect 14331 23962 14361 23996
rect 13968 23928 14361 23962
rect 13968 23925 14297 23928
rect 13968 23891 14122 23925
rect 14156 23894 14297 23925
rect 14331 23894 14361 23928
rect 14156 23891 14361 23894
rect 13968 23860 14361 23891
rect 13968 23853 14297 23860
rect 13968 23819 14122 23853
rect 14156 23826 14297 23853
rect 14331 23826 14361 23860
rect 14156 23819 14361 23826
rect 13968 23792 14361 23819
rect 13968 23781 14297 23792
rect 13968 23747 14122 23781
rect 14156 23758 14297 23781
rect 14331 23758 14361 23792
rect 14156 23747 14361 23758
rect 13968 23724 14361 23747
rect 13968 23709 14297 23724
rect 13968 23675 14122 23709
rect 14156 23690 14297 23709
rect 14331 23690 14361 23724
rect 14156 23675 14361 23690
rect 13968 23656 14361 23675
rect 13968 23637 14297 23656
rect 13968 23603 14122 23637
rect 14156 23622 14297 23637
rect 14331 23622 14361 23656
rect 14156 23603 14361 23622
rect 13968 23588 14361 23603
rect 13968 23565 14297 23588
rect 13968 23531 14122 23565
rect 14156 23554 14297 23565
rect 14331 23554 14361 23588
rect 14156 23531 14361 23554
rect 13968 23520 14361 23531
rect 13968 23493 14297 23520
rect 13968 23459 14122 23493
rect 14156 23486 14297 23493
rect 14331 23486 14361 23520
rect 14156 23459 14361 23486
rect 13968 23452 14361 23459
rect 13968 23421 14297 23452
rect 13968 23387 14122 23421
rect 14156 23418 14297 23421
rect 14331 23418 14361 23452
rect 14156 23387 14361 23418
rect 13968 23384 14361 23387
rect 13968 23350 14297 23384
rect 14331 23350 14361 23384
rect 13968 23349 14361 23350
rect 13968 23315 14122 23349
rect 14156 23316 14361 23349
rect 14156 23315 14297 23316
rect 13968 23282 14297 23315
rect 14331 23282 14361 23316
rect 13968 23277 14361 23282
rect 13968 23243 14122 23277
rect 14156 23248 14361 23277
rect 14156 23243 14297 23248
rect 13968 23214 14297 23243
rect 14331 23214 14361 23248
rect 13968 23205 14361 23214
rect 13968 23171 14122 23205
rect 14156 23180 14361 23205
rect 14156 23171 14297 23180
rect 13968 23146 14297 23171
rect 14331 23146 14361 23180
rect 13968 23133 14361 23146
rect 13968 23099 14122 23133
rect 14156 23112 14361 23133
rect 14156 23099 14297 23112
rect 13968 23078 14297 23099
rect 14331 23078 14361 23112
rect 13968 23061 14361 23078
rect 13968 23027 14122 23061
rect 14156 23044 14361 23061
rect 14156 23027 14297 23044
rect 13968 23010 14297 23027
rect 14331 23010 14361 23044
rect 13968 22989 14361 23010
rect 13968 22955 14122 22989
rect 14156 22976 14361 22989
rect 14156 22955 14297 22976
rect 13968 22942 14297 22955
rect 14331 22942 14361 22976
rect 13968 22917 14361 22942
rect 13968 22883 14122 22917
rect 14156 22908 14361 22917
rect 14156 22883 14297 22908
rect 13968 22874 14297 22883
rect 14331 22874 14361 22908
rect 13968 22845 14361 22874
rect 13968 22811 14122 22845
rect 14156 22840 14361 22845
rect 14156 22811 14297 22840
rect 13968 22806 14297 22811
rect 14331 22806 14361 22840
rect 13968 22773 14361 22806
rect 13968 22739 14122 22773
rect 14156 22772 14361 22773
rect 14156 22739 14297 22772
rect 13968 22738 14297 22739
rect 14331 22738 14361 22772
rect 13968 22704 14361 22738
rect 13968 22701 14297 22704
rect 13968 22667 14122 22701
rect 14156 22670 14297 22701
rect 14331 22670 14361 22704
rect 14156 22667 14361 22670
rect 13968 22636 14361 22667
rect 13968 22629 14297 22636
rect 13968 22595 14122 22629
rect 14156 22602 14297 22629
rect 14331 22602 14361 22636
rect 14156 22595 14361 22602
rect 13968 22568 14361 22595
rect 13968 22557 14297 22568
rect 13968 22523 14122 22557
rect 14156 22534 14297 22557
rect 14331 22534 14361 22568
rect 14156 22523 14361 22534
rect 13968 22500 14361 22523
rect 13968 22485 14297 22500
rect 13968 22451 14122 22485
rect 14156 22466 14297 22485
rect 14331 22466 14361 22500
rect 14156 22451 14361 22466
rect 13968 22432 14361 22451
rect 13968 22413 14297 22432
rect 13968 22379 14122 22413
rect 14156 22398 14297 22413
rect 14331 22398 14361 22432
rect 14156 22379 14361 22398
rect 13968 22364 14361 22379
rect 13968 22341 14297 22364
rect 13968 22307 14122 22341
rect 14156 22330 14297 22341
rect 14331 22330 14361 22364
rect 14156 22307 14361 22330
rect 13968 22296 14361 22307
rect 13968 22269 14297 22296
rect 13968 22235 14122 22269
rect 14156 22262 14297 22269
rect 14331 22262 14361 22296
rect 14156 22235 14361 22262
rect 13968 22228 14361 22235
rect 13968 22197 14297 22228
rect 13968 22163 14122 22197
rect 14156 22194 14297 22197
rect 14331 22194 14361 22228
rect 14156 22163 14361 22194
rect 13968 22160 14361 22163
rect 13968 22126 14297 22160
rect 14331 22126 14361 22160
rect 13968 22125 14361 22126
rect 13968 22091 14122 22125
rect 14156 22092 14361 22125
rect 14156 22091 14297 22092
rect 13968 22058 14297 22091
rect 14331 22058 14361 22092
rect 13968 22053 14361 22058
rect 13968 22019 14122 22053
rect 14156 22024 14361 22053
rect 14156 22019 14297 22024
rect 13968 21990 14297 22019
rect 14331 21990 14361 22024
rect 13968 21981 14361 21990
rect 13968 21947 14122 21981
rect 14156 21956 14361 21981
rect 14156 21947 14297 21956
rect 13968 21922 14297 21947
rect 14331 21922 14361 21956
rect 13968 21909 14361 21922
rect 13968 21875 14122 21909
rect 14156 21888 14361 21909
rect 14156 21875 14297 21888
rect 13968 21854 14297 21875
rect 14331 21854 14361 21888
rect 13968 21837 14361 21854
rect 13968 21803 14122 21837
rect 14156 21820 14361 21837
rect 14156 21803 14297 21820
rect 13968 21786 14297 21803
rect 14331 21786 14361 21820
rect 13968 21765 14361 21786
rect 13968 21731 14122 21765
rect 14156 21752 14361 21765
rect 14156 21731 14297 21752
rect 13968 21718 14297 21731
rect 14331 21718 14361 21752
rect 13968 21693 14361 21718
rect 13968 21659 14122 21693
rect 14156 21684 14361 21693
rect 14156 21659 14297 21684
rect 13968 21650 14297 21659
rect 14331 21650 14361 21684
rect 13968 21621 14361 21650
rect 13968 21587 14122 21621
rect 14156 21616 14361 21621
rect 14156 21587 14297 21616
rect 13968 21582 14297 21587
rect 14331 21582 14361 21616
rect 13968 21549 14361 21582
rect 13968 21515 14122 21549
rect 14156 21548 14361 21549
rect 14156 21515 14297 21548
rect 13968 21514 14297 21515
rect 14331 21514 14361 21548
rect 13968 21480 14361 21514
rect 13968 21477 14297 21480
rect 13968 21443 14122 21477
rect 14156 21446 14297 21477
rect 14331 21446 14361 21480
rect 14156 21443 14361 21446
rect 13968 21412 14361 21443
rect 13968 21405 14297 21412
rect 13968 21371 14122 21405
rect 14156 21378 14297 21405
rect 14331 21378 14361 21412
rect 14156 21371 14361 21378
rect 13968 21344 14361 21371
rect 13968 21333 14297 21344
rect 13968 21299 14122 21333
rect 14156 21310 14297 21333
rect 14331 21310 14361 21344
rect 14156 21299 14361 21310
rect 13968 21276 14361 21299
rect 13968 21261 14297 21276
rect 13968 21227 14122 21261
rect 14156 21242 14297 21261
rect 14331 21242 14361 21276
rect 14156 21227 14361 21242
rect 13968 21208 14361 21227
rect 13968 21189 14297 21208
rect 13968 21155 14122 21189
rect 14156 21174 14297 21189
rect 14331 21174 14361 21208
rect 14156 21155 14361 21174
rect 13968 21140 14361 21155
rect 13968 21117 14297 21140
rect 13968 21083 14122 21117
rect 14156 21106 14297 21117
rect 14331 21106 14361 21140
rect 14156 21083 14361 21106
rect 13968 21072 14361 21083
rect 13968 21045 14297 21072
rect 13968 21011 14122 21045
rect 14156 21038 14297 21045
rect 14331 21038 14361 21072
rect 14156 21011 14361 21038
rect 13968 21004 14361 21011
rect 13968 20973 14297 21004
rect 13968 20939 14122 20973
rect 14156 20970 14297 20973
rect 14331 20970 14361 21004
rect 14156 20939 14361 20970
rect 13968 20936 14361 20939
rect 13968 20902 14297 20936
rect 14331 20902 14361 20936
rect 13968 20901 14361 20902
rect 13968 20867 14122 20901
rect 14156 20868 14361 20901
rect 14156 20867 14297 20868
rect 13968 20834 14297 20867
rect 14331 20834 14361 20868
rect 13968 20829 14361 20834
rect 13968 20795 14122 20829
rect 14156 20800 14361 20829
rect 14156 20795 14297 20800
rect 13968 20766 14297 20795
rect 14331 20766 14361 20800
rect 13968 20757 14361 20766
rect 13968 20723 14122 20757
rect 14156 20732 14361 20757
rect 14156 20723 14297 20732
rect 13968 20698 14297 20723
rect 14331 20698 14361 20732
rect 13968 20685 14361 20698
rect 13968 20651 14122 20685
rect 14156 20664 14361 20685
rect 14156 20651 14297 20664
rect 13968 20630 14297 20651
rect 14331 20630 14361 20664
rect 13968 20613 14361 20630
rect 13968 20579 14122 20613
rect 14156 20596 14361 20613
rect 14156 20579 14297 20596
rect 13968 20562 14297 20579
rect 14331 20562 14361 20596
rect 13968 20541 14361 20562
rect 13968 20507 14122 20541
rect 14156 20528 14361 20541
rect 14156 20507 14297 20528
rect 13968 20494 14297 20507
rect 14331 20494 14361 20528
rect 13968 20469 14361 20494
rect 13968 20435 14122 20469
rect 14156 20460 14361 20469
rect 14156 20435 14297 20460
rect 13968 20426 14297 20435
rect 14331 20426 14361 20460
rect 13968 20397 14361 20426
rect 13968 20363 14122 20397
rect 14156 20392 14361 20397
rect 14156 20363 14297 20392
rect 13968 20358 14297 20363
rect 14331 20358 14361 20392
rect 13968 20325 14361 20358
rect 13968 20291 14122 20325
rect 14156 20324 14361 20325
rect 14156 20291 14297 20324
rect 13968 20290 14297 20291
rect 14331 20290 14361 20324
rect 13968 20256 14361 20290
rect 13968 20253 14297 20256
rect 13968 20219 14122 20253
rect 14156 20222 14297 20253
rect 14331 20222 14361 20256
rect 14156 20219 14361 20222
rect 13968 20188 14361 20219
rect 13968 20181 14297 20188
rect 13968 20147 14122 20181
rect 14156 20154 14297 20181
rect 14331 20154 14361 20188
rect 14156 20147 14361 20154
rect 13968 20120 14361 20147
rect 13968 20109 14297 20120
rect 13968 20075 14122 20109
rect 14156 20086 14297 20109
rect 14331 20086 14361 20120
rect 14156 20075 14361 20086
rect 13968 20052 14361 20075
rect 13968 20037 14297 20052
rect 13968 20003 14122 20037
rect 14156 20018 14297 20037
rect 14331 20018 14361 20052
rect 14156 20003 14361 20018
rect 13968 19984 14361 20003
rect 13968 19965 14297 19984
rect 13968 19931 14122 19965
rect 14156 19950 14297 19965
rect 14331 19950 14361 19984
rect 14156 19931 14361 19950
rect 13968 19916 14361 19931
rect 13968 19893 14297 19916
rect 13968 19859 14122 19893
rect 14156 19882 14297 19893
rect 14331 19882 14361 19916
rect 14156 19859 14361 19882
rect 13968 19848 14361 19859
rect 13968 19821 14297 19848
rect 13968 19787 14122 19821
rect 14156 19814 14297 19821
rect 14331 19814 14361 19848
rect 14156 19787 14361 19814
rect 13968 19780 14361 19787
rect 13968 19749 14297 19780
rect 13968 19715 14122 19749
rect 14156 19746 14297 19749
rect 14331 19746 14361 19780
rect 14156 19715 14361 19746
rect 13968 19712 14361 19715
rect 13968 19678 14297 19712
rect 14331 19678 14361 19712
rect 13968 19677 14361 19678
rect 13968 19643 14122 19677
rect 14156 19644 14361 19677
rect 14156 19643 14297 19644
rect 13968 19610 14297 19643
rect 14331 19610 14361 19644
rect 13968 19605 14361 19610
rect 13968 19571 14122 19605
rect 14156 19576 14361 19605
rect 14156 19571 14297 19576
rect 13968 19542 14297 19571
rect 14331 19542 14361 19576
rect 13968 19533 14361 19542
rect 13968 19499 14122 19533
rect 14156 19508 14361 19533
rect 14156 19499 14297 19508
rect 13968 19474 14297 19499
rect 14331 19474 14361 19508
rect 13968 19461 14361 19474
rect 13968 19427 14122 19461
rect 14156 19440 14361 19461
rect 14156 19427 14297 19440
rect 13968 19406 14297 19427
rect 14331 19406 14361 19440
rect 13968 19389 14361 19406
rect 13968 19355 14122 19389
rect 14156 19372 14361 19389
rect 14156 19355 14297 19372
rect 13968 19338 14297 19355
rect 14331 19338 14361 19372
rect 13968 19317 14361 19338
rect 13968 19283 14122 19317
rect 14156 19304 14361 19317
rect 14156 19283 14297 19304
rect 13968 19270 14297 19283
rect 14331 19270 14361 19304
rect 13968 19245 14361 19270
rect 13968 19211 14122 19245
rect 14156 19236 14361 19245
rect 14156 19211 14297 19236
rect 13968 19202 14297 19211
rect 14331 19202 14361 19236
rect 13968 19173 14361 19202
rect 13968 19139 14122 19173
rect 14156 19168 14361 19173
rect 14156 19139 14297 19168
rect 13968 19134 14297 19139
rect 14331 19134 14361 19168
rect 13968 19101 14361 19134
rect 13968 19067 14122 19101
rect 14156 19100 14361 19101
rect 14156 19067 14297 19100
rect 13968 19066 14297 19067
rect 14331 19066 14361 19100
rect 13968 19032 14361 19066
rect 13968 19029 14297 19032
rect 13968 18995 14122 19029
rect 14156 18998 14297 19029
rect 14331 18998 14361 19032
rect 14156 18995 14361 18998
rect 13968 18964 14361 18995
rect 13968 18957 14297 18964
rect 13968 18923 14122 18957
rect 14156 18930 14297 18957
rect 14331 18930 14361 18964
rect 14156 18923 14361 18930
rect 13968 18896 14361 18923
rect 13968 18885 14297 18896
rect 13968 18851 14122 18885
rect 14156 18862 14297 18885
rect 14331 18862 14361 18896
rect 14156 18851 14361 18862
rect 13968 18828 14361 18851
rect 13968 18813 14297 18828
rect 13968 18779 14122 18813
rect 14156 18794 14297 18813
rect 14331 18794 14361 18828
rect 14156 18779 14361 18794
rect 13968 18760 14361 18779
rect 13968 18741 14297 18760
rect 13968 18707 14122 18741
rect 14156 18726 14297 18741
rect 14331 18726 14361 18760
rect 14156 18707 14361 18726
rect 13968 18692 14361 18707
rect 13968 18669 14297 18692
rect 13968 18635 14122 18669
rect 14156 18658 14297 18669
rect 14331 18658 14361 18692
rect 14156 18635 14361 18658
rect 13968 18624 14361 18635
rect 13968 18597 14297 18624
rect 13968 18563 14122 18597
rect 14156 18590 14297 18597
rect 14331 18590 14361 18624
rect 14156 18563 14361 18590
rect 13968 18556 14361 18563
rect 13968 18525 14297 18556
rect 13968 18491 14122 18525
rect 14156 18522 14297 18525
rect 14331 18522 14361 18556
rect 14156 18491 14361 18522
rect 13968 18488 14361 18491
rect 13968 18454 14297 18488
rect 14331 18454 14361 18488
rect 13968 18453 14361 18454
rect 13968 18419 14122 18453
rect 14156 18420 14361 18453
rect 14156 18419 14297 18420
rect 13968 18386 14297 18419
rect 14331 18386 14361 18420
rect 13968 18381 14361 18386
rect 13968 18347 14122 18381
rect 14156 18352 14361 18381
rect 14156 18347 14297 18352
rect 13968 18318 14297 18347
rect 14331 18318 14361 18352
rect 13968 18309 14361 18318
rect 13968 18275 14122 18309
rect 14156 18284 14361 18309
rect 14156 18275 14297 18284
rect 13968 18250 14297 18275
rect 14331 18250 14361 18284
rect 13968 18237 14361 18250
rect 13968 18203 14122 18237
rect 14156 18216 14361 18237
rect 14156 18203 14297 18216
rect 13968 18182 14297 18203
rect 14331 18182 14361 18216
rect 13968 18165 14361 18182
rect 13968 18131 14122 18165
rect 14156 18148 14361 18165
rect 14156 18131 14297 18148
rect 13968 18114 14297 18131
rect 14331 18114 14361 18148
rect 13968 18093 14361 18114
rect 13968 18059 14122 18093
rect 14156 18080 14361 18093
rect 14156 18059 14297 18080
rect 13968 18046 14297 18059
rect 14331 18046 14361 18080
rect 13968 18021 14361 18046
rect 13968 17987 14122 18021
rect 14156 18012 14361 18021
rect 14156 17987 14297 18012
rect 13968 17978 14297 17987
rect 14331 17978 14361 18012
rect 13968 17949 14361 17978
rect 13968 17915 14122 17949
rect 14156 17944 14361 17949
rect 14156 17915 14297 17944
rect 13968 17910 14297 17915
rect 14331 17910 14361 17944
rect 13968 17877 14361 17910
rect 13968 17843 14122 17877
rect 14156 17876 14361 17877
rect 14156 17843 14297 17876
rect 13968 17842 14297 17843
rect 14331 17842 14361 17876
rect 13968 17808 14361 17842
rect 13968 17805 14297 17808
rect 13968 17771 14122 17805
rect 14156 17774 14297 17805
rect 14331 17774 14361 17808
rect 14156 17771 14361 17774
rect 13968 17740 14361 17771
rect 13968 17733 14297 17740
rect 13968 17699 14122 17733
rect 14156 17706 14297 17733
rect 14331 17706 14361 17740
rect 14156 17699 14361 17706
rect 13968 17672 14361 17699
rect 13968 17661 14297 17672
rect 13968 17627 14122 17661
rect 14156 17638 14297 17661
rect 14331 17638 14361 17672
rect 14156 17627 14361 17638
rect 13968 17604 14361 17627
rect 13968 17589 14297 17604
rect 13968 17555 14122 17589
rect 14156 17570 14297 17589
rect 14331 17570 14361 17604
rect 14156 17555 14361 17570
rect 13968 17536 14361 17555
rect 13968 17517 14297 17536
rect 13968 17483 14122 17517
rect 14156 17502 14297 17517
rect 14331 17502 14361 17536
rect 14156 17483 14361 17502
rect 13968 17468 14361 17483
rect 13968 17445 14297 17468
rect 13968 17411 14122 17445
rect 14156 17434 14297 17445
rect 14331 17434 14361 17468
rect 14156 17411 14361 17434
rect 13968 17400 14361 17411
rect 13968 17373 14297 17400
rect 13968 17339 14122 17373
rect 14156 17366 14297 17373
rect 14331 17366 14361 17400
rect 14156 17339 14361 17366
rect 13968 17332 14361 17339
rect 13968 17301 14297 17332
rect 13968 17267 14122 17301
rect 14156 17298 14297 17301
rect 14331 17298 14361 17332
rect 14156 17267 14361 17298
rect 13968 17264 14361 17267
rect 13968 17230 14297 17264
rect 14331 17230 14361 17264
rect 13968 17229 14361 17230
rect 13968 17195 14122 17229
rect 14156 17196 14361 17229
rect 14156 17195 14297 17196
rect 13968 17162 14297 17195
rect 14331 17162 14361 17196
rect 13968 17157 14361 17162
rect 13968 17123 14122 17157
rect 14156 17128 14361 17157
rect 14156 17123 14297 17128
rect 13968 17094 14297 17123
rect 14331 17094 14361 17128
rect 13968 17085 14361 17094
rect 13968 17051 14122 17085
rect 14156 17060 14361 17085
rect 14156 17051 14297 17060
rect 13968 17026 14297 17051
rect 14331 17026 14361 17060
rect 13968 17013 14361 17026
rect 13968 16979 14122 17013
rect 14156 16992 14361 17013
rect 14156 16979 14297 16992
rect 13968 16958 14297 16979
rect 14331 16958 14361 16992
rect 13968 16941 14361 16958
rect 13968 16907 14122 16941
rect 14156 16924 14361 16941
rect 14156 16907 14297 16924
rect 13968 16890 14297 16907
rect 14331 16890 14361 16924
rect 13968 16869 14361 16890
rect 13968 16835 14122 16869
rect 14156 16856 14361 16869
rect 14156 16835 14297 16856
rect 13968 16822 14297 16835
rect 14331 16822 14361 16856
rect 13968 16797 14361 16822
rect 13968 16763 14122 16797
rect 14156 16788 14361 16797
rect 14156 16763 14297 16788
rect 13968 16754 14297 16763
rect 14331 16754 14361 16788
rect 13968 16725 14361 16754
rect 13968 16691 14122 16725
rect 14156 16720 14361 16725
rect 14156 16691 14297 16720
rect 13968 16686 14297 16691
rect 14331 16686 14361 16720
rect 13968 16653 14361 16686
rect 13968 16619 14122 16653
rect 14156 16652 14361 16653
rect 14156 16619 14297 16652
rect 13968 16618 14297 16619
rect 14331 16618 14361 16652
rect 13968 16584 14361 16618
rect 13968 16581 14297 16584
rect 13968 16547 14122 16581
rect 14156 16550 14297 16581
rect 14331 16550 14361 16584
rect 14156 16547 14361 16550
rect 13968 16516 14361 16547
rect 13968 16509 14297 16516
rect 13968 16475 14122 16509
rect 14156 16482 14297 16509
rect 14331 16482 14361 16516
rect 14156 16475 14361 16482
rect 13968 16448 14361 16475
rect 13968 16437 14297 16448
rect 13968 16403 14122 16437
rect 14156 16414 14297 16437
rect 14331 16414 14361 16448
rect 14156 16403 14361 16414
rect 13968 16380 14361 16403
rect 13968 16365 14297 16380
rect 13968 16331 14122 16365
rect 14156 16346 14297 16365
rect 14331 16346 14361 16380
rect 14156 16331 14361 16346
rect 13968 16312 14361 16331
rect 13968 16293 14297 16312
rect 13968 16259 14122 16293
rect 14156 16278 14297 16293
rect 14331 16278 14361 16312
rect 14156 16259 14361 16278
rect 13968 16244 14361 16259
rect 13968 16221 14297 16244
rect 13968 16187 14122 16221
rect 14156 16210 14297 16221
rect 14331 16210 14361 16244
rect 14156 16187 14361 16210
rect 13968 16176 14361 16187
rect 13968 16149 14297 16176
rect 13968 16115 14122 16149
rect 14156 16142 14297 16149
rect 14331 16142 14361 16176
rect 14156 16115 14361 16142
rect 13968 16108 14361 16115
rect 13968 16077 14297 16108
rect 13968 16043 14122 16077
rect 14156 16074 14297 16077
rect 14331 16074 14361 16108
rect 14156 16043 14361 16074
rect 13968 16040 14361 16043
rect 13968 16006 14297 16040
rect 14331 16006 14361 16040
rect 13968 16005 14361 16006
rect 13968 15971 14122 16005
rect 14156 15972 14361 16005
rect 14156 15971 14297 15972
rect 13968 15938 14297 15971
rect 14331 15938 14361 15972
rect 13968 15933 14361 15938
rect 13968 15899 14122 15933
rect 14156 15904 14361 15933
rect 14156 15899 14297 15904
rect 13968 15870 14297 15899
rect 14331 15870 14361 15904
rect 13968 15861 14361 15870
rect 13968 15827 14122 15861
rect 14156 15836 14361 15861
rect 14156 15827 14297 15836
rect 13968 15802 14297 15827
rect 14331 15802 14361 15836
rect 13968 15789 14361 15802
rect 13968 15755 14122 15789
rect 14156 15768 14361 15789
rect 14156 15755 14297 15768
rect 13968 15734 14297 15755
rect 14331 15734 14361 15768
rect 13968 15717 14361 15734
rect 13968 15683 14122 15717
rect 14156 15700 14361 15717
rect 14156 15683 14297 15700
rect 13968 15666 14297 15683
rect 14331 15666 14361 15700
rect 13968 15645 14361 15666
rect 13968 15611 14122 15645
rect 14156 15632 14361 15645
rect 14156 15611 14297 15632
rect 13968 15598 14297 15611
rect 14331 15598 14361 15632
rect 13968 15573 14361 15598
rect 13968 15539 14122 15573
rect 14156 15564 14361 15573
rect 14156 15539 14297 15564
rect 13968 15530 14297 15539
rect 14331 15530 14361 15564
rect 13968 15501 14361 15530
rect 13968 15467 14122 15501
rect 14156 15496 14361 15501
rect 14156 15467 14297 15496
rect 13968 15462 14297 15467
rect 14331 15462 14361 15496
rect 13968 15429 14361 15462
rect 13968 15395 14122 15429
rect 14156 15428 14361 15429
rect 14156 15395 14297 15428
rect 13968 15394 14297 15395
rect 14331 15394 14361 15428
rect 13968 15360 14361 15394
rect 13968 15357 14297 15360
rect 13968 15323 14122 15357
rect 14156 15326 14297 15357
rect 14331 15326 14361 15360
rect 14156 15323 14361 15326
rect 13968 15292 14361 15323
rect 13968 15285 14297 15292
rect 13968 15251 14122 15285
rect 14156 15258 14297 15285
rect 14331 15258 14361 15292
rect 14156 15251 14361 15258
rect 13968 15224 14361 15251
rect 13968 15213 14297 15224
rect 13968 15179 14122 15213
rect 14156 15190 14297 15213
rect 14331 15190 14361 15224
rect 14156 15179 14361 15190
rect 13968 15156 14361 15179
rect 13968 15141 14297 15156
rect 13968 15107 14122 15141
rect 14156 15122 14297 15141
rect 14331 15122 14361 15156
rect 14156 15107 14361 15122
rect 13968 15088 14361 15107
rect 13968 15069 14297 15088
rect 13968 15035 14122 15069
rect 14156 15054 14297 15069
rect 14331 15054 14361 15088
rect 14156 15035 14361 15054
rect 13968 15020 14361 15035
rect 13968 14997 14297 15020
rect 13968 14963 14122 14997
rect 14156 14986 14297 14997
rect 14331 14986 14361 15020
rect 14156 14963 14361 14986
rect 13968 14952 14361 14963
rect 13968 14925 14297 14952
rect 13968 14891 14122 14925
rect 14156 14918 14297 14925
rect 14331 14918 14361 14952
rect 14156 14891 14361 14918
rect 13968 14884 14361 14891
rect 13968 14853 14297 14884
rect 13968 14819 14122 14853
rect 14156 14850 14297 14853
rect 14331 14850 14361 14884
rect 14156 14819 14361 14850
rect 13968 14816 14361 14819
rect 13968 14782 14297 14816
rect 14331 14782 14361 14816
rect 13968 14781 14361 14782
rect 13968 14747 14122 14781
rect 14156 14748 14361 14781
rect 14156 14747 14297 14748
rect 13968 14714 14297 14747
rect 14331 14714 14361 14748
rect 13968 14709 14361 14714
rect 13968 14675 14122 14709
rect 14156 14680 14361 14709
rect 14156 14675 14297 14680
rect 13968 14646 14297 14675
rect 14331 14646 14361 14680
rect 13968 14637 14361 14646
rect 13968 14603 14122 14637
rect 14156 14612 14361 14637
rect 14156 14603 14297 14612
rect 13968 14578 14297 14603
rect 14331 14578 14361 14612
rect 13968 14565 14361 14578
rect 13968 14531 14122 14565
rect 14156 14544 14361 14565
rect 14156 14531 14297 14544
rect 13968 14510 14297 14531
rect 14331 14510 14361 14544
rect 13968 14493 14361 14510
rect 13968 14459 14122 14493
rect 14156 14476 14361 14493
rect 14156 14459 14297 14476
rect 13968 14442 14297 14459
rect 14331 14442 14361 14476
rect 13968 14421 14361 14442
rect 13968 14387 14122 14421
rect 14156 14408 14361 14421
rect 14156 14387 14297 14408
rect 13968 14374 14297 14387
rect 14331 14374 14361 14408
rect 13968 14349 14361 14374
rect 13968 14315 14122 14349
rect 14156 14340 14361 14349
rect 14156 14315 14297 14340
rect 13968 14306 14297 14315
rect 14331 14306 14361 14340
rect 13968 14277 14361 14306
rect 13968 14243 14122 14277
rect 14156 14272 14361 14277
rect 14156 14243 14297 14272
rect 13968 14238 14297 14243
rect 14331 14238 14361 14272
rect 13968 14205 14361 14238
rect 13968 14171 14122 14205
rect 14156 14204 14361 14205
rect 14156 14171 14297 14204
rect 13968 14170 14297 14171
rect 14331 14170 14361 14204
rect 13968 14136 14361 14170
rect 13968 14133 14297 14136
rect 13968 14099 14122 14133
rect 14156 14102 14297 14133
rect 14331 14102 14361 14136
rect 14156 14099 14361 14102
rect 13968 14068 14361 14099
rect 13968 14061 14297 14068
rect 13968 14027 14122 14061
rect 14156 14034 14297 14061
rect 14331 14034 14361 14068
rect 14156 14027 14361 14034
rect 13968 14000 14361 14027
rect 13968 13989 14297 14000
rect 13968 13955 14122 13989
rect 14156 13966 14297 13989
rect 14331 13966 14361 14000
rect 14156 13955 14361 13966
rect 13968 13932 14361 13955
rect 13968 13917 14297 13932
rect 13968 13883 14122 13917
rect 14156 13898 14297 13917
rect 14331 13898 14361 13932
rect 14156 13883 14361 13898
rect 13968 13864 14361 13883
rect 13968 13845 14297 13864
rect 13968 13811 14122 13845
rect 14156 13830 14297 13845
rect 14331 13830 14361 13864
rect 14156 13811 14361 13830
rect 13968 13796 14361 13811
rect 13968 13773 14297 13796
rect 13968 13739 14122 13773
rect 14156 13762 14297 13773
rect 14331 13762 14361 13796
rect 14156 13739 14361 13762
rect 13968 13728 14361 13739
rect 13968 13701 14297 13728
rect 13968 13667 14122 13701
rect 14156 13694 14297 13701
rect 14331 13694 14361 13728
rect 14156 13667 14361 13694
rect 13968 13660 14361 13667
rect 13968 13629 14297 13660
rect 13968 13595 14122 13629
rect 14156 13626 14297 13629
rect 14331 13626 14361 13660
rect 14156 13595 14361 13626
rect 13968 13592 14361 13595
rect 13968 13558 14297 13592
rect 14331 13558 14361 13592
rect 13968 13557 14361 13558
rect 13968 13523 14122 13557
rect 14156 13524 14361 13557
rect 14156 13523 14297 13524
rect 13968 13490 14297 13523
rect 14331 13490 14361 13524
rect 13968 13485 14361 13490
rect 13968 13451 14122 13485
rect 14156 13456 14361 13485
rect 14156 13451 14297 13456
rect 13968 13422 14297 13451
rect 14331 13422 14361 13456
rect 13968 13413 14361 13422
rect 13968 13379 14122 13413
rect 14156 13388 14361 13413
rect 14156 13379 14297 13388
rect 13968 13354 14297 13379
rect 14331 13354 14361 13388
rect 13968 13341 14361 13354
rect 13968 13307 14122 13341
rect 14156 13320 14361 13341
rect 14156 13307 14297 13320
rect 13968 13286 14297 13307
rect 14331 13286 14361 13320
rect 13968 13269 14361 13286
rect 13968 13235 14122 13269
rect 14156 13252 14361 13269
rect 14156 13235 14297 13252
rect 13968 13218 14297 13235
rect 14331 13218 14361 13252
rect 13968 13197 14361 13218
rect 13968 13163 14122 13197
rect 14156 13184 14361 13197
rect 14156 13163 14297 13184
rect 13968 13150 14297 13163
rect 14331 13150 14361 13184
rect 13968 13125 14361 13150
rect 13968 13091 14122 13125
rect 14156 13116 14361 13125
rect 14156 13091 14297 13116
rect 13968 13082 14297 13091
rect 14331 13082 14361 13116
rect 13968 13053 14361 13082
rect 13968 13019 14122 13053
rect 14156 13048 14361 13053
rect 14156 13019 14297 13048
rect 13968 13014 14297 13019
rect 14331 13014 14361 13048
rect 13968 12981 14361 13014
rect 13968 12947 14122 12981
rect 14156 12980 14361 12981
rect 14156 12947 14297 12980
rect 13968 12946 14297 12947
rect 14331 12946 14361 12980
rect 13968 12912 14361 12946
rect 13968 12909 14297 12912
rect 13968 12875 14122 12909
rect 14156 12878 14297 12909
rect 14331 12878 14361 12912
rect 14156 12875 14361 12878
rect 13968 12844 14361 12875
rect 13968 12837 14297 12844
rect 13968 12803 14122 12837
rect 14156 12810 14297 12837
rect 14331 12810 14361 12844
rect 14156 12803 14361 12810
rect 13968 12776 14361 12803
rect 13968 12765 14297 12776
rect 13968 12731 14122 12765
rect 14156 12742 14297 12765
rect 14331 12742 14361 12776
rect 14156 12731 14361 12742
rect 13968 12708 14361 12731
rect 13968 12693 14297 12708
rect 13968 12659 14122 12693
rect 14156 12674 14297 12693
rect 14331 12674 14361 12708
rect 14156 12659 14361 12674
rect 13968 12640 14361 12659
rect 13968 12621 14297 12640
rect 13968 12587 14122 12621
rect 14156 12606 14297 12621
rect 14331 12606 14361 12640
rect 14156 12587 14361 12606
rect 13968 12572 14361 12587
rect 13968 12549 14297 12572
rect 13968 12515 14122 12549
rect 14156 12538 14297 12549
rect 14331 12538 14361 12572
rect 14156 12515 14361 12538
rect 13968 12504 14361 12515
rect 13968 12477 14297 12504
rect 13968 12443 14122 12477
rect 14156 12470 14297 12477
rect 14331 12470 14361 12504
rect 14156 12443 14361 12470
rect 13968 12436 14361 12443
rect 13968 12405 14297 12436
rect 13968 12371 14122 12405
rect 14156 12402 14297 12405
rect 14331 12402 14361 12436
rect 14156 12371 14361 12402
rect 13968 12368 14361 12371
rect 13968 12334 14297 12368
rect 14331 12334 14361 12368
rect 13968 12333 14361 12334
rect 13968 12299 14122 12333
rect 14156 12300 14361 12333
rect 14156 12299 14297 12300
rect 13968 12266 14297 12299
rect 14331 12266 14361 12300
rect 13968 12261 14361 12266
rect 13968 12227 14122 12261
rect 14156 12232 14361 12261
rect 14156 12227 14297 12232
rect 13968 12198 14297 12227
rect 14331 12198 14361 12232
rect 13968 12189 14361 12198
rect 13968 12155 14122 12189
rect 14156 12164 14361 12189
rect 14156 12155 14297 12164
rect 13968 12130 14297 12155
rect 14331 12130 14361 12164
rect 13968 12117 14361 12130
rect 13968 12083 14122 12117
rect 14156 12096 14361 12117
rect 14156 12083 14297 12096
rect 13968 12062 14297 12083
rect 14331 12062 14361 12096
rect 13968 12045 14361 12062
rect 13968 12011 14122 12045
rect 14156 12028 14361 12045
rect 14156 12011 14297 12028
rect 13968 11994 14297 12011
rect 14331 11994 14361 12028
rect 13968 11973 14361 11994
rect 13968 11939 14122 11973
rect 14156 11960 14361 11973
rect 14156 11939 14297 11960
rect 13968 11926 14297 11939
rect 14331 11926 14361 11960
rect 13968 11901 14361 11926
rect 13968 11867 14122 11901
rect 14156 11892 14361 11901
rect 14156 11867 14297 11892
rect 13968 11858 14297 11867
rect 14331 11858 14361 11892
rect 13968 11829 14361 11858
rect 13968 11795 14122 11829
rect 14156 11824 14361 11829
rect 14156 11795 14297 11824
rect 13968 11790 14297 11795
rect 14331 11790 14361 11824
rect 13968 11757 14361 11790
rect 13968 11723 14122 11757
rect 14156 11756 14361 11757
rect 14156 11723 14297 11756
rect 13968 11722 14297 11723
rect 14331 11722 14361 11756
rect 13968 11688 14361 11722
rect 13968 11685 14297 11688
rect 13968 11651 14122 11685
rect 14156 11654 14297 11685
rect 14331 11654 14361 11688
rect 14156 11651 14361 11654
rect 13968 11620 14361 11651
rect 13968 11613 14297 11620
rect 13968 11579 14122 11613
rect 14156 11586 14297 11613
rect 14331 11586 14361 11620
rect 14156 11579 14361 11586
rect 13968 11552 14361 11579
rect 13968 11541 14297 11552
rect 13968 11507 14122 11541
rect 14156 11518 14297 11541
rect 14331 11518 14361 11552
rect 14156 11507 14361 11518
rect 13968 11484 14361 11507
rect 13968 11469 14297 11484
rect 13968 11435 14122 11469
rect 14156 11450 14297 11469
rect 14331 11450 14361 11484
rect 14156 11435 14361 11450
rect 13968 11416 14361 11435
rect 13968 11397 14297 11416
rect 13968 11363 14122 11397
rect 14156 11382 14297 11397
rect 14331 11382 14361 11416
rect 14156 11363 14361 11382
rect 13968 11348 14361 11363
rect 13968 11325 14297 11348
rect 13968 11291 14122 11325
rect 14156 11314 14297 11325
rect 14331 11314 14361 11348
rect 14156 11291 14361 11314
rect 13968 11280 14361 11291
rect 13968 11253 14297 11280
rect 13968 11219 14122 11253
rect 14156 11246 14297 11253
rect 14331 11246 14361 11280
rect 14156 11219 14361 11246
rect 13968 11212 14361 11219
rect 13968 11181 14297 11212
rect 13968 11147 14122 11181
rect 14156 11178 14297 11181
rect 14331 11178 14361 11212
rect 14156 11147 14361 11178
rect 13968 11144 14361 11147
rect 13968 11110 14297 11144
rect 14331 11110 14361 11144
rect 13968 11109 14361 11110
rect 13968 11075 14122 11109
rect 14156 11076 14361 11109
rect 14156 11075 14297 11076
rect 13968 11042 14297 11075
rect 14331 11042 14361 11076
rect 13968 11037 14361 11042
rect 13968 11003 14122 11037
rect 14156 11008 14361 11037
rect 14156 11003 14297 11008
rect 13968 10974 14297 11003
rect 14331 10974 14361 11008
rect 13968 10965 14361 10974
rect 13968 10931 14122 10965
rect 14156 10940 14361 10965
rect 14156 10931 14297 10940
rect 13968 10906 14297 10931
rect 14331 10906 14361 10940
rect 13968 10893 14361 10906
rect 13968 10859 14122 10893
rect 14156 10872 14361 10893
rect 14156 10859 14297 10872
rect 13968 10838 14297 10859
rect 14331 10838 14361 10872
rect 13968 10821 14361 10838
rect 13968 10787 14122 10821
rect 14156 10804 14361 10821
rect 14156 10787 14297 10804
rect 13968 10770 14297 10787
rect 14331 10770 14361 10804
rect 13968 10749 14361 10770
rect 13968 10715 14122 10749
rect 14156 10736 14361 10749
rect 14156 10715 14297 10736
rect 13968 10702 14297 10715
rect 14331 10702 14361 10736
rect 13968 10677 14361 10702
rect 13968 10643 14122 10677
rect 14156 10668 14361 10677
rect 14156 10643 14297 10668
rect 13968 10634 14297 10643
rect 14331 10634 14361 10668
rect 13968 10605 14361 10634
rect 13968 10571 14122 10605
rect 14156 10600 14361 10605
rect 14156 10571 14297 10600
rect 13968 10566 14297 10571
rect 14331 10566 14361 10600
rect 13968 10533 14361 10566
rect 13968 10499 14122 10533
rect 14156 10532 14361 10533
rect 14156 10499 14297 10532
rect 13968 10498 14297 10499
rect 14331 10498 14361 10532
rect 13968 10464 14361 10498
rect 13968 10461 14297 10464
rect 13968 10427 14122 10461
rect 14156 10430 14297 10461
rect 14331 10430 14361 10464
rect 14156 10427 14361 10430
rect 13968 10396 14361 10427
rect 13968 10389 14297 10396
rect 13968 10355 14122 10389
rect 14156 10362 14297 10389
rect 14331 10362 14361 10396
rect 14156 10355 14361 10362
rect 13968 10328 14361 10355
rect 13968 10317 14297 10328
rect 13968 10283 14122 10317
rect 14156 10294 14297 10317
rect 14331 10294 14361 10328
rect 14156 10283 14361 10294
rect 13968 10260 14361 10283
rect 13968 10245 14297 10260
rect 13968 10211 14122 10245
rect 14156 10226 14297 10245
rect 14331 10226 14361 10260
rect 14156 10211 14361 10226
rect 603 10158 632 10192
rect 666 10180 1026 10192
rect 666 10158 807 10180
rect 603 10146 807 10158
rect 841 10146 1026 10180
rect 603 10124 1026 10146
rect 603 10090 632 10124
rect 666 10108 1026 10124
rect 666 10090 807 10108
rect 603 10074 807 10090
rect 841 10088 1026 10108
rect 13968 10192 14361 10211
rect 13968 10173 14297 10192
rect 13968 10139 14122 10173
rect 14156 10158 14297 10173
rect 14331 10158 14361 10192
rect 14156 10139 14361 10158
rect 13968 10124 14361 10139
rect 13968 10101 14297 10124
rect 13968 10088 14122 10101
rect 841 10074 14122 10088
rect 603 10067 14122 10074
rect 14156 10090 14297 10101
rect 14331 10090 14361 10124
rect 14156 10067 14361 10090
rect 603 10056 14361 10067
rect 603 10022 632 10056
rect 666 10022 14297 10056
rect 14331 10022 14361 10056
rect 603 9988 14361 10022
rect 603 9954 632 9988
rect 666 9954 14297 9988
rect 14331 9954 14361 9988
rect 603 9942 14361 9954
rect 603 9920 891 9942
rect 603 9886 632 9920
rect 666 9908 891 9920
rect 925 9908 963 9942
rect 997 9908 1035 9942
rect 1069 9908 1107 9942
rect 1141 9908 1179 9942
rect 1213 9908 1251 9942
rect 1285 9908 1323 9942
rect 1357 9908 1395 9942
rect 1429 9908 1467 9942
rect 1501 9908 1539 9942
rect 1573 9908 1611 9942
rect 1645 9908 1683 9942
rect 1717 9908 1755 9942
rect 1789 9908 1827 9942
rect 1861 9908 1899 9942
rect 1933 9908 1971 9942
rect 2005 9908 2043 9942
rect 2077 9908 2115 9942
rect 2149 9908 2187 9942
rect 2221 9908 2259 9942
rect 2293 9908 2331 9942
rect 2365 9908 2403 9942
rect 2437 9908 2475 9942
rect 2509 9908 2547 9942
rect 2581 9908 2619 9942
rect 2653 9908 2691 9942
rect 2725 9908 2763 9942
rect 2797 9908 2835 9942
rect 2869 9908 2907 9942
rect 2941 9908 2979 9942
rect 3013 9908 3051 9942
rect 3085 9908 3123 9942
rect 3157 9908 3195 9942
rect 3229 9908 3267 9942
rect 3301 9908 3339 9942
rect 3373 9908 3411 9942
rect 3445 9908 3483 9942
rect 3517 9908 3555 9942
rect 3589 9908 3627 9942
rect 3661 9908 3699 9942
rect 3733 9908 3771 9942
rect 3805 9908 3843 9942
rect 3877 9908 3915 9942
rect 3949 9908 3987 9942
rect 4021 9908 4059 9942
rect 4093 9908 4131 9942
rect 4165 9908 4203 9942
rect 4237 9908 4275 9942
rect 4309 9908 4347 9942
rect 4381 9908 4419 9942
rect 4453 9908 4491 9942
rect 4525 9908 4563 9942
rect 4597 9908 4635 9942
rect 4669 9908 4707 9942
rect 4741 9908 4779 9942
rect 4813 9908 4851 9942
rect 4885 9908 4923 9942
rect 4957 9908 4995 9942
rect 5029 9908 5067 9942
rect 5101 9908 5139 9942
rect 5173 9908 5211 9942
rect 5245 9908 5283 9942
rect 5317 9908 5355 9942
rect 5389 9908 5427 9942
rect 5461 9908 5499 9942
rect 5533 9908 5571 9942
rect 5605 9908 5643 9942
rect 5677 9908 5715 9942
rect 5749 9908 5787 9942
rect 5821 9908 5859 9942
rect 5893 9908 5931 9942
rect 5965 9908 6003 9942
rect 6037 9908 6075 9942
rect 6109 9908 6147 9942
rect 6181 9908 6219 9942
rect 6253 9908 6291 9942
rect 6325 9908 6363 9942
rect 6397 9908 6435 9942
rect 6469 9908 6507 9942
rect 6541 9908 6579 9942
rect 6613 9908 6651 9942
rect 6685 9908 6723 9942
rect 6757 9908 6795 9942
rect 6829 9908 6867 9942
rect 6901 9908 6939 9942
rect 6973 9908 7011 9942
rect 7045 9908 7083 9942
rect 7117 9908 7155 9942
rect 7189 9908 7227 9942
rect 7261 9908 7299 9942
rect 7333 9908 7371 9942
rect 7405 9908 7443 9942
rect 7477 9908 7515 9942
rect 7549 9908 7587 9942
rect 7621 9908 7659 9942
rect 7693 9908 7731 9942
rect 7765 9908 7803 9942
rect 7837 9908 7875 9942
rect 7909 9908 7947 9942
rect 7981 9908 8019 9942
rect 8053 9908 8091 9942
rect 8125 9908 8163 9942
rect 8197 9908 8235 9942
rect 8269 9908 8307 9942
rect 8341 9908 8379 9942
rect 8413 9908 8451 9942
rect 8485 9908 8523 9942
rect 8557 9908 8595 9942
rect 8629 9908 8667 9942
rect 8701 9908 8739 9942
rect 8773 9908 8811 9942
rect 8845 9908 8883 9942
rect 8917 9908 8955 9942
rect 8989 9908 9027 9942
rect 9061 9908 9099 9942
rect 9133 9908 9171 9942
rect 9205 9908 9243 9942
rect 9277 9908 9315 9942
rect 9349 9908 9387 9942
rect 9421 9908 9459 9942
rect 9493 9908 9531 9942
rect 9565 9908 9603 9942
rect 9637 9908 9675 9942
rect 9709 9908 9747 9942
rect 9781 9908 9819 9942
rect 9853 9908 9891 9942
rect 9925 9908 9963 9942
rect 9997 9908 10035 9942
rect 10069 9908 10107 9942
rect 10141 9908 10179 9942
rect 10213 9908 10251 9942
rect 10285 9908 10323 9942
rect 10357 9908 10395 9942
rect 10429 9908 10467 9942
rect 10501 9908 10539 9942
rect 10573 9908 10611 9942
rect 10645 9908 10683 9942
rect 10717 9908 10755 9942
rect 10789 9908 10827 9942
rect 10861 9908 10899 9942
rect 10933 9908 10971 9942
rect 11005 9908 11043 9942
rect 11077 9908 11115 9942
rect 11149 9908 11187 9942
rect 11221 9908 11259 9942
rect 11293 9908 11331 9942
rect 11365 9908 11403 9942
rect 11437 9908 11475 9942
rect 11509 9908 11547 9942
rect 11581 9908 11619 9942
rect 11653 9908 11691 9942
rect 11725 9908 11763 9942
rect 11797 9908 11835 9942
rect 11869 9908 11907 9942
rect 11941 9908 11979 9942
rect 12013 9908 12051 9942
rect 12085 9908 12123 9942
rect 12157 9908 12195 9942
rect 12229 9908 12267 9942
rect 12301 9908 12339 9942
rect 12373 9908 12411 9942
rect 12445 9908 12483 9942
rect 12517 9908 12555 9942
rect 12589 9908 12627 9942
rect 12661 9908 12699 9942
rect 12733 9908 12771 9942
rect 12805 9908 12843 9942
rect 12877 9908 12915 9942
rect 12949 9908 12987 9942
rect 13021 9908 13059 9942
rect 13093 9908 13131 9942
rect 13165 9908 13203 9942
rect 13237 9908 13275 9942
rect 13309 9908 13347 9942
rect 13381 9908 13419 9942
rect 13453 9908 13491 9942
rect 13525 9908 13563 9942
rect 13597 9908 13635 9942
rect 13669 9908 13707 9942
rect 13741 9908 13779 9942
rect 13813 9908 13851 9942
rect 13885 9908 13923 9942
rect 13957 9908 13995 9942
rect 14029 9920 14361 9942
rect 14029 9908 14297 9920
rect 666 9886 14297 9908
rect 14331 9886 14361 9920
rect 603 9775 14361 9886
rect 603 9741 766 9775
rect 800 9741 834 9775
rect 868 9774 902 9775
rect 936 9774 970 9775
rect 1004 9774 1038 9775
rect 1072 9774 1106 9775
rect 1140 9774 1174 9775
rect 868 9741 883 9774
rect 936 9741 955 9774
rect 1004 9741 1027 9774
rect 1072 9741 1099 9774
rect 1140 9741 1171 9774
rect 1208 9741 1242 9775
rect 1276 9774 1310 9775
rect 1344 9774 1378 9775
rect 1412 9774 1446 9775
rect 1480 9774 1514 9775
rect 1548 9774 1582 9775
rect 1616 9774 1650 9775
rect 1684 9774 1718 9775
rect 1752 9774 1786 9775
rect 1820 9774 1854 9775
rect 1277 9741 1310 9774
rect 1349 9741 1378 9774
rect 1421 9741 1446 9774
rect 1493 9741 1514 9774
rect 1565 9741 1582 9774
rect 1637 9741 1650 9774
rect 1709 9741 1718 9774
rect 1781 9741 1786 9774
rect 1853 9741 1854 9774
rect 1888 9774 1922 9775
rect 1956 9774 1990 9775
rect 2024 9774 2058 9775
rect 1888 9741 1891 9774
rect 1956 9741 1963 9774
rect 2024 9741 2035 9774
rect 2092 9741 2126 9775
rect 2160 9741 2194 9775
rect 2228 9741 2262 9775
rect 2296 9741 2330 9775
rect 2364 9741 2398 9775
rect 2432 9741 2466 9775
rect 2500 9741 2534 9775
rect 2568 9741 2602 9775
rect 2636 9741 2670 9775
rect 2704 9741 2738 9775
rect 2772 9741 2806 9775
rect 2840 9741 2874 9775
rect 2908 9741 2942 9775
rect 2976 9741 3010 9775
rect 3044 9741 3078 9775
rect 3112 9741 3146 9775
rect 3180 9741 3214 9775
rect 3248 9741 3282 9775
rect 3316 9741 3350 9775
rect 3384 9741 3418 9775
rect 3452 9741 3486 9775
rect 3520 9741 3554 9775
rect 3588 9741 3622 9775
rect 3656 9741 3690 9775
rect 3724 9741 3758 9775
rect 3792 9741 3826 9775
rect 3860 9741 3894 9775
rect 3928 9741 3962 9775
rect 3996 9741 4030 9775
rect 4064 9741 4098 9775
rect 4132 9741 4166 9775
rect 4200 9741 4234 9775
rect 4268 9741 4302 9775
rect 4336 9741 4370 9775
rect 4404 9741 4438 9775
rect 4472 9741 4506 9775
rect 4540 9741 4574 9775
rect 4608 9741 4642 9775
rect 4676 9741 4710 9775
rect 4744 9741 4778 9775
rect 4812 9741 4846 9775
rect 4880 9741 4914 9775
rect 4948 9741 4982 9775
rect 5016 9741 5050 9775
rect 5084 9741 5118 9775
rect 5152 9741 5186 9775
rect 5220 9741 5254 9775
rect 5288 9741 5322 9775
rect 5356 9741 5390 9775
rect 5424 9741 5458 9775
rect 5492 9741 5526 9775
rect 5560 9741 5594 9775
rect 5628 9741 5662 9775
rect 5696 9741 5730 9775
rect 5764 9741 5798 9775
rect 5832 9741 5866 9775
rect 5900 9741 5934 9775
rect 5968 9741 6002 9775
rect 6036 9741 6070 9775
rect 6104 9741 6138 9775
rect 6172 9741 6206 9775
rect 6240 9741 6274 9775
rect 6308 9741 6342 9775
rect 6376 9741 6410 9775
rect 6444 9741 6478 9775
rect 6512 9741 6546 9775
rect 6580 9741 6614 9775
rect 6648 9741 6682 9775
rect 6716 9741 6750 9775
rect 6784 9741 6818 9775
rect 6852 9741 6886 9775
rect 6920 9741 6954 9775
rect 6988 9741 7022 9775
rect 7056 9741 7090 9775
rect 7124 9741 7158 9775
rect 7192 9741 7226 9775
rect 7260 9741 7294 9775
rect 7328 9741 7362 9775
rect 7396 9741 7430 9775
rect 7464 9741 7498 9775
rect 7532 9741 7566 9775
rect 7600 9741 7634 9775
rect 7668 9741 7702 9775
rect 7736 9741 7770 9775
rect 7804 9741 7838 9775
rect 7872 9741 7906 9775
rect 7940 9741 7974 9775
rect 8008 9741 8042 9775
rect 8076 9741 8110 9775
rect 8144 9741 8178 9775
rect 8212 9741 8246 9775
rect 8280 9741 8314 9775
rect 8348 9741 8382 9775
rect 8416 9741 8450 9775
rect 8484 9741 8518 9775
rect 8552 9741 8586 9775
rect 8620 9741 8654 9775
rect 8688 9741 8722 9775
rect 8756 9741 8790 9775
rect 8824 9741 8858 9775
rect 8892 9741 8926 9775
rect 8960 9741 8994 9775
rect 9028 9741 9062 9775
rect 9096 9741 9130 9775
rect 9164 9741 9198 9775
rect 9232 9741 9266 9775
rect 9300 9741 9334 9775
rect 9368 9741 9402 9775
rect 9436 9741 9470 9775
rect 9504 9741 9538 9775
rect 9572 9741 9606 9775
rect 9640 9741 9674 9775
rect 9708 9741 9742 9775
rect 9776 9741 9810 9775
rect 9844 9741 9878 9775
rect 9912 9741 9946 9775
rect 9980 9741 10014 9775
rect 10048 9741 10082 9775
rect 10116 9741 10150 9775
rect 10184 9741 10218 9775
rect 10252 9741 10286 9775
rect 10320 9741 10354 9775
rect 10388 9741 10422 9775
rect 10456 9741 10490 9775
rect 10524 9741 10558 9775
rect 10592 9741 10626 9775
rect 10660 9741 10694 9775
rect 10728 9741 10762 9775
rect 10796 9741 10830 9775
rect 10864 9741 10898 9775
rect 10932 9741 10966 9775
rect 11000 9741 11034 9775
rect 11068 9741 11102 9775
rect 11136 9741 11170 9775
rect 11204 9741 11238 9775
rect 11272 9741 11306 9775
rect 11340 9741 11374 9775
rect 11408 9741 11442 9775
rect 11476 9741 11510 9775
rect 11544 9741 11578 9775
rect 11612 9741 11646 9775
rect 11680 9741 11714 9775
rect 11748 9741 11782 9775
rect 11816 9741 11850 9775
rect 11884 9741 11918 9775
rect 11952 9741 11986 9775
rect 12020 9741 12054 9775
rect 12088 9741 12122 9775
rect 12156 9741 12190 9775
rect 12224 9741 12258 9775
rect 12292 9741 12326 9775
rect 12360 9741 12394 9775
rect 12428 9741 12462 9775
rect 12496 9741 12530 9775
rect 12564 9741 12598 9775
rect 12632 9741 12666 9775
rect 12700 9741 12734 9775
rect 12768 9741 12802 9775
rect 12836 9741 12870 9775
rect 12904 9774 12938 9775
rect 12972 9774 13006 9775
rect 13040 9774 13074 9775
rect 13108 9774 13142 9775
rect 13176 9774 13210 9775
rect 13244 9774 13278 9775
rect 12917 9741 12938 9774
rect 12989 9741 13006 9774
rect 13061 9741 13074 9774
rect 13133 9741 13142 9774
rect 13205 9741 13210 9774
rect 13277 9741 13278 9774
rect 13312 9774 13346 9775
rect 13380 9774 13414 9775
rect 13448 9774 13482 9775
rect 13516 9774 13550 9775
rect 13584 9774 13618 9775
rect 13652 9774 13686 9775
rect 13720 9774 13754 9775
rect 13788 9774 13822 9775
rect 13312 9741 13315 9774
rect 13380 9741 13387 9774
rect 13448 9741 13459 9774
rect 13516 9741 13531 9774
rect 13584 9741 13603 9774
rect 13652 9741 13675 9774
rect 13720 9741 13747 9774
rect 13788 9741 13819 9774
rect 13856 9741 13890 9775
rect 13924 9774 13958 9775
rect 13992 9774 14026 9775
rect 14060 9774 14094 9775
rect 13925 9741 13958 9774
rect 13997 9741 14026 9774
rect 14069 9741 14094 9774
rect 14128 9741 14162 9775
rect 14196 9741 14361 9775
rect 603 9740 883 9741
rect 917 9740 955 9741
rect 989 9740 1027 9741
rect 1061 9740 1099 9741
rect 1133 9740 1171 9741
rect 1205 9740 1243 9741
rect 1277 9740 1315 9741
rect 1349 9740 1387 9741
rect 1421 9740 1459 9741
rect 1493 9740 1531 9741
rect 1565 9740 1603 9741
rect 1637 9740 1675 9741
rect 1709 9740 1747 9741
rect 1781 9740 1819 9741
rect 1853 9740 1891 9741
rect 1925 9740 1963 9741
rect 1997 9740 2035 9741
rect 2069 9740 12883 9741
rect 12917 9740 12955 9741
rect 12989 9740 13027 9741
rect 13061 9740 13099 9741
rect 13133 9740 13171 9741
rect 13205 9740 13243 9741
rect 13277 9740 13315 9741
rect 13349 9740 13387 9741
rect 13421 9740 13459 9741
rect 13493 9740 13531 9741
rect 13565 9740 13603 9741
rect 13637 9740 13675 9741
rect 13709 9740 13747 9741
rect 13781 9740 13819 9741
rect 13853 9740 13891 9741
rect 13925 9740 13963 9741
rect 13997 9740 14035 9741
rect 14069 9740 14361 9741
rect 603 9711 14361 9740
rect 14539 36174 14607 36208
rect 14641 36190 14724 36208
rect 14539 36156 14614 36174
rect 14648 36156 14724 36190
rect 14539 36140 14724 36156
rect 14539 36106 14607 36140
rect 14641 36118 14724 36140
rect 14539 36084 14614 36106
rect 14648 36084 14724 36118
rect 14539 36072 14724 36084
rect 14539 36038 14607 36072
rect 14641 36046 14724 36072
rect 14539 36012 14614 36038
rect 14648 36012 14724 36046
rect 14539 36004 14724 36012
rect 14539 35970 14607 36004
rect 14641 35974 14724 36004
rect 14539 35940 14614 35970
rect 14648 35940 14724 35974
rect 14539 35936 14724 35940
rect 14539 35902 14607 35936
rect 14641 35902 14724 35936
rect 14539 35868 14614 35902
rect 14648 35868 14724 35902
rect 14539 35834 14607 35868
rect 14641 35834 14724 35868
rect 14539 35830 14724 35834
rect 14539 35800 14614 35830
rect 14539 35766 14607 35800
rect 14648 35796 14724 35830
rect 14641 35766 14724 35796
rect 14539 35758 14724 35766
rect 14539 35732 14614 35758
rect 14539 35698 14607 35732
rect 14648 35724 14724 35758
rect 14641 35698 14724 35724
rect 14539 35686 14724 35698
rect 14539 35664 14614 35686
rect 14539 35630 14607 35664
rect 14648 35652 14724 35686
rect 14641 35630 14724 35652
rect 14539 35614 14724 35630
rect 14539 35596 14614 35614
rect 14539 35562 14607 35596
rect 14648 35580 14724 35614
rect 14641 35562 14724 35580
rect 14539 35542 14724 35562
rect 14539 35528 14614 35542
rect 14539 35494 14607 35528
rect 14648 35508 14724 35542
rect 14641 35494 14724 35508
rect 14539 35470 14724 35494
rect 14539 35460 14614 35470
rect 14539 35426 14607 35460
rect 14648 35436 14724 35470
rect 14641 35426 14724 35436
rect 14539 35398 14724 35426
rect 14539 35392 14614 35398
rect 14539 35358 14607 35392
rect 14648 35364 14724 35398
rect 14641 35358 14724 35364
rect 14539 35326 14724 35358
rect 14539 35324 14614 35326
rect 14539 35290 14607 35324
rect 14648 35292 14724 35326
rect 14641 35290 14724 35292
rect 14539 35256 14724 35290
rect 14539 35222 14607 35256
rect 14641 35254 14724 35256
rect 14539 35220 14614 35222
rect 14648 35220 14724 35254
rect 14539 35188 14724 35220
rect 14539 35154 14607 35188
rect 14641 35182 14724 35188
rect 14539 35148 14614 35154
rect 14648 35148 14724 35182
rect 14539 35120 14724 35148
rect 14539 35086 14607 35120
rect 14641 35110 14724 35120
rect 14539 35076 14614 35086
rect 14648 35076 14724 35110
rect 14539 35052 14724 35076
rect 14539 35018 14607 35052
rect 14641 35038 14724 35052
rect 14539 35004 14614 35018
rect 14648 35004 14724 35038
rect 14539 34984 14724 35004
rect 14539 34950 14607 34984
rect 14641 34966 14724 34984
rect 14539 34932 14614 34950
rect 14648 34932 14724 34966
rect 14539 34916 14724 34932
rect 14539 34882 14607 34916
rect 14641 34894 14724 34916
rect 14539 34860 14614 34882
rect 14648 34860 14724 34894
rect 14539 34848 14724 34860
rect 14539 34814 14607 34848
rect 14641 34822 14724 34848
rect 14539 34788 14614 34814
rect 14648 34788 14724 34822
rect 14539 34780 14724 34788
rect 14539 34746 14607 34780
rect 14641 34750 14724 34780
rect 14539 34716 14614 34746
rect 14648 34716 14724 34750
rect 14539 34712 14724 34716
rect 14539 34678 14607 34712
rect 14641 34678 14724 34712
rect 14539 34644 14614 34678
rect 14648 34644 14724 34678
rect 14539 34610 14607 34644
rect 14641 34610 14724 34644
rect 14539 34606 14724 34610
rect 14539 34576 14614 34606
rect 14539 34542 14607 34576
rect 14648 34572 14724 34606
rect 14641 34542 14724 34572
rect 14539 34534 14724 34542
rect 14539 34508 14614 34534
rect 14539 34474 14607 34508
rect 14648 34500 14724 34534
rect 14641 34474 14724 34500
rect 14539 34462 14724 34474
rect 14539 34440 14614 34462
rect 14539 34406 14607 34440
rect 14648 34428 14724 34462
rect 14641 34406 14724 34428
rect 14539 34390 14724 34406
rect 14539 34372 14614 34390
rect 14539 34338 14607 34372
rect 14648 34356 14724 34390
rect 14641 34338 14724 34356
rect 14539 34318 14724 34338
rect 14539 34304 14614 34318
rect 14539 34270 14607 34304
rect 14648 34284 14724 34318
rect 14641 34270 14724 34284
rect 14539 34246 14724 34270
rect 14539 34236 14614 34246
rect 14539 34202 14607 34236
rect 14648 34212 14724 34246
rect 14641 34202 14724 34212
rect 14539 34174 14724 34202
rect 14539 34168 14614 34174
rect 14539 34134 14607 34168
rect 14648 34140 14724 34174
rect 14641 34134 14724 34140
rect 14539 34102 14724 34134
rect 14539 34100 14614 34102
rect 14539 34066 14607 34100
rect 14648 34068 14724 34102
rect 14641 34066 14724 34068
rect 14539 34032 14724 34066
rect 14539 33998 14607 34032
rect 14641 34030 14724 34032
rect 14539 33996 14614 33998
rect 14648 33996 14724 34030
rect 14539 33964 14724 33996
rect 14539 33930 14607 33964
rect 14641 33958 14724 33964
rect 14539 33924 14614 33930
rect 14648 33924 14724 33958
rect 14539 33896 14724 33924
rect 14539 33862 14607 33896
rect 14641 33886 14724 33896
rect 14539 33852 14614 33862
rect 14648 33852 14724 33886
rect 14539 33828 14724 33852
rect 14539 33794 14607 33828
rect 14641 33814 14724 33828
rect 14539 33780 14614 33794
rect 14648 33780 14724 33814
rect 14539 33760 14724 33780
rect 14539 33726 14607 33760
rect 14641 33742 14724 33760
rect 14539 33708 14614 33726
rect 14648 33708 14724 33742
rect 14539 33692 14724 33708
rect 14539 33658 14607 33692
rect 14641 33670 14724 33692
rect 14539 33636 14614 33658
rect 14648 33636 14724 33670
rect 14539 33624 14724 33636
rect 14539 33590 14607 33624
rect 14641 33598 14724 33624
rect 14539 33564 14614 33590
rect 14648 33564 14724 33598
rect 14539 33556 14724 33564
rect 14539 33522 14607 33556
rect 14641 33526 14724 33556
rect 14539 33492 14614 33522
rect 14648 33492 14724 33526
rect 14539 33488 14724 33492
rect 14539 33454 14607 33488
rect 14641 33454 14724 33488
rect 14539 33420 14614 33454
rect 14648 33420 14724 33454
rect 14539 33386 14607 33420
rect 14641 33386 14724 33420
rect 14539 33382 14724 33386
rect 14539 33352 14614 33382
rect 14539 33318 14607 33352
rect 14648 33348 14724 33382
rect 14641 33318 14724 33348
rect 14539 33310 14724 33318
rect 14539 33284 14614 33310
rect 14539 33250 14607 33284
rect 14648 33276 14724 33310
rect 14641 33250 14724 33276
rect 14539 33238 14724 33250
rect 14539 33216 14614 33238
rect 14539 33182 14607 33216
rect 14648 33204 14724 33238
rect 14641 33182 14724 33204
rect 14539 33166 14724 33182
rect 14539 33148 14614 33166
rect 14539 33114 14607 33148
rect 14648 33132 14724 33166
rect 14641 33114 14724 33132
rect 14539 33094 14724 33114
rect 14539 33080 14614 33094
rect 14539 33046 14607 33080
rect 14648 33060 14724 33094
rect 14641 33046 14724 33060
rect 14539 33022 14724 33046
rect 14539 33012 14614 33022
rect 14539 32978 14607 33012
rect 14648 32988 14724 33022
rect 14641 32978 14724 32988
rect 14539 32950 14724 32978
rect 14539 32944 14614 32950
rect 14539 32910 14607 32944
rect 14648 32916 14724 32950
rect 14641 32910 14724 32916
rect 14539 32878 14724 32910
rect 14539 32876 14614 32878
rect 14539 32842 14607 32876
rect 14648 32844 14724 32878
rect 14641 32842 14724 32844
rect 14539 32808 14724 32842
rect 14539 32774 14607 32808
rect 14641 32806 14724 32808
rect 14539 32772 14614 32774
rect 14648 32772 14724 32806
rect 14539 32740 14724 32772
rect 14539 32706 14607 32740
rect 14641 32734 14724 32740
rect 14539 32700 14614 32706
rect 14648 32700 14724 32734
rect 14539 32672 14724 32700
rect 14539 32638 14607 32672
rect 14641 32662 14724 32672
rect 14539 32628 14614 32638
rect 14648 32628 14724 32662
rect 14539 32604 14724 32628
rect 14539 32570 14607 32604
rect 14641 32590 14724 32604
rect 14539 32556 14614 32570
rect 14648 32556 14724 32590
rect 14539 32536 14724 32556
rect 14539 32502 14607 32536
rect 14641 32518 14724 32536
rect 14539 32484 14614 32502
rect 14648 32484 14724 32518
rect 14539 32468 14724 32484
rect 14539 32434 14607 32468
rect 14641 32446 14724 32468
rect 14539 32412 14614 32434
rect 14648 32412 14724 32446
rect 14539 32400 14724 32412
rect 14539 32366 14607 32400
rect 14641 32374 14724 32400
rect 14539 32340 14614 32366
rect 14648 32340 14724 32374
rect 14539 32332 14724 32340
rect 14539 32298 14607 32332
rect 14641 32302 14724 32332
rect 14539 32268 14614 32298
rect 14648 32268 14724 32302
rect 14539 32264 14724 32268
rect 14539 32230 14607 32264
rect 14641 32230 14724 32264
rect 14539 32196 14614 32230
rect 14648 32196 14724 32230
rect 14539 32162 14607 32196
rect 14641 32162 14724 32196
rect 14539 32158 14724 32162
rect 14539 32128 14614 32158
rect 14539 32094 14607 32128
rect 14648 32124 14724 32158
rect 14641 32094 14724 32124
rect 14539 32086 14724 32094
rect 14539 32060 14614 32086
rect 14539 32026 14607 32060
rect 14648 32052 14724 32086
rect 14641 32026 14724 32052
rect 14539 32014 14724 32026
rect 14539 31992 14614 32014
rect 14539 31958 14607 31992
rect 14648 31980 14724 32014
rect 14641 31958 14724 31980
rect 14539 31942 14724 31958
rect 14539 31924 14614 31942
rect 14539 31890 14607 31924
rect 14648 31908 14724 31942
rect 14641 31890 14724 31908
rect 14539 31870 14724 31890
rect 14539 31856 14614 31870
rect 14539 31822 14607 31856
rect 14648 31836 14724 31870
rect 14641 31822 14724 31836
rect 14539 31798 14724 31822
rect 14539 31788 14614 31798
rect 14539 31754 14607 31788
rect 14648 31764 14724 31798
rect 14641 31754 14724 31764
rect 14539 31726 14724 31754
rect 14539 31720 14614 31726
rect 14539 31686 14607 31720
rect 14648 31692 14724 31726
rect 14641 31686 14724 31692
rect 14539 31654 14724 31686
rect 14539 31652 14614 31654
rect 14539 31618 14607 31652
rect 14648 31620 14724 31654
rect 14641 31618 14724 31620
rect 14539 31584 14724 31618
rect 14539 31550 14607 31584
rect 14641 31582 14724 31584
rect 14539 31548 14614 31550
rect 14648 31548 14724 31582
rect 14539 31516 14724 31548
rect 14539 31482 14607 31516
rect 14641 31510 14724 31516
rect 14539 31476 14614 31482
rect 14648 31476 14724 31510
rect 14539 31448 14724 31476
rect 14539 31414 14607 31448
rect 14641 31438 14724 31448
rect 14539 31404 14614 31414
rect 14648 31404 14724 31438
rect 14539 31380 14724 31404
rect 14539 31346 14607 31380
rect 14641 31366 14724 31380
rect 14539 31332 14614 31346
rect 14648 31332 14724 31366
rect 14539 31312 14724 31332
rect 14539 31278 14607 31312
rect 14641 31294 14724 31312
rect 14539 31260 14614 31278
rect 14648 31260 14724 31294
rect 14539 31244 14724 31260
rect 14539 31210 14607 31244
rect 14641 31222 14724 31244
rect 14539 31188 14614 31210
rect 14648 31188 14724 31222
rect 14539 31176 14724 31188
rect 14539 31142 14607 31176
rect 14641 31150 14724 31176
rect 14539 31116 14614 31142
rect 14648 31116 14724 31150
rect 14539 31108 14724 31116
rect 14539 31074 14607 31108
rect 14641 31078 14724 31108
rect 14539 31044 14614 31074
rect 14648 31044 14724 31078
rect 14539 31040 14724 31044
rect 14539 31006 14607 31040
rect 14641 31006 14724 31040
rect 14539 30972 14614 31006
rect 14648 30972 14724 31006
rect 14539 30938 14607 30972
rect 14641 30938 14724 30972
rect 14539 30934 14724 30938
rect 14539 30904 14614 30934
rect 14539 30870 14607 30904
rect 14648 30900 14724 30934
rect 14641 30870 14724 30900
rect 14539 30862 14724 30870
rect 14539 30836 14614 30862
rect 14539 30802 14607 30836
rect 14648 30828 14724 30862
rect 14641 30802 14724 30828
rect 14539 30790 14724 30802
rect 14539 30768 14614 30790
rect 14539 30734 14607 30768
rect 14648 30756 14724 30790
rect 14641 30734 14724 30756
rect 14539 30718 14724 30734
rect 14539 30700 14614 30718
rect 14539 30666 14607 30700
rect 14648 30684 14724 30718
rect 14641 30666 14724 30684
rect 14539 30646 14724 30666
rect 14539 30632 14614 30646
rect 14539 30598 14607 30632
rect 14648 30612 14724 30646
rect 14641 30598 14724 30612
rect 14539 30574 14724 30598
rect 14539 30564 14614 30574
rect 14539 30530 14607 30564
rect 14648 30540 14724 30574
rect 14641 30530 14724 30540
rect 14539 30502 14724 30530
rect 14539 30496 14614 30502
rect 14539 30462 14607 30496
rect 14648 30468 14724 30502
rect 14641 30462 14724 30468
rect 14539 30430 14724 30462
rect 14539 30428 14614 30430
rect 14539 30394 14607 30428
rect 14648 30396 14724 30430
rect 14641 30394 14724 30396
rect 14539 30360 14724 30394
rect 14539 30326 14607 30360
rect 14641 30358 14724 30360
rect 14539 30324 14614 30326
rect 14648 30324 14724 30358
rect 14539 30292 14724 30324
rect 14539 30258 14607 30292
rect 14641 30286 14724 30292
rect 14539 30252 14614 30258
rect 14648 30252 14724 30286
rect 14539 30224 14724 30252
rect 14539 30190 14607 30224
rect 14641 30214 14724 30224
rect 14539 30180 14614 30190
rect 14648 30180 14724 30214
rect 14539 30156 14724 30180
rect 14539 30122 14607 30156
rect 14641 30142 14724 30156
rect 14539 30108 14614 30122
rect 14648 30108 14724 30142
rect 14539 30088 14724 30108
rect 14539 30054 14607 30088
rect 14641 30070 14724 30088
rect 14539 30036 14614 30054
rect 14648 30036 14724 30070
rect 14539 30020 14724 30036
rect 14539 29986 14607 30020
rect 14641 29998 14724 30020
rect 14539 29964 14614 29986
rect 14648 29964 14724 29998
rect 14539 29952 14724 29964
rect 14539 29918 14607 29952
rect 14641 29926 14724 29952
rect 14539 29892 14614 29918
rect 14648 29892 14724 29926
rect 14539 29884 14724 29892
rect 14539 29850 14607 29884
rect 14641 29854 14724 29884
rect 14539 29820 14614 29850
rect 14648 29820 14724 29854
rect 14539 29816 14724 29820
rect 14539 29782 14607 29816
rect 14641 29782 14724 29816
rect 14539 29748 14614 29782
rect 14648 29748 14724 29782
rect 14539 29714 14607 29748
rect 14641 29714 14724 29748
rect 14539 29710 14724 29714
rect 14539 29680 14614 29710
rect 14539 29646 14607 29680
rect 14648 29676 14724 29710
rect 14641 29646 14724 29676
rect 14539 29638 14724 29646
rect 14539 29612 14614 29638
rect 14539 29578 14607 29612
rect 14648 29604 14724 29638
rect 14641 29578 14724 29604
rect 14539 29566 14724 29578
rect 14539 29544 14614 29566
rect 14539 29510 14607 29544
rect 14648 29532 14724 29566
rect 14641 29510 14724 29532
rect 14539 29494 14724 29510
rect 14539 29476 14614 29494
rect 14539 29442 14607 29476
rect 14648 29460 14724 29494
rect 14641 29442 14724 29460
rect 14539 29422 14724 29442
rect 14539 29408 14614 29422
rect 14539 29374 14607 29408
rect 14648 29388 14724 29422
rect 14641 29374 14724 29388
rect 14539 29350 14724 29374
rect 14539 29340 14614 29350
rect 14539 29306 14607 29340
rect 14648 29316 14724 29350
rect 14641 29306 14724 29316
rect 14539 29278 14724 29306
rect 14539 29272 14614 29278
rect 14539 29238 14607 29272
rect 14648 29244 14724 29278
rect 14641 29238 14724 29244
rect 14539 29206 14724 29238
rect 14539 29204 14614 29206
rect 14539 29170 14607 29204
rect 14648 29172 14724 29206
rect 14641 29170 14724 29172
rect 14539 29136 14724 29170
rect 14539 29102 14607 29136
rect 14641 29134 14724 29136
rect 14539 29100 14614 29102
rect 14648 29100 14724 29134
rect 14539 29068 14724 29100
rect 14539 29034 14607 29068
rect 14641 29062 14724 29068
rect 14539 29028 14614 29034
rect 14648 29028 14724 29062
rect 14539 29000 14724 29028
rect 14539 28966 14607 29000
rect 14641 28990 14724 29000
rect 14539 28956 14614 28966
rect 14648 28956 14724 28990
rect 14539 28932 14724 28956
rect 14539 28898 14607 28932
rect 14641 28918 14724 28932
rect 14539 28884 14614 28898
rect 14648 28884 14724 28918
rect 14539 28864 14724 28884
rect 14539 28830 14607 28864
rect 14641 28846 14724 28864
rect 14539 28812 14614 28830
rect 14648 28812 14724 28846
rect 14539 28796 14724 28812
rect 14539 28762 14607 28796
rect 14641 28774 14724 28796
rect 14539 28740 14614 28762
rect 14648 28740 14724 28774
rect 14539 28728 14724 28740
rect 14539 28694 14607 28728
rect 14641 28702 14724 28728
rect 14539 28668 14614 28694
rect 14648 28668 14724 28702
rect 14539 28660 14724 28668
rect 14539 28626 14607 28660
rect 14641 28630 14724 28660
rect 14539 28596 14614 28626
rect 14648 28596 14724 28630
rect 14539 28592 14724 28596
rect 14539 28558 14607 28592
rect 14641 28558 14724 28592
rect 14539 28524 14614 28558
rect 14648 28524 14724 28558
rect 14539 28490 14607 28524
rect 14641 28490 14724 28524
rect 14539 28486 14724 28490
rect 14539 28456 14614 28486
rect 14539 28422 14607 28456
rect 14648 28452 14724 28486
rect 14641 28422 14724 28452
rect 14539 28414 14724 28422
rect 14539 28388 14614 28414
rect 14539 28354 14607 28388
rect 14648 28380 14724 28414
rect 14641 28354 14724 28380
rect 14539 28342 14724 28354
rect 14539 28320 14614 28342
rect 14539 28286 14607 28320
rect 14648 28308 14724 28342
rect 14641 28286 14724 28308
rect 14539 28270 14724 28286
rect 14539 28252 14614 28270
rect 14539 28218 14607 28252
rect 14648 28236 14724 28270
rect 14641 28218 14724 28236
rect 14539 28198 14724 28218
rect 14539 28184 14614 28198
rect 14539 28150 14607 28184
rect 14648 28164 14724 28198
rect 14641 28150 14724 28164
rect 14539 28126 14724 28150
rect 14539 28116 14614 28126
rect 14539 28082 14607 28116
rect 14648 28092 14724 28126
rect 14641 28082 14724 28092
rect 14539 28054 14724 28082
rect 14539 28048 14614 28054
rect 14539 28014 14607 28048
rect 14648 28020 14724 28054
rect 14641 28014 14724 28020
rect 14539 27982 14724 28014
rect 14539 27980 14614 27982
rect 14539 27946 14607 27980
rect 14648 27948 14724 27982
rect 14641 27946 14724 27948
rect 14539 27912 14724 27946
rect 14539 27878 14607 27912
rect 14641 27910 14724 27912
rect 14539 27876 14614 27878
rect 14648 27876 14724 27910
rect 14539 27844 14724 27876
rect 14539 27810 14607 27844
rect 14641 27838 14724 27844
rect 14539 27804 14614 27810
rect 14648 27804 14724 27838
rect 14539 27776 14724 27804
rect 14539 27742 14607 27776
rect 14641 27766 14724 27776
rect 14539 27732 14614 27742
rect 14648 27732 14724 27766
rect 14539 27708 14724 27732
rect 14539 27674 14607 27708
rect 14641 27694 14724 27708
rect 14539 27660 14614 27674
rect 14648 27660 14724 27694
rect 14539 27640 14724 27660
rect 14539 27606 14607 27640
rect 14641 27622 14724 27640
rect 14539 27588 14614 27606
rect 14648 27588 14724 27622
rect 14539 27572 14724 27588
rect 14539 27538 14607 27572
rect 14641 27550 14724 27572
rect 14539 27516 14614 27538
rect 14648 27516 14724 27550
rect 14539 27504 14724 27516
rect 14539 27470 14607 27504
rect 14641 27478 14724 27504
rect 14539 27444 14614 27470
rect 14648 27444 14724 27478
rect 14539 27436 14724 27444
rect 14539 27402 14607 27436
rect 14641 27406 14724 27436
rect 14539 27372 14614 27402
rect 14648 27372 14724 27406
rect 14539 27368 14724 27372
rect 14539 27334 14607 27368
rect 14641 27334 14724 27368
rect 14539 27300 14614 27334
rect 14648 27300 14724 27334
rect 14539 27266 14607 27300
rect 14641 27266 14724 27300
rect 14539 27262 14724 27266
rect 14539 27232 14614 27262
rect 14539 27198 14607 27232
rect 14648 27228 14724 27262
rect 14641 27198 14724 27228
rect 14539 27190 14724 27198
rect 14539 27164 14614 27190
rect 14539 27130 14607 27164
rect 14648 27156 14724 27190
rect 14641 27130 14724 27156
rect 14539 27118 14724 27130
rect 14539 27096 14614 27118
rect 14539 27062 14607 27096
rect 14648 27084 14724 27118
rect 14641 27062 14724 27084
rect 14539 27046 14724 27062
rect 14539 27028 14614 27046
rect 14539 26994 14607 27028
rect 14648 27012 14724 27046
rect 14641 26994 14724 27012
rect 14539 26974 14724 26994
rect 14539 26960 14614 26974
rect 14539 26926 14607 26960
rect 14648 26940 14724 26974
rect 14641 26926 14724 26940
rect 14539 26902 14724 26926
rect 14539 26892 14614 26902
rect 14539 26858 14607 26892
rect 14648 26868 14724 26902
rect 14641 26858 14724 26868
rect 14539 26830 14724 26858
rect 14539 26824 14614 26830
rect 14539 26790 14607 26824
rect 14648 26796 14724 26830
rect 14641 26790 14724 26796
rect 14539 26758 14724 26790
rect 14539 26756 14614 26758
rect 14539 26722 14607 26756
rect 14648 26724 14724 26758
rect 14641 26722 14724 26724
rect 14539 26688 14724 26722
rect 14539 26654 14607 26688
rect 14641 26686 14724 26688
rect 14539 26652 14614 26654
rect 14648 26652 14724 26686
rect 14539 26620 14724 26652
rect 14539 26586 14607 26620
rect 14641 26614 14724 26620
rect 14539 26580 14614 26586
rect 14648 26580 14724 26614
rect 14539 26552 14724 26580
rect 14539 26518 14607 26552
rect 14641 26542 14724 26552
rect 14539 26508 14614 26518
rect 14648 26508 14724 26542
rect 14539 26484 14724 26508
rect 14539 26450 14607 26484
rect 14641 26470 14724 26484
rect 14539 26436 14614 26450
rect 14648 26436 14724 26470
rect 14539 26416 14724 26436
rect 14539 26382 14607 26416
rect 14641 26398 14724 26416
rect 14539 26364 14614 26382
rect 14648 26364 14724 26398
rect 14539 26348 14724 26364
rect 14539 26314 14607 26348
rect 14641 26326 14724 26348
rect 14539 26292 14614 26314
rect 14648 26292 14724 26326
rect 14539 26280 14724 26292
rect 14539 26246 14607 26280
rect 14641 26254 14724 26280
rect 14539 26220 14614 26246
rect 14648 26220 14724 26254
rect 14539 26212 14724 26220
rect 14539 26178 14607 26212
rect 14641 26182 14724 26212
rect 14539 26148 14614 26178
rect 14648 26148 14724 26182
rect 14539 26144 14724 26148
rect 14539 26110 14607 26144
rect 14641 26110 14724 26144
rect 14539 26076 14614 26110
rect 14648 26076 14724 26110
rect 14539 26042 14607 26076
rect 14641 26042 14724 26076
rect 14539 26038 14724 26042
rect 14539 26008 14614 26038
rect 14539 25974 14607 26008
rect 14648 26004 14724 26038
rect 14641 25974 14724 26004
rect 14539 25966 14724 25974
rect 14539 25940 14614 25966
rect 14539 25906 14607 25940
rect 14648 25932 14724 25966
rect 14641 25906 14724 25932
rect 14539 25894 14724 25906
rect 14539 25872 14614 25894
rect 14539 25838 14607 25872
rect 14648 25860 14724 25894
rect 14641 25838 14724 25860
rect 14539 25822 14724 25838
rect 14539 25804 14614 25822
rect 14539 25770 14607 25804
rect 14648 25788 14724 25822
rect 14641 25770 14724 25788
rect 14539 25750 14724 25770
rect 14539 25736 14614 25750
rect 14539 25702 14607 25736
rect 14648 25716 14724 25750
rect 14641 25702 14724 25716
rect 14539 25678 14724 25702
rect 14539 25668 14614 25678
rect 14539 25634 14607 25668
rect 14648 25644 14724 25678
rect 14641 25634 14724 25644
rect 14539 25606 14724 25634
rect 14539 25600 14614 25606
rect 14539 25566 14607 25600
rect 14648 25572 14724 25606
rect 14641 25566 14724 25572
rect 14539 25534 14724 25566
rect 14539 25532 14614 25534
rect 14539 25498 14607 25532
rect 14648 25500 14724 25534
rect 14641 25498 14724 25500
rect 14539 25464 14724 25498
rect 14539 25430 14607 25464
rect 14641 25462 14724 25464
rect 14539 25428 14614 25430
rect 14648 25428 14724 25462
rect 14539 25396 14724 25428
rect 14539 25362 14607 25396
rect 14641 25390 14724 25396
rect 14539 25356 14614 25362
rect 14648 25356 14724 25390
rect 14539 25328 14724 25356
rect 14539 25294 14607 25328
rect 14641 25318 14724 25328
rect 14539 25284 14614 25294
rect 14648 25284 14724 25318
rect 14539 25260 14724 25284
rect 14539 25226 14607 25260
rect 14641 25246 14724 25260
rect 14539 25212 14614 25226
rect 14648 25212 14724 25246
rect 14539 25192 14724 25212
rect 14539 25158 14607 25192
rect 14641 25174 14724 25192
rect 14539 25140 14614 25158
rect 14648 25140 14724 25174
rect 14539 25124 14724 25140
rect 14539 25090 14607 25124
rect 14641 25102 14724 25124
rect 14539 25068 14614 25090
rect 14648 25068 14724 25102
rect 14539 25056 14724 25068
rect 14539 25022 14607 25056
rect 14641 25030 14724 25056
rect 14539 24996 14614 25022
rect 14648 24996 14724 25030
rect 14539 24988 14724 24996
rect 14539 24954 14607 24988
rect 14641 24958 14724 24988
rect 14539 24924 14614 24954
rect 14648 24924 14724 24958
rect 14539 24920 14724 24924
rect 14539 24886 14607 24920
rect 14641 24886 14724 24920
rect 14539 24852 14614 24886
rect 14648 24852 14724 24886
rect 14539 24818 14607 24852
rect 14641 24818 14724 24852
rect 14539 24814 14724 24818
rect 14539 24784 14614 24814
rect 14539 24750 14607 24784
rect 14648 24780 14724 24814
rect 14641 24750 14724 24780
rect 14539 24742 14724 24750
rect 14539 24716 14614 24742
rect 14539 24682 14607 24716
rect 14648 24708 14724 24742
rect 14641 24682 14724 24708
rect 14539 24670 14724 24682
rect 14539 24648 14614 24670
rect 14539 24614 14607 24648
rect 14648 24636 14724 24670
rect 14641 24614 14724 24636
rect 14539 24598 14724 24614
rect 14539 24580 14614 24598
rect 14539 24546 14607 24580
rect 14648 24564 14724 24598
rect 14641 24546 14724 24564
rect 14539 24526 14724 24546
rect 14539 24512 14614 24526
rect 14539 24478 14607 24512
rect 14648 24492 14724 24526
rect 14641 24478 14724 24492
rect 14539 24454 14724 24478
rect 14539 24444 14614 24454
rect 14539 24410 14607 24444
rect 14648 24420 14724 24454
rect 14641 24410 14724 24420
rect 14539 24382 14724 24410
rect 14539 24376 14614 24382
rect 14539 24342 14607 24376
rect 14648 24348 14724 24382
rect 14641 24342 14724 24348
rect 14539 24310 14724 24342
rect 14539 24308 14614 24310
rect 14539 24274 14607 24308
rect 14648 24276 14724 24310
rect 14641 24274 14724 24276
rect 14539 24240 14724 24274
rect 14539 24206 14607 24240
rect 14641 24238 14724 24240
rect 14539 24204 14614 24206
rect 14648 24204 14724 24238
rect 14539 24172 14724 24204
rect 14539 24138 14607 24172
rect 14641 24166 14724 24172
rect 14539 24132 14614 24138
rect 14648 24132 14724 24166
rect 14539 24104 14724 24132
rect 14539 24070 14607 24104
rect 14641 24094 14724 24104
rect 14539 24060 14614 24070
rect 14648 24060 14724 24094
rect 14539 24036 14724 24060
rect 14539 24002 14607 24036
rect 14641 24022 14724 24036
rect 14539 23988 14614 24002
rect 14648 23988 14724 24022
rect 14539 23968 14724 23988
rect 14539 23934 14607 23968
rect 14641 23950 14724 23968
rect 14539 23916 14614 23934
rect 14648 23916 14724 23950
rect 14539 23900 14724 23916
rect 14539 23866 14607 23900
rect 14641 23878 14724 23900
rect 14539 23844 14614 23866
rect 14648 23844 14724 23878
rect 14539 23832 14724 23844
rect 14539 23798 14607 23832
rect 14641 23806 14724 23832
rect 14539 23772 14614 23798
rect 14648 23772 14724 23806
rect 14539 23764 14724 23772
rect 14539 23730 14607 23764
rect 14641 23734 14724 23764
rect 14539 23700 14614 23730
rect 14648 23700 14724 23734
rect 14539 23696 14724 23700
rect 14539 23662 14607 23696
rect 14641 23662 14724 23696
rect 14539 23628 14614 23662
rect 14648 23628 14724 23662
rect 14539 23594 14607 23628
rect 14641 23594 14724 23628
rect 14539 23590 14724 23594
rect 14539 23560 14614 23590
rect 14539 23526 14607 23560
rect 14648 23556 14724 23590
rect 14641 23526 14724 23556
rect 14539 23518 14724 23526
rect 14539 23492 14614 23518
rect 14539 23458 14607 23492
rect 14648 23484 14724 23518
rect 14641 23458 14724 23484
rect 14539 23446 14724 23458
rect 14539 23424 14614 23446
rect 14539 23390 14607 23424
rect 14648 23412 14724 23446
rect 14641 23390 14724 23412
rect 14539 23374 14724 23390
rect 14539 23356 14614 23374
rect 14539 23322 14607 23356
rect 14648 23340 14724 23374
rect 14641 23322 14724 23340
rect 14539 23302 14724 23322
rect 14539 23288 14614 23302
rect 14539 23254 14607 23288
rect 14648 23268 14724 23302
rect 14641 23254 14724 23268
rect 14539 23230 14724 23254
rect 14539 23220 14614 23230
rect 14539 23186 14607 23220
rect 14648 23196 14724 23230
rect 14641 23186 14724 23196
rect 14539 23158 14724 23186
rect 14539 23152 14614 23158
rect 14539 23118 14607 23152
rect 14648 23124 14724 23158
rect 14641 23118 14724 23124
rect 14539 23086 14724 23118
rect 14539 23084 14614 23086
rect 14539 23050 14607 23084
rect 14648 23052 14724 23086
rect 14641 23050 14724 23052
rect 14539 23016 14724 23050
rect 14539 22982 14607 23016
rect 14641 23014 14724 23016
rect 14539 22980 14614 22982
rect 14648 22980 14724 23014
rect 14539 22948 14724 22980
rect 14539 22914 14607 22948
rect 14641 22942 14724 22948
rect 14539 22908 14614 22914
rect 14648 22908 14724 22942
rect 14539 22880 14724 22908
rect 14539 22846 14607 22880
rect 14641 22870 14724 22880
rect 14539 22836 14614 22846
rect 14648 22836 14724 22870
rect 14539 22812 14724 22836
rect 14539 22778 14607 22812
rect 14641 22798 14724 22812
rect 14539 22764 14614 22778
rect 14648 22764 14724 22798
rect 14539 22744 14724 22764
rect 14539 22710 14607 22744
rect 14641 22726 14724 22744
rect 14539 22692 14614 22710
rect 14648 22692 14724 22726
rect 14539 22676 14724 22692
rect 14539 22642 14607 22676
rect 14641 22654 14724 22676
rect 14539 22620 14614 22642
rect 14648 22620 14724 22654
rect 14539 22608 14724 22620
rect 14539 22574 14607 22608
rect 14641 22582 14724 22608
rect 14539 22548 14614 22574
rect 14648 22548 14724 22582
rect 14539 22540 14724 22548
rect 14539 22506 14607 22540
rect 14641 22510 14724 22540
rect 14539 22476 14614 22506
rect 14648 22476 14724 22510
rect 14539 22472 14724 22476
rect 14539 22438 14607 22472
rect 14641 22438 14724 22472
rect 14539 22404 14614 22438
rect 14648 22404 14724 22438
rect 14539 22370 14607 22404
rect 14641 22370 14724 22404
rect 14539 22366 14724 22370
rect 14539 22336 14614 22366
rect 14539 22302 14607 22336
rect 14648 22332 14724 22366
rect 14641 22302 14724 22332
rect 14539 22294 14724 22302
rect 14539 22268 14614 22294
rect 14539 22234 14607 22268
rect 14648 22260 14724 22294
rect 14641 22234 14724 22260
rect 14539 22222 14724 22234
rect 14539 22200 14614 22222
rect 14539 22166 14607 22200
rect 14648 22188 14724 22222
rect 14641 22166 14724 22188
rect 14539 22150 14724 22166
rect 14539 22132 14614 22150
rect 14539 22098 14607 22132
rect 14648 22116 14724 22150
rect 14641 22098 14724 22116
rect 14539 22078 14724 22098
rect 14539 22064 14614 22078
rect 14539 22030 14607 22064
rect 14648 22044 14724 22078
rect 14641 22030 14724 22044
rect 14539 22006 14724 22030
rect 14539 21996 14614 22006
rect 14539 21962 14607 21996
rect 14648 21972 14724 22006
rect 14641 21962 14724 21972
rect 14539 21934 14724 21962
rect 14539 21928 14614 21934
rect 14539 21894 14607 21928
rect 14648 21900 14724 21934
rect 14641 21894 14724 21900
rect 14539 21862 14724 21894
rect 14539 21860 14614 21862
rect 14539 21826 14607 21860
rect 14648 21828 14724 21862
rect 14641 21826 14724 21828
rect 14539 21792 14724 21826
rect 14539 21758 14607 21792
rect 14641 21790 14724 21792
rect 14539 21756 14614 21758
rect 14648 21756 14724 21790
rect 14539 21724 14724 21756
rect 14539 21690 14607 21724
rect 14641 21718 14724 21724
rect 14539 21684 14614 21690
rect 14648 21684 14724 21718
rect 14539 21656 14724 21684
rect 14539 21622 14607 21656
rect 14641 21646 14724 21656
rect 14539 21612 14614 21622
rect 14648 21612 14724 21646
rect 14539 21588 14724 21612
rect 14539 21554 14607 21588
rect 14641 21574 14724 21588
rect 14539 21540 14614 21554
rect 14648 21540 14724 21574
rect 14539 21520 14724 21540
rect 14539 21486 14607 21520
rect 14641 21502 14724 21520
rect 14539 21468 14614 21486
rect 14648 21468 14724 21502
rect 14539 21452 14724 21468
rect 14539 21418 14607 21452
rect 14641 21430 14724 21452
rect 14539 21396 14614 21418
rect 14648 21396 14724 21430
rect 14539 21384 14724 21396
rect 14539 21350 14607 21384
rect 14641 21358 14724 21384
rect 14539 21324 14614 21350
rect 14648 21324 14724 21358
rect 14539 21316 14724 21324
rect 14539 21282 14607 21316
rect 14641 21286 14724 21316
rect 14539 21252 14614 21282
rect 14648 21252 14724 21286
rect 14539 21248 14724 21252
rect 14539 21214 14607 21248
rect 14641 21214 14724 21248
rect 14539 21180 14614 21214
rect 14648 21180 14724 21214
rect 14539 21146 14607 21180
rect 14641 21146 14724 21180
rect 14539 21142 14724 21146
rect 14539 21112 14614 21142
rect 14539 21078 14607 21112
rect 14648 21108 14724 21142
rect 14641 21078 14724 21108
rect 14539 21070 14724 21078
rect 14539 21044 14614 21070
rect 14539 21010 14607 21044
rect 14648 21036 14724 21070
rect 14641 21010 14724 21036
rect 14539 20998 14724 21010
rect 14539 20976 14614 20998
rect 14539 20942 14607 20976
rect 14648 20964 14724 20998
rect 14641 20942 14724 20964
rect 14539 20926 14724 20942
rect 14539 20908 14614 20926
rect 14539 20874 14607 20908
rect 14648 20892 14724 20926
rect 14641 20874 14724 20892
rect 14539 20854 14724 20874
rect 14539 20840 14614 20854
rect 14539 20806 14607 20840
rect 14648 20820 14724 20854
rect 14641 20806 14724 20820
rect 14539 20782 14724 20806
rect 14539 20772 14614 20782
rect 14539 20738 14607 20772
rect 14648 20748 14724 20782
rect 14641 20738 14724 20748
rect 14539 20710 14724 20738
rect 14539 20704 14614 20710
rect 14539 20670 14607 20704
rect 14648 20676 14724 20710
rect 14641 20670 14724 20676
rect 14539 20638 14724 20670
rect 14539 20636 14614 20638
rect 14539 20602 14607 20636
rect 14648 20604 14724 20638
rect 14641 20602 14724 20604
rect 14539 20568 14724 20602
rect 14539 20534 14607 20568
rect 14641 20566 14724 20568
rect 14539 20532 14614 20534
rect 14648 20532 14724 20566
rect 14539 20500 14724 20532
rect 14539 20466 14607 20500
rect 14641 20494 14724 20500
rect 14539 20460 14614 20466
rect 14648 20460 14724 20494
rect 14539 20432 14724 20460
rect 14539 20398 14607 20432
rect 14641 20422 14724 20432
rect 14539 20388 14614 20398
rect 14648 20388 14724 20422
rect 14539 20364 14724 20388
rect 14539 20330 14607 20364
rect 14641 20350 14724 20364
rect 14539 20316 14614 20330
rect 14648 20316 14724 20350
rect 14539 20296 14724 20316
rect 14539 20262 14607 20296
rect 14641 20278 14724 20296
rect 14539 20244 14614 20262
rect 14648 20244 14724 20278
rect 14539 20228 14724 20244
rect 14539 20194 14607 20228
rect 14641 20206 14724 20228
rect 14539 20172 14614 20194
rect 14648 20172 14724 20206
rect 14539 20160 14724 20172
rect 14539 20126 14607 20160
rect 14641 20134 14724 20160
rect 14539 20100 14614 20126
rect 14648 20100 14724 20134
rect 14539 20092 14724 20100
rect 14539 20058 14607 20092
rect 14641 20062 14724 20092
rect 14539 20028 14614 20058
rect 14648 20028 14724 20062
rect 14539 20024 14724 20028
rect 14539 19990 14607 20024
rect 14641 19990 14724 20024
rect 14539 19956 14614 19990
rect 14648 19956 14724 19990
rect 14539 19922 14607 19956
rect 14641 19922 14724 19956
rect 14539 19918 14724 19922
rect 14539 19888 14614 19918
rect 14539 19854 14607 19888
rect 14648 19884 14724 19918
rect 14641 19854 14724 19884
rect 14539 19846 14724 19854
rect 14539 19820 14614 19846
rect 14539 19786 14607 19820
rect 14648 19812 14724 19846
rect 14641 19786 14724 19812
rect 14539 19774 14724 19786
rect 14539 19752 14614 19774
rect 14539 19718 14607 19752
rect 14648 19740 14724 19774
rect 14641 19718 14724 19740
rect 14539 19702 14724 19718
rect 14539 19684 14614 19702
rect 14539 19650 14607 19684
rect 14648 19668 14724 19702
rect 14641 19650 14724 19668
rect 14539 19630 14724 19650
rect 14539 19616 14614 19630
rect 14539 19582 14607 19616
rect 14648 19596 14724 19630
rect 14641 19582 14724 19596
rect 14539 19558 14724 19582
rect 14539 19548 14614 19558
rect 14539 19514 14607 19548
rect 14648 19524 14724 19558
rect 14641 19514 14724 19524
rect 14539 19486 14724 19514
rect 14539 19480 14614 19486
rect 14539 19446 14607 19480
rect 14648 19452 14724 19486
rect 14641 19446 14724 19452
rect 14539 19414 14724 19446
rect 14539 19412 14614 19414
rect 14539 19378 14607 19412
rect 14648 19380 14724 19414
rect 14641 19378 14724 19380
rect 14539 19344 14724 19378
rect 14539 19310 14607 19344
rect 14641 19342 14724 19344
rect 14539 19308 14614 19310
rect 14648 19308 14724 19342
rect 14539 19276 14724 19308
rect 14539 19242 14607 19276
rect 14641 19270 14724 19276
rect 14539 19236 14614 19242
rect 14648 19236 14724 19270
rect 14539 19208 14724 19236
rect 14539 19174 14607 19208
rect 14641 19198 14724 19208
rect 14539 19164 14614 19174
rect 14648 19164 14724 19198
rect 14539 19140 14724 19164
rect 14539 19106 14607 19140
rect 14641 19126 14724 19140
rect 14539 19092 14614 19106
rect 14648 19092 14724 19126
rect 14539 19072 14724 19092
rect 14539 19038 14607 19072
rect 14641 19054 14724 19072
rect 14539 19020 14614 19038
rect 14648 19020 14724 19054
rect 14539 19004 14724 19020
rect 14539 18970 14607 19004
rect 14641 18982 14724 19004
rect 14539 18948 14614 18970
rect 14648 18948 14724 18982
rect 14539 18936 14724 18948
rect 14539 18902 14607 18936
rect 14641 18910 14724 18936
rect 14539 18876 14614 18902
rect 14648 18876 14724 18910
rect 14539 18868 14724 18876
rect 14539 18834 14607 18868
rect 14641 18838 14724 18868
rect 14539 18804 14614 18834
rect 14648 18804 14724 18838
rect 14539 18800 14724 18804
rect 14539 18766 14607 18800
rect 14641 18766 14724 18800
rect 14539 18732 14614 18766
rect 14648 18732 14724 18766
rect 14539 18698 14607 18732
rect 14641 18698 14724 18732
rect 14539 18694 14724 18698
rect 14539 18664 14614 18694
rect 14539 18630 14607 18664
rect 14648 18660 14724 18694
rect 14641 18630 14724 18660
rect 14539 18622 14724 18630
rect 14539 18596 14614 18622
rect 14539 18562 14607 18596
rect 14648 18588 14724 18622
rect 14641 18562 14724 18588
rect 14539 18550 14724 18562
rect 14539 18528 14614 18550
rect 14539 18494 14607 18528
rect 14648 18516 14724 18550
rect 14641 18494 14724 18516
rect 14539 18478 14724 18494
rect 14539 18460 14614 18478
rect 14539 18426 14607 18460
rect 14648 18444 14724 18478
rect 14641 18426 14724 18444
rect 14539 18406 14724 18426
rect 14539 18392 14614 18406
rect 14539 18358 14607 18392
rect 14648 18372 14724 18406
rect 14641 18358 14724 18372
rect 14539 18334 14724 18358
rect 14539 18324 14614 18334
rect 14539 18290 14607 18324
rect 14648 18300 14724 18334
rect 14641 18290 14724 18300
rect 14539 18262 14724 18290
rect 14539 18256 14614 18262
rect 14539 18222 14607 18256
rect 14648 18228 14724 18262
rect 14641 18222 14724 18228
rect 14539 18190 14724 18222
rect 14539 18188 14614 18190
rect 14539 18154 14607 18188
rect 14648 18156 14724 18190
rect 14641 18154 14724 18156
rect 14539 18120 14724 18154
rect 14539 18086 14607 18120
rect 14641 18118 14724 18120
rect 14539 18084 14614 18086
rect 14648 18084 14724 18118
rect 14539 18052 14724 18084
rect 14539 18018 14607 18052
rect 14641 18046 14724 18052
rect 14539 18012 14614 18018
rect 14648 18012 14724 18046
rect 14539 17984 14724 18012
rect 14539 17950 14607 17984
rect 14641 17974 14724 17984
rect 14539 17940 14614 17950
rect 14648 17940 14724 17974
rect 14539 17916 14724 17940
rect 14539 17882 14607 17916
rect 14641 17902 14724 17916
rect 14539 17868 14614 17882
rect 14648 17868 14724 17902
rect 14539 17848 14724 17868
rect 14539 17814 14607 17848
rect 14641 17830 14724 17848
rect 14539 17796 14614 17814
rect 14648 17796 14724 17830
rect 14539 17780 14724 17796
rect 14539 17746 14607 17780
rect 14641 17758 14724 17780
rect 14539 17724 14614 17746
rect 14648 17724 14724 17758
rect 14539 17712 14724 17724
rect 14539 17678 14607 17712
rect 14641 17686 14724 17712
rect 14539 17652 14614 17678
rect 14648 17652 14724 17686
rect 14539 17644 14724 17652
rect 14539 17610 14607 17644
rect 14641 17614 14724 17644
rect 14539 17580 14614 17610
rect 14648 17580 14724 17614
rect 14539 17576 14724 17580
rect 14539 17542 14607 17576
rect 14641 17542 14724 17576
rect 14539 17508 14614 17542
rect 14648 17508 14724 17542
rect 14539 17474 14607 17508
rect 14641 17474 14724 17508
rect 14539 17470 14724 17474
rect 14539 17440 14614 17470
rect 14539 17406 14607 17440
rect 14648 17436 14724 17470
rect 14641 17406 14724 17436
rect 14539 17398 14724 17406
rect 14539 17372 14614 17398
rect 14539 17338 14607 17372
rect 14648 17364 14724 17398
rect 14641 17338 14724 17364
rect 14539 17326 14724 17338
rect 14539 17304 14614 17326
rect 14539 17270 14607 17304
rect 14648 17292 14724 17326
rect 14641 17270 14724 17292
rect 14539 17254 14724 17270
rect 14539 17236 14614 17254
rect 14539 17202 14607 17236
rect 14648 17220 14724 17254
rect 14641 17202 14724 17220
rect 14539 17182 14724 17202
rect 14539 17168 14614 17182
rect 14539 17134 14607 17168
rect 14648 17148 14724 17182
rect 14641 17134 14724 17148
rect 14539 17110 14724 17134
rect 14539 17100 14614 17110
rect 14539 17066 14607 17100
rect 14648 17076 14724 17110
rect 14641 17066 14724 17076
rect 14539 17038 14724 17066
rect 14539 17032 14614 17038
rect 14539 16998 14607 17032
rect 14648 17004 14724 17038
rect 14641 16998 14724 17004
rect 14539 16966 14724 16998
rect 14539 16964 14614 16966
rect 14539 16930 14607 16964
rect 14648 16932 14724 16966
rect 14641 16930 14724 16932
rect 14539 16896 14724 16930
rect 14539 16862 14607 16896
rect 14641 16894 14724 16896
rect 14539 16860 14614 16862
rect 14648 16860 14724 16894
rect 14539 16828 14724 16860
rect 14539 16794 14607 16828
rect 14641 16822 14724 16828
rect 14539 16788 14614 16794
rect 14648 16788 14724 16822
rect 14539 16760 14724 16788
rect 14539 16726 14607 16760
rect 14641 16750 14724 16760
rect 14539 16716 14614 16726
rect 14648 16716 14724 16750
rect 14539 16692 14724 16716
rect 14539 16658 14607 16692
rect 14641 16678 14724 16692
rect 14539 16644 14614 16658
rect 14648 16644 14724 16678
rect 14539 16624 14724 16644
rect 14539 16590 14607 16624
rect 14641 16606 14724 16624
rect 14539 16572 14614 16590
rect 14648 16572 14724 16606
rect 14539 16556 14724 16572
rect 14539 16522 14607 16556
rect 14641 16534 14724 16556
rect 14539 16500 14614 16522
rect 14648 16500 14724 16534
rect 14539 16488 14724 16500
rect 14539 16454 14607 16488
rect 14641 16462 14724 16488
rect 14539 16428 14614 16454
rect 14648 16428 14724 16462
rect 14539 16420 14724 16428
rect 14539 16386 14607 16420
rect 14641 16390 14724 16420
rect 14539 16356 14614 16386
rect 14648 16356 14724 16390
rect 14539 16352 14724 16356
rect 14539 16318 14607 16352
rect 14641 16318 14724 16352
rect 14539 16284 14614 16318
rect 14648 16284 14724 16318
rect 14539 16250 14607 16284
rect 14641 16250 14724 16284
rect 14539 16246 14724 16250
rect 14539 16216 14614 16246
rect 14539 16182 14607 16216
rect 14648 16212 14724 16246
rect 14641 16182 14724 16212
rect 14539 16174 14724 16182
rect 14539 16148 14614 16174
rect 14539 16114 14607 16148
rect 14648 16140 14724 16174
rect 14641 16114 14724 16140
rect 14539 16102 14724 16114
rect 14539 16080 14614 16102
rect 14539 16046 14607 16080
rect 14648 16068 14724 16102
rect 14641 16046 14724 16068
rect 14539 16030 14724 16046
rect 14539 16012 14614 16030
rect 14539 15978 14607 16012
rect 14648 15996 14724 16030
rect 14641 15978 14724 15996
rect 14539 15958 14724 15978
rect 14539 15944 14614 15958
rect 14539 15910 14607 15944
rect 14648 15924 14724 15958
rect 14641 15910 14724 15924
rect 14539 15886 14724 15910
rect 14539 15876 14614 15886
rect 14539 15842 14607 15876
rect 14648 15852 14724 15886
rect 14641 15842 14724 15852
rect 14539 15814 14724 15842
rect 14539 15808 14614 15814
rect 14539 15774 14607 15808
rect 14648 15780 14724 15814
rect 14641 15774 14724 15780
rect 14539 15742 14724 15774
rect 14539 15740 14614 15742
rect 14539 15706 14607 15740
rect 14648 15708 14724 15742
rect 14641 15706 14724 15708
rect 14539 15672 14724 15706
rect 14539 15638 14607 15672
rect 14641 15670 14724 15672
rect 14539 15636 14614 15638
rect 14648 15636 14724 15670
rect 14539 15604 14724 15636
rect 14539 15570 14607 15604
rect 14641 15598 14724 15604
rect 14539 15564 14614 15570
rect 14648 15564 14724 15598
rect 14539 15536 14724 15564
rect 14539 15502 14607 15536
rect 14641 15526 14724 15536
rect 14539 15492 14614 15502
rect 14648 15492 14724 15526
rect 14539 15468 14724 15492
rect 14539 15434 14607 15468
rect 14641 15454 14724 15468
rect 14539 15420 14614 15434
rect 14648 15420 14724 15454
rect 14539 15400 14724 15420
rect 14539 15366 14607 15400
rect 14641 15382 14724 15400
rect 14539 15348 14614 15366
rect 14648 15348 14724 15382
rect 14539 15332 14724 15348
rect 14539 15298 14607 15332
rect 14641 15310 14724 15332
rect 14539 15276 14614 15298
rect 14648 15276 14724 15310
rect 14539 15264 14724 15276
rect 14539 15230 14607 15264
rect 14641 15238 14724 15264
rect 14539 15204 14614 15230
rect 14648 15204 14724 15238
rect 14539 15196 14724 15204
rect 14539 15162 14607 15196
rect 14641 15166 14724 15196
rect 14539 15132 14614 15162
rect 14648 15132 14724 15166
rect 14539 15128 14724 15132
rect 14539 15094 14607 15128
rect 14641 15094 14724 15128
rect 14539 15060 14614 15094
rect 14648 15060 14724 15094
rect 14539 15026 14607 15060
rect 14641 15026 14724 15060
rect 14539 15022 14724 15026
rect 14539 14992 14614 15022
rect 14539 14958 14607 14992
rect 14648 14988 14724 15022
rect 14641 14958 14724 14988
rect 14539 14950 14724 14958
rect 14539 14924 14614 14950
rect 14539 14890 14607 14924
rect 14648 14916 14724 14950
rect 14641 14890 14724 14916
rect 14539 14878 14724 14890
rect 14539 14856 14614 14878
rect 14539 14822 14607 14856
rect 14648 14844 14724 14878
rect 14641 14822 14724 14844
rect 14539 14806 14724 14822
rect 14539 14788 14614 14806
rect 14539 14754 14607 14788
rect 14648 14772 14724 14806
rect 14641 14754 14724 14772
rect 14539 14734 14724 14754
rect 14539 14720 14614 14734
rect 14539 14686 14607 14720
rect 14648 14700 14724 14734
rect 14641 14686 14724 14700
rect 14539 14662 14724 14686
rect 14539 14652 14614 14662
rect 14539 14618 14607 14652
rect 14648 14628 14724 14662
rect 14641 14618 14724 14628
rect 14539 14590 14724 14618
rect 14539 14584 14614 14590
rect 14539 14550 14607 14584
rect 14648 14556 14724 14590
rect 14641 14550 14724 14556
rect 14539 14518 14724 14550
rect 14539 14516 14614 14518
rect 14539 14482 14607 14516
rect 14648 14484 14724 14518
rect 14641 14482 14724 14484
rect 14539 14448 14724 14482
rect 14539 14414 14607 14448
rect 14641 14446 14724 14448
rect 14539 14412 14614 14414
rect 14648 14412 14724 14446
rect 14539 14380 14724 14412
rect 14539 14346 14607 14380
rect 14641 14374 14724 14380
rect 14539 14340 14614 14346
rect 14648 14340 14724 14374
rect 14539 14312 14724 14340
rect 14539 14278 14607 14312
rect 14641 14302 14724 14312
rect 14539 14268 14614 14278
rect 14648 14268 14724 14302
rect 14539 14244 14724 14268
rect 14539 14210 14607 14244
rect 14641 14230 14724 14244
rect 14539 14196 14614 14210
rect 14648 14196 14724 14230
rect 14539 14176 14724 14196
rect 14539 14142 14607 14176
rect 14641 14158 14724 14176
rect 14539 14124 14614 14142
rect 14648 14124 14724 14158
rect 14539 14108 14724 14124
rect 14539 14074 14607 14108
rect 14641 14086 14724 14108
rect 14539 14052 14614 14074
rect 14648 14052 14724 14086
rect 14539 14040 14724 14052
rect 14539 14006 14607 14040
rect 14641 14014 14724 14040
rect 14539 13980 14614 14006
rect 14648 13980 14724 14014
rect 14539 13972 14724 13980
rect 14539 13938 14607 13972
rect 14641 13942 14724 13972
rect 14539 13908 14614 13938
rect 14648 13908 14724 13942
rect 14539 13904 14724 13908
rect 14539 13870 14607 13904
rect 14641 13870 14724 13904
rect 14539 13836 14614 13870
rect 14648 13836 14724 13870
rect 14539 13802 14607 13836
rect 14641 13802 14724 13836
rect 14539 13798 14724 13802
rect 14539 13768 14614 13798
rect 14539 13734 14607 13768
rect 14648 13764 14724 13798
rect 14641 13734 14724 13764
rect 14539 13726 14724 13734
rect 14539 13700 14614 13726
rect 14539 13666 14607 13700
rect 14648 13692 14724 13726
rect 14641 13666 14724 13692
rect 14539 13654 14724 13666
rect 14539 13632 14614 13654
rect 14539 13598 14607 13632
rect 14648 13620 14724 13654
rect 14641 13598 14724 13620
rect 14539 13582 14724 13598
rect 14539 13564 14614 13582
rect 14539 13530 14607 13564
rect 14648 13548 14724 13582
rect 14641 13530 14724 13548
rect 14539 13510 14724 13530
rect 14539 13496 14614 13510
rect 14539 13462 14607 13496
rect 14648 13476 14724 13510
rect 14641 13462 14724 13476
rect 14539 13438 14724 13462
rect 14539 13428 14614 13438
rect 14539 13394 14607 13428
rect 14648 13404 14724 13438
rect 14641 13394 14724 13404
rect 14539 13366 14724 13394
rect 14539 13360 14614 13366
rect 14539 13326 14607 13360
rect 14648 13332 14724 13366
rect 14641 13326 14724 13332
rect 14539 13294 14724 13326
rect 14539 13292 14614 13294
rect 14539 13258 14607 13292
rect 14648 13260 14724 13294
rect 14641 13258 14724 13260
rect 14539 13224 14724 13258
rect 14539 13190 14607 13224
rect 14641 13222 14724 13224
rect 14539 13188 14614 13190
rect 14648 13188 14724 13222
rect 14539 13156 14724 13188
rect 14539 13122 14607 13156
rect 14641 13150 14724 13156
rect 14539 13116 14614 13122
rect 14648 13116 14724 13150
rect 14539 13088 14724 13116
rect 14539 13054 14607 13088
rect 14641 13078 14724 13088
rect 14539 13044 14614 13054
rect 14648 13044 14724 13078
rect 14539 13020 14724 13044
rect 14539 12986 14607 13020
rect 14641 13006 14724 13020
rect 14539 12972 14614 12986
rect 14648 12972 14724 13006
rect 14539 12952 14724 12972
rect 14539 12918 14607 12952
rect 14641 12934 14724 12952
rect 14539 12900 14614 12918
rect 14648 12900 14724 12934
rect 14539 12884 14724 12900
rect 14539 12850 14607 12884
rect 14641 12862 14724 12884
rect 14539 12828 14614 12850
rect 14648 12828 14724 12862
rect 14539 12816 14724 12828
rect 14539 12782 14607 12816
rect 14641 12790 14724 12816
rect 14539 12756 14614 12782
rect 14648 12756 14724 12790
rect 14539 12748 14724 12756
rect 14539 12714 14607 12748
rect 14641 12718 14724 12748
rect 14539 12684 14614 12714
rect 14648 12684 14724 12718
rect 14539 12680 14724 12684
rect 14539 12646 14607 12680
rect 14641 12646 14724 12680
rect 14539 12612 14614 12646
rect 14648 12612 14724 12646
rect 14539 12578 14607 12612
rect 14641 12578 14724 12612
rect 14539 12574 14724 12578
rect 14539 12544 14614 12574
rect 14539 12510 14607 12544
rect 14648 12540 14724 12574
rect 14641 12510 14724 12540
rect 14539 12502 14724 12510
rect 14539 12476 14614 12502
rect 14539 12442 14607 12476
rect 14648 12468 14724 12502
rect 14641 12442 14724 12468
rect 14539 12430 14724 12442
rect 14539 12408 14614 12430
rect 14539 12374 14607 12408
rect 14648 12396 14724 12430
rect 14641 12374 14724 12396
rect 14539 12358 14724 12374
rect 14539 12340 14614 12358
rect 14539 12306 14607 12340
rect 14648 12324 14724 12358
rect 14641 12306 14724 12324
rect 14539 12286 14724 12306
rect 14539 12272 14614 12286
rect 14539 12238 14607 12272
rect 14648 12252 14724 12286
rect 14641 12238 14724 12252
rect 14539 12214 14724 12238
rect 14539 12204 14614 12214
rect 14539 12170 14607 12204
rect 14648 12180 14724 12214
rect 14641 12170 14724 12180
rect 14539 12142 14724 12170
rect 14539 12136 14614 12142
rect 14539 12102 14607 12136
rect 14648 12108 14724 12142
rect 14641 12102 14724 12108
rect 14539 12070 14724 12102
rect 14539 12068 14614 12070
rect 14539 12034 14607 12068
rect 14648 12036 14724 12070
rect 14641 12034 14724 12036
rect 14539 12000 14724 12034
rect 14539 11966 14607 12000
rect 14641 11998 14724 12000
rect 14539 11964 14614 11966
rect 14648 11964 14724 11998
rect 14539 11932 14724 11964
rect 14539 11898 14607 11932
rect 14641 11926 14724 11932
rect 14539 11892 14614 11898
rect 14648 11892 14724 11926
rect 14539 11864 14724 11892
rect 14539 11830 14607 11864
rect 14641 11854 14724 11864
rect 14539 11820 14614 11830
rect 14648 11820 14724 11854
rect 14539 11796 14724 11820
rect 14539 11762 14607 11796
rect 14641 11782 14724 11796
rect 14539 11748 14614 11762
rect 14648 11748 14724 11782
rect 14539 11728 14724 11748
rect 14539 11694 14607 11728
rect 14641 11710 14724 11728
rect 14539 11676 14614 11694
rect 14648 11676 14724 11710
rect 14539 11660 14724 11676
rect 14539 11626 14607 11660
rect 14641 11638 14724 11660
rect 14539 11604 14614 11626
rect 14648 11604 14724 11638
rect 14539 11592 14724 11604
rect 14539 11558 14607 11592
rect 14641 11566 14724 11592
rect 14539 11532 14614 11558
rect 14648 11532 14724 11566
rect 14539 11524 14724 11532
rect 14539 11490 14607 11524
rect 14641 11494 14724 11524
rect 14539 11460 14614 11490
rect 14648 11460 14724 11494
rect 14539 11456 14724 11460
rect 14539 11422 14607 11456
rect 14641 11422 14724 11456
rect 14539 11388 14614 11422
rect 14648 11388 14724 11422
rect 14539 11354 14607 11388
rect 14641 11354 14724 11388
rect 14539 11350 14724 11354
rect 14539 11320 14614 11350
rect 14539 11286 14607 11320
rect 14648 11316 14724 11350
rect 14641 11286 14724 11316
rect 14539 11278 14724 11286
rect 14539 11252 14614 11278
rect 14539 11218 14607 11252
rect 14648 11244 14724 11278
rect 14641 11218 14724 11244
rect 14539 11206 14724 11218
rect 14539 11184 14614 11206
rect 14539 11150 14607 11184
rect 14648 11172 14724 11206
rect 14641 11150 14724 11172
rect 14539 11134 14724 11150
rect 14539 11116 14614 11134
rect 14539 11082 14607 11116
rect 14648 11100 14724 11134
rect 14641 11082 14724 11100
rect 14539 11062 14724 11082
rect 14539 11048 14614 11062
rect 14539 11014 14607 11048
rect 14648 11028 14724 11062
rect 14641 11014 14724 11028
rect 14539 10990 14724 11014
rect 14539 10980 14614 10990
rect 14539 10946 14607 10980
rect 14648 10956 14724 10990
rect 14641 10946 14724 10956
rect 14539 10918 14724 10946
rect 14539 10912 14614 10918
rect 14539 10878 14607 10912
rect 14648 10884 14724 10918
rect 14641 10878 14724 10884
rect 14539 10846 14724 10878
rect 14539 10844 14614 10846
rect 14539 10810 14607 10844
rect 14648 10812 14724 10846
rect 14641 10810 14724 10812
rect 14539 10776 14724 10810
rect 14539 10742 14607 10776
rect 14641 10774 14724 10776
rect 14539 10740 14614 10742
rect 14648 10740 14724 10774
rect 14539 10708 14724 10740
rect 14539 10674 14607 10708
rect 14641 10702 14724 10708
rect 14539 10668 14614 10674
rect 14648 10668 14724 10702
rect 14539 10640 14724 10668
rect 14539 10606 14607 10640
rect 14641 10630 14724 10640
rect 14539 10596 14614 10606
rect 14648 10596 14724 10630
rect 14539 10572 14724 10596
rect 14539 10538 14607 10572
rect 14641 10558 14724 10572
rect 14539 10524 14614 10538
rect 14648 10524 14724 10558
rect 14539 10504 14724 10524
rect 14539 10470 14607 10504
rect 14641 10486 14724 10504
rect 14539 10452 14614 10470
rect 14648 10452 14724 10486
rect 14539 10436 14724 10452
rect 14539 10402 14607 10436
rect 14641 10414 14724 10436
rect 14539 10380 14614 10402
rect 14648 10380 14724 10414
rect 14539 10368 14724 10380
rect 14539 10334 14607 10368
rect 14641 10342 14724 10368
rect 14539 10308 14614 10334
rect 14648 10308 14724 10342
rect 14539 10300 14724 10308
rect 14539 10266 14607 10300
rect 14641 10270 14724 10300
rect 14539 10236 14614 10266
rect 14648 10236 14724 10270
rect 14539 10232 14724 10236
rect 14539 10198 14607 10232
rect 14641 10198 14724 10232
rect 14539 10164 14614 10198
rect 14648 10164 14724 10198
rect 14539 10130 14607 10164
rect 14641 10130 14724 10164
rect 14539 10126 14724 10130
rect 14539 10096 14614 10126
rect 14539 10062 14607 10096
rect 14648 10092 14724 10126
rect 14641 10062 14724 10092
rect 14539 10054 14724 10062
rect 14539 10028 14614 10054
rect 14539 9994 14607 10028
rect 14648 10020 14724 10054
rect 14641 9994 14724 10020
rect 14539 9982 14724 9994
rect 14539 9960 14614 9982
rect 14539 9926 14607 9960
rect 14648 9948 14724 9982
rect 14641 9926 14724 9948
rect 14539 9910 14724 9926
rect 14539 9892 14614 9910
rect 14539 9858 14607 9892
rect 14648 9876 14724 9910
rect 14641 9858 14724 9876
rect 14539 9838 14724 9858
rect 14539 9824 14614 9838
rect 14539 9790 14607 9824
rect 14648 9804 14724 9838
rect 14641 9790 14724 9804
rect 14539 9766 14724 9790
rect 14539 9756 14614 9766
rect 14539 9722 14607 9756
rect 14648 9732 14724 9766
rect 14641 9722 14724 9732
rect 882 9710 2070 9711
rect 12882 9710 14070 9711
rect 245 9682 320 9697
rect 245 9648 312 9682
rect 354 9663 430 9697
rect 346 9648 430 9663
rect 245 9614 430 9648
rect 245 9580 312 9614
rect 346 9580 430 9614
rect 245 9528 430 9580
rect 14539 9694 14724 9722
rect 14539 9688 14614 9694
rect 14539 9654 14607 9688
rect 14648 9660 14724 9694
rect 14641 9654 14724 9660
rect 14539 9620 14724 9654
rect 14539 9586 14607 9620
rect 14641 9586 14724 9620
rect 14539 9528 14724 9586
rect 245 9452 14724 9528
rect 245 9418 320 9452
rect 354 9451 610 9452
rect 644 9451 2311 9452
rect 2345 9451 2383 9452
rect 2417 9451 2455 9452
rect 2489 9451 2527 9452
rect 2561 9451 2599 9452
rect 2633 9451 2671 9452
rect 2705 9451 2743 9452
rect 2777 9451 2815 9452
rect 2849 9451 2887 9452
rect 2921 9451 2959 9452
rect 2993 9451 3031 9452
rect 3065 9451 3103 9452
rect 3137 9451 3175 9452
rect 3209 9451 3247 9452
rect 3281 9451 3319 9452
rect 3353 9451 3391 9452
rect 3425 9451 3463 9452
rect 3497 9451 3535 9452
rect 3569 9451 3607 9452
rect 3641 9451 3679 9452
rect 3713 9451 3751 9452
rect 3785 9451 3823 9452
rect 3857 9451 3895 9452
rect 3929 9451 3967 9452
rect 4001 9451 4039 9452
rect 4073 9451 4111 9452
rect 4145 9451 4183 9452
rect 4217 9451 4255 9452
rect 4289 9451 4327 9452
rect 4361 9451 4399 9452
rect 4433 9451 4471 9452
rect 4505 9451 4543 9452
rect 4577 9451 4615 9452
rect 4649 9451 4687 9452
rect 4721 9451 4759 9452
rect 4793 9451 4831 9452
rect 4865 9451 4903 9452
rect 4937 9451 4975 9452
rect 5009 9451 5047 9452
rect 5081 9451 5119 9452
rect 5153 9451 5191 9452
rect 5225 9451 5263 9452
rect 5297 9451 5335 9452
rect 5369 9451 5407 9452
rect 5441 9451 5479 9452
rect 5513 9451 5551 9452
rect 5585 9451 5623 9452
rect 5657 9451 5695 9452
rect 5729 9451 5767 9452
rect 5801 9451 5839 9452
rect 5873 9451 5911 9452
rect 5945 9451 5983 9452
rect 6017 9451 6055 9452
rect 6089 9451 6127 9452
rect 6161 9451 6199 9452
rect 6233 9451 6271 9452
rect 6305 9451 6343 9452
rect 6377 9451 6415 9452
rect 6449 9451 6487 9452
rect 6521 9451 6559 9452
rect 6593 9451 6631 9452
rect 6665 9451 6703 9452
rect 6737 9451 6775 9452
rect 6809 9451 6847 9452
rect 6881 9451 6919 9452
rect 6953 9451 6991 9452
rect 7025 9451 7063 9452
rect 7097 9451 7135 9452
rect 7169 9451 7207 9452
rect 7241 9451 7279 9452
rect 7313 9451 7351 9452
rect 7385 9451 7423 9452
rect 7457 9451 7495 9452
rect 7529 9451 7567 9452
rect 7601 9451 7639 9452
rect 7673 9451 7711 9452
rect 7745 9451 7783 9452
rect 7817 9451 7855 9452
rect 7889 9451 7927 9452
rect 7961 9451 7999 9452
rect 8033 9451 8071 9452
rect 8105 9451 8143 9452
rect 8177 9451 8215 9452
rect 8249 9451 8287 9452
rect 8321 9451 8359 9452
rect 8393 9451 8431 9452
rect 8465 9451 8503 9452
rect 8537 9451 8575 9452
rect 8609 9451 8647 9452
rect 8681 9451 8719 9452
rect 8753 9451 8791 9452
rect 8825 9451 8863 9452
rect 8897 9451 8935 9452
rect 8969 9451 9007 9452
rect 9041 9451 9079 9452
rect 9113 9451 9151 9452
rect 9185 9451 9223 9452
rect 9257 9451 9295 9452
rect 9329 9451 9367 9452
rect 9401 9451 9439 9452
rect 9473 9451 9511 9452
rect 9545 9451 9583 9452
rect 9617 9451 9655 9452
rect 9689 9451 9727 9452
rect 9761 9451 9799 9452
rect 9833 9451 9871 9452
rect 9905 9451 9943 9452
rect 9977 9451 10015 9452
rect 10049 9451 10087 9452
rect 10121 9451 10159 9452
rect 10193 9451 10231 9452
rect 10265 9451 10303 9452
rect 10337 9451 10375 9452
rect 10409 9451 10447 9452
rect 10481 9451 10519 9452
rect 10553 9451 10591 9452
rect 10625 9451 10663 9452
rect 10697 9451 10735 9452
rect 10769 9451 10807 9452
rect 10841 9451 10879 9452
rect 10913 9451 10951 9452
rect 10985 9451 11023 9452
rect 11057 9451 11095 9452
rect 11129 9451 11167 9452
rect 11201 9451 11239 9452
rect 11273 9451 11311 9452
rect 11345 9451 11383 9452
rect 11417 9451 11455 9452
rect 11489 9451 11527 9452
rect 11561 9451 11599 9452
rect 11633 9451 11671 9452
rect 11705 9451 11743 9452
rect 11777 9451 11815 9452
rect 11849 9451 11887 9452
rect 11921 9451 11959 9452
rect 11993 9451 12031 9452
rect 12065 9451 12103 9452
rect 12137 9451 12175 9452
rect 12209 9451 12247 9452
rect 12281 9451 12319 9452
rect 12353 9451 12391 9452
rect 12425 9451 12463 9452
rect 12497 9451 12535 9452
rect 12569 9451 12607 9452
rect 12641 9451 14314 9452
rect 354 9418 476 9451
rect 245 9417 476 9418
rect 510 9417 544 9451
rect 578 9418 610 9451
rect 578 9417 612 9418
rect 646 9417 680 9451
rect 714 9417 748 9451
rect 782 9417 816 9451
rect 850 9417 884 9451
rect 918 9417 952 9451
rect 986 9417 1020 9451
rect 1054 9417 1088 9451
rect 1122 9417 1156 9451
rect 1190 9417 1224 9451
rect 1258 9417 1292 9451
rect 1326 9417 1360 9451
rect 1394 9417 1428 9451
rect 1462 9417 1496 9451
rect 1530 9417 1564 9451
rect 1598 9417 1632 9451
rect 1666 9417 1700 9451
rect 1734 9417 1768 9451
rect 1802 9417 1836 9451
rect 1870 9417 1904 9451
rect 1938 9417 1972 9451
rect 2006 9417 2040 9451
rect 2074 9417 2108 9451
rect 2142 9417 2176 9451
rect 2210 9417 2244 9451
rect 2278 9418 2311 9451
rect 2278 9417 2312 9418
rect 2346 9417 2380 9451
rect 2417 9418 2448 9451
rect 2489 9418 2516 9451
rect 2561 9418 2584 9451
rect 2633 9418 2652 9451
rect 2705 9418 2720 9451
rect 2777 9418 2788 9451
rect 2849 9418 2856 9451
rect 2921 9418 2924 9451
rect 2414 9417 2448 9418
rect 2482 9417 2516 9418
rect 2550 9417 2584 9418
rect 2618 9417 2652 9418
rect 2686 9417 2720 9418
rect 2754 9417 2788 9418
rect 2822 9417 2856 9418
rect 2890 9417 2924 9418
rect 2958 9418 2959 9451
rect 3026 9418 3031 9451
rect 3094 9418 3103 9451
rect 3162 9418 3175 9451
rect 3230 9418 3247 9451
rect 3298 9418 3319 9451
rect 3366 9418 3391 9451
rect 3434 9418 3463 9451
rect 3502 9418 3535 9451
rect 2958 9417 2992 9418
rect 3026 9417 3060 9418
rect 3094 9417 3128 9418
rect 3162 9417 3196 9418
rect 3230 9417 3264 9418
rect 3298 9417 3332 9418
rect 3366 9417 3400 9418
rect 3434 9417 3468 9418
rect 3502 9417 3536 9418
rect 3570 9417 3604 9451
rect 3641 9418 3672 9451
rect 3713 9418 3740 9451
rect 3785 9418 3808 9451
rect 3857 9418 3876 9451
rect 3929 9418 3944 9451
rect 4001 9418 4012 9451
rect 4073 9418 4080 9451
rect 4145 9418 4148 9451
rect 3638 9417 3672 9418
rect 3706 9417 3740 9418
rect 3774 9417 3808 9418
rect 3842 9417 3876 9418
rect 3910 9417 3944 9418
rect 3978 9417 4012 9418
rect 4046 9417 4080 9418
rect 4114 9417 4148 9418
rect 4182 9418 4183 9451
rect 4250 9418 4255 9451
rect 4318 9418 4327 9451
rect 4386 9418 4399 9451
rect 4454 9418 4471 9451
rect 4522 9418 4543 9451
rect 4590 9418 4615 9451
rect 4658 9418 4687 9451
rect 4726 9418 4759 9451
rect 4182 9417 4216 9418
rect 4250 9417 4284 9418
rect 4318 9417 4352 9418
rect 4386 9417 4420 9418
rect 4454 9417 4488 9418
rect 4522 9417 4556 9418
rect 4590 9417 4624 9418
rect 4658 9417 4692 9418
rect 4726 9417 4760 9418
rect 4794 9417 4828 9451
rect 4865 9418 4896 9451
rect 4937 9418 4964 9451
rect 5009 9418 5032 9451
rect 5081 9418 5100 9451
rect 5153 9418 5168 9451
rect 5225 9418 5236 9451
rect 5297 9418 5304 9451
rect 5369 9418 5372 9451
rect 4862 9417 4896 9418
rect 4930 9417 4964 9418
rect 4998 9417 5032 9418
rect 5066 9417 5100 9418
rect 5134 9417 5168 9418
rect 5202 9417 5236 9418
rect 5270 9417 5304 9418
rect 5338 9417 5372 9418
rect 5406 9418 5407 9451
rect 5474 9418 5479 9451
rect 5542 9418 5551 9451
rect 5610 9418 5623 9451
rect 5678 9418 5695 9451
rect 5746 9418 5767 9451
rect 5814 9418 5839 9451
rect 5882 9418 5911 9451
rect 5950 9418 5983 9451
rect 5406 9417 5440 9418
rect 5474 9417 5508 9418
rect 5542 9417 5576 9418
rect 5610 9417 5644 9418
rect 5678 9417 5712 9418
rect 5746 9417 5780 9418
rect 5814 9417 5848 9418
rect 5882 9417 5916 9418
rect 5950 9417 5984 9418
rect 6018 9417 6052 9451
rect 6089 9418 6120 9451
rect 6161 9418 6188 9451
rect 6233 9418 6256 9451
rect 6305 9418 6324 9451
rect 6377 9418 6392 9451
rect 6449 9418 6460 9451
rect 6521 9418 6528 9451
rect 6593 9418 6596 9451
rect 6086 9417 6120 9418
rect 6154 9417 6188 9418
rect 6222 9417 6256 9418
rect 6290 9417 6324 9418
rect 6358 9417 6392 9418
rect 6426 9417 6460 9418
rect 6494 9417 6528 9418
rect 6562 9417 6596 9418
rect 6630 9418 6631 9451
rect 6698 9418 6703 9451
rect 6766 9418 6775 9451
rect 6834 9418 6847 9451
rect 6902 9418 6919 9451
rect 6970 9418 6991 9451
rect 7038 9418 7063 9451
rect 7106 9418 7135 9451
rect 7174 9418 7207 9451
rect 6630 9417 6664 9418
rect 6698 9417 6732 9418
rect 6766 9417 6800 9418
rect 6834 9417 6868 9418
rect 6902 9417 6936 9418
rect 6970 9417 7004 9418
rect 7038 9417 7072 9418
rect 7106 9417 7140 9418
rect 7174 9417 7208 9418
rect 7242 9417 7276 9451
rect 7313 9418 7344 9451
rect 7385 9418 7412 9451
rect 7457 9418 7480 9451
rect 7529 9418 7548 9451
rect 7601 9418 7616 9451
rect 7673 9418 7684 9451
rect 7745 9418 7752 9451
rect 7817 9418 7820 9451
rect 7310 9417 7344 9418
rect 7378 9417 7412 9418
rect 7446 9417 7480 9418
rect 7514 9417 7548 9418
rect 7582 9417 7616 9418
rect 7650 9417 7684 9418
rect 7718 9417 7752 9418
rect 7786 9417 7820 9418
rect 7854 9418 7855 9451
rect 7922 9418 7927 9451
rect 7990 9418 7999 9451
rect 8058 9418 8071 9451
rect 8126 9418 8143 9451
rect 8194 9418 8215 9451
rect 8262 9418 8287 9451
rect 8330 9418 8359 9451
rect 8398 9418 8431 9451
rect 7854 9417 7888 9418
rect 7922 9417 7956 9418
rect 7990 9417 8024 9418
rect 8058 9417 8092 9418
rect 8126 9417 8160 9418
rect 8194 9417 8228 9418
rect 8262 9417 8296 9418
rect 8330 9417 8364 9418
rect 8398 9417 8432 9418
rect 8466 9417 8500 9451
rect 8537 9418 8568 9451
rect 8609 9418 8636 9451
rect 8681 9418 8704 9451
rect 8753 9418 8772 9451
rect 8825 9418 8840 9451
rect 8897 9418 8908 9451
rect 8969 9418 8976 9451
rect 9041 9418 9044 9451
rect 8534 9417 8568 9418
rect 8602 9417 8636 9418
rect 8670 9417 8704 9418
rect 8738 9417 8772 9418
rect 8806 9417 8840 9418
rect 8874 9417 8908 9418
rect 8942 9417 8976 9418
rect 9010 9417 9044 9418
rect 9078 9418 9079 9451
rect 9146 9418 9151 9451
rect 9214 9418 9223 9451
rect 9282 9418 9295 9451
rect 9350 9418 9367 9451
rect 9418 9418 9439 9451
rect 9486 9418 9511 9451
rect 9554 9418 9583 9451
rect 9622 9418 9655 9451
rect 9078 9417 9112 9418
rect 9146 9417 9180 9418
rect 9214 9417 9248 9418
rect 9282 9417 9316 9418
rect 9350 9417 9384 9418
rect 9418 9417 9452 9418
rect 9486 9417 9520 9418
rect 9554 9417 9588 9418
rect 9622 9417 9656 9418
rect 9690 9417 9724 9451
rect 9761 9418 9792 9451
rect 9833 9418 9860 9451
rect 9905 9418 9928 9451
rect 9977 9418 9996 9451
rect 10049 9418 10064 9451
rect 10121 9418 10132 9451
rect 10193 9418 10200 9451
rect 10265 9418 10268 9451
rect 9758 9417 9792 9418
rect 9826 9417 9860 9418
rect 9894 9417 9928 9418
rect 9962 9417 9996 9418
rect 10030 9417 10064 9418
rect 10098 9417 10132 9418
rect 10166 9417 10200 9418
rect 10234 9417 10268 9418
rect 10302 9418 10303 9451
rect 10370 9418 10375 9451
rect 10438 9418 10447 9451
rect 10506 9418 10519 9451
rect 10574 9418 10591 9451
rect 10642 9418 10663 9451
rect 10710 9418 10735 9451
rect 10778 9418 10807 9451
rect 10846 9418 10879 9451
rect 10302 9417 10336 9418
rect 10370 9417 10404 9418
rect 10438 9417 10472 9418
rect 10506 9417 10540 9418
rect 10574 9417 10608 9418
rect 10642 9417 10676 9418
rect 10710 9417 10744 9418
rect 10778 9417 10812 9418
rect 10846 9417 10880 9418
rect 10914 9417 10948 9451
rect 10985 9418 11016 9451
rect 11057 9418 11084 9451
rect 11129 9418 11152 9451
rect 11201 9418 11220 9451
rect 11273 9418 11288 9451
rect 11345 9418 11356 9451
rect 11417 9418 11424 9451
rect 11489 9418 11492 9451
rect 10982 9417 11016 9418
rect 11050 9417 11084 9418
rect 11118 9417 11152 9418
rect 11186 9417 11220 9418
rect 11254 9417 11288 9418
rect 11322 9417 11356 9418
rect 11390 9417 11424 9418
rect 11458 9417 11492 9418
rect 11526 9418 11527 9451
rect 11594 9418 11599 9451
rect 11662 9418 11671 9451
rect 11730 9418 11743 9451
rect 11798 9418 11815 9451
rect 11866 9418 11887 9451
rect 11934 9418 11959 9451
rect 12002 9418 12031 9451
rect 12070 9418 12103 9451
rect 11526 9417 11560 9418
rect 11594 9417 11628 9418
rect 11662 9417 11696 9418
rect 11730 9417 11764 9418
rect 11798 9417 11832 9418
rect 11866 9417 11900 9418
rect 11934 9417 11968 9418
rect 12002 9417 12036 9418
rect 12070 9417 12104 9418
rect 12138 9417 12172 9451
rect 12209 9418 12240 9451
rect 12281 9418 12308 9451
rect 12353 9418 12376 9451
rect 12425 9418 12444 9451
rect 12497 9418 12512 9451
rect 12569 9418 12580 9451
rect 12641 9418 12648 9451
rect 12206 9417 12240 9418
rect 12274 9417 12308 9418
rect 12342 9417 12376 9418
rect 12410 9417 12444 9418
rect 12478 9417 12512 9418
rect 12546 9417 12580 9418
rect 12614 9417 12648 9418
rect 12682 9417 12716 9451
rect 12750 9417 12784 9451
rect 12818 9417 12852 9451
rect 12886 9417 12920 9451
rect 12954 9417 12988 9451
rect 13022 9417 13056 9451
rect 13090 9417 13124 9451
rect 13158 9417 13192 9451
rect 13226 9417 13260 9451
rect 13294 9417 13328 9451
rect 13362 9417 13396 9451
rect 13430 9417 13464 9451
rect 13498 9417 13532 9451
rect 13566 9417 13600 9451
rect 13634 9417 13668 9451
rect 13702 9417 13736 9451
rect 13770 9417 13804 9451
rect 13838 9417 13872 9451
rect 13906 9417 13940 9451
rect 13974 9417 14008 9451
rect 14042 9417 14076 9451
rect 14110 9417 14144 9451
rect 14178 9417 14212 9451
rect 14246 9417 14280 9451
rect 14348 9451 14614 9452
rect 14314 9417 14348 9418
rect 14382 9417 14416 9451
rect 14450 9417 14484 9451
rect 14518 9418 14614 9451
rect 14648 9418 14724 9452
rect 14518 9417 14724 9418
rect 245 9343 14724 9417
<< viali >>
rect 320 36500 354 36534
rect 14614 36499 14648 36533
rect 556 36497 590 36498
rect 628 36497 662 36498
rect 700 36497 734 36498
rect 772 36497 806 36498
rect 844 36497 878 36498
rect 916 36497 950 36498
rect 988 36497 1022 36498
rect 1060 36497 1094 36498
rect 1132 36497 1166 36498
rect 1204 36497 1238 36498
rect 1276 36497 1310 36498
rect 1348 36497 1382 36498
rect 1420 36497 1454 36498
rect 1492 36497 1526 36498
rect 1564 36497 1598 36498
rect 1636 36497 1670 36498
rect 1708 36497 1742 36498
rect 1780 36497 1814 36498
rect 1852 36497 1886 36498
rect 1924 36497 1958 36498
rect 1996 36497 2030 36498
rect 2068 36497 2102 36498
rect 2140 36497 2174 36498
rect 2212 36497 2246 36498
rect 2284 36497 2318 36498
rect 2356 36497 2390 36498
rect 2428 36497 2462 36498
rect 2500 36497 2534 36498
rect 2572 36497 2606 36498
rect 2644 36497 2678 36498
rect 2716 36497 2750 36498
rect 2788 36497 2822 36498
rect 2860 36497 2894 36498
rect 2932 36497 2966 36498
rect 3004 36497 3038 36498
rect 3076 36497 3110 36498
rect 3148 36497 3182 36498
rect 3220 36497 3254 36498
rect 3292 36497 3326 36498
rect 3364 36497 3398 36498
rect 3436 36497 3470 36498
rect 3508 36497 3542 36498
rect 3580 36497 3614 36498
rect 3652 36497 3686 36498
rect 3724 36497 3758 36498
rect 3796 36497 3830 36498
rect 3868 36497 3902 36498
rect 3940 36497 3974 36498
rect 4012 36497 4046 36498
rect 4084 36497 4118 36498
rect 4156 36497 4190 36498
rect 4228 36497 4262 36498
rect 4300 36497 4334 36498
rect 4372 36497 4406 36498
rect 4444 36497 4478 36498
rect 4516 36497 4550 36498
rect 4588 36497 4622 36498
rect 4660 36497 4694 36498
rect 4732 36497 4766 36498
rect 4804 36497 4838 36498
rect 4876 36497 4910 36498
rect 4948 36497 4982 36498
rect 5020 36497 5054 36498
rect 5092 36497 5126 36498
rect 5164 36497 5198 36498
rect 5236 36497 5270 36498
rect 5308 36497 5342 36498
rect 5380 36497 5414 36498
rect 5452 36497 5486 36498
rect 5524 36497 5558 36498
rect 5596 36497 5630 36498
rect 5668 36497 5702 36498
rect 5740 36497 5774 36498
rect 5812 36497 5846 36498
rect 5884 36497 5918 36498
rect 5956 36497 5990 36498
rect 6028 36497 6062 36498
rect 6100 36497 6134 36498
rect 6172 36497 6206 36498
rect 6244 36497 6278 36498
rect 6316 36497 6350 36498
rect 6388 36497 6422 36498
rect 6460 36497 6494 36498
rect 6532 36497 6566 36498
rect 6604 36497 6638 36498
rect 6676 36497 6710 36498
rect 6748 36497 6782 36498
rect 6820 36497 6854 36498
rect 6892 36497 6926 36498
rect 6964 36497 6998 36498
rect 7036 36497 7070 36498
rect 7108 36497 7142 36498
rect 7180 36497 7214 36498
rect 7252 36497 7286 36498
rect 7324 36497 7358 36498
rect 7396 36497 7430 36498
rect 7468 36497 7502 36498
rect 7540 36497 7574 36498
rect 7612 36497 7646 36498
rect 7684 36497 7718 36498
rect 7756 36497 7790 36498
rect 7828 36497 7862 36498
rect 7900 36497 7934 36498
rect 7972 36497 8006 36498
rect 8044 36497 8078 36498
rect 8116 36497 8150 36498
rect 8188 36497 8222 36498
rect 8260 36497 8294 36498
rect 8332 36497 8366 36498
rect 8404 36497 8438 36498
rect 8476 36497 8510 36498
rect 8548 36497 8582 36498
rect 8620 36497 8654 36498
rect 8692 36497 8726 36498
rect 8764 36497 8798 36498
rect 8836 36497 8870 36498
rect 8908 36497 8942 36498
rect 8980 36497 9014 36498
rect 9052 36497 9086 36498
rect 9124 36497 9158 36498
rect 9196 36497 9230 36498
rect 9268 36497 9302 36498
rect 9340 36497 9374 36498
rect 9412 36497 9446 36498
rect 9484 36497 9518 36498
rect 9556 36497 9590 36498
rect 9628 36497 9662 36498
rect 9700 36497 9734 36498
rect 9772 36497 9806 36498
rect 9844 36497 9878 36498
rect 9916 36497 9950 36498
rect 9988 36497 10022 36498
rect 10060 36497 10094 36498
rect 10132 36497 10166 36498
rect 10204 36497 10238 36498
rect 10276 36497 10310 36498
rect 10348 36497 10382 36498
rect 10420 36497 10454 36498
rect 10492 36497 10526 36498
rect 10564 36497 10598 36498
rect 10636 36497 10670 36498
rect 10708 36497 10742 36498
rect 10780 36497 10814 36498
rect 10852 36497 10886 36498
rect 10924 36497 10958 36498
rect 10996 36497 11030 36498
rect 11068 36497 11102 36498
rect 11140 36497 11174 36498
rect 11212 36497 11246 36498
rect 11284 36497 11318 36498
rect 11356 36497 11390 36498
rect 11428 36497 11462 36498
rect 11500 36497 11534 36498
rect 11572 36497 11606 36498
rect 11644 36497 11678 36498
rect 11716 36497 11750 36498
rect 11788 36497 11822 36498
rect 11860 36497 11894 36498
rect 11932 36497 11966 36498
rect 12004 36497 12038 36498
rect 12076 36497 12110 36498
rect 12148 36497 12182 36498
rect 12220 36497 12254 36498
rect 12292 36497 12326 36498
rect 12364 36497 12398 36498
rect 12436 36497 12470 36498
rect 12508 36497 12542 36498
rect 12580 36497 12614 36498
rect 12652 36497 12686 36498
rect 12724 36497 12758 36498
rect 12796 36497 12830 36498
rect 12868 36497 12902 36498
rect 12940 36497 12974 36498
rect 13012 36497 13046 36498
rect 13084 36497 13118 36498
rect 13156 36497 13190 36498
rect 13228 36497 13262 36498
rect 13300 36497 13334 36498
rect 13372 36497 13406 36498
rect 13444 36497 13478 36498
rect 13516 36497 13550 36498
rect 13588 36497 13622 36498
rect 13660 36497 13694 36498
rect 13732 36497 13766 36498
rect 13804 36497 13838 36498
rect 13876 36497 13910 36498
rect 13948 36497 13982 36498
rect 14020 36497 14054 36498
rect 14092 36497 14126 36498
rect 14164 36497 14198 36498
rect 14236 36497 14270 36498
rect 14308 36497 14342 36498
rect 14380 36497 14414 36498
rect 556 36464 557 36497
rect 557 36464 590 36497
rect 628 36464 659 36497
rect 659 36464 662 36497
rect 700 36464 727 36497
rect 727 36464 734 36497
rect 772 36464 795 36497
rect 795 36464 806 36497
rect 844 36464 863 36497
rect 863 36464 878 36497
rect 916 36464 931 36497
rect 931 36464 950 36497
rect 988 36464 999 36497
rect 999 36464 1022 36497
rect 1060 36464 1067 36497
rect 1067 36464 1094 36497
rect 1132 36464 1135 36497
rect 1135 36464 1166 36497
rect 1204 36464 1237 36497
rect 1237 36464 1238 36497
rect 1276 36464 1305 36497
rect 1305 36464 1310 36497
rect 1348 36464 1373 36497
rect 1373 36464 1382 36497
rect 1420 36464 1441 36497
rect 1441 36464 1454 36497
rect 1492 36464 1509 36497
rect 1509 36464 1526 36497
rect 1564 36464 1577 36497
rect 1577 36464 1598 36497
rect 1636 36464 1645 36497
rect 1645 36464 1670 36497
rect 1708 36464 1713 36497
rect 1713 36464 1742 36497
rect 1780 36464 1781 36497
rect 1781 36464 1814 36497
rect 1852 36464 1883 36497
rect 1883 36464 1886 36497
rect 1924 36464 1951 36497
rect 1951 36464 1958 36497
rect 1996 36464 2019 36497
rect 2019 36464 2030 36497
rect 2068 36464 2087 36497
rect 2087 36464 2102 36497
rect 2140 36464 2155 36497
rect 2155 36464 2174 36497
rect 2212 36464 2223 36497
rect 2223 36464 2246 36497
rect 2284 36464 2291 36497
rect 2291 36464 2318 36497
rect 2356 36464 2359 36497
rect 2359 36464 2390 36497
rect 2428 36464 2461 36497
rect 2461 36464 2462 36497
rect 2500 36464 2529 36497
rect 2529 36464 2534 36497
rect 2572 36464 2597 36497
rect 2597 36464 2606 36497
rect 2644 36464 2665 36497
rect 2665 36464 2678 36497
rect 2716 36464 2733 36497
rect 2733 36464 2750 36497
rect 2788 36464 2801 36497
rect 2801 36464 2822 36497
rect 2860 36464 2869 36497
rect 2869 36464 2894 36497
rect 2932 36464 2937 36497
rect 2937 36464 2966 36497
rect 3004 36464 3005 36497
rect 3005 36464 3038 36497
rect 3076 36464 3107 36497
rect 3107 36464 3110 36497
rect 3148 36464 3175 36497
rect 3175 36464 3182 36497
rect 3220 36464 3243 36497
rect 3243 36464 3254 36497
rect 3292 36464 3311 36497
rect 3311 36464 3326 36497
rect 3364 36464 3379 36497
rect 3379 36464 3398 36497
rect 3436 36464 3447 36497
rect 3447 36464 3470 36497
rect 3508 36464 3515 36497
rect 3515 36464 3542 36497
rect 3580 36464 3583 36497
rect 3583 36464 3614 36497
rect 3652 36464 3685 36497
rect 3685 36464 3686 36497
rect 3724 36464 3753 36497
rect 3753 36464 3758 36497
rect 3796 36464 3821 36497
rect 3821 36464 3830 36497
rect 3868 36464 3889 36497
rect 3889 36464 3902 36497
rect 3940 36464 3957 36497
rect 3957 36464 3974 36497
rect 4012 36464 4025 36497
rect 4025 36464 4046 36497
rect 4084 36464 4093 36497
rect 4093 36464 4118 36497
rect 4156 36464 4161 36497
rect 4161 36464 4190 36497
rect 4228 36464 4229 36497
rect 4229 36464 4262 36497
rect 4300 36464 4331 36497
rect 4331 36464 4334 36497
rect 4372 36464 4399 36497
rect 4399 36464 4406 36497
rect 4444 36464 4467 36497
rect 4467 36464 4478 36497
rect 4516 36464 4535 36497
rect 4535 36464 4550 36497
rect 4588 36464 4603 36497
rect 4603 36464 4622 36497
rect 4660 36464 4671 36497
rect 4671 36464 4694 36497
rect 4732 36464 4739 36497
rect 4739 36464 4766 36497
rect 4804 36464 4807 36497
rect 4807 36464 4838 36497
rect 4876 36464 4909 36497
rect 4909 36464 4910 36497
rect 4948 36464 4977 36497
rect 4977 36464 4982 36497
rect 5020 36464 5045 36497
rect 5045 36464 5054 36497
rect 5092 36464 5113 36497
rect 5113 36464 5126 36497
rect 5164 36464 5181 36497
rect 5181 36464 5198 36497
rect 5236 36464 5249 36497
rect 5249 36464 5270 36497
rect 5308 36464 5317 36497
rect 5317 36464 5342 36497
rect 5380 36464 5385 36497
rect 5385 36464 5414 36497
rect 5452 36464 5453 36497
rect 5453 36464 5486 36497
rect 5524 36464 5555 36497
rect 5555 36464 5558 36497
rect 5596 36464 5623 36497
rect 5623 36464 5630 36497
rect 5668 36464 5691 36497
rect 5691 36464 5702 36497
rect 5740 36464 5759 36497
rect 5759 36464 5774 36497
rect 5812 36464 5827 36497
rect 5827 36464 5846 36497
rect 5884 36464 5895 36497
rect 5895 36464 5918 36497
rect 5956 36464 5963 36497
rect 5963 36464 5990 36497
rect 6028 36464 6031 36497
rect 6031 36464 6062 36497
rect 6100 36464 6133 36497
rect 6133 36464 6134 36497
rect 6172 36464 6201 36497
rect 6201 36464 6206 36497
rect 6244 36464 6269 36497
rect 6269 36464 6278 36497
rect 6316 36464 6337 36497
rect 6337 36464 6350 36497
rect 6388 36464 6405 36497
rect 6405 36464 6422 36497
rect 6460 36464 6473 36497
rect 6473 36464 6494 36497
rect 6532 36464 6541 36497
rect 6541 36464 6566 36497
rect 6604 36464 6609 36497
rect 6609 36464 6638 36497
rect 6676 36464 6677 36497
rect 6677 36464 6710 36497
rect 6748 36464 6779 36497
rect 6779 36464 6782 36497
rect 6820 36464 6847 36497
rect 6847 36464 6854 36497
rect 6892 36464 6915 36497
rect 6915 36464 6926 36497
rect 6964 36464 6983 36497
rect 6983 36464 6998 36497
rect 7036 36464 7051 36497
rect 7051 36464 7070 36497
rect 7108 36464 7119 36497
rect 7119 36464 7142 36497
rect 7180 36464 7187 36497
rect 7187 36464 7214 36497
rect 7252 36464 7255 36497
rect 7255 36464 7286 36497
rect 7324 36464 7357 36497
rect 7357 36464 7358 36497
rect 7396 36464 7425 36497
rect 7425 36464 7430 36497
rect 7468 36464 7493 36497
rect 7493 36464 7502 36497
rect 7540 36464 7561 36497
rect 7561 36464 7574 36497
rect 7612 36464 7629 36497
rect 7629 36464 7646 36497
rect 7684 36464 7697 36497
rect 7697 36464 7718 36497
rect 7756 36464 7765 36497
rect 7765 36464 7790 36497
rect 7828 36464 7833 36497
rect 7833 36464 7862 36497
rect 7900 36464 7901 36497
rect 7901 36464 7934 36497
rect 7972 36464 8003 36497
rect 8003 36464 8006 36497
rect 8044 36464 8071 36497
rect 8071 36464 8078 36497
rect 8116 36464 8139 36497
rect 8139 36464 8150 36497
rect 8188 36464 8207 36497
rect 8207 36464 8222 36497
rect 8260 36464 8275 36497
rect 8275 36464 8294 36497
rect 8332 36464 8343 36497
rect 8343 36464 8366 36497
rect 8404 36464 8411 36497
rect 8411 36464 8438 36497
rect 8476 36464 8479 36497
rect 8479 36464 8510 36497
rect 8548 36464 8581 36497
rect 8581 36464 8582 36497
rect 8620 36464 8649 36497
rect 8649 36464 8654 36497
rect 8692 36464 8717 36497
rect 8717 36464 8726 36497
rect 8764 36464 8785 36497
rect 8785 36464 8798 36497
rect 8836 36464 8853 36497
rect 8853 36464 8870 36497
rect 8908 36464 8921 36497
rect 8921 36464 8942 36497
rect 8980 36464 8989 36497
rect 8989 36464 9014 36497
rect 9052 36464 9057 36497
rect 9057 36464 9086 36497
rect 9124 36464 9125 36497
rect 9125 36464 9158 36497
rect 9196 36464 9227 36497
rect 9227 36464 9230 36497
rect 9268 36464 9295 36497
rect 9295 36464 9302 36497
rect 9340 36464 9363 36497
rect 9363 36464 9374 36497
rect 9412 36464 9431 36497
rect 9431 36464 9446 36497
rect 9484 36464 9499 36497
rect 9499 36464 9518 36497
rect 9556 36464 9567 36497
rect 9567 36464 9590 36497
rect 9628 36464 9635 36497
rect 9635 36464 9662 36497
rect 9700 36464 9703 36497
rect 9703 36464 9734 36497
rect 9772 36464 9805 36497
rect 9805 36464 9806 36497
rect 9844 36464 9873 36497
rect 9873 36464 9878 36497
rect 9916 36464 9941 36497
rect 9941 36464 9950 36497
rect 9988 36464 10009 36497
rect 10009 36464 10022 36497
rect 10060 36464 10077 36497
rect 10077 36464 10094 36497
rect 10132 36464 10145 36497
rect 10145 36464 10166 36497
rect 10204 36464 10213 36497
rect 10213 36464 10238 36497
rect 10276 36464 10281 36497
rect 10281 36464 10310 36497
rect 10348 36464 10349 36497
rect 10349 36464 10382 36497
rect 10420 36464 10451 36497
rect 10451 36464 10454 36497
rect 10492 36464 10519 36497
rect 10519 36464 10526 36497
rect 10564 36464 10587 36497
rect 10587 36464 10598 36497
rect 10636 36464 10655 36497
rect 10655 36464 10670 36497
rect 10708 36464 10723 36497
rect 10723 36464 10742 36497
rect 10780 36464 10791 36497
rect 10791 36464 10814 36497
rect 10852 36464 10859 36497
rect 10859 36464 10886 36497
rect 10924 36464 10927 36497
rect 10927 36464 10958 36497
rect 10996 36464 11029 36497
rect 11029 36464 11030 36497
rect 11068 36464 11097 36497
rect 11097 36464 11102 36497
rect 11140 36464 11165 36497
rect 11165 36464 11174 36497
rect 11212 36464 11233 36497
rect 11233 36464 11246 36497
rect 11284 36464 11301 36497
rect 11301 36464 11318 36497
rect 11356 36464 11369 36497
rect 11369 36464 11390 36497
rect 11428 36464 11437 36497
rect 11437 36464 11462 36497
rect 11500 36464 11505 36497
rect 11505 36464 11534 36497
rect 11572 36464 11573 36497
rect 11573 36464 11606 36497
rect 11644 36464 11675 36497
rect 11675 36464 11678 36497
rect 11716 36464 11743 36497
rect 11743 36464 11750 36497
rect 11788 36464 11811 36497
rect 11811 36464 11822 36497
rect 11860 36464 11879 36497
rect 11879 36464 11894 36497
rect 11932 36464 11947 36497
rect 11947 36464 11966 36497
rect 12004 36464 12015 36497
rect 12015 36464 12038 36497
rect 12076 36464 12083 36497
rect 12083 36464 12110 36497
rect 12148 36464 12151 36497
rect 12151 36464 12182 36497
rect 12220 36464 12253 36497
rect 12253 36464 12254 36497
rect 12292 36464 12321 36497
rect 12321 36464 12326 36497
rect 12364 36464 12389 36497
rect 12389 36464 12398 36497
rect 12436 36464 12457 36497
rect 12457 36464 12470 36497
rect 12508 36464 12525 36497
rect 12525 36464 12542 36497
rect 12580 36464 12593 36497
rect 12593 36464 12614 36497
rect 12652 36464 12661 36497
rect 12661 36464 12686 36497
rect 12724 36464 12729 36497
rect 12729 36464 12758 36497
rect 12796 36464 12797 36497
rect 12797 36464 12830 36497
rect 12868 36464 12899 36497
rect 12899 36464 12902 36497
rect 12940 36464 12967 36497
rect 12967 36464 12974 36497
rect 13012 36464 13035 36497
rect 13035 36464 13046 36497
rect 13084 36464 13103 36497
rect 13103 36464 13118 36497
rect 13156 36464 13171 36497
rect 13171 36464 13190 36497
rect 13228 36464 13239 36497
rect 13239 36464 13262 36497
rect 13300 36464 13307 36497
rect 13307 36464 13334 36497
rect 13372 36464 13375 36497
rect 13375 36464 13406 36497
rect 13444 36464 13477 36497
rect 13477 36464 13478 36497
rect 13516 36464 13545 36497
rect 13545 36464 13550 36497
rect 13588 36464 13613 36497
rect 13613 36464 13622 36497
rect 13660 36464 13681 36497
rect 13681 36464 13694 36497
rect 13732 36464 13749 36497
rect 13749 36464 13766 36497
rect 13804 36464 13817 36497
rect 13817 36464 13838 36497
rect 13876 36464 13885 36497
rect 13885 36464 13910 36497
rect 13948 36464 13953 36497
rect 13953 36464 13982 36497
rect 14020 36464 14021 36497
rect 14021 36464 14054 36497
rect 14092 36464 14123 36497
rect 14123 36464 14126 36497
rect 14164 36464 14191 36497
rect 14191 36464 14198 36497
rect 14236 36464 14259 36497
rect 14259 36464 14270 36497
rect 14308 36464 14327 36497
rect 14327 36464 14342 36497
rect 14380 36464 14395 36497
rect 14395 36464 14414 36497
rect 320 36428 354 36462
rect 14614 36427 14648 36461
rect 320 36236 346 36265
rect 346 36236 354 36265
rect 320 36231 354 36236
rect 14614 36242 14641 36262
rect 14641 36242 14648 36262
rect 14614 36228 14648 36242
rect 320 36168 346 36193
rect 346 36168 354 36193
rect 320 36159 354 36168
rect 320 36100 346 36121
rect 346 36100 354 36121
rect 320 36087 354 36100
rect 320 36032 346 36049
rect 346 36032 354 36049
rect 320 36015 354 36032
rect 320 35964 346 35977
rect 346 35964 354 35977
rect 320 35943 354 35964
rect 320 35896 346 35905
rect 346 35896 354 35905
rect 320 35871 354 35896
rect 320 35828 346 35833
rect 346 35828 354 35833
rect 320 35799 354 35828
rect 320 35760 346 35761
rect 346 35760 354 35761
rect 320 35727 354 35760
rect 320 35658 354 35689
rect 320 35655 346 35658
rect 346 35655 354 35658
rect 320 35590 354 35617
rect 320 35583 346 35590
rect 346 35583 354 35590
rect 320 35522 354 35545
rect 320 35511 346 35522
rect 346 35511 354 35522
rect 320 35454 354 35473
rect 320 35439 346 35454
rect 346 35439 354 35454
rect 320 35386 354 35401
rect 320 35367 346 35386
rect 346 35367 354 35386
rect 320 35318 354 35329
rect 320 35295 346 35318
rect 346 35295 354 35318
rect 320 35250 354 35257
rect 320 35223 346 35250
rect 346 35223 354 35250
rect 320 35182 354 35185
rect 320 35151 346 35182
rect 346 35151 354 35182
rect 320 35080 346 35113
rect 346 35080 354 35113
rect 320 35079 354 35080
rect 320 35012 346 35041
rect 346 35012 354 35041
rect 320 35007 354 35012
rect 320 34944 346 34969
rect 346 34944 354 34969
rect 320 34935 354 34944
rect 320 34876 346 34897
rect 346 34876 354 34897
rect 320 34863 354 34876
rect 320 34808 346 34825
rect 346 34808 354 34825
rect 320 34791 354 34808
rect 320 34740 346 34753
rect 346 34740 354 34753
rect 320 34719 354 34740
rect 320 34672 346 34681
rect 346 34672 354 34681
rect 320 34647 354 34672
rect 320 34604 346 34609
rect 346 34604 354 34609
rect 320 34575 354 34604
rect 320 34536 346 34537
rect 346 34536 354 34537
rect 320 34503 354 34536
rect 320 34434 354 34465
rect 320 34431 346 34434
rect 346 34431 354 34434
rect 320 34366 354 34393
rect 320 34359 346 34366
rect 346 34359 354 34366
rect 320 34298 354 34321
rect 320 34287 346 34298
rect 346 34287 354 34298
rect 320 34230 354 34249
rect 320 34215 346 34230
rect 346 34215 354 34230
rect 320 34162 354 34177
rect 320 34143 346 34162
rect 346 34143 354 34162
rect 320 34094 354 34105
rect 320 34071 346 34094
rect 346 34071 354 34094
rect 320 34026 354 34033
rect 320 33999 346 34026
rect 346 33999 354 34026
rect 320 33958 354 33961
rect 320 33927 346 33958
rect 346 33927 354 33958
rect 320 33856 346 33889
rect 346 33856 354 33889
rect 320 33855 354 33856
rect 320 33788 346 33817
rect 346 33788 354 33817
rect 320 33783 354 33788
rect 320 33720 346 33745
rect 346 33720 354 33745
rect 320 33711 354 33720
rect 320 33652 346 33673
rect 346 33652 354 33673
rect 320 33639 354 33652
rect 320 33584 346 33601
rect 346 33584 354 33601
rect 320 33567 354 33584
rect 320 33516 346 33529
rect 346 33516 354 33529
rect 320 33495 354 33516
rect 320 33448 346 33457
rect 346 33448 354 33457
rect 320 33423 354 33448
rect 320 33380 346 33385
rect 346 33380 354 33385
rect 320 33351 354 33380
rect 320 33312 346 33313
rect 346 33312 354 33313
rect 320 33279 354 33312
rect 320 33210 354 33241
rect 320 33207 346 33210
rect 346 33207 354 33210
rect 320 33142 354 33169
rect 320 33135 346 33142
rect 346 33135 354 33142
rect 320 33074 354 33097
rect 320 33063 346 33074
rect 346 33063 354 33074
rect 320 33006 354 33025
rect 320 32991 346 33006
rect 346 32991 354 33006
rect 320 32938 354 32953
rect 320 32919 346 32938
rect 346 32919 354 32938
rect 320 32870 354 32881
rect 320 32847 346 32870
rect 346 32847 354 32870
rect 320 32802 354 32809
rect 320 32775 346 32802
rect 346 32775 354 32802
rect 320 32734 354 32737
rect 320 32703 346 32734
rect 346 32703 354 32734
rect 320 32632 346 32665
rect 346 32632 354 32665
rect 320 32631 354 32632
rect 320 32564 346 32593
rect 346 32564 354 32593
rect 320 32559 354 32564
rect 320 32496 346 32521
rect 346 32496 354 32521
rect 320 32487 354 32496
rect 320 32428 346 32449
rect 346 32428 354 32449
rect 320 32415 354 32428
rect 320 32360 346 32377
rect 346 32360 354 32377
rect 320 32343 354 32360
rect 320 32292 346 32305
rect 346 32292 354 32305
rect 320 32271 354 32292
rect 320 32224 346 32233
rect 346 32224 354 32233
rect 320 32199 354 32224
rect 320 32156 346 32161
rect 346 32156 354 32161
rect 320 32127 354 32156
rect 320 32088 346 32089
rect 346 32088 354 32089
rect 320 32055 354 32088
rect 320 31986 354 32017
rect 320 31983 346 31986
rect 346 31983 354 31986
rect 320 31918 354 31945
rect 320 31911 346 31918
rect 346 31911 354 31918
rect 320 31850 354 31873
rect 320 31839 346 31850
rect 346 31839 354 31850
rect 320 31782 354 31801
rect 320 31767 346 31782
rect 346 31767 354 31782
rect 320 31714 354 31729
rect 320 31695 346 31714
rect 346 31695 354 31714
rect 320 31646 354 31657
rect 320 31623 346 31646
rect 346 31623 354 31646
rect 320 31578 354 31585
rect 320 31551 346 31578
rect 346 31551 354 31578
rect 320 31510 354 31513
rect 320 31479 346 31510
rect 346 31479 354 31510
rect 320 31408 346 31441
rect 346 31408 354 31441
rect 320 31407 354 31408
rect 320 31340 346 31369
rect 346 31340 354 31369
rect 320 31335 354 31340
rect 320 31272 346 31297
rect 346 31272 354 31297
rect 320 31263 354 31272
rect 320 31204 346 31225
rect 346 31204 354 31225
rect 320 31191 354 31204
rect 320 31136 346 31153
rect 346 31136 354 31153
rect 320 31119 354 31136
rect 320 31068 346 31081
rect 346 31068 354 31081
rect 320 31047 354 31068
rect 320 31000 346 31009
rect 346 31000 354 31009
rect 320 30975 354 31000
rect 320 30932 346 30937
rect 346 30932 354 30937
rect 320 30903 354 30932
rect 320 30864 346 30865
rect 346 30864 354 30865
rect 320 30831 354 30864
rect 320 30762 354 30793
rect 320 30759 346 30762
rect 346 30759 354 30762
rect 320 30694 354 30721
rect 320 30687 346 30694
rect 346 30687 354 30694
rect 320 30626 354 30649
rect 320 30615 346 30626
rect 346 30615 354 30626
rect 320 30558 354 30577
rect 320 30543 346 30558
rect 346 30543 354 30558
rect 320 30490 354 30505
rect 320 30471 346 30490
rect 346 30471 354 30490
rect 320 30422 354 30433
rect 320 30399 346 30422
rect 346 30399 354 30422
rect 320 30354 354 30361
rect 320 30327 346 30354
rect 346 30327 354 30354
rect 320 30286 354 30289
rect 320 30255 346 30286
rect 346 30255 354 30286
rect 320 30184 346 30217
rect 346 30184 354 30217
rect 320 30183 354 30184
rect 320 30116 346 30145
rect 346 30116 354 30145
rect 320 30111 354 30116
rect 320 30048 346 30073
rect 346 30048 354 30073
rect 320 30039 354 30048
rect 320 29980 346 30001
rect 346 29980 354 30001
rect 320 29967 354 29980
rect 320 29912 346 29929
rect 346 29912 354 29929
rect 320 29895 354 29912
rect 320 29844 346 29857
rect 346 29844 354 29857
rect 320 29823 354 29844
rect 320 29776 346 29785
rect 346 29776 354 29785
rect 320 29751 354 29776
rect 320 29708 346 29713
rect 346 29708 354 29713
rect 320 29679 354 29708
rect 320 29640 346 29641
rect 346 29640 354 29641
rect 320 29607 354 29640
rect 320 29538 354 29569
rect 320 29535 346 29538
rect 346 29535 354 29538
rect 320 29470 354 29497
rect 320 29463 346 29470
rect 346 29463 354 29470
rect 320 29402 354 29425
rect 320 29391 346 29402
rect 346 29391 354 29402
rect 320 29334 354 29353
rect 320 29319 346 29334
rect 346 29319 354 29334
rect 320 29266 354 29281
rect 320 29247 346 29266
rect 346 29247 354 29266
rect 320 29198 354 29209
rect 320 29175 346 29198
rect 346 29175 354 29198
rect 320 29130 354 29137
rect 320 29103 346 29130
rect 346 29103 354 29130
rect 320 29062 354 29065
rect 320 29031 346 29062
rect 346 29031 354 29062
rect 320 28960 346 28993
rect 346 28960 354 28993
rect 320 28959 354 28960
rect 320 28892 346 28921
rect 346 28892 354 28921
rect 320 28887 354 28892
rect 320 28824 346 28849
rect 346 28824 354 28849
rect 320 28815 354 28824
rect 320 28756 346 28777
rect 346 28756 354 28777
rect 320 28743 354 28756
rect 320 28688 346 28705
rect 346 28688 354 28705
rect 320 28671 354 28688
rect 320 28620 346 28633
rect 346 28620 354 28633
rect 320 28599 354 28620
rect 320 28552 346 28561
rect 346 28552 354 28561
rect 320 28527 354 28552
rect 320 28484 346 28489
rect 346 28484 354 28489
rect 320 28455 354 28484
rect 320 28416 346 28417
rect 346 28416 354 28417
rect 320 28383 354 28416
rect 320 28314 354 28345
rect 320 28311 346 28314
rect 346 28311 354 28314
rect 320 28246 354 28273
rect 320 28239 346 28246
rect 346 28239 354 28246
rect 320 28178 354 28201
rect 320 28167 346 28178
rect 346 28167 354 28178
rect 320 28110 354 28129
rect 320 28095 346 28110
rect 346 28095 354 28110
rect 320 28042 354 28057
rect 320 28023 346 28042
rect 346 28023 354 28042
rect 320 27974 354 27985
rect 320 27951 346 27974
rect 346 27951 354 27974
rect 320 27906 354 27913
rect 320 27879 346 27906
rect 346 27879 354 27906
rect 320 27838 354 27841
rect 320 27807 346 27838
rect 346 27807 354 27838
rect 320 27736 346 27769
rect 346 27736 354 27769
rect 320 27735 354 27736
rect 320 27668 346 27697
rect 346 27668 354 27697
rect 320 27663 354 27668
rect 320 27600 346 27625
rect 346 27600 354 27625
rect 320 27591 354 27600
rect 320 27532 346 27553
rect 346 27532 354 27553
rect 320 27519 354 27532
rect 320 27464 346 27481
rect 346 27464 354 27481
rect 320 27447 354 27464
rect 320 27396 346 27409
rect 346 27396 354 27409
rect 320 27375 354 27396
rect 320 27328 346 27337
rect 346 27328 354 27337
rect 320 27303 354 27328
rect 320 27260 346 27265
rect 346 27260 354 27265
rect 320 27231 354 27260
rect 320 27192 346 27193
rect 346 27192 354 27193
rect 320 27159 354 27192
rect 320 27090 354 27121
rect 320 27087 346 27090
rect 346 27087 354 27090
rect 320 27022 354 27049
rect 320 27015 346 27022
rect 346 27015 354 27022
rect 320 26954 354 26977
rect 320 26943 346 26954
rect 346 26943 354 26954
rect 320 26886 354 26905
rect 320 26871 346 26886
rect 346 26871 354 26886
rect 320 26818 354 26833
rect 320 26799 346 26818
rect 346 26799 354 26818
rect 320 26750 354 26761
rect 320 26727 346 26750
rect 346 26727 354 26750
rect 320 26682 354 26689
rect 320 26655 346 26682
rect 346 26655 354 26682
rect 320 26614 354 26617
rect 320 26583 346 26614
rect 346 26583 354 26614
rect 320 26512 346 26545
rect 346 26512 354 26545
rect 320 26511 354 26512
rect 320 26444 346 26473
rect 346 26444 354 26473
rect 320 26439 354 26444
rect 320 26376 346 26401
rect 346 26376 354 26401
rect 320 26367 354 26376
rect 320 26308 346 26329
rect 346 26308 354 26329
rect 320 26295 354 26308
rect 320 26240 346 26257
rect 346 26240 354 26257
rect 320 26223 354 26240
rect 320 26172 346 26185
rect 346 26172 354 26185
rect 320 26151 354 26172
rect 320 26104 346 26113
rect 346 26104 354 26113
rect 320 26079 354 26104
rect 320 26036 346 26041
rect 346 26036 354 26041
rect 320 26007 354 26036
rect 320 25968 346 25969
rect 346 25968 354 25969
rect 320 25935 354 25968
rect 320 25866 354 25897
rect 320 25863 346 25866
rect 346 25863 354 25866
rect 320 25798 354 25825
rect 320 25791 346 25798
rect 346 25791 354 25798
rect 320 25730 354 25753
rect 320 25719 346 25730
rect 346 25719 354 25730
rect 320 25662 354 25681
rect 320 25647 346 25662
rect 346 25647 354 25662
rect 320 25594 354 25609
rect 320 25575 346 25594
rect 346 25575 354 25594
rect 320 25526 354 25537
rect 320 25503 346 25526
rect 346 25503 354 25526
rect 320 25458 354 25465
rect 320 25431 346 25458
rect 346 25431 354 25458
rect 320 25390 354 25393
rect 320 25359 346 25390
rect 346 25359 354 25390
rect 320 25288 346 25321
rect 346 25288 354 25321
rect 320 25287 354 25288
rect 320 25220 346 25249
rect 346 25220 354 25249
rect 320 25215 354 25220
rect 320 25152 346 25177
rect 346 25152 354 25177
rect 320 25143 354 25152
rect 320 25084 346 25105
rect 346 25084 354 25105
rect 320 25071 354 25084
rect 320 25016 346 25033
rect 346 25016 354 25033
rect 320 24999 354 25016
rect 320 24948 346 24961
rect 346 24948 354 24961
rect 320 24927 354 24948
rect 320 24880 346 24889
rect 346 24880 354 24889
rect 320 24855 354 24880
rect 320 24812 346 24817
rect 346 24812 354 24817
rect 320 24783 354 24812
rect 320 24744 346 24745
rect 346 24744 354 24745
rect 320 24711 354 24744
rect 320 24642 354 24673
rect 320 24639 346 24642
rect 346 24639 354 24642
rect 320 24574 354 24601
rect 320 24567 346 24574
rect 346 24567 354 24574
rect 320 24506 354 24529
rect 320 24495 346 24506
rect 346 24495 354 24506
rect 320 24438 354 24457
rect 320 24423 346 24438
rect 346 24423 354 24438
rect 320 24370 354 24385
rect 320 24351 346 24370
rect 346 24351 354 24370
rect 320 24302 354 24313
rect 320 24279 346 24302
rect 346 24279 354 24302
rect 320 24234 354 24241
rect 320 24207 346 24234
rect 346 24207 354 24234
rect 320 24166 354 24169
rect 320 24135 346 24166
rect 346 24135 354 24166
rect 320 24064 346 24097
rect 346 24064 354 24097
rect 320 24063 354 24064
rect 320 23996 346 24025
rect 346 23996 354 24025
rect 320 23991 354 23996
rect 320 23928 346 23953
rect 346 23928 354 23953
rect 320 23919 354 23928
rect 320 23860 346 23881
rect 346 23860 354 23881
rect 320 23847 354 23860
rect 320 23792 346 23809
rect 346 23792 354 23809
rect 320 23775 354 23792
rect 320 23724 346 23737
rect 346 23724 354 23737
rect 320 23703 354 23724
rect 320 23656 346 23665
rect 346 23656 354 23665
rect 320 23631 354 23656
rect 320 23588 346 23593
rect 346 23588 354 23593
rect 320 23559 354 23588
rect 320 23520 346 23521
rect 346 23520 354 23521
rect 320 23487 354 23520
rect 320 23418 354 23449
rect 320 23415 346 23418
rect 346 23415 354 23418
rect 320 23350 354 23377
rect 320 23343 346 23350
rect 346 23343 354 23350
rect 320 23282 354 23305
rect 320 23271 346 23282
rect 346 23271 354 23282
rect 320 23214 354 23233
rect 320 23199 346 23214
rect 346 23199 354 23214
rect 320 23146 354 23161
rect 320 23127 346 23146
rect 346 23127 354 23146
rect 320 23078 354 23089
rect 320 23055 346 23078
rect 346 23055 354 23078
rect 320 23010 354 23017
rect 320 22983 346 23010
rect 346 22983 354 23010
rect 320 22942 354 22945
rect 320 22911 346 22942
rect 346 22911 354 22942
rect 320 22840 346 22873
rect 346 22840 354 22873
rect 320 22839 354 22840
rect 320 22772 346 22801
rect 346 22772 354 22801
rect 320 22767 354 22772
rect 320 22704 346 22729
rect 346 22704 354 22729
rect 320 22695 354 22704
rect 320 22636 346 22657
rect 346 22636 354 22657
rect 320 22623 354 22636
rect 320 22568 346 22585
rect 346 22568 354 22585
rect 320 22551 354 22568
rect 320 22500 346 22513
rect 346 22500 354 22513
rect 320 22479 354 22500
rect 320 22432 346 22441
rect 346 22432 354 22441
rect 320 22407 354 22432
rect 320 22364 346 22369
rect 346 22364 354 22369
rect 320 22335 354 22364
rect 320 22296 346 22297
rect 346 22296 354 22297
rect 320 22263 354 22296
rect 320 22194 354 22225
rect 320 22191 346 22194
rect 346 22191 354 22194
rect 320 22126 354 22153
rect 320 22119 346 22126
rect 346 22119 354 22126
rect 320 22058 354 22081
rect 320 22047 346 22058
rect 346 22047 354 22058
rect 320 21990 354 22009
rect 320 21975 346 21990
rect 346 21975 354 21990
rect 320 21922 354 21937
rect 320 21903 346 21922
rect 346 21903 354 21922
rect 320 21854 354 21865
rect 320 21831 346 21854
rect 346 21831 354 21854
rect 320 21786 354 21793
rect 320 21759 346 21786
rect 346 21759 354 21786
rect 320 21718 354 21721
rect 320 21687 346 21718
rect 346 21687 354 21718
rect 320 21616 346 21649
rect 346 21616 354 21649
rect 320 21615 354 21616
rect 320 21548 346 21577
rect 346 21548 354 21577
rect 320 21543 354 21548
rect 320 21480 346 21505
rect 346 21480 354 21505
rect 320 21471 354 21480
rect 320 21412 346 21433
rect 346 21412 354 21433
rect 320 21399 354 21412
rect 320 21344 346 21361
rect 346 21344 354 21361
rect 320 21327 354 21344
rect 320 21276 346 21289
rect 346 21276 354 21289
rect 320 21255 354 21276
rect 320 21208 346 21217
rect 346 21208 354 21217
rect 320 21183 354 21208
rect 320 21140 346 21145
rect 346 21140 354 21145
rect 320 21111 354 21140
rect 320 21072 346 21073
rect 346 21072 354 21073
rect 320 21039 354 21072
rect 320 20970 354 21001
rect 320 20967 346 20970
rect 346 20967 354 20970
rect 320 20902 354 20929
rect 320 20895 346 20902
rect 346 20895 354 20902
rect 320 20834 354 20857
rect 320 20823 346 20834
rect 346 20823 354 20834
rect 320 20766 354 20785
rect 320 20751 346 20766
rect 346 20751 354 20766
rect 320 20698 354 20713
rect 320 20679 346 20698
rect 346 20679 354 20698
rect 320 20630 354 20641
rect 320 20607 346 20630
rect 346 20607 354 20630
rect 320 20562 354 20569
rect 320 20535 346 20562
rect 346 20535 354 20562
rect 320 20494 354 20497
rect 320 20463 346 20494
rect 346 20463 354 20494
rect 320 20392 346 20425
rect 346 20392 354 20425
rect 320 20391 354 20392
rect 320 20324 346 20353
rect 346 20324 354 20353
rect 320 20319 354 20324
rect 320 20256 346 20281
rect 346 20256 354 20281
rect 320 20247 354 20256
rect 320 20188 346 20209
rect 346 20188 354 20209
rect 320 20175 354 20188
rect 320 20120 346 20137
rect 346 20120 354 20137
rect 320 20103 354 20120
rect 320 20052 346 20065
rect 346 20052 354 20065
rect 320 20031 354 20052
rect 320 19984 346 19993
rect 346 19984 354 19993
rect 320 19959 354 19984
rect 320 19916 346 19921
rect 346 19916 354 19921
rect 320 19887 354 19916
rect 320 19848 346 19849
rect 346 19848 354 19849
rect 320 19815 354 19848
rect 320 19746 354 19777
rect 320 19743 346 19746
rect 346 19743 354 19746
rect 320 19678 354 19705
rect 320 19671 346 19678
rect 346 19671 354 19678
rect 320 19610 354 19633
rect 320 19599 346 19610
rect 346 19599 354 19610
rect 320 19542 354 19561
rect 320 19527 346 19542
rect 346 19527 354 19542
rect 320 19474 354 19489
rect 320 19455 346 19474
rect 346 19455 354 19474
rect 320 19406 354 19417
rect 320 19383 346 19406
rect 346 19383 354 19406
rect 320 19338 354 19345
rect 320 19311 346 19338
rect 346 19311 354 19338
rect 320 19270 354 19273
rect 320 19239 346 19270
rect 346 19239 354 19270
rect 320 19168 346 19201
rect 346 19168 354 19201
rect 320 19167 354 19168
rect 320 19100 346 19129
rect 346 19100 354 19129
rect 320 19095 354 19100
rect 320 19032 346 19057
rect 346 19032 354 19057
rect 320 19023 354 19032
rect 320 18964 346 18985
rect 346 18964 354 18985
rect 320 18951 354 18964
rect 320 18896 346 18913
rect 346 18896 354 18913
rect 320 18879 354 18896
rect 320 18828 346 18841
rect 346 18828 354 18841
rect 320 18807 354 18828
rect 320 18760 346 18769
rect 346 18760 354 18769
rect 320 18735 354 18760
rect 320 18692 346 18697
rect 346 18692 354 18697
rect 320 18663 354 18692
rect 320 18624 346 18625
rect 346 18624 354 18625
rect 320 18591 354 18624
rect 320 18522 354 18553
rect 320 18519 346 18522
rect 346 18519 354 18522
rect 320 18454 354 18481
rect 320 18447 346 18454
rect 346 18447 354 18454
rect 320 18386 354 18409
rect 320 18375 346 18386
rect 346 18375 354 18386
rect 320 18318 354 18337
rect 320 18303 346 18318
rect 346 18303 354 18318
rect 320 18250 354 18265
rect 320 18231 346 18250
rect 346 18231 354 18250
rect 320 18182 354 18193
rect 320 18159 346 18182
rect 346 18159 354 18182
rect 320 18114 354 18121
rect 320 18087 346 18114
rect 346 18087 354 18114
rect 320 18046 354 18049
rect 320 18015 346 18046
rect 346 18015 354 18046
rect 320 17944 346 17977
rect 346 17944 354 17977
rect 320 17943 354 17944
rect 320 17876 346 17905
rect 346 17876 354 17905
rect 320 17871 354 17876
rect 320 17808 346 17833
rect 346 17808 354 17833
rect 320 17799 354 17808
rect 320 17740 346 17761
rect 346 17740 354 17761
rect 320 17727 354 17740
rect 320 17672 346 17689
rect 346 17672 354 17689
rect 320 17655 354 17672
rect 320 17604 346 17617
rect 346 17604 354 17617
rect 320 17583 354 17604
rect 320 17536 346 17545
rect 346 17536 354 17545
rect 320 17511 354 17536
rect 320 17468 346 17473
rect 346 17468 354 17473
rect 320 17439 354 17468
rect 320 17400 346 17401
rect 346 17400 354 17401
rect 320 17367 354 17400
rect 320 17298 354 17329
rect 320 17295 346 17298
rect 346 17295 354 17298
rect 320 17230 354 17257
rect 320 17223 346 17230
rect 346 17223 354 17230
rect 320 17162 354 17185
rect 320 17151 346 17162
rect 346 17151 354 17162
rect 320 17094 354 17113
rect 320 17079 346 17094
rect 346 17079 354 17094
rect 320 17026 354 17041
rect 320 17007 346 17026
rect 346 17007 354 17026
rect 320 16958 354 16969
rect 320 16935 346 16958
rect 346 16935 354 16958
rect 320 16890 354 16897
rect 320 16863 346 16890
rect 346 16863 354 16890
rect 320 16822 354 16825
rect 320 16791 346 16822
rect 346 16791 354 16822
rect 320 16720 346 16753
rect 346 16720 354 16753
rect 320 16719 354 16720
rect 320 16652 346 16681
rect 346 16652 354 16681
rect 320 16647 354 16652
rect 320 16584 346 16609
rect 346 16584 354 16609
rect 320 16575 354 16584
rect 320 16516 346 16537
rect 346 16516 354 16537
rect 320 16503 354 16516
rect 320 16448 346 16465
rect 346 16448 354 16465
rect 320 16431 354 16448
rect 320 16380 346 16393
rect 346 16380 354 16393
rect 320 16359 354 16380
rect 320 16312 346 16321
rect 346 16312 354 16321
rect 320 16287 354 16312
rect 320 16244 346 16249
rect 346 16244 354 16249
rect 320 16215 354 16244
rect 320 16176 346 16177
rect 346 16176 354 16177
rect 320 16143 354 16176
rect 320 16074 354 16105
rect 320 16071 346 16074
rect 346 16071 354 16074
rect 320 16006 354 16033
rect 320 15999 346 16006
rect 346 15999 354 16006
rect 320 15938 354 15961
rect 320 15927 346 15938
rect 346 15927 354 15938
rect 320 15870 354 15889
rect 320 15855 346 15870
rect 346 15855 354 15870
rect 320 15802 354 15817
rect 320 15783 346 15802
rect 346 15783 354 15802
rect 320 15734 354 15745
rect 320 15711 346 15734
rect 346 15711 354 15734
rect 320 15666 354 15673
rect 320 15639 346 15666
rect 346 15639 354 15666
rect 320 15598 354 15601
rect 320 15567 346 15598
rect 346 15567 354 15598
rect 320 15496 346 15529
rect 346 15496 354 15529
rect 320 15495 354 15496
rect 320 15428 346 15457
rect 346 15428 354 15457
rect 320 15423 354 15428
rect 320 15360 346 15385
rect 346 15360 354 15385
rect 320 15351 354 15360
rect 320 15292 346 15313
rect 346 15292 354 15313
rect 320 15279 354 15292
rect 320 15224 346 15241
rect 346 15224 354 15241
rect 320 15207 354 15224
rect 320 15156 346 15169
rect 346 15156 354 15169
rect 320 15135 354 15156
rect 320 15088 346 15097
rect 346 15088 354 15097
rect 320 15063 354 15088
rect 320 15020 346 15025
rect 346 15020 354 15025
rect 320 14991 354 15020
rect 320 14952 346 14953
rect 346 14952 354 14953
rect 320 14919 354 14952
rect 320 14850 354 14881
rect 320 14847 346 14850
rect 346 14847 354 14850
rect 320 14782 354 14809
rect 320 14775 346 14782
rect 346 14775 354 14782
rect 320 14714 354 14737
rect 320 14703 346 14714
rect 346 14703 354 14714
rect 320 14646 354 14665
rect 320 14631 346 14646
rect 346 14631 354 14646
rect 320 14578 354 14593
rect 320 14559 346 14578
rect 346 14559 354 14578
rect 320 14510 354 14521
rect 320 14487 346 14510
rect 346 14487 354 14510
rect 320 14442 354 14449
rect 320 14415 346 14442
rect 346 14415 354 14442
rect 320 14374 354 14377
rect 320 14343 346 14374
rect 346 14343 354 14374
rect 320 14272 346 14305
rect 346 14272 354 14305
rect 320 14271 354 14272
rect 320 14204 346 14233
rect 346 14204 354 14233
rect 320 14199 354 14204
rect 320 14136 346 14161
rect 346 14136 354 14161
rect 320 14127 354 14136
rect 320 14068 346 14089
rect 346 14068 354 14089
rect 320 14055 354 14068
rect 320 14000 346 14017
rect 346 14000 354 14017
rect 320 13983 354 14000
rect 320 13932 346 13945
rect 346 13932 354 13945
rect 320 13911 354 13932
rect 320 13864 346 13873
rect 346 13864 354 13873
rect 320 13839 354 13864
rect 320 13796 346 13801
rect 346 13796 354 13801
rect 320 13767 354 13796
rect 320 13728 346 13729
rect 346 13728 354 13729
rect 320 13695 354 13728
rect 320 13626 354 13657
rect 320 13623 346 13626
rect 346 13623 354 13626
rect 320 13558 354 13585
rect 320 13551 346 13558
rect 346 13551 354 13558
rect 320 13490 354 13513
rect 320 13479 346 13490
rect 346 13479 354 13490
rect 320 13422 354 13441
rect 320 13407 346 13422
rect 346 13407 354 13422
rect 320 13354 354 13369
rect 320 13335 346 13354
rect 346 13335 354 13354
rect 320 13286 354 13297
rect 320 13263 346 13286
rect 346 13263 354 13286
rect 320 13218 354 13225
rect 320 13191 346 13218
rect 346 13191 354 13218
rect 320 13150 354 13153
rect 320 13119 346 13150
rect 346 13119 354 13150
rect 320 13048 346 13081
rect 346 13048 354 13081
rect 320 13047 354 13048
rect 320 12980 346 13009
rect 346 12980 354 13009
rect 320 12975 354 12980
rect 320 12912 346 12937
rect 346 12912 354 12937
rect 320 12903 354 12912
rect 320 12844 346 12865
rect 346 12844 354 12865
rect 320 12831 354 12844
rect 320 12776 346 12793
rect 346 12776 354 12793
rect 320 12759 354 12776
rect 320 12708 346 12721
rect 346 12708 354 12721
rect 320 12687 354 12708
rect 320 12640 346 12649
rect 346 12640 354 12649
rect 320 12615 354 12640
rect 320 12572 346 12577
rect 346 12572 354 12577
rect 320 12543 354 12572
rect 320 12504 346 12505
rect 346 12504 354 12505
rect 320 12471 354 12504
rect 320 12402 354 12433
rect 320 12399 346 12402
rect 346 12399 354 12402
rect 320 12334 354 12361
rect 320 12327 346 12334
rect 346 12327 354 12334
rect 320 12266 354 12289
rect 320 12255 346 12266
rect 346 12255 354 12266
rect 320 12198 354 12217
rect 320 12183 346 12198
rect 346 12183 354 12198
rect 320 12130 354 12145
rect 320 12111 346 12130
rect 346 12111 354 12130
rect 320 12062 354 12073
rect 320 12039 346 12062
rect 346 12039 354 12062
rect 320 11994 354 12001
rect 320 11967 346 11994
rect 346 11967 354 11994
rect 320 11926 354 11929
rect 320 11895 346 11926
rect 346 11895 354 11926
rect 320 11824 346 11857
rect 346 11824 354 11857
rect 320 11823 354 11824
rect 320 11756 346 11785
rect 346 11756 354 11785
rect 320 11751 354 11756
rect 320 11688 346 11713
rect 346 11688 354 11713
rect 320 11679 354 11688
rect 320 11620 346 11641
rect 346 11620 354 11641
rect 320 11607 354 11620
rect 320 11552 346 11569
rect 346 11552 354 11569
rect 320 11535 354 11552
rect 320 11484 346 11497
rect 346 11484 354 11497
rect 320 11463 354 11484
rect 320 11416 346 11425
rect 346 11416 354 11425
rect 320 11391 354 11416
rect 320 11348 346 11353
rect 346 11348 354 11353
rect 320 11319 354 11348
rect 320 11280 346 11281
rect 346 11280 354 11281
rect 320 11247 354 11280
rect 320 11178 354 11209
rect 320 11175 346 11178
rect 346 11175 354 11178
rect 320 11110 354 11137
rect 320 11103 346 11110
rect 346 11103 354 11110
rect 320 11042 354 11065
rect 320 11031 346 11042
rect 346 11031 354 11042
rect 320 10974 354 10993
rect 320 10959 346 10974
rect 346 10959 354 10974
rect 320 10906 354 10921
rect 320 10887 346 10906
rect 346 10887 354 10906
rect 320 10838 354 10849
rect 320 10815 346 10838
rect 346 10815 354 10838
rect 320 10770 354 10777
rect 320 10743 346 10770
rect 346 10743 354 10770
rect 320 10702 354 10705
rect 320 10671 346 10702
rect 346 10671 354 10702
rect 320 10600 346 10633
rect 346 10600 354 10633
rect 320 10599 354 10600
rect 320 10532 346 10561
rect 346 10532 354 10561
rect 320 10527 354 10532
rect 320 10464 346 10489
rect 346 10464 354 10489
rect 320 10455 354 10464
rect 320 10396 346 10417
rect 346 10396 354 10417
rect 320 10383 354 10396
rect 320 10328 346 10345
rect 346 10328 354 10345
rect 320 10311 354 10328
rect 320 10260 346 10273
rect 346 10260 354 10273
rect 320 10239 354 10260
rect 320 10192 346 10201
rect 346 10192 354 10201
rect 320 10167 354 10192
rect 320 10124 346 10129
rect 346 10124 354 10129
rect 320 10095 354 10124
rect 320 10056 346 10057
rect 346 10056 354 10057
rect 320 10023 354 10056
rect 320 9954 354 9985
rect 320 9951 346 9954
rect 346 9951 354 9954
rect 320 9886 354 9913
rect 320 9879 346 9886
rect 346 9879 354 9886
rect 320 9818 354 9841
rect 320 9807 346 9818
rect 346 9807 354 9818
rect 320 9750 354 9769
rect 320 9735 346 9750
rect 346 9735 354 9750
rect 1009 35969 1043 36003
rect 1081 35969 1115 36003
rect 1153 35969 1187 36003
rect 1225 35969 1259 36003
rect 1297 35969 1331 36003
rect 1369 35969 1403 36003
rect 1441 35969 1475 36003
rect 1513 35969 1547 36003
rect 1585 35969 1619 36003
rect 1657 35969 1691 36003
rect 1729 35969 1763 36003
rect 1801 35969 1835 36003
rect 1873 35969 1907 36003
rect 1945 35969 1979 36003
rect 2017 35969 2051 36003
rect 2089 35969 2123 36003
rect 2161 35969 2195 36003
rect 2233 35969 2267 36003
rect 2305 35969 2339 36003
rect 2377 35969 2411 36003
rect 2449 35969 2483 36003
rect 2521 35969 2555 36003
rect 2593 35969 2627 36003
rect 2665 35969 2699 36003
rect 2737 35969 2771 36003
rect 2809 35969 2843 36003
rect 2881 35969 2915 36003
rect 2953 35969 2987 36003
rect 3025 35969 3059 36003
rect 3097 35969 3131 36003
rect 3169 35969 3203 36003
rect 3241 35969 3275 36003
rect 3313 35969 3347 36003
rect 3385 35969 3419 36003
rect 3457 35969 3491 36003
rect 3529 35969 3563 36003
rect 3601 35969 3635 36003
rect 3673 35969 3707 36003
rect 3745 35969 3779 36003
rect 3817 35969 3851 36003
rect 3889 35969 3923 36003
rect 3961 35969 3995 36003
rect 4033 35969 4067 36003
rect 4105 35969 4139 36003
rect 4177 35969 4211 36003
rect 4249 35969 4283 36003
rect 4321 35969 4355 36003
rect 4393 35969 4427 36003
rect 4465 35969 4499 36003
rect 4537 35969 4571 36003
rect 4609 35969 4643 36003
rect 4681 35969 4715 36003
rect 4753 35969 4787 36003
rect 4825 35969 4859 36003
rect 4897 35969 4931 36003
rect 4969 35969 5003 36003
rect 5041 35969 5075 36003
rect 5113 35969 5147 36003
rect 5185 35969 5219 36003
rect 5257 35969 5291 36003
rect 5329 35969 5363 36003
rect 5401 35969 5435 36003
rect 5473 35969 5507 36003
rect 5545 35969 5579 36003
rect 5617 35969 5651 36003
rect 5689 35969 5723 36003
rect 5761 35969 5795 36003
rect 5833 35969 5867 36003
rect 5905 35969 5939 36003
rect 5977 35969 6011 36003
rect 6049 35969 6083 36003
rect 6121 35969 6155 36003
rect 6193 35969 6227 36003
rect 6265 35969 6299 36003
rect 6337 35969 6371 36003
rect 6409 35969 6443 36003
rect 6481 35969 6515 36003
rect 6553 35969 6587 36003
rect 6625 35969 6659 36003
rect 6697 35969 6731 36003
rect 6769 35969 6803 36003
rect 6841 35969 6875 36003
rect 6913 35969 6947 36003
rect 6985 35969 7019 36003
rect 7057 35969 7091 36003
rect 7129 35969 7163 36003
rect 7201 35969 7235 36003
rect 7273 35969 7307 36003
rect 7345 35969 7379 36003
rect 7417 35969 7451 36003
rect 7489 35969 7523 36003
rect 7561 35969 7595 36003
rect 7633 35969 7667 36003
rect 7705 35969 7739 36003
rect 7777 35969 7811 36003
rect 7849 35969 7883 36003
rect 7921 35969 7955 36003
rect 7993 35969 8027 36003
rect 8065 35969 8099 36003
rect 8137 35969 8171 36003
rect 8209 35969 8243 36003
rect 8281 35969 8315 36003
rect 8353 35969 8387 36003
rect 8425 35969 8459 36003
rect 8497 35969 8531 36003
rect 8569 35969 8603 36003
rect 8641 35969 8675 36003
rect 8713 35969 8747 36003
rect 8785 35969 8819 36003
rect 8857 35969 8891 36003
rect 8929 35969 8963 36003
rect 9001 35969 9035 36003
rect 9073 35969 9107 36003
rect 9145 35969 9179 36003
rect 9217 35969 9251 36003
rect 9289 35969 9323 36003
rect 9361 35969 9395 36003
rect 9433 35969 9467 36003
rect 9505 35969 9539 36003
rect 9577 35969 9611 36003
rect 9649 35969 9683 36003
rect 9721 35969 9755 36003
rect 9793 35969 9827 36003
rect 9865 35969 9899 36003
rect 9937 35969 9971 36003
rect 10009 35969 10043 36003
rect 10081 35969 10115 36003
rect 10153 35969 10187 36003
rect 10225 35969 10259 36003
rect 10297 35969 10331 36003
rect 10369 35969 10403 36003
rect 10441 35969 10475 36003
rect 10513 35969 10547 36003
rect 10585 35969 10619 36003
rect 10657 35969 10691 36003
rect 10729 35969 10763 36003
rect 10801 35969 10835 36003
rect 10873 35969 10907 36003
rect 10945 35969 10979 36003
rect 11017 35969 11051 36003
rect 11089 35969 11123 36003
rect 11161 35969 11195 36003
rect 11233 35969 11267 36003
rect 11305 35969 11339 36003
rect 11377 35969 11411 36003
rect 11449 35969 11483 36003
rect 11521 35969 11555 36003
rect 11593 35969 11627 36003
rect 11665 35969 11699 36003
rect 11737 35969 11771 36003
rect 11809 35969 11843 36003
rect 11881 35969 11915 36003
rect 11953 35969 11987 36003
rect 12025 35969 12059 36003
rect 12097 35969 12131 36003
rect 12169 35969 12203 36003
rect 12241 35969 12275 36003
rect 12313 35969 12347 36003
rect 12385 35969 12419 36003
rect 12457 35969 12491 36003
rect 12529 35969 12563 36003
rect 12601 35969 12635 36003
rect 12673 35969 12707 36003
rect 12745 35969 12779 36003
rect 12817 35969 12851 36003
rect 12889 35969 12923 36003
rect 12961 35969 12995 36003
rect 13033 35969 13067 36003
rect 13105 35969 13139 36003
rect 13177 35969 13211 36003
rect 13249 35969 13283 36003
rect 13321 35969 13355 36003
rect 13393 35969 13427 36003
rect 13465 35969 13499 36003
rect 13537 35969 13571 36003
rect 13609 35969 13643 36003
rect 13681 35969 13715 36003
rect 13753 35969 13787 36003
rect 13825 35969 13859 36003
rect 13897 35969 13931 36003
rect 13969 35969 14003 36003
rect 807 35850 841 35884
rect 807 35778 841 35812
rect 14122 35771 14156 35805
rect 807 35706 841 35740
rect 14122 35699 14156 35733
rect 807 35634 841 35668
rect 14122 35627 14156 35661
rect 807 35562 841 35596
rect 14122 35555 14156 35589
rect 807 35490 841 35524
rect 14122 35483 14156 35517
rect 807 35418 841 35452
rect 14122 35411 14156 35445
rect 807 35346 841 35380
rect 14122 35339 14156 35373
rect 807 35274 841 35308
rect 14122 35267 14156 35301
rect 807 35202 841 35236
rect 14122 35195 14156 35229
rect 807 35130 841 35164
rect 14122 35123 14156 35157
rect 807 35058 841 35092
rect 14122 35051 14156 35085
rect 807 34986 841 35020
rect 14122 34979 14156 35013
rect 807 34914 841 34948
rect 14122 34907 14156 34941
rect 807 34842 841 34876
rect 14122 34835 14156 34869
rect 807 34770 841 34804
rect 807 34698 841 34732
rect 14122 34763 14156 34797
rect 807 34626 841 34660
rect 807 34554 841 34588
rect 807 34482 841 34516
rect 807 34410 841 34444
rect 807 34338 841 34372
rect 807 34266 841 34300
rect 807 34194 841 34228
rect 807 34122 841 34156
rect 807 34050 841 34084
rect 807 33978 841 34012
rect 807 33906 841 33940
rect 807 33834 841 33868
rect 807 33762 841 33796
rect 807 33690 841 33724
rect 807 33618 841 33652
rect 807 33546 841 33580
rect 807 33474 841 33508
rect 807 33402 841 33436
rect 807 33330 841 33364
rect 807 33258 841 33292
rect 807 33186 841 33220
rect 807 33114 841 33148
rect 807 33042 841 33076
rect 807 32970 841 33004
rect 807 32898 841 32932
rect 807 32826 841 32860
rect 807 32754 841 32788
rect 807 32682 841 32716
rect 807 32610 841 32644
rect 807 32538 841 32572
rect 807 32466 841 32500
rect 807 32394 841 32428
rect 807 32322 841 32356
rect 807 32250 841 32284
rect 807 32178 841 32212
rect 807 32106 841 32140
rect 807 32034 841 32068
rect 807 31962 841 31996
rect 807 31890 841 31924
rect 807 31818 841 31852
rect 807 31746 841 31780
rect 807 31674 841 31708
rect 807 31602 841 31636
rect 807 31530 841 31564
rect 807 31458 841 31492
rect 807 31386 841 31420
rect 807 31314 841 31348
rect 807 31242 841 31276
rect 807 31170 841 31204
rect 807 31098 841 31132
rect 807 31026 841 31060
rect 807 30954 841 30988
rect 807 30882 841 30916
rect 807 30810 841 30844
rect 807 30738 841 30772
rect 807 30666 841 30700
rect 807 30594 841 30628
rect 807 30522 841 30556
rect 807 30450 841 30484
rect 807 30378 841 30412
rect 807 30306 841 30340
rect 807 30234 841 30268
rect 807 30162 841 30196
rect 807 30090 841 30124
rect 807 30018 841 30052
rect 807 29946 841 29980
rect 807 29874 841 29908
rect 807 29802 841 29836
rect 807 29730 841 29764
rect 807 29658 841 29692
rect 807 29586 841 29620
rect 807 29514 841 29548
rect 807 29442 841 29476
rect 807 29370 841 29404
rect 807 29298 841 29332
rect 807 29226 841 29260
rect 807 29154 841 29188
rect 807 29082 841 29116
rect 807 29010 841 29044
rect 807 28938 841 28972
rect 807 28866 841 28900
rect 807 28794 841 28828
rect 807 28722 841 28756
rect 807 28650 841 28684
rect 807 28578 841 28612
rect 807 28506 841 28540
rect 807 28434 841 28468
rect 807 28362 841 28396
rect 807 28290 841 28324
rect 807 28218 841 28252
rect 807 28146 841 28180
rect 807 28074 841 28108
rect 807 28002 841 28036
rect 807 27930 841 27964
rect 807 27858 841 27892
rect 807 27786 841 27820
rect 807 27714 841 27748
rect 807 27642 841 27676
rect 807 27570 841 27604
rect 807 27498 841 27532
rect 807 27426 841 27460
rect 807 27354 841 27388
rect 807 27282 841 27316
rect 807 27210 841 27244
rect 807 27138 841 27172
rect 807 27066 841 27100
rect 807 26994 841 27028
rect 807 26922 841 26956
rect 807 26850 841 26884
rect 807 26778 841 26812
rect 807 26706 841 26740
rect 807 26634 841 26668
rect 807 26562 841 26596
rect 807 26490 841 26524
rect 807 26418 841 26452
rect 807 26346 841 26380
rect 807 26274 841 26308
rect 807 26202 841 26236
rect 807 26130 841 26164
rect 807 26058 841 26092
rect 807 25986 841 26020
rect 807 25914 841 25948
rect 807 25842 841 25876
rect 807 25770 841 25804
rect 807 25698 841 25732
rect 807 25626 841 25660
rect 807 25554 841 25588
rect 807 25482 841 25516
rect 807 25410 841 25444
rect 807 25338 841 25372
rect 807 25266 841 25300
rect 807 25194 841 25228
rect 807 25122 841 25156
rect 807 25050 841 25084
rect 807 24978 841 25012
rect 807 24906 841 24940
rect 807 24834 841 24868
rect 807 24762 841 24796
rect 807 24690 841 24724
rect 807 24618 841 24652
rect 807 24546 841 24580
rect 807 24474 841 24508
rect 807 24402 841 24436
rect 807 24330 841 24364
rect 807 24258 841 24292
rect 807 24186 841 24220
rect 807 24114 841 24148
rect 807 24042 841 24076
rect 807 23970 841 24004
rect 807 23898 841 23932
rect 807 23826 841 23860
rect 807 23754 841 23788
rect 807 23682 841 23716
rect 807 23610 841 23644
rect 807 23538 841 23572
rect 807 23466 841 23500
rect 807 23394 841 23428
rect 807 23322 841 23356
rect 807 23250 841 23284
rect 807 23178 841 23212
rect 807 23106 841 23140
rect 807 23034 841 23068
rect 807 22962 841 22996
rect 807 22890 841 22924
rect 807 22818 841 22852
rect 807 22746 841 22780
rect 807 22674 841 22708
rect 807 22602 841 22636
rect 807 22530 841 22564
rect 807 22458 841 22492
rect 807 22386 841 22420
rect 807 22314 841 22348
rect 807 22242 841 22276
rect 807 22170 841 22204
rect 807 22098 841 22132
rect 807 22026 841 22060
rect 807 21954 841 21988
rect 807 21882 841 21916
rect 807 21810 841 21844
rect 807 21738 841 21772
rect 807 21666 841 21700
rect 807 21594 841 21628
rect 807 21522 841 21556
rect 807 21450 841 21484
rect 807 21378 841 21412
rect 807 21306 841 21340
rect 807 21234 841 21268
rect 807 21162 841 21196
rect 807 21090 841 21124
rect 807 21018 841 21052
rect 807 20946 841 20980
rect 807 20874 841 20908
rect 807 20802 841 20836
rect 807 20730 841 20764
rect 807 20658 841 20692
rect 807 20586 841 20620
rect 807 20514 841 20548
rect 807 20442 841 20476
rect 807 20370 841 20404
rect 807 20298 841 20332
rect 807 20226 841 20260
rect 807 20154 841 20188
rect 807 20082 841 20116
rect 807 20010 841 20044
rect 807 19938 841 19972
rect 807 19866 841 19900
rect 807 19794 841 19828
rect 807 19722 841 19756
rect 807 19650 841 19684
rect 807 19578 841 19612
rect 807 19506 841 19540
rect 807 19434 841 19468
rect 807 19362 841 19396
rect 807 19290 841 19324
rect 807 19218 841 19252
rect 807 19146 841 19180
rect 807 19074 841 19108
rect 807 19002 841 19036
rect 807 18930 841 18964
rect 807 18858 841 18892
rect 807 18786 841 18820
rect 807 18714 841 18748
rect 807 18642 841 18676
rect 807 18570 841 18604
rect 807 18498 841 18532
rect 807 18426 841 18460
rect 807 18354 841 18388
rect 807 18282 841 18316
rect 807 18210 841 18244
rect 807 18138 841 18172
rect 807 18066 841 18100
rect 807 17994 841 18028
rect 807 17922 841 17956
rect 807 17850 841 17884
rect 807 17778 841 17812
rect 807 17706 841 17740
rect 807 17634 841 17668
rect 807 17562 841 17596
rect 807 17490 841 17524
rect 807 17418 841 17452
rect 807 17346 841 17380
rect 807 17274 841 17308
rect 807 17202 841 17236
rect 807 17130 841 17164
rect 807 17058 841 17092
rect 807 16986 841 17020
rect 807 16914 841 16948
rect 807 16842 841 16876
rect 807 16770 841 16804
rect 807 16698 841 16732
rect 807 16626 841 16660
rect 807 16554 841 16588
rect 807 16482 841 16516
rect 807 16410 841 16444
rect 807 16338 841 16372
rect 807 16266 841 16300
rect 807 16194 841 16228
rect 807 16122 841 16156
rect 807 16050 841 16084
rect 807 15978 841 16012
rect 807 15906 841 15940
rect 807 15834 841 15868
rect 807 15762 841 15796
rect 807 15690 841 15724
rect 807 15618 841 15652
rect 807 15546 841 15580
rect 807 15474 841 15508
rect 807 15402 841 15436
rect 807 15330 841 15364
rect 807 15258 841 15292
rect 807 15186 841 15220
rect 807 15114 841 15148
rect 807 15042 841 15076
rect 807 14970 841 15004
rect 807 14898 841 14932
rect 807 14826 841 14860
rect 807 14754 841 14788
rect 807 14682 841 14716
rect 807 14610 841 14644
rect 807 14538 841 14572
rect 807 14466 841 14500
rect 807 14394 841 14428
rect 807 14322 841 14356
rect 807 14250 841 14284
rect 807 14178 841 14212
rect 807 14106 841 14140
rect 807 14034 841 14068
rect 807 13962 841 13996
rect 807 13890 841 13924
rect 807 13818 841 13852
rect 807 13746 841 13780
rect 807 13674 841 13708
rect 807 13602 841 13636
rect 807 13530 841 13564
rect 807 13458 841 13492
rect 807 13386 841 13420
rect 807 13314 841 13348
rect 807 13242 841 13276
rect 807 13170 841 13204
rect 807 13098 841 13132
rect 807 13026 841 13060
rect 807 12954 841 12988
rect 807 12882 841 12916
rect 807 12810 841 12844
rect 807 12738 841 12772
rect 807 12666 841 12700
rect 807 12594 841 12628
rect 807 12522 841 12556
rect 807 12450 841 12484
rect 807 12378 841 12412
rect 807 12306 841 12340
rect 807 12234 841 12268
rect 807 12162 841 12196
rect 807 12090 841 12124
rect 807 12018 841 12052
rect 807 11946 841 11980
rect 807 11874 841 11908
rect 807 11802 841 11836
rect 807 11730 841 11764
rect 807 11658 841 11692
rect 807 11586 841 11620
rect 807 11514 841 11548
rect 807 11442 841 11476
rect 807 11370 841 11404
rect 807 11298 841 11332
rect 807 11226 841 11260
rect 807 11154 841 11188
rect 807 11082 841 11116
rect 807 11010 841 11044
rect 807 10938 841 10972
rect 807 10866 841 10900
rect 807 10794 841 10828
rect 807 10722 841 10756
rect 807 10650 841 10684
rect 807 10578 841 10612
rect 807 10506 841 10540
rect 807 10434 841 10468
rect 807 10362 841 10396
rect 807 10290 841 10324
rect 807 10218 841 10252
rect 1301 34645 1305 34679
rect 1305 34645 1335 34679
rect 1373 34645 1407 34679
rect 1445 34645 1475 34679
rect 1475 34645 1479 34679
rect 1517 34645 1543 34679
rect 1543 34645 1551 34679
rect 1589 34645 1611 34679
rect 1611 34645 1623 34679
rect 1661 34645 1679 34679
rect 1679 34645 1695 34679
rect 1733 34645 1747 34679
rect 1747 34645 1767 34679
rect 1805 34645 1815 34679
rect 1815 34645 1839 34679
rect 1877 34645 1883 34679
rect 1883 34645 1911 34679
rect 1949 34645 1951 34679
rect 1951 34645 1983 34679
rect 2021 34645 2053 34679
rect 2053 34645 2055 34679
rect 2093 34645 2121 34679
rect 2121 34645 2127 34679
rect 2165 34645 2189 34679
rect 2189 34645 2199 34679
rect 2237 34645 2257 34679
rect 2257 34645 2271 34679
rect 2309 34645 2325 34679
rect 2325 34645 2343 34679
rect 2381 34645 2393 34679
rect 2393 34645 2415 34679
rect 2453 34645 2461 34679
rect 2461 34645 2487 34679
rect 2525 34645 2529 34679
rect 2529 34645 2559 34679
rect 2597 34645 2631 34679
rect 2669 34645 2699 34679
rect 2699 34645 2703 34679
rect 2741 34645 2767 34679
rect 2767 34645 2775 34679
rect 2813 34645 2835 34679
rect 2835 34645 2847 34679
rect 2885 34645 2903 34679
rect 2903 34645 2919 34679
rect 2957 34645 2971 34679
rect 2971 34645 2991 34679
rect 3029 34645 3039 34679
rect 3039 34645 3063 34679
rect 3101 34645 3107 34679
rect 3107 34645 3135 34679
rect 3173 34645 3175 34679
rect 3175 34645 3207 34679
rect 3245 34645 3277 34679
rect 3277 34645 3279 34679
rect 3317 34645 3345 34679
rect 3345 34645 3351 34679
rect 3389 34645 3413 34679
rect 3413 34645 3423 34679
rect 3461 34645 3481 34679
rect 3481 34645 3495 34679
rect 3533 34645 3549 34679
rect 3549 34645 3567 34679
rect 3605 34645 3617 34679
rect 3617 34645 3639 34679
rect 3677 34645 3685 34679
rect 3685 34645 3711 34679
rect 3749 34645 3753 34679
rect 3753 34645 3783 34679
rect 3821 34645 3855 34679
rect 3893 34645 3923 34679
rect 3923 34645 3927 34679
rect 3965 34645 3991 34679
rect 3991 34645 3999 34679
rect 4037 34645 4059 34679
rect 4059 34645 4071 34679
rect 4109 34645 4127 34679
rect 4127 34645 4143 34679
rect 4181 34645 4195 34679
rect 4195 34645 4215 34679
rect 4253 34645 4263 34679
rect 4263 34645 4287 34679
rect 4325 34645 4331 34679
rect 4331 34645 4359 34679
rect 4397 34645 4399 34679
rect 4399 34645 4431 34679
rect 4469 34645 4501 34679
rect 4501 34645 4503 34679
rect 4541 34645 4569 34679
rect 4569 34645 4575 34679
rect 4613 34645 4637 34679
rect 4637 34645 4647 34679
rect 4685 34645 4705 34679
rect 4705 34645 4719 34679
rect 4757 34645 4773 34679
rect 4773 34645 4791 34679
rect 4829 34645 4841 34679
rect 4841 34645 4863 34679
rect 4901 34645 4909 34679
rect 4909 34645 4935 34679
rect 4973 34645 4977 34679
rect 4977 34645 5007 34679
rect 5045 34645 5079 34679
rect 5117 34645 5147 34679
rect 5147 34645 5151 34679
rect 5189 34645 5215 34679
rect 5215 34645 5223 34679
rect 5261 34645 5283 34679
rect 5283 34645 5295 34679
rect 5333 34645 5351 34679
rect 5351 34645 5367 34679
rect 5405 34645 5419 34679
rect 5419 34645 5439 34679
rect 5477 34645 5487 34679
rect 5487 34645 5511 34679
rect 5549 34645 5555 34679
rect 5555 34645 5583 34679
rect 5621 34645 5623 34679
rect 5623 34645 5655 34679
rect 5693 34645 5725 34679
rect 5725 34645 5727 34679
rect 5765 34645 5793 34679
rect 5793 34645 5799 34679
rect 5837 34645 5861 34679
rect 5861 34645 5871 34679
rect 5909 34645 5929 34679
rect 5929 34645 5943 34679
rect 5981 34645 5997 34679
rect 5997 34645 6015 34679
rect 6053 34645 6065 34679
rect 6065 34645 6087 34679
rect 6125 34645 6133 34679
rect 6133 34645 6159 34679
rect 6197 34645 6201 34679
rect 6201 34645 6231 34679
rect 6269 34645 6303 34679
rect 6341 34645 6371 34679
rect 6371 34645 6375 34679
rect 6413 34645 6439 34679
rect 6439 34645 6447 34679
rect 6485 34645 6507 34679
rect 6507 34645 6519 34679
rect 6557 34645 6575 34679
rect 6575 34645 6591 34679
rect 6629 34645 6643 34679
rect 6643 34645 6663 34679
rect 6701 34645 6711 34679
rect 6711 34645 6735 34679
rect 6773 34645 6779 34679
rect 6779 34645 6807 34679
rect 6845 34645 6847 34679
rect 6847 34645 6879 34679
rect 6917 34645 6949 34679
rect 6949 34645 6951 34679
rect 6989 34645 7017 34679
rect 7017 34645 7023 34679
rect 7061 34645 7085 34679
rect 7085 34645 7095 34679
rect 7133 34645 7153 34679
rect 7153 34645 7167 34679
rect 7205 34645 7221 34679
rect 7221 34645 7239 34679
rect 7277 34645 7289 34679
rect 7289 34645 7311 34679
rect 7349 34645 7357 34679
rect 7357 34645 7383 34679
rect 7421 34645 7425 34679
rect 7425 34645 7455 34679
rect 7493 34645 7527 34679
rect 7565 34645 7595 34679
rect 7595 34645 7599 34679
rect 7637 34645 7663 34679
rect 7663 34645 7671 34679
rect 7709 34645 7731 34679
rect 7731 34645 7743 34679
rect 7781 34645 7799 34679
rect 7799 34645 7815 34679
rect 7853 34645 7867 34679
rect 7867 34645 7887 34679
rect 7925 34645 7935 34679
rect 7935 34645 7959 34679
rect 7997 34645 8003 34679
rect 8003 34645 8031 34679
rect 8069 34645 8071 34679
rect 8071 34645 8103 34679
rect 8141 34645 8173 34679
rect 8173 34645 8175 34679
rect 8213 34645 8241 34679
rect 8241 34645 8247 34679
rect 8285 34645 8309 34679
rect 8309 34645 8319 34679
rect 8357 34645 8377 34679
rect 8377 34645 8391 34679
rect 8429 34645 8445 34679
rect 8445 34645 8463 34679
rect 8501 34645 8513 34679
rect 8513 34645 8535 34679
rect 8573 34645 8581 34679
rect 8581 34645 8607 34679
rect 8645 34645 8649 34679
rect 8649 34645 8679 34679
rect 8717 34645 8751 34679
rect 8789 34645 8819 34679
rect 8819 34645 8823 34679
rect 8861 34645 8887 34679
rect 8887 34645 8895 34679
rect 8933 34645 8955 34679
rect 8955 34645 8967 34679
rect 9005 34645 9023 34679
rect 9023 34645 9039 34679
rect 9077 34645 9091 34679
rect 9091 34645 9111 34679
rect 9149 34645 9159 34679
rect 9159 34645 9183 34679
rect 9221 34645 9227 34679
rect 9227 34645 9255 34679
rect 9293 34645 9295 34679
rect 9295 34645 9327 34679
rect 9365 34645 9397 34679
rect 9397 34645 9399 34679
rect 9437 34645 9465 34679
rect 9465 34645 9471 34679
rect 9509 34645 9533 34679
rect 9533 34645 9543 34679
rect 9581 34645 9601 34679
rect 9601 34645 9615 34679
rect 9653 34645 9669 34679
rect 9669 34645 9687 34679
rect 9725 34645 9737 34679
rect 9737 34645 9759 34679
rect 9797 34645 9805 34679
rect 9805 34645 9831 34679
rect 9869 34645 9873 34679
rect 9873 34645 9903 34679
rect 9941 34645 9975 34679
rect 10013 34645 10043 34679
rect 10043 34645 10047 34679
rect 10085 34645 10111 34679
rect 10111 34645 10119 34679
rect 10157 34645 10179 34679
rect 10179 34645 10191 34679
rect 10229 34645 10247 34679
rect 10247 34645 10263 34679
rect 10301 34645 10315 34679
rect 10315 34645 10335 34679
rect 10373 34645 10383 34679
rect 10383 34645 10407 34679
rect 10445 34645 10451 34679
rect 10451 34645 10479 34679
rect 10517 34645 10519 34679
rect 10519 34645 10551 34679
rect 10589 34645 10621 34679
rect 10621 34645 10623 34679
rect 10661 34645 10689 34679
rect 10689 34645 10695 34679
rect 10733 34645 10757 34679
rect 10757 34645 10767 34679
rect 10805 34645 10825 34679
rect 10825 34645 10839 34679
rect 10877 34645 10893 34679
rect 10893 34645 10911 34679
rect 10949 34645 10961 34679
rect 10961 34645 10983 34679
rect 11021 34645 11029 34679
rect 11029 34645 11055 34679
rect 11093 34645 11097 34679
rect 11097 34645 11127 34679
rect 11165 34645 11199 34679
rect 11237 34645 11267 34679
rect 11267 34645 11271 34679
rect 11309 34645 11335 34679
rect 11335 34645 11343 34679
rect 11381 34645 11403 34679
rect 11403 34645 11415 34679
rect 11453 34645 11471 34679
rect 11471 34645 11487 34679
rect 11525 34645 11539 34679
rect 11539 34645 11559 34679
rect 11597 34645 11607 34679
rect 11607 34645 11631 34679
rect 11669 34645 11675 34679
rect 11675 34645 11703 34679
rect 11741 34645 11743 34679
rect 11743 34645 11775 34679
rect 11813 34645 11845 34679
rect 11845 34645 11847 34679
rect 11885 34645 11913 34679
rect 11913 34645 11919 34679
rect 11957 34645 11981 34679
rect 11981 34645 11991 34679
rect 12029 34645 12049 34679
rect 12049 34645 12063 34679
rect 12101 34645 12117 34679
rect 12117 34645 12135 34679
rect 12173 34645 12185 34679
rect 12185 34645 12207 34679
rect 12245 34645 12253 34679
rect 12253 34645 12279 34679
rect 12317 34645 12321 34679
rect 12321 34645 12351 34679
rect 12389 34645 12423 34679
rect 12461 34645 12491 34679
rect 12491 34645 12495 34679
rect 12533 34645 12559 34679
rect 12559 34645 12567 34679
rect 12605 34645 12627 34679
rect 12627 34645 12639 34679
rect 12677 34645 12695 34679
rect 12695 34645 12711 34679
rect 12749 34645 12763 34679
rect 12763 34645 12783 34679
rect 12821 34645 12831 34679
rect 12831 34645 12855 34679
rect 12893 34645 12899 34679
rect 12899 34645 12927 34679
rect 12965 34645 12967 34679
rect 12967 34645 12999 34679
rect 13037 34645 13069 34679
rect 13069 34645 13071 34679
rect 13109 34645 13137 34679
rect 13137 34645 13143 34679
rect 13181 34645 13205 34679
rect 13205 34645 13215 34679
rect 13253 34645 13273 34679
rect 13273 34645 13287 34679
rect 13325 34645 13341 34679
rect 13341 34645 13359 34679
rect 13397 34645 13409 34679
rect 13409 34645 13431 34679
rect 13469 34645 13477 34679
rect 13477 34645 13503 34679
rect 13541 34645 13545 34679
rect 13545 34645 13575 34679
rect 13613 34645 13647 34679
rect 13685 34645 13715 34679
rect 13715 34645 13719 34679
rect 1161 34444 1195 34466
rect 1161 34432 1195 34444
rect 1161 34376 1195 34394
rect 1161 34360 1195 34376
rect 1161 34308 1195 34322
rect 1161 34288 1195 34308
rect 1161 34240 1195 34250
rect 1161 34216 1195 34240
rect 1161 34172 1195 34178
rect 1161 34144 1195 34172
rect 1161 34104 1195 34106
rect 1161 34072 1195 34104
rect 1161 34002 1195 34034
rect 1161 34000 1195 34002
rect 1161 33934 1195 33962
rect 1161 33928 1195 33934
rect 1161 33866 1195 33890
rect 1161 33856 1195 33866
rect 1161 33798 1195 33818
rect 1161 33784 1195 33798
rect 1161 33730 1195 33746
rect 1161 33712 1195 33730
rect 1161 33662 1195 33674
rect 1161 33640 1195 33662
rect 1161 33594 1195 33602
rect 1161 33568 1195 33594
rect 1161 33526 1195 33530
rect 1161 33496 1195 33526
rect 1161 33424 1195 33458
rect 1161 33356 1195 33386
rect 1161 33352 1195 33356
rect 1161 33288 1195 33314
rect 1161 33280 1195 33288
rect 1161 33220 1195 33242
rect 1161 33208 1195 33220
rect 1161 33152 1195 33170
rect 1161 33136 1195 33152
rect 1161 33084 1195 33098
rect 1161 33064 1195 33084
rect 1161 33016 1195 33026
rect 1161 32992 1195 33016
rect 1161 32948 1195 32954
rect 1161 32920 1195 32948
rect 1161 32880 1195 32882
rect 1161 32848 1195 32880
rect 1161 32778 1195 32810
rect 1161 32776 1195 32778
rect 1161 32710 1195 32738
rect 1161 32704 1195 32710
rect 1161 32642 1195 32666
rect 1161 32632 1195 32642
rect 1161 32574 1195 32594
rect 1161 32560 1195 32574
rect 1161 32506 1195 32522
rect 1161 32488 1195 32506
rect 1161 32438 1195 32450
rect 1161 32416 1195 32438
rect 1161 32370 1195 32378
rect 1161 32344 1195 32370
rect 1161 32302 1195 32306
rect 1161 32272 1195 32302
rect 1161 32200 1195 32234
rect 1161 32132 1195 32162
rect 1161 32128 1195 32132
rect 1161 32064 1195 32090
rect 1161 32056 1195 32064
rect 1161 31996 1195 32018
rect 1161 31984 1195 31996
rect 1161 31928 1195 31946
rect 1161 31912 1195 31928
rect 1161 31860 1195 31874
rect 1161 31840 1195 31860
rect 1161 31792 1195 31802
rect 1161 31768 1195 31792
rect 1161 31724 1195 31730
rect 1161 31696 1195 31724
rect 1161 31656 1195 31658
rect 1161 31624 1195 31656
rect 1161 31554 1195 31586
rect 1161 31552 1195 31554
rect 1161 31486 1195 31514
rect 1161 31480 1195 31486
rect 1161 31418 1195 31442
rect 1161 31408 1195 31418
rect 1161 31350 1195 31370
rect 1161 31336 1195 31350
rect 1161 31282 1195 31298
rect 1161 31264 1195 31282
rect 1161 31214 1195 31226
rect 1161 31192 1195 31214
rect 1161 31146 1195 31154
rect 1161 31120 1195 31146
rect 1161 31078 1195 31082
rect 1161 31048 1195 31078
rect 1161 30976 1195 31010
rect 1161 30908 1195 30938
rect 1161 30904 1195 30908
rect 1161 30840 1195 30866
rect 1161 30832 1195 30840
rect 1161 30772 1195 30794
rect 1161 30760 1195 30772
rect 1161 30704 1195 30722
rect 1161 30688 1195 30704
rect 1161 30636 1195 30650
rect 1161 30616 1195 30636
rect 1161 30568 1195 30578
rect 1161 30544 1195 30568
rect 1161 30500 1195 30506
rect 1161 30472 1195 30500
rect 1161 30432 1195 30434
rect 1161 30400 1195 30432
rect 1161 30330 1195 30362
rect 1161 30328 1195 30330
rect 1161 30262 1195 30290
rect 1161 30256 1195 30262
rect 1161 30194 1195 30218
rect 1161 30184 1195 30194
rect 1161 30126 1195 30146
rect 1161 30112 1195 30126
rect 1161 30058 1195 30074
rect 1161 30040 1195 30058
rect 1161 29990 1195 30002
rect 1161 29968 1195 29990
rect 1161 29922 1195 29930
rect 1161 29896 1195 29922
rect 1161 29854 1195 29858
rect 1161 29824 1195 29854
rect 1161 29752 1195 29786
rect 1161 29684 1195 29714
rect 1161 29680 1195 29684
rect 1161 29616 1195 29642
rect 1161 29608 1195 29616
rect 1161 29548 1195 29570
rect 1161 29536 1195 29548
rect 1161 29480 1195 29498
rect 1161 29464 1195 29480
rect 1161 29412 1195 29426
rect 1161 29392 1195 29412
rect 1161 29344 1195 29354
rect 1161 29320 1195 29344
rect 1161 29276 1195 29282
rect 1161 29248 1195 29276
rect 1161 29208 1195 29210
rect 1161 29176 1195 29208
rect 1161 29106 1195 29138
rect 1161 29104 1195 29106
rect 1161 29038 1195 29066
rect 1161 29032 1195 29038
rect 1161 28970 1195 28994
rect 1161 28960 1195 28970
rect 1161 28902 1195 28922
rect 1161 28888 1195 28902
rect 13809 34473 13843 34474
rect 13809 34440 13843 34473
rect 13809 34371 13843 34402
rect 13809 34368 13843 34371
rect 13809 34303 13843 34330
rect 13809 34296 13843 34303
rect 13809 34235 13843 34258
rect 13809 34224 13843 34235
rect 13809 34167 13843 34186
rect 13809 34152 13843 34167
rect 13809 34099 13843 34114
rect 13809 34080 13843 34099
rect 13809 34031 13843 34042
rect 13809 34008 13843 34031
rect 13809 33963 13843 33970
rect 13809 33936 13843 33963
rect 13809 33895 13843 33898
rect 13809 33864 13843 33895
rect 13809 33793 13843 33826
rect 13809 33792 13843 33793
rect 13809 33725 13843 33754
rect 13809 33720 13843 33725
rect 13809 33657 13843 33682
rect 13809 33648 13843 33657
rect 13809 33589 13843 33610
rect 13809 33576 13843 33589
rect 13809 33521 13843 33538
rect 13809 33504 13843 33521
rect 13809 33453 13843 33466
rect 13809 33432 13843 33453
rect 13809 33385 13843 33394
rect 13809 33360 13843 33385
rect 13809 33317 13843 33322
rect 13809 33288 13843 33317
rect 13809 33249 13843 33250
rect 13809 33216 13843 33249
rect 13809 33147 13843 33178
rect 13809 33144 13843 33147
rect 13809 33079 13843 33106
rect 13809 33072 13843 33079
rect 13809 33011 13843 33034
rect 13809 33000 13843 33011
rect 13809 32943 13843 32962
rect 13809 32928 13843 32943
rect 13809 32875 13843 32890
rect 13809 32856 13843 32875
rect 13809 32807 13843 32818
rect 13809 32784 13843 32807
rect 13809 32739 13843 32746
rect 13809 32712 13843 32739
rect 13809 32671 13843 32674
rect 13809 32640 13843 32671
rect 13809 32569 13843 32602
rect 13809 32568 13843 32569
rect 13809 32501 13843 32530
rect 13809 32496 13843 32501
rect 13809 32433 13843 32458
rect 13809 32424 13843 32433
rect 13809 32365 13843 32386
rect 13809 32352 13843 32365
rect 13809 32297 13843 32314
rect 13809 32280 13843 32297
rect 13809 32229 13843 32242
rect 13809 32208 13843 32229
rect 13809 32161 13843 32170
rect 13809 32136 13843 32161
rect 13809 32093 13843 32098
rect 13809 32064 13843 32093
rect 13809 32025 13843 32026
rect 13809 31992 13843 32025
rect 13809 31923 13843 31954
rect 13809 31920 13843 31923
rect 13809 31855 13843 31882
rect 13809 31848 13843 31855
rect 13809 31787 13843 31810
rect 13809 31776 13843 31787
rect 13809 31719 13843 31738
rect 13809 31704 13843 31719
rect 13809 31651 13843 31666
rect 13809 31632 13843 31651
rect 13809 31583 13843 31594
rect 13809 31560 13843 31583
rect 13809 31515 13843 31522
rect 13809 31488 13843 31515
rect 13809 31447 13843 31450
rect 13809 31416 13843 31447
rect 13809 31345 13843 31378
rect 13809 31344 13843 31345
rect 13809 31277 13843 31306
rect 13809 31272 13843 31277
rect 13809 31209 13843 31234
rect 13809 31200 13843 31209
rect 13809 31141 13843 31162
rect 13809 31128 13843 31141
rect 13809 31073 13843 31090
rect 13809 31056 13843 31073
rect 13809 31005 13843 31018
rect 13809 30984 13843 31005
rect 13809 30937 13843 30946
rect 13809 30912 13843 30937
rect 13809 30869 13843 30874
rect 13809 30840 13843 30869
rect 13809 30801 13843 30802
rect 13809 30768 13843 30801
rect 13809 30699 13843 30730
rect 13809 30696 13843 30699
rect 13809 30631 13843 30658
rect 13809 30624 13843 30631
rect 13809 30563 13843 30586
rect 13809 30552 13843 30563
rect 13809 30495 13843 30514
rect 13809 30480 13843 30495
rect 13809 30427 13843 30442
rect 13809 30408 13843 30427
rect 13809 30359 13843 30370
rect 13809 30336 13843 30359
rect 13809 30291 13843 30298
rect 13809 30264 13843 30291
rect 13809 30223 13843 30226
rect 13809 30192 13843 30223
rect 13809 30121 13843 30154
rect 13809 30120 13843 30121
rect 13809 30053 13843 30082
rect 13809 30048 13843 30053
rect 13809 29985 13843 30010
rect 13809 29976 13843 29985
rect 13809 29917 13843 29938
rect 13809 29904 13843 29917
rect 13809 29849 13843 29866
rect 13809 29832 13843 29849
rect 13809 29781 13843 29794
rect 13809 29760 13843 29781
rect 13809 29713 13843 29722
rect 13809 29688 13843 29713
rect 13809 29645 13843 29650
rect 13809 29616 13843 29645
rect 13809 29577 13843 29578
rect 13809 29544 13843 29577
rect 13809 29475 13843 29506
rect 13809 29472 13843 29475
rect 13809 29407 13843 29434
rect 13809 29400 13843 29407
rect 13809 29339 13843 29362
rect 13809 29328 13843 29339
rect 13809 29271 13843 29290
rect 13809 29256 13843 29271
rect 13809 29203 13843 29218
rect 13809 29184 13843 29203
rect 13809 29135 13843 29146
rect 13809 29112 13843 29135
rect 13809 29067 13843 29074
rect 13809 29040 13843 29067
rect 13809 28999 13843 29002
rect 13809 28968 13843 28999
rect 1161 28834 1195 28850
rect 1161 28816 1195 28834
rect 1161 28766 1195 28778
rect 1161 28744 1195 28766
rect 1161 28698 1195 28706
rect 1161 28672 1195 28698
rect 1161 28630 1195 28634
rect 1161 28600 1195 28630
rect 1161 28528 1195 28562
rect 1161 28460 1195 28490
rect 1161 28456 1195 28460
rect 1161 28392 1195 28418
rect 1161 28384 1195 28392
rect 1161 28324 1195 28346
rect 1161 28312 1195 28324
rect 1161 28256 1195 28274
rect 1161 28240 1195 28256
rect 1161 28188 1195 28202
rect 1161 28168 1195 28188
rect 1161 28120 1195 28130
rect 1161 28096 1195 28120
rect 1161 28052 1195 28058
rect 1161 28024 1195 28052
rect 1161 27984 1195 27986
rect 1161 27952 1195 27984
rect 1161 27882 1195 27914
rect 1161 27880 1195 27882
rect 1161 27814 1195 27842
rect 1161 27808 1195 27814
rect 1161 27746 1195 27770
rect 1161 27736 1195 27746
rect 1161 27678 1195 27698
rect 1161 27664 1195 27678
rect 1161 27610 1195 27626
rect 1161 27592 1195 27610
rect 1161 27542 1195 27554
rect 1161 27520 1195 27542
rect 1161 27474 1195 27482
rect 1161 27448 1195 27474
rect 1161 27406 1195 27410
rect 1161 27376 1195 27406
rect 1161 27304 1195 27338
rect 1161 27236 1195 27266
rect 1161 27232 1195 27236
rect 1161 27168 1195 27194
rect 1161 27160 1195 27168
rect 1161 27100 1195 27122
rect 1161 27088 1195 27100
rect 1161 27032 1195 27050
rect 1161 27016 1195 27032
rect 1982 28553 2119 28875
rect 2119 28553 12897 28875
rect 12897 28553 13032 28875
rect 1726 28422 1976 28489
rect 1726 27504 1976 28422
rect 13031 28422 13281 28482
rect 1726 27447 1976 27504
rect 13031 27504 13281 28422
rect 13031 27440 13281 27504
rect 1985 27084 2119 27334
rect 2119 27084 12897 27334
rect 12897 27084 13035 27334
rect 13809 28897 13843 28930
rect 13809 28896 13843 28897
rect 13809 28829 13843 28858
rect 13809 28824 13843 28829
rect 13809 28761 13843 28786
rect 13809 28752 13843 28761
rect 1161 26964 1195 26978
rect 1161 26944 1195 26964
rect 1161 26896 1195 26906
rect 1161 26872 1195 26896
rect 1161 26828 1195 26834
rect 1161 26800 1195 26828
rect 1161 26760 1195 26762
rect 1161 26728 1195 26760
rect 1161 26658 1195 26690
rect 1161 26656 1195 26658
rect 1161 26590 1195 26618
rect 1161 26584 1195 26590
rect 1161 26522 1195 26546
rect 1161 26512 1195 26522
rect 1161 26454 1195 26474
rect 1161 26440 1195 26454
rect 1161 26386 1195 26402
rect 1161 26368 1195 26386
rect 1161 26318 1195 26330
rect 1161 26296 1195 26318
rect 1161 26250 1195 26258
rect 1161 26224 1195 26250
rect 1161 26182 1195 26186
rect 1161 26152 1195 26182
rect 1161 26080 1195 26114
rect 1161 26012 1195 26042
rect 1161 26008 1195 26012
rect 1161 25944 1195 25970
rect 1161 25936 1195 25944
rect 1161 25876 1195 25898
rect 1161 25864 1195 25876
rect 1161 25808 1195 25826
rect 1161 25792 1195 25808
rect 1161 25740 1195 25754
rect 1161 25720 1195 25740
rect 1161 25672 1195 25682
rect 1161 25648 1195 25672
rect 1161 25604 1195 25610
rect 1161 25576 1195 25604
rect 1161 25536 1195 25538
rect 1161 25504 1195 25536
rect 1161 25434 1195 25466
rect 1161 25432 1195 25434
rect 1161 25366 1195 25394
rect 1161 25360 1195 25366
rect 1161 25298 1195 25322
rect 1161 25288 1195 25298
rect 1161 25230 1195 25250
rect 1161 25216 1195 25230
rect 1161 25162 1195 25178
rect 1161 25144 1195 25162
rect 1161 25094 1195 25106
rect 1161 25072 1195 25094
rect 1161 25026 1195 25034
rect 1161 25000 1195 25026
rect 1161 24958 1195 24962
rect 1161 24928 1195 24958
rect 1161 24856 1195 24890
rect 1161 24788 1195 24818
rect 1161 24784 1195 24788
rect 1161 24720 1195 24746
rect 1161 24712 1195 24720
rect 1161 24652 1195 24674
rect 1161 24640 1195 24652
rect 1161 24584 1195 24602
rect 1161 24568 1195 24584
rect 1161 24516 1195 24530
rect 1161 24496 1195 24516
rect 1161 24448 1195 24458
rect 1161 24424 1195 24448
rect 1161 24380 1195 24386
rect 1161 24352 1195 24380
rect 1161 24312 1195 24314
rect 1161 24280 1195 24312
rect 1161 24210 1195 24242
rect 1161 24208 1195 24210
rect 1161 24142 1195 24170
rect 1161 24136 1195 24142
rect 1161 24074 1195 24098
rect 1161 24064 1195 24074
rect 1161 24006 1195 24026
rect 1161 23992 1195 24006
rect 1161 23938 1195 23954
rect 1161 23920 1195 23938
rect 1161 23870 1195 23882
rect 1161 23848 1195 23870
rect 1161 23802 1195 23810
rect 1161 23776 1195 23802
rect 1161 23734 1195 23738
rect 1161 23704 1195 23734
rect 1161 23632 1195 23666
rect 1161 23564 1195 23594
rect 1161 23560 1195 23564
rect 1161 23496 1195 23522
rect 1161 23488 1195 23496
rect 1161 23428 1195 23450
rect 1161 23416 1195 23428
rect 1161 23360 1195 23378
rect 1161 23344 1195 23360
rect 1161 23292 1195 23306
rect 1161 23272 1195 23292
rect 1161 23224 1195 23234
rect 1161 23200 1195 23224
rect 1161 23156 1195 23162
rect 1161 23128 1195 23156
rect 1161 23088 1195 23090
rect 1161 23056 1195 23088
rect 1161 22986 1195 23018
rect 1161 22984 1195 22986
rect 1161 22918 1195 22946
rect 1161 22912 1195 22918
rect 1161 22850 1195 22874
rect 1161 22840 1195 22850
rect 1161 22782 1195 22802
rect 1161 22768 1195 22782
rect 1161 22714 1195 22730
rect 1161 22696 1195 22714
rect 1161 22646 1195 22658
rect 1161 22624 1195 22646
rect 1161 22578 1195 22586
rect 1161 22552 1195 22578
rect 1161 22510 1195 22514
rect 1161 22480 1195 22510
rect 1161 22408 1195 22442
rect 1161 22340 1195 22370
rect 1161 22336 1195 22340
rect 1161 22272 1195 22298
rect 1161 22264 1195 22272
rect 1161 22204 1195 22226
rect 1161 22192 1195 22204
rect 1161 22136 1195 22154
rect 1161 22120 1195 22136
rect 1161 22068 1195 22082
rect 1161 22048 1195 22068
rect 1161 22000 1195 22010
rect 1161 21976 1195 22000
rect 1161 21932 1195 21938
rect 1161 21904 1195 21932
rect 1161 21864 1195 21866
rect 1161 21832 1195 21864
rect 1161 21762 1195 21794
rect 1161 21760 1195 21762
rect 1161 21694 1195 21722
rect 1161 21688 1195 21694
rect 1161 21626 1195 21650
rect 1161 21616 1195 21626
rect 1161 21558 1195 21578
rect 1161 21544 1195 21558
rect 1161 21490 1195 21506
rect 1161 21472 1195 21490
rect 1161 21422 1195 21434
rect 1161 21400 1195 21422
rect 1161 21354 1195 21362
rect 1161 21328 1195 21354
rect 1161 21286 1195 21290
rect 1161 21256 1195 21286
rect 1161 21184 1195 21218
rect 1161 21116 1195 21146
rect 1161 21112 1195 21116
rect 1161 21048 1195 21074
rect 1161 21040 1195 21048
rect 1161 20980 1195 21002
rect 1161 20968 1195 20980
rect 1161 20912 1195 20930
rect 1161 20896 1195 20912
rect 1161 20844 1195 20858
rect 1161 20824 1195 20844
rect 1161 20776 1195 20786
rect 1161 20752 1195 20776
rect 1161 20708 1195 20714
rect 1161 20680 1195 20708
rect 1161 20640 1195 20642
rect 1161 20608 1195 20640
rect 1161 20538 1195 20570
rect 1161 20536 1195 20538
rect 1161 20470 1195 20498
rect 1161 20464 1195 20470
rect 1161 20402 1195 20426
rect 1161 20392 1195 20402
rect 1161 20334 1195 20354
rect 1161 20320 1195 20334
rect 1161 20266 1195 20282
rect 1161 20248 1195 20266
rect 1161 20198 1195 20210
rect 1161 20176 1195 20198
rect 1161 20130 1195 20138
rect 1161 20104 1195 20130
rect 1161 20062 1195 20066
rect 1161 20032 1195 20062
rect 1161 19960 1195 19994
rect 1161 19892 1195 19922
rect 1161 19888 1195 19892
rect 1161 19824 1195 19850
rect 1161 19816 1195 19824
rect 1161 19756 1195 19778
rect 1161 19744 1195 19756
rect 1161 19688 1195 19706
rect 1161 19672 1195 19688
rect 1161 19620 1195 19634
rect 1161 19600 1195 19620
rect 1161 19552 1195 19562
rect 1161 19528 1195 19552
rect 1161 19484 1195 19490
rect 1161 19456 1195 19484
rect 1161 19416 1195 19418
rect 1161 19384 1195 19416
rect 1161 19314 1195 19346
rect 1161 19312 1195 19314
rect 1161 19246 1195 19274
rect 1161 19240 1195 19246
rect 1161 19178 1195 19202
rect 1161 19168 1195 19178
rect 1161 19110 1195 19130
rect 1161 19096 1195 19110
rect 1161 19042 1195 19058
rect 1161 19024 1195 19042
rect 1161 18974 1195 18986
rect 1161 18952 1195 18974
rect 1161 18906 1195 18914
rect 1161 18880 1195 18906
rect 1161 18838 1195 18842
rect 1161 18808 1195 18838
rect 1161 18736 1195 18770
rect 1161 18668 1195 18698
rect 1161 18664 1195 18668
rect 1161 18600 1195 18626
rect 1161 18592 1195 18600
rect 1161 18532 1195 18554
rect 1161 18520 1195 18532
rect 1161 18464 1195 18482
rect 1161 18448 1195 18464
rect 1161 18396 1195 18410
rect 1161 18376 1195 18396
rect 1161 18328 1195 18338
rect 1161 18304 1195 18328
rect 1161 18260 1195 18266
rect 1161 18232 1195 18260
rect 1161 18192 1195 18194
rect 1161 18160 1195 18192
rect 1161 18090 1195 18122
rect 1161 18088 1195 18090
rect 1161 18022 1195 18050
rect 1161 18016 1195 18022
rect 1161 17954 1195 17978
rect 1161 17944 1195 17954
rect 1161 17886 1195 17906
rect 1161 17872 1195 17886
rect 1161 17818 1195 17834
rect 1161 17800 1195 17818
rect 1161 17750 1195 17762
rect 1161 17728 1195 17750
rect 1161 17682 1195 17690
rect 1161 17656 1195 17682
rect 1161 17614 1195 17618
rect 1161 17584 1195 17614
rect 1161 17512 1195 17546
rect 1161 17444 1195 17474
rect 1161 17440 1195 17444
rect 1161 17376 1195 17402
rect 1161 17368 1195 17376
rect 1161 17308 1195 17330
rect 1161 17296 1195 17308
rect 1161 17240 1195 17258
rect 1161 17224 1195 17240
rect 1161 17172 1195 17186
rect 1161 17152 1195 17172
rect 1161 17104 1195 17114
rect 1161 17080 1195 17104
rect 1161 17036 1195 17042
rect 1161 17008 1195 17036
rect 1161 16968 1195 16970
rect 1161 16936 1195 16968
rect 1161 16866 1195 16898
rect 1161 16864 1195 16866
rect 1161 16798 1195 16826
rect 1161 16792 1195 16798
rect 1161 16730 1195 16754
rect 1161 16720 1195 16730
rect 1161 16662 1195 16682
rect 1161 16648 1195 16662
rect 1161 16594 1195 16610
rect 1161 16576 1195 16594
rect 1161 16526 1195 16538
rect 1161 16504 1195 16526
rect 1161 16458 1195 16466
rect 1161 16432 1195 16458
rect 1161 16390 1195 16394
rect 1161 16360 1195 16390
rect 1161 16288 1195 16322
rect 1161 16220 1195 16250
rect 1161 16216 1195 16220
rect 1161 16152 1195 16178
rect 1161 16144 1195 16152
rect 1161 16084 1195 16106
rect 1161 16072 1195 16084
rect 1161 16016 1195 16034
rect 1161 16000 1195 16016
rect 1161 15948 1195 15962
rect 1161 15928 1195 15948
rect 1161 15880 1195 15890
rect 1161 15856 1195 15880
rect 1161 15812 1195 15818
rect 1161 15784 1195 15812
rect 1161 15744 1195 15746
rect 1161 15712 1195 15744
rect 1161 15642 1195 15674
rect 1161 15640 1195 15642
rect 1161 15574 1195 15602
rect 1161 15568 1195 15574
rect 1161 15506 1195 15530
rect 1161 15496 1195 15506
rect 1161 15438 1195 15458
rect 1161 15424 1195 15438
rect 1161 15370 1195 15386
rect 1161 15352 1195 15370
rect 1161 15302 1195 15314
rect 1161 15280 1195 15302
rect 1161 15234 1195 15242
rect 1161 15208 1195 15234
rect 1161 15166 1195 15170
rect 1161 15136 1195 15166
rect 1161 15064 1195 15098
rect 1161 14996 1195 15026
rect 1161 14992 1195 14996
rect 1161 14928 1195 14954
rect 1161 14920 1195 14928
rect 1161 14860 1195 14882
rect 1161 14848 1195 14860
rect 1161 14792 1195 14810
rect 1161 14776 1195 14792
rect 1161 14724 1195 14738
rect 1161 14704 1195 14724
rect 1161 14656 1195 14666
rect 1161 14632 1195 14656
rect 1161 14588 1195 14594
rect 1161 14560 1195 14588
rect 1161 14520 1195 14522
rect 1161 14488 1195 14520
rect 1161 14418 1195 14450
rect 1161 14416 1195 14418
rect 1161 14350 1195 14378
rect 1161 14344 1195 14350
rect 1161 14282 1195 14306
rect 1161 14272 1195 14282
rect 1161 14214 1195 14234
rect 1161 14200 1195 14214
rect 1161 14146 1195 14162
rect 1161 14128 1195 14146
rect 1161 14078 1195 14090
rect 1161 14056 1195 14078
rect 1161 14010 1195 14018
rect 1161 13984 1195 14010
rect 1161 13942 1195 13946
rect 1161 13912 1195 13942
rect 1161 13840 1195 13874
rect 1161 13772 1195 13802
rect 1161 13768 1195 13772
rect 1161 13704 1195 13730
rect 1161 13696 1195 13704
rect 1161 13636 1195 13658
rect 1161 13624 1195 13636
rect 1161 13568 1195 13586
rect 1161 13552 1195 13568
rect 1161 13500 1195 13514
rect 1161 13480 1195 13500
rect 1161 13432 1195 13442
rect 1161 13408 1195 13432
rect 1161 13364 1195 13370
rect 1161 13336 1195 13364
rect 1161 13296 1195 13298
rect 1161 13264 1195 13296
rect 1161 13194 1195 13226
rect 1161 13192 1195 13194
rect 1161 13126 1195 13154
rect 1161 13120 1195 13126
rect 1161 13058 1195 13082
rect 1161 13048 1195 13058
rect 1161 12990 1195 13010
rect 1161 12976 1195 12990
rect 1161 12922 1195 12938
rect 1161 12904 1195 12922
rect 1161 12854 1195 12866
rect 1161 12832 1195 12854
rect 1161 12786 1195 12794
rect 1161 12760 1195 12786
rect 1161 12718 1195 12722
rect 1161 12688 1195 12718
rect 1161 12616 1195 12650
rect 1161 12548 1195 12578
rect 1161 12544 1195 12548
rect 1161 12480 1195 12506
rect 1161 12472 1195 12480
rect 1161 12412 1195 12434
rect 1161 12400 1195 12412
rect 1161 12344 1195 12362
rect 1161 12328 1195 12344
rect 1161 12276 1195 12290
rect 1161 12256 1195 12276
rect 1161 12208 1195 12218
rect 1161 12184 1195 12208
rect 1161 12140 1195 12146
rect 1161 12112 1195 12140
rect 1161 12072 1195 12074
rect 1161 12040 1195 12072
rect 1161 11970 1195 12002
rect 1161 11968 1195 11970
rect 1161 11902 1195 11930
rect 1161 11896 1195 11902
rect 1161 11834 1195 11858
rect 1161 11824 1195 11834
rect 1161 11766 1195 11786
rect 1161 11752 1195 11766
rect 1161 11698 1195 11714
rect 1161 11680 1195 11698
rect 1161 11630 1195 11642
rect 1161 11608 1195 11630
rect 1161 11562 1195 11570
rect 1161 11536 1195 11562
rect 1161 11494 1195 11498
rect 1161 11464 1195 11494
rect 1161 11392 1195 11426
rect 1161 11324 1195 11354
rect 1161 11320 1195 11324
rect 1161 11256 1195 11282
rect 1161 11248 1195 11256
rect 1161 11188 1195 11210
rect 1161 11176 1195 11188
rect 1161 11120 1195 11138
rect 1161 11104 1195 11120
rect 1161 11052 1195 11066
rect 1161 11032 1195 11052
rect 1161 10984 1195 10994
rect 1161 10960 1195 10984
rect 1161 10916 1195 10922
rect 1161 10888 1195 10916
rect 1161 10848 1195 10850
rect 1161 10816 1195 10848
rect 1161 10746 1195 10778
rect 1161 10744 1195 10746
rect 1161 10678 1195 10706
rect 1161 10672 1195 10678
rect 1161 10610 1195 10634
rect 1161 10600 1195 10610
rect 1161 10542 1195 10562
rect 1161 10528 1195 10542
rect 1161 10474 1195 10490
rect 1161 10456 1195 10474
rect 1161 10406 1195 10418
rect 1161 10384 1195 10406
rect 13809 23355 13843 23381
rect 13809 23347 13843 23355
rect 13809 23287 13843 23309
rect 13809 23275 13843 23287
rect 13809 23219 13843 23237
rect 13809 23203 13843 23219
rect 13809 23151 13843 23165
rect 13809 23131 13843 23151
rect 13809 23083 13843 23093
rect 13809 23059 13843 23083
rect 13809 23015 13843 23021
rect 13809 22987 13843 23015
rect 13809 22947 13843 22949
rect 13809 22915 13843 22947
rect 13809 22845 13843 22877
rect 13809 22843 13843 22845
rect 13809 22777 13843 22805
rect 13809 22771 13843 22777
rect 13809 22709 13843 22733
rect 13809 22699 13843 22709
rect 13809 22641 13843 22661
rect 13809 22627 13843 22641
rect 13809 22573 13843 22589
rect 13809 22555 13843 22573
rect 13809 22505 13843 22517
rect 13809 22483 13843 22505
rect 13809 22437 13843 22445
rect 13809 22411 13843 22437
rect 13809 22369 13843 22373
rect 13809 22339 13843 22369
rect 13809 22267 13843 22301
rect 13809 22199 13843 22229
rect 13809 22195 13843 22199
rect 13809 22131 13843 22157
rect 13809 22123 13843 22131
rect 13809 22063 13843 22085
rect 13809 22051 13843 22063
rect 13809 21995 13843 22013
rect 13809 21979 13843 21995
rect 13809 21927 13843 21941
rect 13809 21907 13843 21927
rect 13809 21859 13843 21869
rect 13809 21835 13843 21859
rect 13809 21791 13843 21797
rect 13809 21763 13843 21791
rect 13809 21723 13843 21725
rect 13809 21691 13843 21723
rect 13809 21621 13843 21653
rect 13809 21619 13843 21621
rect 13809 21553 13843 21581
rect 13809 21547 13843 21553
rect 13809 21485 13843 21509
rect 13809 21475 13843 21485
rect 13809 21417 13843 21437
rect 13809 21403 13843 21417
rect 13809 21349 13843 21365
rect 13809 21331 13843 21349
rect 13809 21281 13843 21293
rect 13809 21259 13843 21281
rect 13809 21213 13843 21221
rect 13809 21187 13843 21213
rect 13809 21145 13843 21149
rect 13809 21115 13843 21145
rect 13809 21043 13843 21077
rect 13809 20975 13843 21005
rect 13809 20971 13843 20975
rect 13809 20907 13843 20933
rect 13809 20899 13843 20907
rect 13809 20839 13843 20861
rect 13809 20827 13843 20839
rect 13809 20771 13843 20789
rect 13809 20755 13843 20771
rect 13809 20703 13843 20717
rect 13809 20683 13843 20703
rect 13809 20635 13843 20645
rect 13809 20611 13843 20635
rect 13809 20567 13843 20573
rect 13809 20539 13843 20567
rect 13809 20499 13843 20501
rect 13809 20467 13843 20499
rect 13809 20397 13843 20429
rect 13809 20395 13843 20397
rect 13809 20329 13843 20357
rect 13809 20323 13843 20329
rect 13809 20261 13843 20285
rect 13809 20251 13843 20261
rect 13809 20193 13843 20213
rect 13809 20179 13843 20193
rect 13809 20125 13843 20141
rect 13809 20107 13843 20125
rect 13809 20057 13843 20069
rect 13809 20035 13843 20057
rect 13809 19989 13843 19997
rect 13809 19963 13843 19989
rect 13809 19921 13843 19925
rect 13809 19891 13843 19921
rect 13809 19819 13843 19853
rect 13809 19751 13843 19781
rect 13809 19747 13843 19751
rect 13809 19683 13843 19709
rect 13809 19675 13843 19683
rect 13809 19615 13843 19637
rect 13809 19603 13843 19615
rect 13809 19547 13843 19565
rect 13809 19531 13843 19547
rect 13809 19479 13843 19493
rect 13809 19459 13843 19479
rect 13809 19411 13843 19421
rect 13809 19387 13843 19411
rect 13809 19343 13843 19349
rect 13809 19315 13843 19343
rect 13809 19275 13843 19277
rect 13809 19243 13843 19275
rect 13809 19173 13843 19205
rect 13809 19171 13843 19173
rect 13809 19105 13843 19133
rect 13809 19099 13843 19105
rect 13809 19037 13843 19061
rect 13809 19027 13843 19037
rect 13809 18969 13843 18989
rect 13809 18955 13843 18969
rect 13809 18901 13843 18917
rect 13809 18883 13843 18901
rect 13809 18833 13843 18845
rect 13809 18811 13843 18833
rect 13809 18765 13843 18773
rect 13809 18739 13843 18765
rect 13809 18697 13843 18701
rect 13809 18667 13843 18697
rect 13809 18595 13843 18629
rect 13809 18527 13843 18557
rect 13809 18523 13843 18527
rect 13809 18459 13843 18485
rect 13809 18451 13843 18459
rect 13809 18391 13843 18413
rect 13809 18379 13843 18391
rect 13809 18323 13843 18341
rect 13809 18307 13843 18323
rect 13809 18255 13843 18269
rect 13809 18235 13843 18255
rect 13809 18187 13843 18197
rect 13809 18163 13843 18187
rect 13809 18119 13843 18125
rect 13809 18091 13843 18119
rect 13809 18051 13843 18053
rect 13809 18019 13843 18051
rect 13809 17949 13843 17981
rect 13809 17947 13843 17949
rect 13809 17881 13843 17909
rect 13809 17875 13843 17881
rect 13809 17813 13843 17837
rect 13809 17803 13843 17813
rect 13809 17745 13843 17765
rect 13809 17731 13843 17745
rect 13809 17677 13843 17693
rect 13809 17659 13843 17677
rect 13809 17609 13843 17621
rect 13809 17587 13843 17609
rect 13809 17541 13843 17549
rect 13809 17515 13843 17541
rect 13809 17473 13843 17477
rect 13809 17443 13843 17473
rect 13809 17371 13843 17405
rect 13809 17303 13843 17333
rect 13809 17299 13843 17303
rect 13809 17235 13843 17261
rect 13809 17227 13843 17235
rect 13809 17167 13843 17189
rect 13809 17155 13843 17167
rect 13809 17099 13843 17117
rect 13809 17083 13843 17099
rect 13809 17031 13843 17045
rect 13809 17011 13843 17031
rect 13809 16963 13843 16973
rect 13809 16939 13843 16963
rect 13809 16895 13843 16901
rect 13809 16867 13843 16895
rect 13809 16827 13843 16829
rect 13809 16795 13843 16827
rect 13809 16725 13843 16757
rect 13809 16723 13843 16725
rect 13809 16657 13843 16685
rect 13809 16651 13843 16657
rect 13809 16589 13843 16613
rect 13809 16579 13843 16589
rect 13809 16521 13843 16541
rect 13809 16507 13843 16521
rect 13809 16453 13843 16469
rect 13809 16435 13843 16453
rect 13809 16385 13843 16397
rect 13809 16363 13843 16385
rect 13809 16317 13843 16325
rect 13809 16291 13843 16317
rect 13809 16249 13843 16253
rect 13809 16219 13843 16249
rect 13809 16147 13843 16181
rect 13809 16079 13843 16109
rect 13809 16075 13843 16079
rect 13809 16011 13843 16037
rect 13809 16003 13843 16011
rect 13809 15943 13843 15965
rect 13809 15931 13843 15943
rect 13809 15875 13843 15893
rect 13809 15859 13843 15875
rect 13809 15807 13843 15821
rect 13809 15787 13843 15807
rect 13809 15739 13843 15749
rect 13809 15715 13843 15739
rect 13809 15671 13843 15677
rect 13809 15643 13843 15671
rect 13809 15603 13843 15605
rect 13809 15571 13843 15603
rect 13809 15501 13843 15533
rect 13809 15499 13843 15501
rect 13809 15433 13843 15461
rect 13809 15427 13843 15433
rect 13809 15365 13843 15389
rect 13809 15355 13843 15365
rect 13809 15297 13843 15317
rect 13809 15283 13843 15297
rect 13809 15229 13843 15245
rect 13809 15211 13843 15229
rect 13809 15161 13843 15173
rect 13809 15139 13843 15161
rect 13809 15093 13843 15101
rect 13809 15067 13843 15093
rect 13809 15025 13843 15029
rect 13809 14995 13843 15025
rect 13809 14923 13843 14957
rect 13809 14855 13843 14885
rect 13809 14851 13843 14855
rect 13809 14787 13843 14813
rect 13809 14779 13843 14787
rect 13809 14719 13843 14741
rect 13809 14707 13843 14719
rect 13809 14651 13843 14669
rect 13809 14635 13843 14651
rect 13809 14583 13843 14597
rect 13809 14563 13843 14583
rect 13809 14515 13843 14525
rect 13809 14491 13843 14515
rect 13809 14447 13843 14453
rect 13809 14419 13843 14447
rect 13809 14379 13843 14381
rect 13809 14347 13843 14379
rect 13809 14277 13843 14309
rect 13809 14275 13843 14277
rect 13809 14209 13843 14237
rect 13809 14203 13843 14209
rect 13809 14141 13843 14165
rect 13809 14131 13843 14141
rect 13809 14073 13843 14093
rect 13809 14059 13843 14073
rect 13809 14005 13843 14021
rect 13809 13987 13843 14005
rect 13809 13937 13843 13949
rect 13809 13915 13843 13937
rect 13809 13869 13843 13877
rect 13809 13843 13843 13869
rect 13809 13801 13843 13805
rect 13809 13771 13843 13801
rect 13809 13699 13843 13733
rect 13809 13631 13843 13661
rect 13809 13627 13843 13631
rect 13809 13563 13843 13589
rect 13809 13555 13843 13563
rect 13809 13495 13843 13517
rect 13809 13483 13843 13495
rect 13809 13427 13843 13445
rect 13809 13411 13843 13427
rect 13809 13359 13843 13373
rect 13809 13339 13843 13359
rect 13809 13291 13843 13301
rect 13809 13267 13843 13291
rect 13809 13223 13843 13229
rect 13809 13195 13843 13223
rect 13809 13155 13843 13157
rect 13809 13123 13843 13155
rect 13809 13053 13843 13085
rect 13809 13051 13843 13053
rect 13809 12985 13843 13013
rect 13809 12979 13843 12985
rect 13809 12917 13843 12941
rect 13809 12907 13843 12917
rect 13809 12849 13843 12869
rect 13809 12835 13843 12849
rect 13809 12781 13843 12797
rect 13809 12763 13843 12781
rect 13809 12713 13843 12725
rect 13809 12691 13843 12713
rect 13809 12645 13843 12653
rect 13809 12619 13843 12645
rect 13809 12577 13843 12581
rect 13809 12547 13843 12577
rect 13809 12475 13843 12509
rect 13809 12407 13843 12437
rect 13809 12403 13843 12407
rect 13809 12339 13843 12365
rect 13809 12331 13843 12339
rect 13809 12271 13843 12293
rect 13809 12259 13843 12271
rect 13809 12203 13843 12221
rect 13809 12187 13843 12203
rect 13809 12135 13843 12149
rect 13809 12115 13843 12135
rect 13809 12067 13843 12077
rect 13809 12043 13843 12067
rect 13809 11999 13843 12005
rect 13809 11971 13843 11999
rect 13809 11931 13843 11933
rect 13809 11899 13843 11931
rect 13809 11829 13843 11861
rect 13809 11827 13843 11829
rect 13809 11761 13843 11789
rect 13809 11755 13843 11761
rect 13809 11693 13843 11717
rect 13809 11683 13843 11693
rect 13809 11625 13843 11645
rect 13809 11611 13843 11625
rect 13809 11557 13843 11573
rect 13809 11539 13843 11557
rect 13809 11489 13843 11501
rect 13809 11467 13843 11489
rect 13809 11421 13843 11429
rect 13809 11395 13843 11421
rect 13809 11353 13843 11357
rect 13809 11323 13843 11353
rect 13809 11251 13843 11285
rect 13809 11183 13843 11213
rect 13809 11179 13843 11183
rect 13809 11115 13843 11141
rect 13809 11107 13843 11115
rect 13809 11047 13843 11069
rect 13809 11035 13843 11047
rect 13809 10979 13843 10997
rect 13809 10963 13843 10979
rect 13809 10911 13843 10925
rect 13809 10891 13843 10911
rect 13809 10843 13843 10853
rect 13809 10819 13843 10843
rect 13809 10775 13843 10781
rect 13809 10747 13843 10775
rect 13809 10707 13843 10709
rect 13809 10675 13843 10707
rect 13809 10605 13843 10637
rect 13809 10603 13843 10605
rect 13809 10537 13843 10565
rect 13809 10531 13843 10537
rect 13809 10469 13843 10493
rect 13809 10459 13843 10469
rect 13809 10401 13843 10421
rect 13809 10387 13843 10401
rect 1298 10244 1302 10278
rect 1302 10244 1332 10278
rect 1370 10244 1404 10278
rect 1442 10244 1472 10278
rect 1472 10244 1476 10278
rect 1514 10244 1540 10278
rect 1540 10244 1548 10278
rect 1586 10244 1608 10278
rect 1608 10244 1620 10278
rect 1658 10244 1676 10278
rect 1676 10244 1692 10278
rect 1730 10244 1744 10278
rect 1744 10244 1764 10278
rect 1802 10244 1812 10278
rect 1812 10244 1836 10278
rect 1874 10244 1880 10278
rect 1880 10244 1908 10278
rect 1946 10244 1948 10278
rect 1948 10244 1980 10278
rect 2018 10244 2050 10278
rect 2050 10244 2052 10278
rect 2090 10244 2118 10278
rect 2118 10244 2124 10278
rect 2162 10244 2186 10278
rect 2186 10244 2196 10278
rect 2234 10244 2254 10278
rect 2254 10244 2268 10278
rect 2306 10244 2322 10278
rect 2322 10244 2340 10278
rect 2378 10244 2390 10278
rect 2390 10244 2412 10278
rect 2450 10244 2458 10278
rect 2458 10244 2484 10278
rect 2522 10244 2526 10278
rect 2526 10244 2556 10278
rect 2594 10244 2628 10278
rect 2666 10244 2696 10278
rect 2696 10244 2700 10278
rect 2738 10244 2764 10278
rect 2764 10244 2772 10278
rect 2810 10244 2832 10278
rect 2832 10244 2844 10278
rect 2882 10244 2900 10278
rect 2900 10244 2916 10278
rect 2954 10244 2968 10278
rect 2968 10244 2988 10278
rect 3026 10244 3036 10278
rect 3036 10244 3060 10278
rect 3098 10244 3104 10278
rect 3104 10244 3132 10278
rect 3170 10244 3172 10278
rect 3172 10244 3204 10278
rect 3242 10244 3274 10278
rect 3274 10244 3276 10278
rect 3314 10244 3342 10278
rect 3342 10244 3348 10278
rect 3386 10244 3410 10278
rect 3410 10244 3420 10278
rect 3458 10244 3478 10278
rect 3478 10244 3492 10278
rect 3530 10244 3546 10278
rect 3546 10244 3564 10278
rect 3602 10244 3614 10278
rect 3614 10244 3636 10278
rect 3674 10244 3682 10278
rect 3682 10244 3708 10278
rect 3746 10244 3750 10278
rect 3750 10244 3780 10278
rect 3818 10244 3852 10278
rect 3890 10244 3920 10278
rect 3920 10244 3924 10278
rect 3962 10244 3988 10278
rect 3988 10244 3996 10278
rect 4034 10244 4056 10278
rect 4056 10244 4068 10278
rect 4106 10244 4124 10278
rect 4124 10244 4140 10278
rect 4178 10244 4192 10278
rect 4192 10244 4212 10278
rect 4250 10244 4260 10278
rect 4260 10244 4284 10278
rect 4322 10244 4328 10278
rect 4328 10244 4356 10278
rect 4394 10244 4396 10278
rect 4396 10244 4428 10278
rect 4466 10244 4498 10278
rect 4498 10244 4500 10278
rect 4538 10244 4566 10278
rect 4566 10244 4572 10278
rect 4610 10244 4634 10278
rect 4634 10244 4644 10278
rect 4682 10244 4702 10278
rect 4702 10244 4716 10278
rect 4754 10244 4770 10278
rect 4770 10244 4788 10278
rect 4826 10244 4838 10278
rect 4838 10244 4860 10278
rect 4898 10244 4906 10278
rect 4906 10244 4932 10278
rect 4970 10244 4974 10278
rect 4974 10244 5004 10278
rect 5042 10244 5076 10278
rect 5114 10244 5144 10278
rect 5144 10244 5148 10278
rect 5186 10244 5212 10278
rect 5212 10244 5220 10278
rect 5258 10244 5280 10278
rect 5280 10244 5292 10278
rect 5330 10244 5348 10278
rect 5348 10244 5364 10278
rect 5402 10244 5416 10278
rect 5416 10244 5436 10278
rect 5474 10244 5484 10278
rect 5484 10244 5508 10278
rect 5546 10244 5552 10278
rect 5552 10244 5580 10278
rect 5618 10244 5620 10278
rect 5620 10244 5652 10278
rect 5690 10244 5722 10278
rect 5722 10244 5724 10278
rect 5762 10244 5790 10278
rect 5790 10244 5796 10278
rect 5834 10244 5858 10278
rect 5858 10244 5868 10278
rect 5906 10244 5926 10278
rect 5926 10244 5940 10278
rect 5978 10244 5994 10278
rect 5994 10244 6012 10278
rect 6050 10244 6062 10278
rect 6062 10244 6084 10278
rect 6122 10244 6130 10278
rect 6130 10244 6156 10278
rect 6194 10244 6198 10278
rect 6198 10244 6228 10278
rect 6266 10244 6300 10278
rect 6338 10244 6368 10278
rect 6368 10244 6372 10278
rect 6410 10244 6436 10278
rect 6436 10244 6444 10278
rect 6482 10244 6504 10278
rect 6504 10244 6516 10278
rect 6554 10244 6572 10278
rect 6572 10244 6588 10278
rect 6626 10244 6640 10278
rect 6640 10244 6660 10278
rect 6698 10244 6708 10278
rect 6708 10244 6732 10278
rect 6770 10244 6776 10278
rect 6776 10244 6804 10278
rect 6842 10244 6844 10278
rect 6844 10244 6876 10278
rect 6914 10244 6946 10278
rect 6946 10244 6948 10278
rect 6986 10244 7014 10278
rect 7014 10244 7020 10278
rect 7058 10244 7082 10278
rect 7082 10244 7092 10278
rect 7130 10244 7150 10278
rect 7150 10244 7164 10278
rect 7202 10244 7218 10278
rect 7218 10244 7236 10278
rect 7274 10244 7286 10278
rect 7286 10244 7308 10278
rect 7346 10244 7354 10278
rect 7354 10244 7380 10278
rect 7418 10244 7422 10278
rect 7422 10244 7452 10278
rect 7490 10244 7524 10278
rect 7562 10244 7592 10278
rect 7592 10244 7596 10278
rect 7634 10244 7660 10278
rect 7660 10244 7668 10278
rect 7706 10244 7728 10278
rect 7728 10244 7740 10278
rect 7778 10244 7796 10278
rect 7796 10244 7812 10278
rect 7850 10244 7864 10278
rect 7864 10244 7884 10278
rect 7922 10244 7932 10278
rect 7932 10244 7956 10278
rect 7994 10244 8000 10278
rect 8000 10244 8028 10278
rect 8066 10244 8068 10278
rect 8068 10244 8100 10278
rect 8138 10244 8170 10278
rect 8170 10244 8172 10278
rect 8210 10244 8238 10278
rect 8238 10244 8244 10278
rect 8282 10244 8306 10278
rect 8306 10244 8316 10278
rect 8354 10244 8374 10278
rect 8374 10244 8388 10278
rect 8426 10244 8442 10278
rect 8442 10244 8460 10278
rect 8498 10244 8510 10278
rect 8510 10244 8532 10278
rect 8570 10244 8578 10278
rect 8578 10244 8604 10278
rect 8642 10244 8646 10278
rect 8646 10244 8676 10278
rect 8714 10244 8748 10278
rect 8786 10244 8816 10278
rect 8816 10244 8820 10278
rect 8858 10244 8884 10278
rect 8884 10244 8892 10278
rect 8930 10244 8952 10278
rect 8952 10244 8964 10278
rect 9002 10244 9020 10278
rect 9020 10244 9036 10278
rect 9074 10244 9088 10278
rect 9088 10244 9108 10278
rect 9146 10244 9156 10278
rect 9156 10244 9180 10278
rect 9218 10244 9224 10278
rect 9224 10244 9252 10278
rect 9290 10244 9292 10278
rect 9292 10244 9324 10278
rect 9362 10244 9394 10278
rect 9394 10244 9396 10278
rect 9434 10244 9462 10278
rect 9462 10244 9468 10278
rect 9506 10244 9530 10278
rect 9530 10244 9540 10278
rect 9578 10244 9598 10278
rect 9598 10244 9612 10278
rect 9650 10244 9666 10278
rect 9666 10244 9684 10278
rect 9722 10244 9734 10278
rect 9734 10244 9756 10278
rect 9794 10244 9802 10278
rect 9802 10244 9828 10278
rect 9866 10244 9870 10278
rect 9870 10244 9900 10278
rect 9938 10244 9972 10278
rect 10010 10244 10040 10278
rect 10040 10244 10044 10278
rect 10082 10244 10108 10278
rect 10108 10244 10116 10278
rect 10154 10244 10176 10278
rect 10176 10244 10188 10278
rect 10226 10244 10244 10278
rect 10244 10244 10260 10278
rect 10298 10244 10312 10278
rect 10312 10244 10332 10278
rect 10370 10244 10380 10278
rect 10380 10244 10404 10278
rect 10442 10244 10448 10278
rect 10448 10244 10476 10278
rect 10514 10244 10516 10278
rect 10516 10244 10548 10278
rect 10586 10244 10618 10278
rect 10618 10244 10620 10278
rect 10658 10244 10686 10278
rect 10686 10244 10692 10278
rect 10730 10244 10754 10278
rect 10754 10244 10764 10278
rect 10802 10244 10822 10278
rect 10822 10244 10836 10278
rect 10874 10244 10890 10278
rect 10890 10244 10908 10278
rect 10946 10244 10958 10278
rect 10958 10244 10980 10278
rect 11018 10244 11026 10278
rect 11026 10244 11052 10278
rect 11090 10244 11094 10278
rect 11094 10244 11124 10278
rect 11162 10244 11196 10278
rect 11234 10244 11264 10278
rect 11264 10244 11268 10278
rect 11306 10244 11332 10278
rect 11332 10244 11340 10278
rect 11378 10244 11400 10278
rect 11400 10244 11412 10278
rect 11450 10244 11468 10278
rect 11468 10244 11484 10278
rect 11522 10244 11536 10278
rect 11536 10244 11556 10278
rect 11594 10244 11604 10278
rect 11604 10244 11628 10278
rect 11666 10244 11672 10278
rect 11672 10244 11700 10278
rect 11738 10244 11740 10278
rect 11740 10244 11772 10278
rect 11810 10244 11842 10278
rect 11842 10244 11844 10278
rect 11882 10244 11910 10278
rect 11910 10244 11916 10278
rect 11954 10244 11978 10278
rect 11978 10244 11988 10278
rect 12026 10244 12046 10278
rect 12046 10244 12060 10278
rect 12098 10244 12114 10278
rect 12114 10244 12132 10278
rect 12170 10244 12182 10278
rect 12182 10244 12204 10278
rect 12242 10244 12250 10278
rect 12250 10244 12276 10278
rect 12314 10244 12318 10278
rect 12318 10244 12348 10278
rect 12386 10244 12420 10278
rect 12458 10244 12488 10278
rect 12488 10244 12492 10278
rect 12530 10244 12556 10278
rect 12556 10244 12564 10278
rect 12602 10244 12624 10278
rect 12624 10244 12636 10278
rect 12674 10244 12692 10278
rect 12692 10244 12708 10278
rect 12746 10244 12760 10278
rect 12760 10244 12780 10278
rect 12818 10244 12828 10278
rect 12828 10244 12852 10278
rect 12890 10244 12896 10278
rect 12896 10244 12924 10278
rect 12962 10244 12964 10278
rect 12964 10244 12996 10278
rect 13034 10244 13066 10278
rect 13066 10244 13068 10278
rect 13106 10244 13134 10278
rect 13134 10244 13140 10278
rect 13178 10244 13202 10278
rect 13202 10244 13212 10278
rect 13250 10244 13270 10278
rect 13270 10244 13284 10278
rect 13322 10244 13338 10278
rect 13338 10244 13356 10278
rect 13394 10244 13406 10278
rect 13406 10244 13428 10278
rect 13466 10244 13474 10278
rect 13474 10244 13500 10278
rect 13538 10244 13542 10278
rect 13542 10244 13572 10278
rect 13610 10244 13644 10278
rect 13682 10244 13712 10278
rect 13712 10244 13716 10278
rect 14122 34691 14156 34725
rect 14122 34619 14156 34653
rect 14122 34547 14156 34581
rect 14122 34475 14156 34509
rect 14122 34403 14156 34437
rect 14122 34331 14156 34365
rect 14122 34259 14156 34293
rect 14122 34187 14156 34221
rect 14122 34115 14156 34149
rect 14122 34043 14156 34077
rect 14122 33971 14156 34005
rect 14122 33899 14156 33933
rect 14122 33827 14156 33861
rect 14122 33755 14156 33789
rect 14122 33683 14156 33717
rect 14122 33611 14156 33645
rect 14122 33539 14156 33573
rect 14122 33467 14156 33501
rect 14122 33395 14156 33429
rect 14122 33323 14156 33357
rect 14122 33251 14156 33285
rect 14122 33179 14156 33213
rect 14122 33107 14156 33141
rect 14122 33035 14156 33069
rect 14122 32963 14156 32997
rect 14122 32891 14156 32925
rect 14122 32819 14156 32853
rect 14122 32747 14156 32781
rect 14122 32675 14156 32709
rect 14122 32603 14156 32637
rect 14122 32531 14156 32565
rect 14122 32459 14156 32493
rect 14122 32387 14156 32421
rect 14122 32315 14156 32349
rect 14122 32243 14156 32277
rect 14122 32171 14156 32205
rect 14122 32099 14156 32133
rect 14122 32027 14156 32061
rect 14122 31955 14156 31989
rect 14122 31883 14156 31917
rect 14122 31811 14156 31845
rect 14122 31739 14156 31773
rect 14122 31667 14156 31701
rect 14122 31595 14156 31629
rect 14122 31523 14156 31557
rect 14122 31451 14156 31485
rect 14122 31379 14156 31413
rect 14122 31307 14156 31341
rect 14122 31235 14156 31269
rect 14122 31163 14156 31197
rect 14122 31091 14156 31125
rect 14122 31019 14156 31053
rect 14122 30947 14156 30981
rect 14122 30875 14156 30909
rect 14122 30803 14156 30837
rect 14122 30731 14156 30765
rect 14122 30659 14156 30693
rect 14122 30587 14156 30621
rect 14122 30515 14156 30549
rect 14122 30443 14156 30477
rect 14122 30371 14156 30405
rect 14122 30299 14156 30333
rect 14122 30227 14156 30261
rect 14122 30155 14156 30189
rect 14122 30083 14156 30117
rect 14122 30011 14156 30045
rect 14122 29939 14156 29973
rect 14122 29867 14156 29901
rect 14122 29795 14156 29829
rect 14122 29723 14156 29757
rect 14122 29651 14156 29685
rect 14122 29579 14156 29613
rect 14122 29507 14156 29541
rect 14122 29435 14156 29469
rect 14122 29363 14156 29397
rect 14122 29291 14156 29325
rect 14122 29219 14156 29253
rect 14122 29147 14156 29181
rect 14122 29075 14156 29109
rect 14122 29003 14156 29037
rect 14122 28931 14156 28965
rect 14122 28859 14156 28893
rect 14122 28787 14156 28821
rect 14122 28715 14156 28749
rect 14122 28643 14156 28677
rect 14122 28571 14156 28605
rect 14122 28499 14156 28533
rect 14122 28427 14156 28461
rect 14122 28355 14156 28389
rect 14122 28283 14156 28317
rect 14122 28211 14156 28245
rect 14122 28139 14156 28173
rect 14122 28067 14156 28101
rect 14122 27995 14156 28029
rect 14122 27923 14156 27957
rect 14122 27851 14156 27885
rect 14122 27779 14156 27813
rect 14122 27707 14156 27741
rect 14122 27635 14156 27669
rect 14122 27563 14156 27597
rect 14122 27491 14156 27525
rect 14122 27419 14156 27453
rect 14122 27347 14156 27381
rect 14122 27275 14156 27309
rect 14122 27203 14156 27237
rect 14122 27131 14156 27165
rect 14122 27059 14156 27093
rect 14122 26987 14156 27021
rect 14122 26915 14156 26949
rect 14122 26843 14156 26877
rect 14122 26771 14156 26805
rect 14122 26699 14156 26733
rect 14122 26627 14156 26661
rect 14122 26555 14156 26589
rect 14122 26483 14156 26517
rect 14122 26411 14156 26445
rect 14122 26339 14156 26373
rect 14122 26267 14156 26301
rect 14122 26195 14156 26229
rect 14122 26123 14156 26157
rect 14122 26051 14156 26085
rect 14122 25979 14156 26013
rect 14122 25907 14156 25941
rect 14122 25835 14156 25869
rect 14122 25763 14156 25797
rect 14122 25691 14156 25725
rect 14122 25619 14156 25653
rect 14122 25547 14156 25581
rect 14122 25475 14156 25509
rect 14122 25403 14156 25437
rect 14122 25331 14156 25365
rect 14122 25259 14156 25293
rect 14122 25187 14156 25221
rect 14122 25115 14156 25149
rect 14122 25043 14156 25077
rect 14122 24971 14156 25005
rect 14122 24899 14156 24933
rect 14122 24827 14156 24861
rect 14122 24755 14156 24789
rect 14122 24683 14156 24717
rect 14122 24611 14156 24645
rect 14122 24539 14156 24573
rect 14122 24467 14156 24501
rect 14122 24395 14156 24429
rect 14122 24323 14156 24357
rect 14122 24251 14156 24285
rect 14122 24179 14156 24213
rect 14122 24107 14156 24141
rect 14122 24035 14156 24069
rect 14122 23963 14156 23997
rect 14122 23891 14156 23925
rect 14122 23819 14156 23853
rect 14122 23747 14156 23781
rect 14122 23675 14156 23709
rect 14122 23603 14156 23637
rect 14122 23531 14156 23565
rect 14122 23459 14156 23493
rect 14122 23387 14156 23421
rect 14122 23315 14156 23349
rect 14122 23243 14156 23277
rect 14122 23171 14156 23205
rect 14122 23099 14156 23133
rect 14122 23027 14156 23061
rect 14122 22955 14156 22989
rect 14122 22883 14156 22917
rect 14122 22811 14156 22845
rect 14122 22739 14156 22773
rect 14122 22667 14156 22701
rect 14122 22595 14156 22629
rect 14122 22523 14156 22557
rect 14122 22451 14156 22485
rect 14122 22379 14156 22413
rect 14122 22307 14156 22341
rect 14122 22235 14156 22269
rect 14122 22163 14156 22197
rect 14122 22091 14156 22125
rect 14122 22019 14156 22053
rect 14122 21947 14156 21981
rect 14122 21875 14156 21909
rect 14122 21803 14156 21837
rect 14122 21731 14156 21765
rect 14122 21659 14156 21693
rect 14122 21587 14156 21621
rect 14122 21515 14156 21549
rect 14122 21443 14156 21477
rect 14122 21371 14156 21405
rect 14122 21299 14156 21333
rect 14122 21227 14156 21261
rect 14122 21155 14156 21189
rect 14122 21083 14156 21117
rect 14122 21011 14156 21045
rect 14122 20939 14156 20973
rect 14122 20867 14156 20901
rect 14122 20795 14156 20829
rect 14122 20723 14156 20757
rect 14122 20651 14156 20685
rect 14122 20579 14156 20613
rect 14122 20507 14156 20541
rect 14122 20435 14156 20469
rect 14122 20363 14156 20397
rect 14122 20291 14156 20325
rect 14122 20219 14156 20253
rect 14122 20147 14156 20181
rect 14122 20075 14156 20109
rect 14122 20003 14156 20037
rect 14122 19931 14156 19965
rect 14122 19859 14156 19893
rect 14122 19787 14156 19821
rect 14122 19715 14156 19749
rect 14122 19643 14156 19677
rect 14122 19571 14156 19605
rect 14122 19499 14156 19533
rect 14122 19427 14156 19461
rect 14122 19355 14156 19389
rect 14122 19283 14156 19317
rect 14122 19211 14156 19245
rect 14122 19139 14156 19173
rect 14122 19067 14156 19101
rect 14122 18995 14156 19029
rect 14122 18923 14156 18957
rect 14122 18851 14156 18885
rect 14122 18779 14156 18813
rect 14122 18707 14156 18741
rect 14122 18635 14156 18669
rect 14122 18563 14156 18597
rect 14122 18491 14156 18525
rect 14122 18419 14156 18453
rect 14122 18347 14156 18381
rect 14122 18275 14156 18309
rect 14122 18203 14156 18237
rect 14122 18131 14156 18165
rect 14122 18059 14156 18093
rect 14122 17987 14156 18021
rect 14122 17915 14156 17949
rect 14122 17843 14156 17877
rect 14122 17771 14156 17805
rect 14122 17699 14156 17733
rect 14122 17627 14156 17661
rect 14122 17555 14156 17589
rect 14122 17483 14156 17517
rect 14122 17411 14156 17445
rect 14122 17339 14156 17373
rect 14122 17267 14156 17301
rect 14122 17195 14156 17229
rect 14122 17123 14156 17157
rect 14122 17051 14156 17085
rect 14122 16979 14156 17013
rect 14122 16907 14156 16941
rect 14122 16835 14156 16869
rect 14122 16763 14156 16797
rect 14122 16691 14156 16725
rect 14122 16619 14156 16653
rect 14122 16547 14156 16581
rect 14122 16475 14156 16509
rect 14122 16403 14156 16437
rect 14122 16331 14156 16365
rect 14122 16259 14156 16293
rect 14122 16187 14156 16221
rect 14122 16115 14156 16149
rect 14122 16043 14156 16077
rect 14122 15971 14156 16005
rect 14122 15899 14156 15933
rect 14122 15827 14156 15861
rect 14122 15755 14156 15789
rect 14122 15683 14156 15717
rect 14122 15611 14156 15645
rect 14122 15539 14156 15573
rect 14122 15467 14156 15501
rect 14122 15395 14156 15429
rect 14122 15323 14156 15357
rect 14122 15251 14156 15285
rect 14122 15179 14156 15213
rect 14122 15107 14156 15141
rect 14122 15035 14156 15069
rect 14122 14963 14156 14997
rect 14122 14891 14156 14925
rect 14122 14819 14156 14853
rect 14122 14747 14156 14781
rect 14122 14675 14156 14709
rect 14122 14603 14156 14637
rect 14122 14531 14156 14565
rect 14122 14459 14156 14493
rect 14122 14387 14156 14421
rect 14122 14315 14156 14349
rect 14122 14243 14156 14277
rect 14122 14171 14156 14205
rect 14122 14099 14156 14133
rect 14122 14027 14156 14061
rect 14122 13955 14156 13989
rect 14122 13883 14156 13917
rect 14122 13811 14156 13845
rect 14122 13739 14156 13773
rect 14122 13667 14156 13701
rect 14122 13595 14156 13629
rect 14122 13523 14156 13557
rect 14122 13451 14156 13485
rect 14122 13379 14156 13413
rect 14122 13307 14156 13341
rect 14122 13235 14156 13269
rect 14122 13163 14156 13197
rect 14122 13091 14156 13125
rect 14122 13019 14156 13053
rect 14122 12947 14156 12981
rect 14122 12875 14156 12909
rect 14122 12803 14156 12837
rect 14122 12731 14156 12765
rect 14122 12659 14156 12693
rect 14122 12587 14156 12621
rect 14122 12515 14156 12549
rect 14122 12443 14156 12477
rect 14122 12371 14156 12405
rect 14122 12299 14156 12333
rect 14122 12227 14156 12261
rect 14122 12155 14156 12189
rect 14122 12083 14156 12117
rect 14122 12011 14156 12045
rect 14122 11939 14156 11973
rect 14122 11867 14156 11901
rect 14122 11795 14156 11829
rect 14122 11723 14156 11757
rect 14122 11651 14156 11685
rect 14122 11579 14156 11613
rect 14122 11507 14156 11541
rect 14122 11435 14156 11469
rect 14122 11363 14156 11397
rect 14122 11291 14156 11325
rect 14122 11219 14156 11253
rect 14122 11147 14156 11181
rect 14122 11075 14156 11109
rect 14122 11003 14156 11037
rect 14122 10931 14156 10965
rect 14122 10859 14156 10893
rect 14122 10787 14156 10821
rect 14122 10715 14156 10749
rect 14122 10643 14156 10677
rect 14122 10571 14156 10605
rect 14122 10499 14156 10533
rect 14122 10427 14156 10461
rect 14122 10355 14156 10389
rect 14122 10283 14156 10317
rect 14122 10211 14156 10245
rect 807 10146 841 10180
rect 807 10074 841 10108
rect 14122 10139 14156 10173
rect 14122 10067 14156 10101
rect 891 9908 925 9942
rect 963 9908 997 9942
rect 1035 9908 1069 9942
rect 1107 9908 1141 9942
rect 1179 9908 1213 9942
rect 1251 9908 1285 9942
rect 1323 9908 1357 9942
rect 1395 9908 1429 9942
rect 1467 9908 1501 9942
rect 1539 9908 1573 9942
rect 1611 9908 1645 9942
rect 1683 9908 1717 9942
rect 1755 9908 1789 9942
rect 1827 9908 1861 9942
rect 1899 9908 1933 9942
rect 1971 9908 2005 9942
rect 2043 9908 2077 9942
rect 2115 9908 2149 9942
rect 2187 9908 2221 9942
rect 2259 9908 2293 9942
rect 2331 9908 2365 9942
rect 2403 9908 2437 9942
rect 2475 9908 2509 9942
rect 2547 9908 2581 9942
rect 2619 9908 2653 9942
rect 2691 9908 2725 9942
rect 2763 9908 2797 9942
rect 2835 9908 2869 9942
rect 2907 9908 2941 9942
rect 2979 9908 3013 9942
rect 3051 9908 3085 9942
rect 3123 9908 3157 9942
rect 3195 9908 3229 9942
rect 3267 9908 3301 9942
rect 3339 9908 3373 9942
rect 3411 9908 3445 9942
rect 3483 9908 3517 9942
rect 3555 9908 3589 9942
rect 3627 9908 3661 9942
rect 3699 9908 3733 9942
rect 3771 9908 3805 9942
rect 3843 9908 3877 9942
rect 3915 9908 3949 9942
rect 3987 9908 4021 9942
rect 4059 9908 4093 9942
rect 4131 9908 4165 9942
rect 4203 9908 4237 9942
rect 4275 9908 4309 9942
rect 4347 9908 4381 9942
rect 4419 9908 4453 9942
rect 4491 9908 4525 9942
rect 4563 9908 4597 9942
rect 4635 9908 4669 9942
rect 4707 9908 4741 9942
rect 4779 9908 4813 9942
rect 4851 9908 4885 9942
rect 4923 9908 4957 9942
rect 4995 9908 5029 9942
rect 5067 9908 5101 9942
rect 5139 9908 5173 9942
rect 5211 9908 5245 9942
rect 5283 9908 5317 9942
rect 5355 9908 5389 9942
rect 5427 9908 5461 9942
rect 5499 9908 5533 9942
rect 5571 9908 5605 9942
rect 5643 9908 5677 9942
rect 5715 9908 5749 9942
rect 5787 9908 5821 9942
rect 5859 9908 5893 9942
rect 5931 9908 5965 9942
rect 6003 9908 6037 9942
rect 6075 9908 6109 9942
rect 6147 9908 6181 9942
rect 6219 9908 6253 9942
rect 6291 9908 6325 9942
rect 6363 9908 6397 9942
rect 6435 9908 6469 9942
rect 6507 9908 6541 9942
rect 6579 9908 6613 9942
rect 6651 9908 6685 9942
rect 6723 9908 6757 9942
rect 6795 9908 6829 9942
rect 6867 9908 6901 9942
rect 6939 9908 6973 9942
rect 7011 9908 7045 9942
rect 7083 9908 7117 9942
rect 7155 9908 7189 9942
rect 7227 9908 7261 9942
rect 7299 9908 7333 9942
rect 7371 9908 7405 9942
rect 7443 9908 7477 9942
rect 7515 9908 7549 9942
rect 7587 9908 7621 9942
rect 7659 9908 7693 9942
rect 7731 9908 7765 9942
rect 7803 9908 7837 9942
rect 7875 9908 7909 9942
rect 7947 9908 7981 9942
rect 8019 9908 8053 9942
rect 8091 9908 8125 9942
rect 8163 9908 8197 9942
rect 8235 9908 8269 9942
rect 8307 9908 8341 9942
rect 8379 9908 8413 9942
rect 8451 9908 8485 9942
rect 8523 9908 8557 9942
rect 8595 9908 8629 9942
rect 8667 9908 8701 9942
rect 8739 9908 8773 9942
rect 8811 9908 8845 9942
rect 8883 9908 8917 9942
rect 8955 9908 8989 9942
rect 9027 9908 9061 9942
rect 9099 9908 9133 9942
rect 9171 9908 9205 9942
rect 9243 9908 9277 9942
rect 9315 9908 9349 9942
rect 9387 9908 9421 9942
rect 9459 9908 9493 9942
rect 9531 9908 9565 9942
rect 9603 9908 9637 9942
rect 9675 9908 9709 9942
rect 9747 9908 9781 9942
rect 9819 9908 9853 9942
rect 9891 9908 9925 9942
rect 9963 9908 9997 9942
rect 10035 9908 10069 9942
rect 10107 9908 10141 9942
rect 10179 9908 10213 9942
rect 10251 9908 10285 9942
rect 10323 9908 10357 9942
rect 10395 9908 10429 9942
rect 10467 9908 10501 9942
rect 10539 9908 10573 9942
rect 10611 9908 10645 9942
rect 10683 9908 10717 9942
rect 10755 9908 10789 9942
rect 10827 9908 10861 9942
rect 10899 9908 10933 9942
rect 10971 9908 11005 9942
rect 11043 9908 11077 9942
rect 11115 9908 11149 9942
rect 11187 9908 11221 9942
rect 11259 9908 11293 9942
rect 11331 9908 11365 9942
rect 11403 9908 11437 9942
rect 11475 9908 11509 9942
rect 11547 9908 11581 9942
rect 11619 9908 11653 9942
rect 11691 9908 11725 9942
rect 11763 9908 11797 9942
rect 11835 9908 11869 9942
rect 11907 9908 11941 9942
rect 11979 9908 12013 9942
rect 12051 9908 12085 9942
rect 12123 9908 12157 9942
rect 12195 9908 12229 9942
rect 12267 9908 12301 9942
rect 12339 9908 12373 9942
rect 12411 9908 12445 9942
rect 12483 9908 12517 9942
rect 12555 9908 12589 9942
rect 12627 9908 12661 9942
rect 12699 9908 12733 9942
rect 12771 9908 12805 9942
rect 12843 9908 12877 9942
rect 12915 9908 12949 9942
rect 12987 9908 13021 9942
rect 13059 9908 13093 9942
rect 13131 9908 13165 9942
rect 13203 9908 13237 9942
rect 13275 9908 13309 9942
rect 13347 9908 13381 9942
rect 13419 9908 13453 9942
rect 13491 9908 13525 9942
rect 13563 9908 13597 9942
rect 13635 9908 13669 9942
rect 13707 9908 13741 9942
rect 13779 9908 13813 9942
rect 13851 9908 13885 9942
rect 13923 9908 13957 9942
rect 13995 9908 14029 9942
rect 883 9741 902 9774
rect 902 9741 917 9774
rect 955 9741 970 9774
rect 970 9741 989 9774
rect 1027 9741 1038 9774
rect 1038 9741 1061 9774
rect 1099 9741 1106 9774
rect 1106 9741 1133 9774
rect 1171 9741 1174 9774
rect 1174 9741 1205 9774
rect 1243 9741 1276 9774
rect 1276 9741 1277 9774
rect 1315 9741 1344 9774
rect 1344 9741 1349 9774
rect 1387 9741 1412 9774
rect 1412 9741 1421 9774
rect 1459 9741 1480 9774
rect 1480 9741 1493 9774
rect 1531 9741 1548 9774
rect 1548 9741 1565 9774
rect 1603 9741 1616 9774
rect 1616 9741 1637 9774
rect 1675 9741 1684 9774
rect 1684 9741 1709 9774
rect 1747 9741 1752 9774
rect 1752 9741 1781 9774
rect 1819 9741 1820 9774
rect 1820 9741 1853 9774
rect 1891 9741 1922 9774
rect 1922 9741 1925 9774
rect 1963 9741 1990 9774
rect 1990 9741 1997 9774
rect 2035 9741 2058 9774
rect 2058 9741 2069 9774
rect 12883 9741 12904 9774
rect 12904 9741 12917 9774
rect 12955 9741 12972 9774
rect 12972 9741 12989 9774
rect 13027 9741 13040 9774
rect 13040 9741 13061 9774
rect 13099 9741 13108 9774
rect 13108 9741 13133 9774
rect 13171 9741 13176 9774
rect 13176 9741 13205 9774
rect 13243 9741 13244 9774
rect 13244 9741 13277 9774
rect 13315 9741 13346 9774
rect 13346 9741 13349 9774
rect 13387 9741 13414 9774
rect 13414 9741 13421 9774
rect 13459 9741 13482 9774
rect 13482 9741 13493 9774
rect 13531 9741 13550 9774
rect 13550 9741 13565 9774
rect 13603 9741 13618 9774
rect 13618 9741 13637 9774
rect 13675 9741 13686 9774
rect 13686 9741 13709 9774
rect 13747 9741 13754 9774
rect 13754 9741 13781 9774
rect 13819 9741 13822 9774
rect 13822 9741 13853 9774
rect 13891 9741 13924 9774
rect 13924 9741 13925 9774
rect 13963 9741 13992 9774
rect 13992 9741 13997 9774
rect 14035 9741 14060 9774
rect 14060 9741 14069 9774
rect 883 9740 917 9741
rect 955 9740 989 9741
rect 1027 9740 1061 9741
rect 1099 9740 1133 9741
rect 1171 9740 1205 9741
rect 1243 9740 1277 9741
rect 1315 9740 1349 9741
rect 1387 9740 1421 9741
rect 1459 9740 1493 9741
rect 1531 9740 1565 9741
rect 1603 9740 1637 9741
rect 1675 9740 1709 9741
rect 1747 9740 1781 9741
rect 1819 9740 1853 9741
rect 1891 9740 1925 9741
rect 1963 9740 1997 9741
rect 2035 9740 2069 9741
rect 12883 9740 12917 9741
rect 12955 9740 12989 9741
rect 13027 9740 13061 9741
rect 13099 9740 13133 9741
rect 13171 9740 13205 9741
rect 13243 9740 13277 9741
rect 13315 9740 13349 9741
rect 13387 9740 13421 9741
rect 13459 9740 13493 9741
rect 13531 9740 13565 9741
rect 13603 9740 13637 9741
rect 13675 9740 13709 9741
rect 13747 9740 13781 9741
rect 13819 9740 13853 9741
rect 13891 9740 13925 9741
rect 13963 9740 13997 9741
rect 14035 9740 14069 9741
rect 14614 36174 14641 36190
rect 14641 36174 14648 36190
rect 14614 36156 14648 36174
rect 14614 36106 14641 36118
rect 14641 36106 14648 36118
rect 14614 36084 14648 36106
rect 14614 36038 14641 36046
rect 14641 36038 14648 36046
rect 14614 36012 14648 36038
rect 14614 35970 14641 35974
rect 14641 35970 14648 35974
rect 14614 35940 14648 35970
rect 14614 35868 14648 35902
rect 14614 35800 14648 35830
rect 14614 35796 14641 35800
rect 14641 35796 14648 35800
rect 14614 35732 14648 35758
rect 14614 35724 14641 35732
rect 14641 35724 14648 35732
rect 14614 35664 14648 35686
rect 14614 35652 14641 35664
rect 14641 35652 14648 35664
rect 14614 35596 14648 35614
rect 14614 35580 14641 35596
rect 14641 35580 14648 35596
rect 14614 35528 14648 35542
rect 14614 35508 14641 35528
rect 14641 35508 14648 35528
rect 14614 35460 14648 35470
rect 14614 35436 14641 35460
rect 14641 35436 14648 35460
rect 14614 35392 14648 35398
rect 14614 35364 14641 35392
rect 14641 35364 14648 35392
rect 14614 35324 14648 35326
rect 14614 35292 14641 35324
rect 14641 35292 14648 35324
rect 14614 35222 14641 35254
rect 14641 35222 14648 35254
rect 14614 35220 14648 35222
rect 14614 35154 14641 35182
rect 14641 35154 14648 35182
rect 14614 35148 14648 35154
rect 14614 35086 14641 35110
rect 14641 35086 14648 35110
rect 14614 35076 14648 35086
rect 14614 35018 14641 35038
rect 14641 35018 14648 35038
rect 14614 35004 14648 35018
rect 14614 34950 14641 34966
rect 14641 34950 14648 34966
rect 14614 34932 14648 34950
rect 14614 34882 14641 34894
rect 14641 34882 14648 34894
rect 14614 34860 14648 34882
rect 14614 34814 14641 34822
rect 14641 34814 14648 34822
rect 14614 34788 14648 34814
rect 14614 34746 14641 34750
rect 14641 34746 14648 34750
rect 14614 34716 14648 34746
rect 14614 34644 14648 34678
rect 14614 34576 14648 34606
rect 14614 34572 14641 34576
rect 14641 34572 14648 34576
rect 14614 34508 14648 34534
rect 14614 34500 14641 34508
rect 14641 34500 14648 34508
rect 14614 34440 14648 34462
rect 14614 34428 14641 34440
rect 14641 34428 14648 34440
rect 14614 34372 14648 34390
rect 14614 34356 14641 34372
rect 14641 34356 14648 34372
rect 14614 34304 14648 34318
rect 14614 34284 14641 34304
rect 14641 34284 14648 34304
rect 14614 34236 14648 34246
rect 14614 34212 14641 34236
rect 14641 34212 14648 34236
rect 14614 34168 14648 34174
rect 14614 34140 14641 34168
rect 14641 34140 14648 34168
rect 14614 34100 14648 34102
rect 14614 34068 14641 34100
rect 14641 34068 14648 34100
rect 14614 33998 14641 34030
rect 14641 33998 14648 34030
rect 14614 33996 14648 33998
rect 14614 33930 14641 33958
rect 14641 33930 14648 33958
rect 14614 33924 14648 33930
rect 14614 33862 14641 33886
rect 14641 33862 14648 33886
rect 14614 33852 14648 33862
rect 14614 33794 14641 33814
rect 14641 33794 14648 33814
rect 14614 33780 14648 33794
rect 14614 33726 14641 33742
rect 14641 33726 14648 33742
rect 14614 33708 14648 33726
rect 14614 33658 14641 33670
rect 14641 33658 14648 33670
rect 14614 33636 14648 33658
rect 14614 33590 14641 33598
rect 14641 33590 14648 33598
rect 14614 33564 14648 33590
rect 14614 33522 14641 33526
rect 14641 33522 14648 33526
rect 14614 33492 14648 33522
rect 14614 33420 14648 33454
rect 14614 33352 14648 33382
rect 14614 33348 14641 33352
rect 14641 33348 14648 33352
rect 14614 33284 14648 33310
rect 14614 33276 14641 33284
rect 14641 33276 14648 33284
rect 14614 33216 14648 33238
rect 14614 33204 14641 33216
rect 14641 33204 14648 33216
rect 14614 33148 14648 33166
rect 14614 33132 14641 33148
rect 14641 33132 14648 33148
rect 14614 33080 14648 33094
rect 14614 33060 14641 33080
rect 14641 33060 14648 33080
rect 14614 33012 14648 33022
rect 14614 32988 14641 33012
rect 14641 32988 14648 33012
rect 14614 32944 14648 32950
rect 14614 32916 14641 32944
rect 14641 32916 14648 32944
rect 14614 32876 14648 32878
rect 14614 32844 14641 32876
rect 14641 32844 14648 32876
rect 14614 32774 14641 32806
rect 14641 32774 14648 32806
rect 14614 32772 14648 32774
rect 14614 32706 14641 32734
rect 14641 32706 14648 32734
rect 14614 32700 14648 32706
rect 14614 32638 14641 32662
rect 14641 32638 14648 32662
rect 14614 32628 14648 32638
rect 14614 32570 14641 32590
rect 14641 32570 14648 32590
rect 14614 32556 14648 32570
rect 14614 32502 14641 32518
rect 14641 32502 14648 32518
rect 14614 32484 14648 32502
rect 14614 32434 14641 32446
rect 14641 32434 14648 32446
rect 14614 32412 14648 32434
rect 14614 32366 14641 32374
rect 14641 32366 14648 32374
rect 14614 32340 14648 32366
rect 14614 32298 14641 32302
rect 14641 32298 14648 32302
rect 14614 32268 14648 32298
rect 14614 32196 14648 32230
rect 14614 32128 14648 32158
rect 14614 32124 14641 32128
rect 14641 32124 14648 32128
rect 14614 32060 14648 32086
rect 14614 32052 14641 32060
rect 14641 32052 14648 32060
rect 14614 31992 14648 32014
rect 14614 31980 14641 31992
rect 14641 31980 14648 31992
rect 14614 31924 14648 31942
rect 14614 31908 14641 31924
rect 14641 31908 14648 31924
rect 14614 31856 14648 31870
rect 14614 31836 14641 31856
rect 14641 31836 14648 31856
rect 14614 31788 14648 31798
rect 14614 31764 14641 31788
rect 14641 31764 14648 31788
rect 14614 31720 14648 31726
rect 14614 31692 14641 31720
rect 14641 31692 14648 31720
rect 14614 31652 14648 31654
rect 14614 31620 14641 31652
rect 14641 31620 14648 31652
rect 14614 31550 14641 31582
rect 14641 31550 14648 31582
rect 14614 31548 14648 31550
rect 14614 31482 14641 31510
rect 14641 31482 14648 31510
rect 14614 31476 14648 31482
rect 14614 31414 14641 31438
rect 14641 31414 14648 31438
rect 14614 31404 14648 31414
rect 14614 31346 14641 31366
rect 14641 31346 14648 31366
rect 14614 31332 14648 31346
rect 14614 31278 14641 31294
rect 14641 31278 14648 31294
rect 14614 31260 14648 31278
rect 14614 31210 14641 31222
rect 14641 31210 14648 31222
rect 14614 31188 14648 31210
rect 14614 31142 14641 31150
rect 14641 31142 14648 31150
rect 14614 31116 14648 31142
rect 14614 31074 14641 31078
rect 14641 31074 14648 31078
rect 14614 31044 14648 31074
rect 14614 30972 14648 31006
rect 14614 30904 14648 30934
rect 14614 30900 14641 30904
rect 14641 30900 14648 30904
rect 14614 30836 14648 30862
rect 14614 30828 14641 30836
rect 14641 30828 14648 30836
rect 14614 30768 14648 30790
rect 14614 30756 14641 30768
rect 14641 30756 14648 30768
rect 14614 30700 14648 30718
rect 14614 30684 14641 30700
rect 14641 30684 14648 30700
rect 14614 30632 14648 30646
rect 14614 30612 14641 30632
rect 14641 30612 14648 30632
rect 14614 30564 14648 30574
rect 14614 30540 14641 30564
rect 14641 30540 14648 30564
rect 14614 30496 14648 30502
rect 14614 30468 14641 30496
rect 14641 30468 14648 30496
rect 14614 30428 14648 30430
rect 14614 30396 14641 30428
rect 14641 30396 14648 30428
rect 14614 30326 14641 30358
rect 14641 30326 14648 30358
rect 14614 30324 14648 30326
rect 14614 30258 14641 30286
rect 14641 30258 14648 30286
rect 14614 30252 14648 30258
rect 14614 30190 14641 30214
rect 14641 30190 14648 30214
rect 14614 30180 14648 30190
rect 14614 30122 14641 30142
rect 14641 30122 14648 30142
rect 14614 30108 14648 30122
rect 14614 30054 14641 30070
rect 14641 30054 14648 30070
rect 14614 30036 14648 30054
rect 14614 29986 14641 29998
rect 14641 29986 14648 29998
rect 14614 29964 14648 29986
rect 14614 29918 14641 29926
rect 14641 29918 14648 29926
rect 14614 29892 14648 29918
rect 14614 29850 14641 29854
rect 14641 29850 14648 29854
rect 14614 29820 14648 29850
rect 14614 29748 14648 29782
rect 14614 29680 14648 29710
rect 14614 29676 14641 29680
rect 14641 29676 14648 29680
rect 14614 29612 14648 29638
rect 14614 29604 14641 29612
rect 14641 29604 14648 29612
rect 14614 29544 14648 29566
rect 14614 29532 14641 29544
rect 14641 29532 14648 29544
rect 14614 29476 14648 29494
rect 14614 29460 14641 29476
rect 14641 29460 14648 29476
rect 14614 29408 14648 29422
rect 14614 29388 14641 29408
rect 14641 29388 14648 29408
rect 14614 29340 14648 29350
rect 14614 29316 14641 29340
rect 14641 29316 14648 29340
rect 14614 29272 14648 29278
rect 14614 29244 14641 29272
rect 14641 29244 14648 29272
rect 14614 29204 14648 29206
rect 14614 29172 14641 29204
rect 14641 29172 14648 29204
rect 14614 29102 14641 29134
rect 14641 29102 14648 29134
rect 14614 29100 14648 29102
rect 14614 29034 14641 29062
rect 14641 29034 14648 29062
rect 14614 29028 14648 29034
rect 14614 28966 14641 28990
rect 14641 28966 14648 28990
rect 14614 28956 14648 28966
rect 14614 28898 14641 28918
rect 14641 28898 14648 28918
rect 14614 28884 14648 28898
rect 14614 28830 14641 28846
rect 14641 28830 14648 28846
rect 14614 28812 14648 28830
rect 14614 28762 14641 28774
rect 14641 28762 14648 28774
rect 14614 28740 14648 28762
rect 14614 28694 14641 28702
rect 14641 28694 14648 28702
rect 14614 28668 14648 28694
rect 14614 28626 14641 28630
rect 14641 28626 14648 28630
rect 14614 28596 14648 28626
rect 14614 28524 14648 28558
rect 14614 28456 14648 28486
rect 14614 28452 14641 28456
rect 14641 28452 14648 28456
rect 14614 28388 14648 28414
rect 14614 28380 14641 28388
rect 14641 28380 14648 28388
rect 14614 28320 14648 28342
rect 14614 28308 14641 28320
rect 14641 28308 14648 28320
rect 14614 28252 14648 28270
rect 14614 28236 14641 28252
rect 14641 28236 14648 28252
rect 14614 28184 14648 28198
rect 14614 28164 14641 28184
rect 14641 28164 14648 28184
rect 14614 28116 14648 28126
rect 14614 28092 14641 28116
rect 14641 28092 14648 28116
rect 14614 28048 14648 28054
rect 14614 28020 14641 28048
rect 14641 28020 14648 28048
rect 14614 27980 14648 27982
rect 14614 27948 14641 27980
rect 14641 27948 14648 27980
rect 14614 27878 14641 27910
rect 14641 27878 14648 27910
rect 14614 27876 14648 27878
rect 14614 27810 14641 27838
rect 14641 27810 14648 27838
rect 14614 27804 14648 27810
rect 14614 27742 14641 27766
rect 14641 27742 14648 27766
rect 14614 27732 14648 27742
rect 14614 27674 14641 27694
rect 14641 27674 14648 27694
rect 14614 27660 14648 27674
rect 14614 27606 14641 27622
rect 14641 27606 14648 27622
rect 14614 27588 14648 27606
rect 14614 27538 14641 27550
rect 14641 27538 14648 27550
rect 14614 27516 14648 27538
rect 14614 27470 14641 27478
rect 14641 27470 14648 27478
rect 14614 27444 14648 27470
rect 14614 27402 14641 27406
rect 14641 27402 14648 27406
rect 14614 27372 14648 27402
rect 14614 27300 14648 27334
rect 14614 27232 14648 27262
rect 14614 27228 14641 27232
rect 14641 27228 14648 27232
rect 14614 27164 14648 27190
rect 14614 27156 14641 27164
rect 14641 27156 14648 27164
rect 14614 27096 14648 27118
rect 14614 27084 14641 27096
rect 14641 27084 14648 27096
rect 14614 27028 14648 27046
rect 14614 27012 14641 27028
rect 14641 27012 14648 27028
rect 14614 26960 14648 26974
rect 14614 26940 14641 26960
rect 14641 26940 14648 26960
rect 14614 26892 14648 26902
rect 14614 26868 14641 26892
rect 14641 26868 14648 26892
rect 14614 26824 14648 26830
rect 14614 26796 14641 26824
rect 14641 26796 14648 26824
rect 14614 26756 14648 26758
rect 14614 26724 14641 26756
rect 14641 26724 14648 26756
rect 14614 26654 14641 26686
rect 14641 26654 14648 26686
rect 14614 26652 14648 26654
rect 14614 26586 14641 26614
rect 14641 26586 14648 26614
rect 14614 26580 14648 26586
rect 14614 26518 14641 26542
rect 14641 26518 14648 26542
rect 14614 26508 14648 26518
rect 14614 26450 14641 26470
rect 14641 26450 14648 26470
rect 14614 26436 14648 26450
rect 14614 26382 14641 26398
rect 14641 26382 14648 26398
rect 14614 26364 14648 26382
rect 14614 26314 14641 26326
rect 14641 26314 14648 26326
rect 14614 26292 14648 26314
rect 14614 26246 14641 26254
rect 14641 26246 14648 26254
rect 14614 26220 14648 26246
rect 14614 26178 14641 26182
rect 14641 26178 14648 26182
rect 14614 26148 14648 26178
rect 14614 26076 14648 26110
rect 14614 26008 14648 26038
rect 14614 26004 14641 26008
rect 14641 26004 14648 26008
rect 14614 25940 14648 25966
rect 14614 25932 14641 25940
rect 14641 25932 14648 25940
rect 14614 25872 14648 25894
rect 14614 25860 14641 25872
rect 14641 25860 14648 25872
rect 14614 25804 14648 25822
rect 14614 25788 14641 25804
rect 14641 25788 14648 25804
rect 14614 25736 14648 25750
rect 14614 25716 14641 25736
rect 14641 25716 14648 25736
rect 14614 25668 14648 25678
rect 14614 25644 14641 25668
rect 14641 25644 14648 25668
rect 14614 25600 14648 25606
rect 14614 25572 14641 25600
rect 14641 25572 14648 25600
rect 14614 25532 14648 25534
rect 14614 25500 14641 25532
rect 14641 25500 14648 25532
rect 14614 25430 14641 25462
rect 14641 25430 14648 25462
rect 14614 25428 14648 25430
rect 14614 25362 14641 25390
rect 14641 25362 14648 25390
rect 14614 25356 14648 25362
rect 14614 25294 14641 25318
rect 14641 25294 14648 25318
rect 14614 25284 14648 25294
rect 14614 25226 14641 25246
rect 14641 25226 14648 25246
rect 14614 25212 14648 25226
rect 14614 25158 14641 25174
rect 14641 25158 14648 25174
rect 14614 25140 14648 25158
rect 14614 25090 14641 25102
rect 14641 25090 14648 25102
rect 14614 25068 14648 25090
rect 14614 25022 14641 25030
rect 14641 25022 14648 25030
rect 14614 24996 14648 25022
rect 14614 24954 14641 24958
rect 14641 24954 14648 24958
rect 14614 24924 14648 24954
rect 14614 24852 14648 24886
rect 14614 24784 14648 24814
rect 14614 24780 14641 24784
rect 14641 24780 14648 24784
rect 14614 24716 14648 24742
rect 14614 24708 14641 24716
rect 14641 24708 14648 24716
rect 14614 24648 14648 24670
rect 14614 24636 14641 24648
rect 14641 24636 14648 24648
rect 14614 24580 14648 24598
rect 14614 24564 14641 24580
rect 14641 24564 14648 24580
rect 14614 24512 14648 24526
rect 14614 24492 14641 24512
rect 14641 24492 14648 24512
rect 14614 24444 14648 24454
rect 14614 24420 14641 24444
rect 14641 24420 14648 24444
rect 14614 24376 14648 24382
rect 14614 24348 14641 24376
rect 14641 24348 14648 24376
rect 14614 24308 14648 24310
rect 14614 24276 14641 24308
rect 14641 24276 14648 24308
rect 14614 24206 14641 24238
rect 14641 24206 14648 24238
rect 14614 24204 14648 24206
rect 14614 24138 14641 24166
rect 14641 24138 14648 24166
rect 14614 24132 14648 24138
rect 14614 24070 14641 24094
rect 14641 24070 14648 24094
rect 14614 24060 14648 24070
rect 14614 24002 14641 24022
rect 14641 24002 14648 24022
rect 14614 23988 14648 24002
rect 14614 23934 14641 23950
rect 14641 23934 14648 23950
rect 14614 23916 14648 23934
rect 14614 23866 14641 23878
rect 14641 23866 14648 23878
rect 14614 23844 14648 23866
rect 14614 23798 14641 23806
rect 14641 23798 14648 23806
rect 14614 23772 14648 23798
rect 14614 23730 14641 23734
rect 14641 23730 14648 23734
rect 14614 23700 14648 23730
rect 14614 23628 14648 23662
rect 14614 23560 14648 23590
rect 14614 23556 14641 23560
rect 14641 23556 14648 23560
rect 14614 23492 14648 23518
rect 14614 23484 14641 23492
rect 14641 23484 14648 23492
rect 14614 23424 14648 23446
rect 14614 23412 14641 23424
rect 14641 23412 14648 23424
rect 14614 23356 14648 23374
rect 14614 23340 14641 23356
rect 14641 23340 14648 23356
rect 14614 23288 14648 23302
rect 14614 23268 14641 23288
rect 14641 23268 14648 23288
rect 14614 23220 14648 23230
rect 14614 23196 14641 23220
rect 14641 23196 14648 23220
rect 14614 23152 14648 23158
rect 14614 23124 14641 23152
rect 14641 23124 14648 23152
rect 14614 23084 14648 23086
rect 14614 23052 14641 23084
rect 14641 23052 14648 23084
rect 14614 22982 14641 23014
rect 14641 22982 14648 23014
rect 14614 22980 14648 22982
rect 14614 22914 14641 22942
rect 14641 22914 14648 22942
rect 14614 22908 14648 22914
rect 14614 22846 14641 22870
rect 14641 22846 14648 22870
rect 14614 22836 14648 22846
rect 14614 22778 14641 22798
rect 14641 22778 14648 22798
rect 14614 22764 14648 22778
rect 14614 22710 14641 22726
rect 14641 22710 14648 22726
rect 14614 22692 14648 22710
rect 14614 22642 14641 22654
rect 14641 22642 14648 22654
rect 14614 22620 14648 22642
rect 14614 22574 14641 22582
rect 14641 22574 14648 22582
rect 14614 22548 14648 22574
rect 14614 22506 14641 22510
rect 14641 22506 14648 22510
rect 14614 22476 14648 22506
rect 14614 22404 14648 22438
rect 14614 22336 14648 22366
rect 14614 22332 14641 22336
rect 14641 22332 14648 22336
rect 14614 22268 14648 22294
rect 14614 22260 14641 22268
rect 14641 22260 14648 22268
rect 14614 22200 14648 22222
rect 14614 22188 14641 22200
rect 14641 22188 14648 22200
rect 14614 22132 14648 22150
rect 14614 22116 14641 22132
rect 14641 22116 14648 22132
rect 14614 22064 14648 22078
rect 14614 22044 14641 22064
rect 14641 22044 14648 22064
rect 14614 21996 14648 22006
rect 14614 21972 14641 21996
rect 14641 21972 14648 21996
rect 14614 21928 14648 21934
rect 14614 21900 14641 21928
rect 14641 21900 14648 21928
rect 14614 21860 14648 21862
rect 14614 21828 14641 21860
rect 14641 21828 14648 21860
rect 14614 21758 14641 21790
rect 14641 21758 14648 21790
rect 14614 21756 14648 21758
rect 14614 21690 14641 21718
rect 14641 21690 14648 21718
rect 14614 21684 14648 21690
rect 14614 21622 14641 21646
rect 14641 21622 14648 21646
rect 14614 21612 14648 21622
rect 14614 21554 14641 21574
rect 14641 21554 14648 21574
rect 14614 21540 14648 21554
rect 14614 21486 14641 21502
rect 14641 21486 14648 21502
rect 14614 21468 14648 21486
rect 14614 21418 14641 21430
rect 14641 21418 14648 21430
rect 14614 21396 14648 21418
rect 14614 21350 14641 21358
rect 14641 21350 14648 21358
rect 14614 21324 14648 21350
rect 14614 21282 14641 21286
rect 14641 21282 14648 21286
rect 14614 21252 14648 21282
rect 14614 21180 14648 21214
rect 14614 21112 14648 21142
rect 14614 21108 14641 21112
rect 14641 21108 14648 21112
rect 14614 21044 14648 21070
rect 14614 21036 14641 21044
rect 14641 21036 14648 21044
rect 14614 20976 14648 20998
rect 14614 20964 14641 20976
rect 14641 20964 14648 20976
rect 14614 20908 14648 20926
rect 14614 20892 14641 20908
rect 14641 20892 14648 20908
rect 14614 20840 14648 20854
rect 14614 20820 14641 20840
rect 14641 20820 14648 20840
rect 14614 20772 14648 20782
rect 14614 20748 14641 20772
rect 14641 20748 14648 20772
rect 14614 20704 14648 20710
rect 14614 20676 14641 20704
rect 14641 20676 14648 20704
rect 14614 20636 14648 20638
rect 14614 20604 14641 20636
rect 14641 20604 14648 20636
rect 14614 20534 14641 20566
rect 14641 20534 14648 20566
rect 14614 20532 14648 20534
rect 14614 20466 14641 20494
rect 14641 20466 14648 20494
rect 14614 20460 14648 20466
rect 14614 20398 14641 20422
rect 14641 20398 14648 20422
rect 14614 20388 14648 20398
rect 14614 20330 14641 20350
rect 14641 20330 14648 20350
rect 14614 20316 14648 20330
rect 14614 20262 14641 20278
rect 14641 20262 14648 20278
rect 14614 20244 14648 20262
rect 14614 20194 14641 20206
rect 14641 20194 14648 20206
rect 14614 20172 14648 20194
rect 14614 20126 14641 20134
rect 14641 20126 14648 20134
rect 14614 20100 14648 20126
rect 14614 20058 14641 20062
rect 14641 20058 14648 20062
rect 14614 20028 14648 20058
rect 14614 19956 14648 19990
rect 14614 19888 14648 19918
rect 14614 19884 14641 19888
rect 14641 19884 14648 19888
rect 14614 19820 14648 19846
rect 14614 19812 14641 19820
rect 14641 19812 14648 19820
rect 14614 19752 14648 19774
rect 14614 19740 14641 19752
rect 14641 19740 14648 19752
rect 14614 19684 14648 19702
rect 14614 19668 14641 19684
rect 14641 19668 14648 19684
rect 14614 19616 14648 19630
rect 14614 19596 14641 19616
rect 14641 19596 14648 19616
rect 14614 19548 14648 19558
rect 14614 19524 14641 19548
rect 14641 19524 14648 19548
rect 14614 19480 14648 19486
rect 14614 19452 14641 19480
rect 14641 19452 14648 19480
rect 14614 19412 14648 19414
rect 14614 19380 14641 19412
rect 14641 19380 14648 19412
rect 14614 19310 14641 19342
rect 14641 19310 14648 19342
rect 14614 19308 14648 19310
rect 14614 19242 14641 19270
rect 14641 19242 14648 19270
rect 14614 19236 14648 19242
rect 14614 19174 14641 19198
rect 14641 19174 14648 19198
rect 14614 19164 14648 19174
rect 14614 19106 14641 19126
rect 14641 19106 14648 19126
rect 14614 19092 14648 19106
rect 14614 19038 14641 19054
rect 14641 19038 14648 19054
rect 14614 19020 14648 19038
rect 14614 18970 14641 18982
rect 14641 18970 14648 18982
rect 14614 18948 14648 18970
rect 14614 18902 14641 18910
rect 14641 18902 14648 18910
rect 14614 18876 14648 18902
rect 14614 18834 14641 18838
rect 14641 18834 14648 18838
rect 14614 18804 14648 18834
rect 14614 18732 14648 18766
rect 14614 18664 14648 18694
rect 14614 18660 14641 18664
rect 14641 18660 14648 18664
rect 14614 18596 14648 18622
rect 14614 18588 14641 18596
rect 14641 18588 14648 18596
rect 14614 18528 14648 18550
rect 14614 18516 14641 18528
rect 14641 18516 14648 18528
rect 14614 18460 14648 18478
rect 14614 18444 14641 18460
rect 14641 18444 14648 18460
rect 14614 18392 14648 18406
rect 14614 18372 14641 18392
rect 14641 18372 14648 18392
rect 14614 18324 14648 18334
rect 14614 18300 14641 18324
rect 14641 18300 14648 18324
rect 14614 18256 14648 18262
rect 14614 18228 14641 18256
rect 14641 18228 14648 18256
rect 14614 18188 14648 18190
rect 14614 18156 14641 18188
rect 14641 18156 14648 18188
rect 14614 18086 14641 18118
rect 14641 18086 14648 18118
rect 14614 18084 14648 18086
rect 14614 18018 14641 18046
rect 14641 18018 14648 18046
rect 14614 18012 14648 18018
rect 14614 17950 14641 17974
rect 14641 17950 14648 17974
rect 14614 17940 14648 17950
rect 14614 17882 14641 17902
rect 14641 17882 14648 17902
rect 14614 17868 14648 17882
rect 14614 17814 14641 17830
rect 14641 17814 14648 17830
rect 14614 17796 14648 17814
rect 14614 17746 14641 17758
rect 14641 17746 14648 17758
rect 14614 17724 14648 17746
rect 14614 17678 14641 17686
rect 14641 17678 14648 17686
rect 14614 17652 14648 17678
rect 14614 17610 14641 17614
rect 14641 17610 14648 17614
rect 14614 17580 14648 17610
rect 14614 17508 14648 17542
rect 14614 17440 14648 17470
rect 14614 17436 14641 17440
rect 14641 17436 14648 17440
rect 14614 17372 14648 17398
rect 14614 17364 14641 17372
rect 14641 17364 14648 17372
rect 14614 17304 14648 17326
rect 14614 17292 14641 17304
rect 14641 17292 14648 17304
rect 14614 17236 14648 17254
rect 14614 17220 14641 17236
rect 14641 17220 14648 17236
rect 14614 17168 14648 17182
rect 14614 17148 14641 17168
rect 14641 17148 14648 17168
rect 14614 17100 14648 17110
rect 14614 17076 14641 17100
rect 14641 17076 14648 17100
rect 14614 17032 14648 17038
rect 14614 17004 14641 17032
rect 14641 17004 14648 17032
rect 14614 16964 14648 16966
rect 14614 16932 14641 16964
rect 14641 16932 14648 16964
rect 14614 16862 14641 16894
rect 14641 16862 14648 16894
rect 14614 16860 14648 16862
rect 14614 16794 14641 16822
rect 14641 16794 14648 16822
rect 14614 16788 14648 16794
rect 14614 16726 14641 16750
rect 14641 16726 14648 16750
rect 14614 16716 14648 16726
rect 14614 16658 14641 16678
rect 14641 16658 14648 16678
rect 14614 16644 14648 16658
rect 14614 16590 14641 16606
rect 14641 16590 14648 16606
rect 14614 16572 14648 16590
rect 14614 16522 14641 16534
rect 14641 16522 14648 16534
rect 14614 16500 14648 16522
rect 14614 16454 14641 16462
rect 14641 16454 14648 16462
rect 14614 16428 14648 16454
rect 14614 16386 14641 16390
rect 14641 16386 14648 16390
rect 14614 16356 14648 16386
rect 14614 16284 14648 16318
rect 14614 16216 14648 16246
rect 14614 16212 14641 16216
rect 14641 16212 14648 16216
rect 14614 16148 14648 16174
rect 14614 16140 14641 16148
rect 14641 16140 14648 16148
rect 14614 16080 14648 16102
rect 14614 16068 14641 16080
rect 14641 16068 14648 16080
rect 14614 16012 14648 16030
rect 14614 15996 14641 16012
rect 14641 15996 14648 16012
rect 14614 15944 14648 15958
rect 14614 15924 14641 15944
rect 14641 15924 14648 15944
rect 14614 15876 14648 15886
rect 14614 15852 14641 15876
rect 14641 15852 14648 15876
rect 14614 15808 14648 15814
rect 14614 15780 14641 15808
rect 14641 15780 14648 15808
rect 14614 15740 14648 15742
rect 14614 15708 14641 15740
rect 14641 15708 14648 15740
rect 14614 15638 14641 15670
rect 14641 15638 14648 15670
rect 14614 15636 14648 15638
rect 14614 15570 14641 15598
rect 14641 15570 14648 15598
rect 14614 15564 14648 15570
rect 14614 15502 14641 15526
rect 14641 15502 14648 15526
rect 14614 15492 14648 15502
rect 14614 15434 14641 15454
rect 14641 15434 14648 15454
rect 14614 15420 14648 15434
rect 14614 15366 14641 15382
rect 14641 15366 14648 15382
rect 14614 15348 14648 15366
rect 14614 15298 14641 15310
rect 14641 15298 14648 15310
rect 14614 15276 14648 15298
rect 14614 15230 14641 15238
rect 14641 15230 14648 15238
rect 14614 15204 14648 15230
rect 14614 15162 14641 15166
rect 14641 15162 14648 15166
rect 14614 15132 14648 15162
rect 14614 15060 14648 15094
rect 14614 14992 14648 15022
rect 14614 14988 14641 14992
rect 14641 14988 14648 14992
rect 14614 14924 14648 14950
rect 14614 14916 14641 14924
rect 14641 14916 14648 14924
rect 14614 14856 14648 14878
rect 14614 14844 14641 14856
rect 14641 14844 14648 14856
rect 14614 14788 14648 14806
rect 14614 14772 14641 14788
rect 14641 14772 14648 14788
rect 14614 14720 14648 14734
rect 14614 14700 14641 14720
rect 14641 14700 14648 14720
rect 14614 14652 14648 14662
rect 14614 14628 14641 14652
rect 14641 14628 14648 14652
rect 14614 14584 14648 14590
rect 14614 14556 14641 14584
rect 14641 14556 14648 14584
rect 14614 14516 14648 14518
rect 14614 14484 14641 14516
rect 14641 14484 14648 14516
rect 14614 14414 14641 14446
rect 14641 14414 14648 14446
rect 14614 14412 14648 14414
rect 14614 14346 14641 14374
rect 14641 14346 14648 14374
rect 14614 14340 14648 14346
rect 14614 14278 14641 14302
rect 14641 14278 14648 14302
rect 14614 14268 14648 14278
rect 14614 14210 14641 14230
rect 14641 14210 14648 14230
rect 14614 14196 14648 14210
rect 14614 14142 14641 14158
rect 14641 14142 14648 14158
rect 14614 14124 14648 14142
rect 14614 14074 14641 14086
rect 14641 14074 14648 14086
rect 14614 14052 14648 14074
rect 14614 14006 14641 14014
rect 14641 14006 14648 14014
rect 14614 13980 14648 14006
rect 14614 13938 14641 13942
rect 14641 13938 14648 13942
rect 14614 13908 14648 13938
rect 14614 13836 14648 13870
rect 14614 13768 14648 13798
rect 14614 13764 14641 13768
rect 14641 13764 14648 13768
rect 14614 13700 14648 13726
rect 14614 13692 14641 13700
rect 14641 13692 14648 13700
rect 14614 13632 14648 13654
rect 14614 13620 14641 13632
rect 14641 13620 14648 13632
rect 14614 13564 14648 13582
rect 14614 13548 14641 13564
rect 14641 13548 14648 13564
rect 14614 13496 14648 13510
rect 14614 13476 14641 13496
rect 14641 13476 14648 13496
rect 14614 13428 14648 13438
rect 14614 13404 14641 13428
rect 14641 13404 14648 13428
rect 14614 13360 14648 13366
rect 14614 13332 14641 13360
rect 14641 13332 14648 13360
rect 14614 13292 14648 13294
rect 14614 13260 14641 13292
rect 14641 13260 14648 13292
rect 14614 13190 14641 13222
rect 14641 13190 14648 13222
rect 14614 13188 14648 13190
rect 14614 13122 14641 13150
rect 14641 13122 14648 13150
rect 14614 13116 14648 13122
rect 14614 13054 14641 13078
rect 14641 13054 14648 13078
rect 14614 13044 14648 13054
rect 14614 12986 14641 13006
rect 14641 12986 14648 13006
rect 14614 12972 14648 12986
rect 14614 12918 14641 12934
rect 14641 12918 14648 12934
rect 14614 12900 14648 12918
rect 14614 12850 14641 12862
rect 14641 12850 14648 12862
rect 14614 12828 14648 12850
rect 14614 12782 14641 12790
rect 14641 12782 14648 12790
rect 14614 12756 14648 12782
rect 14614 12714 14641 12718
rect 14641 12714 14648 12718
rect 14614 12684 14648 12714
rect 14614 12612 14648 12646
rect 14614 12544 14648 12574
rect 14614 12540 14641 12544
rect 14641 12540 14648 12544
rect 14614 12476 14648 12502
rect 14614 12468 14641 12476
rect 14641 12468 14648 12476
rect 14614 12408 14648 12430
rect 14614 12396 14641 12408
rect 14641 12396 14648 12408
rect 14614 12340 14648 12358
rect 14614 12324 14641 12340
rect 14641 12324 14648 12340
rect 14614 12272 14648 12286
rect 14614 12252 14641 12272
rect 14641 12252 14648 12272
rect 14614 12204 14648 12214
rect 14614 12180 14641 12204
rect 14641 12180 14648 12204
rect 14614 12136 14648 12142
rect 14614 12108 14641 12136
rect 14641 12108 14648 12136
rect 14614 12068 14648 12070
rect 14614 12036 14641 12068
rect 14641 12036 14648 12068
rect 14614 11966 14641 11998
rect 14641 11966 14648 11998
rect 14614 11964 14648 11966
rect 14614 11898 14641 11926
rect 14641 11898 14648 11926
rect 14614 11892 14648 11898
rect 14614 11830 14641 11854
rect 14641 11830 14648 11854
rect 14614 11820 14648 11830
rect 14614 11762 14641 11782
rect 14641 11762 14648 11782
rect 14614 11748 14648 11762
rect 14614 11694 14641 11710
rect 14641 11694 14648 11710
rect 14614 11676 14648 11694
rect 14614 11626 14641 11638
rect 14641 11626 14648 11638
rect 14614 11604 14648 11626
rect 14614 11558 14641 11566
rect 14641 11558 14648 11566
rect 14614 11532 14648 11558
rect 14614 11490 14641 11494
rect 14641 11490 14648 11494
rect 14614 11460 14648 11490
rect 14614 11388 14648 11422
rect 14614 11320 14648 11350
rect 14614 11316 14641 11320
rect 14641 11316 14648 11320
rect 14614 11252 14648 11278
rect 14614 11244 14641 11252
rect 14641 11244 14648 11252
rect 14614 11184 14648 11206
rect 14614 11172 14641 11184
rect 14641 11172 14648 11184
rect 14614 11116 14648 11134
rect 14614 11100 14641 11116
rect 14641 11100 14648 11116
rect 14614 11048 14648 11062
rect 14614 11028 14641 11048
rect 14641 11028 14648 11048
rect 14614 10980 14648 10990
rect 14614 10956 14641 10980
rect 14641 10956 14648 10980
rect 14614 10912 14648 10918
rect 14614 10884 14641 10912
rect 14641 10884 14648 10912
rect 14614 10844 14648 10846
rect 14614 10812 14641 10844
rect 14641 10812 14648 10844
rect 14614 10742 14641 10774
rect 14641 10742 14648 10774
rect 14614 10740 14648 10742
rect 14614 10674 14641 10702
rect 14641 10674 14648 10702
rect 14614 10668 14648 10674
rect 14614 10606 14641 10630
rect 14641 10606 14648 10630
rect 14614 10596 14648 10606
rect 14614 10538 14641 10558
rect 14641 10538 14648 10558
rect 14614 10524 14648 10538
rect 14614 10470 14641 10486
rect 14641 10470 14648 10486
rect 14614 10452 14648 10470
rect 14614 10402 14641 10414
rect 14641 10402 14648 10414
rect 14614 10380 14648 10402
rect 14614 10334 14641 10342
rect 14641 10334 14648 10342
rect 14614 10308 14648 10334
rect 14614 10266 14641 10270
rect 14641 10266 14648 10270
rect 14614 10236 14648 10266
rect 14614 10164 14648 10198
rect 14614 10096 14648 10126
rect 14614 10092 14641 10096
rect 14641 10092 14648 10096
rect 14614 10028 14648 10054
rect 14614 10020 14641 10028
rect 14641 10020 14648 10028
rect 14614 9960 14648 9982
rect 14614 9948 14641 9960
rect 14641 9948 14648 9960
rect 14614 9892 14648 9910
rect 14614 9876 14641 9892
rect 14641 9876 14648 9892
rect 14614 9824 14648 9838
rect 14614 9804 14641 9824
rect 14641 9804 14648 9824
rect 14614 9756 14648 9766
rect 14614 9732 14641 9756
rect 14641 9732 14648 9756
rect 320 9682 354 9697
rect 320 9663 346 9682
rect 346 9663 354 9682
rect 14614 9688 14648 9694
rect 14614 9660 14641 9688
rect 14641 9660 14648 9688
rect 320 9418 354 9452
rect 610 9451 644 9452
rect 2311 9451 2345 9452
rect 2383 9451 2417 9452
rect 2455 9451 2489 9452
rect 2527 9451 2561 9452
rect 2599 9451 2633 9452
rect 2671 9451 2705 9452
rect 2743 9451 2777 9452
rect 2815 9451 2849 9452
rect 2887 9451 2921 9452
rect 2959 9451 2993 9452
rect 3031 9451 3065 9452
rect 3103 9451 3137 9452
rect 3175 9451 3209 9452
rect 3247 9451 3281 9452
rect 3319 9451 3353 9452
rect 3391 9451 3425 9452
rect 3463 9451 3497 9452
rect 3535 9451 3569 9452
rect 3607 9451 3641 9452
rect 3679 9451 3713 9452
rect 3751 9451 3785 9452
rect 3823 9451 3857 9452
rect 3895 9451 3929 9452
rect 3967 9451 4001 9452
rect 4039 9451 4073 9452
rect 4111 9451 4145 9452
rect 4183 9451 4217 9452
rect 4255 9451 4289 9452
rect 4327 9451 4361 9452
rect 4399 9451 4433 9452
rect 4471 9451 4505 9452
rect 4543 9451 4577 9452
rect 4615 9451 4649 9452
rect 4687 9451 4721 9452
rect 4759 9451 4793 9452
rect 4831 9451 4865 9452
rect 4903 9451 4937 9452
rect 4975 9451 5009 9452
rect 5047 9451 5081 9452
rect 5119 9451 5153 9452
rect 5191 9451 5225 9452
rect 5263 9451 5297 9452
rect 5335 9451 5369 9452
rect 5407 9451 5441 9452
rect 5479 9451 5513 9452
rect 5551 9451 5585 9452
rect 5623 9451 5657 9452
rect 5695 9451 5729 9452
rect 5767 9451 5801 9452
rect 5839 9451 5873 9452
rect 5911 9451 5945 9452
rect 5983 9451 6017 9452
rect 6055 9451 6089 9452
rect 6127 9451 6161 9452
rect 6199 9451 6233 9452
rect 6271 9451 6305 9452
rect 6343 9451 6377 9452
rect 6415 9451 6449 9452
rect 6487 9451 6521 9452
rect 6559 9451 6593 9452
rect 6631 9451 6665 9452
rect 6703 9451 6737 9452
rect 6775 9451 6809 9452
rect 6847 9451 6881 9452
rect 6919 9451 6953 9452
rect 6991 9451 7025 9452
rect 7063 9451 7097 9452
rect 7135 9451 7169 9452
rect 7207 9451 7241 9452
rect 7279 9451 7313 9452
rect 7351 9451 7385 9452
rect 7423 9451 7457 9452
rect 7495 9451 7529 9452
rect 7567 9451 7601 9452
rect 7639 9451 7673 9452
rect 7711 9451 7745 9452
rect 7783 9451 7817 9452
rect 7855 9451 7889 9452
rect 7927 9451 7961 9452
rect 7999 9451 8033 9452
rect 8071 9451 8105 9452
rect 8143 9451 8177 9452
rect 8215 9451 8249 9452
rect 8287 9451 8321 9452
rect 8359 9451 8393 9452
rect 8431 9451 8465 9452
rect 8503 9451 8537 9452
rect 8575 9451 8609 9452
rect 8647 9451 8681 9452
rect 8719 9451 8753 9452
rect 8791 9451 8825 9452
rect 8863 9451 8897 9452
rect 8935 9451 8969 9452
rect 9007 9451 9041 9452
rect 9079 9451 9113 9452
rect 9151 9451 9185 9452
rect 9223 9451 9257 9452
rect 9295 9451 9329 9452
rect 9367 9451 9401 9452
rect 9439 9451 9473 9452
rect 9511 9451 9545 9452
rect 9583 9451 9617 9452
rect 9655 9451 9689 9452
rect 9727 9451 9761 9452
rect 9799 9451 9833 9452
rect 9871 9451 9905 9452
rect 9943 9451 9977 9452
rect 10015 9451 10049 9452
rect 10087 9451 10121 9452
rect 10159 9451 10193 9452
rect 10231 9451 10265 9452
rect 10303 9451 10337 9452
rect 10375 9451 10409 9452
rect 10447 9451 10481 9452
rect 10519 9451 10553 9452
rect 10591 9451 10625 9452
rect 10663 9451 10697 9452
rect 10735 9451 10769 9452
rect 10807 9451 10841 9452
rect 10879 9451 10913 9452
rect 10951 9451 10985 9452
rect 11023 9451 11057 9452
rect 11095 9451 11129 9452
rect 11167 9451 11201 9452
rect 11239 9451 11273 9452
rect 11311 9451 11345 9452
rect 11383 9451 11417 9452
rect 11455 9451 11489 9452
rect 11527 9451 11561 9452
rect 11599 9451 11633 9452
rect 11671 9451 11705 9452
rect 11743 9451 11777 9452
rect 11815 9451 11849 9452
rect 11887 9451 11921 9452
rect 11959 9451 11993 9452
rect 12031 9451 12065 9452
rect 12103 9451 12137 9452
rect 12175 9451 12209 9452
rect 12247 9451 12281 9452
rect 12319 9451 12353 9452
rect 12391 9451 12425 9452
rect 12463 9451 12497 9452
rect 12535 9451 12569 9452
rect 12607 9451 12641 9452
rect 610 9418 612 9451
rect 612 9418 644 9451
rect 2311 9418 2312 9451
rect 2312 9418 2345 9451
rect 2383 9418 2414 9451
rect 2414 9418 2417 9451
rect 2455 9418 2482 9451
rect 2482 9418 2489 9451
rect 2527 9418 2550 9451
rect 2550 9418 2561 9451
rect 2599 9418 2618 9451
rect 2618 9418 2633 9451
rect 2671 9418 2686 9451
rect 2686 9418 2705 9451
rect 2743 9418 2754 9451
rect 2754 9418 2777 9451
rect 2815 9418 2822 9451
rect 2822 9418 2849 9451
rect 2887 9418 2890 9451
rect 2890 9418 2921 9451
rect 2959 9418 2992 9451
rect 2992 9418 2993 9451
rect 3031 9418 3060 9451
rect 3060 9418 3065 9451
rect 3103 9418 3128 9451
rect 3128 9418 3137 9451
rect 3175 9418 3196 9451
rect 3196 9418 3209 9451
rect 3247 9418 3264 9451
rect 3264 9418 3281 9451
rect 3319 9418 3332 9451
rect 3332 9418 3353 9451
rect 3391 9418 3400 9451
rect 3400 9418 3425 9451
rect 3463 9418 3468 9451
rect 3468 9418 3497 9451
rect 3535 9418 3536 9451
rect 3536 9418 3569 9451
rect 3607 9418 3638 9451
rect 3638 9418 3641 9451
rect 3679 9418 3706 9451
rect 3706 9418 3713 9451
rect 3751 9418 3774 9451
rect 3774 9418 3785 9451
rect 3823 9418 3842 9451
rect 3842 9418 3857 9451
rect 3895 9418 3910 9451
rect 3910 9418 3929 9451
rect 3967 9418 3978 9451
rect 3978 9418 4001 9451
rect 4039 9418 4046 9451
rect 4046 9418 4073 9451
rect 4111 9418 4114 9451
rect 4114 9418 4145 9451
rect 4183 9418 4216 9451
rect 4216 9418 4217 9451
rect 4255 9418 4284 9451
rect 4284 9418 4289 9451
rect 4327 9418 4352 9451
rect 4352 9418 4361 9451
rect 4399 9418 4420 9451
rect 4420 9418 4433 9451
rect 4471 9418 4488 9451
rect 4488 9418 4505 9451
rect 4543 9418 4556 9451
rect 4556 9418 4577 9451
rect 4615 9418 4624 9451
rect 4624 9418 4649 9451
rect 4687 9418 4692 9451
rect 4692 9418 4721 9451
rect 4759 9418 4760 9451
rect 4760 9418 4793 9451
rect 4831 9418 4862 9451
rect 4862 9418 4865 9451
rect 4903 9418 4930 9451
rect 4930 9418 4937 9451
rect 4975 9418 4998 9451
rect 4998 9418 5009 9451
rect 5047 9418 5066 9451
rect 5066 9418 5081 9451
rect 5119 9418 5134 9451
rect 5134 9418 5153 9451
rect 5191 9418 5202 9451
rect 5202 9418 5225 9451
rect 5263 9418 5270 9451
rect 5270 9418 5297 9451
rect 5335 9418 5338 9451
rect 5338 9418 5369 9451
rect 5407 9418 5440 9451
rect 5440 9418 5441 9451
rect 5479 9418 5508 9451
rect 5508 9418 5513 9451
rect 5551 9418 5576 9451
rect 5576 9418 5585 9451
rect 5623 9418 5644 9451
rect 5644 9418 5657 9451
rect 5695 9418 5712 9451
rect 5712 9418 5729 9451
rect 5767 9418 5780 9451
rect 5780 9418 5801 9451
rect 5839 9418 5848 9451
rect 5848 9418 5873 9451
rect 5911 9418 5916 9451
rect 5916 9418 5945 9451
rect 5983 9418 5984 9451
rect 5984 9418 6017 9451
rect 6055 9418 6086 9451
rect 6086 9418 6089 9451
rect 6127 9418 6154 9451
rect 6154 9418 6161 9451
rect 6199 9418 6222 9451
rect 6222 9418 6233 9451
rect 6271 9418 6290 9451
rect 6290 9418 6305 9451
rect 6343 9418 6358 9451
rect 6358 9418 6377 9451
rect 6415 9418 6426 9451
rect 6426 9418 6449 9451
rect 6487 9418 6494 9451
rect 6494 9418 6521 9451
rect 6559 9418 6562 9451
rect 6562 9418 6593 9451
rect 6631 9418 6664 9451
rect 6664 9418 6665 9451
rect 6703 9418 6732 9451
rect 6732 9418 6737 9451
rect 6775 9418 6800 9451
rect 6800 9418 6809 9451
rect 6847 9418 6868 9451
rect 6868 9418 6881 9451
rect 6919 9418 6936 9451
rect 6936 9418 6953 9451
rect 6991 9418 7004 9451
rect 7004 9418 7025 9451
rect 7063 9418 7072 9451
rect 7072 9418 7097 9451
rect 7135 9418 7140 9451
rect 7140 9418 7169 9451
rect 7207 9418 7208 9451
rect 7208 9418 7241 9451
rect 7279 9418 7310 9451
rect 7310 9418 7313 9451
rect 7351 9418 7378 9451
rect 7378 9418 7385 9451
rect 7423 9418 7446 9451
rect 7446 9418 7457 9451
rect 7495 9418 7514 9451
rect 7514 9418 7529 9451
rect 7567 9418 7582 9451
rect 7582 9418 7601 9451
rect 7639 9418 7650 9451
rect 7650 9418 7673 9451
rect 7711 9418 7718 9451
rect 7718 9418 7745 9451
rect 7783 9418 7786 9451
rect 7786 9418 7817 9451
rect 7855 9418 7888 9451
rect 7888 9418 7889 9451
rect 7927 9418 7956 9451
rect 7956 9418 7961 9451
rect 7999 9418 8024 9451
rect 8024 9418 8033 9451
rect 8071 9418 8092 9451
rect 8092 9418 8105 9451
rect 8143 9418 8160 9451
rect 8160 9418 8177 9451
rect 8215 9418 8228 9451
rect 8228 9418 8249 9451
rect 8287 9418 8296 9451
rect 8296 9418 8321 9451
rect 8359 9418 8364 9451
rect 8364 9418 8393 9451
rect 8431 9418 8432 9451
rect 8432 9418 8465 9451
rect 8503 9418 8534 9451
rect 8534 9418 8537 9451
rect 8575 9418 8602 9451
rect 8602 9418 8609 9451
rect 8647 9418 8670 9451
rect 8670 9418 8681 9451
rect 8719 9418 8738 9451
rect 8738 9418 8753 9451
rect 8791 9418 8806 9451
rect 8806 9418 8825 9451
rect 8863 9418 8874 9451
rect 8874 9418 8897 9451
rect 8935 9418 8942 9451
rect 8942 9418 8969 9451
rect 9007 9418 9010 9451
rect 9010 9418 9041 9451
rect 9079 9418 9112 9451
rect 9112 9418 9113 9451
rect 9151 9418 9180 9451
rect 9180 9418 9185 9451
rect 9223 9418 9248 9451
rect 9248 9418 9257 9451
rect 9295 9418 9316 9451
rect 9316 9418 9329 9451
rect 9367 9418 9384 9451
rect 9384 9418 9401 9451
rect 9439 9418 9452 9451
rect 9452 9418 9473 9451
rect 9511 9418 9520 9451
rect 9520 9418 9545 9451
rect 9583 9418 9588 9451
rect 9588 9418 9617 9451
rect 9655 9418 9656 9451
rect 9656 9418 9689 9451
rect 9727 9418 9758 9451
rect 9758 9418 9761 9451
rect 9799 9418 9826 9451
rect 9826 9418 9833 9451
rect 9871 9418 9894 9451
rect 9894 9418 9905 9451
rect 9943 9418 9962 9451
rect 9962 9418 9977 9451
rect 10015 9418 10030 9451
rect 10030 9418 10049 9451
rect 10087 9418 10098 9451
rect 10098 9418 10121 9451
rect 10159 9418 10166 9451
rect 10166 9418 10193 9451
rect 10231 9418 10234 9451
rect 10234 9418 10265 9451
rect 10303 9418 10336 9451
rect 10336 9418 10337 9451
rect 10375 9418 10404 9451
rect 10404 9418 10409 9451
rect 10447 9418 10472 9451
rect 10472 9418 10481 9451
rect 10519 9418 10540 9451
rect 10540 9418 10553 9451
rect 10591 9418 10608 9451
rect 10608 9418 10625 9451
rect 10663 9418 10676 9451
rect 10676 9418 10697 9451
rect 10735 9418 10744 9451
rect 10744 9418 10769 9451
rect 10807 9418 10812 9451
rect 10812 9418 10841 9451
rect 10879 9418 10880 9451
rect 10880 9418 10913 9451
rect 10951 9418 10982 9451
rect 10982 9418 10985 9451
rect 11023 9418 11050 9451
rect 11050 9418 11057 9451
rect 11095 9418 11118 9451
rect 11118 9418 11129 9451
rect 11167 9418 11186 9451
rect 11186 9418 11201 9451
rect 11239 9418 11254 9451
rect 11254 9418 11273 9451
rect 11311 9418 11322 9451
rect 11322 9418 11345 9451
rect 11383 9418 11390 9451
rect 11390 9418 11417 9451
rect 11455 9418 11458 9451
rect 11458 9418 11489 9451
rect 11527 9418 11560 9451
rect 11560 9418 11561 9451
rect 11599 9418 11628 9451
rect 11628 9418 11633 9451
rect 11671 9418 11696 9451
rect 11696 9418 11705 9451
rect 11743 9418 11764 9451
rect 11764 9418 11777 9451
rect 11815 9418 11832 9451
rect 11832 9418 11849 9451
rect 11887 9418 11900 9451
rect 11900 9418 11921 9451
rect 11959 9418 11968 9451
rect 11968 9418 11993 9451
rect 12031 9418 12036 9451
rect 12036 9418 12065 9451
rect 12103 9418 12104 9451
rect 12104 9418 12137 9451
rect 12175 9418 12206 9451
rect 12206 9418 12209 9451
rect 12247 9418 12274 9451
rect 12274 9418 12281 9451
rect 12319 9418 12342 9451
rect 12342 9418 12353 9451
rect 12391 9418 12410 9451
rect 12410 9418 12425 9451
rect 12463 9418 12478 9451
rect 12478 9418 12497 9451
rect 12535 9418 12546 9451
rect 12546 9418 12569 9451
rect 12607 9418 12614 9451
rect 12614 9418 12641 9451
rect 14314 9418 14348 9452
rect 14614 9418 14648 9452
<< metal1 >>
rect 245 36534 14724 36574
rect 245 36500 320 36534
rect 354 36533 14724 36534
rect 354 36500 14614 36533
rect 245 36499 14614 36500
rect 14648 36499 14724 36533
rect 245 36498 14724 36499
rect 245 36464 556 36498
rect 590 36464 628 36498
rect 662 36464 700 36498
rect 734 36464 772 36498
rect 806 36464 844 36498
rect 878 36464 916 36498
rect 950 36464 988 36498
rect 1022 36464 1060 36498
rect 1094 36464 1132 36498
rect 1166 36464 1204 36498
rect 1238 36464 1276 36498
rect 1310 36464 1348 36498
rect 1382 36464 1420 36498
rect 1454 36464 1492 36498
rect 1526 36464 1564 36498
rect 1598 36464 1636 36498
rect 1670 36464 1708 36498
rect 1742 36464 1780 36498
rect 1814 36464 1852 36498
rect 1886 36464 1924 36498
rect 1958 36464 1996 36498
rect 2030 36464 2068 36498
rect 2102 36464 2140 36498
rect 2174 36464 2212 36498
rect 2246 36464 2284 36498
rect 2318 36464 2356 36498
rect 2390 36464 2428 36498
rect 2462 36464 2500 36498
rect 2534 36464 2572 36498
rect 2606 36464 2644 36498
rect 2678 36464 2716 36498
rect 2750 36464 2788 36498
rect 2822 36464 2860 36498
rect 2894 36464 2932 36498
rect 2966 36464 3004 36498
rect 3038 36464 3076 36498
rect 3110 36464 3148 36498
rect 3182 36464 3220 36498
rect 3254 36464 3292 36498
rect 3326 36464 3364 36498
rect 3398 36464 3436 36498
rect 3470 36464 3508 36498
rect 3542 36464 3580 36498
rect 3614 36464 3652 36498
rect 3686 36464 3724 36498
rect 3758 36464 3796 36498
rect 3830 36464 3868 36498
rect 3902 36464 3940 36498
rect 3974 36464 4012 36498
rect 4046 36464 4084 36498
rect 4118 36464 4156 36498
rect 4190 36464 4228 36498
rect 4262 36464 4300 36498
rect 4334 36464 4372 36498
rect 4406 36464 4444 36498
rect 4478 36464 4516 36498
rect 4550 36464 4588 36498
rect 4622 36464 4660 36498
rect 4694 36464 4732 36498
rect 4766 36464 4804 36498
rect 4838 36464 4876 36498
rect 4910 36464 4948 36498
rect 4982 36464 5020 36498
rect 5054 36464 5092 36498
rect 5126 36464 5164 36498
rect 5198 36464 5236 36498
rect 5270 36464 5308 36498
rect 5342 36464 5380 36498
rect 5414 36464 5452 36498
rect 5486 36464 5524 36498
rect 5558 36464 5596 36498
rect 5630 36464 5668 36498
rect 5702 36464 5740 36498
rect 5774 36464 5812 36498
rect 5846 36464 5884 36498
rect 5918 36464 5956 36498
rect 5990 36464 6028 36498
rect 6062 36464 6100 36498
rect 6134 36464 6172 36498
rect 6206 36464 6244 36498
rect 6278 36464 6316 36498
rect 6350 36464 6388 36498
rect 6422 36464 6460 36498
rect 6494 36464 6532 36498
rect 6566 36464 6604 36498
rect 6638 36464 6676 36498
rect 6710 36464 6748 36498
rect 6782 36464 6820 36498
rect 6854 36464 6892 36498
rect 6926 36464 6964 36498
rect 6998 36464 7036 36498
rect 7070 36464 7108 36498
rect 7142 36464 7180 36498
rect 7214 36464 7252 36498
rect 7286 36464 7324 36498
rect 7358 36464 7396 36498
rect 7430 36464 7468 36498
rect 7502 36464 7540 36498
rect 7574 36464 7612 36498
rect 7646 36464 7684 36498
rect 7718 36464 7756 36498
rect 7790 36464 7828 36498
rect 7862 36464 7900 36498
rect 7934 36464 7972 36498
rect 8006 36464 8044 36498
rect 8078 36464 8116 36498
rect 8150 36464 8188 36498
rect 8222 36464 8260 36498
rect 8294 36464 8332 36498
rect 8366 36464 8404 36498
rect 8438 36464 8476 36498
rect 8510 36464 8548 36498
rect 8582 36464 8620 36498
rect 8654 36464 8692 36498
rect 8726 36464 8764 36498
rect 8798 36464 8836 36498
rect 8870 36464 8908 36498
rect 8942 36464 8980 36498
rect 9014 36464 9052 36498
rect 9086 36464 9124 36498
rect 9158 36464 9196 36498
rect 9230 36464 9268 36498
rect 9302 36464 9340 36498
rect 9374 36464 9412 36498
rect 9446 36464 9484 36498
rect 9518 36464 9556 36498
rect 9590 36464 9628 36498
rect 9662 36464 9700 36498
rect 9734 36464 9772 36498
rect 9806 36464 9844 36498
rect 9878 36464 9916 36498
rect 9950 36464 9988 36498
rect 10022 36464 10060 36498
rect 10094 36464 10132 36498
rect 10166 36464 10204 36498
rect 10238 36464 10276 36498
rect 10310 36464 10348 36498
rect 10382 36464 10420 36498
rect 10454 36464 10492 36498
rect 10526 36464 10564 36498
rect 10598 36464 10636 36498
rect 10670 36464 10708 36498
rect 10742 36464 10780 36498
rect 10814 36464 10852 36498
rect 10886 36464 10924 36498
rect 10958 36464 10996 36498
rect 11030 36464 11068 36498
rect 11102 36464 11140 36498
rect 11174 36464 11212 36498
rect 11246 36464 11284 36498
rect 11318 36464 11356 36498
rect 11390 36464 11428 36498
rect 11462 36464 11500 36498
rect 11534 36464 11572 36498
rect 11606 36464 11644 36498
rect 11678 36464 11716 36498
rect 11750 36464 11788 36498
rect 11822 36464 11860 36498
rect 11894 36464 11932 36498
rect 11966 36464 12004 36498
rect 12038 36464 12076 36498
rect 12110 36464 12148 36498
rect 12182 36464 12220 36498
rect 12254 36464 12292 36498
rect 12326 36464 12364 36498
rect 12398 36464 12436 36498
rect 12470 36464 12508 36498
rect 12542 36464 12580 36498
rect 12614 36464 12652 36498
rect 12686 36464 12724 36498
rect 12758 36464 12796 36498
rect 12830 36464 12868 36498
rect 12902 36464 12940 36498
rect 12974 36464 13012 36498
rect 13046 36464 13084 36498
rect 13118 36464 13156 36498
rect 13190 36464 13228 36498
rect 13262 36464 13300 36498
rect 13334 36464 13372 36498
rect 13406 36464 13444 36498
rect 13478 36464 13516 36498
rect 13550 36464 13588 36498
rect 13622 36464 13660 36498
rect 13694 36464 13732 36498
rect 13766 36464 13804 36498
rect 13838 36464 13876 36498
rect 13910 36464 13948 36498
rect 13982 36464 14020 36498
rect 14054 36464 14092 36498
rect 14126 36464 14164 36498
rect 14198 36464 14236 36498
rect 14270 36464 14308 36498
rect 14342 36464 14380 36498
rect 14414 36464 14724 36498
rect 245 36462 14724 36464
rect 245 36428 320 36462
rect 354 36461 14724 36462
rect 354 36428 14614 36461
rect 245 36427 14614 36428
rect 14648 36427 14724 36461
rect 245 36389 14724 36427
rect 245 36265 430 36389
rect 245 36231 320 36265
rect 354 36231 430 36265
rect 245 36193 430 36231
rect 245 36159 320 36193
rect 354 36159 430 36193
rect 245 36121 430 36159
rect 245 36087 320 36121
rect 354 36087 430 36121
rect 245 36049 430 36087
rect 14539 36262 14724 36389
rect 14539 36228 14614 36262
rect 14648 36228 14724 36262
rect 14539 36190 14724 36228
rect 14539 36156 14614 36190
rect 14648 36156 14724 36190
rect 14539 36118 14724 36156
rect 14539 36084 14614 36118
rect 14648 36084 14724 36118
rect 245 36015 320 36049
rect 354 36015 430 36049
tri 850 36046 857 36053 se
rect 857 36046 14119 36053
tri 14119 36046 14126 36053 sw
rect 14539 36046 14724 36084
tri 823 36019 850 36046 se
rect 850 36019 14126 36046
rect 245 35977 430 36015
tri 816 36012 823 36019 se
rect 823 36012 14126 36019
tri 14126 36012 14160 36046 sw
rect 14539 36012 14614 36046
rect 14648 36012 14724 36046
tri 807 36003 816 36012 se
rect 816 36003 14160 36012
rect 245 35943 320 35977
rect 354 35943 430 35977
tri 773 35969 807 36003 se
rect 807 35969 1009 36003
rect 1043 35969 1081 36003
rect 1115 35969 1153 36003
rect 1187 35969 1225 36003
rect 1259 35969 1297 36003
rect 1331 35969 1369 36003
rect 1403 35969 1441 36003
rect 1475 35969 1513 36003
rect 1547 35969 1585 36003
rect 1619 35969 1657 36003
rect 1691 35969 1729 36003
rect 1763 35969 1801 36003
rect 1835 35969 1873 36003
rect 1907 35969 1945 36003
rect 1979 35969 2017 36003
rect 2051 35969 2089 36003
rect 2123 35969 2161 36003
rect 2195 35969 2233 36003
rect 2267 35969 2305 36003
rect 2339 35969 2377 36003
rect 2411 35969 2449 36003
rect 2483 35969 2521 36003
rect 2555 35969 2593 36003
rect 2627 35969 2665 36003
rect 2699 35969 2737 36003
rect 2771 35969 2809 36003
rect 2843 35969 2881 36003
rect 2915 35969 2953 36003
rect 2987 35969 3025 36003
rect 3059 35969 3097 36003
rect 3131 35969 3169 36003
rect 3203 35969 3241 36003
rect 3275 35969 3313 36003
rect 3347 35969 3385 36003
rect 3419 35969 3457 36003
rect 3491 35969 3529 36003
rect 3563 35969 3601 36003
rect 3635 35969 3673 36003
rect 3707 35969 3745 36003
rect 3779 35969 3817 36003
rect 3851 35969 3889 36003
rect 3923 35969 3961 36003
rect 3995 35969 4033 36003
rect 4067 35969 4105 36003
rect 4139 35969 4177 36003
rect 4211 35969 4249 36003
rect 4283 35969 4321 36003
rect 4355 35969 4393 36003
rect 4427 35969 4465 36003
rect 4499 35969 4537 36003
rect 4571 35969 4609 36003
rect 4643 35969 4681 36003
rect 4715 35969 4753 36003
rect 4787 35969 4825 36003
rect 4859 35969 4897 36003
rect 4931 35969 4969 36003
rect 5003 35969 5041 36003
rect 5075 35969 5113 36003
rect 5147 35969 5185 36003
rect 5219 35969 5257 36003
rect 5291 35969 5329 36003
rect 5363 35969 5401 36003
rect 5435 35969 5473 36003
rect 5507 35969 5545 36003
rect 5579 35969 5617 36003
rect 5651 35969 5689 36003
rect 5723 35969 5761 36003
rect 5795 35969 5833 36003
rect 5867 35969 5905 36003
rect 5939 35969 5977 36003
rect 6011 35969 6049 36003
rect 6083 35969 6121 36003
rect 6155 35969 6193 36003
rect 6227 35969 6265 36003
rect 6299 35969 6337 36003
rect 6371 35969 6409 36003
rect 6443 35969 6481 36003
rect 6515 35969 6553 36003
rect 6587 35969 6625 36003
rect 6659 35969 6697 36003
rect 6731 35969 6769 36003
rect 6803 35969 6841 36003
rect 6875 35969 6913 36003
rect 6947 35969 6985 36003
rect 7019 35969 7057 36003
rect 7091 35969 7129 36003
rect 7163 35969 7201 36003
rect 7235 35969 7273 36003
rect 7307 35969 7345 36003
rect 7379 35969 7417 36003
rect 7451 35969 7489 36003
rect 7523 35969 7561 36003
rect 7595 35969 7633 36003
rect 7667 35969 7705 36003
rect 7739 35969 7777 36003
rect 7811 35969 7849 36003
rect 7883 35969 7921 36003
rect 7955 35969 7993 36003
rect 8027 35969 8065 36003
rect 8099 35969 8137 36003
rect 8171 35969 8209 36003
rect 8243 35969 8281 36003
rect 8315 35969 8353 36003
rect 8387 35969 8425 36003
rect 8459 35969 8497 36003
rect 8531 35969 8569 36003
rect 8603 35969 8641 36003
rect 8675 35969 8713 36003
rect 8747 35969 8785 36003
rect 8819 35969 8857 36003
rect 8891 35969 8929 36003
rect 8963 35969 9001 36003
rect 9035 35969 9073 36003
rect 9107 35969 9145 36003
rect 9179 35969 9217 36003
rect 9251 35969 9289 36003
rect 9323 35969 9361 36003
rect 9395 35969 9433 36003
rect 9467 35969 9505 36003
rect 9539 35969 9577 36003
rect 9611 35969 9649 36003
rect 9683 35969 9721 36003
rect 9755 35969 9793 36003
rect 9827 35969 9865 36003
rect 9899 35969 9937 36003
rect 9971 35969 10009 36003
rect 10043 35969 10081 36003
rect 10115 35969 10153 36003
rect 10187 35969 10225 36003
rect 10259 35969 10297 36003
rect 10331 35969 10369 36003
rect 10403 35969 10441 36003
rect 10475 35969 10513 36003
rect 10547 35969 10585 36003
rect 10619 35969 10657 36003
rect 10691 35969 10729 36003
rect 10763 35969 10801 36003
rect 10835 35969 10873 36003
rect 10907 35969 10945 36003
rect 10979 35969 11017 36003
rect 11051 35969 11089 36003
rect 11123 35969 11161 36003
rect 11195 35969 11233 36003
rect 11267 35969 11305 36003
rect 11339 35969 11377 36003
rect 11411 35969 11449 36003
rect 11483 35969 11521 36003
rect 11555 35969 11593 36003
rect 11627 35969 11665 36003
rect 11699 35969 11737 36003
rect 11771 35969 11809 36003
rect 11843 35969 11881 36003
rect 11915 35969 11953 36003
rect 11987 35969 12025 36003
rect 12059 35969 12097 36003
rect 12131 35969 12169 36003
rect 12203 35969 12241 36003
rect 12275 35969 12313 36003
rect 12347 35969 12385 36003
rect 12419 35969 12457 36003
rect 12491 35969 12529 36003
rect 12563 35969 12601 36003
rect 12635 35969 12673 36003
rect 12707 35969 12745 36003
rect 12779 35969 12817 36003
rect 12851 35969 12889 36003
rect 12923 35969 12961 36003
rect 12995 35969 13033 36003
rect 13067 35969 13105 36003
rect 13139 35969 13177 36003
rect 13211 35969 13249 36003
rect 13283 35969 13321 36003
rect 13355 35969 13393 36003
rect 13427 35969 13465 36003
rect 13499 35969 13537 36003
rect 13571 35969 13609 36003
rect 13643 35969 13681 36003
rect 13715 35969 13753 36003
rect 13787 35969 13825 36003
rect 13859 35969 13897 36003
rect 13931 35969 13969 36003
rect 14003 35974 14160 36003
tri 14160 35974 14198 36012 sw
rect 14539 35974 14724 36012
rect 14003 35969 14198 35974
rect 245 35905 430 35943
rect 245 35871 320 35905
rect 354 35871 430 35905
rect 245 35833 430 35871
rect 245 35799 320 35833
rect 354 35799 430 35833
rect 245 35761 430 35799
rect 245 35727 320 35761
rect 354 35727 430 35761
rect 245 35689 430 35727
rect 245 35655 320 35689
rect 354 35655 430 35689
rect 245 35617 430 35655
rect 245 35583 320 35617
rect 354 35583 430 35617
rect 245 35545 430 35583
rect 245 35511 320 35545
rect 354 35511 430 35545
rect 245 35473 430 35511
rect 245 35439 320 35473
rect 354 35439 430 35473
rect 245 35401 430 35439
rect 245 35367 320 35401
rect 354 35367 430 35401
rect 245 35329 430 35367
rect 245 35295 320 35329
rect 354 35295 430 35329
rect 245 35257 430 35295
rect 245 35223 320 35257
rect 354 35223 430 35257
rect 245 35185 430 35223
rect 245 35151 320 35185
rect 354 35151 430 35185
rect 245 35113 430 35151
rect 245 35079 320 35113
rect 354 35079 430 35113
rect 245 35041 430 35079
rect 245 35007 320 35041
rect 354 35007 430 35041
rect 245 34969 430 35007
rect 245 34935 320 34969
rect 354 34935 430 34969
rect 245 34897 430 34935
rect 245 34863 320 34897
rect 354 34863 430 34897
rect 245 34825 430 34863
rect 245 34791 320 34825
rect 354 34791 430 34825
rect 245 34753 430 34791
rect 245 34719 320 34753
rect 354 34719 430 34753
rect 245 34681 430 34719
rect 245 34647 320 34681
rect 354 34647 430 34681
rect 245 34609 430 34647
rect 245 34575 320 34609
rect 354 34575 430 34609
rect 245 34537 430 34575
rect 245 34503 320 34537
rect 354 34503 430 34537
rect 245 34465 430 34503
rect 245 34431 320 34465
rect 354 34431 430 34465
rect 245 34393 430 34431
rect 245 34359 320 34393
rect 354 34359 430 34393
rect 245 34321 430 34359
rect 245 34287 320 34321
rect 354 34287 430 34321
rect 245 34249 430 34287
rect 245 34215 320 34249
rect 354 34215 430 34249
rect 245 34177 430 34215
rect 245 34143 320 34177
rect 354 34143 430 34177
rect 245 34105 430 34143
rect 245 34071 320 34105
rect 354 34071 430 34105
rect 245 34033 430 34071
rect 245 33999 320 34033
rect 354 33999 430 34033
rect 245 33961 430 33999
rect 245 33927 320 33961
rect 354 33927 430 33961
rect 245 33889 430 33927
rect 245 33855 320 33889
rect 354 33855 430 33889
rect 245 33817 430 33855
rect 245 33783 320 33817
rect 354 33783 430 33817
rect 245 33745 430 33783
rect 245 33711 320 33745
rect 354 33711 430 33745
rect 245 33673 430 33711
rect 245 33639 320 33673
rect 354 33639 430 33673
rect 245 33601 430 33639
rect 245 33567 320 33601
rect 354 33567 430 33601
rect 245 33529 430 33567
rect 245 33495 320 33529
rect 354 33495 430 33529
rect 245 33457 430 33495
rect 245 33423 320 33457
rect 354 33423 430 33457
rect 245 33385 430 33423
rect 245 33351 320 33385
rect 354 33351 430 33385
rect 245 33313 430 33351
rect 245 33279 320 33313
rect 354 33279 430 33313
rect 245 33241 430 33279
rect 245 33207 320 33241
rect 354 33207 430 33241
rect 245 33169 430 33207
rect 245 33135 320 33169
rect 354 33135 430 33169
rect 245 33097 430 33135
rect 245 33063 320 33097
rect 354 33063 430 33097
rect 245 33025 430 33063
rect 245 32991 320 33025
rect 354 32991 430 33025
rect 245 32953 430 32991
rect 245 32919 320 32953
rect 354 32919 430 32953
rect 245 32881 430 32919
rect 245 32847 320 32881
rect 354 32847 430 32881
rect 245 32809 430 32847
rect 245 32775 320 32809
rect 354 32775 430 32809
rect 245 32737 430 32775
rect 245 32703 320 32737
rect 354 32703 430 32737
rect 245 32665 430 32703
rect 245 32631 320 32665
rect 354 32631 430 32665
rect 245 32593 430 32631
rect 245 32559 320 32593
rect 354 32559 430 32593
rect 245 32521 430 32559
rect 245 32487 320 32521
rect 354 32487 430 32521
rect 245 32449 430 32487
rect 245 32415 320 32449
rect 354 32415 430 32449
rect 245 32377 430 32415
rect 245 32343 320 32377
rect 354 32343 430 32377
rect 245 32305 430 32343
rect 245 32271 320 32305
rect 354 32271 430 32305
rect 245 32233 430 32271
rect 245 32199 320 32233
rect 354 32199 430 32233
rect 245 32161 430 32199
rect 245 32127 320 32161
rect 354 32127 430 32161
rect 245 32089 430 32127
rect 245 32055 320 32089
rect 354 32055 430 32089
rect 245 32017 430 32055
rect 245 31983 320 32017
rect 354 31983 430 32017
rect 245 31945 430 31983
rect 245 31911 320 31945
rect 354 31911 430 31945
rect 245 31873 430 31911
rect 245 31839 320 31873
rect 354 31839 430 31873
rect 245 31801 430 31839
rect 245 31767 320 31801
rect 354 31767 430 31801
rect 245 31729 430 31767
rect 245 31695 320 31729
rect 354 31695 430 31729
rect 245 31657 430 31695
rect 245 31623 320 31657
rect 354 31623 430 31657
rect 245 31585 430 31623
rect 245 31551 320 31585
rect 354 31551 430 31585
rect 245 31513 430 31551
rect 245 31479 320 31513
rect 354 31479 430 31513
rect 245 31441 430 31479
rect 245 31407 320 31441
rect 354 31407 430 31441
rect 245 31369 430 31407
rect 245 31335 320 31369
rect 354 31335 430 31369
rect 245 31297 430 31335
rect 245 31263 320 31297
rect 354 31263 430 31297
rect 245 31225 430 31263
rect 245 31191 320 31225
rect 354 31191 430 31225
rect 245 31153 430 31191
rect 245 31119 320 31153
rect 354 31119 430 31153
rect 245 31081 430 31119
rect 245 31047 320 31081
rect 354 31047 430 31081
rect 245 31009 430 31047
rect 245 30975 320 31009
rect 354 30975 430 31009
rect 245 30937 430 30975
rect 245 30903 320 30937
rect 354 30903 430 30937
rect 245 30865 430 30903
rect 245 30831 320 30865
rect 354 30831 430 30865
rect 245 30793 430 30831
rect 245 30759 320 30793
rect 354 30759 430 30793
rect 245 30721 430 30759
rect 245 30687 320 30721
rect 354 30687 430 30721
rect 245 30649 430 30687
rect 245 30615 320 30649
rect 354 30615 430 30649
rect 245 30577 430 30615
rect 245 30543 320 30577
rect 354 30543 430 30577
rect 245 30505 430 30543
rect 245 30471 320 30505
rect 354 30471 430 30505
rect 245 30433 430 30471
rect 245 30399 320 30433
rect 354 30399 430 30433
rect 245 30361 430 30399
rect 245 30327 320 30361
rect 354 30327 430 30361
rect 245 30289 430 30327
rect 245 30255 320 30289
rect 354 30255 430 30289
rect 245 30217 430 30255
rect 245 30183 320 30217
rect 354 30183 430 30217
rect 245 30145 430 30183
rect 245 30111 320 30145
rect 354 30111 430 30145
rect 245 30073 430 30111
rect 245 30039 320 30073
rect 354 30039 430 30073
rect 245 30001 430 30039
rect 245 29967 320 30001
rect 354 29967 430 30001
rect 245 29929 430 29967
rect 245 29895 320 29929
rect 354 29895 430 29929
rect 245 29857 430 29895
rect 245 29823 320 29857
rect 354 29823 430 29857
rect 245 29785 430 29823
rect 245 29751 320 29785
rect 354 29751 430 29785
rect 245 29713 430 29751
rect 245 29679 320 29713
rect 354 29679 430 29713
rect 245 29641 430 29679
rect 245 29607 320 29641
rect 354 29607 430 29641
rect 245 29569 430 29607
rect 245 29535 320 29569
rect 354 29535 430 29569
rect 245 29497 430 29535
rect 245 29463 320 29497
rect 354 29463 430 29497
rect 245 29425 430 29463
rect 245 29391 320 29425
rect 354 29391 430 29425
rect 245 29353 430 29391
rect 245 29319 320 29353
rect 354 29319 430 29353
rect 245 29281 430 29319
rect 245 29247 320 29281
rect 354 29247 430 29281
rect 245 29209 430 29247
rect 245 29175 320 29209
rect 354 29175 430 29209
rect 245 29137 430 29175
rect 245 29103 320 29137
rect 354 29103 430 29137
rect 245 29065 430 29103
rect 245 29031 320 29065
rect 354 29031 430 29065
rect 245 28993 430 29031
rect 245 28959 320 28993
rect 354 28959 430 28993
rect 245 28921 430 28959
rect 245 28887 320 28921
rect 354 28887 430 28921
rect 245 28849 430 28887
rect 245 28815 320 28849
rect 354 28815 430 28849
rect 245 28777 430 28815
rect 245 28743 320 28777
rect 354 28743 430 28777
rect 245 28705 430 28743
rect 245 28671 320 28705
rect 354 28671 430 28705
rect 245 28633 430 28671
rect 245 28599 320 28633
rect 354 28599 430 28633
rect 245 28561 430 28599
rect 245 28527 320 28561
rect 354 28527 430 28561
rect 245 28489 430 28527
rect 245 28455 320 28489
rect 354 28455 430 28489
rect 245 28417 430 28455
rect 245 28383 320 28417
rect 354 28383 430 28417
rect 245 28345 430 28383
rect 245 28311 320 28345
rect 354 28311 430 28345
rect 245 28273 430 28311
rect 245 28239 320 28273
rect 354 28239 430 28273
rect 245 28201 430 28239
rect 245 28167 320 28201
rect 354 28167 430 28201
rect 245 28129 430 28167
rect 245 28095 320 28129
rect 354 28095 430 28129
rect 245 28057 430 28095
rect 245 28023 320 28057
rect 354 28023 430 28057
rect 245 27985 430 28023
rect 245 27951 320 27985
rect 354 27951 430 27985
rect 245 27913 430 27951
rect 245 27879 320 27913
rect 354 27879 430 27913
rect 245 27841 430 27879
rect 245 27807 320 27841
rect 354 27807 430 27841
rect 245 27769 430 27807
rect 245 27735 320 27769
rect 354 27735 430 27769
rect 245 27697 430 27735
rect 245 27663 320 27697
rect 354 27663 430 27697
rect 245 27625 430 27663
rect 245 27591 320 27625
rect 354 27591 430 27625
rect 245 27553 430 27591
rect 245 27519 320 27553
rect 354 27519 430 27553
rect 245 27481 430 27519
rect 245 27447 320 27481
rect 354 27447 430 27481
rect 245 27409 430 27447
rect 245 27375 320 27409
rect 354 27375 430 27409
rect 245 27337 430 27375
rect 245 27303 320 27337
rect 354 27303 430 27337
rect 245 27265 430 27303
rect 245 27231 320 27265
rect 354 27231 430 27265
rect 245 27193 430 27231
rect 245 27159 320 27193
rect 354 27159 430 27193
rect 245 27121 430 27159
rect 245 27087 320 27121
rect 354 27087 430 27121
rect 245 27049 430 27087
rect 245 27015 320 27049
rect 354 27015 430 27049
rect 245 26977 430 27015
rect 245 26943 320 26977
rect 354 26943 430 26977
rect 245 26905 430 26943
rect 245 26871 320 26905
rect 354 26871 430 26905
rect 245 26833 430 26871
rect 245 26799 320 26833
rect 354 26799 430 26833
rect 245 26761 430 26799
rect 245 26727 320 26761
rect 354 26727 430 26761
rect 245 26689 430 26727
rect 245 26655 320 26689
rect 354 26655 430 26689
rect 245 26617 430 26655
rect 245 26583 320 26617
rect 354 26583 430 26617
rect 245 26545 430 26583
rect 245 26511 320 26545
rect 354 26511 430 26545
rect 245 26473 430 26511
rect 245 26439 320 26473
rect 354 26439 430 26473
rect 245 26401 430 26439
rect 245 26367 320 26401
rect 354 26367 430 26401
rect 245 26329 430 26367
rect 245 26295 320 26329
rect 354 26295 430 26329
rect 245 26257 430 26295
rect 245 26223 320 26257
rect 354 26223 430 26257
rect 245 26185 430 26223
rect 245 26151 320 26185
rect 354 26151 430 26185
rect 245 26113 430 26151
rect 245 26079 320 26113
rect 354 26079 430 26113
rect 245 26041 430 26079
rect 245 26007 320 26041
rect 354 26007 430 26041
rect 245 25969 430 26007
rect 245 25935 320 25969
rect 354 25935 430 25969
rect 245 25897 430 25935
rect 245 25863 320 25897
rect 354 25863 430 25897
rect 245 25825 430 25863
rect 245 25791 320 25825
rect 354 25791 430 25825
rect 245 25753 430 25791
rect 245 25719 320 25753
rect 354 25719 430 25753
rect 245 25681 430 25719
rect 245 25647 320 25681
rect 354 25647 430 25681
rect 245 25609 430 25647
rect 245 25575 320 25609
rect 354 25575 430 25609
rect 245 25537 430 25575
rect 245 25503 320 25537
rect 354 25503 430 25537
rect 245 25465 430 25503
rect 245 25431 320 25465
rect 354 25431 430 25465
rect 245 25393 430 25431
rect 245 25359 320 25393
rect 354 25359 430 25393
rect 245 25321 430 25359
rect 245 25287 320 25321
rect 354 25287 430 25321
rect 245 25249 430 25287
rect 245 25215 320 25249
rect 354 25215 430 25249
rect 245 25177 430 25215
rect 245 25143 320 25177
rect 354 25143 430 25177
rect 245 25105 430 25143
rect 245 25071 320 25105
rect 354 25071 430 25105
rect 245 25033 430 25071
rect 245 24999 320 25033
rect 354 24999 430 25033
rect 245 24961 430 24999
rect 245 24927 320 24961
rect 354 24927 430 24961
rect 245 24889 430 24927
rect 245 24855 320 24889
rect 354 24855 430 24889
rect 245 24817 430 24855
rect 245 24783 320 24817
rect 354 24783 430 24817
rect 245 24745 430 24783
rect 245 24711 320 24745
rect 354 24711 430 24745
rect 245 24673 430 24711
rect 245 24639 320 24673
rect 354 24639 430 24673
rect 245 24601 430 24639
rect 245 24567 320 24601
rect 354 24567 430 24601
rect 245 24529 430 24567
rect 245 24495 320 24529
rect 354 24495 430 24529
rect 245 24457 430 24495
rect 245 24423 320 24457
rect 354 24423 430 24457
rect 245 24385 430 24423
rect 245 24351 320 24385
rect 354 24351 430 24385
rect 245 24313 430 24351
rect 245 24279 320 24313
rect 354 24279 430 24313
rect 245 24241 430 24279
rect 245 24207 320 24241
rect 354 24207 430 24241
rect 245 24169 430 24207
rect 245 24135 320 24169
rect 354 24135 430 24169
rect 245 24097 430 24135
rect 245 24063 320 24097
rect 354 24063 430 24097
rect 245 24025 430 24063
rect 245 23991 320 24025
rect 354 23991 430 24025
rect 245 23953 430 23991
rect 245 23919 320 23953
rect 354 23919 430 23953
rect 245 23881 430 23919
rect 245 23847 320 23881
rect 354 23847 430 23881
rect 245 23809 430 23847
rect 245 23775 320 23809
rect 354 23775 430 23809
rect 245 23737 430 23775
rect 245 23703 320 23737
rect 354 23703 430 23737
rect 245 23665 430 23703
rect 245 23631 320 23665
rect 354 23631 430 23665
rect 245 23593 430 23631
rect 245 23559 320 23593
rect 354 23559 430 23593
rect 245 23521 430 23559
rect 245 23487 320 23521
rect 354 23487 430 23521
rect 245 23449 430 23487
rect 245 23415 320 23449
rect 354 23415 430 23449
rect 245 23377 430 23415
rect 245 23343 320 23377
rect 354 23343 430 23377
rect 245 23305 430 23343
rect 245 23271 320 23305
rect 354 23271 430 23305
rect 245 23233 430 23271
rect 245 23199 320 23233
rect 354 23199 430 23233
rect 245 23161 430 23199
rect 245 23127 320 23161
rect 354 23127 430 23161
rect 245 23089 430 23127
rect 245 23055 320 23089
rect 354 23055 430 23089
rect 245 23017 430 23055
rect 245 22983 320 23017
rect 354 22983 430 23017
rect 245 22945 430 22983
rect 245 22911 320 22945
rect 354 22911 430 22945
rect 245 22873 430 22911
rect 245 22839 320 22873
rect 354 22839 430 22873
rect 245 22801 430 22839
rect 245 22767 320 22801
rect 354 22767 430 22801
rect 245 22729 430 22767
rect 245 22695 320 22729
rect 354 22695 430 22729
rect 245 22657 430 22695
rect 245 22623 320 22657
rect 354 22623 430 22657
rect 245 22585 430 22623
rect 245 22551 320 22585
rect 354 22551 430 22585
rect 245 22513 430 22551
rect 245 22479 320 22513
rect 354 22479 430 22513
rect 245 22441 430 22479
rect 245 22407 320 22441
rect 354 22407 430 22441
rect 245 22369 430 22407
rect 245 22335 320 22369
rect 354 22335 430 22369
rect 245 22297 430 22335
rect 245 22263 320 22297
rect 354 22263 430 22297
rect 245 22225 430 22263
rect 245 22191 320 22225
rect 354 22191 430 22225
rect 245 22153 430 22191
rect 245 22119 320 22153
rect 354 22119 430 22153
rect 245 22081 430 22119
rect 245 22047 320 22081
rect 354 22047 430 22081
rect 245 22009 430 22047
rect 245 21975 320 22009
rect 354 21975 430 22009
rect 245 21937 430 21975
rect 245 21903 320 21937
rect 354 21903 430 21937
rect 245 21865 430 21903
rect 245 21831 320 21865
rect 354 21831 430 21865
rect 245 21793 430 21831
rect 245 21759 320 21793
rect 354 21759 430 21793
rect 245 21721 430 21759
rect 245 21687 320 21721
rect 354 21687 430 21721
rect 245 21649 430 21687
rect 245 21615 320 21649
rect 354 21615 430 21649
rect 245 21577 430 21615
rect 245 21543 320 21577
rect 354 21543 430 21577
rect 245 21505 430 21543
rect 245 21471 320 21505
rect 354 21471 430 21505
rect 245 21433 430 21471
rect 245 21399 320 21433
rect 354 21399 430 21433
rect 245 21361 430 21399
rect 245 21327 320 21361
rect 354 21327 430 21361
rect 245 21289 430 21327
rect 245 21255 320 21289
rect 354 21255 430 21289
rect 245 21217 430 21255
rect 245 21183 320 21217
rect 354 21183 430 21217
rect 245 21145 430 21183
rect 245 21111 320 21145
rect 354 21111 430 21145
rect 245 21073 430 21111
rect 245 21039 320 21073
rect 354 21039 430 21073
rect 245 21001 430 21039
rect 245 20967 320 21001
rect 354 20967 430 21001
rect 245 20929 430 20967
rect 245 20895 320 20929
rect 354 20895 430 20929
rect 245 20857 430 20895
rect 245 20823 320 20857
rect 354 20823 430 20857
rect 245 20785 430 20823
rect 245 20751 320 20785
rect 354 20751 430 20785
rect 245 20713 430 20751
rect 245 20679 320 20713
rect 354 20679 430 20713
rect 245 20641 430 20679
rect 245 20607 320 20641
rect 354 20607 430 20641
rect 245 20569 430 20607
rect 245 20535 320 20569
rect 354 20535 430 20569
rect 245 20497 430 20535
rect 245 20463 320 20497
rect 354 20463 430 20497
rect 245 20425 430 20463
rect 245 20391 320 20425
rect 354 20391 430 20425
rect 245 20353 430 20391
rect 245 20319 320 20353
rect 354 20319 430 20353
rect 245 20281 430 20319
rect 245 20247 320 20281
rect 354 20247 430 20281
rect 245 20209 430 20247
rect 245 20175 320 20209
rect 354 20175 430 20209
rect 245 20137 430 20175
rect 245 20103 320 20137
rect 354 20103 430 20137
rect 245 20065 430 20103
rect 245 20031 320 20065
rect 354 20031 430 20065
rect 245 19993 430 20031
rect 245 19959 320 19993
rect 354 19959 430 19993
rect 245 19921 430 19959
rect 245 19887 320 19921
rect 354 19887 430 19921
rect 245 19849 430 19887
rect 245 19815 320 19849
rect 354 19815 430 19849
rect 245 19777 430 19815
rect 245 19743 320 19777
rect 354 19743 430 19777
rect 245 19705 430 19743
rect 245 19671 320 19705
rect 354 19671 430 19705
rect 245 19633 430 19671
rect 245 19599 320 19633
rect 354 19599 430 19633
rect 245 19561 430 19599
rect 245 19527 320 19561
rect 354 19527 430 19561
rect 245 19489 430 19527
rect 245 19455 320 19489
rect 354 19455 430 19489
rect 245 19417 430 19455
rect 245 19383 320 19417
rect 354 19383 430 19417
rect 245 19345 430 19383
rect 245 19311 320 19345
rect 354 19311 430 19345
rect 245 19273 430 19311
rect 245 19239 320 19273
rect 354 19239 430 19273
rect 245 19201 430 19239
rect 245 19167 320 19201
rect 354 19167 430 19201
rect 245 19129 430 19167
rect 245 19095 320 19129
rect 354 19095 430 19129
rect 245 19057 430 19095
rect 245 19023 320 19057
rect 354 19023 430 19057
rect 245 18985 430 19023
rect 245 18951 320 18985
rect 354 18951 430 18985
rect 245 18913 430 18951
rect 245 18879 320 18913
rect 354 18879 430 18913
rect 245 18841 430 18879
rect 245 18807 320 18841
rect 354 18807 430 18841
rect 245 18769 430 18807
rect 245 18735 320 18769
rect 354 18735 430 18769
rect 245 18697 430 18735
rect 245 18663 320 18697
rect 354 18663 430 18697
rect 245 18625 430 18663
rect 245 18591 320 18625
rect 354 18591 430 18625
rect 245 18553 430 18591
rect 245 18519 320 18553
rect 354 18519 430 18553
rect 245 18481 430 18519
rect 245 18447 320 18481
rect 354 18447 430 18481
rect 245 18409 430 18447
rect 245 18375 320 18409
rect 354 18375 430 18409
rect 245 18337 430 18375
rect 245 18303 320 18337
rect 354 18303 430 18337
rect 245 18265 430 18303
rect 245 18231 320 18265
rect 354 18231 430 18265
rect 245 18193 430 18231
rect 245 18159 320 18193
rect 354 18159 430 18193
rect 245 18121 430 18159
rect 245 18087 320 18121
rect 354 18087 430 18121
rect 245 18049 430 18087
rect 245 18015 320 18049
rect 354 18015 430 18049
rect 245 17977 430 18015
rect 245 17943 320 17977
rect 354 17943 430 17977
rect 245 17905 430 17943
rect 245 17871 320 17905
rect 354 17871 430 17905
rect 245 17833 430 17871
rect 245 17799 320 17833
rect 354 17799 430 17833
rect 245 17761 430 17799
rect 245 17727 320 17761
rect 354 17727 430 17761
rect 245 17689 430 17727
rect 245 17655 320 17689
rect 354 17655 430 17689
rect 245 17617 430 17655
rect 245 17583 320 17617
rect 354 17583 430 17617
rect 245 17545 430 17583
rect 245 17511 320 17545
rect 354 17511 430 17545
rect 245 17473 430 17511
rect 245 17439 320 17473
rect 354 17439 430 17473
rect 245 17401 430 17439
rect 245 17367 320 17401
rect 354 17367 430 17401
rect 245 17329 430 17367
rect 245 17295 320 17329
rect 354 17295 430 17329
rect 245 17257 430 17295
rect 245 17223 320 17257
rect 354 17223 430 17257
rect 245 17185 430 17223
rect 245 17151 320 17185
rect 354 17151 430 17185
rect 245 17113 430 17151
rect 245 17079 320 17113
rect 354 17079 430 17113
rect 245 17041 430 17079
rect 245 17007 320 17041
rect 354 17007 430 17041
rect 245 16969 430 17007
rect 245 16935 320 16969
rect 354 16935 430 16969
rect 245 16897 430 16935
rect 245 16863 320 16897
rect 354 16863 430 16897
rect 245 16825 430 16863
rect 245 16791 320 16825
rect 354 16791 430 16825
rect 245 16753 430 16791
rect 245 16719 320 16753
rect 354 16719 430 16753
rect 245 16681 430 16719
rect 245 16647 320 16681
rect 354 16647 430 16681
rect 245 16609 430 16647
rect 245 16575 320 16609
rect 354 16575 430 16609
rect 245 16537 430 16575
rect 245 16503 320 16537
rect 354 16503 430 16537
rect 245 16465 430 16503
rect 245 16431 320 16465
rect 354 16431 430 16465
rect 245 16393 430 16431
rect 245 16359 320 16393
rect 354 16359 430 16393
rect 245 16321 430 16359
rect 245 16287 320 16321
rect 354 16287 430 16321
rect 245 16249 430 16287
rect 245 16215 320 16249
rect 354 16215 430 16249
rect 245 16177 430 16215
rect 245 16143 320 16177
rect 354 16143 430 16177
rect 245 16105 430 16143
rect 245 16071 320 16105
rect 354 16071 430 16105
rect 245 16033 430 16071
rect 245 15999 320 16033
rect 354 15999 430 16033
rect 245 15961 430 15999
rect 245 15927 320 15961
rect 354 15927 430 15961
rect 245 15889 430 15927
rect 245 15855 320 15889
rect 354 15855 430 15889
rect 245 15817 430 15855
rect 245 15783 320 15817
rect 354 15783 430 15817
rect 245 15745 430 15783
rect 245 15711 320 15745
rect 354 15711 430 15745
rect 245 15673 430 15711
rect 245 15639 320 15673
rect 354 15639 430 15673
rect 245 15601 430 15639
rect 245 15567 320 15601
rect 354 15567 430 15601
rect 245 15529 430 15567
rect 245 15495 320 15529
rect 354 15495 430 15529
rect 245 15457 430 15495
rect 245 15423 320 15457
rect 354 15423 430 15457
rect 245 15385 430 15423
rect 245 15351 320 15385
rect 354 15351 430 15385
rect 245 15313 430 15351
rect 245 15279 320 15313
rect 354 15279 430 15313
rect 245 15241 430 15279
rect 245 15207 320 15241
rect 354 15207 430 15241
rect 245 15169 430 15207
rect 245 15135 320 15169
rect 354 15135 430 15169
rect 245 15097 430 15135
rect 245 15063 320 15097
rect 354 15063 430 15097
rect 245 15025 430 15063
rect 245 14991 320 15025
rect 354 14991 430 15025
rect 245 14953 430 14991
rect 245 14919 320 14953
rect 354 14919 430 14953
rect 245 14881 430 14919
rect 245 14847 320 14881
rect 354 14847 430 14881
rect 245 14809 430 14847
rect 245 14775 320 14809
rect 354 14775 430 14809
rect 245 14737 430 14775
rect 245 14703 320 14737
rect 354 14703 430 14737
rect 245 14665 430 14703
rect 245 14631 320 14665
rect 354 14631 430 14665
rect 245 14593 430 14631
rect 245 14559 320 14593
rect 354 14559 430 14593
rect 245 14521 430 14559
rect 245 14487 320 14521
rect 354 14487 430 14521
rect 245 14449 430 14487
rect 245 14415 320 14449
rect 354 14415 430 14449
rect 245 14377 430 14415
rect 245 14343 320 14377
rect 354 14343 430 14377
rect 245 14305 430 14343
rect 245 14271 320 14305
rect 354 14271 430 14305
rect 245 14233 430 14271
rect 245 14199 320 14233
rect 354 14199 430 14233
rect 245 14161 430 14199
rect 245 14127 320 14161
rect 354 14127 430 14161
rect 245 14089 430 14127
rect 245 14055 320 14089
rect 354 14055 430 14089
rect 245 14017 430 14055
rect 245 13983 320 14017
rect 354 13983 430 14017
rect 245 13945 430 13983
rect 245 13911 320 13945
rect 354 13911 430 13945
rect 245 13873 430 13911
rect 245 13839 320 13873
rect 354 13839 430 13873
rect 245 13801 430 13839
rect 245 13767 320 13801
rect 354 13767 430 13801
rect 245 13729 430 13767
rect 245 13695 320 13729
rect 354 13695 430 13729
rect 245 13657 430 13695
rect 245 13623 320 13657
rect 354 13623 430 13657
rect 245 13585 430 13623
rect 245 13551 320 13585
rect 354 13551 430 13585
rect 245 13513 430 13551
rect 245 13479 320 13513
rect 354 13479 430 13513
rect 245 13441 430 13479
rect 245 13407 320 13441
rect 354 13407 430 13441
rect 245 13369 430 13407
rect 245 13335 320 13369
rect 354 13335 430 13369
rect 245 13297 430 13335
rect 245 13263 320 13297
rect 354 13263 430 13297
rect 245 13225 430 13263
rect 245 13191 320 13225
rect 354 13191 430 13225
rect 245 13153 430 13191
rect 245 13119 320 13153
rect 354 13119 430 13153
rect 245 13081 430 13119
rect 245 13047 320 13081
rect 354 13047 430 13081
rect 245 13009 430 13047
rect 245 12975 320 13009
rect 354 12975 430 13009
rect 245 12937 430 12975
rect 245 12903 320 12937
rect 354 12903 430 12937
rect 245 12865 430 12903
rect 245 12831 320 12865
rect 354 12831 430 12865
rect 245 12793 430 12831
rect 245 12759 320 12793
rect 354 12759 430 12793
rect 245 12721 430 12759
rect 245 12687 320 12721
rect 354 12687 430 12721
rect 245 12649 430 12687
rect 245 12615 320 12649
rect 354 12615 430 12649
rect 245 12577 430 12615
rect 245 12543 320 12577
rect 354 12543 430 12577
rect 245 12505 430 12543
rect 245 12471 320 12505
rect 354 12471 430 12505
rect 245 12433 430 12471
rect 245 12399 320 12433
rect 354 12399 430 12433
rect 245 12361 430 12399
rect 245 12327 320 12361
rect 354 12327 430 12361
rect 245 12289 430 12327
rect 245 12255 320 12289
rect 354 12255 430 12289
rect 245 12217 430 12255
rect 245 12183 320 12217
rect 354 12183 430 12217
rect 245 12145 430 12183
rect 245 12111 320 12145
rect 354 12111 430 12145
rect 245 12073 430 12111
rect 245 12039 320 12073
rect 354 12039 430 12073
rect 245 12001 430 12039
rect 245 11967 320 12001
rect 354 11967 430 12001
rect 245 11929 430 11967
rect 245 11895 320 11929
rect 354 11895 430 11929
rect 245 11857 430 11895
rect 245 11823 320 11857
rect 354 11823 430 11857
rect 245 11785 430 11823
rect 245 11751 320 11785
rect 354 11751 430 11785
rect 245 11713 430 11751
rect 245 11679 320 11713
rect 354 11679 430 11713
rect 245 11641 430 11679
rect 245 11607 320 11641
rect 354 11607 430 11641
rect 245 11569 430 11607
rect 245 11535 320 11569
rect 354 11535 430 11569
rect 245 11497 430 11535
rect 245 11463 320 11497
rect 354 11463 430 11497
rect 245 11425 430 11463
rect 245 11391 320 11425
rect 354 11391 430 11425
rect 245 11353 430 11391
rect 245 11319 320 11353
rect 354 11319 430 11353
rect 245 11281 430 11319
rect 245 11247 320 11281
rect 354 11247 430 11281
rect 245 11209 430 11247
rect 245 11175 320 11209
rect 354 11175 430 11209
rect 245 11137 430 11175
rect 245 11103 320 11137
rect 354 11103 430 11137
rect 245 11065 430 11103
rect 245 11031 320 11065
rect 354 11031 430 11065
rect 245 10993 430 11031
rect 245 10959 320 10993
rect 354 10959 430 10993
rect 245 10921 430 10959
rect 245 10887 320 10921
rect 354 10887 430 10921
rect 245 10849 430 10887
rect 245 10815 320 10849
rect 354 10815 430 10849
rect 245 10777 430 10815
rect 245 10743 320 10777
rect 354 10743 430 10777
rect 245 10705 430 10743
rect 245 10671 320 10705
rect 354 10671 430 10705
rect 245 10633 430 10671
rect 245 10599 320 10633
rect 354 10599 430 10633
rect 245 10561 430 10599
rect 245 10527 320 10561
rect 354 10527 430 10561
rect 245 10489 430 10527
rect 245 10455 320 10489
rect 354 10455 430 10489
rect 245 10417 430 10455
rect 245 10383 320 10417
rect 354 10383 430 10417
rect 245 10345 430 10383
rect 245 10311 320 10345
rect 354 10311 430 10345
rect 245 10273 430 10311
rect 245 10239 320 10273
rect 354 10239 430 10273
rect 245 10201 430 10239
rect 245 10167 320 10201
rect 354 10167 430 10201
rect 245 10129 430 10167
rect 245 10095 320 10129
rect 354 10095 430 10129
rect 245 10057 430 10095
rect 245 10023 320 10057
rect 354 10023 430 10057
rect 245 9985 430 10023
rect 245 9951 320 9985
rect 354 9951 430 9985
rect 245 9913 430 9951
tri 757 35953 773 35969 se
rect 773 35953 14198 35969
tri 14198 35953 14219 35974 sw
rect 757 35933 14219 35953
rect 757 35902 886 35933
tri 886 35902 917 35933 nw
tri 14059 35902 14090 35933 ne
rect 14090 35902 14219 35933
rect 757 35884 877 35902
tri 877 35893 886 35902 nw
tri 14090 35893 14099 35902 ne
rect 757 35850 807 35884
rect 841 35850 877 35884
rect 757 35812 877 35850
rect 757 35778 807 35812
rect 841 35778 877 35812
rect 757 35740 877 35778
rect 757 35706 807 35740
rect 841 35706 877 35740
rect 757 35668 877 35706
rect 757 35634 807 35668
rect 841 35634 877 35668
rect 757 35596 877 35634
rect 757 35562 807 35596
rect 841 35562 877 35596
rect 757 35524 877 35562
rect 757 35490 807 35524
rect 841 35490 877 35524
rect 757 35452 877 35490
rect 757 35418 807 35452
rect 841 35418 877 35452
rect 757 35380 877 35418
rect 757 35346 807 35380
rect 841 35346 877 35380
rect 757 35308 877 35346
rect 757 35274 807 35308
rect 841 35274 877 35308
rect 757 35236 877 35274
rect 757 35202 807 35236
rect 841 35202 877 35236
rect 757 35164 877 35202
rect 757 35130 807 35164
rect 841 35130 877 35164
rect 757 35092 877 35130
rect 757 35058 807 35092
rect 841 35058 877 35092
rect 757 35020 877 35058
rect 757 34986 807 35020
rect 841 34986 877 35020
rect 757 34948 877 34986
rect 757 34914 807 34948
rect 841 34914 877 34948
rect 757 34876 877 34914
rect 757 34842 807 34876
rect 841 34842 877 34876
rect 757 34804 877 34842
rect 757 34770 807 34804
rect 841 34770 877 34804
rect 757 34732 877 34770
rect 757 34698 807 34732
rect 841 34698 877 34732
rect 14099 35805 14219 35902
rect 14099 35771 14122 35805
rect 14156 35771 14219 35805
rect 14099 35733 14219 35771
rect 14099 35699 14122 35733
rect 14156 35699 14219 35733
rect 14099 35661 14219 35699
rect 14099 35627 14122 35661
rect 14156 35627 14219 35661
rect 14099 35589 14219 35627
rect 14099 35555 14122 35589
rect 14156 35555 14219 35589
rect 14099 35517 14219 35555
rect 14099 35483 14122 35517
rect 14156 35483 14219 35517
rect 14099 35445 14219 35483
rect 14099 35411 14122 35445
rect 14156 35411 14219 35445
rect 14099 35373 14219 35411
rect 14099 35339 14122 35373
rect 14156 35339 14219 35373
rect 14099 35301 14219 35339
rect 14099 35267 14122 35301
rect 14156 35267 14219 35301
rect 14099 35229 14219 35267
rect 14099 35195 14122 35229
rect 14156 35195 14219 35229
rect 14099 35157 14219 35195
rect 14099 35123 14122 35157
rect 14156 35123 14219 35157
rect 14099 35085 14219 35123
rect 14099 35051 14122 35085
rect 14156 35051 14219 35085
rect 14099 35013 14219 35051
rect 14099 34979 14122 35013
rect 14156 34979 14219 35013
rect 14099 34941 14219 34979
rect 14099 34907 14122 34941
rect 14156 34907 14219 34941
rect 14099 34869 14219 34907
rect 14099 34835 14122 34869
rect 14156 34835 14219 34869
rect 14099 34797 14219 34835
rect 14099 34763 14122 34797
rect 14156 34763 14219 34797
rect 14099 34725 14219 34763
rect 757 34660 877 34698
rect 757 34626 807 34660
rect 841 34626 877 34660
rect 757 34588 877 34626
rect 757 34554 807 34588
rect 841 34554 877 34588
rect 757 34516 877 34554
rect 757 34482 807 34516
rect 841 34482 877 34516
rect 757 34444 877 34482
rect 757 34410 807 34444
rect 841 34410 877 34444
rect 757 34372 877 34410
rect 757 34338 807 34372
rect 841 34338 877 34372
rect 757 34300 877 34338
rect 757 34266 807 34300
rect 841 34266 877 34300
rect 757 34228 877 34266
rect 757 34194 807 34228
rect 841 34194 877 34228
rect 757 34156 877 34194
rect 757 34122 807 34156
rect 841 34122 877 34156
rect 757 34084 877 34122
rect 757 34050 807 34084
rect 841 34050 877 34084
rect 757 34012 877 34050
rect 757 33978 807 34012
rect 841 33978 877 34012
rect 757 33940 877 33978
rect 757 33906 807 33940
rect 841 33906 877 33940
rect 757 33868 877 33906
rect 757 33834 807 33868
rect 841 33834 877 33868
rect 757 33796 877 33834
rect 757 33762 807 33796
rect 841 33762 877 33796
rect 757 33724 877 33762
rect 757 33690 807 33724
rect 841 33690 877 33724
rect 757 33652 877 33690
rect 757 33618 807 33652
rect 841 33618 877 33652
rect 757 33580 877 33618
rect 757 33546 807 33580
rect 841 33546 877 33580
rect 757 33508 877 33546
rect 757 33474 807 33508
rect 841 33474 877 33508
rect 757 33436 877 33474
rect 757 33402 807 33436
rect 841 33402 877 33436
rect 757 33364 877 33402
rect 757 33330 807 33364
rect 841 33330 877 33364
rect 757 33292 877 33330
rect 757 33258 807 33292
rect 841 33258 877 33292
rect 757 33220 877 33258
rect 757 33186 807 33220
rect 841 33186 877 33220
rect 757 33148 877 33186
rect 757 33114 807 33148
rect 841 33114 877 33148
rect 757 33076 877 33114
rect 757 33042 807 33076
rect 841 33042 877 33076
rect 757 33004 877 33042
rect 757 32970 807 33004
rect 841 32970 877 33004
rect 757 32932 877 32970
rect 757 32898 807 32932
rect 841 32898 877 32932
rect 757 32860 877 32898
rect 757 32826 807 32860
rect 841 32826 877 32860
rect 757 32788 877 32826
rect 757 32754 807 32788
rect 841 32754 877 32788
rect 757 32716 877 32754
rect 757 32682 807 32716
rect 841 32682 877 32716
rect 757 32644 877 32682
rect 757 32610 807 32644
rect 841 32610 877 32644
rect 757 32572 877 32610
rect 757 32538 807 32572
rect 841 32538 877 32572
rect 757 32500 877 32538
rect 757 32466 807 32500
rect 841 32466 877 32500
rect 757 32428 877 32466
rect 757 32394 807 32428
rect 841 32394 877 32428
rect 757 32356 877 32394
rect 757 32322 807 32356
rect 841 32322 877 32356
rect 757 32284 877 32322
rect 757 32250 807 32284
rect 841 32250 877 32284
rect 757 32212 877 32250
rect 757 32178 807 32212
rect 841 32178 877 32212
rect 757 32140 877 32178
rect 757 32106 807 32140
rect 841 32106 877 32140
rect 757 32068 877 32106
rect 757 32034 807 32068
rect 841 32034 877 32068
rect 757 31996 877 32034
rect 757 31962 807 31996
rect 841 31962 877 31996
rect 757 31924 877 31962
rect 757 31890 807 31924
rect 841 31890 877 31924
rect 757 31852 877 31890
rect 757 31818 807 31852
rect 841 31818 877 31852
rect 757 31780 877 31818
rect 757 31746 807 31780
rect 841 31746 877 31780
rect 757 31708 877 31746
rect 757 31674 807 31708
rect 841 31674 877 31708
rect 757 31636 877 31674
rect 757 31602 807 31636
rect 841 31602 877 31636
rect 757 31564 877 31602
rect 757 31530 807 31564
rect 841 31530 877 31564
rect 757 31492 877 31530
rect 757 31458 807 31492
rect 841 31458 877 31492
rect 757 31420 877 31458
rect 757 31386 807 31420
rect 841 31386 877 31420
rect 757 31348 877 31386
rect 757 31314 807 31348
rect 841 31314 877 31348
rect 757 31276 877 31314
rect 757 31242 807 31276
rect 841 31242 877 31276
rect 757 31204 877 31242
rect 757 31170 807 31204
rect 841 31170 877 31204
rect 757 31132 877 31170
rect 757 31098 807 31132
rect 841 31098 877 31132
rect 757 31060 877 31098
rect 757 31026 807 31060
rect 841 31026 877 31060
rect 757 30988 877 31026
rect 757 30954 807 30988
rect 841 30954 877 30988
rect 757 30916 877 30954
rect 757 30882 807 30916
rect 841 30882 877 30916
rect 757 30844 877 30882
rect 757 30810 807 30844
rect 841 30810 877 30844
rect 757 30772 877 30810
rect 757 30738 807 30772
rect 841 30738 877 30772
rect 757 30700 877 30738
rect 757 30666 807 30700
rect 841 30666 877 30700
rect 757 30628 877 30666
rect 757 30594 807 30628
rect 841 30594 877 30628
rect 757 30556 877 30594
rect 757 30522 807 30556
rect 841 30522 877 30556
rect 757 30484 877 30522
rect 757 30450 807 30484
rect 841 30450 877 30484
rect 757 30412 877 30450
rect 757 30378 807 30412
rect 841 30378 877 30412
rect 757 30340 877 30378
rect 757 30306 807 30340
rect 841 30306 877 30340
rect 757 30268 877 30306
rect 757 30234 807 30268
rect 841 30234 877 30268
rect 757 30196 877 30234
rect 757 30162 807 30196
rect 841 30162 877 30196
rect 757 30124 877 30162
rect 757 30090 807 30124
rect 841 30090 877 30124
rect 757 30052 877 30090
rect 757 30018 807 30052
rect 841 30018 877 30052
rect 757 29980 877 30018
rect 757 29946 807 29980
rect 841 29946 877 29980
rect 757 29908 877 29946
rect 757 29874 807 29908
rect 841 29874 877 29908
rect 757 29836 877 29874
rect 757 29802 807 29836
rect 841 29802 877 29836
rect 757 29764 877 29802
rect 757 29730 807 29764
rect 841 29730 877 29764
rect 757 29692 877 29730
rect 757 29658 807 29692
rect 841 29658 877 29692
rect 757 29620 877 29658
rect 757 29586 807 29620
rect 841 29586 877 29620
rect 757 29548 877 29586
rect 757 29514 807 29548
rect 841 29514 877 29548
rect 757 29476 877 29514
rect 757 29442 807 29476
rect 841 29442 877 29476
rect 757 29404 877 29442
rect 757 29370 807 29404
rect 841 29370 877 29404
rect 757 29332 877 29370
rect 757 29298 807 29332
rect 841 29298 877 29332
rect 757 29260 877 29298
rect 757 29226 807 29260
rect 841 29226 877 29260
rect 757 29188 877 29226
rect 757 29154 807 29188
rect 841 29154 877 29188
rect 757 29116 877 29154
rect 757 29082 807 29116
rect 841 29082 877 29116
rect 757 29044 877 29082
rect 757 29010 807 29044
rect 841 29010 877 29044
rect 757 28972 877 29010
rect 757 28938 807 28972
rect 841 28938 877 28972
rect 757 28900 877 28938
rect 757 28866 807 28900
rect 841 28866 877 28900
rect 757 28828 877 28866
rect 757 28794 807 28828
rect 841 28794 877 28828
rect 757 28756 877 28794
rect 757 28722 807 28756
rect 841 28722 877 28756
rect 757 28684 877 28722
rect 757 28650 807 28684
rect 841 28650 877 28684
rect 757 28612 877 28650
rect 757 28578 807 28612
rect 841 28578 877 28612
rect 757 28540 877 28578
rect 757 28506 807 28540
rect 841 28506 877 28540
rect 757 28468 877 28506
rect 757 28434 807 28468
rect 841 28434 877 28468
rect 757 28396 877 28434
rect 757 28362 807 28396
rect 841 28362 877 28396
rect 757 28324 877 28362
rect 757 28290 807 28324
rect 841 28290 877 28324
rect 757 28252 877 28290
rect 757 28218 807 28252
rect 841 28218 877 28252
rect 757 28180 877 28218
rect 757 28146 807 28180
rect 841 28146 877 28180
rect 757 28108 877 28146
rect 757 28074 807 28108
rect 841 28074 877 28108
rect 757 28036 877 28074
rect 757 28002 807 28036
rect 841 28002 877 28036
rect 757 27964 877 28002
rect 757 27930 807 27964
rect 841 27930 877 27964
rect 757 27892 877 27930
rect 757 27858 807 27892
rect 841 27858 877 27892
rect 757 27820 877 27858
rect 757 27786 807 27820
rect 841 27786 877 27820
rect 757 27748 877 27786
rect 757 27714 807 27748
rect 841 27714 877 27748
rect 757 27676 877 27714
rect 757 27642 807 27676
rect 841 27642 877 27676
rect 757 27604 877 27642
rect 757 27570 807 27604
rect 841 27570 877 27604
rect 757 27532 877 27570
rect 757 27498 807 27532
rect 841 27498 877 27532
rect 757 27460 877 27498
rect 757 27426 807 27460
rect 841 27426 877 27460
rect 757 27388 877 27426
rect 757 27354 807 27388
rect 841 27354 877 27388
rect 757 27316 877 27354
rect 757 27282 807 27316
rect 841 27282 877 27316
rect 757 27244 877 27282
rect 757 27210 807 27244
rect 841 27210 877 27244
rect 757 27172 877 27210
rect 757 27138 807 27172
rect 841 27138 877 27172
rect 757 27100 877 27138
rect 757 27066 807 27100
rect 841 27066 877 27100
rect 757 27028 877 27066
rect 757 26994 807 27028
rect 841 26994 877 27028
rect 757 26956 877 26994
rect 757 26922 807 26956
rect 841 26922 877 26956
rect 757 26884 877 26922
rect 757 26850 807 26884
rect 841 26850 877 26884
rect 757 26812 877 26850
rect 757 26778 807 26812
rect 841 26778 877 26812
rect 757 26740 877 26778
rect 757 26706 807 26740
rect 841 26706 877 26740
rect 757 26668 877 26706
rect 757 26634 807 26668
rect 841 26634 877 26668
rect 757 26596 877 26634
rect 757 26562 807 26596
rect 841 26562 877 26596
rect 757 26524 877 26562
rect 757 26490 807 26524
rect 841 26490 877 26524
rect 757 26452 877 26490
rect 757 26418 807 26452
rect 841 26418 877 26452
rect 757 26380 877 26418
rect 757 26346 807 26380
rect 841 26346 877 26380
rect 757 26308 877 26346
rect 757 26274 807 26308
rect 841 26274 877 26308
rect 757 26236 877 26274
rect 757 26202 807 26236
rect 841 26202 877 26236
rect 757 26164 877 26202
rect 757 26130 807 26164
rect 841 26130 877 26164
rect 757 26092 877 26130
rect 757 26058 807 26092
rect 841 26058 877 26092
rect 757 26020 877 26058
rect 757 25986 807 26020
rect 841 25986 877 26020
rect 757 25948 877 25986
rect 757 25914 807 25948
rect 841 25914 877 25948
rect 757 25876 877 25914
rect 757 25842 807 25876
rect 841 25842 877 25876
rect 757 25804 877 25842
rect 757 25770 807 25804
rect 841 25770 877 25804
rect 757 25732 877 25770
rect 757 25698 807 25732
rect 841 25698 877 25732
rect 757 25660 877 25698
rect 757 25626 807 25660
rect 841 25626 877 25660
rect 757 25588 877 25626
rect 757 25554 807 25588
rect 841 25554 877 25588
rect 757 25516 877 25554
rect 757 25482 807 25516
rect 841 25482 877 25516
rect 757 25444 877 25482
rect 757 25410 807 25444
rect 841 25410 877 25444
rect 757 25372 877 25410
rect 757 25338 807 25372
rect 841 25338 877 25372
rect 757 25300 877 25338
rect 757 25266 807 25300
rect 841 25266 877 25300
rect 757 25228 877 25266
rect 757 25194 807 25228
rect 841 25194 877 25228
rect 757 25156 877 25194
rect 757 25122 807 25156
rect 841 25122 877 25156
rect 757 25084 877 25122
rect 757 25050 807 25084
rect 841 25050 877 25084
rect 757 25012 877 25050
rect 757 24978 807 25012
rect 841 24978 877 25012
rect 757 24940 877 24978
rect 757 24906 807 24940
rect 841 24906 877 24940
rect 757 24868 877 24906
rect 757 24834 807 24868
rect 841 24834 877 24868
rect 757 24796 877 24834
rect 757 24762 807 24796
rect 841 24762 877 24796
rect 757 24724 877 24762
rect 757 24690 807 24724
rect 841 24690 877 24724
rect 757 24652 877 24690
rect 757 24618 807 24652
rect 841 24618 877 24652
rect 757 24580 877 24618
rect 757 24546 807 24580
rect 841 24546 877 24580
rect 757 24508 877 24546
rect 757 24474 807 24508
rect 841 24474 877 24508
rect 757 24436 877 24474
rect 757 24402 807 24436
rect 841 24402 877 24436
rect 757 24364 877 24402
rect 757 24330 807 24364
rect 841 24330 877 24364
rect 757 24292 877 24330
rect 757 24258 807 24292
rect 841 24258 877 24292
rect 757 24220 877 24258
rect 757 24186 807 24220
rect 841 24186 877 24220
rect 757 24148 877 24186
rect 757 24114 807 24148
rect 841 24114 877 24148
rect 757 24076 877 24114
rect 757 24042 807 24076
rect 841 24042 877 24076
rect 757 24004 877 24042
rect 757 23970 807 24004
rect 841 23970 877 24004
rect 757 23932 877 23970
rect 757 23898 807 23932
rect 841 23898 877 23932
rect 757 23860 877 23898
rect 757 23826 807 23860
rect 841 23826 877 23860
rect 757 23788 877 23826
rect 757 23754 807 23788
rect 841 23754 877 23788
rect 757 23716 877 23754
rect 757 23682 807 23716
rect 841 23682 877 23716
rect 757 23644 877 23682
rect 757 23610 807 23644
rect 841 23610 877 23644
rect 757 23572 877 23610
rect 757 23538 807 23572
rect 841 23538 877 23572
rect 757 23500 877 23538
rect 757 23466 807 23500
rect 841 23466 877 23500
rect 757 23428 877 23466
rect 757 23394 807 23428
rect 841 23394 877 23428
rect 757 23356 877 23394
rect 757 23322 807 23356
rect 841 23322 877 23356
rect 757 23284 877 23322
rect 757 23250 807 23284
rect 841 23250 877 23284
rect 757 23212 877 23250
rect 757 23178 807 23212
rect 841 23178 877 23212
rect 757 23140 877 23178
rect 757 23106 807 23140
rect 841 23106 877 23140
rect 757 23068 877 23106
rect 757 23034 807 23068
rect 841 23034 877 23068
rect 757 22996 877 23034
rect 757 22962 807 22996
rect 841 22962 877 22996
rect 757 22924 877 22962
rect 757 22890 807 22924
rect 841 22890 877 22924
rect 757 22852 877 22890
rect 757 22818 807 22852
rect 841 22818 877 22852
rect 757 22780 877 22818
rect 757 22746 807 22780
rect 841 22746 877 22780
rect 757 22708 877 22746
rect 757 22674 807 22708
rect 841 22674 877 22708
rect 757 22636 877 22674
rect 757 22602 807 22636
rect 841 22602 877 22636
rect 757 22564 877 22602
rect 757 22530 807 22564
rect 841 22530 877 22564
rect 757 22492 877 22530
rect 757 22458 807 22492
rect 841 22458 877 22492
rect 757 22420 877 22458
rect 757 22386 807 22420
rect 841 22386 877 22420
rect 757 22348 877 22386
rect 757 22314 807 22348
rect 841 22314 877 22348
rect 757 22276 877 22314
rect 757 22242 807 22276
rect 841 22242 877 22276
rect 757 22204 877 22242
rect 757 22170 807 22204
rect 841 22170 877 22204
rect 757 22132 877 22170
rect 757 22098 807 22132
rect 841 22098 877 22132
rect 757 22060 877 22098
rect 757 22026 807 22060
rect 841 22026 877 22060
rect 757 21988 877 22026
rect 757 21954 807 21988
rect 841 21954 877 21988
rect 757 21916 877 21954
rect 757 21882 807 21916
rect 841 21882 877 21916
rect 757 21844 877 21882
rect 757 21810 807 21844
rect 841 21810 877 21844
rect 757 21772 877 21810
rect 757 21738 807 21772
rect 841 21738 877 21772
rect 757 21700 877 21738
rect 757 21666 807 21700
rect 841 21666 877 21700
rect 757 21628 877 21666
rect 757 21594 807 21628
rect 841 21594 877 21628
rect 757 21556 877 21594
rect 757 21522 807 21556
rect 841 21522 877 21556
rect 757 21484 877 21522
rect 757 21450 807 21484
rect 841 21450 877 21484
rect 757 21412 877 21450
rect 757 21378 807 21412
rect 841 21378 877 21412
rect 757 21340 877 21378
rect 757 21306 807 21340
rect 841 21306 877 21340
rect 757 21268 877 21306
rect 757 21234 807 21268
rect 841 21234 877 21268
rect 757 21196 877 21234
rect 757 21162 807 21196
rect 841 21162 877 21196
rect 757 21124 877 21162
rect 757 21090 807 21124
rect 841 21090 877 21124
rect 757 21052 877 21090
rect 757 21018 807 21052
rect 841 21018 877 21052
rect 757 20980 877 21018
rect 757 20946 807 20980
rect 841 20946 877 20980
rect 757 20908 877 20946
rect 757 20874 807 20908
rect 841 20874 877 20908
rect 757 20836 877 20874
rect 757 20802 807 20836
rect 841 20802 877 20836
rect 757 20764 877 20802
rect 757 20730 807 20764
rect 841 20730 877 20764
rect 757 20692 877 20730
rect 757 20658 807 20692
rect 841 20658 877 20692
rect 757 20620 877 20658
rect 757 20586 807 20620
rect 841 20586 877 20620
rect 757 20548 877 20586
rect 757 20514 807 20548
rect 841 20514 877 20548
rect 757 20476 877 20514
rect 757 20442 807 20476
rect 841 20442 877 20476
rect 757 20404 877 20442
rect 757 20370 807 20404
rect 841 20370 877 20404
rect 757 20332 877 20370
rect 757 20298 807 20332
rect 841 20298 877 20332
rect 757 20260 877 20298
rect 757 20226 807 20260
rect 841 20226 877 20260
rect 757 20188 877 20226
rect 757 20154 807 20188
rect 841 20154 877 20188
rect 757 20116 877 20154
rect 757 20082 807 20116
rect 841 20082 877 20116
rect 757 20044 877 20082
rect 757 20010 807 20044
rect 841 20010 877 20044
rect 757 19972 877 20010
rect 757 19938 807 19972
rect 841 19938 877 19972
rect 757 19900 877 19938
rect 757 19866 807 19900
rect 841 19866 877 19900
rect 757 19828 877 19866
rect 757 19794 807 19828
rect 841 19794 877 19828
rect 757 19756 877 19794
rect 757 19722 807 19756
rect 841 19722 877 19756
rect 757 19684 877 19722
rect 757 19650 807 19684
rect 841 19650 877 19684
rect 757 19612 877 19650
rect 757 19578 807 19612
rect 841 19578 877 19612
rect 757 19540 877 19578
rect 757 19506 807 19540
rect 841 19506 877 19540
rect 757 19468 877 19506
rect 757 19434 807 19468
rect 841 19434 877 19468
rect 757 19396 877 19434
rect 757 19362 807 19396
rect 841 19362 877 19396
rect 757 19324 877 19362
rect 757 19290 807 19324
rect 841 19290 877 19324
rect 757 19252 877 19290
rect 757 19218 807 19252
rect 841 19218 877 19252
rect 757 19180 877 19218
rect 757 19146 807 19180
rect 841 19146 877 19180
rect 757 19108 877 19146
rect 757 19074 807 19108
rect 841 19074 877 19108
rect 757 19036 877 19074
rect 757 19002 807 19036
rect 841 19002 877 19036
rect 757 18964 877 19002
rect 757 18930 807 18964
rect 841 18930 877 18964
rect 757 18892 877 18930
rect 757 18858 807 18892
rect 841 18858 877 18892
rect 757 18820 877 18858
rect 757 18786 807 18820
rect 841 18786 877 18820
rect 757 18748 877 18786
rect 757 18714 807 18748
rect 841 18714 877 18748
rect 757 18676 877 18714
rect 757 18642 807 18676
rect 841 18642 877 18676
rect 757 18604 877 18642
rect 757 18570 807 18604
rect 841 18570 877 18604
rect 757 18532 877 18570
rect 757 18498 807 18532
rect 841 18498 877 18532
rect 757 18460 877 18498
rect 757 18426 807 18460
rect 841 18426 877 18460
rect 757 18388 877 18426
rect 757 18354 807 18388
rect 841 18354 877 18388
rect 757 18316 877 18354
rect 757 18282 807 18316
rect 841 18282 877 18316
rect 757 18244 877 18282
rect 757 18210 807 18244
rect 841 18210 877 18244
rect 757 18172 877 18210
rect 757 18138 807 18172
rect 841 18138 877 18172
rect 757 18100 877 18138
rect 757 18066 807 18100
rect 841 18066 877 18100
rect 757 18028 877 18066
rect 757 17994 807 18028
rect 841 17994 877 18028
rect 757 17956 877 17994
rect 757 17922 807 17956
rect 841 17922 877 17956
rect 757 17884 877 17922
rect 757 17850 807 17884
rect 841 17850 877 17884
rect 757 17812 877 17850
rect 757 17778 807 17812
rect 841 17778 877 17812
rect 757 17740 877 17778
rect 757 17706 807 17740
rect 841 17706 877 17740
rect 757 17668 877 17706
rect 757 17634 807 17668
rect 841 17634 877 17668
rect 757 17596 877 17634
rect 757 17562 807 17596
rect 841 17562 877 17596
rect 757 17524 877 17562
rect 757 17490 807 17524
rect 841 17490 877 17524
rect 757 17452 877 17490
rect 757 17418 807 17452
rect 841 17418 877 17452
rect 757 17380 877 17418
rect 757 17346 807 17380
rect 841 17346 877 17380
rect 757 17308 877 17346
rect 757 17274 807 17308
rect 841 17274 877 17308
rect 757 17236 877 17274
rect 757 17202 807 17236
rect 841 17202 877 17236
rect 757 17164 877 17202
rect 757 17130 807 17164
rect 841 17130 877 17164
rect 757 17092 877 17130
rect 757 17058 807 17092
rect 841 17058 877 17092
rect 757 17020 877 17058
rect 757 16986 807 17020
rect 841 16986 877 17020
rect 757 16948 877 16986
rect 757 16914 807 16948
rect 841 16914 877 16948
rect 757 16876 877 16914
rect 757 16842 807 16876
rect 841 16842 877 16876
rect 757 16804 877 16842
rect 757 16770 807 16804
rect 841 16770 877 16804
rect 757 16732 877 16770
rect 757 16698 807 16732
rect 841 16698 877 16732
rect 757 16660 877 16698
rect 757 16626 807 16660
rect 841 16626 877 16660
rect 757 16588 877 16626
rect 757 16554 807 16588
rect 841 16554 877 16588
rect 757 16516 877 16554
rect 757 16482 807 16516
rect 841 16482 877 16516
rect 757 16444 877 16482
rect 757 16410 807 16444
rect 841 16410 877 16444
rect 757 16372 877 16410
rect 757 16338 807 16372
rect 841 16338 877 16372
rect 757 16300 877 16338
rect 757 16266 807 16300
rect 841 16266 877 16300
rect 757 16228 877 16266
rect 757 16194 807 16228
rect 841 16194 877 16228
rect 757 16156 877 16194
rect 757 16122 807 16156
rect 841 16122 877 16156
rect 757 16084 877 16122
rect 757 16050 807 16084
rect 841 16050 877 16084
rect 757 16012 877 16050
rect 757 15978 807 16012
rect 841 15978 877 16012
rect 757 15940 877 15978
rect 757 15906 807 15940
rect 841 15906 877 15940
rect 757 15868 877 15906
rect 757 15834 807 15868
rect 841 15834 877 15868
rect 757 15796 877 15834
rect 757 15762 807 15796
rect 841 15762 877 15796
rect 757 15724 877 15762
rect 757 15690 807 15724
rect 841 15690 877 15724
rect 757 15652 877 15690
rect 757 15618 807 15652
rect 841 15618 877 15652
rect 757 15580 877 15618
rect 757 15546 807 15580
rect 841 15546 877 15580
rect 757 15508 877 15546
rect 757 15474 807 15508
rect 841 15474 877 15508
rect 757 15436 877 15474
rect 757 15402 807 15436
rect 841 15402 877 15436
rect 757 15364 877 15402
rect 757 15330 807 15364
rect 841 15330 877 15364
rect 757 15292 877 15330
rect 757 15258 807 15292
rect 841 15258 877 15292
rect 757 15220 877 15258
rect 757 15186 807 15220
rect 841 15186 877 15220
rect 757 15148 877 15186
rect 757 15114 807 15148
rect 841 15114 877 15148
rect 757 15076 877 15114
rect 757 15042 807 15076
rect 841 15042 877 15076
rect 757 15004 877 15042
rect 757 14970 807 15004
rect 841 14970 877 15004
rect 757 14932 877 14970
rect 757 14898 807 14932
rect 841 14898 877 14932
rect 757 14860 877 14898
rect 757 14826 807 14860
rect 841 14826 877 14860
rect 757 14788 877 14826
rect 757 14754 807 14788
rect 841 14754 877 14788
rect 757 14716 877 14754
rect 757 14682 807 14716
rect 841 14682 877 14716
rect 757 14644 877 14682
rect 757 14610 807 14644
rect 841 14610 877 14644
rect 757 14572 877 14610
rect 757 14538 807 14572
rect 841 14538 877 14572
rect 757 14500 877 14538
rect 757 14466 807 14500
rect 841 14466 877 14500
rect 757 14428 877 14466
rect 757 14394 807 14428
rect 841 14394 877 14428
rect 757 14356 877 14394
rect 757 14322 807 14356
rect 841 14322 877 14356
rect 757 14284 877 14322
rect 757 14250 807 14284
rect 841 14250 877 14284
rect 757 14212 877 14250
rect 757 14178 807 14212
rect 841 14178 877 14212
rect 757 14140 877 14178
rect 757 14106 807 14140
rect 841 14106 877 14140
rect 757 14068 877 14106
rect 757 14034 807 14068
rect 841 14034 877 14068
rect 757 13996 877 14034
rect 757 13962 807 13996
rect 841 13962 877 13996
rect 757 13924 877 13962
rect 757 13890 807 13924
rect 841 13890 877 13924
rect 757 13852 877 13890
rect 757 13818 807 13852
rect 841 13818 877 13852
rect 757 13780 877 13818
rect 757 13746 807 13780
rect 841 13746 877 13780
rect 757 13708 877 13746
rect 757 13674 807 13708
rect 841 13674 877 13708
rect 757 13636 877 13674
rect 757 13602 807 13636
rect 841 13602 877 13636
rect 757 13564 877 13602
rect 757 13530 807 13564
rect 841 13530 877 13564
rect 757 13492 877 13530
rect 757 13458 807 13492
rect 841 13458 877 13492
rect 757 13420 877 13458
rect 757 13386 807 13420
rect 841 13386 877 13420
rect 757 13348 877 13386
rect 757 13314 807 13348
rect 841 13314 877 13348
rect 757 13276 877 13314
rect 757 13242 807 13276
rect 841 13242 877 13276
rect 757 13204 877 13242
rect 757 13170 807 13204
rect 841 13170 877 13204
rect 757 13132 877 13170
rect 757 13098 807 13132
rect 841 13098 877 13132
rect 757 13060 877 13098
rect 757 13026 807 13060
rect 841 13026 877 13060
rect 757 12988 877 13026
rect 757 12954 807 12988
rect 841 12954 877 12988
rect 757 12916 877 12954
rect 757 12882 807 12916
rect 841 12882 877 12916
rect 757 12844 877 12882
rect 757 12810 807 12844
rect 841 12810 877 12844
rect 757 12772 877 12810
rect 757 12738 807 12772
rect 841 12738 877 12772
rect 757 12700 877 12738
rect 757 12666 807 12700
rect 841 12666 877 12700
rect 757 12628 877 12666
rect 757 12594 807 12628
rect 841 12594 877 12628
rect 757 12556 877 12594
rect 757 12522 807 12556
rect 841 12522 877 12556
rect 757 12484 877 12522
rect 757 12450 807 12484
rect 841 12450 877 12484
rect 757 12412 877 12450
rect 757 12378 807 12412
rect 841 12378 877 12412
rect 757 12340 877 12378
rect 757 12306 807 12340
rect 841 12306 877 12340
rect 757 12268 877 12306
rect 757 12234 807 12268
rect 841 12234 877 12268
rect 757 12196 877 12234
rect 757 12162 807 12196
rect 841 12162 877 12196
rect 757 12124 877 12162
rect 757 12090 807 12124
rect 841 12090 877 12124
rect 757 12052 877 12090
rect 757 12018 807 12052
rect 841 12018 877 12052
rect 757 11980 877 12018
rect 757 11946 807 11980
rect 841 11946 877 11980
rect 757 11908 877 11946
rect 757 11874 807 11908
rect 841 11874 877 11908
rect 757 11836 877 11874
rect 757 11802 807 11836
rect 841 11802 877 11836
rect 757 11764 877 11802
rect 757 11730 807 11764
rect 841 11730 877 11764
rect 757 11692 877 11730
rect 757 11658 807 11692
rect 841 11658 877 11692
rect 757 11620 877 11658
rect 757 11586 807 11620
rect 841 11586 877 11620
rect 757 11548 877 11586
rect 757 11514 807 11548
rect 841 11514 877 11548
rect 757 11476 877 11514
rect 757 11442 807 11476
rect 841 11442 877 11476
rect 757 11404 877 11442
rect 757 11370 807 11404
rect 841 11370 877 11404
rect 757 11332 877 11370
rect 757 11298 807 11332
rect 841 11298 877 11332
rect 757 11260 877 11298
rect 757 11226 807 11260
rect 841 11226 877 11260
rect 757 11188 877 11226
rect 757 11154 807 11188
rect 841 11154 877 11188
rect 757 11116 877 11154
rect 757 11082 807 11116
rect 841 11082 877 11116
rect 757 11044 877 11082
rect 757 11010 807 11044
rect 841 11010 877 11044
rect 757 10972 877 11010
rect 757 10938 807 10972
rect 841 10938 877 10972
rect 757 10900 877 10938
rect 757 10866 807 10900
rect 841 10866 877 10900
rect 757 10828 877 10866
rect 757 10794 807 10828
rect 841 10794 877 10828
rect 757 10756 877 10794
rect 757 10722 807 10756
rect 841 10722 877 10756
rect 757 10684 877 10722
rect 757 10650 807 10684
rect 841 10650 877 10684
rect 757 10612 877 10650
rect 757 10578 807 10612
rect 841 10578 877 10612
rect 757 10540 877 10578
rect 757 10506 807 10540
rect 841 10506 877 10540
rect 757 10468 877 10506
rect 757 10434 807 10468
rect 841 10434 877 10468
rect 757 10396 877 10434
rect 757 10362 807 10396
rect 841 10362 877 10396
rect 757 10324 877 10362
rect 757 10290 807 10324
rect 841 10290 877 10324
rect 757 10252 877 10290
rect 757 10218 807 10252
rect 841 10218 877 10252
rect 757 10180 877 10218
rect 1119 34679 13887 34721
rect 1119 34645 1301 34679
rect 1335 34645 1373 34679
rect 1407 34645 1445 34679
rect 1479 34645 1517 34679
rect 1551 34645 1589 34679
rect 1623 34645 1661 34679
rect 1695 34645 1733 34679
rect 1767 34645 1805 34679
rect 1839 34645 1877 34679
rect 1911 34645 1949 34679
rect 1983 34645 2021 34679
rect 2055 34645 2093 34679
rect 2127 34645 2165 34679
rect 2199 34645 2237 34679
rect 2271 34645 2309 34679
rect 2343 34645 2381 34679
rect 2415 34645 2453 34679
rect 2487 34645 2525 34679
rect 2559 34645 2597 34679
rect 2631 34645 2669 34679
rect 2703 34645 2741 34679
rect 2775 34645 2813 34679
rect 2847 34645 2885 34679
rect 2919 34645 2957 34679
rect 2991 34645 3029 34679
rect 3063 34645 3101 34679
rect 3135 34645 3173 34679
rect 3207 34645 3245 34679
rect 3279 34645 3317 34679
rect 3351 34645 3389 34679
rect 3423 34645 3461 34679
rect 3495 34645 3533 34679
rect 3567 34645 3605 34679
rect 3639 34645 3677 34679
rect 3711 34645 3749 34679
rect 3783 34645 3821 34679
rect 3855 34645 3893 34679
rect 3927 34645 3965 34679
rect 3999 34645 4037 34679
rect 4071 34645 4109 34679
rect 4143 34645 4181 34679
rect 4215 34645 4253 34679
rect 4287 34645 4325 34679
rect 4359 34645 4397 34679
rect 4431 34645 4469 34679
rect 4503 34645 4541 34679
rect 4575 34645 4613 34679
rect 4647 34645 4685 34679
rect 4719 34645 4757 34679
rect 4791 34645 4829 34679
rect 4863 34645 4901 34679
rect 4935 34645 4973 34679
rect 5007 34645 5045 34679
rect 5079 34645 5117 34679
rect 5151 34645 5189 34679
rect 5223 34645 5261 34679
rect 5295 34645 5333 34679
rect 5367 34645 5405 34679
rect 5439 34645 5477 34679
rect 5511 34645 5549 34679
rect 5583 34645 5621 34679
rect 5655 34645 5693 34679
rect 5727 34645 5765 34679
rect 5799 34645 5837 34679
rect 5871 34645 5909 34679
rect 5943 34645 5981 34679
rect 6015 34645 6053 34679
rect 6087 34645 6125 34679
rect 6159 34645 6197 34679
rect 6231 34645 6269 34679
rect 6303 34645 6341 34679
rect 6375 34645 6413 34679
rect 6447 34645 6485 34679
rect 6519 34645 6557 34679
rect 6591 34645 6629 34679
rect 6663 34645 6701 34679
rect 6735 34645 6773 34679
rect 6807 34645 6845 34679
rect 6879 34645 6917 34679
rect 6951 34645 6989 34679
rect 7023 34645 7061 34679
rect 7095 34645 7133 34679
rect 7167 34645 7205 34679
rect 7239 34645 7277 34679
rect 7311 34645 7349 34679
rect 7383 34645 7421 34679
rect 7455 34645 7493 34679
rect 7527 34645 7565 34679
rect 7599 34645 7637 34679
rect 7671 34645 7709 34679
rect 7743 34645 7781 34679
rect 7815 34645 7853 34679
rect 7887 34645 7925 34679
rect 7959 34645 7997 34679
rect 8031 34645 8069 34679
rect 8103 34645 8141 34679
rect 8175 34645 8213 34679
rect 8247 34645 8285 34679
rect 8319 34645 8357 34679
rect 8391 34645 8429 34679
rect 8463 34645 8501 34679
rect 8535 34645 8573 34679
rect 8607 34645 8645 34679
rect 8679 34645 8717 34679
rect 8751 34645 8789 34679
rect 8823 34645 8861 34679
rect 8895 34645 8933 34679
rect 8967 34645 9005 34679
rect 9039 34645 9077 34679
rect 9111 34645 9149 34679
rect 9183 34645 9221 34679
rect 9255 34645 9293 34679
rect 9327 34645 9365 34679
rect 9399 34645 9437 34679
rect 9471 34645 9509 34679
rect 9543 34645 9581 34679
rect 9615 34645 9653 34679
rect 9687 34645 9725 34679
rect 9759 34645 9797 34679
rect 9831 34645 9869 34679
rect 9903 34645 9941 34679
rect 9975 34645 10013 34679
rect 10047 34645 10085 34679
rect 10119 34645 10157 34679
rect 10191 34645 10229 34679
rect 10263 34645 10301 34679
rect 10335 34645 10373 34679
rect 10407 34645 10445 34679
rect 10479 34645 10517 34679
rect 10551 34645 10589 34679
rect 10623 34645 10661 34679
rect 10695 34645 10733 34679
rect 10767 34645 10805 34679
rect 10839 34645 10877 34679
rect 10911 34645 10949 34679
rect 10983 34645 11021 34679
rect 11055 34645 11093 34679
rect 11127 34645 11165 34679
rect 11199 34645 11237 34679
rect 11271 34645 11309 34679
rect 11343 34645 11381 34679
rect 11415 34645 11453 34679
rect 11487 34645 11525 34679
rect 11559 34645 11597 34679
rect 11631 34645 11669 34679
rect 11703 34645 11741 34679
rect 11775 34645 11813 34679
rect 11847 34645 11885 34679
rect 11919 34645 11957 34679
rect 11991 34645 12029 34679
rect 12063 34645 12101 34679
rect 12135 34645 12173 34679
rect 12207 34645 12245 34679
rect 12279 34645 12317 34679
rect 12351 34645 12389 34679
rect 12423 34645 12461 34679
rect 12495 34645 12533 34679
rect 12567 34645 12605 34679
rect 12639 34645 12677 34679
rect 12711 34645 12749 34679
rect 12783 34645 12821 34679
rect 12855 34645 12893 34679
rect 12927 34645 12965 34679
rect 12999 34645 13037 34679
rect 13071 34645 13109 34679
rect 13143 34645 13181 34679
rect 13215 34645 13253 34679
rect 13287 34645 13325 34679
rect 13359 34645 13397 34679
rect 13431 34645 13469 34679
rect 13503 34645 13541 34679
rect 13575 34645 13613 34679
rect 13647 34645 13685 34679
rect 13719 34645 13887 34679
rect 1119 34603 13887 34645
rect 1119 34466 1237 34603
rect 1119 34432 1161 34466
rect 1195 34432 1237 34466
rect 1119 34394 1237 34432
rect 1119 34360 1161 34394
rect 1195 34360 1237 34394
rect 1119 34322 1237 34360
rect 1119 34288 1161 34322
rect 1195 34288 1237 34322
rect 1119 34250 1237 34288
rect 1119 34216 1161 34250
rect 1195 34216 1237 34250
rect 1119 34178 1237 34216
rect 1119 34144 1161 34178
rect 1195 34144 1237 34178
rect 1119 34106 1237 34144
rect 1119 34072 1161 34106
rect 1195 34072 1237 34106
rect 1119 34034 1237 34072
rect 1119 34000 1161 34034
rect 1195 34000 1237 34034
rect 1119 33962 1237 34000
rect 1119 33928 1161 33962
rect 1195 33928 1237 33962
rect 1119 33890 1237 33928
rect 1119 33856 1161 33890
rect 1195 33856 1237 33890
rect 1119 33818 1237 33856
rect 1119 33784 1161 33818
rect 1195 33784 1237 33818
rect 1119 33746 1237 33784
rect 1119 33712 1161 33746
rect 1195 33712 1237 33746
rect 1119 33674 1237 33712
rect 1119 33640 1161 33674
rect 1195 33640 1237 33674
rect 1119 33602 1237 33640
rect 1119 33568 1161 33602
rect 1195 33568 1237 33602
rect 1119 33530 1237 33568
rect 1119 33496 1161 33530
rect 1195 33496 1237 33530
rect 1119 33458 1237 33496
rect 1119 33424 1161 33458
rect 1195 33424 1237 33458
rect 1119 33386 1237 33424
rect 1119 33352 1161 33386
rect 1195 33352 1237 33386
rect 1119 33314 1237 33352
rect 1119 33280 1161 33314
rect 1195 33280 1237 33314
rect 1119 33242 1237 33280
rect 1119 33208 1161 33242
rect 1195 33208 1237 33242
rect 1119 33170 1237 33208
rect 1119 33136 1161 33170
rect 1195 33136 1237 33170
rect 1119 33098 1237 33136
rect 1119 33064 1161 33098
rect 1195 33064 1237 33098
rect 1119 33026 1237 33064
rect 1119 32992 1161 33026
rect 1195 32992 1237 33026
rect 1119 32954 1237 32992
rect 1119 32920 1161 32954
rect 1195 32920 1237 32954
rect 1119 32882 1237 32920
rect 1119 32848 1161 32882
rect 1195 32848 1237 32882
rect 1119 32810 1237 32848
rect 1119 32776 1161 32810
rect 1195 32776 1237 32810
rect 1119 32738 1237 32776
rect 1119 32704 1161 32738
rect 1195 32704 1237 32738
rect 1119 32666 1237 32704
rect 1119 32632 1161 32666
rect 1195 32632 1237 32666
rect 1119 32594 1237 32632
rect 1119 32560 1161 32594
rect 1195 32560 1237 32594
rect 1119 32522 1237 32560
rect 1119 32488 1161 32522
rect 1195 32488 1237 32522
rect 1119 32450 1237 32488
rect 1119 32416 1161 32450
rect 1195 32416 1237 32450
rect 1119 32378 1237 32416
rect 1119 32344 1161 32378
rect 1195 32344 1237 32378
rect 1119 32306 1237 32344
rect 1119 32272 1161 32306
rect 1195 32272 1237 32306
rect 1119 32234 1237 32272
rect 1119 32200 1161 32234
rect 1195 32200 1237 32234
rect 1119 32162 1237 32200
rect 1119 32128 1161 32162
rect 1195 32128 1237 32162
rect 1119 32090 1237 32128
rect 1119 32056 1161 32090
rect 1195 32056 1237 32090
rect 1119 32018 1237 32056
rect 1119 31984 1161 32018
rect 1195 31984 1237 32018
rect 1119 31946 1237 31984
rect 1119 31912 1161 31946
rect 1195 31912 1237 31946
rect 1119 31874 1237 31912
rect 1119 31840 1161 31874
rect 1195 31840 1237 31874
rect 1119 31802 1237 31840
rect 1119 31768 1161 31802
rect 1195 31768 1237 31802
rect 1119 31730 1237 31768
rect 1119 31696 1161 31730
rect 1195 31696 1237 31730
rect 1119 31658 1237 31696
rect 1119 31624 1161 31658
rect 1195 31624 1237 31658
rect 1119 31586 1237 31624
rect 1119 31552 1161 31586
rect 1195 31552 1237 31586
rect 1119 31514 1237 31552
rect 1119 31480 1161 31514
rect 1195 31480 1237 31514
rect 1119 31442 1237 31480
rect 1119 31408 1161 31442
rect 1195 31408 1237 31442
rect 1119 31370 1237 31408
rect 1119 31336 1161 31370
rect 1195 31336 1237 31370
rect 1119 31298 1237 31336
rect 1119 31264 1161 31298
rect 1195 31264 1237 31298
rect 1119 31226 1237 31264
rect 1119 31192 1161 31226
rect 1195 31192 1237 31226
rect 1119 31154 1237 31192
rect 1119 31120 1161 31154
rect 1195 31120 1237 31154
rect 1119 31082 1237 31120
rect 1119 31048 1161 31082
rect 1195 31048 1237 31082
rect 1119 31010 1237 31048
rect 1119 30976 1161 31010
rect 1195 30976 1237 31010
rect 1119 30938 1237 30976
rect 1119 30904 1161 30938
rect 1195 30904 1237 30938
rect 1119 30866 1237 30904
rect 1119 30832 1161 30866
rect 1195 30832 1237 30866
rect 1119 30794 1237 30832
rect 1119 30760 1161 30794
rect 1195 30760 1237 30794
rect 1119 30722 1237 30760
rect 1119 30688 1161 30722
rect 1195 30688 1237 30722
rect 1119 30650 1237 30688
rect 1119 30616 1161 30650
rect 1195 30616 1237 30650
rect 1119 30578 1237 30616
rect 1119 30544 1161 30578
rect 1195 30544 1237 30578
rect 1119 30506 1237 30544
rect 1119 30472 1161 30506
rect 1195 30472 1237 30506
rect 1119 30434 1237 30472
rect 1119 30400 1161 30434
rect 1195 30400 1237 30434
rect 1119 30362 1237 30400
rect 1119 30328 1161 30362
rect 1195 30328 1237 30362
rect 1119 30290 1237 30328
rect 1119 30256 1161 30290
rect 1195 30281 1237 30290
rect 13769 34474 13887 34603
rect 13769 34440 13809 34474
rect 13843 34440 13887 34474
rect 13769 34402 13887 34440
rect 13769 34368 13809 34402
rect 13843 34368 13887 34402
rect 13769 34330 13887 34368
rect 13769 34296 13809 34330
rect 13843 34296 13887 34330
rect 13769 34258 13887 34296
rect 13769 34224 13809 34258
rect 13843 34224 13887 34258
rect 13769 34186 13887 34224
rect 13769 34152 13809 34186
rect 13843 34152 13887 34186
rect 13769 34114 13887 34152
rect 13769 34080 13809 34114
rect 13843 34080 13887 34114
rect 13769 34042 13887 34080
rect 13769 34008 13809 34042
rect 13843 34008 13887 34042
rect 13769 33970 13887 34008
rect 13769 33936 13809 33970
rect 13843 33936 13887 33970
rect 13769 33898 13887 33936
rect 13769 33864 13809 33898
rect 13843 33864 13887 33898
rect 13769 33826 13887 33864
rect 13769 33792 13809 33826
rect 13843 33792 13887 33826
rect 13769 33754 13887 33792
rect 13769 33720 13809 33754
rect 13843 33720 13887 33754
rect 13769 33682 13887 33720
rect 13769 33648 13809 33682
rect 13843 33648 13887 33682
rect 13769 33610 13887 33648
rect 13769 33576 13809 33610
rect 13843 33576 13887 33610
rect 13769 33538 13887 33576
rect 13769 33504 13809 33538
rect 13843 33504 13887 33538
rect 13769 33466 13887 33504
rect 13769 33432 13809 33466
rect 13843 33432 13887 33466
rect 13769 33394 13887 33432
rect 13769 33360 13809 33394
rect 13843 33360 13887 33394
rect 13769 33322 13887 33360
rect 13769 33288 13809 33322
rect 13843 33288 13887 33322
rect 13769 33250 13887 33288
rect 13769 33216 13809 33250
rect 13843 33216 13887 33250
rect 13769 33178 13887 33216
rect 13769 33144 13809 33178
rect 13843 33144 13887 33178
rect 13769 33106 13887 33144
rect 13769 33072 13809 33106
rect 13843 33072 13887 33106
rect 13769 33034 13887 33072
rect 13769 33000 13809 33034
rect 13843 33000 13887 33034
rect 13769 32962 13887 33000
rect 13769 32928 13809 32962
rect 13843 32928 13887 32962
rect 13769 32890 13887 32928
rect 13769 32856 13809 32890
rect 13843 32856 13887 32890
rect 13769 32818 13887 32856
rect 13769 32784 13809 32818
rect 13843 32784 13887 32818
rect 13769 32746 13887 32784
rect 13769 32712 13809 32746
rect 13843 32712 13887 32746
rect 13769 32674 13887 32712
rect 13769 32640 13809 32674
rect 13843 32640 13887 32674
rect 13769 32602 13887 32640
rect 13769 32568 13809 32602
rect 13843 32568 13887 32602
rect 13769 32530 13887 32568
rect 13769 32496 13809 32530
rect 13843 32496 13887 32530
rect 13769 32458 13887 32496
rect 13769 32424 13809 32458
rect 13843 32424 13887 32458
rect 13769 32386 13887 32424
rect 13769 32352 13809 32386
rect 13843 32352 13887 32386
rect 13769 32314 13887 32352
rect 13769 32280 13809 32314
rect 13843 32280 13887 32314
rect 13769 32242 13887 32280
rect 13769 32208 13809 32242
rect 13843 32208 13887 32242
rect 13769 32170 13887 32208
rect 13769 32136 13809 32170
rect 13843 32136 13887 32170
rect 13769 32098 13887 32136
rect 13769 32064 13809 32098
rect 13843 32064 13887 32098
rect 13769 32026 13887 32064
rect 13769 31992 13809 32026
rect 13843 31992 13887 32026
rect 13769 31954 13887 31992
rect 13769 31920 13809 31954
rect 13843 31920 13887 31954
rect 13769 31882 13887 31920
rect 13769 31848 13809 31882
rect 13843 31848 13887 31882
rect 13769 31810 13887 31848
rect 13769 31776 13809 31810
rect 13843 31776 13887 31810
rect 13769 31738 13887 31776
rect 13769 31704 13809 31738
rect 13843 31704 13887 31738
rect 13769 31666 13887 31704
rect 13769 31632 13809 31666
rect 13843 31632 13887 31666
rect 13769 31594 13887 31632
rect 13769 31560 13809 31594
rect 13843 31560 13887 31594
rect 13769 31522 13887 31560
rect 13769 31488 13809 31522
rect 13843 31488 13887 31522
rect 13769 31450 13887 31488
rect 13769 31416 13809 31450
rect 13843 31416 13887 31450
rect 13769 31378 13887 31416
rect 13769 31344 13809 31378
rect 13843 31344 13887 31378
rect 13769 31306 13887 31344
rect 13769 31272 13809 31306
rect 13843 31272 13887 31306
rect 13769 31234 13887 31272
rect 13769 31200 13809 31234
rect 13843 31200 13887 31234
rect 13769 31162 13887 31200
rect 13769 31128 13809 31162
rect 13843 31128 13887 31162
rect 13769 31090 13887 31128
rect 13769 31056 13809 31090
rect 13843 31056 13887 31090
rect 13769 31018 13887 31056
rect 13769 30984 13809 31018
rect 13843 30984 13887 31018
rect 13769 30946 13887 30984
rect 13769 30912 13809 30946
rect 13843 30912 13887 30946
rect 13769 30874 13887 30912
rect 13769 30840 13809 30874
rect 13843 30840 13887 30874
rect 13769 30802 13887 30840
rect 13769 30768 13809 30802
rect 13843 30768 13887 30802
rect 13769 30730 13887 30768
rect 13769 30696 13809 30730
rect 13843 30696 13887 30730
rect 13769 30658 13887 30696
rect 13769 30624 13809 30658
rect 13843 30624 13887 30658
rect 13769 30586 13887 30624
rect 13769 30552 13809 30586
rect 13843 30552 13887 30586
rect 13769 30514 13887 30552
rect 13769 30480 13809 30514
rect 13843 30480 13887 30514
rect 13769 30442 13887 30480
rect 13769 30408 13809 30442
rect 13843 30408 13887 30442
rect 13769 30370 13887 30408
rect 13769 30336 13809 30370
rect 13843 30336 13887 30370
rect 13769 30298 13887 30336
rect 1195 30264 10091 30281
tri 10091 30264 10108 30281 sw
rect 13769 30264 13809 30298
rect 13843 30264 13887 30298
rect 1195 30261 10108 30264
tri 10108 30261 10111 30264 sw
rect 1195 30256 10111 30261
rect 1119 30227 10111 30256
tri 10111 30227 10145 30261 sw
rect 1119 30218 4944 30227
rect 1119 30184 1161 30218
rect 1195 30184 4944 30218
rect 1119 30146 4944 30184
rect 1119 30112 1161 30146
rect 1195 30112 4944 30146
rect 1119 30074 4944 30112
rect 1119 30040 1161 30074
rect 1195 30040 4944 30074
rect 1119 30002 4944 30040
rect 1119 29968 1161 30002
rect 1195 29968 4944 30002
rect 1119 29930 4944 29968
rect 1119 29896 1161 29930
rect 1195 29896 4944 29930
rect 1119 29858 4944 29896
rect 1119 29824 1161 29858
rect 1195 29824 4944 29858
rect 1119 29786 4944 29824
rect 1119 29752 1161 29786
rect 1195 29752 4944 29786
rect 1119 29714 4944 29752
rect 1119 29680 1161 29714
rect 1195 29680 4944 29714
rect 1119 29642 4944 29680
rect 1119 29608 1161 29642
rect 1195 29608 4944 29642
rect 1119 29570 4944 29608
rect 1119 29536 1161 29570
rect 1195 29536 4944 29570
rect 1119 29498 4944 29536
rect 1119 29464 1161 29498
rect 1195 29464 4944 29498
rect 1119 29426 4944 29464
rect 1119 29392 1161 29426
rect 1195 29407 4944 29426
rect 7236 29407 7745 30227
rect 10037 30226 10145 30227
tri 10145 30226 10146 30227 sw
rect 13769 30226 13887 30264
rect 10037 30192 10146 30226
tri 10146 30192 10180 30226 sw
rect 13769 30192 13809 30226
rect 13843 30192 13887 30226
rect 10037 30189 10180 30192
tri 10180 30189 10183 30192 sw
rect 10037 30155 10183 30189
tri 10183 30155 10217 30189 sw
rect 10037 30154 10217 30155
tri 10217 30154 10218 30155 sw
rect 13769 30154 13887 30192
rect 10037 30120 10218 30154
tri 10218 30120 10252 30154 sw
rect 13769 30120 13809 30154
rect 13843 30120 13887 30154
rect 10037 30117 10252 30120
tri 10252 30117 10255 30120 sw
rect 10037 30083 10255 30117
tri 10255 30083 10289 30117 sw
rect 10037 30082 10289 30083
tri 10289 30082 10290 30083 sw
rect 13769 30082 13887 30120
rect 10037 30081 10290 30082
tri 10290 30081 10291 30082 sw
rect 10037 29553 10291 30081
rect 10037 29544 10282 29553
tri 10282 29544 10291 29553 nw
rect 13769 30048 13809 30082
rect 13843 30048 13887 30082
rect 13769 30010 13887 30048
rect 13769 29976 13809 30010
rect 13843 29976 13887 30010
rect 13769 29938 13887 29976
rect 13769 29904 13809 29938
rect 13843 29904 13887 29938
rect 13769 29866 13887 29904
rect 13769 29832 13809 29866
rect 13843 29832 13887 29866
rect 13769 29794 13887 29832
rect 13769 29760 13809 29794
rect 13843 29760 13887 29794
rect 13769 29722 13887 29760
rect 13769 29688 13809 29722
rect 13843 29688 13887 29722
rect 13769 29650 13887 29688
rect 13769 29616 13809 29650
rect 13843 29616 13887 29650
rect 13769 29578 13887 29616
rect 13769 29544 13809 29578
rect 13843 29544 13887 29578
rect 10037 29541 10279 29544
tri 10279 29541 10282 29544 nw
rect 10037 29507 10245 29541
tri 10245 29507 10279 29541 nw
rect 10037 29506 10244 29507
tri 10244 29506 10245 29507 nw
rect 13769 29506 13887 29544
rect 10037 29472 10210 29506
tri 10210 29472 10244 29506 nw
rect 13769 29472 13809 29506
rect 13843 29472 13887 29506
rect 10037 29469 10207 29472
tri 10207 29469 10210 29472 nw
rect 10037 29435 10173 29469
tri 10173 29435 10207 29469 nw
rect 10037 29434 10172 29435
tri 10172 29434 10173 29435 nw
rect 13769 29434 13887 29472
rect 10037 29407 10138 29434
rect 1195 29400 10138 29407
tri 10138 29400 10172 29434 nw
rect 13769 29400 13809 29434
rect 13843 29400 13887 29434
rect 1195 29397 10135 29400
tri 10135 29397 10138 29400 nw
rect 1195 29392 10101 29397
rect 1119 29363 10101 29392
tri 10101 29363 10135 29397 nw
rect 1119 29362 10100 29363
tri 10100 29362 10101 29363 nw
rect 13769 29362 13887 29400
rect 1119 29354 10091 29362
rect 1119 29320 1161 29354
rect 1195 29353 10091 29354
tri 10091 29353 10100 29362 nw
rect 1195 29320 1442 29353
rect 1119 29282 1442 29320
rect 1119 29248 1161 29282
rect 1195 29248 1442 29282
rect 1119 29210 1442 29248
rect 1119 29176 1161 29210
rect 1195 29176 1442 29210
rect 1119 29138 1442 29176
rect 1119 29104 1161 29138
rect 1195 29104 1442 29138
rect 1119 29066 1442 29104
rect 1119 29032 1161 29066
rect 1195 29032 1442 29066
rect 1119 28994 1442 29032
rect 1119 28960 1161 28994
rect 1195 28960 1442 28994
rect 1119 28922 1442 28960
rect 1119 28888 1161 28922
rect 1195 28888 1442 28922
rect 13769 29328 13809 29362
rect 13843 29328 13887 29362
rect 13769 29290 13887 29328
rect 13769 29256 13809 29290
rect 13843 29256 13887 29290
rect 13769 29218 13887 29256
rect 13769 29184 13809 29218
rect 13843 29184 13887 29218
rect 13769 29146 13887 29184
rect 13769 29112 13809 29146
rect 13843 29112 13887 29146
rect 13769 29074 13887 29112
rect 13769 29040 13809 29074
rect 13843 29040 13887 29074
rect 13769 29002 13887 29040
rect 13769 28968 13809 29002
rect 13843 28968 13887 29002
rect 13769 28930 13887 28968
tri 1846 28896 1859 28909 se
rect 1859 28896 13157 28909
tri 13157 28896 13170 28909 sw
rect 13769 28896 13809 28930
rect 13843 28896 13887 28930
tri 1843 28893 1846 28896 se
rect 1846 28893 13170 28896
tri 13170 28893 13173 28896 sw
rect 1119 28850 1442 28888
tri 1831 28881 1843 28893 se
rect 1843 28881 13173 28893
tri 1825 28875 1831 28881 se
rect 1831 28875 13173 28881
rect 1119 28816 1161 28850
rect 1195 28816 1442 28850
rect 1119 28778 1442 28816
rect 1119 28744 1161 28778
rect 1195 28744 1442 28778
rect 1119 28706 1442 28744
rect 1119 28672 1161 28706
rect 1195 28672 1442 28706
rect 1119 28634 1442 28672
rect 1119 28600 1161 28634
rect 1195 28600 1442 28634
rect 1119 28562 1442 28600
rect 1119 28528 1161 28562
rect 1195 28528 1442 28562
rect 1119 28490 1442 28528
rect 1119 28456 1161 28490
rect 1195 28456 1442 28490
rect 1119 28418 1442 28456
rect 1119 28384 1161 28418
rect 1195 28384 1442 28418
rect 1119 28346 1442 28384
rect 1119 28312 1161 28346
rect 1195 28312 1442 28346
rect 1119 28274 1442 28312
rect 1119 28240 1161 28274
rect 1195 28240 1442 28274
rect 1119 28202 1442 28240
rect 1119 28168 1161 28202
rect 1195 28168 1442 28202
rect 1119 28130 1442 28168
rect 1119 28096 1161 28130
rect 1195 28096 1442 28130
rect 1119 28058 1442 28096
rect 1119 28024 1161 28058
rect 1195 28024 1442 28058
rect 1119 27986 1442 28024
rect 1119 27952 1161 27986
rect 1195 27952 1442 27986
rect 1119 27914 1442 27952
rect 1119 27880 1161 27914
rect 1195 27880 1442 27914
rect 1119 27842 1442 27880
rect 1119 27808 1161 27842
rect 1195 27808 1442 27842
rect 1119 27770 1442 27808
rect 1119 27736 1161 27770
rect 1195 27736 1442 27770
rect 1119 27698 1442 27736
rect 1119 27664 1161 27698
rect 1195 27664 1442 27698
rect 1119 27626 1442 27664
rect 1119 27592 1161 27626
rect 1195 27592 1442 27626
rect 1119 27554 1442 27592
rect 1119 27520 1161 27554
rect 1195 27520 1442 27554
rect 1119 27482 1442 27520
rect 1119 27448 1161 27482
rect 1195 27448 1442 27482
rect 1119 27410 1442 27448
rect 1119 27376 1161 27410
rect 1195 27376 1442 27410
rect 1119 27338 1442 27376
rect 1119 27304 1161 27338
rect 1195 27304 1442 27338
rect 1119 27266 1442 27304
rect 1119 27232 1161 27266
rect 1195 27232 1442 27266
rect 1119 27194 1442 27232
rect 1119 27160 1161 27194
rect 1195 27160 1442 27194
rect 1119 27122 1442 27160
rect 1119 27088 1161 27122
rect 1195 27088 1442 27122
rect 1119 27050 1442 27088
tri 1659 28709 1825 28875 se
rect 1825 28709 1982 28875
rect 1659 28553 1982 28709
rect 13032 28859 13173 28875
tri 13173 28859 13207 28893 sw
rect 13032 28858 13207 28859
tri 13207 28858 13208 28859 sw
rect 13769 28858 13887 28896
rect 13032 28824 13208 28858
tri 13208 28824 13242 28858 sw
rect 13769 28824 13809 28858
rect 13843 28824 13887 28858
rect 13032 28821 13242 28824
tri 13242 28821 13245 28824 sw
rect 13032 28787 13245 28821
tri 13245 28787 13279 28821 sw
rect 13032 28786 13279 28787
tri 13279 28786 13280 28787 sw
rect 13769 28786 13887 28824
rect 13032 28752 13280 28786
tri 13280 28752 13314 28786 sw
rect 13769 28752 13809 28786
rect 13843 28752 13887 28786
rect 13032 28749 13314 28752
tri 13314 28749 13317 28752 sw
rect 13032 28744 13317 28749
tri 13317 28744 13322 28749 sw
rect 13032 28715 13322 28744
tri 13322 28715 13351 28744 sw
rect 13769 28727 13887 28752
rect 14099 34691 14122 34725
rect 14156 34691 14219 34725
rect 14099 34653 14219 34691
rect 14099 34619 14122 34653
rect 14156 34619 14219 34653
rect 14099 34581 14219 34619
rect 14099 34547 14122 34581
rect 14156 34547 14219 34581
rect 14099 34509 14219 34547
rect 14099 34475 14122 34509
rect 14156 34475 14219 34509
rect 14099 34437 14219 34475
rect 14099 34403 14122 34437
rect 14156 34403 14219 34437
rect 14099 34365 14219 34403
rect 14099 34331 14122 34365
rect 14156 34331 14219 34365
rect 14099 34293 14219 34331
rect 14099 34259 14122 34293
rect 14156 34259 14219 34293
rect 14099 34221 14219 34259
rect 14099 34187 14122 34221
rect 14156 34187 14219 34221
rect 14099 34149 14219 34187
rect 14099 34115 14122 34149
rect 14156 34115 14219 34149
rect 14099 34077 14219 34115
rect 14099 34043 14122 34077
rect 14156 34043 14219 34077
rect 14099 34005 14219 34043
rect 14099 33971 14122 34005
rect 14156 33971 14219 34005
rect 14099 33933 14219 33971
rect 14099 33899 14122 33933
rect 14156 33899 14219 33933
rect 14099 33861 14219 33899
rect 14099 33827 14122 33861
rect 14156 33827 14219 33861
rect 14099 33789 14219 33827
rect 14099 33755 14122 33789
rect 14156 33755 14219 33789
rect 14099 33717 14219 33755
rect 14099 33683 14122 33717
rect 14156 33683 14219 33717
rect 14099 33645 14219 33683
rect 14099 33611 14122 33645
rect 14156 33611 14219 33645
rect 14099 33573 14219 33611
rect 14099 33539 14122 33573
rect 14156 33539 14219 33573
rect 14099 33501 14219 33539
rect 14099 33467 14122 33501
rect 14156 33467 14219 33501
rect 14099 33429 14219 33467
rect 14099 33395 14122 33429
rect 14156 33395 14219 33429
rect 14099 33357 14219 33395
rect 14099 33323 14122 33357
rect 14156 33323 14219 33357
rect 14099 33285 14219 33323
rect 14099 33251 14122 33285
rect 14156 33251 14219 33285
rect 14099 33213 14219 33251
rect 14099 33179 14122 33213
rect 14156 33179 14219 33213
rect 14099 33141 14219 33179
rect 14099 33107 14122 33141
rect 14156 33107 14219 33141
rect 14099 33069 14219 33107
rect 14099 33035 14122 33069
rect 14156 33035 14219 33069
rect 14099 32997 14219 33035
rect 14099 32963 14122 32997
rect 14156 32963 14219 32997
rect 14099 32925 14219 32963
rect 14099 32891 14122 32925
rect 14156 32891 14219 32925
rect 14099 32853 14219 32891
rect 14099 32819 14122 32853
rect 14156 32819 14219 32853
rect 14099 32781 14219 32819
rect 14099 32747 14122 32781
rect 14156 32747 14219 32781
rect 14099 32709 14219 32747
rect 14099 32675 14122 32709
rect 14156 32675 14219 32709
rect 14099 32637 14219 32675
rect 14099 32603 14122 32637
rect 14156 32603 14219 32637
rect 14099 32565 14219 32603
rect 14099 32531 14122 32565
rect 14156 32531 14219 32565
rect 14099 32493 14219 32531
rect 14099 32459 14122 32493
rect 14156 32459 14219 32493
rect 14099 32421 14219 32459
rect 14099 32387 14122 32421
rect 14156 32387 14219 32421
rect 14099 32349 14219 32387
rect 14099 32315 14122 32349
rect 14156 32315 14219 32349
rect 14099 32277 14219 32315
rect 14099 32243 14122 32277
rect 14156 32243 14219 32277
rect 14099 32205 14219 32243
rect 14099 32171 14122 32205
rect 14156 32171 14219 32205
rect 14099 32133 14219 32171
rect 14099 32099 14122 32133
rect 14156 32099 14219 32133
rect 14099 32061 14219 32099
rect 14099 32027 14122 32061
rect 14156 32027 14219 32061
rect 14099 31989 14219 32027
rect 14099 31955 14122 31989
rect 14156 31955 14219 31989
rect 14099 31917 14219 31955
rect 14099 31883 14122 31917
rect 14156 31883 14219 31917
rect 14099 31845 14219 31883
rect 14099 31811 14122 31845
rect 14156 31811 14219 31845
rect 14099 31773 14219 31811
rect 14099 31739 14122 31773
rect 14156 31739 14219 31773
rect 14099 31701 14219 31739
rect 14099 31667 14122 31701
rect 14156 31667 14219 31701
rect 14099 31629 14219 31667
rect 14099 31595 14122 31629
rect 14156 31595 14219 31629
rect 14099 31557 14219 31595
rect 14099 31523 14122 31557
rect 14156 31523 14219 31557
rect 14099 31485 14219 31523
rect 14099 31451 14122 31485
rect 14156 31451 14219 31485
rect 14099 31413 14219 31451
rect 14099 31379 14122 31413
rect 14156 31379 14219 31413
rect 14099 31341 14219 31379
rect 14099 31307 14122 31341
rect 14156 31307 14219 31341
rect 14099 31269 14219 31307
rect 14099 31235 14122 31269
rect 14156 31235 14219 31269
rect 14099 31197 14219 31235
rect 14099 31163 14122 31197
rect 14156 31163 14219 31197
rect 14099 31125 14219 31163
rect 14099 31091 14122 31125
rect 14156 31091 14219 31125
rect 14099 31053 14219 31091
rect 14099 31019 14122 31053
rect 14156 31019 14219 31053
rect 14099 30981 14219 31019
rect 14099 30947 14122 30981
rect 14156 30947 14219 30981
rect 14099 30909 14219 30947
rect 14099 30875 14122 30909
rect 14156 30875 14219 30909
rect 14099 30837 14219 30875
rect 14099 30803 14122 30837
rect 14156 30803 14219 30837
rect 14099 30765 14219 30803
rect 14099 30731 14122 30765
rect 14156 30731 14219 30765
rect 14099 30693 14219 30731
rect 14099 30659 14122 30693
rect 14156 30659 14219 30693
rect 14099 30621 14219 30659
rect 14099 30587 14122 30621
rect 14156 30587 14219 30621
rect 14099 30549 14219 30587
rect 14099 30515 14122 30549
rect 14156 30515 14219 30549
rect 14099 30477 14219 30515
rect 14099 30443 14122 30477
rect 14156 30443 14219 30477
rect 14099 30405 14219 30443
rect 14099 30371 14122 30405
rect 14156 30371 14219 30405
rect 14099 30333 14219 30371
rect 14099 30299 14122 30333
rect 14156 30299 14219 30333
rect 14099 30261 14219 30299
rect 14099 30227 14122 30261
rect 14156 30227 14219 30261
rect 14099 30189 14219 30227
rect 14099 30155 14122 30189
rect 14156 30155 14219 30189
rect 14099 30117 14219 30155
rect 14099 30083 14122 30117
rect 14156 30083 14219 30117
rect 14099 30045 14219 30083
rect 14099 30011 14122 30045
rect 14156 30011 14219 30045
rect 14099 29973 14219 30011
rect 14099 29939 14122 29973
rect 14156 29939 14219 29973
rect 14099 29901 14219 29939
rect 14099 29867 14122 29901
rect 14156 29867 14219 29901
rect 14099 29829 14219 29867
rect 14099 29795 14122 29829
rect 14156 29795 14219 29829
rect 14099 29757 14219 29795
rect 14099 29723 14122 29757
rect 14156 29723 14219 29757
rect 14099 29685 14219 29723
rect 14099 29651 14122 29685
rect 14156 29651 14219 29685
rect 14099 29613 14219 29651
rect 14099 29579 14122 29613
rect 14156 29579 14219 29613
rect 14099 29541 14219 29579
rect 14099 29507 14122 29541
rect 14156 29507 14219 29541
rect 14099 29469 14219 29507
rect 14099 29435 14122 29469
rect 14156 29435 14219 29469
rect 14099 29397 14219 29435
rect 14099 29363 14122 29397
rect 14156 29363 14219 29397
rect 14099 29325 14219 29363
rect 14099 29291 14122 29325
rect 14156 29291 14219 29325
rect 14099 29253 14219 29291
rect 14099 29219 14122 29253
rect 14156 29219 14219 29253
rect 14099 29181 14219 29219
rect 14099 29147 14122 29181
rect 14156 29147 14219 29181
rect 14099 29109 14219 29147
rect 14099 29075 14122 29109
rect 14156 29075 14219 29109
rect 14099 29037 14219 29075
rect 14099 29003 14122 29037
rect 14156 29003 14219 29037
rect 14099 28965 14219 29003
rect 14099 28931 14122 28965
rect 14156 28931 14219 28965
rect 14099 28893 14219 28931
rect 14099 28859 14122 28893
rect 14156 28859 14219 28893
rect 14099 28821 14219 28859
rect 14099 28787 14122 28821
rect 14156 28787 14219 28821
rect 14099 28749 14219 28787
rect 14099 28715 14122 28749
rect 14156 28715 14219 28749
rect 13032 28702 13351 28715
tri 13351 28702 13364 28715 sw
rect 13032 28677 13364 28702
tri 13364 28677 13389 28702 sw
rect 14099 28677 14219 28715
rect 13032 28643 13389 28677
tri 13389 28643 13423 28677 sw
rect 14099 28643 14122 28677
rect 14156 28643 14219 28677
rect 13032 28630 13423 28643
tri 13423 28630 13436 28643 sw
rect 13032 28605 13436 28630
tri 13436 28605 13461 28630 sw
rect 14099 28605 14219 28643
rect 13032 28590 13461 28605
tri 13461 28590 13476 28605 sw
rect 13032 28571 13476 28590
tri 13476 28571 13495 28590 sw
rect 14099 28571 14122 28605
rect 14156 28571 14219 28605
rect 13032 28558 13495 28571
tri 13495 28558 13508 28571 sw
rect 13032 28553 13508 28558
rect 1659 28533 13508 28553
tri 13508 28533 13533 28558 sw
rect 14099 28533 14219 28571
rect 1659 28515 13533 28533
rect 1659 28499 2117 28515
tri 2117 28499 2133 28515 nw
tri 12883 28499 12899 28515 ne
rect 12899 28499 13533 28515
tri 13533 28499 13567 28533 sw
rect 14099 28499 14122 28533
rect 14156 28499 14219 28533
rect 1659 28489 2104 28499
rect 1659 27447 1726 28489
rect 1976 28486 2104 28489
tri 2104 28486 2117 28499 nw
tri 12899 28486 12912 28499 ne
rect 12912 28486 13567 28499
tri 13567 28486 13580 28499 sw
rect 1976 28485 2103 28486
tri 2103 28485 2104 28486 nw
tri 12912 28485 12913 28486 ne
rect 12913 28485 13580 28486
rect 1976 28482 2100 28485
tri 2100 28482 2103 28485 nw
tri 12913 28482 12916 28485 ne
rect 12916 28482 13580 28485
rect 1976 27447 2093 28482
tri 2093 28475 2100 28482 nw
tri 12916 28475 12923 28482 ne
tri 2320 28276 2412 28368 se
rect 2412 28335 12604 28368
rect 2412 28276 4939 28335
rect 2319 28219 4939 28276
rect 7231 28219 7750 28335
rect 10042 28276 12604 28335
tri 12604 28276 12696 28368 sw
rect 10042 28219 12696 28276
rect 2319 28168 12696 28219
rect 2509 28022 4482 28048
rect 4481 27906 4482 28022
rect 2509 27880 4482 27906
rect 10500 28022 12473 28048
rect 12472 27906 12473 28022
rect 10500 27880 12473 27906
rect 2320 27719 12696 27764
rect 2320 27652 4939 27719
tri 2320 27552 2420 27652 ne
rect 2420 27603 4939 27652
rect 7231 27603 7750 27719
rect 10042 27652 12696 27719
rect 10042 27603 12596 27652
rect 2420 27552 12596 27603
tri 12596 27552 12696 27652 nw
rect 1659 27440 2093 27447
tri 2093 27440 2104 27451 sw
tri 12912 27440 12923 27451 se
rect 12923 27440 13031 28482
rect 13281 28461 13580 28482
tri 13580 28461 13605 28486 sw
rect 14099 28461 14219 28499
rect 13281 28427 13605 28461
tri 13605 28427 13639 28461 sw
rect 14099 28427 14122 28461
rect 14156 28427 14219 28461
rect 13281 28414 13639 28427
tri 13639 28414 13652 28427 sw
rect 13281 28389 13652 28414
tri 13652 28389 13677 28414 sw
rect 14099 28389 14219 28427
rect 13281 28355 13677 28389
tri 13677 28355 13711 28389 sw
rect 14099 28355 14122 28389
rect 14156 28355 14219 28389
rect 13281 28342 13711 28355
tri 13711 28342 13724 28355 sw
rect 13281 28317 13724 28342
tri 13724 28317 13749 28342 sw
rect 14099 28317 14219 28355
rect 13281 28283 13749 28317
tri 13749 28283 13783 28317 sw
rect 13281 27440 13783 28283
rect 1659 27437 2104 27440
tri 2104 27437 2107 27440 sw
tri 12909 27437 12912 27440 se
rect 12912 27437 13783 27440
rect 1659 27419 2107 27437
tri 2107 27419 2125 27437 sw
tri 12891 27419 12909 27437 se
rect 12909 27419 13783 27437
rect 1659 27411 2125 27419
tri 2125 27411 2133 27419 sw
tri 12883 27411 12891 27419 se
rect 12891 27411 13783 27419
rect 1659 27334 13783 27411
rect 1659 27217 1985 27334
tri 1659 27084 1792 27217 ne
rect 1792 27084 1985 27217
rect 13035 27217 13783 27334
rect 13035 27203 13343 27217
tri 13343 27203 13357 27217 nw
rect 13035 27190 13330 27203
tri 13330 27190 13343 27203 nw
rect 13035 27165 13305 27190
tri 13305 27165 13330 27190 nw
rect 13035 27131 13271 27165
tri 13271 27131 13305 27165 nw
rect 13035 27118 13258 27131
tri 13258 27118 13271 27131 nw
rect 13035 27093 13233 27118
tri 13233 27093 13258 27118 nw
rect 13035 27084 13199 27093
tri 1792 27059 1817 27084 ne
rect 1817 27059 13199 27084
tri 13199 27059 13233 27093 nw
tri 1817 27053 1823 27059 ne
rect 1823 27053 13186 27059
rect 1119 27016 1161 27050
rect 1195 27016 1442 27050
tri 1823 27046 1830 27053 ne
rect 1830 27046 13186 27053
tri 13186 27046 13199 27059 nw
tri 1830 27021 1855 27046 ne
rect 1855 27021 13161 27046
tri 13161 27021 13186 27046 nw
tri 1855 27017 1859 27021 ne
rect 1859 27017 13157 27021
tri 13157 27017 13161 27021 nw
rect 1119 26978 1442 27016
rect 1119 26944 1161 26978
rect 1195 26944 1442 26978
rect 1119 26906 1442 26944
rect 1119 26872 1161 26906
rect 1195 26872 1442 26906
rect 1119 26834 1442 26872
rect 1119 26800 1161 26834
rect 1195 26800 1442 26834
rect 1119 26762 1442 26800
rect 1119 26728 1161 26762
rect 1195 26728 1442 26762
rect 1119 26690 1442 26728
rect 1119 26656 1161 26690
rect 1195 26656 1442 26690
rect 1119 26618 1442 26656
rect 1119 26584 1161 26618
rect 1195 26584 1442 26618
rect 1119 26546 1442 26584
rect 1119 26512 1161 26546
rect 1195 26512 1442 26546
rect 1119 26474 1442 26512
rect 1119 26440 1161 26474
rect 1195 26440 1442 26474
rect 1119 26402 1442 26440
rect 1119 26368 1161 26402
rect 1195 26368 1442 26402
rect 1119 26330 1442 26368
rect 1119 26296 1161 26330
rect 1195 26296 1442 26330
rect 1119 26258 1442 26296
rect 1119 26224 1161 26258
rect 1195 26224 1442 26258
rect 1119 26192 1442 26224
rect 1119 26186 1736 26192
rect 1119 26152 1161 26186
rect 1195 26152 1736 26186
rect 1119 26114 1736 26152
rect 1119 26080 1161 26114
rect 1195 26080 1736 26114
rect 1119 26042 1736 26080
tri 2413 26051 2414 26052 se
rect 2414 26051 12578 26052
tri 12578 26051 12579 26052 sw
rect 1119 26008 1161 26042
rect 1195 26008 1736 26042
tri 2400 26038 2413 26051 se
rect 2413 26038 12579 26051
tri 12579 26038 12592 26051 sw
tri 2375 26013 2400 26038 se
rect 2400 26025 12592 26038
rect 2400 26013 4933 26025
rect 1119 25970 1736 26008
tri 2341 25979 2375 26013 se
rect 2375 25979 4933 26013
rect 1119 25936 1161 25970
rect 1195 25936 1736 25970
rect 1119 25898 1736 25936
rect 1119 25864 1161 25898
rect 1195 25864 1736 25898
tri 2328 25966 2341 25979 se
rect 2341 25966 4933 25979
rect 2328 25909 4933 25966
rect 7225 25909 7757 26025
rect 10049 26013 12592 26025
tri 12592 26013 12617 26038 sw
rect 10049 25979 12617 26013
tri 12617 25979 12651 26013 sw
rect 10049 25966 12651 25979
tri 12651 25966 12664 25979 sw
rect 10049 25909 12664 25966
rect 2328 25880 12664 25909
rect 1119 25826 1736 25864
rect 1119 25792 1161 25826
rect 1195 25792 1736 25826
rect 1119 25754 1736 25792
rect 1119 25720 1161 25754
rect 1195 25720 1736 25754
rect 1119 25682 1736 25720
rect 1119 25648 1161 25682
rect 1195 25648 1736 25682
rect 1119 25610 1736 25648
rect 2528 25759 4472 25781
rect 2528 25643 2546 25759
rect 4454 25643 4472 25759
rect 2528 25621 4472 25643
rect 10510 25759 12454 25781
rect 10510 25643 10528 25759
rect 12436 25643 12454 25759
rect 10510 25621 12454 25643
rect 1119 25576 1161 25610
rect 1195 25576 1736 25610
rect 1119 25538 1736 25576
rect 1119 25504 1161 25538
rect 1195 25504 1736 25538
rect 1119 25466 1736 25504
rect 1119 25432 1161 25466
rect 1195 25432 1736 25466
rect 1119 25394 1736 25432
rect 2326 25493 12662 25520
rect 2326 25428 4933 25493
tri 2326 25403 2351 25428 ne
rect 2351 25403 4933 25428
rect 1119 25360 1161 25394
rect 1195 25360 1736 25394
tri 2351 25390 2364 25403 ne
rect 2364 25390 4933 25403
tri 2364 25365 2389 25390 ne
rect 2389 25377 4933 25390
rect 7225 25377 7757 25493
rect 10049 25428 12662 25493
rect 10049 25403 12637 25428
tri 12637 25403 12662 25428 nw
rect 10049 25390 12624 25403
tri 12624 25390 12637 25403 nw
rect 10049 25377 12599 25390
rect 2389 25365 12599 25377
tri 12599 25365 12624 25390 nw
rect 1119 25322 1736 25360
tri 2389 25348 2406 25365 ne
rect 2406 25348 12582 25365
tri 12582 25348 12599 25365 nw
rect 1119 25288 1161 25322
rect 1195 25288 1736 25322
rect 1119 25250 1736 25288
rect 1119 25216 1161 25250
rect 1195 25216 1736 25250
rect 1119 25202 1736 25216
rect 1119 25178 1237 25202
rect 1119 25144 1161 25178
rect 1195 25144 1237 25178
rect 1119 25106 1237 25144
rect 1119 25072 1161 25106
rect 1195 25072 1237 25106
rect 1119 25034 1237 25072
rect 1119 25000 1161 25034
rect 1195 25000 1237 25034
rect 1119 24962 1237 25000
rect 1119 24928 1161 24962
rect 1195 24928 1237 24962
rect 1119 24890 1237 24928
rect 1119 24856 1161 24890
rect 1195 24856 1237 24890
rect 1119 24818 1237 24856
rect 1119 24784 1161 24818
rect 1195 24784 1237 24818
rect 1119 24746 1237 24784
rect 1119 24712 1161 24746
rect 1195 24712 1237 24746
rect 1119 24674 1237 24712
rect 1119 24640 1161 24674
rect 1195 24640 1237 24674
rect 1119 24602 1237 24640
rect 1119 24568 1161 24602
rect 1195 24568 1237 24602
rect 1119 24530 1237 24568
rect 13527 24543 13783 27217
tri 4887 24539 4891 24543 se
rect 4891 24539 13783 24543
rect 1119 24496 1161 24530
rect 1195 24496 1237 24530
tri 4874 24526 4887 24539 se
rect 4887 24526 13783 24539
tri 4849 24501 4874 24526 se
rect 4874 24501 13783 24526
rect 1119 24458 1237 24496
tri 4815 24467 4849 24501 se
rect 4849 24489 13783 24501
rect 4849 24467 4945 24489
rect 1119 24424 1161 24458
rect 1195 24424 1237 24458
tri 4802 24454 4815 24467 se
rect 4815 24454 4945 24467
tri 4777 24429 4802 24454 se
rect 4802 24429 4945 24454
rect 1119 24386 1237 24424
tri 4743 24395 4777 24429 se
rect 4777 24395 4945 24429
rect 1119 24352 1161 24386
rect 1195 24352 1237 24386
tri 4730 24382 4743 24395 se
rect 4743 24382 4945 24395
tri 4705 24357 4730 24382 se
rect 4730 24357 4945 24382
rect 1119 24314 1237 24352
rect 1119 24280 1161 24314
rect 1195 24280 1237 24314
rect 1119 24242 1237 24280
rect 1119 24208 1161 24242
rect 1195 24208 1237 24242
rect 1119 24170 1237 24208
rect 1119 24136 1161 24170
rect 1195 24136 1237 24170
rect 1119 24098 1237 24136
rect 1119 24064 1161 24098
rect 1195 24064 1237 24098
rect 1119 24026 1237 24064
rect 1119 23992 1161 24026
rect 1195 23992 1237 24026
rect 1119 23954 1237 23992
rect 1119 23920 1161 23954
rect 1195 23920 1237 23954
rect 1119 23882 1237 23920
rect 1119 23848 1161 23882
rect 1195 23848 1237 23882
rect 1119 23810 1237 23848
rect 1119 23776 1161 23810
rect 1195 23776 1237 23810
tri 4691 24343 4705 24357 se
rect 4705 24343 4945 24357
rect 4691 23815 4945 24343
tri 4691 23806 4700 23815 ne
rect 4700 23806 4945 23815
tri 4700 23781 4725 23806 ne
rect 4725 23781 4945 23806
rect 1119 23738 1237 23776
tri 4725 23747 4759 23781 ne
rect 4759 23747 4945 23781
rect 1119 23704 1161 23738
rect 1195 23704 1237 23738
tri 4759 23734 4772 23747 ne
rect 4772 23734 4945 23747
tri 4772 23709 4797 23734 ne
rect 4797 23709 4945 23734
rect 1119 23666 1237 23704
tri 4797 23675 4831 23709 ne
rect 4831 23675 4945 23709
rect 1119 23632 1161 23666
rect 1195 23632 1237 23666
tri 4831 23662 4844 23675 ne
rect 4844 23669 4945 23675
rect 7237 23669 7744 24489
rect 10036 24041 13783 24489
rect 10036 24035 13777 24041
tri 13777 24035 13783 24041 nw
rect 14099 28283 14122 28317
rect 14156 28283 14219 28317
rect 14099 28245 14219 28283
rect 14099 28211 14122 28245
rect 14156 28211 14219 28245
rect 14099 28173 14219 28211
rect 14099 28139 14122 28173
rect 14156 28139 14219 28173
rect 14099 28101 14219 28139
rect 14099 28067 14122 28101
rect 14156 28067 14219 28101
rect 14099 28029 14219 28067
rect 14099 27995 14122 28029
rect 14156 27995 14219 28029
rect 14099 27957 14219 27995
rect 14099 27923 14122 27957
rect 14156 27923 14219 27957
rect 14099 27885 14219 27923
rect 14099 27851 14122 27885
rect 14156 27851 14219 27885
rect 14099 27813 14219 27851
rect 14099 27779 14122 27813
rect 14156 27779 14219 27813
rect 14099 27741 14219 27779
rect 14099 27707 14122 27741
rect 14156 27707 14219 27741
rect 14099 27669 14219 27707
rect 14099 27635 14122 27669
rect 14156 27635 14219 27669
rect 14099 27597 14219 27635
rect 14099 27563 14122 27597
rect 14156 27563 14219 27597
rect 14099 27525 14219 27563
rect 14099 27491 14122 27525
rect 14156 27491 14219 27525
rect 14099 27453 14219 27491
rect 14099 27419 14122 27453
rect 14156 27419 14219 27453
rect 14099 27381 14219 27419
rect 14099 27347 14122 27381
rect 14156 27347 14219 27381
rect 14099 27309 14219 27347
rect 14099 27275 14122 27309
rect 14156 27275 14219 27309
rect 14099 27237 14219 27275
rect 14099 27203 14122 27237
rect 14156 27203 14219 27237
rect 14099 27165 14219 27203
rect 14099 27131 14122 27165
rect 14156 27131 14219 27165
rect 14099 27093 14219 27131
rect 14099 27059 14122 27093
rect 14156 27059 14219 27093
rect 14099 27021 14219 27059
rect 14099 26987 14122 27021
rect 14156 26987 14219 27021
rect 14099 26949 14219 26987
rect 14099 26915 14122 26949
rect 14156 26915 14219 26949
rect 14099 26877 14219 26915
rect 14099 26843 14122 26877
rect 14156 26843 14219 26877
rect 14099 26805 14219 26843
rect 14099 26771 14122 26805
rect 14156 26771 14219 26805
rect 14099 26733 14219 26771
rect 14099 26699 14122 26733
rect 14156 26699 14219 26733
rect 14099 26661 14219 26699
rect 14099 26627 14122 26661
rect 14156 26627 14219 26661
rect 14099 26589 14219 26627
rect 14099 26555 14122 26589
rect 14156 26555 14219 26589
rect 14099 26517 14219 26555
rect 14099 26483 14122 26517
rect 14156 26483 14219 26517
rect 14099 26445 14219 26483
rect 14099 26411 14122 26445
rect 14156 26411 14219 26445
rect 14099 26373 14219 26411
rect 14099 26339 14122 26373
rect 14156 26339 14219 26373
rect 14099 26301 14219 26339
rect 14099 26267 14122 26301
rect 14156 26267 14219 26301
rect 14099 26229 14219 26267
rect 14099 26195 14122 26229
rect 14156 26195 14219 26229
rect 14099 26157 14219 26195
rect 14099 26123 14122 26157
rect 14156 26123 14219 26157
rect 14099 26085 14219 26123
rect 14099 26051 14122 26085
rect 14156 26051 14219 26085
rect 14099 26013 14219 26051
rect 14099 25979 14122 26013
rect 14156 25979 14219 26013
rect 14099 25941 14219 25979
rect 14099 25907 14122 25941
rect 14156 25907 14219 25941
rect 14099 25869 14219 25907
rect 14099 25835 14122 25869
rect 14156 25835 14219 25869
rect 14099 25797 14219 25835
rect 14099 25763 14122 25797
rect 14156 25763 14219 25797
rect 14099 25725 14219 25763
rect 14099 25691 14122 25725
rect 14156 25691 14219 25725
rect 14099 25653 14219 25691
rect 14099 25619 14122 25653
rect 14156 25619 14219 25653
rect 14099 25581 14219 25619
rect 14099 25547 14122 25581
rect 14156 25547 14219 25581
rect 14099 25509 14219 25547
rect 14099 25475 14122 25509
rect 14156 25475 14219 25509
rect 14099 25437 14219 25475
rect 14099 25403 14122 25437
rect 14156 25403 14219 25437
rect 14099 25365 14219 25403
rect 14099 25331 14122 25365
rect 14156 25331 14219 25365
rect 14099 25293 14219 25331
rect 14099 25259 14122 25293
rect 14156 25259 14219 25293
rect 14099 25221 14219 25259
rect 14099 25187 14122 25221
rect 14156 25187 14219 25221
rect 14099 25149 14219 25187
rect 14099 25115 14122 25149
rect 14156 25115 14219 25149
rect 14099 25077 14219 25115
rect 14099 25043 14122 25077
rect 14156 25043 14219 25077
rect 14099 25005 14219 25043
rect 14099 24971 14122 25005
rect 14156 24971 14219 25005
rect 14099 24933 14219 24971
rect 14099 24899 14122 24933
rect 14156 24899 14219 24933
rect 14099 24861 14219 24899
rect 14099 24827 14122 24861
rect 14156 24827 14219 24861
rect 14099 24789 14219 24827
rect 14099 24755 14122 24789
rect 14156 24755 14219 24789
rect 14099 24717 14219 24755
rect 14099 24683 14122 24717
rect 14156 24683 14219 24717
rect 14099 24645 14219 24683
rect 14099 24611 14122 24645
rect 14156 24611 14219 24645
rect 14099 24573 14219 24611
rect 14099 24539 14122 24573
rect 14156 24539 14219 24573
rect 14099 24501 14219 24539
rect 14099 24467 14122 24501
rect 14156 24467 14219 24501
rect 14099 24429 14219 24467
rect 14099 24395 14122 24429
rect 14156 24395 14219 24429
rect 14099 24357 14219 24395
rect 14099 24323 14122 24357
rect 14156 24323 14219 24357
rect 14099 24285 14219 24323
rect 14099 24251 14122 24285
rect 14156 24251 14219 24285
rect 14099 24213 14219 24251
rect 14099 24179 14122 24213
rect 14156 24179 14219 24213
rect 14099 24141 14219 24179
rect 14099 24107 14122 24141
rect 14156 24107 14219 24141
rect 14099 24069 14219 24107
rect 14099 24035 14122 24069
rect 14156 24035 14219 24069
rect 10036 24022 13764 24035
tri 13764 24022 13777 24035 nw
rect 10036 23997 13739 24022
tri 13739 23997 13764 24022 nw
rect 14099 23997 14219 24035
rect 10036 23963 13705 23997
tri 13705 23963 13739 23997 nw
rect 14099 23963 14122 23997
rect 14156 23963 14219 23997
rect 10036 23950 13692 23963
tri 13692 23950 13705 23963 nw
rect 10036 23925 13667 23950
tri 13667 23925 13692 23950 nw
rect 14099 23925 14219 23963
rect 10036 23891 13633 23925
tri 13633 23891 13667 23925 nw
rect 14099 23891 14122 23925
rect 14156 23891 14219 23925
rect 10036 23878 13620 23891
tri 13620 23878 13633 23891 nw
rect 10036 23853 13595 23878
tri 13595 23853 13620 23878 nw
rect 14099 23853 14219 23891
rect 10036 23819 13561 23853
tri 13561 23819 13595 23853 nw
rect 14099 23819 14122 23853
rect 14156 23819 14219 23853
rect 10036 23806 13548 23819
tri 13548 23806 13561 23819 nw
rect 10036 23781 13523 23806
tri 13523 23781 13548 23806 nw
rect 14099 23781 14219 23819
rect 10036 23747 13489 23781
tri 13489 23747 13523 23781 nw
rect 14099 23747 14122 23781
rect 14156 23747 14219 23781
rect 10036 23734 13476 23747
tri 13476 23734 13489 23747 nw
rect 10036 23709 13451 23734
tri 13451 23709 13476 23734 nw
rect 14099 23709 14219 23747
rect 10036 23675 13417 23709
tri 13417 23675 13451 23709 nw
rect 14099 23675 14122 23709
rect 14156 23675 14219 23709
rect 10036 23669 13404 23675
rect 4844 23662 13404 23669
tri 13404 23662 13417 23675 nw
tri 4844 23637 4869 23662 ne
rect 4869 23637 13379 23662
tri 13379 23637 13404 23662 nw
rect 14099 23637 14219 23675
rect 1119 23594 1237 23632
tri 4869 23615 4891 23637 ne
rect 4891 23615 13357 23637
tri 13357 23615 13379 23637 nw
rect 1119 23560 1161 23594
rect 1195 23560 1237 23594
rect 1119 23522 1237 23560
rect 1119 23488 1161 23522
rect 1195 23488 1237 23522
rect 1119 23450 1237 23488
rect 1119 23416 1161 23450
rect 1195 23416 1237 23450
rect 14099 23603 14122 23637
rect 14156 23603 14219 23637
rect 14099 23565 14219 23603
rect 14099 23531 14122 23565
rect 14156 23531 14219 23565
rect 14099 23493 14219 23531
rect 14099 23459 14122 23493
rect 14156 23459 14219 23493
rect 1119 23378 1237 23416
rect 1119 23344 1161 23378
rect 1195 23344 1237 23378
rect 1119 23306 1237 23344
rect 1119 23272 1161 23306
rect 1195 23272 1237 23306
rect 1119 23234 1237 23272
rect 1119 23200 1161 23234
rect 1195 23200 1237 23234
rect 1119 23162 1237 23200
rect 1119 23128 1161 23162
rect 1195 23128 1237 23162
rect 1119 23090 1237 23128
rect 1119 23056 1161 23090
rect 1195 23056 1237 23090
rect 1119 23018 1237 23056
rect 1119 22984 1161 23018
rect 1195 22984 1237 23018
rect 1119 22946 1237 22984
rect 1119 22912 1161 22946
rect 1195 22912 1237 22946
rect 1119 22874 1237 22912
rect 1119 22840 1161 22874
rect 1195 22840 1237 22874
rect 1119 22802 1237 22840
rect 1119 22768 1161 22802
rect 1195 22768 1237 22802
rect 1119 22730 1237 22768
rect 1119 22696 1161 22730
rect 1195 22696 1237 22730
rect 1119 22658 1237 22696
rect 1119 22624 1161 22658
rect 1195 22624 1237 22658
rect 1119 22586 1237 22624
rect 1119 22552 1161 22586
rect 1195 22552 1237 22586
rect 1119 22514 1237 22552
rect 1119 22480 1161 22514
rect 1195 22480 1237 22514
rect 1119 22442 1237 22480
rect 1119 22408 1161 22442
rect 1195 22408 1237 22442
rect 1119 22370 1237 22408
rect 1119 22336 1161 22370
rect 1195 22336 1237 22370
rect 1119 22298 1237 22336
rect 1119 22264 1161 22298
rect 1195 22264 1237 22298
rect 1119 22226 1237 22264
rect 1119 22192 1161 22226
rect 1195 22192 1237 22226
rect 1119 22154 1237 22192
rect 1119 22120 1161 22154
rect 1195 22120 1237 22154
rect 1119 22082 1237 22120
rect 1119 22048 1161 22082
rect 1195 22048 1237 22082
rect 1119 22010 1237 22048
rect 1119 21976 1161 22010
rect 1195 21976 1237 22010
rect 1119 21938 1237 21976
rect 1119 21904 1161 21938
rect 1195 21904 1237 21938
rect 1119 21866 1237 21904
rect 1119 21832 1161 21866
rect 1195 21832 1237 21866
rect 1119 21794 1237 21832
rect 1119 21760 1161 21794
rect 1195 21760 1237 21794
rect 1119 21722 1237 21760
rect 1119 21688 1161 21722
rect 1195 21688 1237 21722
rect 1119 21650 1237 21688
rect 1119 21616 1161 21650
rect 1195 21616 1237 21650
rect 1119 21578 1237 21616
rect 1119 21544 1161 21578
rect 1195 21544 1237 21578
rect 1119 21506 1237 21544
rect 1119 21472 1161 21506
rect 1195 21472 1237 21506
rect 1119 21434 1237 21472
rect 1119 21400 1161 21434
rect 1195 21400 1237 21434
rect 1119 21362 1237 21400
rect 1119 21328 1161 21362
rect 1195 21328 1237 21362
rect 1119 21290 1237 21328
rect 1119 21256 1161 21290
rect 1195 21256 1237 21290
rect 1119 21218 1237 21256
rect 1119 21184 1161 21218
rect 1195 21184 1237 21218
rect 1119 21146 1237 21184
rect 1119 21112 1161 21146
rect 1195 21112 1237 21146
rect 1119 21074 1237 21112
rect 1119 21040 1161 21074
rect 1195 21040 1237 21074
rect 1119 21002 1237 21040
rect 1119 20968 1161 21002
rect 1195 20968 1237 21002
rect 1119 20930 1237 20968
rect 1119 20896 1161 20930
rect 1195 20896 1237 20930
rect 1119 20858 1237 20896
rect 1119 20824 1161 20858
rect 1195 20824 1237 20858
rect 1119 20786 1237 20824
rect 1119 20752 1161 20786
rect 1195 20752 1237 20786
rect 1119 20714 1237 20752
rect 1119 20680 1161 20714
rect 1195 20680 1237 20714
rect 1119 20642 1237 20680
rect 1119 20608 1161 20642
rect 1195 20608 1237 20642
rect 1119 20570 1237 20608
rect 1119 20536 1161 20570
rect 1195 20536 1237 20570
rect 1119 20498 1237 20536
rect 1119 20464 1161 20498
rect 1195 20464 1237 20498
rect 1119 20426 1237 20464
rect 1119 20392 1161 20426
rect 1195 20392 1237 20426
rect 1119 20354 1237 20392
rect 1119 20320 1161 20354
rect 1195 20320 1237 20354
rect 1119 20282 1237 20320
rect 1119 20248 1161 20282
rect 1195 20248 1237 20282
rect 1119 20210 1237 20248
rect 1119 20176 1161 20210
rect 1195 20176 1237 20210
rect 1119 20138 1237 20176
rect 1119 20104 1161 20138
rect 1195 20104 1237 20138
rect 1119 20066 1237 20104
rect 1119 20032 1161 20066
rect 1195 20032 1237 20066
rect 1119 19994 1237 20032
rect 1119 19960 1161 19994
rect 1195 19960 1237 19994
rect 1119 19922 1237 19960
rect 1119 19888 1161 19922
rect 1195 19888 1237 19922
rect 1119 19850 1237 19888
rect 1119 19816 1161 19850
rect 1195 19816 1237 19850
rect 1119 19778 1237 19816
rect 1119 19744 1161 19778
rect 1195 19744 1237 19778
rect 1119 19706 1237 19744
rect 1119 19672 1161 19706
rect 1195 19672 1237 19706
rect 1119 19634 1237 19672
rect 1119 19600 1161 19634
rect 1195 19600 1237 19634
rect 1119 19562 1237 19600
rect 1119 19528 1161 19562
rect 1195 19528 1237 19562
rect 1119 19490 1237 19528
rect 1119 19456 1161 19490
rect 1195 19456 1237 19490
rect 1119 19418 1237 19456
rect 1119 19384 1161 19418
rect 1195 19384 1237 19418
rect 1119 19346 1237 19384
rect 1119 19312 1161 19346
rect 1195 19312 1237 19346
rect 1119 19274 1237 19312
rect 1119 19240 1161 19274
rect 1195 19240 1237 19274
rect 1119 19202 1237 19240
rect 1119 19168 1161 19202
rect 1195 19168 1237 19202
rect 1119 19130 1237 19168
rect 1119 19096 1161 19130
rect 1195 19096 1237 19130
rect 1119 19058 1237 19096
rect 1119 19024 1161 19058
rect 1195 19024 1237 19058
rect 1119 18986 1237 19024
rect 1119 18952 1161 18986
rect 1195 18952 1237 18986
rect 1119 18914 1237 18952
rect 1119 18880 1161 18914
rect 1195 18880 1237 18914
rect 1119 18842 1237 18880
rect 1119 18808 1161 18842
rect 1195 18808 1237 18842
rect 1119 18770 1237 18808
rect 1119 18736 1161 18770
rect 1195 18736 1237 18770
rect 1119 18698 1237 18736
rect 1119 18664 1161 18698
rect 1195 18664 1237 18698
rect 1119 18626 1237 18664
rect 1119 18592 1161 18626
rect 1195 18592 1237 18626
rect 1119 18554 1237 18592
rect 1119 18520 1161 18554
rect 1195 18520 1237 18554
rect 1119 18482 1237 18520
rect 1119 18448 1161 18482
rect 1195 18448 1237 18482
rect 1119 18410 1237 18448
rect 1119 18376 1161 18410
rect 1195 18376 1237 18410
rect 1119 18338 1237 18376
rect 1119 18304 1161 18338
rect 1195 18304 1237 18338
rect 1119 18266 1237 18304
rect 1119 18232 1161 18266
rect 1195 18232 1237 18266
rect 1119 18194 1237 18232
rect 1119 18160 1161 18194
rect 1195 18160 1237 18194
rect 1119 18122 1237 18160
rect 1119 18088 1161 18122
rect 1195 18088 1237 18122
rect 1119 18050 1237 18088
rect 1119 18016 1161 18050
rect 1195 18016 1237 18050
rect 1119 17978 1237 18016
rect 1119 17944 1161 17978
rect 1195 17944 1237 17978
rect 1119 17906 1237 17944
rect 1119 17872 1161 17906
rect 1195 17872 1237 17906
rect 1119 17834 1237 17872
rect 1119 17800 1161 17834
rect 1195 17800 1237 17834
rect 1119 17762 1237 17800
rect 1119 17728 1161 17762
rect 1195 17728 1237 17762
rect 1119 17690 1237 17728
rect 1119 17656 1161 17690
rect 1195 17656 1237 17690
rect 1119 17618 1237 17656
rect 1119 17584 1161 17618
rect 1195 17584 1237 17618
rect 1119 17546 1237 17584
rect 1119 17512 1161 17546
rect 1195 17512 1237 17546
rect 1119 17474 1237 17512
rect 1119 17440 1161 17474
rect 1195 17440 1237 17474
rect 1119 17402 1237 17440
rect 1119 17368 1161 17402
rect 1195 17368 1237 17402
rect 1119 17330 1237 17368
rect 1119 17296 1161 17330
rect 1195 17296 1237 17330
rect 1119 17258 1237 17296
rect 1119 17224 1161 17258
rect 1195 17224 1237 17258
rect 1119 17186 1237 17224
rect 1119 17152 1161 17186
rect 1195 17152 1237 17186
rect 1119 17114 1237 17152
rect 1119 17080 1161 17114
rect 1195 17080 1237 17114
rect 1119 17042 1237 17080
rect 1119 17008 1161 17042
rect 1195 17008 1237 17042
rect 1119 16970 1237 17008
rect 1119 16936 1161 16970
rect 1195 16936 1237 16970
rect 1119 16898 1237 16936
rect 1119 16864 1161 16898
rect 1195 16864 1237 16898
rect 1119 16826 1237 16864
rect 1119 16792 1161 16826
rect 1195 16792 1237 16826
rect 1119 16754 1237 16792
rect 1119 16720 1161 16754
rect 1195 16720 1237 16754
rect 1119 16682 1237 16720
rect 1119 16648 1161 16682
rect 1195 16648 1237 16682
rect 1119 16610 1237 16648
rect 1119 16576 1161 16610
rect 1195 16576 1237 16610
rect 1119 16538 1237 16576
rect 1119 16504 1161 16538
rect 1195 16504 1237 16538
rect 1119 16466 1237 16504
rect 1119 16432 1161 16466
rect 1195 16432 1237 16466
rect 1119 16394 1237 16432
rect 1119 16360 1161 16394
rect 1195 16360 1237 16394
rect 1119 16322 1237 16360
rect 1119 16288 1161 16322
rect 1195 16288 1237 16322
rect 1119 16250 1237 16288
rect 1119 16216 1161 16250
rect 1195 16216 1237 16250
rect 1119 16178 1237 16216
rect 1119 16144 1161 16178
rect 1195 16144 1237 16178
rect 1119 16106 1237 16144
rect 1119 16072 1161 16106
rect 1195 16072 1237 16106
rect 1119 16034 1237 16072
rect 1119 16000 1161 16034
rect 1195 16000 1237 16034
rect 1119 15962 1237 16000
rect 1119 15928 1161 15962
rect 1195 15928 1237 15962
rect 1119 15890 1237 15928
rect 1119 15856 1161 15890
rect 1195 15856 1237 15890
rect 1119 15818 1237 15856
rect 1119 15784 1161 15818
rect 1195 15784 1237 15818
rect 1119 15746 1237 15784
rect 1119 15712 1161 15746
rect 1195 15712 1237 15746
rect 1119 15674 1237 15712
rect 1119 15640 1161 15674
rect 1195 15640 1237 15674
rect 1119 15602 1237 15640
rect 1119 15568 1161 15602
rect 1195 15568 1237 15602
rect 1119 15530 1237 15568
rect 1119 15496 1161 15530
rect 1195 15496 1237 15530
rect 1119 15458 1237 15496
rect 1119 15424 1161 15458
rect 1195 15424 1237 15458
rect 1119 15386 1237 15424
rect 1119 15352 1161 15386
rect 1195 15352 1237 15386
rect 1119 15314 1237 15352
rect 1119 15280 1161 15314
rect 1195 15280 1237 15314
rect 1119 15242 1237 15280
rect 1119 15208 1161 15242
rect 1195 15208 1237 15242
rect 1119 15170 1237 15208
rect 1119 15136 1161 15170
rect 1195 15136 1237 15170
rect 1119 15098 1237 15136
rect 1119 15064 1161 15098
rect 1195 15064 1237 15098
rect 1119 15026 1237 15064
rect 1119 14992 1161 15026
rect 1195 14992 1237 15026
rect 1119 14954 1237 14992
rect 1119 14920 1161 14954
rect 1195 14920 1237 14954
rect 1119 14882 1237 14920
rect 1119 14848 1161 14882
rect 1195 14848 1237 14882
rect 1119 14810 1237 14848
rect 1119 14776 1161 14810
rect 1195 14776 1237 14810
rect 1119 14738 1237 14776
rect 1119 14704 1161 14738
rect 1195 14704 1237 14738
rect 1119 14666 1237 14704
rect 1119 14632 1161 14666
rect 1195 14632 1237 14666
rect 1119 14594 1237 14632
rect 1119 14560 1161 14594
rect 1195 14560 1237 14594
rect 1119 14522 1237 14560
rect 1119 14488 1161 14522
rect 1195 14488 1237 14522
rect 1119 14450 1237 14488
rect 1119 14416 1161 14450
rect 1195 14416 1237 14450
rect 1119 14378 1237 14416
rect 1119 14344 1161 14378
rect 1195 14344 1237 14378
rect 1119 14306 1237 14344
rect 1119 14272 1161 14306
rect 1195 14272 1237 14306
rect 1119 14234 1237 14272
rect 1119 14200 1161 14234
rect 1195 14200 1237 14234
rect 1119 14162 1237 14200
rect 1119 14128 1161 14162
rect 1195 14128 1237 14162
rect 1119 14090 1237 14128
rect 1119 14056 1161 14090
rect 1195 14056 1237 14090
rect 1119 14018 1237 14056
rect 1119 13984 1161 14018
rect 1195 13984 1237 14018
rect 1119 13946 1237 13984
rect 1119 13912 1161 13946
rect 1195 13912 1237 13946
rect 1119 13874 1237 13912
rect 1119 13840 1161 13874
rect 1195 13840 1237 13874
rect 1119 13802 1237 13840
rect 1119 13768 1161 13802
rect 1195 13768 1237 13802
rect 1119 13730 1237 13768
rect 1119 13696 1161 13730
rect 1195 13696 1237 13730
rect 1119 13658 1237 13696
rect 1119 13624 1161 13658
rect 1195 13624 1237 13658
rect 1119 13586 1237 13624
rect 1119 13552 1161 13586
rect 1195 13552 1237 13586
rect 1119 13514 1237 13552
rect 1119 13480 1161 13514
rect 1195 13480 1237 13514
rect 1119 13442 1237 13480
rect 1119 13408 1161 13442
rect 1195 13408 1237 13442
rect 1119 13370 1237 13408
rect 1119 13336 1161 13370
rect 1195 13336 1237 13370
rect 1119 13298 1237 13336
rect 1119 13264 1161 13298
rect 1195 13264 1237 13298
rect 1119 13226 1237 13264
rect 1119 13192 1161 13226
rect 1195 13192 1237 13226
rect 1119 13154 1237 13192
rect 1119 13120 1161 13154
rect 1195 13120 1237 13154
rect 1119 13082 1237 13120
rect 1119 13048 1161 13082
rect 1195 13048 1237 13082
rect 1119 13010 1237 13048
rect 1119 12976 1161 13010
rect 1195 12976 1237 13010
rect 1119 12938 1237 12976
rect 1119 12904 1161 12938
rect 1195 12904 1237 12938
rect 1119 12866 1237 12904
rect 1119 12832 1161 12866
rect 1195 12832 1237 12866
rect 1119 12794 1237 12832
rect 1119 12760 1161 12794
rect 1195 12760 1237 12794
rect 1119 12722 1237 12760
rect 1119 12688 1161 12722
rect 1195 12688 1237 12722
rect 1119 12650 1237 12688
rect 1119 12616 1161 12650
rect 1195 12616 1237 12650
rect 1119 12578 1237 12616
rect 1119 12544 1161 12578
rect 1195 12544 1237 12578
rect 1119 12506 1237 12544
rect 1119 12472 1161 12506
rect 1195 12472 1237 12506
rect 1119 12434 1237 12472
rect 1119 12400 1161 12434
rect 1195 12400 1237 12434
rect 1119 12362 1237 12400
rect 1119 12328 1161 12362
rect 1195 12328 1237 12362
rect 1119 12290 1237 12328
rect 1119 12256 1161 12290
rect 1195 12256 1237 12290
rect 1119 12218 1237 12256
rect 1119 12184 1161 12218
rect 1195 12184 1237 12218
rect 1119 12146 1237 12184
rect 1119 12112 1161 12146
rect 1195 12112 1237 12146
rect 1119 12074 1237 12112
rect 1119 12040 1161 12074
rect 1195 12040 1237 12074
rect 1119 12002 1237 12040
rect 1119 11968 1161 12002
rect 1195 11968 1237 12002
rect 1119 11930 1237 11968
rect 1119 11896 1161 11930
rect 1195 11896 1237 11930
rect 1119 11858 1237 11896
rect 1119 11824 1161 11858
rect 1195 11824 1237 11858
rect 1119 11786 1237 11824
rect 1119 11752 1161 11786
rect 1195 11752 1237 11786
rect 1119 11714 1237 11752
rect 1119 11680 1161 11714
rect 1195 11680 1237 11714
rect 1119 11642 1237 11680
rect 1119 11608 1161 11642
rect 1195 11608 1237 11642
rect 1119 11570 1237 11608
rect 1119 11536 1161 11570
rect 1195 11536 1237 11570
rect 1119 11498 1237 11536
rect 1119 11464 1161 11498
rect 1195 11464 1237 11498
rect 1119 11426 1237 11464
rect 1119 11392 1161 11426
rect 1195 11392 1237 11426
rect 1119 11354 1237 11392
rect 1119 11320 1161 11354
rect 1195 11320 1237 11354
rect 1119 11282 1237 11320
rect 1119 11248 1161 11282
rect 1195 11248 1237 11282
rect 1119 11210 1237 11248
rect 1119 11176 1161 11210
rect 1195 11176 1237 11210
rect 1119 11138 1237 11176
rect 1119 11104 1161 11138
rect 1195 11104 1237 11138
rect 1119 11066 1237 11104
rect 1119 11032 1161 11066
rect 1195 11032 1237 11066
rect 1119 10994 1237 11032
rect 1119 10960 1161 10994
rect 1195 10960 1237 10994
rect 1119 10922 1237 10960
rect 1119 10888 1161 10922
rect 1195 10888 1237 10922
rect 1119 10850 1237 10888
rect 1119 10816 1161 10850
rect 1195 10816 1237 10850
rect 1119 10778 1237 10816
rect 1119 10744 1161 10778
rect 1195 10744 1237 10778
rect 1119 10706 1237 10744
rect 1119 10672 1161 10706
rect 1195 10672 1237 10706
rect 1119 10634 1237 10672
rect 1119 10600 1161 10634
rect 1195 10600 1237 10634
rect 1119 10562 1237 10600
rect 1119 10528 1161 10562
rect 1195 10528 1237 10562
rect 1119 10490 1237 10528
rect 1119 10456 1161 10490
rect 1195 10456 1237 10490
rect 1119 10418 1237 10456
rect 1119 10384 1161 10418
rect 1195 10384 1237 10418
rect 1119 10319 1237 10384
rect 13769 23381 13888 23428
rect 13769 23347 13809 23381
rect 13843 23347 13888 23381
rect 13769 23309 13888 23347
rect 13769 23275 13809 23309
rect 13843 23275 13888 23309
rect 13769 23237 13888 23275
rect 13769 23203 13809 23237
rect 13843 23203 13888 23237
rect 13769 23165 13888 23203
rect 13769 23131 13809 23165
rect 13843 23131 13888 23165
rect 13769 23093 13888 23131
rect 13769 23059 13809 23093
rect 13843 23059 13888 23093
rect 13769 23021 13888 23059
rect 13769 22987 13809 23021
rect 13843 22987 13888 23021
rect 13769 22949 13888 22987
rect 13769 22915 13809 22949
rect 13843 22915 13888 22949
rect 13769 22877 13888 22915
rect 13769 22843 13809 22877
rect 13843 22843 13888 22877
rect 13769 22805 13888 22843
rect 13769 22771 13809 22805
rect 13843 22771 13888 22805
rect 13769 22733 13888 22771
rect 13769 22699 13809 22733
rect 13843 22699 13888 22733
rect 13769 22661 13888 22699
rect 13769 22627 13809 22661
rect 13843 22627 13888 22661
rect 13769 22589 13888 22627
rect 13769 22555 13809 22589
rect 13843 22555 13888 22589
rect 13769 22517 13888 22555
rect 13769 22483 13809 22517
rect 13843 22483 13888 22517
rect 13769 22445 13888 22483
rect 13769 22411 13809 22445
rect 13843 22411 13888 22445
rect 13769 22373 13888 22411
rect 13769 22339 13809 22373
rect 13843 22339 13888 22373
rect 13769 22301 13888 22339
rect 13769 22267 13809 22301
rect 13843 22267 13888 22301
rect 13769 22229 13888 22267
rect 13769 22195 13809 22229
rect 13843 22195 13888 22229
rect 13769 22157 13888 22195
rect 13769 22123 13809 22157
rect 13843 22123 13888 22157
rect 13769 22085 13888 22123
rect 13769 22051 13809 22085
rect 13843 22051 13888 22085
rect 13769 22013 13888 22051
rect 13769 21979 13809 22013
rect 13843 21979 13888 22013
rect 13769 21941 13888 21979
rect 13769 21907 13809 21941
rect 13843 21907 13888 21941
rect 13769 21869 13888 21907
rect 13769 21835 13809 21869
rect 13843 21835 13888 21869
rect 13769 21797 13888 21835
rect 13769 21763 13809 21797
rect 13843 21763 13888 21797
rect 13769 21725 13888 21763
rect 13769 21691 13809 21725
rect 13843 21691 13888 21725
rect 13769 21653 13888 21691
rect 13769 21619 13809 21653
rect 13843 21619 13888 21653
rect 13769 21581 13888 21619
rect 13769 21547 13809 21581
rect 13843 21547 13888 21581
rect 13769 21509 13888 21547
rect 13769 21475 13809 21509
rect 13843 21475 13888 21509
rect 13769 21437 13888 21475
rect 13769 21403 13809 21437
rect 13843 21403 13888 21437
rect 13769 21365 13888 21403
rect 13769 21331 13809 21365
rect 13843 21331 13888 21365
rect 13769 21293 13888 21331
rect 13769 21259 13809 21293
rect 13843 21259 13888 21293
rect 13769 21221 13888 21259
rect 13769 21187 13809 21221
rect 13843 21187 13888 21221
rect 13769 21149 13888 21187
rect 13769 21115 13809 21149
rect 13843 21115 13888 21149
rect 13769 21077 13888 21115
rect 13769 21043 13809 21077
rect 13843 21043 13888 21077
rect 13769 21005 13888 21043
rect 13769 20971 13809 21005
rect 13843 20971 13888 21005
rect 13769 20933 13888 20971
rect 13769 20899 13809 20933
rect 13843 20899 13888 20933
rect 13769 20861 13888 20899
rect 13769 20827 13809 20861
rect 13843 20827 13888 20861
rect 13769 20789 13888 20827
rect 13769 20755 13809 20789
rect 13843 20755 13888 20789
rect 13769 20717 13888 20755
rect 13769 20683 13809 20717
rect 13843 20683 13888 20717
rect 13769 20645 13888 20683
rect 13769 20611 13809 20645
rect 13843 20611 13888 20645
rect 13769 20573 13888 20611
rect 13769 20539 13809 20573
rect 13843 20539 13888 20573
rect 13769 20501 13888 20539
rect 13769 20467 13809 20501
rect 13843 20467 13888 20501
rect 13769 20429 13888 20467
rect 13769 20395 13809 20429
rect 13843 20395 13888 20429
rect 13769 20357 13888 20395
rect 13769 20323 13809 20357
rect 13843 20323 13888 20357
rect 13769 20285 13888 20323
rect 13769 20251 13809 20285
rect 13843 20251 13888 20285
rect 13769 20213 13888 20251
rect 13769 20179 13809 20213
rect 13843 20179 13888 20213
rect 13769 20141 13888 20179
rect 13769 20107 13809 20141
rect 13843 20107 13888 20141
rect 13769 20069 13888 20107
rect 13769 20035 13809 20069
rect 13843 20035 13888 20069
rect 13769 19997 13888 20035
rect 13769 19963 13809 19997
rect 13843 19963 13888 19997
rect 13769 19925 13888 19963
rect 13769 19891 13809 19925
rect 13843 19891 13888 19925
rect 13769 19853 13888 19891
rect 13769 19819 13809 19853
rect 13843 19819 13888 19853
rect 13769 19781 13888 19819
rect 13769 19747 13809 19781
rect 13843 19747 13888 19781
rect 13769 19709 13888 19747
rect 13769 19675 13809 19709
rect 13843 19675 13888 19709
rect 13769 19637 13888 19675
rect 13769 19603 13809 19637
rect 13843 19603 13888 19637
rect 13769 19565 13888 19603
rect 13769 19531 13809 19565
rect 13843 19531 13888 19565
rect 13769 19493 13888 19531
rect 13769 19459 13809 19493
rect 13843 19459 13888 19493
rect 13769 19421 13888 19459
rect 13769 19387 13809 19421
rect 13843 19387 13888 19421
rect 13769 19349 13888 19387
rect 13769 19315 13809 19349
rect 13843 19315 13888 19349
rect 13769 19277 13888 19315
rect 13769 19243 13809 19277
rect 13843 19243 13888 19277
rect 13769 19205 13888 19243
rect 13769 19171 13809 19205
rect 13843 19171 13888 19205
rect 13769 19133 13888 19171
rect 13769 19099 13809 19133
rect 13843 19099 13888 19133
rect 13769 19061 13888 19099
rect 13769 19027 13809 19061
rect 13843 19027 13888 19061
rect 13769 18989 13888 19027
rect 13769 18955 13809 18989
rect 13843 18955 13888 18989
rect 13769 18917 13888 18955
rect 13769 18883 13809 18917
rect 13843 18883 13888 18917
rect 13769 18845 13888 18883
rect 13769 18811 13809 18845
rect 13843 18811 13888 18845
rect 13769 18773 13888 18811
rect 13769 18739 13809 18773
rect 13843 18739 13888 18773
rect 13769 18701 13888 18739
rect 13769 18667 13809 18701
rect 13843 18667 13888 18701
rect 13769 18629 13888 18667
rect 13769 18595 13809 18629
rect 13843 18595 13888 18629
rect 13769 18557 13888 18595
rect 13769 18523 13809 18557
rect 13843 18523 13888 18557
rect 13769 18485 13888 18523
rect 13769 18451 13809 18485
rect 13843 18451 13888 18485
rect 13769 18413 13888 18451
rect 13769 18379 13809 18413
rect 13843 18379 13888 18413
rect 13769 18341 13888 18379
rect 13769 18307 13809 18341
rect 13843 18307 13888 18341
rect 13769 18269 13888 18307
rect 13769 18235 13809 18269
rect 13843 18235 13888 18269
rect 13769 18197 13888 18235
rect 13769 18163 13809 18197
rect 13843 18163 13888 18197
rect 13769 18125 13888 18163
rect 13769 18091 13809 18125
rect 13843 18091 13888 18125
rect 13769 18053 13888 18091
rect 13769 18019 13809 18053
rect 13843 18019 13888 18053
rect 13769 17981 13888 18019
rect 13769 17947 13809 17981
rect 13843 17947 13888 17981
rect 13769 17909 13888 17947
rect 13769 17875 13809 17909
rect 13843 17875 13888 17909
rect 13769 17837 13888 17875
rect 13769 17803 13809 17837
rect 13843 17803 13888 17837
rect 13769 17765 13888 17803
rect 13769 17731 13809 17765
rect 13843 17731 13888 17765
rect 13769 17693 13888 17731
rect 13769 17659 13809 17693
rect 13843 17659 13888 17693
rect 13769 17621 13888 17659
rect 13769 17587 13809 17621
rect 13843 17587 13888 17621
rect 13769 17549 13888 17587
rect 13769 17515 13809 17549
rect 13843 17515 13888 17549
rect 13769 17477 13888 17515
rect 13769 17443 13809 17477
rect 13843 17443 13888 17477
rect 13769 17405 13888 17443
rect 13769 17371 13809 17405
rect 13843 17371 13888 17405
rect 13769 17333 13888 17371
rect 13769 17299 13809 17333
rect 13843 17299 13888 17333
rect 13769 17261 13888 17299
rect 13769 17227 13809 17261
rect 13843 17227 13888 17261
rect 13769 17189 13888 17227
rect 13769 17155 13809 17189
rect 13843 17155 13888 17189
rect 13769 17117 13888 17155
rect 13769 17083 13809 17117
rect 13843 17083 13888 17117
rect 13769 17045 13888 17083
rect 13769 17011 13809 17045
rect 13843 17011 13888 17045
rect 13769 16973 13888 17011
rect 13769 16939 13809 16973
rect 13843 16939 13888 16973
rect 13769 16901 13888 16939
rect 13769 16867 13809 16901
rect 13843 16867 13888 16901
rect 13769 16829 13888 16867
rect 13769 16795 13809 16829
rect 13843 16795 13888 16829
rect 13769 16757 13888 16795
rect 13769 16723 13809 16757
rect 13843 16723 13888 16757
rect 13769 16685 13888 16723
rect 13769 16651 13809 16685
rect 13843 16651 13888 16685
rect 13769 16613 13888 16651
rect 13769 16579 13809 16613
rect 13843 16579 13888 16613
rect 13769 16541 13888 16579
rect 13769 16507 13809 16541
rect 13843 16507 13888 16541
rect 13769 16469 13888 16507
rect 13769 16435 13809 16469
rect 13843 16435 13888 16469
rect 13769 16397 13888 16435
rect 13769 16363 13809 16397
rect 13843 16363 13888 16397
rect 13769 16325 13888 16363
rect 13769 16291 13809 16325
rect 13843 16291 13888 16325
rect 13769 16253 13888 16291
rect 13769 16219 13809 16253
rect 13843 16219 13888 16253
rect 13769 16181 13888 16219
rect 13769 16147 13809 16181
rect 13843 16147 13888 16181
rect 13769 16109 13888 16147
rect 13769 16075 13809 16109
rect 13843 16075 13888 16109
rect 13769 16037 13888 16075
rect 13769 16003 13809 16037
rect 13843 16003 13888 16037
rect 13769 15965 13888 16003
rect 13769 15931 13809 15965
rect 13843 15931 13888 15965
rect 13769 15893 13888 15931
rect 13769 15859 13809 15893
rect 13843 15859 13888 15893
rect 13769 15821 13888 15859
rect 13769 15787 13809 15821
rect 13843 15787 13888 15821
rect 13769 15749 13888 15787
rect 13769 15715 13809 15749
rect 13843 15715 13888 15749
rect 13769 15677 13888 15715
rect 13769 15643 13809 15677
rect 13843 15643 13888 15677
rect 13769 15605 13888 15643
rect 13769 15571 13809 15605
rect 13843 15571 13888 15605
rect 13769 15533 13888 15571
rect 13769 15499 13809 15533
rect 13843 15499 13888 15533
rect 13769 15461 13888 15499
rect 13769 15427 13809 15461
rect 13843 15427 13888 15461
rect 13769 15389 13888 15427
rect 13769 15355 13809 15389
rect 13843 15355 13888 15389
rect 13769 15317 13888 15355
rect 13769 15283 13809 15317
rect 13843 15283 13888 15317
rect 13769 15245 13888 15283
rect 13769 15211 13809 15245
rect 13843 15211 13888 15245
rect 13769 15173 13888 15211
rect 13769 15139 13809 15173
rect 13843 15139 13888 15173
rect 13769 15101 13888 15139
rect 13769 15067 13809 15101
rect 13843 15067 13888 15101
rect 13769 15029 13888 15067
rect 13769 14995 13809 15029
rect 13843 14995 13888 15029
rect 13769 14957 13888 14995
rect 13769 14923 13809 14957
rect 13843 14923 13888 14957
rect 13769 14885 13888 14923
rect 13769 14851 13809 14885
rect 13843 14851 13888 14885
rect 13769 14813 13888 14851
rect 13769 14779 13809 14813
rect 13843 14779 13888 14813
rect 13769 14741 13888 14779
rect 13769 14707 13809 14741
rect 13843 14707 13888 14741
rect 13769 14669 13888 14707
rect 13769 14635 13809 14669
rect 13843 14635 13888 14669
rect 13769 14597 13888 14635
rect 13769 14563 13809 14597
rect 13843 14563 13888 14597
rect 13769 14525 13888 14563
rect 13769 14491 13809 14525
rect 13843 14491 13888 14525
rect 13769 14453 13888 14491
rect 13769 14419 13809 14453
rect 13843 14419 13888 14453
rect 13769 14381 13888 14419
rect 13769 14347 13809 14381
rect 13843 14347 13888 14381
rect 13769 14309 13888 14347
rect 13769 14275 13809 14309
rect 13843 14275 13888 14309
rect 13769 14237 13888 14275
rect 13769 14203 13809 14237
rect 13843 14203 13888 14237
rect 13769 14165 13888 14203
rect 13769 14131 13809 14165
rect 13843 14131 13888 14165
rect 13769 14093 13888 14131
rect 13769 14059 13809 14093
rect 13843 14059 13888 14093
rect 13769 14021 13888 14059
rect 13769 13987 13809 14021
rect 13843 13987 13888 14021
rect 13769 13949 13888 13987
rect 13769 13915 13809 13949
rect 13843 13915 13888 13949
rect 13769 13877 13888 13915
rect 13769 13843 13809 13877
rect 13843 13843 13888 13877
rect 13769 13805 13888 13843
rect 13769 13771 13809 13805
rect 13843 13771 13888 13805
rect 13769 13733 13888 13771
rect 13769 13699 13809 13733
rect 13843 13699 13888 13733
rect 13769 13661 13888 13699
rect 13769 13627 13809 13661
rect 13843 13627 13888 13661
rect 13769 13589 13888 13627
rect 13769 13555 13809 13589
rect 13843 13555 13888 13589
rect 13769 13517 13888 13555
rect 13769 13483 13809 13517
rect 13843 13483 13888 13517
rect 13769 13445 13888 13483
rect 13769 13411 13809 13445
rect 13843 13411 13888 13445
rect 13769 13373 13888 13411
rect 13769 13339 13809 13373
rect 13843 13339 13888 13373
rect 13769 13301 13888 13339
rect 13769 13267 13809 13301
rect 13843 13267 13888 13301
rect 13769 13229 13888 13267
rect 13769 13195 13809 13229
rect 13843 13195 13888 13229
rect 13769 13157 13888 13195
rect 13769 13123 13809 13157
rect 13843 13123 13888 13157
rect 13769 13085 13888 13123
rect 13769 13051 13809 13085
rect 13843 13051 13888 13085
rect 13769 13013 13888 13051
rect 13769 12979 13809 13013
rect 13843 12979 13888 13013
rect 13769 12941 13888 12979
rect 13769 12907 13809 12941
rect 13843 12907 13888 12941
rect 13769 12869 13888 12907
rect 13769 12835 13809 12869
rect 13843 12835 13888 12869
rect 13769 12797 13888 12835
rect 13769 12763 13809 12797
rect 13843 12763 13888 12797
rect 13769 12725 13888 12763
rect 13769 12691 13809 12725
rect 13843 12691 13888 12725
rect 13769 12653 13888 12691
rect 13769 12619 13809 12653
rect 13843 12619 13888 12653
rect 13769 12581 13888 12619
rect 13769 12547 13809 12581
rect 13843 12547 13888 12581
rect 13769 12509 13888 12547
rect 13769 12475 13809 12509
rect 13843 12475 13888 12509
rect 13769 12437 13888 12475
rect 13769 12403 13809 12437
rect 13843 12403 13888 12437
rect 13769 12365 13888 12403
rect 13769 12331 13809 12365
rect 13843 12331 13888 12365
rect 13769 12293 13888 12331
rect 13769 12259 13809 12293
rect 13843 12259 13888 12293
rect 13769 12221 13888 12259
rect 13769 12187 13809 12221
rect 13843 12187 13888 12221
rect 13769 12149 13888 12187
rect 13769 12115 13809 12149
rect 13843 12115 13888 12149
rect 13769 12077 13888 12115
rect 13769 12043 13809 12077
rect 13843 12043 13888 12077
rect 13769 12005 13888 12043
rect 13769 11971 13809 12005
rect 13843 11971 13888 12005
rect 13769 11933 13888 11971
rect 13769 11899 13809 11933
rect 13843 11899 13888 11933
rect 13769 11861 13888 11899
rect 13769 11827 13809 11861
rect 13843 11827 13888 11861
rect 13769 11789 13888 11827
rect 13769 11755 13809 11789
rect 13843 11755 13888 11789
rect 13769 11717 13888 11755
rect 13769 11683 13809 11717
rect 13843 11683 13888 11717
rect 13769 11645 13888 11683
rect 13769 11611 13809 11645
rect 13843 11611 13888 11645
rect 13769 11573 13888 11611
rect 13769 11539 13809 11573
rect 13843 11539 13888 11573
rect 13769 11501 13888 11539
rect 13769 11467 13809 11501
rect 13843 11467 13888 11501
rect 13769 11429 13888 11467
rect 13769 11395 13809 11429
rect 13843 11395 13888 11429
rect 13769 11357 13888 11395
rect 13769 11323 13809 11357
rect 13843 11323 13888 11357
rect 13769 11285 13888 11323
rect 13769 11251 13809 11285
rect 13843 11251 13888 11285
rect 13769 11213 13888 11251
rect 13769 11179 13809 11213
rect 13843 11179 13888 11213
rect 13769 11141 13888 11179
rect 13769 11107 13809 11141
rect 13843 11107 13888 11141
rect 13769 11069 13888 11107
rect 13769 11035 13809 11069
rect 13843 11035 13888 11069
rect 13769 10997 13888 11035
rect 13769 10963 13809 10997
rect 13843 10963 13888 10997
rect 13769 10925 13888 10963
rect 13769 10891 13809 10925
rect 13843 10891 13888 10925
rect 13769 10853 13888 10891
rect 13769 10819 13809 10853
rect 13843 10819 13888 10853
rect 13769 10781 13888 10819
rect 13769 10747 13809 10781
rect 13843 10747 13888 10781
rect 13769 10709 13888 10747
rect 13769 10675 13809 10709
rect 13843 10675 13888 10709
rect 13769 10637 13888 10675
rect 13769 10603 13809 10637
rect 13843 10603 13888 10637
rect 13769 10565 13888 10603
rect 13769 10531 13809 10565
rect 13843 10531 13888 10565
rect 13769 10493 13888 10531
rect 13769 10459 13809 10493
rect 13843 10459 13888 10493
rect 13769 10421 13888 10459
rect 13769 10387 13809 10421
rect 13843 10387 13888 10421
rect 13769 10319 13888 10387
rect 1119 10278 13888 10319
rect 1119 10244 1298 10278
rect 1332 10244 1370 10278
rect 1404 10244 1442 10278
rect 1476 10244 1514 10278
rect 1548 10244 1586 10278
rect 1620 10244 1658 10278
rect 1692 10244 1730 10278
rect 1764 10244 1802 10278
rect 1836 10244 1874 10278
rect 1908 10244 1946 10278
rect 1980 10244 2018 10278
rect 2052 10244 2090 10278
rect 2124 10244 2162 10278
rect 2196 10244 2234 10278
rect 2268 10244 2306 10278
rect 2340 10244 2378 10278
rect 2412 10244 2450 10278
rect 2484 10244 2522 10278
rect 2556 10244 2594 10278
rect 2628 10244 2666 10278
rect 2700 10244 2738 10278
rect 2772 10244 2810 10278
rect 2844 10244 2882 10278
rect 2916 10244 2954 10278
rect 2988 10244 3026 10278
rect 3060 10244 3098 10278
rect 3132 10244 3170 10278
rect 3204 10244 3242 10278
rect 3276 10244 3314 10278
rect 3348 10244 3386 10278
rect 3420 10244 3458 10278
rect 3492 10244 3530 10278
rect 3564 10244 3602 10278
rect 3636 10244 3674 10278
rect 3708 10244 3746 10278
rect 3780 10244 3818 10278
rect 3852 10244 3890 10278
rect 3924 10244 3962 10278
rect 3996 10244 4034 10278
rect 4068 10244 4106 10278
rect 4140 10244 4178 10278
rect 4212 10244 4250 10278
rect 4284 10244 4322 10278
rect 4356 10244 4394 10278
rect 4428 10244 4466 10278
rect 4500 10244 4538 10278
rect 4572 10244 4610 10278
rect 4644 10244 4682 10278
rect 4716 10244 4754 10278
rect 4788 10244 4826 10278
rect 4860 10244 4898 10278
rect 4932 10244 4970 10278
rect 5004 10244 5042 10278
rect 5076 10244 5114 10278
rect 5148 10244 5186 10278
rect 5220 10244 5258 10278
rect 5292 10244 5330 10278
rect 5364 10244 5402 10278
rect 5436 10244 5474 10278
rect 5508 10244 5546 10278
rect 5580 10244 5618 10278
rect 5652 10244 5690 10278
rect 5724 10244 5762 10278
rect 5796 10244 5834 10278
rect 5868 10244 5906 10278
rect 5940 10244 5978 10278
rect 6012 10244 6050 10278
rect 6084 10244 6122 10278
rect 6156 10244 6194 10278
rect 6228 10244 6266 10278
rect 6300 10244 6338 10278
rect 6372 10244 6410 10278
rect 6444 10244 6482 10278
rect 6516 10244 6554 10278
rect 6588 10244 6626 10278
rect 6660 10244 6698 10278
rect 6732 10244 6770 10278
rect 6804 10244 6842 10278
rect 6876 10244 6914 10278
rect 6948 10244 6986 10278
rect 7020 10244 7058 10278
rect 7092 10244 7130 10278
rect 7164 10244 7202 10278
rect 7236 10244 7274 10278
rect 7308 10244 7346 10278
rect 7380 10244 7418 10278
rect 7452 10244 7490 10278
rect 7524 10244 7562 10278
rect 7596 10244 7634 10278
rect 7668 10244 7706 10278
rect 7740 10244 7778 10278
rect 7812 10244 7850 10278
rect 7884 10244 7922 10278
rect 7956 10244 7994 10278
rect 8028 10244 8066 10278
rect 8100 10244 8138 10278
rect 8172 10244 8210 10278
rect 8244 10244 8282 10278
rect 8316 10244 8354 10278
rect 8388 10244 8426 10278
rect 8460 10244 8498 10278
rect 8532 10244 8570 10278
rect 8604 10244 8642 10278
rect 8676 10244 8714 10278
rect 8748 10244 8786 10278
rect 8820 10244 8858 10278
rect 8892 10244 8930 10278
rect 8964 10244 9002 10278
rect 9036 10244 9074 10278
rect 9108 10244 9146 10278
rect 9180 10244 9218 10278
rect 9252 10244 9290 10278
rect 9324 10244 9362 10278
rect 9396 10244 9434 10278
rect 9468 10244 9506 10278
rect 9540 10244 9578 10278
rect 9612 10244 9650 10278
rect 9684 10244 9722 10278
rect 9756 10244 9794 10278
rect 9828 10244 9866 10278
rect 9900 10244 9938 10278
rect 9972 10244 10010 10278
rect 10044 10244 10082 10278
rect 10116 10244 10154 10278
rect 10188 10244 10226 10278
rect 10260 10244 10298 10278
rect 10332 10244 10370 10278
rect 10404 10244 10442 10278
rect 10476 10244 10514 10278
rect 10548 10244 10586 10278
rect 10620 10244 10658 10278
rect 10692 10244 10730 10278
rect 10764 10244 10802 10278
rect 10836 10244 10874 10278
rect 10908 10244 10946 10278
rect 10980 10244 11018 10278
rect 11052 10244 11090 10278
rect 11124 10244 11162 10278
rect 11196 10244 11234 10278
rect 11268 10244 11306 10278
rect 11340 10244 11378 10278
rect 11412 10244 11450 10278
rect 11484 10244 11522 10278
rect 11556 10244 11594 10278
rect 11628 10244 11666 10278
rect 11700 10244 11738 10278
rect 11772 10244 11810 10278
rect 11844 10244 11882 10278
rect 11916 10244 11954 10278
rect 11988 10244 12026 10278
rect 12060 10244 12098 10278
rect 12132 10244 12170 10278
rect 12204 10244 12242 10278
rect 12276 10244 12314 10278
rect 12348 10244 12386 10278
rect 12420 10244 12458 10278
rect 12492 10244 12530 10278
rect 12564 10244 12602 10278
rect 12636 10244 12674 10278
rect 12708 10244 12746 10278
rect 12780 10244 12818 10278
rect 12852 10244 12890 10278
rect 12924 10244 12962 10278
rect 12996 10244 13034 10278
rect 13068 10244 13106 10278
rect 13140 10244 13178 10278
rect 13212 10244 13250 10278
rect 13284 10244 13322 10278
rect 13356 10244 13394 10278
rect 13428 10244 13466 10278
rect 13500 10244 13538 10278
rect 13572 10244 13610 10278
rect 13644 10244 13682 10278
rect 13716 10244 13888 10278
rect 1119 10201 13888 10244
rect 14099 23421 14219 23459
rect 14099 23387 14122 23421
rect 14156 23387 14219 23421
rect 14099 23349 14219 23387
rect 14099 23315 14122 23349
rect 14156 23315 14219 23349
rect 14099 23277 14219 23315
rect 14099 23243 14122 23277
rect 14156 23243 14219 23277
rect 14099 23205 14219 23243
rect 14099 23171 14122 23205
rect 14156 23171 14219 23205
rect 14099 23133 14219 23171
rect 14099 23099 14122 23133
rect 14156 23099 14219 23133
rect 14099 23061 14219 23099
rect 14099 23027 14122 23061
rect 14156 23027 14219 23061
rect 14099 22989 14219 23027
rect 14099 22955 14122 22989
rect 14156 22955 14219 22989
rect 14099 22917 14219 22955
rect 14099 22883 14122 22917
rect 14156 22883 14219 22917
rect 14099 22845 14219 22883
rect 14099 22811 14122 22845
rect 14156 22811 14219 22845
rect 14099 22773 14219 22811
rect 14099 22739 14122 22773
rect 14156 22739 14219 22773
rect 14099 22701 14219 22739
rect 14099 22667 14122 22701
rect 14156 22667 14219 22701
rect 14099 22629 14219 22667
rect 14099 22595 14122 22629
rect 14156 22595 14219 22629
rect 14099 22557 14219 22595
rect 14099 22523 14122 22557
rect 14156 22523 14219 22557
rect 14099 22485 14219 22523
rect 14099 22451 14122 22485
rect 14156 22451 14219 22485
rect 14099 22413 14219 22451
rect 14099 22379 14122 22413
rect 14156 22379 14219 22413
rect 14099 22341 14219 22379
rect 14099 22307 14122 22341
rect 14156 22307 14219 22341
rect 14099 22269 14219 22307
rect 14099 22235 14122 22269
rect 14156 22235 14219 22269
rect 14099 22197 14219 22235
rect 14099 22163 14122 22197
rect 14156 22163 14219 22197
rect 14099 22125 14219 22163
rect 14099 22091 14122 22125
rect 14156 22091 14219 22125
rect 14099 22053 14219 22091
rect 14099 22019 14122 22053
rect 14156 22019 14219 22053
rect 14099 21981 14219 22019
rect 14099 21947 14122 21981
rect 14156 21947 14219 21981
rect 14099 21909 14219 21947
rect 14099 21875 14122 21909
rect 14156 21875 14219 21909
rect 14099 21837 14219 21875
rect 14099 21803 14122 21837
rect 14156 21803 14219 21837
rect 14099 21765 14219 21803
rect 14099 21731 14122 21765
rect 14156 21731 14219 21765
rect 14099 21693 14219 21731
rect 14099 21659 14122 21693
rect 14156 21659 14219 21693
rect 14099 21621 14219 21659
rect 14099 21587 14122 21621
rect 14156 21587 14219 21621
rect 14099 21549 14219 21587
rect 14099 21515 14122 21549
rect 14156 21515 14219 21549
rect 14099 21477 14219 21515
rect 14099 21443 14122 21477
rect 14156 21443 14219 21477
rect 14099 21405 14219 21443
rect 14099 21371 14122 21405
rect 14156 21371 14219 21405
rect 14099 21333 14219 21371
rect 14099 21299 14122 21333
rect 14156 21299 14219 21333
rect 14099 21261 14219 21299
rect 14099 21227 14122 21261
rect 14156 21227 14219 21261
rect 14099 21189 14219 21227
rect 14099 21155 14122 21189
rect 14156 21155 14219 21189
rect 14099 21117 14219 21155
rect 14099 21083 14122 21117
rect 14156 21083 14219 21117
rect 14099 21045 14219 21083
rect 14099 21011 14122 21045
rect 14156 21011 14219 21045
rect 14099 20973 14219 21011
rect 14099 20939 14122 20973
rect 14156 20939 14219 20973
rect 14099 20901 14219 20939
rect 14099 20867 14122 20901
rect 14156 20867 14219 20901
rect 14099 20829 14219 20867
rect 14099 20795 14122 20829
rect 14156 20795 14219 20829
rect 14099 20757 14219 20795
rect 14099 20723 14122 20757
rect 14156 20723 14219 20757
rect 14099 20685 14219 20723
rect 14099 20651 14122 20685
rect 14156 20651 14219 20685
rect 14099 20613 14219 20651
rect 14099 20579 14122 20613
rect 14156 20579 14219 20613
rect 14099 20541 14219 20579
rect 14099 20507 14122 20541
rect 14156 20507 14219 20541
rect 14099 20469 14219 20507
rect 14099 20435 14122 20469
rect 14156 20435 14219 20469
rect 14099 20397 14219 20435
rect 14099 20363 14122 20397
rect 14156 20363 14219 20397
rect 14099 20325 14219 20363
rect 14099 20291 14122 20325
rect 14156 20291 14219 20325
rect 14099 20253 14219 20291
rect 14099 20219 14122 20253
rect 14156 20219 14219 20253
rect 14099 20181 14219 20219
rect 14099 20147 14122 20181
rect 14156 20147 14219 20181
rect 14099 20109 14219 20147
rect 14099 20075 14122 20109
rect 14156 20075 14219 20109
rect 14099 20037 14219 20075
rect 14099 20003 14122 20037
rect 14156 20003 14219 20037
rect 14099 19965 14219 20003
rect 14099 19931 14122 19965
rect 14156 19931 14219 19965
rect 14099 19893 14219 19931
rect 14099 19859 14122 19893
rect 14156 19859 14219 19893
rect 14099 19821 14219 19859
rect 14099 19787 14122 19821
rect 14156 19787 14219 19821
rect 14099 19749 14219 19787
rect 14099 19715 14122 19749
rect 14156 19715 14219 19749
rect 14099 19677 14219 19715
rect 14099 19643 14122 19677
rect 14156 19643 14219 19677
rect 14099 19605 14219 19643
rect 14099 19571 14122 19605
rect 14156 19571 14219 19605
rect 14099 19533 14219 19571
rect 14099 19499 14122 19533
rect 14156 19499 14219 19533
rect 14099 19461 14219 19499
rect 14099 19427 14122 19461
rect 14156 19427 14219 19461
rect 14099 19389 14219 19427
rect 14099 19355 14122 19389
rect 14156 19355 14219 19389
rect 14099 19317 14219 19355
rect 14099 19283 14122 19317
rect 14156 19283 14219 19317
rect 14099 19245 14219 19283
rect 14099 19211 14122 19245
rect 14156 19211 14219 19245
rect 14099 19173 14219 19211
rect 14099 19139 14122 19173
rect 14156 19139 14219 19173
rect 14099 19101 14219 19139
rect 14099 19067 14122 19101
rect 14156 19067 14219 19101
rect 14099 19029 14219 19067
rect 14099 18995 14122 19029
rect 14156 18995 14219 19029
rect 14099 18957 14219 18995
rect 14099 18923 14122 18957
rect 14156 18923 14219 18957
rect 14099 18885 14219 18923
rect 14099 18851 14122 18885
rect 14156 18851 14219 18885
rect 14099 18813 14219 18851
rect 14099 18779 14122 18813
rect 14156 18779 14219 18813
rect 14099 18741 14219 18779
rect 14099 18707 14122 18741
rect 14156 18707 14219 18741
rect 14099 18669 14219 18707
rect 14099 18635 14122 18669
rect 14156 18635 14219 18669
rect 14099 18597 14219 18635
rect 14099 18563 14122 18597
rect 14156 18563 14219 18597
rect 14099 18525 14219 18563
rect 14099 18491 14122 18525
rect 14156 18491 14219 18525
rect 14099 18453 14219 18491
rect 14099 18419 14122 18453
rect 14156 18419 14219 18453
rect 14099 18381 14219 18419
rect 14099 18347 14122 18381
rect 14156 18347 14219 18381
rect 14099 18309 14219 18347
rect 14099 18275 14122 18309
rect 14156 18275 14219 18309
rect 14099 18237 14219 18275
rect 14099 18203 14122 18237
rect 14156 18203 14219 18237
rect 14099 18165 14219 18203
rect 14099 18131 14122 18165
rect 14156 18131 14219 18165
rect 14099 18093 14219 18131
rect 14099 18059 14122 18093
rect 14156 18059 14219 18093
rect 14099 18021 14219 18059
rect 14099 17987 14122 18021
rect 14156 17987 14219 18021
rect 14099 17949 14219 17987
rect 14099 17915 14122 17949
rect 14156 17915 14219 17949
rect 14099 17877 14219 17915
rect 14099 17843 14122 17877
rect 14156 17843 14219 17877
rect 14099 17805 14219 17843
rect 14099 17771 14122 17805
rect 14156 17771 14219 17805
rect 14099 17733 14219 17771
rect 14099 17699 14122 17733
rect 14156 17699 14219 17733
rect 14099 17661 14219 17699
rect 14099 17627 14122 17661
rect 14156 17627 14219 17661
rect 14099 17589 14219 17627
rect 14099 17555 14122 17589
rect 14156 17555 14219 17589
rect 14099 17517 14219 17555
rect 14099 17483 14122 17517
rect 14156 17483 14219 17517
rect 14099 17445 14219 17483
rect 14099 17411 14122 17445
rect 14156 17411 14219 17445
rect 14099 17373 14219 17411
rect 14099 17339 14122 17373
rect 14156 17339 14219 17373
rect 14099 17301 14219 17339
rect 14099 17267 14122 17301
rect 14156 17267 14219 17301
rect 14099 17229 14219 17267
rect 14099 17195 14122 17229
rect 14156 17195 14219 17229
rect 14099 17157 14219 17195
rect 14099 17123 14122 17157
rect 14156 17123 14219 17157
rect 14099 17085 14219 17123
rect 14099 17051 14122 17085
rect 14156 17051 14219 17085
rect 14099 17013 14219 17051
rect 14099 16979 14122 17013
rect 14156 16979 14219 17013
rect 14099 16941 14219 16979
rect 14099 16907 14122 16941
rect 14156 16907 14219 16941
rect 14099 16869 14219 16907
rect 14099 16835 14122 16869
rect 14156 16835 14219 16869
rect 14099 16797 14219 16835
rect 14099 16763 14122 16797
rect 14156 16763 14219 16797
rect 14099 16725 14219 16763
rect 14099 16691 14122 16725
rect 14156 16691 14219 16725
rect 14099 16653 14219 16691
rect 14099 16619 14122 16653
rect 14156 16619 14219 16653
rect 14099 16581 14219 16619
rect 14099 16547 14122 16581
rect 14156 16547 14219 16581
rect 14099 16509 14219 16547
rect 14099 16475 14122 16509
rect 14156 16475 14219 16509
rect 14099 16437 14219 16475
rect 14099 16403 14122 16437
rect 14156 16403 14219 16437
rect 14099 16365 14219 16403
rect 14099 16331 14122 16365
rect 14156 16331 14219 16365
rect 14099 16293 14219 16331
rect 14099 16259 14122 16293
rect 14156 16259 14219 16293
rect 14099 16221 14219 16259
rect 14099 16187 14122 16221
rect 14156 16187 14219 16221
rect 14099 16149 14219 16187
rect 14099 16115 14122 16149
rect 14156 16115 14219 16149
rect 14099 16077 14219 16115
rect 14099 16043 14122 16077
rect 14156 16043 14219 16077
rect 14099 16005 14219 16043
rect 14099 15971 14122 16005
rect 14156 15971 14219 16005
rect 14099 15933 14219 15971
rect 14099 15899 14122 15933
rect 14156 15899 14219 15933
rect 14099 15861 14219 15899
rect 14099 15827 14122 15861
rect 14156 15827 14219 15861
rect 14099 15789 14219 15827
rect 14099 15755 14122 15789
rect 14156 15755 14219 15789
rect 14099 15717 14219 15755
rect 14099 15683 14122 15717
rect 14156 15683 14219 15717
rect 14099 15645 14219 15683
rect 14099 15611 14122 15645
rect 14156 15611 14219 15645
rect 14099 15573 14219 15611
rect 14099 15539 14122 15573
rect 14156 15539 14219 15573
rect 14099 15501 14219 15539
rect 14099 15467 14122 15501
rect 14156 15467 14219 15501
rect 14099 15429 14219 15467
rect 14099 15395 14122 15429
rect 14156 15395 14219 15429
rect 14099 15357 14219 15395
rect 14099 15323 14122 15357
rect 14156 15323 14219 15357
rect 14099 15285 14219 15323
rect 14099 15251 14122 15285
rect 14156 15251 14219 15285
rect 14099 15213 14219 15251
rect 14099 15179 14122 15213
rect 14156 15179 14219 15213
rect 14099 15141 14219 15179
rect 14099 15107 14122 15141
rect 14156 15107 14219 15141
rect 14099 15069 14219 15107
rect 14099 15035 14122 15069
rect 14156 15035 14219 15069
rect 14099 14997 14219 15035
rect 14099 14963 14122 14997
rect 14156 14963 14219 14997
rect 14099 14925 14219 14963
rect 14099 14891 14122 14925
rect 14156 14891 14219 14925
rect 14099 14853 14219 14891
rect 14099 14819 14122 14853
rect 14156 14819 14219 14853
rect 14099 14781 14219 14819
rect 14099 14747 14122 14781
rect 14156 14747 14219 14781
rect 14099 14709 14219 14747
rect 14099 14675 14122 14709
rect 14156 14675 14219 14709
rect 14099 14637 14219 14675
rect 14099 14603 14122 14637
rect 14156 14603 14219 14637
rect 14099 14565 14219 14603
rect 14099 14531 14122 14565
rect 14156 14531 14219 14565
rect 14099 14493 14219 14531
rect 14099 14459 14122 14493
rect 14156 14459 14219 14493
rect 14099 14421 14219 14459
rect 14099 14387 14122 14421
rect 14156 14387 14219 14421
rect 14099 14349 14219 14387
rect 14099 14315 14122 14349
rect 14156 14315 14219 14349
rect 14099 14277 14219 14315
rect 14099 14243 14122 14277
rect 14156 14243 14219 14277
rect 14099 14205 14219 14243
rect 14099 14171 14122 14205
rect 14156 14171 14219 14205
rect 14099 14133 14219 14171
rect 14099 14099 14122 14133
rect 14156 14099 14219 14133
rect 14099 14061 14219 14099
rect 14099 14027 14122 14061
rect 14156 14027 14219 14061
rect 14099 13989 14219 14027
rect 14099 13955 14122 13989
rect 14156 13955 14219 13989
rect 14099 13917 14219 13955
rect 14099 13883 14122 13917
rect 14156 13883 14219 13917
rect 14099 13845 14219 13883
rect 14099 13811 14122 13845
rect 14156 13811 14219 13845
rect 14099 13773 14219 13811
rect 14099 13739 14122 13773
rect 14156 13739 14219 13773
rect 14099 13701 14219 13739
rect 14099 13667 14122 13701
rect 14156 13667 14219 13701
rect 14099 13629 14219 13667
rect 14099 13595 14122 13629
rect 14156 13595 14219 13629
rect 14099 13557 14219 13595
rect 14099 13523 14122 13557
rect 14156 13523 14219 13557
rect 14099 13485 14219 13523
rect 14099 13451 14122 13485
rect 14156 13451 14219 13485
rect 14099 13413 14219 13451
rect 14099 13379 14122 13413
rect 14156 13379 14219 13413
rect 14099 13341 14219 13379
rect 14099 13307 14122 13341
rect 14156 13307 14219 13341
rect 14099 13269 14219 13307
rect 14099 13235 14122 13269
rect 14156 13235 14219 13269
rect 14099 13197 14219 13235
rect 14099 13163 14122 13197
rect 14156 13163 14219 13197
rect 14099 13125 14219 13163
rect 14099 13091 14122 13125
rect 14156 13091 14219 13125
rect 14099 13053 14219 13091
rect 14099 13019 14122 13053
rect 14156 13019 14219 13053
rect 14099 12981 14219 13019
rect 14099 12947 14122 12981
rect 14156 12947 14219 12981
rect 14099 12909 14219 12947
rect 14099 12875 14122 12909
rect 14156 12875 14219 12909
rect 14099 12837 14219 12875
rect 14099 12803 14122 12837
rect 14156 12803 14219 12837
rect 14099 12765 14219 12803
rect 14099 12731 14122 12765
rect 14156 12731 14219 12765
rect 14099 12693 14219 12731
rect 14099 12659 14122 12693
rect 14156 12659 14219 12693
rect 14099 12621 14219 12659
rect 14099 12587 14122 12621
rect 14156 12587 14219 12621
rect 14099 12549 14219 12587
rect 14099 12515 14122 12549
rect 14156 12515 14219 12549
rect 14099 12477 14219 12515
rect 14099 12443 14122 12477
rect 14156 12443 14219 12477
rect 14099 12405 14219 12443
rect 14099 12371 14122 12405
rect 14156 12371 14219 12405
rect 14099 12333 14219 12371
rect 14099 12299 14122 12333
rect 14156 12299 14219 12333
rect 14099 12261 14219 12299
rect 14099 12227 14122 12261
rect 14156 12227 14219 12261
rect 14099 12189 14219 12227
rect 14099 12155 14122 12189
rect 14156 12155 14219 12189
rect 14099 12117 14219 12155
rect 14099 12083 14122 12117
rect 14156 12083 14219 12117
rect 14099 12045 14219 12083
rect 14099 12011 14122 12045
rect 14156 12011 14219 12045
rect 14099 11973 14219 12011
rect 14099 11939 14122 11973
rect 14156 11939 14219 11973
rect 14099 11901 14219 11939
rect 14099 11867 14122 11901
rect 14156 11867 14219 11901
rect 14099 11829 14219 11867
rect 14099 11795 14122 11829
rect 14156 11795 14219 11829
rect 14099 11757 14219 11795
rect 14099 11723 14122 11757
rect 14156 11723 14219 11757
rect 14099 11685 14219 11723
rect 14099 11651 14122 11685
rect 14156 11651 14219 11685
rect 14099 11613 14219 11651
rect 14099 11579 14122 11613
rect 14156 11579 14219 11613
rect 14099 11541 14219 11579
rect 14099 11507 14122 11541
rect 14156 11507 14219 11541
rect 14099 11469 14219 11507
rect 14099 11435 14122 11469
rect 14156 11435 14219 11469
rect 14099 11397 14219 11435
rect 14099 11363 14122 11397
rect 14156 11363 14219 11397
rect 14099 11325 14219 11363
rect 14099 11291 14122 11325
rect 14156 11291 14219 11325
rect 14099 11253 14219 11291
rect 14099 11219 14122 11253
rect 14156 11219 14219 11253
rect 14099 11181 14219 11219
rect 14099 11147 14122 11181
rect 14156 11147 14219 11181
rect 14099 11109 14219 11147
rect 14099 11075 14122 11109
rect 14156 11075 14219 11109
rect 14099 11037 14219 11075
rect 14099 11003 14122 11037
rect 14156 11003 14219 11037
rect 14099 10965 14219 11003
rect 14099 10931 14122 10965
rect 14156 10931 14219 10965
rect 14099 10893 14219 10931
rect 14099 10859 14122 10893
rect 14156 10859 14219 10893
rect 14099 10821 14219 10859
rect 14099 10787 14122 10821
rect 14156 10787 14219 10821
rect 14099 10749 14219 10787
rect 14099 10715 14122 10749
rect 14156 10715 14219 10749
rect 14099 10677 14219 10715
rect 14099 10643 14122 10677
rect 14156 10643 14219 10677
rect 14099 10605 14219 10643
rect 14099 10571 14122 10605
rect 14156 10571 14219 10605
rect 14099 10533 14219 10571
rect 14099 10499 14122 10533
rect 14156 10499 14219 10533
rect 14099 10461 14219 10499
rect 14099 10427 14122 10461
rect 14156 10427 14219 10461
rect 14099 10389 14219 10427
rect 14099 10355 14122 10389
rect 14156 10355 14219 10389
rect 14099 10317 14219 10355
rect 14099 10283 14122 10317
rect 14156 10283 14219 10317
rect 14099 10245 14219 10283
rect 14099 10211 14122 10245
rect 14156 10211 14219 10245
rect 757 10146 807 10180
rect 841 10146 877 10180
rect 757 10108 877 10146
rect 757 10074 807 10108
rect 841 10074 877 10108
rect 757 9982 877 10074
rect 14099 10173 14219 10211
rect 14099 10139 14122 10173
rect 14156 10139 14219 10173
rect 14099 10101 14219 10139
rect 14099 10067 14122 10101
rect 14156 10067 14219 10101
tri 877 9982 898 10003 sw
tri 14078 9982 14099 10003 se
rect 14099 9982 14219 10067
rect 757 9963 898 9982
tri 898 9963 917 9982 sw
tri 14059 9963 14078 9982 se
rect 14078 9963 14219 9982
rect 757 9943 14219 9963
tri 757 9942 758 9943 ne
rect 758 9942 14186 9943
rect 245 9879 320 9913
rect 354 9879 430 9913
tri 758 9908 792 9942 ne
rect 792 9908 891 9942
rect 925 9908 963 9942
rect 997 9908 1035 9942
rect 1069 9908 1107 9942
rect 1141 9908 1179 9942
rect 1213 9908 1251 9942
rect 1285 9908 1323 9942
rect 1357 9908 1395 9942
rect 1429 9908 1467 9942
rect 1501 9908 1539 9942
rect 1573 9908 1611 9942
rect 1645 9908 1683 9942
rect 1717 9908 1755 9942
rect 1789 9908 1827 9942
rect 1861 9908 1899 9942
rect 1933 9908 1971 9942
rect 2005 9908 2043 9942
rect 2077 9908 2115 9942
rect 2149 9908 2187 9942
rect 2221 9908 2259 9942
rect 2293 9908 2331 9942
rect 2365 9908 2403 9942
rect 2437 9908 2475 9942
rect 2509 9908 2547 9942
rect 2581 9908 2619 9942
rect 2653 9908 2691 9942
rect 2725 9908 2763 9942
rect 2797 9908 2835 9942
rect 2869 9908 2907 9942
rect 2941 9908 2979 9942
rect 3013 9908 3051 9942
rect 3085 9908 3123 9942
rect 3157 9908 3195 9942
rect 3229 9908 3267 9942
rect 3301 9908 3339 9942
rect 3373 9908 3411 9942
rect 3445 9908 3483 9942
rect 3517 9908 3555 9942
rect 3589 9908 3627 9942
rect 3661 9908 3699 9942
rect 3733 9908 3771 9942
rect 3805 9908 3843 9942
rect 3877 9908 3915 9942
rect 3949 9908 3987 9942
rect 4021 9908 4059 9942
rect 4093 9908 4131 9942
rect 4165 9908 4203 9942
rect 4237 9908 4275 9942
rect 4309 9908 4347 9942
rect 4381 9908 4419 9942
rect 4453 9908 4491 9942
rect 4525 9908 4563 9942
rect 4597 9908 4635 9942
rect 4669 9908 4707 9942
rect 4741 9908 4779 9942
rect 4813 9908 4851 9942
rect 4885 9908 4923 9942
rect 4957 9908 4995 9942
rect 5029 9908 5067 9942
rect 5101 9908 5139 9942
rect 5173 9908 5211 9942
rect 5245 9908 5283 9942
rect 5317 9908 5355 9942
rect 5389 9908 5427 9942
rect 5461 9908 5499 9942
rect 5533 9908 5571 9942
rect 5605 9908 5643 9942
rect 5677 9908 5715 9942
rect 5749 9908 5787 9942
rect 5821 9908 5859 9942
rect 5893 9908 5931 9942
rect 5965 9908 6003 9942
rect 6037 9908 6075 9942
rect 6109 9908 6147 9942
rect 6181 9908 6219 9942
rect 6253 9908 6291 9942
rect 6325 9908 6363 9942
rect 6397 9908 6435 9942
rect 6469 9908 6507 9942
rect 6541 9908 6579 9942
rect 6613 9908 6651 9942
rect 6685 9908 6723 9942
rect 6757 9908 6795 9942
rect 6829 9908 6867 9942
rect 6901 9908 6939 9942
rect 6973 9908 7011 9942
rect 7045 9908 7083 9942
rect 7117 9908 7155 9942
rect 7189 9908 7227 9942
rect 7261 9908 7299 9942
rect 7333 9908 7371 9942
rect 7405 9908 7443 9942
rect 7477 9908 7515 9942
rect 7549 9908 7587 9942
rect 7621 9908 7659 9942
rect 7693 9908 7731 9942
rect 7765 9908 7803 9942
rect 7837 9908 7875 9942
rect 7909 9908 7947 9942
rect 7981 9908 8019 9942
rect 8053 9908 8091 9942
rect 8125 9908 8163 9942
rect 8197 9908 8235 9942
rect 8269 9908 8307 9942
rect 8341 9908 8379 9942
rect 8413 9908 8451 9942
rect 8485 9908 8523 9942
rect 8557 9908 8595 9942
rect 8629 9908 8667 9942
rect 8701 9908 8739 9942
rect 8773 9908 8811 9942
rect 8845 9908 8883 9942
rect 8917 9908 8955 9942
rect 8989 9908 9027 9942
rect 9061 9908 9099 9942
rect 9133 9908 9171 9942
rect 9205 9908 9243 9942
rect 9277 9908 9315 9942
rect 9349 9908 9387 9942
rect 9421 9908 9459 9942
rect 9493 9908 9531 9942
rect 9565 9908 9603 9942
rect 9637 9908 9675 9942
rect 9709 9908 9747 9942
rect 9781 9908 9819 9942
rect 9853 9908 9891 9942
rect 9925 9908 9963 9942
rect 9997 9908 10035 9942
rect 10069 9908 10107 9942
rect 10141 9908 10179 9942
rect 10213 9908 10251 9942
rect 10285 9908 10323 9942
rect 10357 9908 10395 9942
rect 10429 9908 10467 9942
rect 10501 9908 10539 9942
rect 10573 9908 10611 9942
rect 10645 9908 10683 9942
rect 10717 9908 10755 9942
rect 10789 9908 10827 9942
rect 10861 9908 10899 9942
rect 10933 9908 10971 9942
rect 11005 9908 11043 9942
rect 11077 9908 11115 9942
rect 11149 9908 11187 9942
rect 11221 9908 11259 9942
rect 11293 9908 11331 9942
rect 11365 9908 11403 9942
rect 11437 9908 11475 9942
rect 11509 9908 11547 9942
rect 11581 9908 11619 9942
rect 11653 9908 11691 9942
rect 11725 9908 11763 9942
rect 11797 9908 11835 9942
rect 11869 9908 11907 9942
rect 11941 9908 11979 9942
rect 12013 9908 12051 9942
rect 12085 9908 12123 9942
rect 12157 9908 12195 9942
rect 12229 9908 12267 9942
rect 12301 9908 12339 9942
rect 12373 9908 12411 9942
rect 12445 9908 12483 9942
rect 12517 9908 12555 9942
rect 12589 9908 12627 9942
rect 12661 9908 12699 9942
rect 12733 9908 12771 9942
rect 12805 9908 12843 9942
rect 12877 9908 12915 9942
rect 12949 9908 12987 9942
rect 13021 9908 13059 9942
rect 13093 9908 13131 9942
rect 13165 9908 13203 9942
rect 13237 9908 13275 9942
rect 13309 9908 13347 9942
rect 13381 9908 13419 9942
rect 13453 9908 13491 9942
rect 13525 9908 13563 9942
rect 13597 9908 13635 9942
rect 13669 9908 13707 9942
rect 13741 9908 13779 9942
rect 13813 9908 13851 9942
rect 13885 9908 13923 9942
rect 13957 9908 13995 9942
rect 14029 9910 14186 9942
tri 14186 9910 14219 9943 nw
rect 14539 35940 14614 35974
rect 14648 35940 14724 35974
rect 14539 35902 14724 35940
rect 14539 35868 14614 35902
rect 14648 35868 14724 35902
rect 14539 35830 14724 35868
rect 14539 35796 14614 35830
rect 14648 35796 14724 35830
rect 14539 35758 14724 35796
rect 14539 35724 14614 35758
rect 14648 35724 14724 35758
rect 14539 35686 14724 35724
rect 14539 35652 14614 35686
rect 14648 35652 14724 35686
rect 14539 35614 14724 35652
rect 14539 35580 14614 35614
rect 14648 35580 14724 35614
rect 14539 35542 14724 35580
rect 14539 35508 14614 35542
rect 14648 35508 14724 35542
rect 14539 35470 14724 35508
rect 14539 35436 14614 35470
rect 14648 35436 14724 35470
rect 14539 35398 14724 35436
rect 14539 35364 14614 35398
rect 14648 35364 14724 35398
rect 14539 35326 14724 35364
rect 14539 35292 14614 35326
rect 14648 35292 14724 35326
rect 14539 35254 14724 35292
rect 14539 35220 14614 35254
rect 14648 35220 14724 35254
rect 14539 35182 14724 35220
rect 14539 35148 14614 35182
rect 14648 35148 14724 35182
rect 14539 35110 14724 35148
rect 14539 35076 14614 35110
rect 14648 35076 14724 35110
rect 14539 35038 14724 35076
rect 14539 35004 14614 35038
rect 14648 35004 14724 35038
rect 14539 34966 14724 35004
rect 14539 34932 14614 34966
rect 14648 34932 14724 34966
rect 14539 34894 14724 34932
rect 14539 34860 14614 34894
rect 14648 34860 14724 34894
rect 14539 34822 14724 34860
rect 14539 34788 14614 34822
rect 14648 34788 14724 34822
rect 14539 34750 14724 34788
rect 14539 34716 14614 34750
rect 14648 34716 14724 34750
rect 14539 34678 14724 34716
rect 14539 34644 14614 34678
rect 14648 34644 14724 34678
rect 14539 34606 14724 34644
rect 14539 34572 14614 34606
rect 14648 34572 14724 34606
rect 14539 34534 14724 34572
rect 14539 34500 14614 34534
rect 14648 34500 14724 34534
rect 14539 34462 14724 34500
rect 14539 34428 14614 34462
rect 14648 34428 14724 34462
rect 14539 34390 14724 34428
rect 14539 34356 14614 34390
rect 14648 34356 14724 34390
rect 14539 34318 14724 34356
rect 14539 34284 14614 34318
rect 14648 34284 14724 34318
rect 14539 34246 14724 34284
rect 14539 34212 14614 34246
rect 14648 34212 14724 34246
rect 14539 34174 14724 34212
rect 14539 34140 14614 34174
rect 14648 34140 14724 34174
rect 14539 34102 14724 34140
rect 14539 34068 14614 34102
rect 14648 34068 14724 34102
rect 14539 34030 14724 34068
rect 14539 33996 14614 34030
rect 14648 33996 14724 34030
rect 14539 33958 14724 33996
rect 14539 33924 14614 33958
rect 14648 33924 14724 33958
rect 14539 33886 14724 33924
rect 14539 33852 14614 33886
rect 14648 33852 14724 33886
rect 14539 33814 14724 33852
rect 14539 33780 14614 33814
rect 14648 33780 14724 33814
rect 14539 33742 14724 33780
rect 14539 33708 14614 33742
rect 14648 33708 14724 33742
rect 14539 33670 14724 33708
rect 14539 33636 14614 33670
rect 14648 33636 14724 33670
rect 14539 33598 14724 33636
rect 14539 33564 14614 33598
rect 14648 33564 14724 33598
rect 14539 33526 14724 33564
rect 14539 33492 14614 33526
rect 14648 33492 14724 33526
rect 14539 33454 14724 33492
rect 14539 33420 14614 33454
rect 14648 33420 14724 33454
rect 14539 33382 14724 33420
rect 14539 33348 14614 33382
rect 14648 33348 14724 33382
rect 14539 33310 14724 33348
rect 14539 33276 14614 33310
rect 14648 33276 14724 33310
rect 14539 33238 14724 33276
rect 14539 33204 14614 33238
rect 14648 33204 14724 33238
rect 14539 33166 14724 33204
rect 14539 33132 14614 33166
rect 14648 33132 14724 33166
rect 14539 33094 14724 33132
rect 14539 33060 14614 33094
rect 14648 33060 14724 33094
rect 14539 33022 14724 33060
rect 14539 32988 14614 33022
rect 14648 32988 14724 33022
rect 14539 32950 14724 32988
rect 14539 32916 14614 32950
rect 14648 32916 14724 32950
rect 14539 32878 14724 32916
rect 14539 32844 14614 32878
rect 14648 32844 14724 32878
rect 14539 32806 14724 32844
rect 14539 32772 14614 32806
rect 14648 32772 14724 32806
rect 14539 32734 14724 32772
rect 14539 32700 14614 32734
rect 14648 32700 14724 32734
rect 14539 32662 14724 32700
rect 14539 32628 14614 32662
rect 14648 32628 14724 32662
rect 14539 32590 14724 32628
rect 14539 32556 14614 32590
rect 14648 32556 14724 32590
rect 14539 32518 14724 32556
rect 14539 32484 14614 32518
rect 14648 32484 14724 32518
rect 14539 32446 14724 32484
rect 14539 32412 14614 32446
rect 14648 32412 14724 32446
rect 14539 32374 14724 32412
rect 14539 32340 14614 32374
rect 14648 32340 14724 32374
rect 14539 32302 14724 32340
rect 14539 32268 14614 32302
rect 14648 32268 14724 32302
rect 14539 32230 14724 32268
rect 14539 32196 14614 32230
rect 14648 32196 14724 32230
rect 14539 32158 14724 32196
rect 14539 32124 14614 32158
rect 14648 32124 14724 32158
rect 14539 32086 14724 32124
rect 14539 32052 14614 32086
rect 14648 32052 14724 32086
rect 14539 32014 14724 32052
rect 14539 31980 14614 32014
rect 14648 31980 14724 32014
rect 14539 31942 14724 31980
rect 14539 31908 14614 31942
rect 14648 31908 14724 31942
rect 14539 31870 14724 31908
rect 14539 31836 14614 31870
rect 14648 31836 14724 31870
rect 14539 31798 14724 31836
rect 14539 31764 14614 31798
rect 14648 31764 14724 31798
rect 14539 31726 14724 31764
rect 14539 31692 14614 31726
rect 14648 31692 14724 31726
rect 14539 31654 14724 31692
rect 14539 31620 14614 31654
rect 14648 31620 14724 31654
rect 14539 31582 14724 31620
rect 14539 31548 14614 31582
rect 14648 31548 14724 31582
rect 14539 31510 14724 31548
rect 14539 31476 14614 31510
rect 14648 31476 14724 31510
rect 14539 31438 14724 31476
rect 14539 31404 14614 31438
rect 14648 31404 14724 31438
rect 14539 31366 14724 31404
rect 14539 31332 14614 31366
rect 14648 31332 14724 31366
rect 14539 31294 14724 31332
rect 14539 31260 14614 31294
rect 14648 31260 14724 31294
rect 14539 31222 14724 31260
rect 14539 31188 14614 31222
rect 14648 31188 14724 31222
rect 14539 31150 14724 31188
rect 14539 31116 14614 31150
rect 14648 31116 14724 31150
rect 14539 31078 14724 31116
rect 14539 31044 14614 31078
rect 14648 31044 14724 31078
rect 14539 31006 14724 31044
rect 14539 30972 14614 31006
rect 14648 30972 14724 31006
rect 14539 30934 14724 30972
rect 14539 30900 14614 30934
rect 14648 30900 14724 30934
rect 14539 30862 14724 30900
rect 14539 30828 14614 30862
rect 14648 30828 14724 30862
rect 14539 30790 14724 30828
rect 14539 30756 14614 30790
rect 14648 30756 14724 30790
rect 14539 30718 14724 30756
rect 14539 30684 14614 30718
rect 14648 30684 14724 30718
rect 14539 30646 14724 30684
rect 14539 30612 14614 30646
rect 14648 30612 14724 30646
rect 14539 30574 14724 30612
rect 14539 30540 14614 30574
rect 14648 30540 14724 30574
rect 14539 30502 14724 30540
rect 14539 30468 14614 30502
rect 14648 30468 14724 30502
rect 14539 30430 14724 30468
rect 14539 30396 14614 30430
rect 14648 30396 14724 30430
rect 14539 30358 14724 30396
rect 14539 30324 14614 30358
rect 14648 30324 14724 30358
rect 14539 30286 14724 30324
rect 14539 30252 14614 30286
rect 14648 30252 14724 30286
rect 14539 30214 14724 30252
rect 14539 30180 14614 30214
rect 14648 30180 14724 30214
rect 14539 30142 14724 30180
rect 14539 30108 14614 30142
rect 14648 30108 14724 30142
rect 14539 30070 14724 30108
rect 14539 30036 14614 30070
rect 14648 30036 14724 30070
rect 14539 29998 14724 30036
rect 14539 29964 14614 29998
rect 14648 29964 14724 29998
rect 14539 29926 14724 29964
rect 14539 29892 14614 29926
rect 14648 29892 14724 29926
rect 14539 29854 14724 29892
rect 14539 29820 14614 29854
rect 14648 29820 14724 29854
rect 14539 29782 14724 29820
rect 14539 29748 14614 29782
rect 14648 29748 14724 29782
rect 14539 29710 14724 29748
rect 14539 29676 14614 29710
rect 14648 29676 14724 29710
rect 14539 29638 14724 29676
rect 14539 29604 14614 29638
rect 14648 29604 14724 29638
rect 14539 29566 14724 29604
rect 14539 29532 14614 29566
rect 14648 29532 14724 29566
rect 14539 29494 14724 29532
rect 14539 29460 14614 29494
rect 14648 29460 14724 29494
rect 14539 29422 14724 29460
rect 14539 29388 14614 29422
rect 14648 29388 14724 29422
rect 14539 29350 14724 29388
rect 14539 29316 14614 29350
rect 14648 29316 14724 29350
rect 14539 29278 14724 29316
rect 14539 29244 14614 29278
rect 14648 29244 14724 29278
rect 14539 29206 14724 29244
rect 14539 29172 14614 29206
rect 14648 29172 14724 29206
rect 14539 29134 14724 29172
rect 14539 29100 14614 29134
rect 14648 29100 14724 29134
rect 14539 29062 14724 29100
rect 14539 29028 14614 29062
rect 14648 29028 14724 29062
rect 14539 28990 14724 29028
rect 14539 28956 14614 28990
rect 14648 28956 14724 28990
rect 14539 28918 14724 28956
rect 14539 28884 14614 28918
rect 14648 28884 14724 28918
rect 14539 28846 14724 28884
rect 14539 28812 14614 28846
rect 14648 28812 14724 28846
rect 14539 28774 14724 28812
rect 14539 28740 14614 28774
rect 14648 28740 14724 28774
rect 14539 28702 14724 28740
rect 14539 28668 14614 28702
rect 14648 28668 14724 28702
rect 14539 28630 14724 28668
rect 14539 28596 14614 28630
rect 14648 28596 14724 28630
rect 14539 28558 14724 28596
rect 14539 28524 14614 28558
rect 14648 28524 14724 28558
rect 14539 28486 14724 28524
rect 14539 28452 14614 28486
rect 14648 28452 14724 28486
rect 14539 28414 14724 28452
rect 14539 28380 14614 28414
rect 14648 28380 14724 28414
rect 14539 28342 14724 28380
rect 14539 28308 14614 28342
rect 14648 28308 14724 28342
rect 14539 28270 14724 28308
rect 14539 28236 14614 28270
rect 14648 28236 14724 28270
rect 14539 28198 14724 28236
rect 14539 28164 14614 28198
rect 14648 28164 14724 28198
rect 14539 28126 14724 28164
rect 14539 28092 14614 28126
rect 14648 28092 14724 28126
rect 14539 28054 14724 28092
rect 14539 28020 14614 28054
rect 14648 28020 14724 28054
rect 14539 27982 14724 28020
rect 14539 27948 14614 27982
rect 14648 27948 14724 27982
rect 14539 27910 14724 27948
rect 14539 27876 14614 27910
rect 14648 27876 14724 27910
rect 14539 27838 14724 27876
rect 14539 27804 14614 27838
rect 14648 27804 14724 27838
rect 14539 27766 14724 27804
rect 14539 27732 14614 27766
rect 14648 27732 14724 27766
rect 14539 27694 14724 27732
rect 14539 27660 14614 27694
rect 14648 27660 14724 27694
rect 14539 27622 14724 27660
rect 14539 27588 14614 27622
rect 14648 27588 14724 27622
rect 14539 27550 14724 27588
rect 14539 27516 14614 27550
rect 14648 27516 14724 27550
rect 14539 27478 14724 27516
rect 14539 27444 14614 27478
rect 14648 27444 14724 27478
rect 14539 27406 14724 27444
rect 14539 27372 14614 27406
rect 14648 27372 14724 27406
rect 14539 27334 14724 27372
rect 14539 27300 14614 27334
rect 14648 27300 14724 27334
rect 14539 27262 14724 27300
rect 14539 27228 14614 27262
rect 14648 27228 14724 27262
rect 14539 27190 14724 27228
rect 14539 27156 14614 27190
rect 14648 27156 14724 27190
rect 14539 27118 14724 27156
rect 14539 27084 14614 27118
rect 14648 27084 14724 27118
rect 14539 27046 14724 27084
rect 14539 27012 14614 27046
rect 14648 27012 14724 27046
rect 14539 26974 14724 27012
rect 14539 26940 14614 26974
rect 14648 26940 14724 26974
rect 14539 26902 14724 26940
rect 14539 26868 14614 26902
rect 14648 26868 14724 26902
rect 14539 26830 14724 26868
rect 14539 26796 14614 26830
rect 14648 26796 14724 26830
rect 14539 26758 14724 26796
rect 14539 26724 14614 26758
rect 14648 26724 14724 26758
rect 14539 26686 14724 26724
rect 14539 26652 14614 26686
rect 14648 26652 14724 26686
rect 14539 26614 14724 26652
rect 14539 26580 14614 26614
rect 14648 26580 14724 26614
rect 14539 26542 14724 26580
rect 14539 26508 14614 26542
rect 14648 26508 14724 26542
rect 14539 26470 14724 26508
rect 14539 26436 14614 26470
rect 14648 26436 14724 26470
rect 14539 26398 14724 26436
rect 14539 26364 14614 26398
rect 14648 26364 14724 26398
rect 14539 26326 14724 26364
rect 14539 26292 14614 26326
rect 14648 26292 14724 26326
rect 14539 26254 14724 26292
rect 14539 26220 14614 26254
rect 14648 26220 14724 26254
rect 14539 26182 14724 26220
rect 14539 26148 14614 26182
rect 14648 26148 14724 26182
rect 14539 26110 14724 26148
rect 14539 26076 14614 26110
rect 14648 26076 14724 26110
rect 14539 26038 14724 26076
rect 14539 26004 14614 26038
rect 14648 26004 14724 26038
rect 14539 25966 14724 26004
rect 14539 25932 14614 25966
rect 14648 25932 14724 25966
rect 14539 25894 14724 25932
rect 14539 25860 14614 25894
rect 14648 25860 14724 25894
rect 14539 25822 14724 25860
rect 14539 25788 14614 25822
rect 14648 25788 14724 25822
rect 14539 25750 14724 25788
rect 14539 25716 14614 25750
rect 14648 25716 14724 25750
rect 14539 25678 14724 25716
rect 14539 25644 14614 25678
rect 14648 25644 14724 25678
rect 14539 25606 14724 25644
rect 14539 25572 14614 25606
rect 14648 25572 14724 25606
rect 14539 25534 14724 25572
rect 14539 25500 14614 25534
rect 14648 25500 14724 25534
rect 14539 25462 14724 25500
rect 14539 25428 14614 25462
rect 14648 25428 14724 25462
rect 14539 25390 14724 25428
rect 14539 25356 14614 25390
rect 14648 25356 14724 25390
rect 14539 25318 14724 25356
rect 14539 25284 14614 25318
rect 14648 25284 14724 25318
rect 14539 25246 14724 25284
rect 14539 25212 14614 25246
rect 14648 25212 14724 25246
rect 14539 25174 14724 25212
rect 14539 25140 14614 25174
rect 14648 25140 14724 25174
rect 14539 25102 14724 25140
rect 14539 25068 14614 25102
rect 14648 25068 14724 25102
rect 14539 25030 14724 25068
rect 14539 24996 14614 25030
rect 14648 24996 14724 25030
rect 14539 24958 14724 24996
rect 14539 24924 14614 24958
rect 14648 24924 14724 24958
rect 14539 24886 14724 24924
rect 14539 24852 14614 24886
rect 14648 24852 14724 24886
rect 14539 24814 14724 24852
rect 14539 24780 14614 24814
rect 14648 24780 14724 24814
rect 14539 24742 14724 24780
rect 14539 24708 14614 24742
rect 14648 24708 14724 24742
rect 14539 24670 14724 24708
rect 14539 24636 14614 24670
rect 14648 24636 14724 24670
rect 14539 24598 14724 24636
rect 14539 24564 14614 24598
rect 14648 24564 14724 24598
rect 14539 24526 14724 24564
rect 14539 24492 14614 24526
rect 14648 24492 14724 24526
rect 14539 24454 14724 24492
rect 14539 24420 14614 24454
rect 14648 24420 14724 24454
rect 14539 24382 14724 24420
rect 14539 24348 14614 24382
rect 14648 24348 14724 24382
rect 14539 24310 14724 24348
rect 14539 24276 14614 24310
rect 14648 24276 14724 24310
rect 14539 24238 14724 24276
rect 14539 24204 14614 24238
rect 14648 24204 14724 24238
rect 14539 24166 14724 24204
rect 14539 24132 14614 24166
rect 14648 24132 14724 24166
rect 14539 24094 14724 24132
rect 14539 24060 14614 24094
rect 14648 24060 14724 24094
rect 14539 24022 14724 24060
rect 14539 23988 14614 24022
rect 14648 23988 14724 24022
rect 14539 23950 14724 23988
rect 14539 23916 14614 23950
rect 14648 23916 14724 23950
rect 14539 23878 14724 23916
rect 14539 23844 14614 23878
rect 14648 23844 14724 23878
rect 14539 23806 14724 23844
rect 14539 23772 14614 23806
rect 14648 23772 14724 23806
rect 14539 23734 14724 23772
rect 14539 23700 14614 23734
rect 14648 23700 14724 23734
rect 14539 23662 14724 23700
rect 14539 23628 14614 23662
rect 14648 23628 14724 23662
rect 14539 23590 14724 23628
rect 14539 23556 14614 23590
rect 14648 23556 14724 23590
rect 14539 23518 14724 23556
rect 14539 23484 14614 23518
rect 14648 23484 14724 23518
rect 14539 23446 14724 23484
rect 14539 23412 14614 23446
rect 14648 23412 14724 23446
rect 14539 23374 14724 23412
rect 14539 23340 14614 23374
rect 14648 23340 14724 23374
rect 14539 23302 14724 23340
rect 14539 23268 14614 23302
rect 14648 23268 14724 23302
rect 14539 23230 14724 23268
rect 14539 23196 14614 23230
rect 14648 23196 14724 23230
rect 14539 23158 14724 23196
rect 14539 23124 14614 23158
rect 14648 23124 14724 23158
rect 14539 23086 14724 23124
rect 14539 23052 14614 23086
rect 14648 23052 14724 23086
rect 14539 23014 14724 23052
rect 14539 22980 14614 23014
rect 14648 22980 14724 23014
rect 14539 22942 14724 22980
rect 14539 22908 14614 22942
rect 14648 22908 14724 22942
rect 14539 22870 14724 22908
rect 14539 22836 14614 22870
rect 14648 22836 14724 22870
rect 14539 22798 14724 22836
rect 14539 22764 14614 22798
rect 14648 22764 14724 22798
rect 14539 22726 14724 22764
rect 14539 22692 14614 22726
rect 14648 22692 14724 22726
rect 14539 22654 14724 22692
rect 14539 22620 14614 22654
rect 14648 22620 14724 22654
rect 14539 22582 14724 22620
rect 14539 22548 14614 22582
rect 14648 22548 14724 22582
rect 14539 22510 14724 22548
rect 14539 22476 14614 22510
rect 14648 22476 14724 22510
rect 14539 22438 14724 22476
rect 14539 22404 14614 22438
rect 14648 22404 14724 22438
rect 14539 22366 14724 22404
rect 14539 22332 14614 22366
rect 14648 22332 14724 22366
rect 14539 22294 14724 22332
rect 14539 22260 14614 22294
rect 14648 22260 14724 22294
rect 14539 22222 14724 22260
rect 14539 22188 14614 22222
rect 14648 22188 14724 22222
rect 14539 22150 14724 22188
rect 14539 22116 14614 22150
rect 14648 22116 14724 22150
rect 14539 22078 14724 22116
rect 14539 22044 14614 22078
rect 14648 22044 14724 22078
rect 14539 22006 14724 22044
rect 14539 21972 14614 22006
rect 14648 21972 14724 22006
rect 14539 21934 14724 21972
rect 14539 21900 14614 21934
rect 14648 21900 14724 21934
rect 14539 21862 14724 21900
rect 14539 21828 14614 21862
rect 14648 21828 14724 21862
rect 14539 21790 14724 21828
rect 14539 21756 14614 21790
rect 14648 21756 14724 21790
rect 14539 21718 14724 21756
rect 14539 21684 14614 21718
rect 14648 21684 14724 21718
rect 14539 21646 14724 21684
rect 14539 21612 14614 21646
rect 14648 21612 14724 21646
rect 14539 21574 14724 21612
rect 14539 21540 14614 21574
rect 14648 21540 14724 21574
rect 14539 21502 14724 21540
rect 14539 21468 14614 21502
rect 14648 21468 14724 21502
rect 14539 21430 14724 21468
rect 14539 21396 14614 21430
rect 14648 21396 14724 21430
rect 14539 21358 14724 21396
rect 14539 21324 14614 21358
rect 14648 21324 14724 21358
rect 14539 21286 14724 21324
rect 14539 21252 14614 21286
rect 14648 21252 14724 21286
rect 14539 21214 14724 21252
rect 14539 21180 14614 21214
rect 14648 21180 14724 21214
rect 14539 21142 14724 21180
rect 14539 21108 14614 21142
rect 14648 21108 14724 21142
rect 14539 21070 14724 21108
rect 14539 21036 14614 21070
rect 14648 21036 14724 21070
rect 14539 20998 14724 21036
rect 14539 20964 14614 20998
rect 14648 20964 14724 20998
rect 14539 20926 14724 20964
rect 14539 20892 14614 20926
rect 14648 20892 14724 20926
rect 14539 20854 14724 20892
rect 14539 20820 14614 20854
rect 14648 20820 14724 20854
rect 14539 20782 14724 20820
rect 14539 20748 14614 20782
rect 14648 20748 14724 20782
rect 14539 20710 14724 20748
rect 14539 20676 14614 20710
rect 14648 20676 14724 20710
rect 14539 20638 14724 20676
rect 14539 20604 14614 20638
rect 14648 20604 14724 20638
rect 14539 20566 14724 20604
rect 14539 20532 14614 20566
rect 14648 20532 14724 20566
rect 14539 20494 14724 20532
rect 14539 20460 14614 20494
rect 14648 20460 14724 20494
rect 14539 20422 14724 20460
rect 14539 20388 14614 20422
rect 14648 20388 14724 20422
rect 14539 20350 14724 20388
rect 14539 20316 14614 20350
rect 14648 20316 14724 20350
rect 14539 20278 14724 20316
rect 14539 20244 14614 20278
rect 14648 20244 14724 20278
rect 14539 20206 14724 20244
rect 14539 20172 14614 20206
rect 14648 20172 14724 20206
rect 14539 20134 14724 20172
rect 14539 20100 14614 20134
rect 14648 20100 14724 20134
rect 14539 20062 14724 20100
rect 14539 20028 14614 20062
rect 14648 20028 14724 20062
rect 14539 19990 14724 20028
rect 14539 19956 14614 19990
rect 14648 19956 14724 19990
rect 14539 19918 14724 19956
rect 14539 19884 14614 19918
rect 14648 19884 14724 19918
rect 14539 19846 14724 19884
rect 14539 19812 14614 19846
rect 14648 19812 14724 19846
rect 14539 19774 14724 19812
rect 14539 19740 14614 19774
rect 14648 19740 14724 19774
rect 14539 19702 14724 19740
rect 14539 19668 14614 19702
rect 14648 19668 14724 19702
rect 14539 19630 14724 19668
rect 14539 19596 14614 19630
rect 14648 19596 14724 19630
rect 14539 19558 14724 19596
rect 14539 19524 14614 19558
rect 14648 19524 14724 19558
rect 14539 19486 14724 19524
rect 14539 19452 14614 19486
rect 14648 19452 14724 19486
rect 14539 19414 14724 19452
rect 14539 19380 14614 19414
rect 14648 19380 14724 19414
rect 14539 19342 14724 19380
rect 14539 19308 14614 19342
rect 14648 19308 14724 19342
rect 14539 19270 14724 19308
rect 14539 19236 14614 19270
rect 14648 19236 14724 19270
rect 14539 19198 14724 19236
rect 14539 19164 14614 19198
rect 14648 19164 14724 19198
rect 14539 19126 14724 19164
rect 14539 19092 14614 19126
rect 14648 19092 14724 19126
rect 14539 19054 14724 19092
rect 14539 19020 14614 19054
rect 14648 19020 14724 19054
rect 14539 18982 14724 19020
rect 14539 18948 14614 18982
rect 14648 18948 14724 18982
rect 14539 18910 14724 18948
rect 14539 18876 14614 18910
rect 14648 18876 14724 18910
rect 14539 18838 14724 18876
rect 14539 18804 14614 18838
rect 14648 18804 14724 18838
rect 14539 18766 14724 18804
rect 14539 18732 14614 18766
rect 14648 18732 14724 18766
rect 14539 18694 14724 18732
rect 14539 18660 14614 18694
rect 14648 18660 14724 18694
rect 14539 18622 14724 18660
rect 14539 18588 14614 18622
rect 14648 18588 14724 18622
rect 14539 18550 14724 18588
rect 14539 18516 14614 18550
rect 14648 18516 14724 18550
rect 14539 18478 14724 18516
rect 14539 18444 14614 18478
rect 14648 18444 14724 18478
rect 14539 18406 14724 18444
rect 14539 18372 14614 18406
rect 14648 18372 14724 18406
rect 14539 18334 14724 18372
rect 14539 18300 14614 18334
rect 14648 18300 14724 18334
rect 14539 18262 14724 18300
rect 14539 18228 14614 18262
rect 14648 18228 14724 18262
rect 14539 18190 14724 18228
rect 14539 18156 14614 18190
rect 14648 18156 14724 18190
rect 14539 18118 14724 18156
rect 14539 18084 14614 18118
rect 14648 18084 14724 18118
rect 14539 18046 14724 18084
rect 14539 18012 14614 18046
rect 14648 18012 14724 18046
rect 14539 17974 14724 18012
rect 14539 17940 14614 17974
rect 14648 17940 14724 17974
rect 14539 17902 14724 17940
rect 14539 17868 14614 17902
rect 14648 17868 14724 17902
rect 14539 17830 14724 17868
rect 14539 17796 14614 17830
rect 14648 17796 14724 17830
rect 14539 17758 14724 17796
rect 14539 17724 14614 17758
rect 14648 17724 14724 17758
rect 14539 17686 14724 17724
rect 14539 17652 14614 17686
rect 14648 17652 14724 17686
rect 14539 17614 14724 17652
rect 14539 17580 14614 17614
rect 14648 17580 14724 17614
rect 14539 17542 14724 17580
rect 14539 17508 14614 17542
rect 14648 17508 14724 17542
rect 14539 17470 14724 17508
rect 14539 17436 14614 17470
rect 14648 17436 14724 17470
rect 14539 17398 14724 17436
rect 14539 17364 14614 17398
rect 14648 17364 14724 17398
rect 14539 17326 14724 17364
rect 14539 17292 14614 17326
rect 14648 17292 14724 17326
rect 14539 17254 14724 17292
rect 14539 17220 14614 17254
rect 14648 17220 14724 17254
rect 14539 17182 14724 17220
rect 14539 17148 14614 17182
rect 14648 17148 14724 17182
rect 14539 17110 14724 17148
rect 14539 17076 14614 17110
rect 14648 17076 14724 17110
rect 14539 17038 14724 17076
rect 14539 17004 14614 17038
rect 14648 17004 14724 17038
rect 14539 16966 14724 17004
rect 14539 16932 14614 16966
rect 14648 16932 14724 16966
rect 14539 16894 14724 16932
rect 14539 16860 14614 16894
rect 14648 16860 14724 16894
rect 14539 16822 14724 16860
rect 14539 16788 14614 16822
rect 14648 16788 14724 16822
rect 14539 16750 14724 16788
rect 14539 16716 14614 16750
rect 14648 16716 14724 16750
rect 14539 16678 14724 16716
rect 14539 16644 14614 16678
rect 14648 16644 14724 16678
rect 14539 16606 14724 16644
rect 14539 16572 14614 16606
rect 14648 16572 14724 16606
rect 14539 16534 14724 16572
rect 14539 16500 14614 16534
rect 14648 16500 14724 16534
rect 14539 16462 14724 16500
rect 14539 16428 14614 16462
rect 14648 16428 14724 16462
rect 14539 16390 14724 16428
rect 14539 16356 14614 16390
rect 14648 16356 14724 16390
rect 14539 16318 14724 16356
rect 14539 16284 14614 16318
rect 14648 16284 14724 16318
rect 14539 16246 14724 16284
rect 14539 16212 14614 16246
rect 14648 16212 14724 16246
rect 14539 16174 14724 16212
rect 14539 16140 14614 16174
rect 14648 16140 14724 16174
rect 14539 16102 14724 16140
rect 14539 16068 14614 16102
rect 14648 16068 14724 16102
rect 14539 16030 14724 16068
rect 14539 15996 14614 16030
rect 14648 15996 14724 16030
rect 14539 15958 14724 15996
rect 14539 15924 14614 15958
rect 14648 15924 14724 15958
rect 14539 15886 14724 15924
rect 14539 15852 14614 15886
rect 14648 15852 14724 15886
rect 14539 15814 14724 15852
rect 14539 15780 14614 15814
rect 14648 15780 14724 15814
rect 14539 15742 14724 15780
rect 14539 15708 14614 15742
rect 14648 15708 14724 15742
rect 14539 15670 14724 15708
rect 14539 15636 14614 15670
rect 14648 15636 14724 15670
rect 14539 15598 14724 15636
rect 14539 15564 14614 15598
rect 14648 15564 14724 15598
rect 14539 15526 14724 15564
rect 14539 15492 14614 15526
rect 14648 15492 14724 15526
rect 14539 15454 14724 15492
rect 14539 15420 14614 15454
rect 14648 15420 14724 15454
rect 14539 15382 14724 15420
rect 14539 15348 14614 15382
rect 14648 15348 14724 15382
rect 14539 15310 14724 15348
rect 14539 15276 14614 15310
rect 14648 15276 14724 15310
rect 14539 15238 14724 15276
rect 14539 15204 14614 15238
rect 14648 15204 14724 15238
rect 14539 15166 14724 15204
rect 14539 15132 14614 15166
rect 14648 15132 14724 15166
rect 14539 15094 14724 15132
rect 14539 15060 14614 15094
rect 14648 15060 14724 15094
rect 14539 15022 14724 15060
rect 14539 14988 14614 15022
rect 14648 14988 14724 15022
rect 14539 14950 14724 14988
rect 14539 14916 14614 14950
rect 14648 14916 14724 14950
rect 14539 14878 14724 14916
rect 14539 14844 14614 14878
rect 14648 14844 14724 14878
rect 14539 14806 14724 14844
rect 14539 14772 14614 14806
rect 14648 14772 14724 14806
rect 14539 14734 14724 14772
rect 14539 14700 14614 14734
rect 14648 14700 14724 14734
rect 14539 14662 14724 14700
rect 14539 14628 14614 14662
rect 14648 14628 14724 14662
rect 14539 14590 14724 14628
rect 14539 14556 14614 14590
rect 14648 14556 14724 14590
rect 14539 14518 14724 14556
rect 14539 14484 14614 14518
rect 14648 14484 14724 14518
rect 14539 14446 14724 14484
rect 14539 14412 14614 14446
rect 14648 14412 14724 14446
rect 14539 14374 14724 14412
rect 14539 14340 14614 14374
rect 14648 14340 14724 14374
rect 14539 14302 14724 14340
rect 14539 14268 14614 14302
rect 14648 14268 14724 14302
rect 14539 14230 14724 14268
rect 14539 14196 14614 14230
rect 14648 14196 14724 14230
rect 14539 14158 14724 14196
rect 14539 14124 14614 14158
rect 14648 14124 14724 14158
rect 14539 14086 14724 14124
rect 14539 14052 14614 14086
rect 14648 14052 14724 14086
rect 14539 14014 14724 14052
rect 14539 13980 14614 14014
rect 14648 13980 14724 14014
rect 14539 13942 14724 13980
rect 14539 13908 14614 13942
rect 14648 13908 14724 13942
rect 14539 13870 14724 13908
rect 14539 13836 14614 13870
rect 14648 13836 14724 13870
rect 14539 13798 14724 13836
rect 14539 13764 14614 13798
rect 14648 13764 14724 13798
rect 14539 13726 14724 13764
rect 14539 13692 14614 13726
rect 14648 13692 14724 13726
rect 14539 13654 14724 13692
rect 14539 13620 14614 13654
rect 14648 13620 14724 13654
rect 14539 13582 14724 13620
rect 14539 13548 14614 13582
rect 14648 13548 14724 13582
rect 14539 13510 14724 13548
rect 14539 13476 14614 13510
rect 14648 13476 14724 13510
rect 14539 13438 14724 13476
rect 14539 13404 14614 13438
rect 14648 13404 14724 13438
rect 14539 13366 14724 13404
rect 14539 13332 14614 13366
rect 14648 13332 14724 13366
rect 14539 13294 14724 13332
rect 14539 13260 14614 13294
rect 14648 13260 14724 13294
rect 14539 13222 14724 13260
rect 14539 13188 14614 13222
rect 14648 13188 14724 13222
rect 14539 13150 14724 13188
rect 14539 13116 14614 13150
rect 14648 13116 14724 13150
rect 14539 13078 14724 13116
rect 14539 13044 14614 13078
rect 14648 13044 14724 13078
rect 14539 13006 14724 13044
rect 14539 12972 14614 13006
rect 14648 12972 14724 13006
rect 14539 12934 14724 12972
rect 14539 12900 14614 12934
rect 14648 12900 14724 12934
rect 14539 12862 14724 12900
rect 14539 12828 14614 12862
rect 14648 12828 14724 12862
rect 14539 12790 14724 12828
rect 14539 12756 14614 12790
rect 14648 12756 14724 12790
rect 14539 12718 14724 12756
rect 14539 12684 14614 12718
rect 14648 12684 14724 12718
rect 14539 12646 14724 12684
rect 14539 12612 14614 12646
rect 14648 12612 14724 12646
rect 14539 12574 14724 12612
rect 14539 12540 14614 12574
rect 14648 12540 14724 12574
rect 14539 12502 14724 12540
rect 14539 12468 14614 12502
rect 14648 12468 14724 12502
rect 14539 12430 14724 12468
rect 14539 12396 14614 12430
rect 14648 12396 14724 12430
rect 14539 12358 14724 12396
rect 14539 12324 14614 12358
rect 14648 12324 14724 12358
rect 14539 12286 14724 12324
rect 14539 12252 14614 12286
rect 14648 12252 14724 12286
rect 14539 12214 14724 12252
rect 14539 12180 14614 12214
rect 14648 12180 14724 12214
rect 14539 12142 14724 12180
rect 14539 12108 14614 12142
rect 14648 12108 14724 12142
rect 14539 12070 14724 12108
rect 14539 12036 14614 12070
rect 14648 12036 14724 12070
rect 14539 11998 14724 12036
rect 14539 11964 14614 11998
rect 14648 11964 14724 11998
rect 14539 11926 14724 11964
rect 14539 11892 14614 11926
rect 14648 11892 14724 11926
rect 14539 11854 14724 11892
rect 14539 11820 14614 11854
rect 14648 11820 14724 11854
rect 14539 11782 14724 11820
rect 14539 11748 14614 11782
rect 14648 11748 14724 11782
rect 14539 11710 14724 11748
rect 14539 11676 14614 11710
rect 14648 11676 14724 11710
rect 14539 11638 14724 11676
rect 14539 11604 14614 11638
rect 14648 11604 14724 11638
rect 14539 11566 14724 11604
rect 14539 11532 14614 11566
rect 14648 11532 14724 11566
rect 14539 11494 14724 11532
rect 14539 11460 14614 11494
rect 14648 11460 14724 11494
rect 14539 11422 14724 11460
rect 14539 11388 14614 11422
rect 14648 11388 14724 11422
rect 14539 11350 14724 11388
rect 14539 11316 14614 11350
rect 14648 11316 14724 11350
rect 14539 11278 14724 11316
rect 14539 11244 14614 11278
rect 14648 11244 14724 11278
rect 14539 11206 14724 11244
rect 14539 11172 14614 11206
rect 14648 11172 14724 11206
rect 14539 11134 14724 11172
rect 14539 11100 14614 11134
rect 14648 11100 14724 11134
rect 14539 11062 14724 11100
rect 14539 11028 14614 11062
rect 14648 11028 14724 11062
rect 14539 10990 14724 11028
rect 14539 10956 14614 10990
rect 14648 10956 14724 10990
rect 14539 10918 14724 10956
rect 14539 10884 14614 10918
rect 14648 10884 14724 10918
rect 14539 10846 14724 10884
rect 14539 10812 14614 10846
rect 14648 10812 14724 10846
rect 14539 10774 14724 10812
rect 14539 10740 14614 10774
rect 14648 10740 14724 10774
rect 14539 10702 14724 10740
rect 14539 10668 14614 10702
rect 14648 10668 14724 10702
rect 14539 10630 14724 10668
rect 14539 10596 14614 10630
rect 14648 10596 14724 10630
rect 14539 10558 14724 10596
rect 14539 10524 14614 10558
rect 14648 10524 14724 10558
rect 14539 10486 14724 10524
rect 14539 10452 14614 10486
rect 14648 10452 14724 10486
rect 14539 10414 14724 10452
rect 14539 10380 14614 10414
rect 14648 10380 14724 10414
rect 14539 10342 14724 10380
rect 14539 10308 14614 10342
rect 14648 10308 14724 10342
rect 14539 10270 14724 10308
rect 14539 10236 14614 10270
rect 14648 10236 14724 10270
rect 14539 10198 14724 10236
rect 14539 10164 14614 10198
rect 14648 10164 14724 10198
rect 14539 10126 14724 10164
rect 14539 10092 14614 10126
rect 14648 10092 14724 10126
rect 14539 10054 14724 10092
rect 14539 10020 14614 10054
rect 14648 10020 14724 10054
rect 14539 9982 14724 10020
rect 14539 9948 14614 9982
rect 14648 9948 14724 9982
rect 14539 9910 14724 9948
rect 14029 9908 14152 9910
rect 245 9841 430 9879
tri 792 9876 824 9908 ne
rect 824 9876 14152 9908
tri 14152 9876 14186 9910 nw
rect 14539 9876 14614 9910
rect 14648 9876 14724 9910
tri 824 9843 857 9876 ne
rect 857 9843 14119 9876
tri 14119 9843 14152 9876 nw
rect 245 9807 320 9841
rect 354 9807 430 9841
rect 245 9769 430 9807
rect 245 9735 320 9769
rect 354 9735 430 9769
rect 245 9697 430 9735
rect 245 9663 320 9697
rect 354 9663 430 9697
rect 245 9528 430 9663
rect 858 9774 2096 9843
rect 858 9740 883 9774
rect 917 9740 955 9774
rect 989 9740 1027 9774
rect 1061 9740 1099 9774
rect 1133 9740 1171 9774
rect 1205 9740 1243 9774
rect 1277 9740 1315 9774
rect 1349 9740 1387 9774
rect 1421 9740 1459 9774
rect 1493 9740 1531 9774
rect 1565 9740 1603 9774
rect 1637 9740 1675 9774
rect 1709 9740 1747 9774
rect 1781 9740 1819 9774
rect 1853 9740 1891 9774
rect 1925 9740 1963 9774
rect 1997 9740 2035 9774
rect 2069 9740 2096 9774
rect 858 9731 2096 9740
rect 245 9452 720 9528
rect 245 9418 320 9452
rect 354 9418 610 9452
rect 644 9418 720 9452
rect 245 9343 720 9418
rect 858 9295 908 9731
rect 2048 9295 2096 9731
rect 12858 9774 14096 9843
rect 12858 9740 12883 9774
rect 12917 9740 12955 9774
rect 12989 9740 13027 9774
rect 13061 9740 13099 9774
rect 13133 9740 13171 9774
rect 13205 9740 13243 9774
rect 13277 9740 13315 9774
rect 13349 9740 13387 9774
rect 13421 9740 13459 9774
rect 13493 9740 13531 9774
rect 13565 9740 13603 9774
rect 13637 9740 13675 9774
rect 13709 9740 13747 9774
rect 13781 9740 13819 9774
rect 13853 9740 13891 9774
rect 13925 9740 13963 9774
rect 13997 9740 14035 9774
rect 14069 9740 14096 9774
rect 12858 9731 14096 9740
rect 11273 9528 12512 9529
rect 2248 9484 12705 9528
rect 2248 9483 11322 9484
rect 2248 9452 2445 9483
rect 3585 9452 11322 9483
rect 12462 9452 12705 9484
rect 2248 9418 2311 9452
rect 2345 9418 2383 9452
rect 2417 9418 2445 9452
rect 3585 9418 3607 9452
rect 3641 9418 3679 9452
rect 3713 9418 3751 9452
rect 3785 9418 3823 9452
rect 3857 9418 3895 9452
rect 3929 9418 3967 9452
rect 4001 9418 4039 9452
rect 4073 9418 4111 9452
rect 4145 9418 4183 9452
rect 4217 9418 4255 9452
rect 4289 9418 4327 9452
rect 4361 9418 4399 9452
rect 4433 9418 4471 9452
rect 4505 9418 4543 9452
rect 4577 9418 4615 9452
rect 4649 9418 4687 9452
rect 4721 9418 4759 9452
rect 4793 9418 4831 9452
rect 4865 9418 4903 9452
rect 4937 9418 4975 9452
rect 5009 9418 5047 9452
rect 5081 9418 5119 9452
rect 5153 9418 5191 9452
rect 5225 9418 5263 9452
rect 5297 9418 5335 9452
rect 5369 9418 5407 9452
rect 5441 9418 5479 9452
rect 5513 9418 5551 9452
rect 5585 9418 5623 9452
rect 5657 9418 5695 9452
rect 5729 9418 5767 9452
rect 5801 9418 5839 9452
rect 5873 9418 5911 9452
rect 5945 9418 5983 9452
rect 6017 9418 6055 9452
rect 6089 9418 6127 9452
rect 6161 9418 6199 9452
rect 6233 9418 6271 9452
rect 6305 9418 6343 9452
rect 6377 9418 6415 9452
rect 6449 9418 6487 9452
rect 6521 9418 6559 9452
rect 6593 9418 6631 9452
rect 6665 9418 6703 9452
rect 6737 9418 6775 9452
rect 6809 9418 6847 9452
rect 6881 9418 6919 9452
rect 6953 9418 6991 9452
rect 7025 9418 7063 9452
rect 7097 9418 7135 9452
rect 7169 9418 7207 9452
rect 7241 9418 7279 9452
rect 7313 9418 7351 9452
rect 7385 9418 7423 9452
rect 7457 9418 7495 9452
rect 7529 9418 7567 9452
rect 7601 9418 7639 9452
rect 7673 9418 7711 9452
rect 7745 9418 7783 9452
rect 7817 9418 7855 9452
rect 7889 9418 7927 9452
rect 7961 9418 7999 9452
rect 8033 9418 8071 9452
rect 8105 9418 8143 9452
rect 8177 9418 8215 9452
rect 8249 9418 8287 9452
rect 8321 9418 8359 9452
rect 8393 9418 8431 9452
rect 8465 9418 8503 9452
rect 8537 9418 8575 9452
rect 8609 9418 8647 9452
rect 8681 9418 8719 9452
rect 8753 9418 8791 9452
rect 8825 9418 8863 9452
rect 8897 9418 8935 9452
rect 8969 9418 9007 9452
rect 9041 9418 9079 9452
rect 9113 9418 9151 9452
rect 9185 9418 9223 9452
rect 9257 9418 9295 9452
rect 9329 9418 9367 9452
rect 9401 9418 9439 9452
rect 9473 9418 9511 9452
rect 9545 9418 9583 9452
rect 9617 9418 9655 9452
rect 9689 9418 9727 9452
rect 9761 9418 9799 9452
rect 9833 9418 9871 9452
rect 9905 9418 9943 9452
rect 9977 9418 10015 9452
rect 10049 9418 10087 9452
rect 10121 9418 10159 9452
rect 10193 9418 10231 9452
rect 10265 9418 10303 9452
rect 10337 9418 10375 9452
rect 10409 9418 10447 9452
rect 10481 9418 10519 9452
rect 10553 9418 10591 9452
rect 10625 9418 10663 9452
rect 10697 9418 10735 9452
rect 10769 9418 10807 9452
rect 10841 9418 10879 9452
rect 10913 9418 10951 9452
rect 10985 9418 11023 9452
rect 11057 9418 11095 9452
rect 11129 9418 11167 9452
rect 11201 9418 11239 9452
rect 11273 9418 11311 9452
rect 12462 9418 12463 9452
rect 12497 9418 12535 9452
rect 12569 9418 12607 9452
rect 12641 9418 12705 9452
rect 2248 9343 2445 9418
rect 858 9252 2096 9295
rect 2396 8983 2445 9343
rect 3585 9343 11322 9418
rect 3585 8983 3635 9343
rect 2396 8939 3635 8983
rect 11273 8984 11322 9343
rect 12462 9343 12705 9418
rect 12462 8984 12512 9343
rect 12858 9295 12908 9731
rect 14048 9295 14096 9731
rect 14539 9838 14724 9876
rect 14539 9804 14614 9838
rect 14648 9804 14724 9838
rect 14539 9766 14724 9804
rect 14539 9732 14614 9766
rect 14648 9732 14724 9766
rect 14539 9694 14724 9732
rect 14539 9660 14614 9694
rect 14648 9660 14724 9694
rect 14539 9528 14724 9660
rect 14232 9452 14724 9528
rect 14232 9418 14314 9452
rect 14348 9418 14614 9452
rect 14648 9418 14724 9452
rect 14232 9343 14724 9418
rect 12858 9252 14096 9295
rect 11273 8940 12512 8984
<< via1 >>
rect 4944 29407 7236 30227
rect 7745 29407 10037 30227
rect 4939 28219 7231 28335
rect 7750 28219 10042 28335
rect 2509 27906 4481 28022
rect 10500 27906 12472 28022
rect 4939 27603 7231 27719
rect 7750 27603 10042 27719
rect 4933 25909 7225 26025
rect 7757 25909 10049 26025
rect 2546 25643 4454 25759
rect 10528 25643 12436 25759
rect 4933 25377 7225 25493
rect 7757 25377 10049 25493
rect 4945 23669 7237 24489
rect 7744 23669 10036 24489
rect 908 9295 2048 9731
rect 2445 9452 3585 9483
rect 11322 9452 12462 9484
rect 2445 9418 2455 9452
rect 2455 9418 2489 9452
rect 2489 9418 2527 9452
rect 2527 9418 2561 9452
rect 2561 9418 2599 9452
rect 2599 9418 2633 9452
rect 2633 9418 2671 9452
rect 2671 9418 2705 9452
rect 2705 9418 2743 9452
rect 2743 9418 2777 9452
rect 2777 9418 2815 9452
rect 2815 9418 2849 9452
rect 2849 9418 2887 9452
rect 2887 9418 2921 9452
rect 2921 9418 2959 9452
rect 2959 9418 2993 9452
rect 2993 9418 3031 9452
rect 3031 9418 3065 9452
rect 3065 9418 3103 9452
rect 3103 9418 3137 9452
rect 3137 9418 3175 9452
rect 3175 9418 3209 9452
rect 3209 9418 3247 9452
rect 3247 9418 3281 9452
rect 3281 9418 3319 9452
rect 3319 9418 3353 9452
rect 3353 9418 3391 9452
rect 3391 9418 3425 9452
rect 3425 9418 3463 9452
rect 3463 9418 3497 9452
rect 3497 9418 3535 9452
rect 3535 9418 3569 9452
rect 3569 9418 3585 9452
rect 11322 9418 11345 9452
rect 11345 9418 11383 9452
rect 11383 9418 11417 9452
rect 11417 9418 11455 9452
rect 11455 9418 11489 9452
rect 11489 9418 11527 9452
rect 11527 9418 11561 9452
rect 11561 9418 11599 9452
rect 11599 9418 11633 9452
rect 11633 9418 11671 9452
rect 11671 9418 11705 9452
rect 11705 9418 11743 9452
rect 11743 9418 11777 9452
rect 11777 9418 11815 9452
rect 11815 9418 11849 9452
rect 11849 9418 11887 9452
rect 11887 9418 11921 9452
rect 11921 9418 11959 9452
rect 11959 9418 11993 9452
rect 11993 9418 12031 9452
rect 12031 9418 12065 9452
rect 12065 9418 12103 9452
rect 12103 9418 12137 9452
rect 12137 9418 12175 9452
rect 12175 9418 12209 9452
rect 12209 9418 12247 9452
rect 12247 9418 12281 9452
rect 12281 9418 12319 9452
rect 12319 9418 12353 9452
rect 12353 9418 12391 9452
rect 12391 9418 12425 9452
rect 12425 9418 12462 9452
rect 2445 8983 3585 9418
rect 11322 8984 12462 9418
rect 12908 9295 14048 9731
<< metal2 >>
tri 4891 39322 4991 39422 se
rect 4991 39322 7191 39422
tri 7191 39322 7291 39422 sw
rect 4891 39213 7291 39322
rect 4891 35317 4979 39213
rect 7195 35317 7291 39213
rect 4891 30227 7291 35317
rect 4891 29407 4944 30227
rect 7236 29407 7291 30227
tri 301 28975 501 29175 se
rect 501 28975 4291 29175
tri 4291 28975 4491 29175 sw
rect 301 28869 4491 28975
rect 301 23293 466 28869
rect 2442 28022 4491 28869
rect 2442 27906 2509 28022
rect 4481 27906 4491 28022
rect 2442 25759 4491 27906
rect 4891 28335 7291 29407
rect 4891 28219 4939 28335
rect 7231 28219 7291 28335
rect 4891 27719 7291 28219
rect 4891 27603 4939 27719
rect 7231 27603 7291 27719
rect 4891 27317 7291 27603
tri 4891 27117 5091 27317 ne
rect 5091 27117 7091 27317
tri 7091 27117 7291 27317 nw
tri 7691 39322 7791 39422 se
rect 7791 39322 9991 39422
tri 9991 39322 10091 39422 sw
rect 7691 39213 10091 39322
rect 7691 35317 7779 39213
rect 9995 35317 10091 39213
rect 7691 30227 10091 35317
rect 7691 29407 7745 30227
rect 10037 29407 10091 30227
rect 7691 28335 10091 29407
rect 7691 28219 7750 28335
rect 10042 28219 10091 28335
rect 7691 27719 10091 28219
rect 7691 27603 7750 27719
rect 10042 27603 10091 27719
rect 7691 27317 10091 27603
tri 7691 27117 7891 27317 ne
rect 7891 27117 9891 27317
tri 9891 27117 10091 27317 nw
tri 10491 28975 10691 29175 se
rect 10691 28975 14431 29175
tri 14431 28975 14631 29175 sw
rect 10491 28917 14631 28975
rect 10491 28022 12455 28917
rect 10491 27906 10500 28022
rect 2442 25643 2546 25759
rect 4454 25643 4491 25759
rect 2442 23293 4491 25643
rect 301 23016 4491 23293
tri 301 22816 501 23016 ne
rect 501 22816 4291 23016
tri 4291 22816 4491 23016 nw
tri 4891 26278 5091 26478 se
rect 5091 26278 7091 26478
tri 7091 26278 7291 26478 sw
rect 4891 26025 7291 26278
rect 4891 25909 4933 26025
rect 7225 25909 7291 26025
rect 4891 25493 7291 25909
rect 4891 25377 4933 25493
rect 7225 25377 7291 25493
rect 4891 24489 7291 25377
rect 4891 23669 4945 24489
rect 7237 23669 7291 24489
rect 4891 18931 7291 23669
rect 4891 17275 4942 18931
rect 7238 17275 7291 18931
rect 4891 17214 7291 17275
rect 4891 17086 5103 17214
tri 4891 16986 4991 17086 ne
rect 4991 17078 5103 17086
rect 7239 17078 7291 17214
rect 4991 17056 7291 17078
rect 4991 16986 7221 17056
tri 7221 16986 7291 17056 nw
tri 7691 26278 7891 26478 se
rect 7891 26278 9891 26478
tri 9891 26278 10091 26478 sw
rect 7691 26025 10091 26278
rect 7691 25909 7757 26025
rect 10049 25909 10091 26025
rect 7691 25493 10091 25909
rect 7691 25377 7757 25493
rect 10049 25377 10091 25493
rect 7691 24489 10091 25377
rect 7691 23669 7744 24489
rect 10036 23669 10091 24489
rect 7691 18931 10091 23669
rect 10491 25759 12455 27906
rect 10491 25643 10528 25759
rect 12436 25643 12455 25759
rect 10491 23341 12455 25643
rect 14431 23341 14631 28917
rect 10491 23016 14631 23341
tri 10491 22816 10691 23016 ne
rect 10691 22816 14431 23016
tri 14431 22816 14631 23016 nw
rect 7691 17275 7742 18931
rect 10038 17275 10091 18931
rect 7691 17214 10091 17275
rect 7691 17078 7739 17214
rect 9875 17086 10091 17214
rect 9875 17078 9991 17086
rect 7691 17056 9991 17078
tri 7691 16986 7761 17056 ne
rect 7761 16986 9991 17056
tri 9991 16986 10091 17086 nw
rect 858 9741 2096 9772
rect 858 9285 890 9741
rect 2066 9285 2096 9741
rect 12858 9741 14096 9772
rect 858 9252 2096 9285
rect 2396 9501 3635 9528
rect 2396 8965 2427 9501
rect 3603 8965 3635 9501
rect 2396 8939 3635 8965
rect 11273 9502 12512 9529
rect 11273 8966 11304 9502
rect 12480 8966 12512 9502
rect 12858 9285 12890 9741
rect 14066 9285 14096 9741
rect 12858 9252 14096 9285
rect 11273 8940 12512 8966
<< via2 >>
rect 4979 35317 7195 39213
rect 466 23293 2442 28869
rect 7779 35317 9995 39213
rect 12455 28022 14431 28917
rect 12455 27906 12472 28022
rect 12472 27906 14431 28022
rect 4942 17275 7238 18931
rect 5103 17078 7239 17214
rect 12455 23341 14431 27906
rect 7742 17275 10038 18931
rect 7739 17078 9875 17214
rect 890 9731 2066 9741
rect 890 9295 908 9731
rect 908 9295 2048 9731
rect 2048 9295 2066 9731
rect 890 9285 2066 9295
rect 2427 9483 3603 9501
rect 2427 8983 2445 9483
rect 2445 8983 3585 9483
rect 3585 8983 3603 9483
rect 2427 8965 3603 8983
rect 11304 9484 12480 9502
rect 11304 8984 11322 9484
rect 11322 8984 12462 9484
rect 12462 8984 12480 9484
rect 11304 8966 12480 8984
rect 12890 9731 14066 9741
rect 12890 9295 12908 9731
rect 12908 9295 14048 9731
rect 14048 9295 14066 9731
rect 12890 9285 14066 9295
<< metal3 >>
tri 4805 39522 5205 39922 se
rect 5205 39522 9786 39922
tri 9786 39522 10186 39922 sw
rect 4805 39217 10186 39522
rect 4805 35313 4975 39217
rect 7199 35313 7775 39217
rect 9999 35313 10186 39217
rect 4805 35266 10186 35313
tri 4805 35166 4905 35266 ne
rect 4905 35166 10086 35266
tri 10086 35166 10186 35266 nw
tri 99 33575 1155 34631 se
rect 1155 34604 3100 34631
rect 1155 34540 2276 34604
rect 2340 34540 2359 34604
rect 2423 34540 2443 34604
rect 2507 34540 2527 34604
rect 2591 34540 2611 34604
rect 2675 34540 3100 34604
rect 1155 34510 3100 34540
rect 1155 34446 2276 34510
rect 2340 34446 2359 34510
rect 2423 34446 2443 34510
rect 2507 34446 2527 34510
rect 2591 34446 2611 34510
rect 2675 34446 3100 34510
rect 1155 34427 3100 34446
rect 1155 34363 2148 34427
rect 2212 34416 3100 34427
rect 2212 34363 2276 34416
rect 1155 34352 2276 34363
rect 2340 34352 2359 34416
rect 2423 34352 2443 34416
rect 2507 34352 2527 34416
rect 2591 34352 2611 34416
rect 2675 34352 3100 34416
rect 1155 34322 3100 34352
rect 1155 34302 2276 34322
rect 1155 34238 2004 34302
rect 2068 34238 2084 34302
rect 2148 34238 2164 34302
rect 2228 34258 2276 34302
rect 2340 34258 2359 34322
rect 2423 34258 2443 34322
rect 2507 34258 2527 34322
rect 2591 34258 2611 34322
rect 2675 34258 3100 34322
rect 2228 34238 3100 34258
rect 1155 34228 3100 34238
rect 1155 34206 2276 34228
rect 1155 34169 2004 34206
rect 1155 34105 1890 34169
rect 1954 34142 2004 34169
rect 2068 34142 2084 34206
rect 2148 34142 2164 34206
rect 2228 34164 2276 34206
rect 2340 34164 2359 34228
rect 2423 34164 2443 34228
rect 2507 34164 2527 34228
rect 2591 34164 2611 34228
rect 2675 34164 3100 34228
rect 2228 34142 3100 34164
rect 1954 34134 3100 34142
rect 1954 34105 2276 34134
rect 1155 34070 2276 34105
rect 2340 34070 2359 34134
rect 2423 34070 2443 34134
rect 2507 34070 2527 34134
rect 2591 34070 2611 34134
rect 2675 34070 3100 34134
rect 1155 34064 3100 34070
rect 1155 34000 1748 34064
rect 1812 34000 1837 34064
rect 1901 34000 1927 34064
rect 1991 34000 2017 34064
rect 2081 34000 2107 34064
rect 2171 34000 3100 34064
rect 1155 33995 3100 34000
rect 1155 33948 2247 33995
rect 1155 33884 1748 33948
rect 1812 33884 1837 33948
rect 1901 33884 1927 33948
rect 1991 33884 2017 33948
rect 2081 33884 2107 33948
rect 2171 33931 2247 33948
rect 2311 33931 3100 33995
rect 2171 33884 3100 33931
rect 1155 33872 3100 33884
rect 1155 33808 1644 33872
rect 1708 33848 3100 33872
rect 1708 33832 2700 33848
rect 1708 33808 1748 33832
rect 1155 33768 1748 33808
rect 1812 33768 1837 33832
rect 1901 33768 1927 33832
rect 1991 33768 2017 33832
rect 2081 33768 2107 33832
rect 2171 33768 2700 33832
rect 1155 33740 2700 33768
rect 1155 33676 1424 33740
rect 1488 33676 1513 33740
rect 1577 33676 1603 33740
rect 1667 33676 1693 33740
rect 1757 33676 1783 33740
rect 1847 33707 2700 33740
rect 1847 33676 1929 33707
rect 1155 33643 1929 33676
rect 1993 33643 2700 33707
rect 1155 33624 2700 33643
rect 1155 33575 1424 33624
rect 99 33560 1424 33575
rect 1488 33560 1513 33624
rect 1577 33560 1603 33624
rect 1667 33560 1693 33624
rect 1757 33560 1783 33624
rect 1847 33560 2700 33624
rect 99 33544 2700 33560
rect 99 33480 1316 33544
rect 1380 33508 2700 33544
rect 1380 33480 1424 33508
rect 99 33444 1424 33480
rect 1488 33444 1513 33508
rect 1577 33444 1603 33508
rect 1667 33444 1693 33508
rect 1757 33444 1783 33508
rect 1847 33444 2700 33508
tri 2700 33448 3100 33848 nw
rect 11900 34604 13835 34631
rect 11900 34540 12341 34604
rect 12405 34540 12425 34604
rect 12489 34540 12509 34604
rect 12573 34540 12593 34604
rect 12657 34540 12677 34604
rect 12741 34540 13835 34604
rect 11900 34510 13835 34540
rect 11900 34446 12341 34510
rect 12405 34446 12425 34510
rect 12489 34446 12509 34510
rect 12573 34446 12593 34510
rect 12657 34446 12677 34510
rect 12741 34446 13835 34510
rect 11900 34427 13835 34446
rect 11900 34416 12804 34427
rect 11900 34352 12341 34416
rect 12405 34352 12425 34416
rect 12489 34352 12509 34416
rect 12573 34352 12593 34416
rect 12657 34352 12677 34416
rect 12741 34363 12804 34416
rect 12868 34363 13835 34427
rect 12741 34352 13835 34363
rect 11900 34322 13835 34352
rect 11900 34258 12341 34322
rect 12405 34258 12425 34322
rect 12489 34258 12509 34322
rect 12573 34258 12593 34322
rect 12657 34258 12677 34322
rect 12741 34302 13835 34322
rect 12741 34258 12788 34302
rect 11900 34238 12788 34258
rect 12852 34238 12868 34302
rect 12932 34238 12948 34302
rect 13012 34238 13835 34302
rect 11900 34228 13835 34238
rect 11900 34164 12341 34228
rect 12405 34164 12425 34228
rect 12489 34164 12509 34228
rect 12573 34164 12593 34228
rect 12657 34164 12677 34228
rect 12741 34206 13835 34228
rect 12741 34164 12788 34206
rect 11900 34142 12788 34164
rect 12852 34142 12868 34206
rect 12932 34142 12948 34206
rect 13012 34169 13835 34206
rect 13012 34142 13062 34169
rect 11900 34134 13062 34142
rect 11900 34070 12341 34134
rect 12405 34070 12425 34134
rect 12489 34070 12509 34134
rect 12573 34070 12593 34134
rect 12657 34070 12677 34134
rect 12741 34105 13062 34134
rect 13126 34105 13835 34169
rect 12741 34070 13835 34105
rect 11900 34064 13835 34070
rect 11900 34000 12845 34064
rect 12909 34000 12935 34064
rect 12999 34000 13025 34064
rect 13089 34000 13115 34064
rect 13179 34000 13204 34064
rect 13268 34000 13835 34064
rect 11900 33995 13835 34000
rect 11900 33931 12705 33995
rect 12769 33948 13835 33995
rect 12769 33931 12845 33948
rect 11900 33884 12845 33931
rect 12909 33884 12935 33948
rect 12999 33884 13025 33948
rect 13089 33884 13115 33948
rect 13179 33884 13204 33948
rect 13268 33884 13835 33948
rect 11900 33872 13835 33884
rect 11900 33848 13308 33872
tri 11900 33448 12300 33848 ne
rect 12300 33832 13308 33848
rect 12300 33768 12845 33832
rect 12909 33768 12935 33832
rect 12999 33768 13025 33832
rect 13089 33768 13115 33832
rect 13179 33768 13204 33832
rect 13268 33808 13308 33832
rect 13372 33808 13835 33872
rect 13268 33768 13835 33808
rect 12300 33740 13835 33768
rect 12300 33707 13169 33740
rect 12300 33643 13023 33707
rect 13087 33676 13169 33707
rect 13233 33676 13259 33740
rect 13323 33676 13349 33740
rect 13413 33676 13439 33740
rect 13503 33676 13528 33740
rect 13592 33676 13835 33740
rect 13087 33643 13835 33676
rect 12300 33624 13835 33643
rect 12300 33560 13169 33624
rect 13233 33560 13259 33624
rect 13323 33560 13349 33624
rect 13413 33560 13439 33624
rect 13503 33560 13528 33624
rect 13592 33608 13835 33624
tri 13835 33608 14858 34631 sw
rect 13592 33560 14858 33608
rect 12300 33544 14858 33560
rect 12300 33508 13636 33544
rect 99 33420 2700 33444
rect 99 33356 1104 33420
rect 1168 33356 1193 33420
rect 1257 33356 1283 33420
rect 1347 33356 1373 33420
rect 1437 33356 1463 33420
rect 1527 33382 2700 33420
rect 1527 33356 1604 33382
rect 99 33318 1604 33356
rect 1668 33318 2700 33382
rect 99 33304 2700 33318
rect 99 33240 1104 33304
rect 1168 33240 1193 33304
rect 1257 33240 1283 33304
rect 1347 33240 1373 33304
rect 1437 33240 1463 33304
rect 1527 33240 2700 33304
rect 99 33188 2700 33240
rect 99 33124 1104 33188
rect 1168 33124 1193 33188
rect 1257 33124 1283 33188
rect 1347 33124 1373 33188
rect 1437 33124 1463 33188
rect 1527 33124 2700 33188
rect 99 33095 2700 33124
rect 99 33031 982 33095
rect 1046 33031 1072 33095
rect 1136 33031 1162 33095
rect 1226 33031 1252 33095
rect 1316 33031 1342 33095
rect 1406 33031 1432 33095
rect 1496 33031 2700 33095
rect 99 33015 2700 33031
rect 99 32951 982 33015
rect 1046 32951 1072 33015
rect 1136 32951 1162 33015
rect 1226 32951 1252 33015
rect 1316 32951 1342 33015
rect 1406 32951 1432 33015
rect 1496 32951 2700 33015
rect 99 32935 2700 32951
rect 99 32871 982 32935
rect 1046 32871 1072 32935
rect 1136 32871 1162 32935
rect 1226 32871 1252 32935
rect 1316 32871 1342 32935
rect 1406 32871 1432 32935
rect 1496 32871 2700 32935
rect 99 32855 2700 32871
rect 99 32791 982 32855
rect 1046 32791 1072 32855
rect 1136 32791 1162 32855
rect 1226 32791 1252 32855
rect 1316 32791 1342 32855
rect 1406 32791 1432 32855
rect 1496 32791 2700 32855
rect 99 32775 2700 32791
rect 99 32711 982 32775
rect 1046 32711 1072 32775
rect 1136 32711 1162 32775
rect 1226 32711 1252 32775
rect 1316 32711 1342 32775
rect 1406 32711 1432 32775
rect 1496 32711 2700 32775
rect 99 32695 2700 32711
rect 99 32631 982 32695
rect 1046 32631 1072 32695
rect 1136 32631 1162 32695
rect 1226 32631 1252 32695
rect 1316 32631 1342 32695
rect 1406 32631 1432 32695
rect 1496 32631 2700 32695
rect 99 32615 2700 32631
rect 99 32551 982 32615
rect 1046 32551 1072 32615
rect 1136 32551 1162 32615
rect 1226 32551 1252 32615
rect 1316 32551 1342 32615
rect 1406 32551 1432 32615
rect 1496 32551 2700 32615
rect 99 32535 2700 32551
rect 99 32471 982 32535
rect 1046 32471 1072 32535
rect 1136 32471 1162 32535
rect 1226 32471 1252 32535
rect 1316 32471 1342 32535
rect 1406 32471 1432 32535
rect 1496 32471 2700 32535
rect 99 32455 2700 32471
rect 99 32391 982 32455
rect 1046 32391 1072 32455
rect 1136 32391 1162 32455
rect 1226 32391 1252 32455
rect 1316 32391 1342 32455
rect 1406 32391 1432 32455
rect 1496 32391 2700 32455
rect 99 32375 2700 32391
rect 99 32311 982 32375
rect 1046 32311 1072 32375
rect 1136 32311 1162 32375
rect 1226 32311 1252 32375
rect 1316 32311 1342 32375
rect 1406 32311 1432 32375
rect 1496 32311 2700 32375
rect 99 32295 2700 32311
rect 99 32231 982 32295
rect 1046 32231 1072 32295
rect 1136 32231 1162 32295
rect 1226 32231 1252 32295
rect 1316 32231 1342 32295
rect 1406 32231 1432 32295
rect 1496 32231 2700 32295
rect 99 32215 2700 32231
rect 99 32151 982 32215
rect 1046 32151 1072 32215
rect 1136 32151 1162 32215
rect 1226 32151 1252 32215
rect 1316 32151 1342 32215
rect 1406 32151 1432 32215
rect 1496 32151 2700 32215
rect 99 32135 2700 32151
rect 99 32071 982 32135
rect 1046 32071 1072 32135
rect 1136 32071 1162 32135
rect 1226 32071 1252 32135
rect 1316 32071 1342 32135
rect 1406 32071 1432 32135
rect 1496 32071 2700 32135
rect 99 32055 2700 32071
rect 99 31991 982 32055
rect 1046 31991 1072 32055
rect 1136 31991 1162 32055
rect 1226 31991 1252 32055
rect 1316 31991 1342 32055
rect 1406 31991 1432 32055
rect 1496 31991 2700 32055
rect 99 31975 2700 31991
rect 99 31911 982 31975
rect 1046 31911 1072 31975
rect 1136 31911 1162 31975
rect 1226 31911 1252 31975
rect 1316 31911 1342 31975
rect 1406 31911 1432 31975
rect 1496 31911 2700 31975
rect 99 31895 2700 31911
rect 99 31831 982 31895
rect 1046 31831 1072 31895
rect 1136 31831 1162 31895
rect 1226 31831 1252 31895
rect 1316 31831 1342 31895
rect 1406 31831 1432 31895
rect 1496 31831 2700 31895
rect 99 31815 2700 31831
rect 99 31751 982 31815
rect 1046 31751 1072 31815
rect 1136 31751 1162 31815
rect 1226 31751 1252 31815
rect 1316 31751 1342 31815
rect 1406 31751 1432 31815
rect 1496 31751 2700 31815
rect 99 31735 2700 31751
rect 99 31671 982 31735
rect 1046 31671 1072 31735
rect 1136 31671 1162 31735
rect 1226 31671 1252 31735
rect 1316 31671 1342 31735
rect 1406 31671 1432 31735
rect 1496 31671 2700 31735
rect 99 31655 2700 31671
rect 99 31591 982 31655
rect 1046 31591 1072 31655
rect 1136 31591 1162 31655
rect 1226 31591 1252 31655
rect 1316 31591 1342 31655
rect 1406 31591 1432 31655
rect 1496 31591 2700 31655
rect 99 31575 2700 31591
rect 99 31511 982 31575
rect 1046 31511 1072 31575
rect 1136 31511 1162 31575
rect 1226 31511 1252 31575
rect 1316 31511 1342 31575
rect 1406 31511 1432 31575
rect 1496 31511 2700 31575
rect 99 31495 2700 31511
rect 99 31431 982 31495
rect 1046 31431 1072 31495
rect 1136 31431 1162 31495
rect 1226 31431 1252 31495
rect 1316 31431 1342 31495
rect 1406 31431 1432 31495
rect 1496 31431 2700 31495
rect 99 31415 2700 31431
rect 99 31351 982 31415
rect 1046 31351 1072 31415
rect 1136 31351 1162 31415
rect 1226 31351 1252 31415
rect 1316 31351 1342 31415
rect 1406 31351 1432 31415
rect 1496 31351 2700 31415
rect 99 31335 2700 31351
rect 99 31271 982 31335
rect 1046 31271 1072 31335
rect 1136 31271 1162 31335
rect 1226 31271 1252 31335
rect 1316 31271 1342 31335
rect 1406 31271 1432 31335
rect 1496 31271 2700 31335
rect 99 31255 2700 31271
rect 99 31191 982 31255
rect 1046 31191 1072 31255
rect 1136 31191 1162 31255
rect 1226 31191 1252 31255
rect 1316 31191 1342 31255
rect 1406 31191 1432 31255
rect 1496 31191 2700 31255
rect 99 31175 2700 31191
rect 99 31111 982 31175
rect 1046 31111 1072 31175
rect 1136 31111 1162 31175
rect 1226 31111 1252 31175
rect 1316 31111 1342 31175
rect 1406 31111 1432 31175
rect 1496 31111 2700 31175
rect 99 31095 2700 31111
rect 99 31031 982 31095
rect 1046 31031 1072 31095
rect 1136 31031 1162 31095
rect 1226 31031 1252 31095
rect 1316 31031 1342 31095
rect 1406 31031 1432 31095
rect 1496 31031 2700 31095
rect 99 31015 2700 31031
rect 99 30951 982 31015
rect 1046 30951 1072 31015
rect 1136 30951 1162 31015
rect 1226 30951 1252 31015
rect 1316 30951 1342 31015
rect 1406 30951 1432 31015
rect 1496 30951 2700 31015
rect 99 30935 2700 30951
rect 99 30871 982 30935
rect 1046 30871 1072 30935
rect 1136 30871 1162 30935
rect 1226 30871 1252 30935
rect 1316 30871 1342 30935
rect 1406 30871 1432 30935
rect 1496 30871 2700 30935
rect 99 30855 2700 30871
rect 99 30791 982 30855
rect 1046 30791 1072 30855
rect 1136 30791 1162 30855
rect 1226 30791 1252 30855
rect 1316 30791 1342 30855
rect 1406 30791 1432 30855
rect 1496 30791 2700 30855
rect 99 30775 2700 30791
rect 99 30711 982 30775
rect 1046 30711 1072 30775
rect 1136 30711 1162 30775
rect 1226 30711 1252 30775
rect 1316 30711 1342 30775
rect 1406 30711 1432 30775
rect 1496 30711 2700 30775
rect 99 30695 2700 30711
rect 99 30631 982 30695
rect 1046 30631 1072 30695
rect 1136 30631 1162 30695
rect 1226 30631 1252 30695
rect 1316 30631 1342 30695
rect 1406 30631 1432 30695
rect 1496 30631 2700 30695
rect 99 30615 2700 30631
rect 99 30551 982 30615
rect 1046 30551 1072 30615
rect 1136 30551 1162 30615
rect 1226 30551 1252 30615
rect 1316 30551 1342 30615
rect 1406 30551 1432 30615
rect 1496 30551 2700 30615
rect 99 30535 2700 30551
rect 99 30471 982 30535
rect 1046 30471 1072 30535
rect 1136 30471 1162 30535
rect 1226 30471 1252 30535
rect 1316 30471 1342 30535
rect 1406 30471 1432 30535
rect 1496 30471 2700 30535
rect 99 30455 2700 30471
rect 99 30391 982 30455
rect 1046 30391 1072 30455
rect 1136 30391 1162 30455
rect 1226 30391 1252 30455
rect 1316 30391 1342 30455
rect 1406 30391 1432 30455
rect 1496 30391 2700 30455
rect 99 30375 2700 30391
rect 99 30311 982 30375
rect 1046 30311 1072 30375
rect 1136 30311 1162 30375
rect 1226 30311 1252 30375
rect 1316 30311 1342 30375
rect 1406 30311 1432 30375
rect 1496 30311 2700 30375
rect 99 30295 2700 30311
rect 99 30231 982 30295
rect 1046 30231 1072 30295
rect 1136 30231 1162 30295
rect 1226 30231 1252 30295
rect 1316 30231 1342 30295
rect 1406 30231 1432 30295
rect 1496 30231 2700 30295
rect 99 30215 2700 30231
rect 99 30151 982 30215
rect 1046 30151 1072 30215
rect 1136 30151 1162 30215
rect 1226 30151 1252 30215
rect 1316 30151 1342 30215
rect 1406 30151 1432 30215
rect 1496 30151 2700 30215
rect 99 30135 2700 30151
rect 99 30071 982 30135
rect 1046 30071 1072 30135
rect 1136 30071 1162 30135
rect 1226 30071 1252 30135
rect 1316 30071 1342 30135
rect 1406 30071 1432 30135
rect 1496 30071 2700 30135
rect 99 30055 2700 30071
rect 99 29991 982 30055
rect 1046 29991 1072 30055
rect 1136 29991 1162 30055
rect 1226 29991 1252 30055
rect 1316 29991 1342 30055
rect 1406 29991 1432 30055
rect 1496 29991 2700 30055
rect 99 29975 2700 29991
rect 99 29911 982 29975
rect 1046 29911 1072 29975
rect 1136 29911 1162 29975
rect 1226 29911 1252 29975
rect 1316 29911 1342 29975
rect 1406 29911 1432 29975
rect 1496 29911 2700 29975
rect 99 29895 2700 29911
rect 99 29831 982 29895
rect 1046 29831 1072 29895
rect 1136 29831 1162 29895
rect 1226 29831 1252 29895
rect 1316 29831 1342 29895
rect 1406 29831 1432 29895
rect 1496 29831 2700 29895
rect 99 29815 2700 29831
rect 99 29751 982 29815
rect 1046 29751 1072 29815
rect 1136 29751 1162 29815
rect 1226 29751 1252 29815
rect 1316 29751 1342 29815
rect 1406 29751 1432 29815
rect 1496 29751 2700 29815
rect 99 29735 2700 29751
rect 99 29671 982 29735
rect 1046 29671 1072 29735
rect 1136 29671 1162 29735
rect 1226 29671 1252 29735
rect 1316 29671 1342 29735
rect 1406 29671 1432 29735
rect 1496 29671 2700 29735
rect 99 29655 2700 29671
rect 99 29591 982 29655
rect 1046 29591 1072 29655
rect 1136 29591 1162 29655
rect 1226 29591 1252 29655
rect 1316 29591 1342 29655
rect 1406 29591 1432 29655
rect 1496 29591 2700 29655
rect 99 29575 2700 29591
rect 99 29511 982 29575
rect 1046 29511 1072 29575
rect 1136 29511 1162 29575
rect 1226 29511 1252 29575
rect 1316 29511 1342 29575
rect 1406 29511 1432 29575
rect 1496 29511 2700 29575
rect 99 29495 2700 29511
rect 99 29431 982 29495
rect 1046 29431 1072 29495
rect 1136 29431 1162 29495
rect 1226 29431 1252 29495
rect 1316 29431 1342 29495
rect 1406 29431 1432 29495
rect 1496 29431 2700 29495
rect 99 29415 2700 29431
rect 99 29351 982 29415
rect 1046 29351 1072 29415
rect 1136 29351 1162 29415
rect 1226 29351 1252 29415
rect 1316 29351 1342 29415
rect 1406 29351 1432 29415
rect 1496 29351 2700 29415
rect 99 29335 2700 29351
rect 99 29271 982 29335
rect 1046 29271 1072 29335
rect 1136 29271 1162 29335
rect 1226 29271 1252 29335
rect 1316 29271 1342 29335
rect 1406 29271 1432 29335
rect 1496 29271 2700 29335
rect 99 29255 2700 29271
rect 99 29191 982 29255
rect 1046 29191 1072 29255
rect 1136 29191 1162 29255
rect 1226 29191 1252 29255
rect 1316 29191 1342 29255
rect 1406 29191 1432 29255
rect 1496 29191 2700 29255
rect 99 29175 2700 29191
rect 99 29111 982 29175
rect 1046 29111 1072 29175
rect 1136 29111 1162 29175
rect 1226 29111 1252 29175
rect 1316 29111 1342 29175
rect 1406 29111 1432 29175
rect 1496 29111 2700 29175
rect 99 29095 2700 29111
rect 99 29031 982 29095
rect 1046 29031 1072 29095
rect 1136 29031 1162 29095
rect 1226 29031 1252 29095
rect 1316 29031 1342 29095
rect 1406 29031 1432 29095
rect 1496 29031 2700 29095
rect 99 29015 2700 29031
rect 99 28951 982 29015
rect 1046 28951 1072 29015
rect 1136 28951 1162 29015
rect 1226 28951 1252 29015
rect 1316 28951 1342 29015
rect 1406 28951 1432 29015
rect 1496 28951 2700 29015
rect 99 28935 2700 28951
rect 99 28871 982 28935
rect 1046 28871 1072 28935
rect 1136 28871 1162 28935
rect 1226 28871 1252 28935
rect 1316 28871 1342 28935
rect 1406 28871 1432 28935
rect 1496 28871 2700 28935
rect 99 28869 2700 28871
rect 99 23293 466 28869
rect 2442 23293 2700 28869
rect 99 23271 982 23293
rect 1046 23271 1072 23293
rect 1136 23271 1162 23293
rect 1226 23271 1252 23293
rect 1316 23271 1342 23293
rect 1406 23271 1432 23293
rect 1496 23271 2700 23293
rect 99 23254 2700 23271
rect 99 23190 982 23254
rect 1046 23190 1072 23254
rect 1136 23190 1162 23254
rect 1226 23190 1252 23254
rect 1316 23190 1342 23254
rect 1406 23190 1432 23254
rect 1496 23190 2700 23254
rect 99 23173 2700 23190
rect 99 23109 982 23173
rect 1046 23109 1072 23173
rect 1136 23109 1162 23173
rect 1226 23109 1252 23173
rect 1316 23109 1342 23173
rect 1406 23109 1432 23173
rect 1496 23109 2700 23173
rect 99 23092 2700 23109
rect 99 23028 982 23092
rect 1046 23028 1072 23092
rect 1136 23028 1162 23092
rect 1226 23028 1252 23092
rect 1316 23028 1342 23092
rect 1406 23028 1432 23092
rect 1496 23028 2700 23092
rect 99 23011 2700 23028
rect 99 22947 982 23011
rect 1046 22947 1072 23011
rect 1136 22947 1162 23011
rect 1226 22947 1252 23011
rect 1316 22947 1342 23011
rect 1406 22947 1432 23011
rect 1496 22947 2700 23011
rect 99 22930 2700 22947
rect 99 22866 982 22930
rect 1046 22866 1072 22930
rect 1136 22866 1162 22930
rect 1226 22866 1252 22930
rect 1316 22866 1342 22930
rect 1406 22866 1432 22930
rect 1496 22866 2700 22930
rect 99 22849 2700 22866
rect 99 22785 982 22849
rect 1046 22785 1072 22849
rect 1136 22785 1162 22849
rect 1226 22785 1252 22849
rect 1316 22785 1342 22849
rect 1406 22785 1432 22849
rect 1496 22785 2700 22849
rect 99 22768 2700 22785
rect 99 22704 982 22768
rect 1046 22704 1072 22768
rect 1136 22704 1162 22768
rect 1226 22704 1252 22768
rect 1316 22704 1342 22768
rect 1406 22704 1432 22768
rect 1496 22704 2700 22768
rect 99 22687 2700 22704
rect 99 22623 982 22687
rect 1046 22623 1072 22687
rect 1136 22623 1162 22687
rect 1226 22623 1252 22687
rect 1316 22623 1342 22687
rect 1406 22623 1432 22687
rect 1496 22623 2700 22687
rect 99 22606 2700 22623
rect 99 22542 982 22606
rect 1046 22542 1072 22606
rect 1136 22542 1162 22606
rect 1226 22542 1252 22606
rect 1316 22542 1342 22606
rect 1406 22542 1432 22606
rect 1496 22542 2700 22606
rect 99 22525 2700 22542
rect 99 22461 982 22525
rect 1046 22461 1072 22525
rect 1136 22461 1162 22525
rect 1226 22461 1252 22525
rect 1316 22461 1342 22525
rect 1406 22461 1432 22525
rect 1496 22461 2700 22525
rect 99 22444 2700 22461
rect 99 22380 982 22444
rect 1046 22380 1072 22444
rect 1136 22380 1162 22444
rect 1226 22380 1252 22444
rect 1316 22380 1342 22444
rect 1406 22380 1432 22444
rect 1496 22380 2700 22444
rect 99 22363 2700 22380
rect 99 22299 982 22363
rect 1046 22299 1072 22363
rect 1136 22299 1162 22363
rect 1226 22299 1252 22363
rect 1316 22299 1342 22363
rect 1406 22299 1432 22363
rect 1496 22299 2700 22363
rect 99 22282 2700 22299
rect 99 22218 982 22282
rect 1046 22218 1072 22282
rect 1136 22218 1162 22282
rect 1226 22218 1252 22282
rect 1316 22218 1342 22282
rect 1406 22218 1432 22282
rect 1496 22218 2700 22282
rect 99 22201 2700 22218
rect 99 22137 982 22201
rect 1046 22137 1072 22201
rect 1136 22137 1162 22201
rect 1226 22137 1252 22201
rect 1316 22137 1342 22201
rect 1406 22137 1432 22201
rect 1496 22137 2700 22201
rect 99 22120 2700 22137
rect 99 22056 982 22120
rect 1046 22056 1072 22120
rect 1136 22056 1162 22120
rect 1226 22056 1252 22120
rect 1316 22056 1342 22120
rect 1406 22056 1432 22120
rect 1496 22056 2700 22120
rect 99 22039 2700 22056
rect 99 21975 982 22039
rect 1046 21975 1072 22039
rect 1136 21975 1162 22039
rect 1226 21975 1252 22039
rect 1316 21975 1342 22039
rect 1406 21975 1432 22039
rect 1496 21975 2700 22039
rect 99 21958 2700 21975
rect 99 21894 982 21958
rect 1046 21894 1072 21958
rect 1136 21894 1162 21958
rect 1226 21894 1252 21958
rect 1316 21894 1342 21958
rect 1406 21894 1432 21958
rect 1496 21894 2700 21958
rect 99 21877 2700 21894
rect 99 21813 982 21877
rect 1046 21813 1072 21877
rect 1136 21813 1162 21877
rect 1226 21813 1252 21877
rect 1316 21813 1342 21877
rect 1406 21813 1432 21877
rect 1496 21813 2700 21877
rect 99 21796 2700 21813
rect 99 21732 982 21796
rect 1046 21732 1072 21796
rect 1136 21732 1162 21796
rect 1226 21732 1252 21796
rect 1316 21732 1342 21796
rect 1406 21732 1432 21796
rect 1496 21732 2700 21796
rect 99 21715 2700 21732
rect 99 21651 982 21715
rect 1046 21651 1072 21715
rect 1136 21651 1162 21715
rect 1226 21651 1252 21715
rect 1316 21651 1342 21715
rect 1406 21651 1432 21715
rect 1496 21651 2700 21715
rect 99 21634 2700 21651
rect 99 21570 982 21634
rect 1046 21570 1072 21634
rect 1136 21570 1162 21634
rect 1226 21570 1252 21634
rect 1316 21570 1342 21634
rect 1406 21570 1432 21634
rect 1496 21570 2700 21634
rect 99 21553 2700 21570
rect 99 21489 982 21553
rect 1046 21489 1072 21553
rect 1136 21489 1162 21553
rect 1226 21489 1252 21553
rect 1316 21489 1342 21553
rect 1406 21489 1432 21553
rect 1496 21489 2700 21553
rect 99 21472 2700 21489
rect 99 21408 982 21472
rect 1046 21408 1072 21472
rect 1136 21408 1162 21472
rect 1226 21408 1252 21472
rect 1316 21408 1342 21472
rect 1406 21408 1432 21472
rect 1496 21408 2700 21472
rect 99 21391 2700 21408
rect 99 21327 982 21391
rect 1046 21327 1072 21391
rect 1136 21327 1162 21391
rect 1226 21327 1252 21391
rect 1316 21327 1342 21391
rect 1406 21327 1432 21391
rect 1496 21327 2700 21391
rect 99 21310 2700 21327
rect 99 21246 982 21310
rect 1046 21246 1072 21310
rect 1136 21246 1162 21310
rect 1226 21246 1252 21310
rect 1316 21246 1342 21310
rect 1406 21246 1432 21310
rect 1496 21246 2700 21310
rect 99 21229 2700 21246
rect 99 21165 982 21229
rect 1046 21165 1072 21229
rect 1136 21165 1162 21229
rect 1226 21165 1252 21229
rect 1316 21165 1342 21229
rect 1406 21165 1432 21229
rect 1496 21165 2700 21229
rect 99 21148 2700 21165
rect 99 21084 982 21148
rect 1046 21084 1072 21148
rect 1136 21084 1162 21148
rect 1226 21084 1252 21148
rect 1316 21084 1342 21148
rect 1406 21084 1432 21148
rect 1496 21084 2700 21148
rect 99 21067 2700 21084
rect 99 21003 982 21067
rect 1046 21003 1072 21067
rect 1136 21003 1162 21067
rect 1226 21003 1252 21067
rect 1316 21003 1342 21067
rect 1406 21003 1432 21067
rect 1496 21003 2700 21067
rect 99 20986 2700 21003
rect 99 20922 982 20986
rect 1046 20922 1072 20986
rect 1136 20922 1162 20986
rect 1226 20922 1252 20986
rect 1316 20922 1342 20986
rect 1406 20922 1432 20986
rect 1496 20925 2700 20986
rect 1496 20922 1531 20925
rect 99 20905 1531 20922
rect 99 20841 982 20905
rect 1046 20841 1072 20905
rect 1136 20841 1162 20905
rect 1226 20841 1252 20905
rect 1316 20841 1342 20905
rect 1406 20841 1432 20905
rect 1496 20861 1531 20905
rect 1595 20861 2700 20925
rect 1496 20841 2700 20861
rect 99 20811 2700 20841
rect 99 20769 1312 20811
rect 99 20705 1141 20769
rect 1205 20747 1312 20769
rect 1376 20747 1401 20811
rect 1465 20747 1491 20811
rect 1555 20747 1581 20811
rect 1645 20747 1671 20811
rect 1735 20747 2700 20811
rect 1205 20705 2700 20747
rect 99 20695 2700 20705
rect 99 20631 1312 20695
rect 1376 20631 1401 20695
rect 1465 20631 1491 20695
rect 1555 20631 1581 20695
rect 1645 20631 1671 20695
rect 1735 20631 2700 20695
rect 99 20617 2700 20631
rect 99 20579 1812 20617
rect 99 20515 1312 20579
rect 1376 20515 1401 20579
rect 1465 20515 1491 20579
rect 1555 20515 1581 20579
rect 1645 20515 1671 20579
rect 1735 20553 1812 20579
rect 1876 20553 2700 20617
rect 1735 20515 2700 20553
rect 99 20491 2700 20515
rect 99 20455 1632 20491
rect 99 20391 1524 20455
rect 1588 20427 1632 20455
rect 1696 20427 1721 20491
rect 1785 20427 1811 20491
rect 1875 20427 1901 20491
rect 1965 20427 1991 20491
rect 2055 20427 2700 20491
rect 1588 20391 2700 20427
rect 99 20375 2700 20391
rect 99 20311 1632 20375
rect 1696 20311 1721 20375
rect 1785 20311 1811 20375
rect 1875 20311 1901 20375
rect 1965 20311 1991 20375
rect 2055 20311 2700 20375
rect 99 20292 2700 20311
rect 99 20259 2137 20292
rect 99 20195 1632 20259
rect 1696 20195 1721 20259
rect 1785 20195 1811 20259
rect 1875 20195 1901 20259
rect 1965 20195 1991 20259
rect 2055 20228 2137 20259
rect 2201 20228 2700 20292
rect 12300 33444 13169 33508
rect 13233 33444 13259 33508
rect 13323 33444 13349 33508
rect 13413 33444 13439 33508
rect 13503 33444 13528 33508
rect 13592 33480 13636 33508
rect 13700 33480 14858 33544
rect 13592 33444 14858 33480
rect 12300 33420 14858 33444
rect 12300 33382 13489 33420
rect 12300 33318 13348 33382
rect 13412 33356 13489 33382
rect 13553 33356 13579 33420
rect 13643 33356 13669 33420
rect 13733 33356 13759 33420
rect 13823 33356 13848 33420
rect 13912 33356 14858 33420
rect 13412 33318 14858 33356
rect 12300 33304 14858 33318
rect 12300 33240 13489 33304
rect 13553 33240 13579 33304
rect 13643 33240 13669 33304
rect 13733 33240 13759 33304
rect 13823 33240 13848 33304
rect 13912 33240 14858 33304
rect 12300 33188 14858 33240
rect 12300 33124 13489 33188
rect 13553 33124 13579 33188
rect 13643 33124 13669 33188
rect 13733 33124 13759 33188
rect 13823 33124 13848 33188
rect 13912 33124 14858 33188
rect 12300 33095 14858 33124
rect 12300 33031 13520 33095
rect 13584 33031 13610 33095
rect 13674 33031 13700 33095
rect 13764 33031 13790 33095
rect 13854 33031 13880 33095
rect 13944 33031 13970 33095
rect 14034 33031 14858 33095
rect 12300 33015 14858 33031
rect 12300 32951 13520 33015
rect 13584 32951 13610 33015
rect 13674 32951 13700 33015
rect 13764 32951 13790 33015
rect 13854 32951 13880 33015
rect 13944 32951 13970 33015
rect 14034 32951 14858 33015
rect 12300 32935 14858 32951
rect 12300 32871 13520 32935
rect 13584 32871 13610 32935
rect 13674 32871 13700 32935
rect 13764 32871 13790 32935
rect 13854 32871 13880 32935
rect 13944 32871 13970 32935
rect 14034 32871 14858 32935
rect 12300 32855 14858 32871
rect 12300 32791 13520 32855
rect 13584 32791 13610 32855
rect 13674 32791 13700 32855
rect 13764 32791 13790 32855
rect 13854 32791 13880 32855
rect 13944 32791 13970 32855
rect 14034 32791 14858 32855
rect 12300 32775 14858 32791
rect 12300 32711 13520 32775
rect 13584 32711 13610 32775
rect 13674 32711 13700 32775
rect 13764 32711 13790 32775
rect 13854 32711 13880 32775
rect 13944 32711 13970 32775
rect 14034 32711 14858 32775
rect 12300 32695 14858 32711
rect 12300 32631 13520 32695
rect 13584 32631 13610 32695
rect 13674 32631 13700 32695
rect 13764 32631 13790 32695
rect 13854 32631 13880 32695
rect 13944 32631 13970 32695
rect 14034 32631 14858 32695
rect 12300 32615 14858 32631
rect 12300 32551 13520 32615
rect 13584 32551 13610 32615
rect 13674 32551 13700 32615
rect 13764 32551 13790 32615
rect 13854 32551 13880 32615
rect 13944 32551 13970 32615
rect 14034 32551 14858 32615
rect 12300 32535 14858 32551
rect 12300 32471 13520 32535
rect 13584 32471 13610 32535
rect 13674 32471 13700 32535
rect 13764 32471 13790 32535
rect 13854 32471 13880 32535
rect 13944 32471 13970 32535
rect 14034 32471 14858 32535
rect 12300 32455 14858 32471
rect 12300 32391 13520 32455
rect 13584 32391 13610 32455
rect 13674 32391 13700 32455
rect 13764 32391 13790 32455
rect 13854 32391 13880 32455
rect 13944 32391 13970 32455
rect 14034 32391 14858 32455
rect 12300 32375 14858 32391
rect 12300 32311 13520 32375
rect 13584 32311 13610 32375
rect 13674 32311 13700 32375
rect 13764 32311 13790 32375
rect 13854 32311 13880 32375
rect 13944 32311 13970 32375
rect 14034 32311 14858 32375
rect 12300 32295 14858 32311
rect 12300 32231 13520 32295
rect 13584 32231 13610 32295
rect 13674 32231 13700 32295
rect 13764 32231 13790 32295
rect 13854 32231 13880 32295
rect 13944 32231 13970 32295
rect 14034 32231 14858 32295
rect 12300 32215 14858 32231
rect 12300 32151 13520 32215
rect 13584 32151 13610 32215
rect 13674 32151 13700 32215
rect 13764 32151 13790 32215
rect 13854 32151 13880 32215
rect 13944 32151 13970 32215
rect 14034 32151 14858 32215
rect 12300 32135 14858 32151
rect 12300 32071 13520 32135
rect 13584 32071 13610 32135
rect 13674 32071 13700 32135
rect 13764 32071 13790 32135
rect 13854 32071 13880 32135
rect 13944 32071 13970 32135
rect 14034 32071 14858 32135
rect 12300 32055 14858 32071
rect 12300 31991 13520 32055
rect 13584 31991 13610 32055
rect 13674 31991 13700 32055
rect 13764 31991 13790 32055
rect 13854 31991 13880 32055
rect 13944 31991 13970 32055
rect 14034 31991 14858 32055
rect 12300 31975 14858 31991
rect 12300 31911 13520 31975
rect 13584 31911 13610 31975
rect 13674 31911 13700 31975
rect 13764 31911 13790 31975
rect 13854 31911 13880 31975
rect 13944 31911 13970 31975
rect 14034 31911 14858 31975
rect 12300 31895 14858 31911
rect 12300 31831 13520 31895
rect 13584 31831 13610 31895
rect 13674 31831 13700 31895
rect 13764 31831 13790 31895
rect 13854 31831 13880 31895
rect 13944 31831 13970 31895
rect 14034 31831 14858 31895
rect 12300 31815 14858 31831
rect 12300 31751 13520 31815
rect 13584 31751 13610 31815
rect 13674 31751 13700 31815
rect 13764 31751 13790 31815
rect 13854 31751 13880 31815
rect 13944 31751 13970 31815
rect 14034 31751 14858 31815
rect 12300 31735 14858 31751
rect 12300 31671 13520 31735
rect 13584 31671 13610 31735
rect 13674 31671 13700 31735
rect 13764 31671 13790 31735
rect 13854 31671 13880 31735
rect 13944 31671 13970 31735
rect 14034 31671 14858 31735
rect 12300 31655 14858 31671
rect 12300 31591 13520 31655
rect 13584 31591 13610 31655
rect 13674 31591 13700 31655
rect 13764 31591 13790 31655
rect 13854 31591 13880 31655
rect 13944 31591 13970 31655
rect 14034 31591 14858 31655
rect 12300 31575 14858 31591
rect 12300 31511 13520 31575
rect 13584 31511 13610 31575
rect 13674 31511 13700 31575
rect 13764 31511 13790 31575
rect 13854 31511 13880 31575
rect 13944 31511 13970 31575
rect 14034 31511 14858 31575
rect 12300 31495 14858 31511
rect 12300 31431 13520 31495
rect 13584 31431 13610 31495
rect 13674 31431 13700 31495
rect 13764 31431 13790 31495
rect 13854 31431 13880 31495
rect 13944 31431 13970 31495
rect 14034 31431 14858 31495
rect 12300 31415 14858 31431
rect 12300 31351 13520 31415
rect 13584 31351 13610 31415
rect 13674 31351 13700 31415
rect 13764 31351 13790 31415
rect 13854 31351 13880 31415
rect 13944 31351 13970 31415
rect 14034 31351 14858 31415
rect 12300 31335 14858 31351
rect 12300 31271 13520 31335
rect 13584 31271 13610 31335
rect 13674 31271 13700 31335
rect 13764 31271 13790 31335
rect 13854 31271 13880 31335
rect 13944 31271 13970 31335
rect 14034 31271 14858 31335
rect 12300 31255 14858 31271
rect 12300 31191 13520 31255
rect 13584 31191 13610 31255
rect 13674 31191 13700 31255
rect 13764 31191 13790 31255
rect 13854 31191 13880 31255
rect 13944 31191 13970 31255
rect 14034 31191 14858 31255
rect 12300 31175 14858 31191
rect 12300 31111 13520 31175
rect 13584 31111 13610 31175
rect 13674 31111 13700 31175
rect 13764 31111 13790 31175
rect 13854 31111 13880 31175
rect 13944 31111 13970 31175
rect 14034 31111 14858 31175
rect 12300 31095 14858 31111
rect 12300 31031 13520 31095
rect 13584 31031 13610 31095
rect 13674 31031 13700 31095
rect 13764 31031 13790 31095
rect 13854 31031 13880 31095
rect 13944 31031 13970 31095
rect 14034 31031 14858 31095
rect 12300 31015 14858 31031
rect 12300 30951 13520 31015
rect 13584 30951 13610 31015
rect 13674 30951 13700 31015
rect 13764 30951 13790 31015
rect 13854 30951 13880 31015
rect 13944 30951 13970 31015
rect 14034 30951 14858 31015
rect 12300 30935 14858 30951
rect 12300 30871 13520 30935
rect 13584 30871 13610 30935
rect 13674 30871 13700 30935
rect 13764 30871 13790 30935
rect 13854 30871 13880 30935
rect 13944 30871 13970 30935
rect 14034 30871 14858 30935
rect 12300 30855 14858 30871
rect 12300 30791 13520 30855
rect 13584 30791 13610 30855
rect 13674 30791 13700 30855
rect 13764 30791 13790 30855
rect 13854 30791 13880 30855
rect 13944 30791 13970 30855
rect 14034 30791 14858 30855
rect 12300 30775 14858 30791
rect 12300 30711 13520 30775
rect 13584 30711 13610 30775
rect 13674 30711 13700 30775
rect 13764 30711 13790 30775
rect 13854 30711 13880 30775
rect 13944 30711 13970 30775
rect 14034 30711 14858 30775
rect 12300 30695 14858 30711
rect 12300 30631 13520 30695
rect 13584 30631 13610 30695
rect 13674 30631 13700 30695
rect 13764 30631 13790 30695
rect 13854 30631 13880 30695
rect 13944 30631 13970 30695
rect 14034 30631 14858 30695
rect 12300 30615 14858 30631
rect 12300 30551 13520 30615
rect 13584 30551 13610 30615
rect 13674 30551 13700 30615
rect 13764 30551 13790 30615
rect 13854 30551 13880 30615
rect 13944 30551 13970 30615
rect 14034 30551 14858 30615
rect 12300 30535 14858 30551
rect 12300 30471 13520 30535
rect 13584 30471 13610 30535
rect 13674 30471 13700 30535
rect 13764 30471 13790 30535
rect 13854 30471 13880 30535
rect 13944 30471 13970 30535
rect 14034 30471 14858 30535
rect 12300 30455 14858 30471
rect 12300 30391 13520 30455
rect 13584 30391 13610 30455
rect 13674 30391 13700 30455
rect 13764 30391 13790 30455
rect 13854 30391 13880 30455
rect 13944 30391 13970 30455
rect 14034 30391 14858 30455
rect 12300 30375 14858 30391
rect 12300 30311 13520 30375
rect 13584 30311 13610 30375
rect 13674 30311 13700 30375
rect 13764 30311 13790 30375
rect 13854 30311 13880 30375
rect 13944 30311 13970 30375
rect 14034 30311 14858 30375
rect 12300 30295 14858 30311
rect 12300 30231 13520 30295
rect 13584 30231 13610 30295
rect 13674 30231 13700 30295
rect 13764 30231 13790 30295
rect 13854 30231 13880 30295
rect 13944 30231 13970 30295
rect 14034 30231 14858 30295
rect 12300 30215 14858 30231
rect 12300 30151 13520 30215
rect 13584 30151 13610 30215
rect 13674 30151 13700 30215
rect 13764 30151 13790 30215
rect 13854 30151 13880 30215
rect 13944 30151 13970 30215
rect 14034 30151 14858 30215
rect 12300 30135 14858 30151
rect 12300 30071 13520 30135
rect 13584 30071 13610 30135
rect 13674 30071 13700 30135
rect 13764 30071 13790 30135
rect 13854 30071 13880 30135
rect 13944 30071 13970 30135
rect 14034 30071 14858 30135
rect 12300 30055 14858 30071
rect 12300 29991 13520 30055
rect 13584 29991 13610 30055
rect 13674 29991 13700 30055
rect 13764 29991 13790 30055
rect 13854 29991 13880 30055
rect 13944 29991 13970 30055
rect 14034 29991 14858 30055
rect 12300 29975 14858 29991
rect 12300 29911 13520 29975
rect 13584 29911 13610 29975
rect 13674 29911 13700 29975
rect 13764 29911 13790 29975
rect 13854 29911 13880 29975
rect 13944 29911 13970 29975
rect 14034 29911 14858 29975
rect 12300 29895 14858 29911
rect 12300 29831 13520 29895
rect 13584 29831 13610 29895
rect 13674 29831 13700 29895
rect 13764 29831 13790 29895
rect 13854 29831 13880 29895
rect 13944 29831 13970 29895
rect 14034 29831 14858 29895
rect 12300 29815 14858 29831
rect 12300 29751 13520 29815
rect 13584 29751 13610 29815
rect 13674 29751 13700 29815
rect 13764 29751 13790 29815
rect 13854 29751 13880 29815
rect 13944 29751 13970 29815
rect 14034 29751 14858 29815
rect 12300 29735 14858 29751
rect 12300 29671 13520 29735
rect 13584 29671 13610 29735
rect 13674 29671 13700 29735
rect 13764 29671 13790 29735
rect 13854 29671 13880 29735
rect 13944 29671 13970 29735
rect 14034 29671 14858 29735
rect 12300 29655 14858 29671
rect 12300 29591 13520 29655
rect 13584 29591 13610 29655
rect 13674 29591 13700 29655
rect 13764 29591 13790 29655
rect 13854 29591 13880 29655
rect 13944 29591 13970 29655
rect 14034 29591 14858 29655
rect 12300 29575 14858 29591
rect 12300 29511 13520 29575
rect 13584 29511 13610 29575
rect 13674 29511 13700 29575
rect 13764 29511 13790 29575
rect 13854 29511 13880 29575
rect 13944 29511 13970 29575
rect 14034 29511 14858 29575
rect 12300 29495 14858 29511
rect 12300 29431 13520 29495
rect 13584 29431 13610 29495
rect 13674 29431 13700 29495
rect 13764 29431 13790 29495
rect 13854 29431 13880 29495
rect 13944 29431 13970 29495
rect 14034 29431 14858 29495
rect 12300 29415 14858 29431
rect 12300 29351 13520 29415
rect 13584 29351 13610 29415
rect 13674 29351 13700 29415
rect 13764 29351 13790 29415
rect 13854 29351 13880 29415
rect 13944 29351 13970 29415
rect 14034 29351 14858 29415
rect 12300 29335 14858 29351
rect 12300 29271 13520 29335
rect 13584 29271 13610 29335
rect 13674 29271 13700 29335
rect 13764 29271 13790 29335
rect 13854 29271 13880 29335
rect 13944 29271 13970 29335
rect 14034 29271 14858 29335
rect 12300 29255 14858 29271
rect 12300 29191 13520 29255
rect 13584 29191 13610 29255
rect 13674 29191 13700 29255
rect 13764 29191 13790 29255
rect 13854 29191 13880 29255
rect 13944 29191 13970 29255
rect 14034 29191 14858 29255
rect 12300 29175 14858 29191
rect 12300 29111 13520 29175
rect 13584 29111 13610 29175
rect 13674 29111 13700 29175
rect 13764 29111 13790 29175
rect 13854 29111 13880 29175
rect 13944 29111 13970 29175
rect 14034 29111 14858 29175
rect 12300 29095 14858 29111
rect 12300 29031 13520 29095
rect 13584 29031 13610 29095
rect 13674 29031 13700 29095
rect 13764 29031 13790 29095
rect 13854 29031 13880 29095
rect 13944 29031 13970 29095
rect 14034 29031 14858 29095
rect 12300 29015 14858 29031
rect 12300 28951 13520 29015
rect 13584 28951 13610 29015
rect 13674 28951 13700 29015
rect 13764 28951 13790 29015
rect 13854 28951 13880 29015
rect 13944 28951 13970 29015
rect 14034 28951 14858 29015
rect 12300 28935 14858 28951
rect 12300 28917 13520 28935
rect 13584 28917 13610 28935
rect 13674 28917 13700 28935
rect 13764 28917 13790 28935
rect 13854 28917 13880 28935
rect 13944 28917 13970 28935
rect 14034 28917 14858 28935
rect 12300 23341 12455 28917
rect 14431 23341 14858 28917
rect 12300 23335 14858 23341
rect 12300 23271 13520 23335
rect 13584 23271 13610 23335
rect 13674 23271 13700 23335
rect 13764 23271 13790 23335
rect 13854 23271 13880 23335
rect 13944 23271 13970 23335
rect 14034 23271 14858 23335
rect 12300 23254 14858 23271
rect 12300 23190 13520 23254
rect 13584 23190 13610 23254
rect 13674 23190 13700 23254
rect 13764 23190 13790 23254
rect 13854 23190 13880 23254
rect 13944 23190 13970 23254
rect 14034 23190 14858 23254
rect 12300 23173 14858 23190
rect 12300 23109 13520 23173
rect 13584 23109 13610 23173
rect 13674 23109 13700 23173
rect 13764 23109 13790 23173
rect 13854 23109 13880 23173
rect 13944 23109 13970 23173
rect 14034 23109 14858 23173
rect 12300 23092 14858 23109
rect 12300 23028 13520 23092
rect 13584 23028 13610 23092
rect 13674 23028 13700 23092
rect 13764 23028 13790 23092
rect 13854 23028 13880 23092
rect 13944 23028 13970 23092
rect 14034 23028 14858 23092
rect 12300 23011 14858 23028
rect 12300 22947 13520 23011
rect 13584 22947 13610 23011
rect 13674 22947 13700 23011
rect 13764 22947 13790 23011
rect 13854 22947 13880 23011
rect 13944 22947 13970 23011
rect 14034 22947 14858 23011
rect 12300 22930 14858 22947
rect 12300 22866 13520 22930
rect 13584 22866 13610 22930
rect 13674 22866 13700 22930
rect 13764 22866 13790 22930
rect 13854 22866 13880 22930
rect 13944 22866 13970 22930
rect 14034 22866 14858 22930
rect 12300 22849 14858 22866
rect 12300 22785 13520 22849
rect 13584 22785 13610 22849
rect 13674 22785 13700 22849
rect 13764 22785 13790 22849
rect 13854 22785 13880 22849
rect 13944 22785 13970 22849
rect 14034 22785 14858 22849
rect 12300 22768 14858 22785
rect 12300 22704 13520 22768
rect 13584 22704 13610 22768
rect 13674 22704 13700 22768
rect 13764 22704 13790 22768
rect 13854 22704 13880 22768
rect 13944 22704 13970 22768
rect 14034 22704 14858 22768
rect 12300 22687 14858 22704
rect 12300 22623 13520 22687
rect 13584 22623 13610 22687
rect 13674 22623 13700 22687
rect 13764 22623 13790 22687
rect 13854 22623 13880 22687
rect 13944 22623 13970 22687
rect 14034 22623 14858 22687
rect 12300 22606 14858 22623
rect 12300 22542 13520 22606
rect 13584 22542 13610 22606
rect 13674 22542 13700 22606
rect 13764 22542 13790 22606
rect 13854 22542 13880 22606
rect 13944 22542 13970 22606
rect 14034 22542 14858 22606
rect 12300 22525 14858 22542
rect 12300 22461 13520 22525
rect 13584 22461 13610 22525
rect 13674 22461 13700 22525
rect 13764 22461 13790 22525
rect 13854 22461 13880 22525
rect 13944 22461 13970 22525
rect 14034 22461 14858 22525
rect 12300 22444 14858 22461
rect 12300 22380 13520 22444
rect 13584 22380 13610 22444
rect 13674 22380 13700 22444
rect 13764 22380 13790 22444
rect 13854 22380 13880 22444
rect 13944 22380 13970 22444
rect 14034 22380 14858 22444
rect 12300 22363 14858 22380
rect 12300 22299 13520 22363
rect 13584 22299 13610 22363
rect 13674 22299 13700 22363
rect 13764 22299 13790 22363
rect 13854 22299 13880 22363
rect 13944 22299 13970 22363
rect 14034 22299 14858 22363
rect 12300 22282 14858 22299
rect 12300 22218 13520 22282
rect 13584 22218 13610 22282
rect 13674 22218 13700 22282
rect 13764 22218 13790 22282
rect 13854 22218 13880 22282
rect 13944 22218 13970 22282
rect 14034 22218 14858 22282
rect 12300 22201 14858 22218
rect 12300 22137 13520 22201
rect 13584 22137 13610 22201
rect 13674 22137 13700 22201
rect 13764 22137 13790 22201
rect 13854 22137 13880 22201
rect 13944 22137 13970 22201
rect 14034 22137 14858 22201
rect 12300 22120 14858 22137
rect 12300 22056 13520 22120
rect 13584 22056 13610 22120
rect 13674 22056 13700 22120
rect 13764 22056 13790 22120
rect 13854 22056 13880 22120
rect 13944 22056 13970 22120
rect 14034 22056 14858 22120
rect 12300 22039 14858 22056
rect 12300 21975 13520 22039
rect 13584 21975 13610 22039
rect 13674 21975 13700 22039
rect 13764 21975 13790 22039
rect 13854 21975 13880 22039
rect 13944 21975 13970 22039
rect 14034 21975 14858 22039
rect 12300 21958 14858 21975
rect 12300 21894 13520 21958
rect 13584 21894 13610 21958
rect 13674 21894 13700 21958
rect 13764 21894 13790 21958
rect 13854 21894 13880 21958
rect 13944 21894 13970 21958
rect 14034 21894 14858 21958
rect 12300 21877 14858 21894
rect 12300 21813 13520 21877
rect 13584 21813 13610 21877
rect 13674 21813 13700 21877
rect 13764 21813 13790 21877
rect 13854 21813 13880 21877
rect 13944 21813 13970 21877
rect 14034 21813 14858 21877
rect 12300 21796 14858 21813
rect 12300 21732 13520 21796
rect 13584 21732 13610 21796
rect 13674 21732 13700 21796
rect 13764 21732 13790 21796
rect 13854 21732 13880 21796
rect 13944 21732 13970 21796
rect 14034 21732 14858 21796
rect 12300 21715 14858 21732
rect 12300 21651 13520 21715
rect 13584 21651 13610 21715
rect 13674 21651 13700 21715
rect 13764 21651 13790 21715
rect 13854 21651 13880 21715
rect 13944 21651 13970 21715
rect 14034 21651 14858 21715
rect 12300 21634 14858 21651
rect 12300 21570 13520 21634
rect 13584 21570 13610 21634
rect 13674 21570 13700 21634
rect 13764 21570 13790 21634
rect 13854 21570 13880 21634
rect 13944 21570 13970 21634
rect 14034 21570 14858 21634
rect 12300 21553 14858 21570
rect 12300 21489 13520 21553
rect 13584 21489 13610 21553
rect 13674 21489 13700 21553
rect 13764 21489 13790 21553
rect 13854 21489 13880 21553
rect 13944 21489 13970 21553
rect 14034 21489 14858 21553
rect 12300 21472 14858 21489
rect 12300 21408 13520 21472
rect 13584 21408 13610 21472
rect 13674 21408 13700 21472
rect 13764 21408 13790 21472
rect 13854 21408 13880 21472
rect 13944 21408 13970 21472
rect 14034 21408 14858 21472
rect 12300 21391 14858 21408
rect 12300 21327 13520 21391
rect 13584 21327 13610 21391
rect 13674 21327 13700 21391
rect 13764 21327 13790 21391
rect 13854 21327 13880 21391
rect 13944 21327 13970 21391
rect 14034 21327 14858 21391
rect 12300 21310 14858 21327
rect 12300 21246 13520 21310
rect 13584 21246 13610 21310
rect 13674 21246 13700 21310
rect 13764 21246 13790 21310
rect 13854 21246 13880 21310
rect 13944 21246 13970 21310
rect 14034 21246 14858 21310
rect 12300 21229 14858 21246
rect 12300 21165 13520 21229
rect 13584 21165 13610 21229
rect 13674 21165 13700 21229
rect 13764 21165 13790 21229
rect 13854 21165 13880 21229
rect 13944 21165 13970 21229
rect 14034 21165 14858 21229
rect 12300 21148 14858 21165
rect 12300 21084 13520 21148
rect 13584 21084 13610 21148
rect 13674 21084 13700 21148
rect 13764 21084 13790 21148
rect 13854 21084 13880 21148
rect 13944 21084 13970 21148
rect 14034 21084 14858 21148
rect 12300 21067 14858 21084
rect 12300 21003 13520 21067
rect 13584 21003 13610 21067
rect 13674 21003 13700 21067
rect 13764 21003 13790 21067
rect 13854 21003 13880 21067
rect 13944 21003 13970 21067
rect 14034 21003 14858 21067
rect 12300 20986 14858 21003
rect 12300 20925 13520 20986
rect 12300 20861 13421 20925
rect 13485 20922 13520 20925
rect 13584 20922 13610 20986
rect 13674 20922 13700 20986
rect 13764 20922 13790 20986
rect 13854 20922 13880 20986
rect 13944 20922 13970 20986
rect 14034 20922 14858 20986
rect 13485 20905 14858 20922
rect 13485 20861 13520 20905
rect 12300 20841 13520 20861
rect 13584 20841 13610 20905
rect 13674 20841 13700 20905
rect 13764 20841 13790 20905
rect 13854 20841 13880 20905
rect 13944 20841 13970 20905
rect 14034 20841 14858 20905
rect 12300 20811 14858 20841
rect 12300 20747 13281 20811
rect 13345 20747 13371 20811
rect 13435 20747 13461 20811
rect 13525 20747 13551 20811
rect 13615 20747 13640 20811
rect 13704 20809 14858 20811
rect 13704 20747 13749 20809
rect 12300 20745 13749 20747
rect 13813 20802 14858 20809
rect 13813 20745 13851 20802
rect 12300 20738 13851 20745
rect 13915 20738 14858 20802
rect 12300 20698 14858 20738
rect 12300 20695 13749 20698
rect 12300 20631 13281 20695
rect 13345 20631 13371 20695
rect 13435 20631 13461 20695
rect 13525 20631 13551 20695
rect 13615 20631 13640 20695
rect 13704 20634 13749 20695
rect 13813 20634 14858 20698
rect 13704 20631 14858 20634
rect 12300 20617 14858 20631
rect 12300 20553 13140 20617
rect 13204 20579 14858 20617
rect 13204 20553 13281 20579
rect 12300 20515 13281 20553
rect 13345 20515 13371 20579
rect 13435 20515 13461 20579
rect 13525 20515 13551 20579
rect 13615 20515 13640 20579
rect 13704 20515 14858 20579
rect 12300 20491 14858 20515
rect 12300 20427 12961 20491
rect 13025 20427 13051 20491
rect 13115 20427 13141 20491
rect 13205 20427 13231 20491
rect 13295 20427 13320 20491
rect 13384 20455 14858 20491
rect 13384 20427 13428 20455
rect 12300 20391 13428 20427
rect 13492 20391 14858 20455
rect 12300 20375 14858 20391
rect 12300 20311 12961 20375
rect 13025 20311 13051 20375
rect 13115 20311 13141 20375
rect 13205 20311 13231 20375
rect 13295 20311 13320 20375
rect 13384 20311 14858 20375
rect 12300 20292 14858 20311
rect 2055 20195 2700 20228
rect 99 20167 2700 20195
rect 99 20127 1956 20167
rect 99 20063 1852 20127
rect 1916 20103 1956 20127
rect 2020 20103 2045 20167
rect 2109 20103 2135 20167
rect 2199 20103 2225 20167
rect 2289 20103 2315 20167
rect 2379 20103 2700 20167
rect 1916 20063 2700 20103
rect 99 20056 2700 20063
tri 2700 20056 2923 20279 sw
tri 12110 20069 12300 20259 se
rect 12300 20228 12815 20292
rect 12879 20259 14858 20292
rect 12879 20228 12961 20259
rect 12300 20195 12961 20228
rect 13025 20195 13051 20259
rect 13115 20195 13141 20259
rect 13205 20195 13231 20259
rect 13295 20195 13320 20259
rect 13384 20195 14858 20259
rect 12300 20167 14858 20195
rect 12300 20103 12637 20167
rect 12701 20103 12727 20167
rect 12791 20103 12817 20167
rect 12881 20103 12907 20167
rect 12971 20103 12996 20167
rect 13060 20127 14858 20167
rect 13060 20103 13100 20127
rect 12300 20069 13100 20103
tri 12097 20056 12110 20069 se
rect 12110 20063 13100 20069
rect 13164 20063 14858 20127
rect 12110 20056 14858 20063
rect 99 20051 2456 20056
rect 99 19987 1956 20051
rect 2020 19987 2045 20051
rect 2109 19987 2135 20051
rect 2199 19987 2225 20051
rect 2289 19987 2315 20051
rect 2379 19992 2456 20051
rect 2520 19992 2571 20056
rect 2635 19992 2686 20056
rect 2750 19992 2802 20056
rect 2866 19992 2923 20056
rect 2379 19987 2923 19992
rect 99 19941 2923 19987
tri 2923 19941 3038 20056 sw
tri 12027 19986 12097 20056 se
rect 12097 19992 12150 20056
rect 12214 19992 12266 20056
rect 12330 19992 12381 20056
rect 12445 19992 12496 20056
rect 12560 20051 14858 20056
rect 12560 19992 12637 20051
rect 12097 19987 12637 19992
rect 12701 19987 12727 20051
rect 12791 19987 12817 20051
rect 12881 19987 12907 20051
rect 12971 19987 12996 20051
rect 13060 19987 14858 20051
rect 12097 19986 14858 19987
tri 11982 19941 12027 19986 se
rect 12027 19941 14858 19986
rect 99 19936 2906 19941
rect 99 19935 2456 19936
rect 99 19871 1956 19935
rect 2020 19871 2045 19935
rect 2109 19871 2135 19935
rect 2199 19871 2225 19935
rect 2289 19871 2315 19935
rect 2379 19872 2456 19935
rect 2520 19872 2571 19936
rect 2635 19872 2686 19936
rect 2750 19872 2802 19936
rect 2866 19877 2906 19936
rect 2970 19877 3038 19941
rect 2866 19872 3038 19877
rect 2379 19871 3038 19872
rect 99 19830 3038 19871
tri 3038 19830 3149 19941 sw
tri 11885 19844 11982 19941 se
rect 11982 19877 12046 19941
rect 12110 19936 14858 19941
rect 12110 19877 12150 19936
rect 11982 19872 12150 19877
rect 12214 19872 12266 19936
rect 12330 19872 12381 19936
rect 12445 19872 12496 19936
rect 12560 19935 14858 19936
rect 12560 19872 12637 19935
rect 11982 19871 12637 19872
rect 12701 19871 12727 19935
rect 12791 19871 12817 19935
rect 12881 19871 12907 19935
rect 12971 19871 12996 19935
rect 13060 19871 14858 19935
rect 11982 19844 14858 19871
tri 11871 19830 11885 19844 se
rect 11885 19830 14858 19844
rect 99 19786 2293 19830
rect 99 19722 2193 19786
rect 2257 19766 2293 19786
rect 2357 19766 2377 19830
rect 2441 19766 2461 19830
rect 2525 19766 2545 19830
rect 2609 19766 2629 19830
rect 2693 19766 2713 19830
rect 2777 19766 2797 19830
rect 2861 19766 2881 19830
rect 2945 19766 2965 19830
rect 3029 19766 3049 19830
rect 3113 19766 3149 19830
rect 2257 19722 3149 19766
rect 99 19714 3149 19722
rect 99 19650 2293 19714
rect 2357 19650 2377 19714
rect 2441 19650 2461 19714
rect 2525 19650 2545 19714
rect 2609 19650 2629 19714
rect 2693 19650 2713 19714
rect 2777 19650 2797 19714
rect 2861 19650 2881 19714
rect 2945 19650 2965 19714
rect 3029 19650 3049 19714
rect 3113 19693 3149 19714
tri 3149 19693 3286 19830 sw
tri 11753 19712 11871 19830 se
rect 11871 19766 11903 19830
rect 11967 19766 11987 19830
rect 12051 19766 12071 19830
rect 12135 19766 12155 19830
rect 12219 19766 12239 19830
rect 12303 19766 12323 19830
rect 12387 19766 12407 19830
rect 12471 19766 12491 19830
rect 12555 19766 12575 19830
rect 12639 19766 12659 19830
rect 12723 19786 14858 19830
rect 12723 19766 12759 19786
rect 11871 19722 12759 19766
rect 12823 19722 14858 19786
rect 11871 19714 14858 19722
rect 11871 19712 11903 19714
tri 11734 19693 11753 19712 se
rect 11753 19693 11903 19712
rect 3113 19650 3153 19693
rect 99 19629 3153 19650
rect 3217 19629 3286 19693
rect 99 19600 3286 19629
rect 99 19598 3153 19600
rect 99 19534 2293 19598
rect 2357 19534 2377 19598
rect 2441 19534 2461 19598
rect 2525 19534 2545 19598
rect 2609 19534 2629 19598
rect 2693 19534 2713 19598
rect 2777 19534 2797 19598
rect 2861 19534 2881 19598
rect 2945 19534 2965 19598
rect 3029 19534 3049 19598
rect 3113 19536 3153 19598
rect 3217 19536 3286 19600
rect 3113 19534 3286 19536
rect 99 19524 3286 19534
tri 99 18934 689 19524 ne
rect 689 18934 3286 19524
tri 3286 18934 4045 19693 sw
tri 11237 19196 11734 19693 se
rect 11734 19629 11799 19693
rect 11863 19650 11903 19693
rect 11967 19650 11987 19714
rect 12051 19650 12071 19714
rect 12135 19650 12155 19714
rect 12219 19650 12239 19714
rect 12303 19650 12323 19714
rect 12387 19650 12407 19714
rect 12471 19650 12491 19714
rect 12555 19650 12575 19714
rect 12639 19650 12659 19714
rect 12723 19650 14858 19714
rect 11863 19629 14858 19650
rect 11734 19600 14858 19629
rect 11734 19536 11799 19600
rect 11863 19598 14858 19600
rect 11863 19536 11903 19598
rect 11734 19534 11903 19536
rect 11967 19534 11987 19598
rect 12051 19534 12071 19598
rect 12135 19534 12155 19598
rect 12219 19534 12239 19598
rect 12303 19534 12323 19598
rect 12387 19534 12407 19598
rect 12471 19534 12491 19598
rect 12555 19534 12575 19598
rect 12639 19534 12659 19598
rect 12723 19574 14858 19598
rect 12723 19534 14696 19574
rect 11734 19412 14696 19534
tri 14696 19412 14858 19574 nw
rect 11734 19196 12260 19412
tri 4842 18996 5042 19196 se
rect 5042 18996 9935 19196
tri 9935 18996 10135 19196 sw
tri 689 18931 692 18934 ne
rect 692 18931 4045 18934
tri 4045 18931 4048 18934 sw
rect 4842 18931 10135 18996
tri 692 17275 2348 18931 ne
rect 2348 18871 4048 18931
tri 4048 18871 4108 18931 sw
rect 2348 17275 4108 18871
tri 2348 17273 2350 17275 ne
rect 2350 17273 4108 17275
tri 2350 17231 2392 17273 ne
rect 2392 17231 4108 17273
tri 2392 17214 2409 17231 ne
rect 2409 17214 4108 17231
rect 4842 18895 4942 18931
rect 7238 18895 7742 18931
rect 10038 18895 10135 18931
rect 4842 17311 4938 18895
rect 7242 17311 7738 18895
rect 10042 17311 10135 18895
rect 4842 17275 4942 17311
rect 7238 17275 7742 17311
rect 10038 17275 10135 17311
rect 4842 17230 10135 17275
tri 4842 17214 4858 17230 ne
rect 4858 17218 9935 17230
rect 4858 17214 5099 17218
tri 2409 17078 2545 17214 ne
rect 2545 17078 4108 17214
tri 4858 17078 4994 17214 ne
rect 4994 17078 5099 17214
tri 2545 17061 2562 17078 ne
rect 2562 17061 4108 17078
tri 4994 17071 5001 17078 ne
rect 5001 17074 5099 17078
rect 7243 17074 7735 17218
rect 9879 17074 9935 17218
rect 5001 17071 9935 17074
tri 4108 17061 4118 17071 sw
tri 5001 17061 5011 17071 ne
rect 5011 17061 9935 17071
tri 2562 16924 2699 17061 ne
rect 2699 16924 4118 17061
tri 2699 15671 3952 16924 ne
rect 3952 16471 4118 16924
tri 4118 16471 4708 17061 sw
tri 5011 17030 5042 17061 ne
rect 5042 17030 9935 17061
tri 9935 17030 10135 17230 nw
tri 10912 18871 11237 19196 se
rect 11237 18871 12260 19196
tri 10872 17030 10912 17070 se
rect 10912 17030 12260 18871
tri 10313 16471 10872 17030 se
rect 10872 16976 12260 17030
tri 12260 16976 14696 19412 nw
rect 10872 16974 12258 16976
rect 10872 16572 11858 16974
tri 11858 16574 12258 16974 nw
rect 10872 16471 10955 16572
rect 3952 15671 4708 16471
tri 4708 15671 5508 16471 sw
tri 9513 15671 10313 16471 se
rect 10313 15671 10955 16471
tri 3952 14871 4752 15671 ne
rect 4752 14871 5508 15671
tri 5508 14871 6308 15671 sw
tri 8713 14871 9513 15671 se
rect 9513 15669 10955 15671
tri 10955 15669 11858 16572 nw
rect 9513 14871 10157 15669
tri 10157 14871 10955 15669 nw
tri 4752 14071 5552 14871 ne
rect 5552 14071 6308 14871
tri 6308 14071 7108 14871 sw
tri 7913 14071 8713 14871 se
rect 8713 14071 9357 14871
tri 9357 14071 10157 14871 nw
tri 5552 12871 6752 14071 ne
rect 6752 12870 8156 14071
tri 8156 12870 9357 14071 nw
rect 858 9741 2098 9774
rect 858 9285 890 9741
rect 2066 9285 2098 9741
rect 858 4811 2098 9285
rect 2396 9501 3635 9528
rect 2396 8965 2427 9501
rect 3603 8965 3635 9501
rect 2396 6025 3635 8965
rect 2396 5241 2423 6025
rect 3607 5241 3635 6025
rect 2396 5122 3635 5241
rect 858 4027 887 4811
rect 2071 4027 2098 4811
rect 858 3955 2098 4027
rect 6752 1 8153 12870
rect 12858 9741 14098 9774
rect 11273 9502 12512 9529
rect 11273 8966 11304 9502
rect 12480 8966 12512 9502
rect 11273 6024 12512 8966
rect 11273 5240 11297 6024
rect 12481 5240 12512 6024
rect 11273 5122 12512 5240
rect 12858 9285 12890 9741
rect 14066 9285 14098 9741
rect 12858 4811 14098 9285
rect 12858 4027 12887 4811
rect 14071 4027 14098 4811
rect 12858 3955 14098 4027
<< via3 >>
rect 4975 39213 7199 39217
rect 4975 35317 4979 39213
rect 4979 35317 7195 39213
rect 7195 35317 7199 39213
rect 4975 35313 7199 35317
rect 7775 39213 9999 39217
rect 7775 35317 7779 39213
rect 7779 35317 9995 39213
rect 9995 35317 9999 39213
rect 7775 35313 9999 35317
rect 2276 34540 2340 34604
rect 2359 34540 2423 34604
rect 2443 34540 2507 34604
rect 2527 34540 2591 34604
rect 2611 34540 2675 34604
rect 2276 34446 2340 34510
rect 2359 34446 2423 34510
rect 2443 34446 2507 34510
rect 2527 34446 2591 34510
rect 2611 34446 2675 34510
rect 2148 34363 2212 34427
rect 2276 34352 2340 34416
rect 2359 34352 2423 34416
rect 2443 34352 2507 34416
rect 2527 34352 2591 34416
rect 2611 34352 2675 34416
rect 2004 34238 2068 34302
rect 2084 34238 2148 34302
rect 2164 34238 2228 34302
rect 2276 34258 2340 34322
rect 2359 34258 2423 34322
rect 2443 34258 2507 34322
rect 2527 34258 2591 34322
rect 2611 34258 2675 34322
rect 1890 34105 1954 34169
rect 2004 34142 2068 34206
rect 2084 34142 2148 34206
rect 2164 34142 2228 34206
rect 2276 34164 2340 34228
rect 2359 34164 2423 34228
rect 2443 34164 2507 34228
rect 2527 34164 2591 34228
rect 2611 34164 2675 34228
rect 2276 34070 2340 34134
rect 2359 34070 2423 34134
rect 2443 34070 2507 34134
rect 2527 34070 2591 34134
rect 2611 34070 2675 34134
rect 1748 34000 1812 34064
rect 1837 34000 1901 34064
rect 1927 34000 1991 34064
rect 2017 34000 2081 34064
rect 2107 34000 2171 34064
rect 1748 33884 1812 33948
rect 1837 33884 1901 33948
rect 1927 33884 1991 33948
rect 2017 33884 2081 33948
rect 2107 33884 2171 33948
rect 2247 33931 2311 33995
rect 1644 33808 1708 33872
rect 1748 33768 1812 33832
rect 1837 33768 1901 33832
rect 1927 33768 1991 33832
rect 2017 33768 2081 33832
rect 2107 33768 2171 33832
rect 1424 33676 1488 33740
rect 1513 33676 1577 33740
rect 1603 33676 1667 33740
rect 1693 33676 1757 33740
rect 1783 33676 1847 33740
rect 1929 33643 1993 33707
rect 1424 33560 1488 33624
rect 1513 33560 1577 33624
rect 1603 33560 1667 33624
rect 1693 33560 1757 33624
rect 1783 33560 1847 33624
rect 1316 33480 1380 33544
rect 1424 33444 1488 33508
rect 1513 33444 1577 33508
rect 1603 33444 1667 33508
rect 1693 33444 1757 33508
rect 1783 33444 1847 33508
rect 12341 34540 12405 34604
rect 12425 34540 12489 34604
rect 12509 34540 12573 34604
rect 12593 34540 12657 34604
rect 12677 34540 12741 34604
rect 12341 34446 12405 34510
rect 12425 34446 12489 34510
rect 12509 34446 12573 34510
rect 12593 34446 12657 34510
rect 12677 34446 12741 34510
rect 12341 34352 12405 34416
rect 12425 34352 12489 34416
rect 12509 34352 12573 34416
rect 12593 34352 12657 34416
rect 12677 34352 12741 34416
rect 12804 34363 12868 34427
rect 12341 34258 12405 34322
rect 12425 34258 12489 34322
rect 12509 34258 12573 34322
rect 12593 34258 12657 34322
rect 12677 34258 12741 34322
rect 12788 34238 12852 34302
rect 12868 34238 12932 34302
rect 12948 34238 13012 34302
rect 12341 34164 12405 34228
rect 12425 34164 12489 34228
rect 12509 34164 12573 34228
rect 12593 34164 12657 34228
rect 12677 34164 12741 34228
rect 12788 34142 12852 34206
rect 12868 34142 12932 34206
rect 12948 34142 13012 34206
rect 12341 34070 12405 34134
rect 12425 34070 12489 34134
rect 12509 34070 12573 34134
rect 12593 34070 12657 34134
rect 12677 34070 12741 34134
rect 13062 34105 13126 34169
rect 12845 34000 12909 34064
rect 12935 34000 12999 34064
rect 13025 34000 13089 34064
rect 13115 34000 13179 34064
rect 13204 34000 13268 34064
rect 12705 33931 12769 33995
rect 12845 33884 12909 33948
rect 12935 33884 12999 33948
rect 13025 33884 13089 33948
rect 13115 33884 13179 33948
rect 13204 33884 13268 33948
rect 12845 33768 12909 33832
rect 12935 33768 12999 33832
rect 13025 33768 13089 33832
rect 13115 33768 13179 33832
rect 13204 33768 13268 33832
rect 13308 33808 13372 33872
rect 13023 33643 13087 33707
rect 13169 33676 13233 33740
rect 13259 33676 13323 33740
rect 13349 33676 13413 33740
rect 13439 33676 13503 33740
rect 13528 33676 13592 33740
rect 13169 33560 13233 33624
rect 13259 33560 13323 33624
rect 13349 33560 13413 33624
rect 13439 33560 13503 33624
rect 13528 33560 13592 33624
rect 1104 33356 1168 33420
rect 1193 33356 1257 33420
rect 1283 33356 1347 33420
rect 1373 33356 1437 33420
rect 1463 33356 1527 33420
rect 1604 33318 1668 33382
rect 1104 33240 1168 33304
rect 1193 33240 1257 33304
rect 1283 33240 1347 33304
rect 1373 33240 1437 33304
rect 1463 33240 1527 33304
rect 1104 33124 1168 33188
rect 1193 33124 1257 33188
rect 1283 33124 1347 33188
rect 1373 33124 1437 33188
rect 1463 33124 1527 33188
rect 982 33031 1046 33095
rect 1072 33031 1136 33095
rect 1162 33031 1226 33095
rect 1252 33031 1316 33095
rect 1342 33031 1406 33095
rect 1432 33031 1496 33095
rect 982 32951 1046 33015
rect 1072 32951 1136 33015
rect 1162 32951 1226 33015
rect 1252 32951 1316 33015
rect 1342 32951 1406 33015
rect 1432 32951 1496 33015
rect 982 32871 1046 32935
rect 1072 32871 1136 32935
rect 1162 32871 1226 32935
rect 1252 32871 1316 32935
rect 1342 32871 1406 32935
rect 1432 32871 1496 32935
rect 982 32791 1046 32855
rect 1072 32791 1136 32855
rect 1162 32791 1226 32855
rect 1252 32791 1316 32855
rect 1342 32791 1406 32855
rect 1432 32791 1496 32855
rect 982 32711 1046 32775
rect 1072 32711 1136 32775
rect 1162 32711 1226 32775
rect 1252 32711 1316 32775
rect 1342 32711 1406 32775
rect 1432 32711 1496 32775
rect 982 32631 1046 32695
rect 1072 32631 1136 32695
rect 1162 32631 1226 32695
rect 1252 32631 1316 32695
rect 1342 32631 1406 32695
rect 1432 32631 1496 32695
rect 982 32551 1046 32615
rect 1072 32551 1136 32615
rect 1162 32551 1226 32615
rect 1252 32551 1316 32615
rect 1342 32551 1406 32615
rect 1432 32551 1496 32615
rect 982 32471 1046 32535
rect 1072 32471 1136 32535
rect 1162 32471 1226 32535
rect 1252 32471 1316 32535
rect 1342 32471 1406 32535
rect 1432 32471 1496 32535
rect 982 32391 1046 32455
rect 1072 32391 1136 32455
rect 1162 32391 1226 32455
rect 1252 32391 1316 32455
rect 1342 32391 1406 32455
rect 1432 32391 1496 32455
rect 982 32311 1046 32375
rect 1072 32311 1136 32375
rect 1162 32311 1226 32375
rect 1252 32311 1316 32375
rect 1342 32311 1406 32375
rect 1432 32311 1496 32375
rect 982 32231 1046 32295
rect 1072 32231 1136 32295
rect 1162 32231 1226 32295
rect 1252 32231 1316 32295
rect 1342 32231 1406 32295
rect 1432 32231 1496 32295
rect 982 32151 1046 32215
rect 1072 32151 1136 32215
rect 1162 32151 1226 32215
rect 1252 32151 1316 32215
rect 1342 32151 1406 32215
rect 1432 32151 1496 32215
rect 982 32071 1046 32135
rect 1072 32071 1136 32135
rect 1162 32071 1226 32135
rect 1252 32071 1316 32135
rect 1342 32071 1406 32135
rect 1432 32071 1496 32135
rect 982 31991 1046 32055
rect 1072 31991 1136 32055
rect 1162 31991 1226 32055
rect 1252 31991 1316 32055
rect 1342 31991 1406 32055
rect 1432 31991 1496 32055
rect 982 31911 1046 31975
rect 1072 31911 1136 31975
rect 1162 31911 1226 31975
rect 1252 31911 1316 31975
rect 1342 31911 1406 31975
rect 1432 31911 1496 31975
rect 982 31831 1046 31895
rect 1072 31831 1136 31895
rect 1162 31831 1226 31895
rect 1252 31831 1316 31895
rect 1342 31831 1406 31895
rect 1432 31831 1496 31895
rect 982 31751 1046 31815
rect 1072 31751 1136 31815
rect 1162 31751 1226 31815
rect 1252 31751 1316 31815
rect 1342 31751 1406 31815
rect 1432 31751 1496 31815
rect 982 31671 1046 31735
rect 1072 31671 1136 31735
rect 1162 31671 1226 31735
rect 1252 31671 1316 31735
rect 1342 31671 1406 31735
rect 1432 31671 1496 31735
rect 982 31591 1046 31655
rect 1072 31591 1136 31655
rect 1162 31591 1226 31655
rect 1252 31591 1316 31655
rect 1342 31591 1406 31655
rect 1432 31591 1496 31655
rect 982 31511 1046 31575
rect 1072 31511 1136 31575
rect 1162 31511 1226 31575
rect 1252 31511 1316 31575
rect 1342 31511 1406 31575
rect 1432 31511 1496 31575
rect 982 31431 1046 31495
rect 1072 31431 1136 31495
rect 1162 31431 1226 31495
rect 1252 31431 1316 31495
rect 1342 31431 1406 31495
rect 1432 31431 1496 31495
rect 982 31351 1046 31415
rect 1072 31351 1136 31415
rect 1162 31351 1226 31415
rect 1252 31351 1316 31415
rect 1342 31351 1406 31415
rect 1432 31351 1496 31415
rect 982 31271 1046 31335
rect 1072 31271 1136 31335
rect 1162 31271 1226 31335
rect 1252 31271 1316 31335
rect 1342 31271 1406 31335
rect 1432 31271 1496 31335
rect 982 31191 1046 31255
rect 1072 31191 1136 31255
rect 1162 31191 1226 31255
rect 1252 31191 1316 31255
rect 1342 31191 1406 31255
rect 1432 31191 1496 31255
rect 982 31111 1046 31175
rect 1072 31111 1136 31175
rect 1162 31111 1226 31175
rect 1252 31111 1316 31175
rect 1342 31111 1406 31175
rect 1432 31111 1496 31175
rect 982 31031 1046 31095
rect 1072 31031 1136 31095
rect 1162 31031 1226 31095
rect 1252 31031 1316 31095
rect 1342 31031 1406 31095
rect 1432 31031 1496 31095
rect 982 30951 1046 31015
rect 1072 30951 1136 31015
rect 1162 30951 1226 31015
rect 1252 30951 1316 31015
rect 1342 30951 1406 31015
rect 1432 30951 1496 31015
rect 982 30871 1046 30935
rect 1072 30871 1136 30935
rect 1162 30871 1226 30935
rect 1252 30871 1316 30935
rect 1342 30871 1406 30935
rect 1432 30871 1496 30935
rect 982 30791 1046 30855
rect 1072 30791 1136 30855
rect 1162 30791 1226 30855
rect 1252 30791 1316 30855
rect 1342 30791 1406 30855
rect 1432 30791 1496 30855
rect 982 30711 1046 30775
rect 1072 30711 1136 30775
rect 1162 30711 1226 30775
rect 1252 30711 1316 30775
rect 1342 30711 1406 30775
rect 1432 30711 1496 30775
rect 982 30631 1046 30695
rect 1072 30631 1136 30695
rect 1162 30631 1226 30695
rect 1252 30631 1316 30695
rect 1342 30631 1406 30695
rect 1432 30631 1496 30695
rect 982 30551 1046 30615
rect 1072 30551 1136 30615
rect 1162 30551 1226 30615
rect 1252 30551 1316 30615
rect 1342 30551 1406 30615
rect 1432 30551 1496 30615
rect 982 30471 1046 30535
rect 1072 30471 1136 30535
rect 1162 30471 1226 30535
rect 1252 30471 1316 30535
rect 1342 30471 1406 30535
rect 1432 30471 1496 30535
rect 982 30391 1046 30455
rect 1072 30391 1136 30455
rect 1162 30391 1226 30455
rect 1252 30391 1316 30455
rect 1342 30391 1406 30455
rect 1432 30391 1496 30455
rect 982 30311 1046 30375
rect 1072 30311 1136 30375
rect 1162 30311 1226 30375
rect 1252 30311 1316 30375
rect 1342 30311 1406 30375
rect 1432 30311 1496 30375
rect 982 30231 1046 30295
rect 1072 30231 1136 30295
rect 1162 30231 1226 30295
rect 1252 30231 1316 30295
rect 1342 30231 1406 30295
rect 1432 30231 1496 30295
rect 982 30151 1046 30215
rect 1072 30151 1136 30215
rect 1162 30151 1226 30215
rect 1252 30151 1316 30215
rect 1342 30151 1406 30215
rect 1432 30151 1496 30215
rect 982 30071 1046 30135
rect 1072 30071 1136 30135
rect 1162 30071 1226 30135
rect 1252 30071 1316 30135
rect 1342 30071 1406 30135
rect 1432 30071 1496 30135
rect 982 29991 1046 30055
rect 1072 29991 1136 30055
rect 1162 29991 1226 30055
rect 1252 29991 1316 30055
rect 1342 29991 1406 30055
rect 1432 29991 1496 30055
rect 982 29911 1046 29975
rect 1072 29911 1136 29975
rect 1162 29911 1226 29975
rect 1252 29911 1316 29975
rect 1342 29911 1406 29975
rect 1432 29911 1496 29975
rect 982 29831 1046 29895
rect 1072 29831 1136 29895
rect 1162 29831 1226 29895
rect 1252 29831 1316 29895
rect 1342 29831 1406 29895
rect 1432 29831 1496 29895
rect 982 29751 1046 29815
rect 1072 29751 1136 29815
rect 1162 29751 1226 29815
rect 1252 29751 1316 29815
rect 1342 29751 1406 29815
rect 1432 29751 1496 29815
rect 982 29671 1046 29735
rect 1072 29671 1136 29735
rect 1162 29671 1226 29735
rect 1252 29671 1316 29735
rect 1342 29671 1406 29735
rect 1432 29671 1496 29735
rect 982 29591 1046 29655
rect 1072 29591 1136 29655
rect 1162 29591 1226 29655
rect 1252 29591 1316 29655
rect 1342 29591 1406 29655
rect 1432 29591 1496 29655
rect 982 29511 1046 29575
rect 1072 29511 1136 29575
rect 1162 29511 1226 29575
rect 1252 29511 1316 29575
rect 1342 29511 1406 29575
rect 1432 29511 1496 29575
rect 982 29431 1046 29495
rect 1072 29431 1136 29495
rect 1162 29431 1226 29495
rect 1252 29431 1316 29495
rect 1342 29431 1406 29495
rect 1432 29431 1496 29495
rect 982 29351 1046 29415
rect 1072 29351 1136 29415
rect 1162 29351 1226 29415
rect 1252 29351 1316 29415
rect 1342 29351 1406 29415
rect 1432 29351 1496 29415
rect 982 29271 1046 29335
rect 1072 29271 1136 29335
rect 1162 29271 1226 29335
rect 1252 29271 1316 29335
rect 1342 29271 1406 29335
rect 1432 29271 1496 29335
rect 982 29191 1046 29255
rect 1072 29191 1136 29255
rect 1162 29191 1226 29255
rect 1252 29191 1316 29255
rect 1342 29191 1406 29255
rect 1432 29191 1496 29255
rect 982 29111 1046 29175
rect 1072 29111 1136 29175
rect 1162 29111 1226 29175
rect 1252 29111 1316 29175
rect 1342 29111 1406 29175
rect 1432 29111 1496 29175
rect 982 29031 1046 29095
rect 1072 29031 1136 29095
rect 1162 29031 1226 29095
rect 1252 29031 1316 29095
rect 1342 29031 1406 29095
rect 1432 29031 1496 29095
rect 982 28951 1046 29015
rect 1072 28951 1136 29015
rect 1162 28951 1226 29015
rect 1252 28951 1316 29015
rect 1342 28951 1406 29015
rect 1432 28951 1496 29015
rect 982 28871 1046 28935
rect 1072 28871 1136 28935
rect 1162 28871 1226 28935
rect 1252 28871 1316 28935
rect 1342 28871 1406 28935
rect 1432 28871 1496 28935
rect 982 28791 1046 28855
rect 1072 28791 1136 28855
rect 1162 28791 1226 28855
rect 1252 28791 1316 28855
rect 1342 28791 1406 28855
rect 1432 28791 1496 28855
rect 982 28711 1046 28775
rect 1072 28711 1136 28775
rect 1162 28711 1226 28775
rect 1252 28711 1316 28775
rect 1342 28711 1406 28775
rect 1432 28711 1496 28775
rect 982 28631 1046 28695
rect 1072 28631 1136 28695
rect 1162 28631 1226 28695
rect 1252 28631 1316 28695
rect 1342 28631 1406 28695
rect 1432 28631 1496 28695
rect 982 28551 1046 28615
rect 1072 28551 1136 28615
rect 1162 28551 1226 28615
rect 1252 28551 1316 28615
rect 1342 28551 1406 28615
rect 1432 28551 1496 28615
rect 982 28471 1046 28535
rect 1072 28471 1136 28535
rect 1162 28471 1226 28535
rect 1252 28471 1316 28535
rect 1342 28471 1406 28535
rect 1432 28471 1496 28535
rect 982 28391 1046 28455
rect 1072 28391 1136 28455
rect 1162 28391 1226 28455
rect 1252 28391 1316 28455
rect 1342 28391 1406 28455
rect 1432 28391 1496 28455
rect 982 28311 1046 28375
rect 1072 28311 1136 28375
rect 1162 28311 1226 28375
rect 1252 28311 1316 28375
rect 1342 28311 1406 28375
rect 1432 28311 1496 28375
rect 982 28231 1046 28295
rect 1072 28231 1136 28295
rect 1162 28231 1226 28295
rect 1252 28231 1316 28295
rect 1342 28231 1406 28295
rect 1432 28231 1496 28295
rect 982 28151 1046 28215
rect 1072 28151 1136 28215
rect 1162 28151 1226 28215
rect 1252 28151 1316 28215
rect 1342 28151 1406 28215
rect 1432 28151 1496 28215
rect 982 28071 1046 28135
rect 1072 28071 1136 28135
rect 1162 28071 1226 28135
rect 1252 28071 1316 28135
rect 1342 28071 1406 28135
rect 1432 28071 1496 28135
rect 982 27991 1046 28055
rect 1072 27991 1136 28055
rect 1162 27991 1226 28055
rect 1252 27991 1316 28055
rect 1342 27991 1406 28055
rect 1432 27991 1496 28055
rect 982 27911 1046 27975
rect 1072 27911 1136 27975
rect 1162 27911 1226 27975
rect 1252 27911 1316 27975
rect 1342 27911 1406 27975
rect 1432 27911 1496 27975
rect 982 27831 1046 27895
rect 1072 27831 1136 27895
rect 1162 27831 1226 27895
rect 1252 27831 1316 27895
rect 1342 27831 1406 27895
rect 1432 27831 1496 27895
rect 982 27751 1046 27815
rect 1072 27751 1136 27815
rect 1162 27751 1226 27815
rect 1252 27751 1316 27815
rect 1342 27751 1406 27815
rect 1432 27751 1496 27815
rect 982 27671 1046 27735
rect 1072 27671 1136 27735
rect 1162 27671 1226 27735
rect 1252 27671 1316 27735
rect 1342 27671 1406 27735
rect 1432 27671 1496 27735
rect 982 27591 1046 27655
rect 1072 27591 1136 27655
rect 1162 27591 1226 27655
rect 1252 27591 1316 27655
rect 1342 27591 1406 27655
rect 1432 27591 1496 27655
rect 982 27511 1046 27575
rect 1072 27511 1136 27575
rect 1162 27511 1226 27575
rect 1252 27511 1316 27575
rect 1342 27511 1406 27575
rect 1432 27511 1496 27575
rect 982 27431 1046 27495
rect 1072 27431 1136 27495
rect 1162 27431 1226 27495
rect 1252 27431 1316 27495
rect 1342 27431 1406 27495
rect 1432 27431 1496 27495
rect 982 27351 1046 27415
rect 1072 27351 1136 27415
rect 1162 27351 1226 27415
rect 1252 27351 1316 27415
rect 1342 27351 1406 27415
rect 1432 27351 1496 27415
rect 982 27271 1046 27335
rect 1072 27271 1136 27335
rect 1162 27271 1226 27335
rect 1252 27271 1316 27335
rect 1342 27271 1406 27335
rect 1432 27271 1496 27335
rect 982 27191 1046 27255
rect 1072 27191 1136 27255
rect 1162 27191 1226 27255
rect 1252 27191 1316 27255
rect 1342 27191 1406 27255
rect 1432 27191 1496 27255
rect 982 27111 1046 27175
rect 1072 27111 1136 27175
rect 1162 27111 1226 27175
rect 1252 27111 1316 27175
rect 1342 27111 1406 27175
rect 1432 27111 1496 27175
rect 982 27031 1046 27095
rect 1072 27031 1136 27095
rect 1162 27031 1226 27095
rect 1252 27031 1316 27095
rect 1342 27031 1406 27095
rect 1432 27031 1496 27095
rect 982 26951 1046 27015
rect 1072 26951 1136 27015
rect 1162 26951 1226 27015
rect 1252 26951 1316 27015
rect 1342 26951 1406 27015
rect 1432 26951 1496 27015
rect 982 26871 1046 26935
rect 1072 26871 1136 26935
rect 1162 26871 1226 26935
rect 1252 26871 1316 26935
rect 1342 26871 1406 26935
rect 1432 26871 1496 26935
rect 982 26791 1046 26855
rect 1072 26791 1136 26855
rect 1162 26791 1226 26855
rect 1252 26791 1316 26855
rect 1342 26791 1406 26855
rect 1432 26791 1496 26855
rect 982 26711 1046 26775
rect 1072 26711 1136 26775
rect 1162 26711 1226 26775
rect 1252 26711 1316 26775
rect 1342 26711 1406 26775
rect 1432 26711 1496 26775
rect 982 26631 1046 26695
rect 1072 26631 1136 26695
rect 1162 26631 1226 26695
rect 1252 26631 1316 26695
rect 1342 26631 1406 26695
rect 1432 26631 1496 26695
rect 982 26551 1046 26615
rect 1072 26551 1136 26615
rect 1162 26551 1226 26615
rect 1252 26551 1316 26615
rect 1342 26551 1406 26615
rect 1432 26551 1496 26615
rect 982 26471 1046 26535
rect 1072 26471 1136 26535
rect 1162 26471 1226 26535
rect 1252 26471 1316 26535
rect 1342 26471 1406 26535
rect 1432 26471 1496 26535
rect 982 26391 1046 26455
rect 1072 26391 1136 26455
rect 1162 26391 1226 26455
rect 1252 26391 1316 26455
rect 1342 26391 1406 26455
rect 1432 26391 1496 26455
rect 982 26311 1046 26375
rect 1072 26311 1136 26375
rect 1162 26311 1226 26375
rect 1252 26311 1316 26375
rect 1342 26311 1406 26375
rect 1432 26311 1496 26375
rect 982 26231 1046 26295
rect 1072 26231 1136 26295
rect 1162 26231 1226 26295
rect 1252 26231 1316 26295
rect 1342 26231 1406 26295
rect 1432 26231 1496 26295
rect 982 26151 1046 26215
rect 1072 26151 1136 26215
rect 1162 26151 1226 26215
rect 1252 26151 1316 26215
rect 1342 26151 1406 26215
rect 1432 26151 1496 26215
rect 982 26071 1046 26135
rect 1072 26071 1136 26135
rect 1162 26071 1226 26135
rect 1252 26071 1316 26135
rect 1342 26071 1406 26135
rect 1432 26071 1496 26135
rect 982 25991 1046 26055
rect 1072 25991 1136 26055
rect 1162 25991 1226 26055
rect 1252 25991 1316 26055
rect 1342 25991 1406 26055
rect 1432 25991 1496 26055
rect 982 25911 1046 25975
rect 1072 25911 1136 25975
rect 1162 25911 1226 25975
rect 1252 25911 1316 25975
rect 1342 25911 1406 25975
rect 1432 25911 1496 25975
rect 982 25831 1046 25895
rect 1072 25831 1136 25895
rect 1162 25831 1226 25895
rect 1252 25831 1316 25895
rect 1342 25831 1406 25895
rect 1432 25831 1496 25895
rect 982 25751 1046 25815
rect 1072 25751 1136 25815
rect 1162 25751 1226 25815
rect 1252 25751 1316 25815
rect 1342 25751 1406 25815
rect 1432 25751 1496 25815
rect 982 25671 1046 25735
rect 1072 25671 1136 25735
rect 1162 25671 1226 25735
rect 1252 25671 1316 25735
rect 1342 25671 1406 25735
rect 1432 25671 1496 25735
rect 982 25591 1046 25655
rect 1072 25591 1136 25655
rect 1162 25591 1226 25655
rect 1252 25591 1316 25655
rect 1342 25591 1406 25655
rect 1432 25591 1496 25655
rect 982 25511 1046 25575
rect 1072 25511 1136 25575
rect 1162 25511 1226 25575
rect 1252 25511 1316 25575
rect 1342 25511 1406 25575
rect 1432 25511 1496 25575
rect 982 25431 1046 25495
rect 1072 25431 1136 25495
rect 1162 25431 1226 25495
rect 1252 25431 1316 25495
rect 1342 25431 1406 25495
rect 1432 25431 1496 25495
rect 982 25351 1046 25415
rect 1072 25351 1136 25415
rect 1162 25351 1226 25415
rect 1252 25351 1316 25415
rect 1342 25351 1406 25415
rect 1432 25351 1496 25415
rect 982 25271 1046 25335
rect 1072 25271 1136 25335
rect 1162 25271 1226 25335
rect 1252 25271 1316 25335
rect 1342 25271 1406 25335
rect 1432 25271 1496 25335
rect 982 25191 1046 25255
rect 1072 25191 1136 25255
rect 1162 25191 1226 25255
rect 1252 25191 1316 25255
rect 1342 25191 1406 25255
rect 1432 25191 1496 25255
rect 982 25111 1046 25175
rect 1072 25111 1136 25175
rect 1162 25111 1226 25175
rect 1252 25111 1316 25175
rect 1342 25111 1406 25175
rect 1432 25111 1496 25175
rect 982 25031 1046 25095
rect 1072 25031 1136 25095
rect 1162 25031 1226 25095
rect 1252 25031 1316 25095
rect 1342 25031 1406 25095
rect 1432 25031 1496 25095
rect 982 24951 1046 25015
rect 1072 24951 1136 25015
rect 1162 24951 1226 25015
rect 1252 24951 1316 25015
rect 1342 24951 1406 25015
rect 1432 24951 1496 25015
rect 982 24871 1046 24935
rect 1072 24871 1136 24935
rect 1162 24871 1226 24935
rect 1252 24871 1316 24935
rect 1342 24871 1406 24935
rect 1432 24871 1496 24935
rect 982 24791 1046 24855
rect 1072 24791 1136 24855
rect 1162 24791 1226 24855
rect 1252 24791 1316 24855
rect 1342 24791 1406 24855
rect 1432 24791 1496 24855
rect 982 24711 1046 24775
rect 1072 24711 1136 24775
rect 1162 24711 1226 24775
rect 1252 24711 1316 24775
rect 1342 24711 1406 24775
rect 1432 24711 1496 24775
rect 982 24631 1046 24695
rect 1072 24631 1136 24695
rect 1162 24631 1226 24695
rect 1252 24631 1316 24695
rect 1342 24631 1406 24695
rect 1432 24631 1496 24695
rect 982 24551 1046 24615
rect 1072 24551 1136 24615
rect 1162 24551 1226 24615
rect 1252 24551 1316 24615
rect 1342 24551 1406 24615
rect 1432 24551 1496 24615
rect 982 24471 1046 24535
rect 1072 24471 1136 24535
rect 1162 24471 1226 24535
rect 1252 24471 1316 24535
rect 1342 24471 1406 24535
rect 1432 24471 1496 24535
rect 982 24391 1046 24455
rect 1072 24391 1136 24455
rect 1162 24391 1226 24455
rect 1252 24391 1316 24455
rect 1342 24391 1406 24455
rect 1432 24391 1496 24455
rect 982 24311 1046 24375
rect 1072 24311 1136 24375
rect 1162 24311 1226 24375
rect 1252 24311 1316 24375
rect 1342 24311 1406 24375
rect 1432 24311 1496 24375
rect 982 24231 1046 24295
rect 1072 24231 1136 24295
rect 1162 24231 1226 24295
rect 1252 24231 1316 24295
rect 1342 24231 1406 24295
rect 1432 24231 1496 24295
rect 982 24151 1046 24215
rect 1072 24151 1136 24215
rect 1162 24151 1226 24215
rect 1252 24151 1316 24215
rect 1342 24151 1406 24215
rect 1432 24151 1496 24215
rect 982 24071 1046 24135
rect 1072 24071 1136 24135
rect 1162 24071 1226 24135
rect 1252 24071 1316 24135
rect 1342 24071 1406 24135
rect 1432 24071 1496 24135
rect 982 23991 1046 24055
rect 1072 23991 1136 24055
rect 1162 23991 1226 24055
rect 1252 23991 1316 24055
rect 1342 23991 1406 24055
rect 1432 23991 1496 24055
rect 982 23911 1046 23975
rect 1072 23911 1136 23975
rect 1162 23911 1226 23975
rect 1252 23911 1316 23975
rect 1342 23911 1406 23975
rect 1432 23911 1496 23975
rect 982 23831 1046 23895
rect 1072 23831 1136 23895
rect 1162 23831 1226 23895
rect 1252 23831 1316 23895
rect 1342 23831 1406 23895
rect 1432 23831 1496 23895
rect 982 23751 1046 23815
rect 1072 23751 1136 23815
rect 1162 23751 1226 23815
rect 1252 23751 1316 23815
rect 1342 23751 1406 23815
rect 1432 23751 1496 23815
rect 982 23671 1046 23735
rect 1072 23671 1136 23735
rect 1162 23671 1226 23735
rect 1252 23671 1316 23735
rect 1342 23671 1406 23735
rect 1432 23671 1496 23735
rect 982 23591 1046 23655
rect 1072 23591 1136 23655
rect 1162 23591 1226 23655
rect 1252 23591 1316 23655
rect 1342 23591 1406 23655
rect 1432 23591 1496 23655
rect 982 23511 1046 23575
rect 1072 23511 1136 23575
rect 1162 23511 1226 23575
rect 1252 23511 1316 23575
rect 1342 23511 1406 23575
rect 1432 23511 1496 23575
rect 982 23431 1046 23495
rect 1072 23431 1136 23495
rect 1162 23431 1226 23495
rect 1252 23431 1316 23495
rect 1342 23431 1406 23495
rect 1432 23431 1496 23495
rect 982 23351 1046 23415
rect 1072 23351 1136 23415
rect 1162 23351 1226 23415
rect 1252 23351 1316 23415
rect 1342 23351 1406 23415
rect 1432 23351 1496 23415
rect 982 23293 1046 23335
rect 1072 23293 1136 23335
rect 1162 23293 1226 23335
rect 1252 23293 1316 23335
rect 1342 23293 1406 23335
rect 1432 23293 1496 23335
rect 982 23271 1046 23293
rect 1072 23271 1136 23293
rect 1162 23271 1226 23293
rect 1252 23271 1316 23293
rect 1342 23271 1406 23293
rect 1432 23271 1496 23293
rect 982 23190 1046 23254
rect 1072 23190 1136 23254
rect 1162 23190 1226 23254
rect 1252 23190 1316 23254
rect 1342 23190 1406 23254
rect 1432 23190 1496 23254
rect 982 23109 1046 23173
rect 1072 23109 1136 23173
rect 1162 23109 1226 23173
rect 1252 23109 1316 23173
rect 1342 23109 1406 23173
rect 1432 23109 1496 23173
rect 982 23028 1046 23092
rect 1072 23028 1136 23092
rect 1162 23028 1226 23092
rect 1252 23028 1316 23092
rect 1342 23028 1406 23092
rect 1432 23028 1496 23092
rect 982 22947 1046 23011
rect 1072 22947 1136 23011
rect 1162 22947 1226 23011
rect 1252 22947 1316 23011
rect 1342 22947 1406 23011
rect 1432 22947 1496 23011
rect 982 22866 1046 22930
rect 1072 22866 1136 22930
rect 1162 22866 1226 22930
rect 1252 22866 1316 22930
rect 1342 22866 1406 22930
rect 1432 22866 1496 22930
rect 982 22785 1046 22849
rect 1072 22785 1136 22849
rect 1162 22785 1226 22849
rect 1252 22785 1316 22849
rect 1342 22785 1406 22849
rect 1432 22785 1496 22849
rect 982 22704 1046 22768
rect 1072 22704 1136 22768
rect 1162 22704 1226 22768
rect 1252 22704 1316 22768
rect 1342 22704 1406 22768
rect 1432 22704 1496 22768
rect 982 22623 1046 22687
rect 1072 22623 1136 22687
rect 1162 22623 1226 22687
rect 1252 22623 1316 22687
rect 1342 22623 1406 22687
rect 1432 22623 1496 22687
rect 982 22542 1046 22606
rect 1072 22542 1136 22606
rect 1162 22542 1226 22606
rect 1252 22542 1316 22606
rect 1342 22542 1406 22606
rect 1432 22542 1496 22606
rect 982 22461 1046 22525
rect 1072 22461 1136 22525
rect 1162 22461 1226 22525
rect 1252 22461 1316 22525
rect 1342 22461 1406 22525
rect 1432 22461 1496 22525
rect 982 22380 1046 22444
rect 1072 22380 1136 22444
rect 1162 22380 1226 22444
rect 1252 22380 1316 22444
rect 1342 22380 1406 22444
rect 1432 22380 1496 22444
rect 982 22299 1046 22363
rect 1072 22299 1136 22363
rect 1162 22299 1226 22363
rect 1252 22299 1316 22363
rect 1342 22299 1406 22363
rect 1432 22299 1496 22363
rect 982 22218 1046 22282
rect 1072 22218 1136 22282
rect 1162 22218 1226 22282
rect 1252 22218 1316 22282
rect 1342 22218 1406 22282
rect 1432 22218 1496 22282
rect 982 22137 1046 22201
rect 1072 22137 1136 22201
rect 1162 22137 1226 22201
rect 1252 22137 1316 22201
rect 1342 22137 1406 22201
rect 1432 22137 1496 22201
rect 982 22056 1046 22120
rect 1072 22056 1136 22120
rect 1162 22056 1226 22120
rect 1252 22056 1316 22120
rect 1342 22056 1406 22120
rect 1432 22056 1496 22120
rect 982 21975 1046 22039
rect 1072 21975 1136 22039
rect 1162 21975 1226 22039
rect 1252 21975 1316 22039
rect 1342 21975 1406 22039
rect 1432 21975 1496 22039
rect 982 21894 1046 21958
rect 1072 21894 1136 21958
rect 1162 21894 1226 21958
rect 1252 21894 1316 21958
rect 1342 21894 1406 21958
rect 1432 21894 1496 21958
rect 982 21813 1046 21877
rect 1072 21813 1136 21877
rect 1162 21813 1226 21877
rect 1252 21813 1316 21877
rect 1342 21813 1406 21877
rect 1432 21813 1496 21877
rect 982 21732 1046 21796
rect 1072 21732 1136 21796
rect 1162 21732 1226 21796
rect 1252 21732 1316 21796
rect 1342 21732 1406 21796
rect 1432 21732 1496 21796
rect 982 21651 1046 21715
rect 1072 21651 1136 21715
rect 1162 21651 1226 21715
rect 1252 21651 1316 21715
rect 1342 21651 1406 21715
rect 1432 21651 1496 21715
rect 982 21570 1046 21634
rect 1072 21570 1136 21634
rect 1162 21570 1226 21634
rect 1252 21570 1316 21634
rect 1342 21570 1406 21634
rect 1432 21570 1496 21634
rect 982 21489 1046 21553
rect 1072 21489 1136 21553
rect 1162 21489 1226 21553
rect 1252 21489 1316 21553
rect 1342 21489 1406 21553
rect 1432 21489 1496 21553
rect 982 21408 1046 21472
rect 1072 21408 1136 21472
rect 1162 21408 1226 21472
rect 1252 21408 1316 21472
rect 1342 21408 1406 21472
rect 1432 21408 1496 21472
rect 982 21327 1046 21391
rect 1072 21327 1136 21391
rect 1162 21327 1226 21391
rect 1252 21327 1316 21391
rect 1342 21327 1406 21391
rect 1432 21327 1496 21391
rect 982 21246 1046 21310
rect 1072 21246 1136 21310
rect 1162 21246 1226 21310
rect 1252 21246 1316 21310
rect 1342 21246 1406 21310
rect 1432 21246 1496 21310
rect 982 21165 1046 21229
rect 1072 21165 1136 21229
rect 1162 21165 1226 21229
rect 1252 21165 1316 21229
rect 1342 21165 1406 21229
rect 1432 21165 1496 21229
rect 982 21084 1046 21148
rect 1072 21084 1136 21148
rect 1162 21084 1226 21148
rect 1252 21084 1316 21148
rect 1342 21084 1406 21148
rect 1432 21084 1496 21148
rect 982 21003 1046 21067
rect 1072 21003 1136 21067
rect 1162 21003 1226 21067
rect 1252 21003 1316 21067
rect 1342 21003 1406 21067
rect 1432 21003 1496 21067
rect 982 20922 1046 20986
rect 1072 20922 1136 20986
rect 1162 20922 1226 20986
rect 1252 20922 1316 20986
rect 1342 20922 1406 20986
rect 1432 20922 1496 20986
rect 982 20841 1046 20905
rect 1072 20841 1136 20905
rect 1162 20841 1226 20905
rect 1252 20841 1316 20905
rect 1342 20841 1406 20905
rect 1432 20841 1496 20905
rect 1531 20861 1595 20925
rect 1141 20705 1205 20769
rect 1312 20747 1376 20811
rect 1401 20747 1465 20811
rect 1491 20747 1555 20811
rect 1581 20747 1645 20811
rect 1671 20747 1735 20811
rect 1312 20631 1376 20695
rect 1401 20631 1465 20695
rect 1491 20631 1555 20695
rect 1581 20631 1645 20695
rect 1671 20631 1735 20695
rect 1312 20515 1376 20579
rect 1401 20515 1465 20579
rect 1491 20515 1555 20579
rect 1581 20515 1645 20579
rect 1671 20515 1735 20579
rect 1812 20553 1876 20617
rect 1524 20391 1588 20455
rect 1632 20427 1696 20491
rect 1721 20427 1785 20491
rect 1811 20427 1875 20491
rect 1901 20427 1965 20491
rect 1991 20427 2055 20491
rect 1632 20311 1696 20375
rect 1721 20311 1785 20375
rect 1811 20311 1875 20375
rect 1901 20311 1965 20375
rect 1991 20311 2055 20375
rect 1632 20195 1696 20259
rect 1721 20195 1785 20259
rect 1811 20195 1875 20259
rect 1901 20195 1965 20259
rect 1991 20195 2055 20259
rect 2137 20228 2201 20292
rect 13169 33444 13233 33508
rect 13259 33444 13323 33508
rect 13349 33444 13413 33508
rect 13439 33444 13503 33508
rect 13528 33444 13592 33508
rect 13636 33480 13700 33544
rect 13348 33318 13412 33382
rect 13489 33356 13553 33420
rect 13579 33356 13643 33420
rect 13669 33356 13733 33420
rect 13759 33356 13823 33420
rect 13848 33356 13912 33420
rect 13489 33240 13553 33304
rect 13579 33240 13643 33304
rect 13669 33240 13733 33304
rect 13759 33240 13823 33304
rect 13848 33240 13912 33304
rect 13489 33124 13553 33188
rect 13579 33124 13643 33188
rect 13669 33124 13733 33188
rect 13759 33124 13823 33188
rect 13848 33124 13912 33188
rect 13520 33031 13584 33095
rect 13610 33031 13674 33095
rect 13700 33031 13764 33095
rect 13790 33031 13854 33095
rect 13880 33031 13944 33095
rect 13970 33031 14034 33095
rect 13520 32951 13584 33015
rect 13610 32951 13674 33015
rect 13700 32951 13764 33015
rect 13790 32951 13854 33015
rect 13880 32951 13944 33015
rect 13970 32951 14034 33015
rect 13520 32871 13584 32935
rect 13610 32871 13674 32935
rect 13700 32871 13764 32935
rect 13790 32871 13854 32935
rect 13880 32871 13944 32935
rect 13970 32871 14034 32935
rect 13520 32791 13584 32855
rect 13610 32791 13674 32855
rect 13700 32791 13764 32855
rect 13790 32791 13854 32855
rect 13880 32791 13944 32855
rect 13970 32791 14034 32855
rect 13520 32711 13584 32775
rect 13610 32711 13674 32775
rect 13700 32711 13764 32775
rect 13790 32711 13854 32775
rect 13880 32711 13944 32775
rect 13970 32711 14034 32775
rect 13520 32631 13584 32695
rect 13610 32631 13674 32695
rect 13700 32631 13764 32695
rect 13790 32631 13854 32695
rect 13880 32631 13944 32695
rect 13970 32631 14034 32695
rect 13520 32551 13584 32615
rect 13610 32551 13674 32615
rect 13700 32551 13764 32615
rect 13790 32551 13854 32615
rect 13880 32551 13944 32615
rect 13970 32551 14034 32615
rect 13520 32471 13584 32535
rect 13610 32471 13674 32535
rect 13700 32471 13764 32535
rect 13790 32471 13854 32535
rect 13880 32471 13944 32535
rect 13970 32471 14034 32535
rect 13520 32391 13584 32455
rect 13610 32391 13674 32455
rect 13700 32391 13764 32455
rect 13790 32391 13854 32455
rect 13880 32391 13944 32455
rect 13970 32391 14034 32455
rect 13520 32311 13584 32375
rect 13610 32311 13674 32375
rect 13700 32311 13764 32375
rect 13790 32311 13854 32375
rect 13880 32311 13944 32375
rect 13970 32311 14034 32375
rect 13520 32231 13584 32295
rect 13610 32231 13674 32295
rect 13700 32231 13764 32295
rect 13790 32231 13854 32295
rect 13880 32231 13944 32295
rect 13970 32231 14034 32295
rect 13520 32151 13584 32215
rect 13610 32151 13674 32215
rect 13700 32151 13764 32215
rect 13790 32151 13854 32215
rect 13880 32151 13944 32215
rect 13970 32151 14034 32215
rect 13520 32071 13584 32135
rect 13610 32071 13674 32135
rect 13700 32071 13764 32135
rect 13790 32071 13854 32135
rect 13880 32071 13944 32135
rect 13970 32071 14034 32135
rect 13520 31991 13584 32055
rect 13610 31991 13674 32055
rect 13700 31991 13764 32055
rect 13790 31991 13854 32055
rect 13880 31991 13944 32055
rect 13970 31991 14034 32055
rect 13520 31911 13584 31975
rect 13610 31911 13674 31975
rect 13700 31911 13764 31975
rect 13790 31911 13854 31975
rect 13880 31911 13944 31975
rect 13970 31911 14034 31975
rect 13520 31831 13584 31895
rect 13610 31831 13674 31895
rect 13700 31831 13764 31895
rect 13790 31831 13854 31895
rect 13880 31831 13944 31895
rect 13970 31831 14034 31895
rect 13520 31751 13584 31815
rect 13610 31751 13674 31815
rect 13700 31751 13764 31815
rect 13790 31751 13854 31815
rect 13880 31751 13944 31815
rect 13970 31751 14034 31815
rect 13520 31671 13584 31735
rect 13610 31671 13674 31735
rect 13700 31671 13764 31735
rect 13790 31671 13854 31735
rect 13880 31671 13944 31735
rect 13970 31671 14034 31735
rect 13520 31591 13584 31655
rect 13610 31591 13674 31655
rect 13700 31591 13764 31655
rect 13790 31591 13854 31655
rect 13880 31591 13944 31655
rect 13970 31591 14034 31655
rect 13520 31511 13584 31575
rect 13610 31511 13674 31575
rect 13700 31511 13764 31575
rect 13790 31511 13854 31575
rect 13880 31511 13944 31575
rect 13970 31511 14034 31575
rect 13520 31431 13584 31495
rect 13610 31431 13674 31495
rect 13700 31431 13764 31495
rect 13790 31431 13854 31495
rect 13880 31431 13944 31495
rect 13970 31431 14034 31495
rect 13520 31351 13584 31415
rect 13610 31351 13674 31415
rect 13700 31351 13764 31415
rect 13790 31351 13854 31415
rect 13880 31351 13944 31415
rect 13970 31351 14034 31415
rect 13520 31271 13584 31335
rect 13610 31271 13674 31335
rect 13700 31271 13764 31335
rect 13790 31271 13854 31335
rect 13880 31271 13944 31335
rect 13970 31271 14034 31335
rect 13520 31191 13584 31255
rect 13610 31191 13674 31255
rect 13700 31191 13764 31255
rect 13790 31191 13854 31255
rect 13880 31191 13944 31255
rect 13970 31191 14034 31255
rect 13520 31111 13584 31175
rect 13610 31111 13674 31175
rect 13700 31111 13764 31175
rect 13790 31111 13854 31175
rect 13880 31111 13944 31175
rect 13970 31111 14034 31175
rect 13520 31031 13584 31095
rect 13610 31031 13674 31095
rect 13700 31031 13764 31095
rect 13790 31031 13854 31095
rect 13880 31031 13944 31095
rect 13970 31031 14034 31095
rect 13520 30951 13584 31015
rect 13610 30951 13674 31015
rect 13700 30951 13764 31015
rect 13790 30951 13854 31015
rect 13880 30951 13944 31015
rect 13970 30951 14034 31015
rect 13520 30871 13584 30935
rect 13610 30871 13674 30935
rect 13700 30871 13764 30935
rect 13790 30871 13854 30935
rect 13880 30871 13944 30935
rect 13970 30871 14034 30935
rect 13520 30791 13584 30855
rect 13610 30791 13674 30855
rect 13700 30791 13764 30855
rect 13790 30791 13854 30855
rect 13880 30791 13944 30855
rect 13970 30791 14034 30855
rect 13520 30711 13584 30775
rect 13610 30711 13674 30775
rect 13700 30711 13764 30775
rect 13790 30711 13854 30775
rect 13880 30711 13944 30775
rect 13970 30711 14034 30775
rect 13520 30631 13584 30695
rect 13610 30631 13674 30695
rect 13700 30631 13764 30695
rect 13790 30631 13854 30695
rect 13880 30631 13944 30695
rect 13970 30631 14034 30695
rect 13520 30551 13584 30615
rect 13610 30551 13674 30615
rect 13700 30551 13764 30615
rect 13790 30551 13854 30615
rect 13880 30551 13944 30615
rect 13970 30551 14034 30615
rect 13520 30471 13584 30535
rect 13610 30471 13674 30535
rect 13700 30471 13764 30535
rect 13790 30471 13854 30535
rect 13880 30471 13944 30535
rect 13970 30471 14034 30535
rect 13520 30391 13584 30455
rect 13610 30391 13674 30455
rect 13700 30391 13764 30455
rect 13790 30391 13854 30455
rect 13880 30391 13944 30455
rect 13970 30391 14034 30455
rect 13520 30311 13584 30375
rect 13610 30311 13674 30375
rect 13700 30311 13764 30375
rect 13790 30311 13854 30375
rect 13880 30311 13944 30375
rect 13970 30311 14034 30375
rect 13520 30231 13584 30295
rect 13610 30231 13674 30295
rect 13700 30231 13764 30295
rect 13790 30231 13854 30295
rect 13880 30231 13944 30295
rect 13970 30231 14034 30295
rect 13520 30151 13584 30215
rect 13610 30151 13674 30215
rect 13700 30151 13764 30215
rect 13790 30151 13854 30215
rect 13880 30151 13944 30215
rect 13970 30151 14034 30215
rect 13520 30071 13584 30135
rect 13610 30071 13674 30135
rect 13700 30071 13764 30135
rect 13790 30071 13854 30135
rect 13880 30071 13944 30135
rect 13970 30071 14034 30135
rect 13520 29991 13584 30055
rect 13610 29991 13674 30055
rect 13700 29991 13764 30055
rect 13790 29991 13854 30055
rect 13880 29991 13944 30055
rect 13970 29991 14034 30055
rect 13520 29911 13584 29975
rect 13610 29911 13674 29975
rect 13700 29911 13764 29975
rect 13790 29911 13854 29975
rect 13880 29911 13944 29975
rect 13970 29911 14034 29975
rect 13520 29831 13584 29895
rect 13610 29831 13674 29895
rect 13700 29831 13764 29895
rect 13790 29831 13854 29895
rect 13880 29831 13944 29895
rect 13970 29831 14034 29895
rect 13520 29751 13584 29815
rect 13610 29751 13674 29815
rect 13700 29751 13764 29815
rect 13790 29751 13854 29815
rect 13880 29751 13944 29815
rect 13970 29751 14034 29815
rect 13520 29671 13584 29735
rect 13610 29671 13674 29735
rect 13700 29671 13764 29735
rect 13790 29671 13854 29735
rect 13880 29671 13944 29735
rect 13970 29671 14034 29735
rect 13520 29591 13584 29655
rect 13610 29591 13674 29655
rect 13700 29591 13764 29655
rect 13790 29591 13854 29655
rect 13880 29591 13944 29655
rect 13970 29591 14034 29655
rect 13520 29511 13584 29575
rect 13610 29511 13674 29575
rect 13700 29511 13764 29575
rect 13790 29511 13854 29575
rect 13880 29511 13944 29575
rect 13970 29511 14034 29575
rect 13520 29431 13584 29495
rect 13610 29431 13674 29495
rect 13700 29431 13764 29495
rect 13790 29431 13854 29495
rect 13880 29431 13944 29495
rect 13970 29431 14034 29495
rect 13520 29351 13584 29415
rect 13610 29351 13674 29415
rect 13700 29351 13764 29415
rect 13790 29351 13854 29415
rect 13880 29351 13944 29415
rect 13970 29351 14034 29415
rect 13520 29271 13584 29335
rect 13610 29271 13674 29335
rect 13700 29271 13764 29335
rect 13790 29271 13854 29335
rect 13880 29271 13944 29335
rect 13970 29271 14034 29335
rect 13520 29191 13584 29255
rect 13610 29191 13674 29255
rect 13700 29191 13764 29255
rect 13790 29191 13854 29255
rect 13880 29191 13944 29255
rect 13970 29191 14034 29255
rect 13520 29111 13584 29175
rect 13610 29111 13674 29175
rect 13700 29111 13764 29175
rect 13790 29111 13854 29175
rect 13880 29111 13944 29175
rect 13970 29111 14034 29175
rect 13520 29031 13584 29095
rect 13610 29031 13674 29095
rect 13700 29031 13764 29095
rect 13790 29031 13854 29095
rect 13880 29031 13944 29095
rect 13970 29031 14034 29095
rect 13520 28951 13584 29015
rect 13610 28951 13674 29015
rect 13700 28951 13764 29015
rect 13790 28951 13854 29015
rect 13880 28951 13944 29015
rect 13970 28951 14034 29015
rect 13520 28917 13584 28935
rect 13610 28917 13674 28935
rect 13700 28917 13764 28935
rect 13790 28917 13854 28935
rect 13880 28917 13944 28935
rect 13970 28917 14034 28935
rect 13520 28871 13584 28917
rect 13610 28871 13674 28917
rect 13700 28871 13764 28917
rect 13790 28871 13854 28917
rect 13880 28871 13944 28917
rect 13970 28871 14034 28917
rect 13520 28791 13584 28855
rect 13610 28791 13674 28855
rect 13700 28791 13764 28855
rect 13790 28791 13854 28855
rect 13880 28791 13944 28855
rect 13970 28791 14034 28855
rect 13520 28711 13584 28775
rect 13610 28711 13674 28775
rect 13700 28711 13764 28775
rect 13790 28711 13854 28775
rect 13880 28711 13944 28775
rect 13970 28711 14034 28775
rect 13520 28631 13584 28695
rect 13610 28631 13674 28695
rect 13700 28631 13764 28695
rect 13790 28631 13854 28695
rect 13880 28631 13944 28695
rect 13970 28631 14034 28695
rect 13520 28551 13584 28615
rect 13610 28551 13674 28615
rect 13700 28551 13764 28615
rect 13790 28551 13854 28615
rect 13880 28551 13944 28615
rect 13970 28551 14034 28615
rect 13520 28471 13584 28535
rect 13610 28471 13674 28535
rect 13700 28471 13764 28535
rect 13790 28471 13854 28535
rect 13880 28471 13944 28535
rect 13970 28471 14034 28535
rect 13520 28391 13584 28455
rect 13610 28391 13674 28455
rect 13700 28391 13764 28455
rect 13790 28391 13854 28455
rect 13880 28391 13944 28455
rect 13970 28391 14034 28455
rect 13520 28311 13584 28375
rect 13610 28311 13674 28375
rect 13700 28311 13764 28375
rect 13790 28311 13854 28375
rect 13880 28311 13944 28375
rect 13970 28311 14034 28375
rect 13520 28231 13584 28295
rect 13610 28231 13674 28295
rect 13700 28231 13764 28295
rect 13790 28231 13854 28295
rect 13880 28231 13944 28295
rect 13970 28231 14034 28295
rect 13520 28151 13584 28215
rect 13610 28151 13674 28215
rect 13700 28151 13764 28215
rect 13790 28151 13854 28215
rect 13880 28151 13944 28215
rect 13970 28151 14034 28215
rect 13520 28071 13584 28135
rect 13610 28071 13674 28135
rect 13700 28071 13764 28135
rect 13790 28071 13854 28135
rect 13880 28071 13944 28135
rect 13970 28071 14034 28135
rect 13520 27991 13584 28055
rect 13610 27991 13674 28055
rect 13700 27991 13764 28055
rect 13790 27991 13854 28055
rect 13880 27991 13944 28055
rect 13970 27991 14034 28055
rect 13520 27911 13584 27975
rect 13610 27911 13674 27975
rect 13700 27911 13764 27975
rect 13790 27911 13854 27975
rect 13880 27911 13944 27975
rect 13970 27911 14034 27975
rect 13520 27831 13584 27895
rect 13610 27831 13674 27895
rect 13700 27831 13764 27895
rect 13790 27831 13854 27895
rect 13880 27831 13944 27895
rect 13970 27831 14034 27895
rect 13520 27751 13584 27815
rect 13610 27751 13674 27815
rect 13700 27751 13764 27815
rect 13790 27751 13854 27815
rect 13880 27751 13944 27815
rect 13970 27751 14034 27815
rect 13520 27671 13584 27735
rect 13610 27671 13674 27735
rect 13700 27671 13764 27735
rect 13790 27671 13854 27735
rect 13880 27671 13944 27735
rect 13970 27671 14034 27735
rect 13520 27591 13584 27655
rect 13610 27591 13674 27655
rect 13700 27591 13764 27655
rect 13790 27591 13854 27655
rect 13880 27591 13944 27655
rect 13970 27591 14034 27655
rect 13520 27511 13584 27575
rect 13610 27511 13674 27575
rect 13700 27511 13764 27575
rect 13790 27511 13854 27575
rect 13880 27511 13944 27575
rect 13970 27511 14034 27575
rect 13520 27431 13584 27495
rect 13610 27431 13674 27495
rect 13700 27431 13764 27495
rect 13790 27431 13854 27495
rect 13880 27431 13944 27495
rect 13970 27431 14034 27495
rect 13520 27351 13584 27415
rect 13610 27351 13674 27415
rect 13700 27351 13764 27415
rect 13790 27351 13854 27415
rect 13880 27351 13944 27415
rect 13970 27351 14034 27415
rect 13520 27271 13584 27335
rect 13610 27271 13674 27335
rect 13700 27271 13764 27335
rect 13790 27271 13854 27335
rect 13880 27271 13944 27335
rect 13970 27271 14034 27335
rect 13520 27191 13584 27255
rect 13610 27191 13674 27255
rect 13700 27191 13764 27255
rect 13790 27191 13854 27255
rect 13880 27191 13944 27255
rect 13970 27191 14034 27255
rect 13520 27111 13584 27175
rect 13610 27111 13674 27175
rect 13700 27111 13764 27175
rect 13790 27111 13854 27175
rect 13880 27111 13944 27175
rect 13970 27111 14034 27175
rect 13520 27031 13584 27095
rect 13610 27031 13674 27095
rect 13700 27031 13764 27095
rect 13790 27031 13854 27095
rect 13880 27031 13944 27095
rect 13970 27031 14034 27095
rect 13520 26951 13584 27015
rect 13610 26951 13674 27015
rect 13700 26951 13764 27015
rect 13790 26951 13854 27015
rect 13880 26951 13944 27015
rect 13970 26951 14034 27015
rect 13520 26871 13584 26935
rect 13610 26871 13674 26935
rect 13700 26871 13764 26935
rect 13790 26871 13854 26935
rect 13880 26871 13944 26935
rect 13970 26871 14034 26935
rect 13520 26791 13584 26855
rect 13610 26791 13674 26855
rect 13700 26791 13764 26855
rect 13790 26791 13854 26855
rect 13880 26791 13944 26855
rect 13970 26791 14034 26855
rect 13520 26711 13584 26775
rect 13610 26711 13674 26775
rect 13700 26711 13764 26775
rect 13790 26711 13854 26775
rect 13880 26711 13944 26775
rect 13970 26711 14034 26775
rect 13520 26631 13584 26695
rect 13610 26631 13674 26695
rect 13700 26631 13764 26695
rect 13790 26631 13854 26695
rect 13880 26631 13944 26695
rect 13970 26631 14034 26695
rect 13520 26551 13584 26615
rect 13610 26551 13674 26615
rect 13700 26551 13764 26615
rect 13790 26551 13854 26615
rect 13880 26551 13944 26615
rect 13970 26551 14034 26615
rect 13520 26471 13584 26535
rect 13610 26471 13674 26535
rect 13700 26471 13764 26535
rect 13790 26471 13854 26535
rect 13880 26471 13944 26535
rect 13970 26471 14034 26535
rect 13520 26391 13584 26455
rect 13610 26391 13674 26455
rect 13700 26391 13764 26455
rect 13790 26391 13854 26455
rect 13880 26391 13944 26455
rect 13970 26391 14034 26455
rect 13520 26311 13584 26375
rect 13610 26311 13674 26375
rect 13700 26311 13764 26375
rect 13790 26311 13854 26375
rect 13880 26311 13944 26375
rect 13970 26311 14034 26375
rect 13520 26231 13584 26295
rect 13610 26231 13674 26295
rect 13700 26231 13764 26295
rect 13790 26231 13854 26295
rect 13880 26231 13944 26295
rect 13970 26231 14034 26295
rect 13520 26151 13584 26215
rect 13610 26151 13674 26215
rect 13700 26151 13764 26215
rect 13790 26151 13854 26215
rect 13880 26151 13944 26215
rect 13970 26151 14034 26215
rect 13520 26071 13584 26135
rect 13610 26071 13674 26135
rect 13700 26071 13764 26135
rect 13790 26071 13854 26135
rect 13880 26071 13944 26135
rect 13970 26071 14034 26135
rect 13520 25991 13584 26055
rect 13610 25991 13674 26055
rect 13700 25991 13764 26055
rect 13790 25991 13854 26055
rect 13880 25991 13944 26055
rect 13970 25991 14034 26055
rect 13520 25911 13584 25975
rect 13610 25911 13674 25975
rect 13700 25911 13764 25975
rect 13790 25911 13854 25975
rect 13880 25911 13944 25975
rect 13970 25911 14034 25975
rect 13520 25831 13584 25895
rect 13610 25831 13674 25895
rect 13700 25831 13764 25895
rect 13790 25831 13854 25895
rect 13880 25831 13944 25895
rect 13970 25831 14034 25895
rect 13520 25751 13584 25815
rect 13610 25751 13674 25815
rect 13700 25751 13764 25815
rect 13790 25751 13854 25815
rect 13880 25751 13944 25815
rect 13970 25751 14034 25815
rect 13520 25671 13584 25735
rect 13610 25671 13674 25735
rect 13700 25671 13764 25735
rect 13790 25671 13854 25735
rect 13880 25671 13944 25735
rect 13970 25671 14034 25735
rect 13520 25591 13584 25655
rect 13610 25591 13674 25655
rect 13700 25591 13764 25655
rect 13790 25591 13854 25655
rect 13880 25591 13944 25655
rect 13970 25591 14034 25655
rect 13520 25511 13584 25575
rect 13610 25511 13674 25575
rect 13700 25511 13764 25575
rect 13790 25511 13854 25575
rect 13880 25511 13944 25575
rect 13970 25511 14034 25575
rect 13520 25431 13584 25495
rect 13610 25431 13674 25495
rect 13700 25431 13764 25495
rect 13790 25431 13854 25495
rect 13880 25431 13944 25495
rect 13970 25431 14034 25495
rect 13520 25351 13584 25415
rect 13610 25351 13674 25415
rect 13700 25351 13764 25415
rect 13790 25351 13854 25415
rect 13880 25351 13944 25415
rect 13970 25351 14034 25415
rect 13520 25271 13584 25335
rect 13610 25271 13674 25335
rect 13700 25271 13764 25335
rect 13790 25271 13854 25335
rect 13880 25271 13944 25335
rect 13970 25271 14034 25335
rect 13520 25191 13584 25255
rect 13610 25191 13674 25255
rect 13700 25191 13764 25255
rect 13790 25191 13854 25255
rect 13880 25191 13944 25255
rect 13970 25191 14034 25255
rect 13520 25111 13584 25175
rect 13610 25111 13674 25175
rect 13700 25111 13764 25175
rect 13790 25111 13854 25175
rect 13880 25111 13944 25175
rect 13970 25111 14034 25175
rect 13520 25031 13584 25095
rect 13610 25031 13674 25095
rect 13700 25031 13764 25095
rect 13790 25031 13854 25095
rect 13880 25031 13944 25095
rect 13970 25031 14034 25095
rect 13520 24951 13584 25015
rect 13610 24951 13674 25015
rect 13700 24951 13764 25015
rect 13790 24951 13854 25015
rect 13880 24951 13944 25015
rect 13970 24951 14034 25015
rect 13520 24871 13584 24935
rect 13610 24871 13674 24935
rect 13700 24871 13764 24935
rect 13790 24871 13854 24935
rect 13880 24871 13944 24935
rect 13970 24871 14034 24935
rect 13520 24791 13584 24855
rect 13610 24791 13674 24855
rect 13700 24791 13764 24855
rect 13790 24791 13854 24855
rect 13880 24791 13944 24855
rect 13970 24791 14034 24855
rect 13520 24711 13584 24775
rect 13610 24711 13674 24775
rect 13700 24711 13764 24775
rect 13790 24711 13854 24775
rect 13880 24711 13944 24775
rect 13970 24711 14034 24775
rect 13520 24631 13584 24695
rect 13610 24631 13674 24695
rect 13700 24631 13764 24695
rect 13790 24631 13854 24695
rect 13880 24631 13944 24695
rect 13970 24631 14034 24695
rect 13520 24551 13584 24615
rect 13610 24551 13674 24615
rect 13700 24551 13764 24615
rect 13790 24551 13854 24615
rect 13880 24551 13944 24615
rect 13970 24551 14034 24615
rect 13520 24471 13584 24535
rect 13610 24471 13674 24535
rect 13700 24471 13764 24535
rect 13790 24471 13854 24535
rect 13880 24471 13944 24535
rect 13970 24471 14034 24535
rect 13520 24391 13584 24455
rect 13610 24391 13674 24455
rect 13700 24391 13764 24455
rect 13790 24391 13854 24455
rect 13880 24391 13944 24455
rect 13970 24391 14034 24455
rect 13520 24311 13584 24375
rect 13610 24311 13674 24375
rect 13700 24311 13764 24375
rect 13790 24311 13854 24375
rect 13880 24311 13944 24375
rect 13970 24311 14034 24375
rect 13520 24231 13584 24295
rect 13610 24231 13674 24295
rect 13700 24231 13764 24295
rect 13790 24231 13854 24295
rect 13880 24231 13944 24295
rect 13970 24231 14034 24295
rect 13520 24151 13584 24215
rect 13610 24151 13674 24215
rect 13700 24151 13764 24215
rect 13790 24151 13854 24215
rect 13880 24151 13944 24215
rect 13970 24151 14034 24215
rect 13520 24071 13584 24135
rect 13610 24071 13674 24135
rect 13700 24071 13764 24135
rect 13790 24071 13854 24135
rect 13880 24071 13944 24135
rect 13970 24071 14034 24135
rect 13520 23991 13584 24055
rect 13610 23991 13674 24055
rect 13700 23991 13764 24055
rect 13790 23991 13854 24055
rect 13880 23991 13944 24055
rect 13970 23991 14034 24055
rect 13520 23911 13584 23975
rect 13610 23911 13674 23975
rect 13700 23911 13764 23975
rect 13790 23911 13854 23975
rect 13880 23911 13944 23975
rect 13970 23911 14034 23975
rect 13520 23831 13584 23895
rect 13610 23831 13674 23895
rect 13700 23831 13764 23895
rect 13790 23831 13854 23895
rect 13880 23831 13944 23895
rect 13970 23831 14034 23895
rect 13520 23751 13584 23815
rect 13610 23751 13674 23815
rect 13700 23751 13764 23815
rect 13790 23751 13854 23815
rect 13880 23751 13944 23815
rect 13970 23751 14034 23815
rect 13520 23671 13584 23735
rect 13610 23671 13674 23735
rect 13700 23671 13764 23735
rect 13790 23671 13854 23735
rect 13880 23671 13944 23735
rect 13970 23671 14034 23735
rect 13520 23591 13584 23655
rect 13610 23591 13674 23655
rect 13700 23591 13764 23655
rect 13790 23591 13854 23655
rect 13880 23591 13944 23655
rect 13970 23591 14034 23655
rect 13520 23511 13584 23575
rect 13610 23511 13674 23575
rect 13700 23511 13764 23575
rect 13790 23511 13854 23575
rect 13880 23511 13944 23575
rect 13970 23511 14034 23575
rect 13520 23431 13584 23495
rect 13610 23431 13674 23495
rect 13700 23431 13764 23495
rect 13790 23431 13854 23495
rect 13880 23431 13944 23495
rect 13970 23431 14034 23495
rect 13520 23351 13584 23415
rect 13610 23351 13674 23415
rect 13700 23351 13764 23415
rect 13790 23351 13854 23415
rect 13880 23351 13944 23415
rect 13970 23351 14034 23415
rect 13520 23271 13584 23335
rect 13610 23271 13674 23335
rect 13700 23271 13764 23335
rect 13790 23271 13854 23335
rect 13880 23271 13944 23335
rect 13970 23271 14034 23335
rect 13520 23190 13584 23254
rect 13610 23190 13674 23254
rect 13700 23190 13764 23254
rect 13790 23190 13854 23254
rect 13880 23190 13944 23254
rect 13970 23190 14034 23254
rect 13520 23109 13584 23173
rect 13610 23109 13674 23173
rect 13700 23109 13764 23173
rect 13790 23109 13854 23173
rect 13880 23109 13944 23173
rect 13970 23109 14034 23173
rect 13520 23028 13584 23092
rect 13610 23028 13674 23092
rect 13700 23028 13764 23092
rect 13790 23028 13854 23092
rect 13880 23028 13944 23092
rect 13970 23028 14034 23092
rect 13520 22947 13584 23011
rect 13610 22947 13674 23011
rect 13700 22947 13764 23011
rect 13790 22947 13854 23011
rect 13880 22947 13944 23011
rect 13970 22947 14034 23011
rect 13520 22866 13584 22930
rect 13610 22866 13674 22930
rect 13700 22866 13764 22930
rect 13790 22866 13854 22930
rect 13880 22866 13944 22930
rect 13970 22866 14034 22930
rect 13520 22785 13584 22849
rect 13610 22785 13674 22849
rect 13700 22785 13764 22849
rect 13790 22785 13854 22849
rect 13880 22785 13944 22849
rect 13970 22785 14034 22849
rect 13520 22704 13584 22768
rect 13610 22704 13674 22768
rect 13700 22704 13764 22768
rect 13790 22704 13854 22768
rect 13880 22704 13944 22768
rect 13970 22704 14034 22768
rect 13520 22623 13584 22687
rect 13610 22623 13674 22687
rect 13700 22623 13764 22687
rect 13790 22623 13854 22687
rect 13880 22623 13944 22687
rect 13970 22623 14034 22687
rect 13520 22542 13584 22606
rect 13610 22542 13674 22606
rect 13700 22542 13764 22606
rect 13790 22542 13854 22606
rect 13880 22542 13944 22606
rect 13970 22542 14034 22606
rect 13520 22461 13584 22525
rect 13610 22461 13674 22525
rect 13700 22461 13764 22525
rect 13790 22461 13854 22525
rect 13880 22461 13944 22525
rect 13970 22461 14034 22525
rect 13520 22380 13584 22444
rect 13610 22380 13674 22444
rect 13700 22380 13764 22444
rect 13790 22380 13854 22444
rect 13880 22380 13944 22444
rect 13970 22380 14034 22444
rect 13520 22299 13584 22363
rect 13610 22299 13674 22363
rect 13700 22299 13764 22363
rect 13790 22299 13854 22363
rect 13880 22299 13944 22363
rect 13970 22299 14034 22363
rect 13520 22218 13584 22282
rect 13610 22218 13674 22282
rect 13700 22218 13764 22282
rect 13790 22218 13854 22282
rect 13880 22218 13944 22282
rect 13970 22218 14034 22282
rect 13520 22137 13584 22201
rect 13610 22137 13674 22201
rect 13700 22137 13764 22201
rect 13790 22137 13854 22201
rect 13880 22137 13944 22201
rect 13970 22137 14034 22201
rect 13520 22056 13584 22120
rect 13610 22056 13674 22120
rect 13700 22056 13764 22120
rect 13790 22056 13854 22120
rect 13880 22056 13944 22120
rect 13970 22056 14034 22120
rect 13520 21975 13584 22039
rect 13610 21975 13674 22039
rect 13700 21975 13764 22039
rect 13790 21975 13854 22039
rect 13880 21975 13944 22039
rect 13970 21975 14034 22039
rect 13520 21894 13584 21958
rect 13610 21894 13674 21958
rect 13700 21894 13764 21958
rect 13790 21894 13854 21958
rect 13880 21894 13944 21958
rect 13970 21894 14034 21958
rect 13520 21813 13584 21877
rect 13610 21813 13674 21877
rect 13700 21813 13764 21877
rect 13790 21813 13854 21877
rect 13880 21813 13944 21877
rect 13970 21813 14034 21877
rect 13520 21732 13584 21796
rect 13610 21732 13674 21796
rect 13700 21732 13764 21796
rect 13790 21732 13854 21796
rect 13880 21732 13944 21796
rect 13970 21732 14034 21796
rect 13520 21651 13584 21715
rect 13610 21651 13674 21715
rect 13700 21651 13764 21715
rect 13790 21651 13854 21715
rect 13880 21651 13944 21715
rect 13970 21651 14034 21715
rect 13520 21570 13584 21634
rect 13610 21570 13674 21634
rect 13700 21570 13764 21634
rect 13790 21570 13854 21634
rect 13880 21570 13944 21634
rect 13970 21570 14034 21634
rect 13520 21489 13584 21553
rect 13610 21489 13674 21553
rect 13700 21489 13764 21553
rect 13790 21489 13854 21553
rect 13880 21489 13944 21553
rect 13970 21489 14034 21553
rect 13520 21408 13584 21472
rect 13610 21408 13674 21472
rect 13700 21408 13764 21472
rect 13790 21408 13854 21472
rect 13880 21408 13944 21472
rect 13970 21408 14034 21472
rect 13520 21327 13584 21391
rect 13610 21327 13674 21391
rect 13700 21327 13764 21391
rect 13790 21327 13854 21391
rect 13880 21327 13944 21391
rect 13970 21327 14034 21391
rect 13520 21246 13584 21310
rect 13610 21246 13674 21310
rect 13700 21246 13764 21310
rect 13790 21246 13854 21310
rect 13880 21246 13944 21310
rect 13970 21246 14034 21310
rect 13520 21165 13584 21229
rect 13610 21165 13674 21229
rect 13700 21165 13764 21229
rect 13790 21165 13854 21229
rect 13880 21165 13944 21229
rect 13970 21165 14034 21229
rect 13520 21084 13584 21148
rect 13610 21084 13674 21148
rect 13700 21084 13764 21148
rect 13790 21084 13854 21148
rect 13880 21084 13944 21148
rect 13970 21084 14034 21148
rect 13520 21003 13584 21067
rect 13610 21003 13674 21067
rect 13700 21003 13764 21067
rect 13790 21003 13854 21067
rect 13880 21003 13944 21067
rect 13970 21003 14034 21067
rect 13421 20861 13485 20925
rect 13520 20922 13584 20986
rect 13610 20922 13674 20986
rect 13700 20922 13764 20986
rect 13790 20922 13854 20986
rect 13880 20922 13944 20986
rect 13970 20922 14034 20986
rect 13520 20841 13584 20905
rect 13610 20841 13674 20905
rect 13700 20841 13764 20905
rect 13790 20841 13854 20905
rect 13880 20841 13944 20905
rect 13970 20841 14034 20905
rect 13281 20747 13345 20811
rect 13371 20747 13435 20811
rect 13461 20747 13525 20811
rect 13551 20747 13615 20811
rect 13640 20747 13704 20811
rect 13749 20745 13813 20809
rect 13851 20738 13915 20802
rect 13281 20631 13345 20695
rect 13371 20631 13435 20695
rect 13461 20631 13525 20695
rect 13551 20631 13615 20695
rect 13640 20631 13704 20695
rect 13749 20634 13813 20698
rect 13140 20553 13204 20617
rect 13281 20515 13345 20579
rect 13371 20515 13435 20579
rect 13461 20515 13525 20579
rect 13551 20515 13615 20579
rect 13640 20515 13704 20579
rect 12961 20427 13025 20491
rect 13051 20427 13115 20491
rect 13141 20427 13205 20491
rect 13231 20427 13295 20491
rect 13320 20427 13384 20491
rect 13428 20391 13492 20455
rect 12961 20311 13025 20375
rect 13051 20311 13115 20375
rect 13141 20311 13205 20375
rect 13231 20311 13295 20375
rect 13320 20311 13384 20375
rect 1852 20063 1916 20127
rect 1956 20103 2020 20167
rect 2045 20103 2109 20167
rect 2135 20103 2199 20167
rect 2225 20103 2289 20167
rect 2315 20103 2379 20167
rect 12815 20228 12879 20292
rect 12961 20195 13025 20259
rect 13051 20195 13115 20259
rect 13141 20195 13205 20259
rect 13231 20195 13295 20259
rect 13320 20195 13384 20259
rect 12637 20103 12701 20167
rect 12727 20103 12791 20167
rect 12817 20103 12881 20167
rect 12907 20103 12971 20167
rect 12996 20103 13060 20167
rect 13100 20063 13164 20127
rect 1956 19987 2020 20051
rect 2045 19987 2109 20051
rect 2135 19987 2199 20051
rect 2225 19987 2289 20051
rect 2315 19987 2379 20051
rect 2456 19992 2520 20056
rect 2571 19992 2635 20056
rect 2686 19992 2750 20056
rect 2802 19992 2866 20056
rect 12150 19992 12214 20056
rect 12266 19992 12330 20056
rect 12381 19992 12445 20056
rect 12496 19992 12560 20056
rect 12637 19987 12701 20051
rect 12727 19987 12791 20051
rect 12817 19987 12881 20051
rect 12907 19987 12971 20051
rect 12996 19987 13060 20051
rect 1956 19871 2020 19935
rect 2045 19871 2109 19935
rect 2135 19871 2199 19935
rect 2225 19871 2289 19935
rect 2315 19871 2379 19935
rect 2456 19872 2520 19936
rect 2571 19872 2635 19936
rect 2686 19872 2750 19936
rect 2802 19872 2866 19936
rect 2906 19877 2970 19941
rect 12046 19877 12110 19941
rect 12150 19872 12214 19936
rect 12266 19872 12330 19936
rect 12381 19872 12445 19936
rect 12496 19872 12560 19936
rect 12637 19871 12701 19935
rect 12727 19871 12791 19935
rect 12817 19871 12881 19935
rect 12907 19871 12971 19935
rect 12996 19871 13060 19935
rect 2193 19722 2257 19786
rect 2293 19766 2357 19830
rect 2377 19766 2441 19830
rect 2461 19766 2525 19830
rect 2545 19766 2609 19830
rect 2629 19766 2693 19830
rect 2713 19766 2777 19830
rect 2797 19766 2861 19830
rect 2881 19766 2945 19830
rect 2965 19766 3029 19830
rect 3049 19766 3113 19830
rect 2293 19650 2357 19714
rect 2377 19650 2441 19714
rect 2461 19650 2525 19714
rect 2545 19650 2609 19714
rect 2629 19650 2693 19714
rect 2713 19650 2777 19714
rect 2797 19650 2861 19714
rect 2881 19650 2945 19714
rect 2965 19650 3029 19714
rect 3049 19650 3113 19714
rect 11903 19766 11967 19830
rect 11987 19766 12051 19830
rect 12071 19766 12135 19830
rect 12155 19766 12219 19830
rect 12239 19766 12303 19830
rect 12323 19766 12387 19830
rect 12407 19766 12471 19830
rect 12491 19766 12555 19830
rect 12575 19766 12639 19830
rect 12659 19766 12723 19830
rect 12759 19722 12823 19786
rect 3153 19629 3217 19693
rect 2293 19534 2357 19598
rect 2377 19534 2441 19598
rect 2461 19534 2525 19598
rect 2545 19534 2609 19598
rect 2629 19534 2693 19598
rect 2713 19534 2777 19598
rect 2797 19534 2861 19598
rect 2881 19534 2945 19598
rect 2965 19534 3029 19598
rect 3049 19534 3113 19598
rect 3153 19536 3217 19600
rect 11799 19629 11863 19693
rect 11903 19650 11967 19714
rect 11987 19650 12051 19714
rect 12071 19650 12135 19714
rect 12155 19650 12219 19714
rect 12239 19650 12303 19714
rect 12323 19650 12387 19714
rect 12407 19650 12471 19714
rect 12491 19650 12555 19714
rect 12575 19650 12639 19714
rect 12659 19650 12723 19714
rect 11799 19536 11863 19600
rect 11903 19534 11967 19598
rect 11987 19534 12051 19598
rect 12071 19534 12135 19598
rect 12155 19534 12219 19598
rect 12239 19534 12303 19598
rect 12323 19534 12387 19598
rect 12407 19534 12471 19598
rect 12491 19534 12555 19598
rect 12575 19534 12639 19598
rect 12659 19534 12723 19598
rect 4938 17311 4942 18895
rect 4942 17311 7238 18895
rect 7238 17311 7242 18895
rect 7738 17311 7742 18895
rect 7742 17311 10038 18895
rect 10038 17311 10042 18895
rect 5099 17214 7243 17218
rect 5099 17078 5103 17214
rect 5103 17078 7239 17214
rect 7239 17078 7243 17214
rect 5099 17074 7243 17078
rect 7735 17214 9879 17218
rect 7735 17078 7739 17214
rect 7739 17078 9875 17214
rect 9875 17078 9879 17214
rect 7735 17074 9879 17078
rect 2423 5241 3607 6025
rect 887 4027 2071 4811
rect 11297 5240 12481 6024
rect 12887 4027 14071 4811
<< metal4 >>
rect 4949 39217 7225 39241
rect 767 36409 1727 37008
rect 4949 35313 4975 39217
rect 7199 35313 7225 39217
rect 4949 35290 7225 35313
rect 7749 39217 10025 39241
rect 7749 35313 7775 39217
rect 9999 35313 10025 39217
rect 13204 36409 14164 37008
rect 7749 35290 10025 35313
rect 2275 34604 2676 34607
rect 2275 34540 2276 34604
rect 2340 34540 2359 34604
rect 2423 34540 2443 34604
rect 2507 34540 2527 34604
rect 2591 34540 2611 34604
rect 2675 34540 2676 34604
rect 2275 34510 2676 34540
rect 2131 34427 2213 34460
rect 2131 34363 2148 34427
rect 2212 34363 2213 34427
rect 2131 34330 2213 34363
rect 2275 34446 2276 34510
rect 2340 34446 2359 34510
rect 2423 34446 2443 34510
rect 2507 34446 2527 34510
rect 2591 34446 2611 34510
rect 2675 34446 2676 34510
rect 2275 34416 2676 34446
rect 2275 34352 2276 34416
rect 2340 34352 2359 34416
rect 2423 34352 2443 34416
rect 2507 34352 2527 34416
rect 2591 34352 2611 34416
rect 2675 34352 2676 34416
rect 2275 34322 2676 34352
rect 2002 34302 2230 34303
rect 2002 34238 2004 34302
rect 2068 34238 2084 34302
rect 2148 34238 2164 34302
rect 2228 34238 2230 34302
rect 2002 34206 2230 34238
rect 1873 34169 1955 34202
rect 1873 34105 1890 34169
rect 1954 34105 1955 34169
rect 2002 34142 2004 34206
rect 2068 34142 2084 34206
rect 2148 34142 2164 34206
rect 2228 34142 2230 34206
rect 2002 34141 2230 34142
rect 2275 34258 2276 34322
rect 2340 34258 2359 34322
rect 2423 34258 2443 34322
rect 2507 34258 2527 34322
rect 2591 34258 2611 34322
rect 2675 34258 2676 34322
rect 2275 34228 2676 34258
rect 2275 34164 2276 34228
rect 2340 34164 2359 34228
rect 2423 34164 2443 34228
rect 2507 34164 2527 34228
rect 2591 34164 2611 34228
rect 2675 34164 2676 34228
rect 1873 34072 1955 34105
rect 2275 34134 2676 34164
rect 2275 34070 2276 34134
rect 2340 34070 2359 34134
rect 2423 34070 2443 34134
rect 2507 34070 2527 34134
rect 2591 34070 2611 34134
rect 2675 34070 2676 34134
rect 2275 34067 2676 34070
rect 12340 34604 12742 34607
rect 12340 34540 12341 34604
rect 12405 34540 12425 34604
rect 12489 34540 12509 34604
rect 12573 34540 12593 34604
rect 12657 34540 12677 34604
rect 12741 34540 12742 34604
rect 12340 34510 12742 34540
rect 12340 34446 12341 34510
rect 12405 34446 12425 34510
rect 12489 34446 12509 34510
rect 12573 34446 12593 34510
rect 12657 34446 12677 34510
rect 12741 34446 12742 34510
rect 12340 34416 12742 34446
rect 12340 34352 12341 34416
rect 12405 34352 12425 34416
rect 12489 34352 12509 34416
rect 12573 34352 12593 34416
rect 12657 34352 12677 34416
rect 12741 34352 12742 34416
rect 12340 34322 12742 34352
rect 12803 34427 12885 34460
rect 12803 34363 12804 34427
rect 12868 34363 12885 34427
rect 12803 34330 12885 34363
rect 12340 34258 12341 34322
rect 12405 34258 12425 34322
rect 12489 34258 12509 34322
rect 12573 34258 12593 34322
rect 12657 34258 12677 34322
rect 12741 34258 12742 34322
rect 12340 34228 12742 34258
rect 12340 34164 12341 34228
rect 12405 34164 12425 34228
rect 12489 34164 12509 34228
rect 12573 34164 12593 34228
rect 12657 34164 12677 34228
rect 12741 34164 12742 34228
rect 12340 34134 12742 34164
rect 12786 34302 13014 34303
rect 12786 34238 12788 34302
rect 12852 34238 12868 34302
rect 12932 34238 12948 34302
rect 13012 34238 13014 34302
rect 12786 34206 13014 34238
rect 12786 34142 12788 34206
rect 12852 34142 12868 34206
rect 12932 34142 12948 34206
rect 13012 34142 13014 34206
rect 12786 34141 13014 34142
rect 13061 34169 13143 34202
rect 12340 34070 12341 34134
rect 12405 34070 12425 34134
rect 12489 34070 12509 34134
rect 12573 34070 12593 34134
rect 12657 34070 12677 34134
rect 12741 34070 12742 34134
rect 13061 34105 13062 34169
rect 13126 34105 13143 34169
rect 13061 34072 13143 34105
rect 12340 34067 12742 34070
rect 1747 34064 2172 34066
rect 1747 34000 1748 34064
rect 1812 34000 1837 34064
rect 1901 34000 1927 34064
rect 1991 34000 2017 34064
rect 2081 34000 2107 34064
rect 2171 34000 2172 34064
rect 12844 34064 13269 34066
rect 1747 33948 2172 34000
rect 1584 33872 1709 33905
rect 1584 33808 1644 33872
rect 1708 33808 1709 33872
rect 1584 33775 1709 33808
rect 1747 33884 1748 33948
rect 1812 33884 1837 33948
rect 1901 33884 1927 33948
rect 1991 33884 2017 33948
rect 2081 33884 2107 33948
rect 2171 33884 2172 33948
rect 2187 33995 2312 34028
rect 2187 33931 2247 33995
rect 2311 33931 2312 33995
rect 2187 33898 2312 33931
rect 12704 33995 12829 34028
rect 12704 33931 12705 33995
rect 12769 33931 12829 33995
rect 12704 33898 12829 33931
rect 12844 34000 12845 34064
rect 12909 34000 12935 34064
rect 12999 34000 13025 34064
rect 13089 34000 13115 34064
rect 13179 34000 13204 34064
rect 13268 34000 13269 34064
rect 12844 33948 13269 34000
rect 1747 33832 2172 33884
rect 1747 33768 1748 33832
rect 1812 33768 1837 33832
rect 1901 33768 1927 33832
rect 1991 33768 2017 33832
rect 2081 33768 2107 33832
rect 2171 33768 2172 33832
rect 1747 33766 2172 33768
rect 12844 33884 12845 33948
rect 12909 33884 12935 33948
rect 12999 33884 13025 33948
rect 13089 33884 13115 33948
rect 13179 33884 13204 33948
rect 13268 33884 13269 33948
rect 12844 33832 13269 33884
rect 12844 33768 12845 33832
rect 12909 33768 12935 33832
rect 12999 33768 13025 33832
rect 13089 33768 13115 33832
rect 13179 33768 13204 33832
rect 13268 33768 13269 33832
rect 13307 33872 13432 33905
rect 13307 33808 13308 33872
rect 13372 33808 13432 33872
rect 13307 33775 13432 33808
rect 12844 33766 13269 33768
rect 1423 33740 1848 33742
rect 13168 33740 13593 33742
rect 1423 33676 1424 33740
rect 1488 33676 1513 33740
rect 1577 33676 1603 33740
rect 1667 33676 1693 33740
rect 1757 33676 1783 33740
rect 1847 33676 1848 33740
rect 1423 33624 1848 33676
rect 1256 33544 1381 33577
rect 1256 33480 1316 33544
rect 1380 33480 1381 33544
rect 1256 33447 1381 33480
rect 1423 33560 1424 33624
rect 1488 33560 1513 33624
rect 1577 33560 1603 33624
rect 1667 33560 1693 33624
rect 1757 33560 1783 33624
rect 1847 33560 1848 33624
rect 1869 33707 1994 33740
rect 1869 33643 1929 33707
rect 1993 33643 1994 33707
rect 1869 33610 1994 33643
rect 13022 33707 13147 33740
rect 13022 33643 13023 33707
rect 13087 33643 13147 33707
rect 13022 33610 13147 33643
rect 13168 33676 13169 33740
rect 13233 33676 13259 33740
rect 13323 33676 13349 33740
rect 13413 33676 13439 33740
rect 13503 33676 13528 33740
rect 13592 33676 13593 33740
rect 13168 33624 13593 33676
rect 1423 33508 1848 33560
rect 1423 33444 1424 33508
rect 1488 33444 1513 33508
rect 1577 33444 1603 33508
rect 1667 33444 1693 33508
rect 1757 33444 1783 33508
rect 1847 33444 1848 33508
rect 1423 33442 1848 33444
rect 13168 33560 13169 33624
rect 13233 33560 13259 33624
rect 13323 33560 13349 33624
rect 13413 33560 13439 33624
rect 13503 33560 13528 33624
rect 13592 33560 13593 33624
rect 13168 33508 13593 33560
rect 13168 33444 13169 33508
rect 13233 33444 13259 33508
rect 13323 33444 13349 33508
rect 13413 33444 13439 33508
rect 13503 33444 13528 33508
rect 13592 33444 13593 33508
rect 13635 33544 13760 33577
rect 13635 33480 13636 33544
rect 13700 33480 13760 33544
rect 13635 33447 13760 33480
rect 13168 33442 13593 33444
rect 1103 33420 1528 33422
rect 1103 33356 1104 33420
rect 1168 33356 1193 33420
rect 1257 33356 1283 33420
rect 1347 33356 1373 33420
rect 1437 33356 1463 33420
rect 1527 33356 1528 33420
rect 13488 33420 13913 33422
rect 1103 33304 1528 33356
rect 1103 33240 1104 33304
rect 1168 33240 1193 33304
rect 1257 33240 1283 33304
rect 1347 33240 1373 33304
rect 1437 33240 1463 33304
rect 1527 33240 1528 33304
rect 1544 33382 1669 33415
rect 1544 33318 1604 33382
rect 1668 33318 1669 33382
rect 1544 33285 1669 33318
rect 13347 33382 13472 33415
rect 13347 33318 13348 33382
rect 13412 33318 13472 33382
rect 13347 33285 13472 33318
rect 13488 33356 13489 33420
rect 13553 33356 13579 33420
rect 13643 33356 13669 33420
rect 13733 33356 13759 33420
rect 13823 33356 13848 33420
rect 13912 33356 13913 33420
rect 13488 33304 13913 33356
rect 1103 33188 1528 33240
rect 1103 33124 1104 33188
rect 1168 33124 1193 33188
rect 1257 33124 1283 33188
rect 1347 33124 1373 33188
rect 1437 33124 1463 33188
rect 1527 33124 1528 33188
rect 1103 33122 1528 33124
rect 13488 33240 13489 33304
rect 13553 33240 13579 33304
rect 13643 33240 13669 33304
rect 13733 33240 13759 33304
rect 13823 33240 13848 33304
rect 13912 33240 13913 33304
rect 13488 33188 13913 33240
rect 13488 33124 13489 33188
rect 13553 33124 13579 33188
rect 13643 33124 13669 33188
rect 13733 33124 13759 33188
rect 13823 33124 13848 33188
rect 13912 33124 13913 33188
rect 13488 33122 13913 33124
rect 977 33095 1501 33096
rect 977 33031 982 33095
rect 1046 33031 1072 33095
rect 1136 33031 1162 33095
rect 1226 33031 1252 33095
rect 1316 33031 1342 33095
rect 1406 33031 1432 33095
rect 1496 33031 1501 33095
rect 977 33015 1501 33031
rect 977 32951 982 33015
rect 1046 32951 1072 33015
rect 1136 32951 1162 33015
rect 1226 32951 1252 33015
rect 1316 32951 1342 33015
rect 1406 32951 1432 33015
rect 1496 32951 1501 33015
rect 977 32935 1501 32951
rect 977 32871 982 32935
rect 1046 32871 1072 32935
rect 1136 32871 1162 32935
rect 1226 32871 1252 32935
rect 1316 32871 1342 32935
rect 1406 32871 1432 32935
rect 1496 32871 1501 32935
rect 977 32855 1501 32871
rect 977 32791 982 32855
rect 1046 32791 1072 32855
rect 1136 32791 1162 32855
rect 1226 32791 1252 32855
rect 1316 32791 1342 32855
rect 1406 32791 1432 32855
rect 1496 32791 1501 32855
rect 977 32775 1501 32791
rect 977 32711 982 32775
rect 1046 32711 1072 32775
rect 1136 32711 1162 32775
rect 1226 32711 1252 32775
rect 1316 32711 1342 32775
rect 1406 32711 1432 32775
rect 1496 32711 1501 32775
rect 977 32695 1501 32711
rect 977 32631 982 32695
rect 1046 32631 1072 32695
rect 1136 32631 1162 32695
rect 1226 32631 1252 32695
rect 1316 32631 1342 32695
rect 1406 32631 1432 32695
rect 1496 32631 1501 32695
rect 977 32615 1501 32631
rect 977 32551 982 32615
rect 1046 32551 1072 32615
rect 1136 32551 1162 32615
rect 1226 32551 1252 32615
rect 1316 32551 1342 32615
rect 1406 32551 1432 32615
rect 1496 32551 1501 32615
rect 977 32535 1501 32551
rect 977 32471 982 32535
rect 1046 32471 1072 32535
rect 1136 32471 1162 32535
rect 1226 32471 1252 32535
rect 1316 32471 1342 32535
rect 1406 32471 1432 32535
rect 1496 32471 1501 32535
rect 977 32455 1501 32471
rect 977 32391 982 32455
rect 1046 32391 1072 32455
rect 1136 32391 1162 32455
rect 1226 32391 1252 32455
rect 1316 32391 1342 32455
rect 1406 32391 1432 32455
rect 1496 32391 1501 32455
rect 977 32375 1501 32391
rect 977 32311 982 32375
rect 1046 32311 1072 32375
rect 1136 32311 1162 32375
rect 1226 32311 1252 32375
rect 1316 32311 1342 32375
rect 1406 32311 1432 32375
rect 1496 32311 1501 32375
rect 977 32295 1501 32311
rect 977 32231 982 32295
rect 1046 32231 1072 32295
rect 1136 32231 1162 32295
rect 1226 32231 1252 32295
rect 1316 32231 1342 32295
rect 1406 32231 1432 32295
rect 1496 32231 1501 32295
rect 977 32215 1501 32231
rect 977 32151 982 32215
rect 1046 32151 1072 32215
rect 1136 32151 1162 32215
rect 1226 32151 1252 32215
rect 1316 32151 1342 32215
rect 1406 32151 1432 32215
rect 1496 32151 1501 32215
rect 977 32135 1501 32151
rect 977 32071 982 32135
rect 1046 32071 1072 32135
rect 1136 32071 1162 32135
rect 1226 32071 1252 32135
rect 1316 32071 1342 32135
rect 1406 32071 1432 32135
rect 1496 32071 1501 32135
rect 977 32055 1501 32071
rect 977 31991 982 32055
rect 1046 31991 1072 32055
rect 1136 31991 1162 32055
rect 1226 31991 1252 32055
rect 1316 31991 1342 32055
rect 1406 31991 1432 32055
rect 1496 31991 1501 32055
rect 977 31975 1501 31991
rect 977 31911 982 31975
rect 1046 31911 1072 31975
rect 1136 31911 1162 31975
rect 1226 31911 1252 31975
rect 1316 31911 1342 31975
rect 1406 31911 1432 31975
rect 1496 31911 1501 31975
rect 977 31895 1501 31911
rect 977 31831 982 31895
rect 1046 31831 1072 31895
rect 1136 31831 1162 31895
rect 1226 31831 1252 31895
rect 1316 31831 1342 31895
rect 1406 31831 1432 31895
rect 1496 31831 1501 31895
rect 977 31815 1501 31831
rect 977 31751 982 31815
rect 1046 31751 1072 31815
rect 1136 31751 1162 31815
rect 1226 31751 1252 31815
rect 1316 31751 1342 31815
rect 1406 31751 1432 31815
rect 1496 31751 1501 31815
rect 977 31735 1501 31751
rect 977 31671 982 31735
rect 1046 31671 1072 31735
rect 1136 31671 1162 31735
rect 1226 31671 1252 31735
rect 1316 31671 1342 31735
rect 1406 31671 1432 31735
rect 1496 31671 1501 31735
rect 977 31655 1501 31671
rect 977 31591 982 31655
rect 1046 31591 1072 31655
rect 1136 31591 1162 31655
rect 1226 31591 1252 31655
rect 1316 31591 1342 31655
rect 1406 31591 1432 31655
rect 1496 31591 1501 31655
rect 977 31575 1501 31591
rect 977 31511 982 31575
rect 1046 31511 1072 31575
rect 1136 31511 1162 31575
rect 1226 31511 1252 31575
rect 1316 31511 1342 31575
rect 1406 31511 1432 31575
rect 1496 31511 1501 31575
rect 977 31495 1501 31511
rect 977 31431 982 31495
rect 1046 31431 1072 31495
rect 1136 31431 1162 31495
rect 1226 31431 1252 31495
rect 1316 31431 1342 31495
rect 1406 31431 1432 31495
rect 1496 31431 1501 31495
rect 977 31415 1501 31431
rect 977 31351 982 31415
rect 1046 31351 1072 31415
rect 1136 31351 1162 31415
rect 1226 31351 1252 31415
rect 1316 31351 1342 31415
rect 1406 31351 1432 31415
rect 1496 31351 1501 31415
rect 977 31335 1501 31351
rect 977 31271 982 31335
rect 1046 31271 1072 31335
rect 1136 31271 1162 31335
rect 1226 31271 1252 31335
rect 1316 31271 1342 31335
rect 1406 31271 1432 31335
rect 1496 31271 1501 31335
rect 977 31255 1501 31271
rect 977 31191 982 31255
rect 1046 31191 1072 31255
rect 1136 31191 1162 31255
rect 1226 31191 1252 31255
rect 1316 31191 1342 31255
rect 1406 31191 1432 31255
rect 1496 31191 1501 31255
rect 977 31175 1501 31191
rect 977 31111 982 31175
rect 1046 31111 1072 31175
rect 1136 31111 1162 31175
rect 1226 31111 1252 31175
rect 1316 31111 1342 31175
rect 1406 31111 1432 31175
rect 1496 31111 1501 31175
rect 977 31095 1501 31111
rect 977 31031 982 31095
rect 1046 31031 1072 31095
rect 1136 31031 1162 31095
rect 1226 31031 1252 31095
rect 1316 31031 1342 31095
rect 1406 31031 1432 31095
rect 1496 31031 1501 31095
rect 977 31015 1501 31031
rect 977 30951 982 31015
rect 1046 30951 1072 31015
rect 1136 30951 1162 31015
rect 1226 30951 1252 31015
rect 1316 30951 1342 31015
rect 1406 30951 1432 31015
rect 1496 30951 1501 31015
rect 977 30935 1501 30951
rect 977 30871 982 30935
rect 1046 30871 1072 30935
rect 1136 30871 1162 30935
rect 1226 30871 1252 30935
rect 1316 30871 1342 30935
rect 1406 30871 1432 30935
rect 1496 30871 1501 30935
rect 977 30855 1501 30871
rect 977 30791 982 30855
rect 1046 30791 1072 30855
rect 1136 30791 1162 30855
rect 1226 30791 1252 30855
rect 1316 30791 1342 30855
rect 1406 30791 1432 30855
rect 1496 30791 1501 30855
rect 977 30775 1501 30791
rect 977 30711 982 30775
rect 1046 30711 1072 30775
rect 1136 30711 1162 30775
rect 1226 30711 1252 30775
rect 1316 30711 1342 30775
rect 1406 30711 1432 30775
rect 1496 30711 1501 30775
rect 977 30695 1501 30711
rect 977 30631 982 30695
rect 1046 30631 1072 30695
rect 1136 30631 1162 30695
rect 1226 30631 1252 30695
rect 1316 30631 1342 30695
rect 1406 30631 1432 30695
rect 1496 30631 1501 30695
rect 977 30615 1501 30631
rect 977 30551 982 30615
rect 1046 30551 1072 30615
rect 1136 30551 1162 30615
rect 1226 30551 1252 30615
rect 1316 30551 1342 30615
rect 1406 30551 1432 30615
rect 1496 30551 1501 30615
rect 977 30535 1501 30551
rect 977 30471 982 30535
rect 1046 30471 1072 30535
rect 1136 30471 1162 30535
rect 1226 30471 1252 30535
rect 1316 30471 1342 30535
rect 1406 30471 1432 30535
rect 1496 30471 1501 30535
rect 977 30455 1501 30471
rect 977 30391 982 30455
rect 1046 30391 1072 30455
rect 1136 30391 1162 30455
rect 1226 30391 1252 30455
rect 1316 30391 1342 30455
rect 1406 30391 1432 30455
rect 1496 30391 1501 30455
rect 977 30375 1501 30391
rect 977 30311 982 30375
rect 1046 30311 1072 30375
rect 1136 30311 1162 30375
rect 1226 30311 1252 30375
rect 1316 30311 1342 30375
rect 1406 30311 1432 30375
rect 1496 30311 1501 30375
rect 977 30295 1501 30311
rect 977 30231 982 30295
rect 1046 30231 1072 30295
rect 1136 30231 1162 30295
rect 1226 30231 1252 30295
rect 1316 30231 1342 30295
rect 1406 30231 1432 30295
rect 1496 30231 1501 30295
rect 977 30215 1501 30231
rect 977 30151 982 30215
rect 1046 30151 1072 30215
rect 1136 30151 1162 30215
rect 1226 30151 1252 30215
rect 1316 30151 1342 30215
rect 1406 30151 1432 30215
rect 1496 30151 1501 30215
rect 977 30135 1501 30151
rect 977 30071 982 30135
rect 1046 30071 1072 30135
rect 1136 30071 1162 30135
rect 1226 30071 1252 30135
rect 1316 30071 1342 30135
rect 1406 30071 1432 30135
rect 1496 30071 1501 30135
rect 977 30055 1501 30071
rect 977 29991 982 30055
rect 1046 29991 1072 30055
rect 1136 29991 1162 30055
rect 1226 29991 1252 30055
rect 1316 29991 1342 30055
rect 1406 29991 1432 30055
rect 1496 29991 1501 30055
rect 977 29975 1501 29991
rect 977 29911 982 29975
rect 1046 29911 1072 29975
rect 1136 29911 1162 29975
rect 1226 29911 1252 29975
rect 1316 29911 1342 29975
rect 1406 29911 1432 29975
rect 1496 29911 1501 29975
rect 977 29895 1501 29911
rect 977 29831 982 29895
rect 1046 29831 1072 29895
rect 1136 29831 1162 29895
rect 1226 29831 1252 29895
rect 1316 29831 1342 29895
rect 1406 29831 1432 29895
rect 1496 29831 1501 29895
rect 977 29815 1501 29831
rect 977 29751 982 29815
rect 1046 29751 1072 29815
rect 1136 29751 1162 29815
rect 1226 29751 1252 29815
rect 1316 29751 1342 29815
rect 1406 29751 1432 29815
rect 1496 29751 1501 29815
rect 977 29735 1501 29751
rect 977 29671 982 29735
rect 1046 29671 1072 29735
rect 1136 29671 1162 29735
rect 1226 29671 1252 29735
rect 1316 29671 1342 29735
rect 1406 29671 1432 29735
rect 1496 29671 1501 29735
rect 977 29655 1501 29671
rect 977 29591 982 29655
rect 1046 29591 1072 29655
rect 1136 29591 1162 29655
rect 1226 29591 1252 29655
rect 1316 29591 1342 29655
rect 1406 29591 1432 29655
rect 1496 29591 1501 29655
rect 977 29575 1501 29591
rect 977 29511 982 29575
rect 1046 29511 1072 29575
rect 1136 29511 1162 29575
rect 1226 29511 1252 29575
rect 1316 29511 1342 29575
rect 1406 29511 1432 29575
rect 1496 29511 1501 29575
rect 977 29495 1501 29511
rect 977 29431 982 29495
rect 1046 29431 1072 29495
rect 1136 29431 1162 29495
rect 1226 29431 1252 29495
rect 1316 29431 1342 29495
rect 1406 29431 1432 29495
rect 1496 29431 1501 29495
rect 977 29415 1501 29431
rect 977 29351 982 29415
rect 1046 29351 1072 29415
rect 1136 29351 1162 29415
rect 1226 29351 1252 29415
rect 1316 29351 1342 29415
rect 1406 29351 1432 29415
rect 1496 29351 1501 29415
rect 977 29335 1501 29351
rect 977 29271 982 29335
rect 1046 29271 1072 29335
rect 1136 29271 1162 29335
rect 1226 29271 1252 29335
rect 1316 29271 1342 29335
rect 1406 29271 1432 29335
rect 1496 29271 1501 29335
rect 977 29255 1501 29271
rect 977 29191 982 29255
rect 1046 29191 1072 29255
rect 1136 29191 1162 29255
rect 1226 29191 1252 29255
rect 1316 29191 1342 29255
rect 1406 29191 1432 29255
rect 1496 29191 1501 29255
rect 977 29175 1501 29191
rect 977 29111 982 29175
rect 1046 29111 1072 29175
rect 1136 29111 1162 29175
rect 1226 29111 1252 29175
rect 1316 29111 1342 29175
rect 1406 29111 1432 29175
rect 1496 29111 1501 29175
rect 977 29095 1501 29111
rect 977 29031 982 29095
rect 1046 29031 1072 29095
rect 1136 29031 1162 29095
rect 1226 29031 1252 29095
rect 1316 29031 1342 29095
rect 1406 29031 1432 29095
rect 1496 29031 1501 29095
rect 977 29015 1501 29031
rect 977 28951 982 29015
rect 1046 28951 1072 29015
rect 1136 28951 1162 29015
rect 1226 28951 1252 29015
rect 1316 28951 1342 29015
rect 1406 28951 1432 29015
rect 1496 28951 1501 29015
rect 977 28935 1501 28951
rect 977 28871 982 28935
rect 1046 28871 1072 28935
rect 1136 28871 1162 28935
rect 1226 28871 1252 28935
rect 1316 28871 1342 28935
rect 1406 28871 1432 28935
rect 1496 28871 1501 28935
rect 977 28855 1501 28871
rect 977 28791 982 28855
rect 1046 28791 1072 28855
rect 1136 28791 1162 28855
rect 1226 28791 1252 28855
rect 1316 28791 1342 28855
rect 1406 28791 1432 28855
rect 1496 28791 1501 28855
rect 977 28775 1501 28791
rect 977 28711 982 28775
rect 1046 28711 1072 28775
rect 1136 28711 1162 28775
rect 1226 28711 1252 28775
rect 1316 28711 1342 28775
rect 1406 28711 1432 28775
rect 1496 28711 1501 28775
rect 977 28695 1501 28711
rect 977 28631 982 28695
rect 1046 28631 1072 28695
rect 1136 28631 1162 28695
rect 1226 28631 1252 28695
rect 1316 28631 1342 28695
rect 1406 28631 1432 28695
rect 1496 28631 1501 28695
rect 977 28615 1501 28631
rect 977 28551 982 28615
rect 1046 28551 1072 28615
rect 1136 28551 1162 28615
rect 1226 28551 1252 28615
rect 1316 28551 1342 28615
rect 1406 28551 1432 28615
rect 1496 28551 1501 28615
rect 977 28535 1501 28551
rect 977 28471 982 28535
rect 1046 28471 1072 28535
rect 1136 28471 1162 28535
rect 1226 28471 1252 28535
rect 1316 28471 1342 28535
rect 1406 28471 1432 28535
rect 1496 28471 1501 28535
rect 977 28455 1501 28471
rect 977 28391 982 28455
rect 1046 28391 1072 28455
rect 1136 28391 1162 28455
rect 1226 28391 1252 28455
rect 1316 28391 1342 28455
rect 1406 28391 1432 28455
rect 1496 28391 1501 28455
rect 977 28375 1501 28391
rect 977 28311 982 28375
rect 1046 28311 1072 28375
rect 1136 28311 1162 28375
rect 1226 28311 1252 28375
rect 1316 28311 1342 28375
rect 1406 28311 1432 28375
rect 1496 28311 1501 28375
rect 977 28295 1501 28311
rect 977 28231 982 28295
rect 1046 28231 1072 28295
rect 1136 28231 1162 28295
rect 1226 28231 1252 28295
rect 1316 28231 1342 28295
rect 1406 28231 1432 28295
rect 1496 28231 1501 28295
rect 977 28215 1501 28231
rect 977 28151 982 28215
rect 1046 28151 1072 28215
rect 1136 28151 1162 28215
rect 1226 28151 1252 28215
rect 1316 28151 1342 28215
rect 1406 28151 1432 28215
rect 1496 28151 1501 28215
rect 977 28135 1501 28151
rect 977 28071 982 28135
rect 1046 28071 1072 28135
rect 1136 28071 1162 28135
rect 1226 28071 1252 28135
rect 1316 28071 1342 28135
rect 1406 28071 1432 28135
rect 1496 28071 1501 28135
rect 977 28055 1501 28071
rect 977 27991 982 28055
rect 1046 27991 1072 28055
rect 1136 27991 1162 28055
rect 1226 27991 1252 28055
rect 1316 27991 1342 28055
rect 1406 27991 1432 28055
rect 1496 27991 1501 28055
rect 977 27975 1501 27991
rect 977 27911 982 27975
rect 1046 27911 1072 27975
rect 1136 27911 1162 27975
rect 1226 27911 1252 27975
rect 1316 27911 1342 27975
rect 1406 27911 1432 27975
rect 1496 27911 1501 27975
rect 977 27895 1501 27911
rect 977 27831 982 27895
rect 1046 27831 1072 27895
rect 1136 27831 1162 27895
rect 1226 27831 1252 27895
rect 1316 27831 1342 27895
rect 1406 27831 1432 27895
rect 1496 27831 1501 27895
rect 977 27815 1501 27831
rect 977 27751 982 27815
rect 1046 27751 1072 27815
rect 1136 27751 1162 27815
rect 1226 27751 1252 27815
rect 1316 27751 1342 27815
rect 1406 27751 1432 27815
rect 1496 27751 1501 27815
rect 977 27735 1501 27751
rect 977 27671 982 27735
rect 1046 27671 1072 27735
rect 1136 27671 1162 27735
rect 1226 27671 1252 27735
rect 1316 27671 1342 27735
rect 1406 27671 1432 27735
rect 1496 27671 1501 27735
rect 977 27655 1501 27671
rect 977 27591 982 27655
rect 1046 27591 1072 27655
rect 1136 27591 1162 27655
rect 1226 27591 1252 27655
rect 1316 27591 1342 27655
rect 1406 27591 1432 27655
rect 1496 27591 1501 27655
rect 977 27575 1501 27591
rect 977 27511 982 27575
rect 1046 27511 1072 27575
rect 1136 27511 1162 27575
rect 1226 27511 1252 27575
rect 1316 27511 1342 27575
rect 1406 27511 1432 27575
rect 1496 27511 1501 27575
rect 977 27495 1501 27511
rect 977 27431 982 27495
rect 1046 27431 1072 27495
rect 1136 27431 1162 27495
rect 1226 27431 1252 27495
rect 1316 27431 1342 27495
rect 977 27415 1384 27431
rect 977 27351 982 27415
rect 1046 27351 1072 27415
rect 1136 27351 1162 27415
rect 1226 27351 1252 27415
rect 1316 27351 1342 27415
rect 977 27335 1384 27351
rect 977 27271 982 27335
rect 1046 27271 1072 27335
rect 1136 27271 1162 27335
rect 1226 27271 1252 27335
rect 1316 27271 1342 27335
rect 977 27255 1384 27271
rect 977 27191 982 27255
rect 1046 27191 1072 27255
rect 1136 27191 1162 27255
rect 1226 27191 1252 27255
rect 1316 27191 1342 27255
rect 977 27175 1384 27191
rect 977 27111 982 27175
rect 1046 27111 1072 27175
rect 1136 27111 1162 27175
rect 1226 27111 1252 27175
rect 1316 27111 1342 27175
rect 977 27095 1384 27111
rect 977 27031 982 27095
rect 1046 27031 1072 27095
rect 1136 27031 1162 27095
rect 1226 27031 1252 27095
rect 1316 27031 1342 27095
rect 977 27015 1384 27031
rect 977 26951 982 27015
rect 1046 26951 1072 27015
rect 1136 26951 1162 27015
rect 1226 26951 1252 27015
rect 1316 26951 1342 27015
rect 977 26935 1384 26951
rect 977 26871 982 26935
rect 1046 26871 1072 26935
rect 1136 26871 1162 26935
rect 1226 26871 1252 26935
rect 1316 26871 1342 26935
rect 977 26855 1384 26871
rect 977 26791 982 26855
rect 1046 26791 1072 26855
rect 1136 26791 1162 26855
rect 1226 26791 1252 26855
rect 1316 26791 1342 26855
rect 977 26775 1384 26791
rect 977 26711 982 26775
rect 1046 26711 1072 26775
rect 1136 26711 1162 26775
rect 1226 26711 1252 26775
rect 1316 26711 1342 26775
rect 977 26695 1384 26711
rect 977 26631 982 26695
rect 1046 26631 1072 26695
rect 1136 26631 1162 26695
rect 1226 26631 1252 26695
rect 1316 26631 1342 26695
rect 1406 26631 1432 27495
rect 1496 26631 1501 27495
rect 977 26615 1501 26631
rect 977 26551 982 26615
rect 1046 26551 1072 26615
rect 1136 26551 1162 26615
rect 1226 26551 1252 26615
rect 1316 26551 1342 26615
rect 1406 26551 1432 26615
rect 1496 26551 1501 26615
rect 977 26535 1501 26551
rect 977 26471 982 26535
rect 1046 26471 1072 26535
rect 1136 26471 1162 26535
rect 1226 26471 1252 26535
rect 1316 26471 1342 26535
rect 1406 26471 1432 26535
rect 1496 26471 1501 26535
rect 977 26455 1501 26471
rect 977 26391 982 26455
rect 1046 26391 1072 26455
rect 1136 26391 1162 26455
rect 1226 26391 1252 26455
rect 1316 26391 1342 26455
rect 1406 26391 1432 26455
rect 1496 26391 1501 26455
rect 977 26375 1501 26391
rect 977 26311 982 26375
rect 1046 26311 1072 26375
rect 1136 26311 1162 26375
rect 1226 26311 1252 26375
rect 1316 26311 1342 26375
rect 1406 26311 1432 26375
rect 1496 26311 1501 26375
rect 977 26295 1501 26311
rect 977 26231 982 26295
rect 1046 26231 1072 26295
rect 1136 26231 1162 26295
rect 1226 26231 1252 26295
rect 1316 26231 1342 26295
rect 1406 26231 1432 26295
rect 1496 26231 1501 26295
rect 977 26215 1501 26231
rect 977 26151 982 26215
rect 1046 26151 1072 26215
rect 1136 26151 1162 26215
rect 1226 26151 1252 26215
rect 1316 26151 1342 26215
rect 1406 26151 1432 26215
rect 1496 26151 1501 26215
rect 977 26135 1501 26151
rect 977 26071 982 26135
rect 1046 26071 1072 26135
rect 1136 26071 1162 26135
rect 1226 26071 1252 26135
rect 1316 26071 1342 26135
rect 1406 26071 1432 26135
rect 1496 26071 1501 26135
rect 977 26055 1501 26071
rect 977 25991 982 26055
rect 1046 25991 1072 26055
rect 1136 25991 1162 26055
rect 1226 25991 1252 26055
rect 1316 25991 1342 26055
rect 1406 25991 1432 26055
rect 1496 25991 1501 26055
rect 977 25975 1501 25991
rect 977 25911 982 25975
rect 1046 25911 1072 25975
rect 1136 25911 1162 25975
rect 1226 25911 1252 25975
rect 1316 25911 1342 25975
rect 1406 25911 1432 25975
rect 1496 25911 1501 25975
rect 977 25895 1501 25911
rect 977 25831 982 25895
rect 1046 25831 1072 25895
rect 1136 25831 1162 25895
rect 1226 25831 1252 25895
rect 1316 25831 1342 25895
rect 1406 25831 1432 25895
rect 1496 25831 1501 25895
rect 977 25815 1501 25831
rect 977 25751 982 25815
rect 1046 25751 1072 25815
rect 1136 25751 1162 25815
rect 1226 25751 1252 25815
rect 1316 25751 1342 25815
rect 1406 25751 1432 25815
rect 1496 25751 1501 25815
rect 977 25735 1501 25751
rect 977 25671 982 25735
rect 1046 25671 1072 25735
rect 1136 25671 1162 25735
rect 1226 25671 1252 25735
rect 1316 25671 1342 25735
rect 1406 25671 1432 25735
rect 1496 25671 1501 25735
rect 977 25655 1501 25671
rect 977 25591 982 25655
rect 1046 25591 1072 25655
rect 1136 25591 1162 25655
rect 1226 25591 1252 25655
rect 1316 25591 1342 25655
rect 1406 25591 1432 25655
rect 1496 25591 1501 25655
rect 977 25575 1501 25591
rect 977 25511 982 25575
rect 1046 25511 1072 25575
rect 1136 25511 1162 25575
rect 1226 25511 1252 25575
rect 1316 25511 1342 25575
rect 1406 25511 1432 25575
rect 1496 25511 1501 25575
rect 977 25495 1501 25511
rect 977 25431 982 25495
rect 1046 25431 1072 25495
rect 1136 25431 1162 25495
rect 1226 25431 1252 25495
rect 1316 25431 1342 25495
rect 1406 25431 1432 25495
rect 1496 25431 1501 25495
rect 977 25415 1501 25431
rect 977 25351 982 25415
rect 1046 25351 1072 25415
rect 1136 25351 1162 25415
rect 1226 25351 1252 25415
rect 1316 25351 1342 25415
rect 1406 25351 1432 25415
rect 1496 25351 1501 25415
rect 977 25335 1501 25351
rect 977 25271 982 25335
rect 1046 25271 1072 25335
rect 1136 25271 1162 25335
rect 1226 25271 1252 25335
rect 1316 25271 1342 25335
rect 1406 25271 1432 25335
rect 1496 25271 1501 25335
rect 977 25255 1501 25271
rect 977 25191 982 25255
rect 1046 25191 1072 25255
rect 1136 25191 1162 25255
rect 1226 25191 1252 25255
rect 1316 25191 1342 25255
rect 1406 25191 1432 25255
rect 1496 25191 1501 25255
rect 977 25175 1501 25191
rect 977 25111 982 25175
rect 1046 25111 1072 25175
rect 1136 25111 1162 25175
rect 1226 25111 1252 25175
rect 1316 25111 1342 25175
rect 1406 25111 1432 25175
rect 1496 25111 1501 25175
rect 977 25095 1501 25111
rect 977 25031 982 25095
rect 1046 25031 1072 25095
rect 1136 25031 1162 25095
rect 1226 25031 1252 25095
rect 1316 25031 1342 25095
rect 1406 25031 1432 25095
rect 1496 25031 1501 25095
rect 977 25015 1501 25031
rect 977 24951 982 25015
rect 1046 24951 1072 25015
rect 1136 24951 1162 25015
rect 1226 24951 1252 25015
rect 1316 24951 1342 25015
rect 1406 24951 1432 25015
rect 1496 24951 1501 25015
rect 977 24935 1501 24951
rect 977 24871 982 24935
rect 1046 24871 1072 24935
rect 1136 24871 1162 24935
rect 1226 24871 1252 24935
rect 1316 24871 1342 24935
rect 1406 24871 1432 24935
rect 1496 24871 1501 24935
rect 977 24855 1501 24871
rect 977 24791 982 24855
rect 1046 24791 1072 24855
rect 1136 24791 1162 24855
rect 1226 24791 1252 24855
rect 1316 24791 1342 24855
rect 1406 24791 1432 24855
rect 1496 24791 1501 24855
rect 977 24775 1501 24791
rect 977 24711 982 24775
rect 1046 24711 1072 24775
rect 1136 24711 1162 24775
rect 1226 24711 1252 24775
rect 1316 24711 1342 24775
rect 1406 24711 1432 24775
rect 1496 24711 1501 24775
rect 977 24695 1501 24711
rect 977 24631 982 24695
rect 1046 24631 1072 24695
rect 1136 24631 1162 24695
rect 1226 24631 1252 24695
rect 1316 24631 1342 24695
rect 1406 24631 1432 24695
rect 1496 24631 1501 24695
rect 977 24615 1501 24631
rect 977 24551 982 24615
rect 1046 24551 1072 24615
rect 1136 24551 1162 24615
rect 1226 24551 1252 24615
rect 1316 24551 1342 24615
rect 1406 24551 1432 24615
rect 1496 24551 1501 24615
rect 977 24535 1501 24551
rect 977 24471 982 24535
rect 1046 24471 1072 24535
rect 1136 24471 1162 24535
rect 1226 24471 1252 24535
rect 1316 24471 1342 24535
rect 1406 24471 1432 24535
rect 1496 24471 1501 24535
rect 977 24455 1501 24471
rect 977 24391 982 24455
rect 1046 24391 1072 24455
rect 1136 24391 1162 24455
rect 1226 24391 1252 24455
rect 1316 24391 1342 24455
rect 1406 24391 1432 24455
rect 1496 24391 1501 24455
rect 977 24375 1501 24391
rect 977 24311 982 24375
rect 1046 24311 1072 24375
rect 1136 24311 1162 24375
rect 1226 24311 1252 24375
rect 1316 24311 1342 24375
rect 1406 24311 1432 24375
rect 1496 24311 1501 24375
rect 977 24295 1501 24311
rect 977 24231 982 24295
rect 1046 24231 1072 24295
rect 1136 24231 1162 24295
rect 1226 24231 1252 24295
rect 1316 24231 1342 24295
rect 1406 24231 1432 24295
rect 1496 24231 1501 24295
rect 977 24215 1501 24231
rect 977 24151 982 24215
rect 1046 24151 1072 24215
rect 1136 24151 1162 24215
rect 1226 24151 1252 24215
rect 1316 24151 1342 24215
rect 1406 24151 1432 24215
rect 1496 24151 1501 24215
rect 977 24135 1501 24151
rect 977 24071 982 24135
rect 1046 24071 1072 24135
rect 1136 24071 1162 24135
rect 1226 24071 1252 24135
rect 1316 24071 1342 24135
rect 1406 24071 1432 24135
rect 1496 24071 1501 24135
rect 977 24055 1501 24071
rect 977 23991 982 24055
rect 1046 23991 1072 24055
rect 1136 23991 1162 24055
rect 1226 23991 1252 24055
rect 1316 23991 1342 24055
rect 1406 23991 1432 24055
rect 1496 23991 1501 24055
rect 977 23975 1501 23991
rect 977 23911 982 23975
rect 1046 23911 1072 23975
rect 1136 23911 1162 23975
rect 1226 23911 1252 23975
rect 1316 23911 1342 23975
rect 1406 23911 1432 23975
rect 1496 23911 1501 23975
rect 977 23895 1501 23911
rect 977 23831 982 23895
rect 1046 23831 1072 23895
rect 1136 23831 1162 23895
rect 1226 23831 1252 23895
rect 1316 23831 1342 23895
rect 1406 23831 1432 23895
rect 1496 23831 1501 23895
rect 977 23815 1501 23831
rect 977 23751 982 23815
rect 1046 23751 1072 23815
rect 1136 23751 1162 23815
rect 1226 23751 1252 23815
rect 1316 23751 1342 23815
rect 1406 23751 1432 23815
rect 1496 23751 1501 23815
rect 977 23735 1501 23751
rect 977 23671 982 23735
rect 1046 23671 1072 23735
rect 1136 23671 1162 23735
rect 1226 23671 1252 23735
rect 1316 23671 1342 23735
rect 1406 23671 1432 23735
rect 1496 23671 1501 23735
rect 977 23655 1501 23671
rect 977 23591 982 23655
rect 1046 23591 1072 23655
rect 1136 23591 1162 23655
rect 1226 23591 1252 23655
rect 1316 23591 1342 23655
rect 1406 23591 1432 23655
rect 1496 23591 1501 23655
rect 977 23575 1501 23591
rect 977 23511 982 23575
rect 1046 23511 1072 23575
rect 1136 23511 1162 23575
rect 1226 23511 1252 23575
rect 1316 23511 1342 23575
rect 1406 23511 1432 23575
rect 1496 23511 1501 23575
rect 977 23495 1501 23511
rect 977 23431 982 23495
rect 1046 23431 1072 23495
rect 1136 23431 1162 23495
rect 1226 23431 1252 23495
rect 1316 23431 1342 23495
rect 1406 23431 1432 23495
rect 1496 23431 1501 23495
rect 977 23415 1501 23431
rect 977 23351 982 23415
rect 1046 23351 1072 23415
rect 1136 23351 1162 23415
rect 1226 23351 1252 23415
rect 1316 23351 1342 23415
rect 1406 23351 1432 23415
rect 1496 23351 1501 23415
rect 977 23335 1501 23351
rect 977 23271 982 23335
rect 1046 23271 1072 23335
rect 1136 23271 1162 23335
rect 1226 23271 1252 23335
rect 1316 23271 1342 23335
rect 1406 23271 1432 23335
rect 1496 23271 1501 23335
rect 977 23254 1501 23271
rect 977 23190 982 23254
rect 1046 23190 1072 23254
rect 1136 23190 1162 23254
rect 1226 23190 1252 23254
rect 1316 23190 1342 23254
rect 1406 23190 1432 23254
rect 1496 23190 1501 23254
rect 977 23173 1501 23190
rect 977 23109 982 23173
rect 1046 23109 1072 23173
rect 1136 23109 1162 23173
rect 1226 23109 1252 23173
rect 1316 23109 1342 23173
rect 1406 23109 1432 23173
rect 1496 23109 1501 23173
rect 977 23092 1501 23109
rect 977 23028 982 23092
rect 1046 23028 1072 23092
rect 1136 23028 1162 23092
rect 1226 23028 1252 23092
rect 1316 23028 1342 23092
rect 1406 23028 1432 23092
rect 1496 23028 1501 23092
rect 977 23011 1501 23028
rect 977 22947 982 23011
rect 1046 22947 1072 23011
rect 1136 22947 1162 23011
rect 1226 22947 1252 23011
rect 1316 22947 1342 23011
rect 1406 22947 1432 23011
rect 1496 22947 1501 23011
rect 977 22930 1501 22947
rect 977 22866 982 22930
rect 1046 22866 1072 22930
rect 1136 22866 1162 22930
rect 1226 22866 1252 22930
rect 1316 22866 1342 22930
rect 1406 22866 1432 22930
rect 1496 22866 1501 22930
rect 977 22849 1501 22866
rect 977 22785 982 22849
rect 1046 22785 1072 22849
rect 1136 22785 1162 22849
rect 1226 22785 1252 22849
rect 1316 22785 1342 22849
rect 1406 22785 1432 22849
rect 1496 22785 1501 22849
rect 977 22768 1501 22785
rect 977 22704 982 22768
rect 1046 22704 1072 22768
rect 1136 22704 1162 22768
rect 1226 22704 1252 22768
rect 1316 22704 1342 22768
rect 1406 22704 1432 22768
rect 1496 22704 1501 22768
rect 977 22687 1501 22704
rect 977 22623 982 22687
rect 1046 22623 1072 22687
rect 1136 22623 1162 22687
rect 1226 22623 1252 22687
rect 1316 22623 1342 22687
rect 1406 22623 1432 22687
rect 1496 22623 1501 22687
rect 977 22606 1501 22623
rect 977 22542 982 22606
rect 1046 22542 1072 22606
rect 1136 22542 1162 22606
rect 1226 22542 1252 22606
rect 1316 22542 1342 22606
rect 1406 22542 1432 22606
rect 1496 22542 1501 22606
rect 977 22525 1501 22542
rect 977 22461 982 22525
rect 1046 22461 1072 22525
rect 1136 22461 1162 22525
rect 1226 22461 1252 22525
rect 1316 22461 1342 22525
rect 1406 22461 1432 22525
rect 1496 22461 1501 22525
rect 977 22444 1501 22461
rect 977 22380 982 22444
rect 1046 22380 1072 22444
rect 1136 22380 1162 22444
rect 1226 22380 1252 22444
rect 1316 22380 1342 22444
rect 1406 22380 1432 22444
rect 1496 22380 1501 22444
rect 977 22363 1501 22380
rect 977 22299 982 22363
rect 1046 22299 1072 22363
rect 1136 22299 1162 22363
rect 1226 22299 1252 22363
rect 1316 22299 1342 22363
rect 1406 22299 1432 22363
rect 1496 22299 1501 22363
rect 977 22282 1501 22299
rect 977 22218 982 22282
rect 1046 22218 1072 22282
rect 1136 22218 1162 22282
rect 1226 22218 1252 22282
rect 1316 22218 1342 22282
rect 1406 22218 1432 22282
rect 1496 22218 1501 22282
rect 977 22201 1501 22218
rect 977 22137 982 22201
rect 1046 22137 1072 22201
rect 1136 22137 1162 22201
rect 1226 22137 1252 22201
rect 1316 22137 1342 22201
rect 1406 22137 1432 22201
rect 1496 22137 1501 22201
rect 977 22120 1501 22137
rect 977 22056 982 22120
rect 1046 22056 1072 22120
rect 1136 22056 1162 22120
rect 1226 22056 1252 22120
rect 1316 22056 1342 22120
rect 1406 22056 1432 22120
rect 1496 22056 1501 22120
rect 977 22039 1501 22056
rect 977 21975 982 22039
rect 1046 21975 1072 22039
rect 1136 21975 1162 22039
rect 1226 21975 1252 22039
rect 1316 21975 1342 22039
rect 1406 21975 1432 22039
rect 1496 21975 1501 22039
rect 977 21958 1501 21975
rect 977 21894 982 21958
rect 1046 21894 1072 21958
rect 1136 21894 1162 21958
rect 1226 21894 1252 21958
rect 1316 21894 1342 21958
rect 1406 21894 1432 21958
rect 1496 21894 1501 21958
rect 977 21877 1501 21894
rect 977 21813 982 21877
rect 1046 21813 1072 21877
rect 1136 21813 1162 21877
rect 1226 21813 1252 21877
rect 1316 21813 1342 21877
rect 1406 21813 1432 21877
rect 1496 21813 1501 21877
rect 977 21796 1501 21813
rect 977 21732 982 21796
rect 1046 21732 1072 21796
rect 1136 21732 1162 21796
rect 1226 21732 1252 21796
rect 1316 21732 1342 21796
rect 1406 21732 1432 21796
rect 1496 21732 1501 21796
rect 977 21715 1501 21732
rect 977 21651 982 21715
rect 1046 21651 1072 21715
rect 1136 21651 1162 21715
rect 1226 21651 1252 21715
rect 1316 21651 1342 21715
rect 1406 21651 1432 21715
rect 1496 21651 1501 21715
rect 977 21634 1501 21651
rect 977 21570 982 21634
rect 1046 21570 1072 21634
rect 1136 21570 1162 21634
rect 1226 21570 1252 21634
rect 1316 21570 1342 21634
rect 1406 21570 1432 21634
rect 1496 21570 1501 21634
rect 977 21553 1501 21570
rect 977 21489 982 21553
rect 1046 21489 1072 21553
rect 1136 21489 1162 21553
rect 1226 21489 1252 21553
rect 1316 21489 1342 21553
rect 1406 21489 1432 21553
rect 1496 21489 1501 21553
rect 977 21472 1501 21489
rect 977 21408 982 21472
rect 1046 21408 1072 21472
rect 1136 21408 1162 21472
rect 1226 21408 1252 21472
rect 1316 21408 1342 21472
rect 1406 21408 1432 21472
rect 1496 21408 1501 21472
rect 977 21391 1501 21408
rect 977 21327 982 21391
rect 1046 21327 1072 21391
rect 1136 21327 1162 21391
rect 1226 21327 1252 21391
rect 1316 21327 1342 21391
rect 1406 21327 1432 21391
rect 1496 21327 1501 21391
rect 977 21310 1501 21327
rect 977 21246 982 21310
rect 1046 21246 1072 21310
rect 1136 21246 1162 21310
rect 1226 21246 1252 21310
rect 1316 21246 1342 21310
rect 1406 21246 1432 21310
rect 1496 21246 1501 21310
rect 977 21229 1501 21246
rect 977 21165 982 21229
rect 1046 21165 1072 21229
rect 1136 21165 1162 21229
rect 1226 21165 1252 21229
rect 1316 21165 1342 21229
rect 1406 21165 1432 21229
rect 1496 21165 1501 21229
rect 977 21148 1501 21165
rect 977 21084 982 21148
rect 1046 21084 1072 21148
rect 1136 21084 1162 21148
rect 1226 21084 1252 21148
rect 1316 21084 1342 21148
rect 1406 21084 1432 21148
rect 1496 21084 1501 21148
rect 977 21067 1501 21084
rect 977 21003 982 21067
rect 1046 21003 1072 21067
rect 1136 21003 1162 21067
rect 1226 21003 1252 21067
rect 1316 21003 1342 21067
rect 1406 21003 1432 21067
rect 1496 21003 1501 21067
rect 977 20986 1501 21003
rect 977 20922 982 20986
rect 1046 20922 1072 20986
rect 1136 20922 1162 20986
rect 1226 20922 1252 20986
rect 1316 20922 1342 20986
rect 1406 20922 1432 20986
rect 1496 20958 1501 20986
rect 13515 33095 14039 33096
rect 13515 33031 13520 33095
rect 13584 33031 13610 33095
rect 13674 33031 13700 33095
rect 13764 33031 13790 33095
rect 13854 33031 13880 33095
rect 13944 33031 13970 33095
rect 14034 33031 14039 33095
rect 13515 33015 14039 33031
rect 13515 32951 13520 33015
rect 13584 32951 13610 33015
rect 13674 32951 13700 33015
rect 13764 32951 13790 33015
rect 13854 32951 13880 33015
rect 13944 32951 13970 33015
rect 14034 32951 14039 33015
rect 13515 32935 14039 32951
rect 13515 32871 13520 32935
rect 13584 32871 13610 32935
rect 13674 32871 13700 32935
rect 13764 32871 13790 32935
rect 13854 32871 13880 32935
rect 13944 32871 13970 32935
rect 14034 32871 14039 32935
rect 13515 32855 14039 32871
rect 13515 32791 13520 32855
rect 13584 32791 13610 32855
rect 13674 32791 13700 32855
rect 13764 32791 13790 32855
rect 13854 32791 13880 32855
rect 13944 32791 13970 32855
rect 14034 32791 14039 32855
rect 13515 32775 14039 32791
rect 13515 32711 13520 32775
rect 13584 32711 13610 32775
rect 13674 32711 13700 32775
rect 13764 32711 13790 32775
rect 13854 32711 13880 32775
rect 13944 32711 13970 32775
rect 14034 32711 14039 32775
rect 13515 32695 14039 32711
rect 13515 32631 13520 32695
rect 13584 32631 13610 32695
rect 13674 32631 13700 32695
rect 13764 32631 13790 32695
rect 13854 32631 13880 32695
rect 13944 32631 13970 32695
rect 14034 32631 14039 32695
rect 13515 32615 14039 32631
rect 13515 32551 13520 32615
rect 13584 32551 13610 32615
rect 13674 32551 13700 32615
rect 13764 32551 13790 32615
rect 13854 32551 13880 32615
rect 13944 32551 13970 32615
rect 14034 32551 14039 32615
rect 13515 32535 14039 32551
rect 13515 32471 13520 32535
rect 13584 32471 13610 32535
rect 13674 32471 13700 32535
rect 13764 32471 13790 32535
rect 13854 32471 13880 32535
rect 13944 32471 13970 32535
rect 14034 32471 14039 32535
rect 13515 32455 14039 32471
rect 13515 32391 13520 32455
rect 13584 32391 13610 32455
rect 13674 32391 13700 32455
rect 13764 32391 13790 32455
rect 13854 32391 13880 32455
rect 13944 32391 13970 32455
rect 14034 32391 14039 32455
rect 13515 32375 14039 32391
rect 13515 32311 13520 32375
rect 13584 32311 13610 32375
rect 13674 32311 13700 32375
rect 13764 32311 13790 32375
rect 13854 32311 13880 32375
rect 13944 32311 13970 32375
rect 14034 32311 14039 32375
rect 13515 32295 14039 32311
rect 13515 32231 13520 32295
rect 13584 32231 13610 32295
rect 13674 32231 13700 32295
rect 13764 32231 13790 32295
rect 13854 32231 13880 32295
rect 13944 32231 13970 32295
rect 14034 32231 14039 32295
rect 13515 32215 14039 32231
rect 13515 32151 13520 32215
rect 13584 32151 13610 32215
rect 13674 32151 13700 32215
rect 13764 32151 13790 32215
rect 13854 32151 13880 32215
rect 13944 32151 13970 32215
rect 14034 32151 14039 32215
rect 13515 32135 14039 32151
rect 13515 32071 13520 32135
rect 13584 32071 13610 32135
rect 13674 32071 13700 32135
rect 13764 32071 13790 32135
rect 13854 32071 13880 32135
rect 13944 32071 13970 32135
rect 14034 32071 14039 32135
rect 13515 32055 14039 32071
rect 13515 31991 13520 32055
rect 13584 31991 13610 32055
rect 13674 31991 13700 32055
rect 13764 31991 13790 32055
rect 13854 31991 13880 32055
rect 13944 31991 13970 32055
rect 14034 31991 14039 32055
rect 13515 31975 14039 31991
rect 13515 31911 13520 31975
rect 13584 31911 13610 31975
rect 13674 31911 13700 31975
rect 13764 31911 13790 31975
rect 13854 31911 13880 31975
rect 13944 31911 13970 31975
rect 14034 31911 14039 31975
rect 13515 31895 14039 31911
rect 13515 31831 13520 31895
rect 13584 31831 13610 31895
rect 13674 31831 13700 31895
rect 13764 31831 13790 31895
rect 13854 31831 13880 31895
rect 13944 31831 13970 31895
rect 14034 31831 14039 31895
rect 13515 31815 14039 31831
rect 13515 31751 13520 31815
rect 13584 31751 13610 31815
rect 13674 31751 13700 31815
rect 13764 31751 13790 31815
rect 13854 31751 13880 31815
rect 13944 31751 13970 31815
rect 14034 31751 14039 31815
rect 13515 31735 14039 31751
rect 13515 31671 13520 31735
rect 13584 31671 13610 31735
rect 13674 31671 13700 31735
rect 13764 31671 13790 31735
rect 13854 31671 13880 31735
rect 13944 31671 13970 31735
rect 14034 31671 14039 31735
rect 13515 31655 14039 31671
rect 13515 31591 13520 31655
rect 13584 31591 13610 31655
rect 13674 31591 13700 31655
rect 13764 31591 13790 31655
rect 13854 31591 13880 31655
rect 13944 31591 13970 31655
rect 14034 31591 14039 31655
rect 13515 31575 14039 31591
rect 13515 31511 13520 31575
rect 13584 31511 13610 31575
rect 13674 31511 13700 31575
rect 13764 31511 13790 31575
rect 13854 31511 13880 31575
rect 13944 31511 13970 31575
rect 14034 31511 14039 31575
rect 13515 31495 14039 31511
rect 13515 31431 13520 31495
rect 13584 31431 13610 31495
rect 13674 31431 13700 31495
rect 13764 31431 13790 31495
rect 13854 31431 13880 31495
rect 13944 31431 13970 31495
rect 14034 31431 14039 31495
rect 13515 31415 14039 31431
rect 13515 31351 13520 31415
rect 13584 31351 13610 31415
rect 13674 31351 13700 31415
rect 13764 31351 13790 31415
rect 13854 31351 13880 31415
rect 13944 31351 13970 31415
rect 14034 31351 14039 31415
rect 13515 31335 14039 31351
rect 13515 31271 13520 31335
rect 13584 31271 13610 31335
rect 13674 31271 13700 31335
rect 13764 31271 13790 31335
rect 13854 31271 13880 31335
rect 13944 31271 13970 31335
rect 14034 31271 14039 31335
rect 13515 31255 14039 31271
rect 13515 31191 13520 31255
rect 13584 31191 13610 31255
rect 13674 31191 13700 31255
rect 13764 31191 13790 31255
rect 13854 31191 13880 31255
rect 13944 31191 13970 31255
rect 14034 31191 14039 31255
rect 13515 31175 14039 31191
rect 13515 31111 13520 31175
rect 13584 31111 13610 31175
rect 13674 31111 13700 31175
rect 13764 31111 13790 31175
rect 13854 31111 13880 31175
rect 13944 31111 13970 31175
rect 14034 31111 14039 31175
rect 13515 31095 14039 31111
rect 13515 31031 13520 31095
rect 13584 31031 13610 31095
rect 13674 31031 13700 31095
rect 13764 31031 13790 31095
rect 13854 31031 13880 31095
rect 13944 31031 13970 31095
rect 14034 31031 14039 31095
rect 13515 31015 14039 31031
rect 13515 30951 13520 31015
rect 13584 30951 13610 31015
rect 13674 30951 13700 31015
rect 13764 30951 13790 31015
rect 13854 30951 13880 31015
rect 13944 30951 13970 31015
rect 14034 30951 14039 31015
rect 13515 30935 14039 30951
rect 13515 30871 13520 30935
rect 13584 30871 13610 30935
rect 13674 30871 13700 30935
rect 13764 30871 13790 30935
rect 13854 30871 13880 30935
rect 13944 30871 13970 30935
rect 14034 30871 14039 30935
rect 13515 30855 14039 30871
rect 13515 30791 13520 30855
rect 13584 30791 13610 30855
rect 13674 30791 13700 30855
rect 13764 30791 13790 30855
rect 13854 30791 13880 30855
rect 13944 30791 13970 30855
rect 14034 30791 14039 30855
rect 13515 30775 14039 30791
rect 13515 30711 13520 30775
rect 13584 30711 13610 30775
rect 13674 30711 13700 30775
rect 13764 30711 13790 30775
rect 13854 30711 13880 30775
rect 13944 30711 13970 30775
rect 14034 30711 14039 30775
rect 13515 30695 14039 30711
rect 13515 30631 13520 30695
rect 13584 30631 13610 30695
rect 13674 30631 13700 30695
rect 13764 30631 13790 30695
rect 13854 30631 13880 30695
rect 13944 30631 13970 30695
rect 14034 30631 14039 30695
rect 13515 30615 14039 30631
rect 13515 30551 13520 30615
rect 13584 30551 13610 30615
rect 13674 30551 13700 30615
rect 13764 30551 13790 30615
rect 13854 30551 13880 30615
rect 13944 30551 13970 30615
rect 14034 30551 14039 30615
rect 13515 30535 14039 30551
rect 13515 30471 13520 30535
rect 13584 30471 13610 30535
rect 13674 30471 13700 30535
rect 13764 30471 13790 30535
rect 13854 30471 13880 30535
rect 13944 30471 13970 30535
rect 14034 30471 14039 30535
rect 13515 30455 14039 30471
rect 13515 30391 13520 30455
rect 13584 30391 13610 30455
rect 13674 30391 13700 30455
rect 13764 30391 13790 30455
rect 13854 30391 13880 30455
rect 13944 30391 13970 30455
rect 14034 30391 14039 30455
rect 13515 30375 14039 30391
rect 13515 30311 13520 30375
rect 13584 30311 13610 30375
rect 13674 30311 13700 30375
rect 13764 30311 13790 30375
rect 13854 30311 13880 30375
rect 13944 30311 13970 30375
rect 14034 30311 14039 30375
rect 13515 30295 14039 30311
rect 13515 30231 13520 30295
rect 13584 30231 13610 30295
rect 13674 30231 13700 30295
rect 13764 30231 13790 30295
rect 13854 30231 13880 30295
rect 13944 30231 13970 30295
rect 14034 30231 14039 30295
rect 13515 30215 14039 30231
rect 13515 30151 13520 30215
rect 13584 30151 13610 30215
rect 13674 30151 13700 30215
rect 13764 30151 13790 30215
rect 13854 30151 13880 30215
rect 13944 30151 13970 30215
rect 14034 30151 14039 30215
rect 13515 30135 14039 30151
rect 13515 30071 13520 30135
rect 13584 30071 13610 30135
rect 13674 30071 13700 30135
rect 13764 30071 13790 30135
rect 13854 30071 13880 30135
rect 13944 30071 13970 30135
rect 14034 30071 14039 30135
rect 13515 30055 14039 30071
rect 13515 29991 13520 30055
rect 13584 29991 13610 30055
rect 13674 29991 13700 30055
rect 13764 29991 13790 30055
rect 13854 29991 13880 30055
rect 13944 29991 13970 30055
rect 14034 29991 14039 30055
rect 13515 29975 14039 29991
rect 13515 29911 13520 29975
rect 13584 29911 13610 29975
rect 13674 29911 13700 29975
rect 13764 29911 13790 29975
rect 13854 29911 13880 29975
rect 13944 29911 13970 29975
rect 14034 29911 14039 29975
rect 13515 29895 14039 29911
rect 13515 29831 13520 29895
rect 13584 29831 13610 29895
rect 13674 29831 13700 29895
rect 13764 29831 13790 29895
rect 13854 29831 13880 29895
rect 13944 29831 13970 29895
rect 14034 29831 14039 29895
rect 13515 29815 14039 29831
rect 13515 29751 13520 29815
rect 13584 29751 13610 29815
rect 13674 29751 13700 29815
rect 13764 29751 13790 29815
rect 13854 29751 13880 29815
rect 13944 29751 13970 29815
rect 14034 29751 14039 29815
rect 13515 29735 14039 29751
rect 13515 29671 13520 29735
rect 13584 29671 13610 29735
rect 13674 29671 13700 29735
rect 13764 29671 13790 29735
rect 13854 29671 13880 29735
rect 13944 29671 13970 29735
rect 14034 29671 14039 29735
rect 13515 29655 14039 29671
rect 13515 29591 13520 29655
rect 13584 29591 13610 29655
rect 13674 29591 13700 29655
rect 13764 29591 13790 29655
rect 13854 29591 13880 29655
rect 13944 29591 13970 29655
rect 14034 29591 14039 29655
rect 13515 29575 14039 29591
rect 13515 29511 13520 29575
rect 13584 29511 13610 29575
rect 13674 29511 13700 29575
rect 13764 29511 13790 29575
rect 13854 29511 13880 29575
rect 13944 29511 13970 29575
rect 14034 29511 14039 29575
rect 13515 29495 14039 29511
rect 13515 29431 13520 29495
rect 13584 29431 13610 29495
rect 13674 29431 13700 29495
rect 13764 29431 13790 29495
rect 13854 29431 13880 29495
rect 13944 29431 13970 29495
rect 14034 29431 14039 29495
rect 13515 29415 14039 29431
rect 13515 29351 13520 29415
rect 13584 29351 13610 29415
rect 13674 29351 13700 29415
rect 13764 29351 13790 29415
rect 13854 29351 13880 29415
rect 13944 29351 13970 29415
rect 14034 29351 14039 29415
rect 13515 29335 14039 29351
rect 13515 29271 13520 29335
rect 13584 29271 13610 29335
rect 13674 29271 13700 29335
rect 13764 29271 13790 29335
rect 13854 29271 13880 29335
rect 13944 29271 13970 29335
rect 14034 29271 14039 29335
rect 13515 29255 14039 29271
rect 13515 29191 13520 29255
rect 13584 29191 13610 29255
rect 13674 29191 13700 29255
rect 13764 29191 13790 29255
rect 13854 29191 13880 29255
rect 13944 29191 13970 29255
rect 14034 29191 14039 29255
rect 13515 29175 14039 29191
rect 13515 29111 13520 29175
rect 13584 29111 13610 29175
rect 13674 29111 13700 29175
rect 13764 29111 13790 29175
rect 13854 29111 13880 29175
rect 13944 29111 13970 29175
rect 14034 29111 14039 29175
rect 13515 29095 14039 29111
rect 13515 29031 13520 29095
rect 13584 29031 13610 29095
rect 13674 29031 13700 29095
rect 13764 29031 13790 29095
rect 13854 29031 13880 29095
rect 13944 29031 13970 29095
rect 14034 29031 14039 29095
rect 13515 29015 14039 29031
rect 13515 28951 13520 29015
rect 13584 28951 13610 29015
rect 13674 28951 13700 29015
rect 13764 28951 13790 29015
rect 13854 28951 13880 29015
rect 13944 28951 13970 29015
rect 14034 28951 14039 29015
rect 13515 28935 14039 28951
rect 13515 28871 13520 28935
rect 13584 28871 13610 28935
rect 13674 28871 13700 28935
rect 13764 28871 13790 28935
rect 13854 28871 13880 28935
rect 13944 28871 13970 28935
rect 14034 28871 14039 28935
rect 13515 28855 14039 28871
rect 13515 28791 13520 28855
rect 13584 28791 13610 28855
rect 13674 28791 13700 28855
rect 13764 28791 13790 28855
rect 13854 28791 13880 28855
rect 13944 28791 13970 28855
rect 14034 28791 14039 28855
rect 13515 28775 14039 28791
rect 13515 28711 13520 28775
rect 13584 28711 13610 28775
rect 13674 28711 13700 28775
rect 13764 28711 13790 28775
rect 13854 28711 13880 28775
rect 13944 28711 13970 28775
rect 14034 28711 14039 28775
rect 13515 28695 14039 28711
rect 13515 28631 13520 28695
rect 13584 28631 13610 28695
rect 13674 28631 13700 28695
rect 13764 28631 13790 28695
rect 13854 28631 13880 28695
rect 13944 28631 13970 28695
rect 14034 28631 14039 28695
rect 13515 28615 14039 28631
rect 13515 28551 13520 28615
rect 13584 28551 13610 28615
rect 13674 28551 13700 28615
rect 13764 28551 13790 28615
rect 13854 28551 13880 28615
rect 13944 28551 13970 28615
rect 14034 28551 14039 28615
rect 13515 28535 14039 28551
rect 13515 28471 13520 28535
rect 13584 28471 13610 28535
rect 13674 28471 13700 28535
rect 13764 28471 13790 28535
rect 13854 28471 13880 28535
rect 13944 28471 13970 28535
rect 14034 28471 14039 28535
rect 13515 28455 14039 28471
rect 13515 28391 13520 28455
rect 13584 28391 13610 28455
rect 13674 28391 13700 28455
rect 13764 28391 13790 28455
rect 13854 28391 13880 28455
rect 13944 28391 13970 28455
rect 14034 28391 14039 28455
rect 13515 28375 14039 28391
rect 13515 28311 13520 28375
rect 13584 28311 13610 28375
rect 13674 28311 13700 28375
rect 13764 28311 13790 28375
rect 13854 28311 13880 28375
rect 13944 28311 13970 28375
rect 14034 28311 14039 28375
rect 13515 28295 14039 28311
rect 13515 28231 13520 28295
rect 13584 28231 13610 28295
rect 13674 28231 13700 28295
rect 13764 28231 13790 28295
rect 13854 28231 13880 28295
rect 13944 28231 13970 28295
rect 14034 28231 14039 28295
rect 13515 28215 14039 28231
rect 13515 28151 13520 28215
rect 13584 28151 13610 28215
rect 13674 28151 13700 28215
rect 13764 28151 13790 28215
rect 13854 28151 13880 28215
rect 13944 28151 13970 28215
rect 14034 28151 14039 28215
rect 13515 28135 14039 28151
rect 13515 28071 13520 28135
rect 13584 28071 13610 28135
rect 13674 28071 13700 28135
rect 13764 28071 13790 28135
rect 13854 28071 13880 28135
rect 13944 28071 13970 28135
rect 14034 28071 14039 28135
rect 13515 28055 14039 28071
rect 13515 27991 13520 28055
rect 13584 27991 13610 28055
rect 13674 27991 13700 28055
rect 13764 27991 13790 28055
rect 13854 27991 13880 28055
rect 13944 27991 13970 28055
rect 14034 27991 14039 28055
rect 13515 27975 14039 27991
rect 13515 27911 13520 27975
rect 13584 27911 13610 27975
rect 13674 27911 13700 27975
rect 13764 27911 13790 27975
rect 13854 27911 13880 27975
rect 13944 27911 13970 27975
rect 14034 27911 14039 27975
rect 13515 27895 14039 27911
rect 13515 27831 13520 27895
rect 13584 27831 13610 27895
rect 13674 27831 13700 27895
rect 13764 27831 13790 27895
rect 13854 27831 13880 27895
rect 13944 27831 13970 27895
rect 14034 27831 14039 27895
rect 13515 27815 14039 27831
rect 13515 27751 13520 27815
rect 13584 27751 13610 27815
rect 13674 27751 13700 27815
rect 13764 27751 13790 27815
rect 13854 27751 13880 27815
rect 13944 27751 13970 27815
rect 14034 27751 14039 27815
rect 13515 27735 14039 27751
rect 13515 27671 13520 27735
rect 13584 27671 13610 27735
rect 13674 27671 13700 27735
rect 13764 27671 13790 27735
rect 13854 27671 13880 27735
rect 13944 27671 13970 27735
rect 14034 27671 14039 27735
rect 13515 27655 14039 27671
rect 13515 27591 13520 27655
rect 13584 27591 13610 27655
rect 13674 27591 13700 27655
rect 13764 27591 13790 27655
rect 13854 27591 13880 27655
rect 13944 27591 13970 27655
rect 14034 27591 14039 27655
rect 13515 27575 14039 27591
rect 13515 27511 13520 27575
rect 13584 27511 13610 27575
rect 13674 27511 13700 27575
rect 13764 27511 13790 27575
rect 13854 27511 13880 27575
rect 13944 27511 13970 27575
rect 14034 27511 14039 27575
rect 13515 27495 14039 27511
rect 13515 27431 13520 27495
rect 13584 27431 13610 27495
rect 13674 27431 13700 27495
rect 13764 27431 13790 27495
rect 13854 27431 13880 27495
rect 13944 27431 13970 27495
rect 14034 27431 14039 27495
rect 13515 27415 14039 27431
rect 13515 27351 13520 27415
rect 13584 27351 13610 27415
rect 13674 27351 13700 27415
rect 13764 27351 13790 27415
rect 13854 27351 13880 27415
rect 13944 27351 13970 27415
rect 14034 27351 14039 27415
rect 13515 27335 14039 27351
rect 13515 27271 13520 27335
rect 13584 27271 13610 27335
rect 13674 27271 13700 27335
rect 13764 27271 13790 27335
rect 13854 27271 13880 27335
rect 13944 27271 13970 27335
rect 14034 27271 14039 27335
rect 13515 27255 14039 27271
rect 13515 27191 13520 27255
rect 13584 27191 13610 27255
rect 13674 27191 13700 27255
rect 13764 27191 13790 27255
rect 13854 27191 13880 27255
rect 13944 27191 13970 27255
rect 14034 27191 14039 27255
rect 13515 27175 14039 27191
rect 13515 27111 13520 27175
rect 13584 27111 13610 27175
rect 13674 27111 13700 27175
rect 13764 27111 13790 27175
rect 13854 27111 13880 27175
rect 13944 27111 13970 27175
rect 14034 27111 14039 27175
rect 13515 27095 14039 27111
rect 13515 27031 13520 27095
rect 13584 27031 13610 27095
rect 13674 27031 13700 27095
rect 13764 27031 13790 27095
rect 13854 27031 13880 27095
rect 13944 27031 13970 27095
rect 14034 27031 14039 27095
rect 13515 27015 14039 27031
rect 13515 26951 13520 27015
rect 13584 26951 13610 27015
rect 13674 26951 13700 27015
rect 13764 26951 13790 27015
rect 13854 26951 13880 27015
rect 13944 26951 13970 27015
rect 14034 26951 14039 27015
rect 13515 26935 14039 26951
rect 13515 26871 13520 26935
rect 13584 26871 13610 26935
rect 13674 26871 13700 26935
rect 13764 26871 13790 26935
rect 13854 26871 13880 26935
rect 13944 26871 13970 26935
rect 14034 26871 14039 26935
rect 13515 26855 14039 26871
rect 13515 26791 13520 26855
rect 13584 26791 13610 26855
rect 13674 26791 13700 26855
rect 13764 26791 13790 26855
rect 13854 26791 13880 26855
rect 13944 26791 13970 26855
rect 14034 26791 14039 26855
rect 13515 26775 14039 26791
rect 13515 26711 13520 26775
rect 13584 26711 13610 26775
rect 13674 26711 13700 26775
rect 13764 26711 13790 26775
rect 13854 26711 13880 26775
rect 13944 26711 13970 26775
rect 14034 26711 14039 26775
rect 13515 26695 14039 26711
rect 13515 26631 13520 26695
rect 13584 26631 13610 26695
rect 13674 26631 13700 26695
rect 13764 26631 13790 26695
rect 13854 26631 13880 26695
rect 13944 26631 13970 26695
rect 14034 26631 14039 26695
rect 13515 26615 14039 26631
rect 13515 26551 13520 26615
rect 13584 26551 13610 26615
rect 13674 26551 13700 26615
rect 13764 26551 13790 26615
rect 13854 26551 13880 26615
rect 13944 26551 13970 26615
rect 14034 26551 14039 26615
rect 13515 26535 14039 26551
rect 13515 26471 13520 26535
rect 13584 26471 13610 26535
rect 13674 26471 13700 26535
rect 13764 26471 13790 26535
rect 13854 26471 13880 26535
rect 13944 26471 13970 26535
rect 14034 26471 14039 26535
rect 13515 26455 14039 26471
rect 13515 26391 13520 26455
rect 13584 26391 13610 26455
rect 13674 26391 13700 26455
rect 13764 26391 13790 26455
rect 13854 26391 13880 26455
rect 13944 26391 13970 26455
rect 14034 26391 14039 26455
rect 13515 26375 14039 26391
rect 13515 26311 13520 26375
rect 13584 26311 13610 26375
rect 13674 26311 13700 26375
rect 13764 26311 13790 26375
rect 13854 26311 13880 26375
rect 13944 26311 13970 26375
rect 14034 26311 14039 26375
rect 13515 26295 14039 26311
rect 13515 26231 13520 26295
rect 13584 26231 13610 26295
rect 13674 26231 13700 26295
rect 13764 26231 13790 26295
rect 13854 26231 13880 26295
rect 13944 26231 13970 26295
rect 14034 26231 14039 26295
rect 13515 26215 14039 26231
rect 13515 26151 13520 26215
rect 13584 26151 13610 26215
rect 13674 26151 13700 26215
rect 13764 26151 13790 26215
rect 13854 26151 13880 26215
rect 13944 26151 13970 26215
rect 14034 26151 14039 26215
rect 13515 26135 14039 26151
rect 13515 26071 13520 26135
rect 13584 26071 13610 26135
rect 13674 26071 13700 26135
rect 13764 26071 13790 26135
rect 13854 26071 13880 26135
rect 13944 26071 13970 26135
rect 14034 26071 14039 26135
rect 13515 26055 14039 26071
rect 13515 25991 13520 26055
rect 13584 25991 13610 26055
rect 13674 25991 13700 26055
rect 13764 25991 13790 26055
rect 13854 25991 13880 26055
rect 13944 25991 13970 26055
rect 14034 25991 14039 26055
rect 13515 25975 14039 25991
rect 13515 25911 13520 25975
rect 13584 25911 13610 25975
rect 13674 25911 13700 25975
rect 13764 25911 13790 25975
rect 13854 25911 13880 25975
rect 13944 25911 13970 25975
rect 14034 25911 14039 25975
rect 13515 25895 14039 25911
rect 13515 25831 13520 25895
rect 13584 25831 13610 25895
rect 13674 25831 13700 25895
rect 13764 25831 13790 25895
rect 13854 25831 13880 25895
rect 13944 25831 13970 25895
rect 14034 25831 14039 25895
rect 13515 25815 14039 25831
rect 13515 25751 13520 25815
rect 13584 25751 13610 25815
rect 13674 25751 13700 25815
rect 13764 25751 13790 25815
rect 13854 25751 13880 25815
rect 13944 25751 13970 25815
rect 14034 25751 14039 25815
rect 13515 25735 14039 25751
rect 13515 25671 13520 25735
rect 13584 25671 13610 25735
rect 13674 25671 13700 25735
rect 13764 25671 13790 25735
rect 13854 25671 13880 25735
rect 13944 25671 13970 25735
rect 14034 25671 14039 25735
rect 13515 25655 14039 25671
rect 13515 25591 13520 25655
rect 13584 25591 13610 25655
rect 13674 25591 13700 25655
rect 13764 25591 13790 25655
rect 13854 25591 13880 25655
rect 13944 25591 13970 25655
rect 14034 25591 14039 25655
rect 13515 25575 14039 25591
rect 13515 25511 13520 25575
rect 13584 25511 13610 25575
rect 13674 25511 13700 25575
rect 13764 25511 13790 25575
rect 13854 25511 13880 25575
rect 13944 25511 13970 25575
rect 14034 25511 14039 25575
rect 13515 25495 14039 25511
rect 13515 25431 13520 25495
rect 13584 25431 13610 25495
rect 13674 25431 13700 25495
rect 13764 25431 13790 25495
rect 13854 25431 13880 25495
rect 13944 25431 13970 25495
rect 14034 25431 14039 25495
rect 13515 25415 14039 25431
rect 13515 25351 13520 25415
rect 13584 25351 13610 25415
rect 13674 25351 13700 25415
rect 13764 25351 13790 25415
rect 13854 25351 13880 25415
rect 13944 25351 13970 25415
rect 14034 25351 14039 25415
rect 13515 25335 14039 25351
rect 13515 25271 13520 25335
rect 13584 25271 13610 25335
rect 13674 25271 13700 25335
rect 13764 25271 13790 25335
rect 13854 25271 13880 25335
rect 13944 25271 13970 25335
rect 14034 25271 14039 25335
rect 13515 25255 14039 25271
rect 13515 25191 13520 25255
rect 13584 25191 13610 25255
rect 13674 25191 13700 25255
rect 13764 25191 13790 25255
rect 13854 25191 13880 25255
rect 13944 25191 13970 25255
rect 14034 25191 14039 25255
rect 13515 25175 14039 25191
rect 13515 25111 13520 25175
rect 13584 25111 13610 25175
rect 13674 25111 13700 25175
rect 13764 25111 13790 25175
rect 13854 25111 13880 25175
rect 13944 25111 13970 25175
rect 14034 25111 14039 25175
rect 13515 25095 14039 25111
rect 13515 25031 13520 25095
rect 13584 25031 13610 25095
rect 13674 25031 13700 25095
rect 13764 25031 13790 25095
rect 13854 25031 13880 25095
rect 13944 25031 13970 25095
rect 14034 25031 14039 25095
rect 13515 25015 14039 25031
rect 13515 24951 13520 25015
rect 13584 24951 13610 25015
rect 13674 24951 13700 25015
rect 13764 24951 13790 25015
rect 13854 24951 13880 25015
rect 13944 24951 13970 25015
rect 14034 24951 14039 25015
rect 13515 24935 14039 24951
rect 13515 24871 13520 24935
rect 13584 24871 13610 24935
rect 13674 24871 13700 24935
rect 13764 24871 13790 24935
rect 13854 24871 13880 24935
rect 13944 24871 13970 24935
rect 14034 24871 14039 24935
rect 13515 24855 14039 24871
rect 13515 24791 13520 24855
rect 13584 24791 13610 24855
rect 13674 24791 13700 24855
rect 13764 24791 13790 24855
rect 13854 24791 13880 24855
rect 13944 24791 13970 24855
rect 14034 24791 14039 24855
rect 13515 24775 14039 24791
rect 13515 24711 13520 24775
rect 13584 24711 13610 24775
rect 13674 24711 13700 24775
rect 13764 24711 13790 24775
rect 13854 24711 13880 24775
rect 13944 24711 13970 24775
rect 14034 24711 14039 24775
rect 13515 24695 14039 24711
rect 13515 24631 13520 24695
rect 13584 24631 13610 24695
rect 13674 24631 13700 24695
rect 13764 24631 13790 24695
rect 13854 24631 13880 24695
rect 13944 24631 13970 24695
rect 14034 24631 14039 24695
rect 13515 24615 14039 24631
rect 13515 24551 13520 24615
rect 13584 24551 13610 24615
rect 13674 24551 13700 24615
rect 13764 24551 13790 24615
rect 13854 24551 13880 24615
rect 13944 24551 13970 24615
rect 14034 24551 14039 24615
rect 13515 24535 14039 24551
rect 13515 24471 13520 24535
rect 13584 24471 13610 24535
rect 13674 24471 13700 24535
rect 13764 24471 13790 24535
rect 13854 24471 13880 24535
rect 13944 24471 13970 24535
rect 14034 24471 14039 24535
rect 13515 24455 14039 24471
rect 13515 24391 13520 24455
rect 13584 24391 13610 24455
rect 13674 24391 13700 24455
rect 13764 24391 13790 24455
rect 13854 24391 13880 24455
rect 13944 24391 13970 24455
rect 14034 24391 14039 24455
rect 13515 24375 14039 24391
rect 13515 24311 13520 24375
rect 13584 24311 13610 24375
rect 13674 24311 13700 24375
rect 13764 24311 13790 24375
rect 13854 24311 13880 24375
rect 13944 24311 13970 24375
rect 14034 24311 14039 24375
rect 13515 24295 14039 24311
rect 13515 24231 13520 24295
rect 13584 24231 13610 24295
rect 13674 24231 13700 24295
rect 13764 24231 13790 24295
rect 13854 24231 13880 24295
rect 13944 24231 13970 24295
rect 14034 24231 14039 24295
rect 13515 24215 14039 24231
rect 13515 24151 13520 24215
rect 13584 24151 13610 24215
rect 13674 24151 13700 24215
rect 13764 24151 13790 24215
rect 13854 24151 13880 24215
rect 13944 24151 13970 24215
rect 14034 24151 14039 24215
rect 13515 24135 14039 24151
rect 13515 24071 13520 24135
rect 13584 24071 13610 24135
rect 13674 24071 13700 24135
rect 13764 24071 13790 24135
rect 13854 24071 13880 24135
rect 13944 24071 13970 24135
rect 14034 24071 14039 24135
rect 13515 24055 14039 24071
rect 13515 23991 13520 24055
rect 13584 23991 13610 24055
rect 13674 23991 13700 24055
rect 13764 23991 13790 24055
rect 13854 23991 13880 24055
rect 13944 23991 13970 24055
rect 14034 23991 14039 24055
rect 13515 23975 14039 23991
rect 13515 23911 13520 23975
rect 13584 23911 13610 23975
rect 13674 23911 13700 23975
rect 13764 23911 13790 23975
rect 13854 23911 13880 23975
rect 13944 23911 13970 23975
rect 14034 23911 14039 23975
rect 13515 23895 14039 23911
rect 13515 23831 13520 23895
rect 13584 23831 13610 23895
rect 13674 23831 13700 23895
rect 13764 23831 13790 23895
rect 13854 23831 13880 23895
rect 13944 23831 13970 23895
rect 14034 23831 14039 23895
rect 13515 23815 14039 23831
rect 13515 23751 13520 23815
rect 13584 23751 13610 23815
rect 13674 23751 13700 23815
rect 13764 23751 13790 23815
rect 13854 23751 13880 23815
rect 13944 23751 13970 23815
rect 14034 23751 14039 23815
rect 13515 23735 14039 23751
rect 13515 23671 13520 23735
rect 13584 23671 13610 23735
rect 13674 23671 13700 23735
rect 13764 23671 13790 23735
rect 13854 23671 13880 23735
rect 13944 23671 13970 23735
rect 14034 23671 14039 23735
rect 13515 23655 14039 23671
rect 13515 23591 13520 23655
rect 13584 23591 13610 23655
rect 13674 23591 13700 23655
rect 13764 23591 13790 23655
rect 13854 23591 13880 23655
rect 13944 23591 13970 23655
rect 14034 23591 14039 23655
rect 13515 23575 14039 23591
rect 13515 23511 13520 23575
rect 13584 23511 13610 23575
rect 13674 23511 13700 23575
rect 13764 23511 13790 23575
rect 13854 23511 13880 23575
rect 13944 23511 13970 23575
rect 14034 23511 14039 23575
rect 13515 23495 14039 23511
rect 13515 23431 13520 23495
rect 13584 23431 13610 23495
rect 13674 23431 13700 23495
rect 13764 23431 13790 23495
rect 13854 23431 13880 23495
rect 13944 23431 13970 23495
rect 14034 23431 14039 23495
rect 13515 23415 14039 23431
rect 13515 23351 13520 23415
rect 13584 23351 13610 23415
rect 13674 23351 13700 23415
rect 13764 23351 13790 23415
rect 13854 23351 13880 23415
rect 13944 23351 13970 23415
rect 14034 23351 14039 23415
rect 13515 23335 14039 23351
rect 13515 23271 13520 23335
rect 13584 23271 13610 23335
rect 13674 23271 13700 23335
rect 13764 23271 13790 23335
rect 13854 23271 13880 23335
rect 13944 23271 13970 23335
rect 14034 23271 14039 23335
rect 13515 23254 14039 23271
rect 13515 23190 13520 23254
rect 13584 23190 13610 23254
rect 13674 23190 13700 23254
rect 13764 23190 13790 23254
rect 13854 23190 13880 23254
rect 13944 23190 13970 23254
rect 14034 23190 14039 23254
rect 13515 23173 14039 23190
rect 13515 23109 13520 23173
rect 13584 23109 13610 23173
rect 13674 23109 13700 23173
rect 13764 23109 13790 23173
rect 13854 23109 13880 23173
rect 13944 23109 13970 23173
rect 14034 23109 14039 23173
rect 13515 23092 14039 23109
rect 13515 23028 13520 23092
rect 13584 23028 13610 23092
rect 13674 23028 13700 23092
rect 13764 23028 13790 23092
rect 13854 23028 13880 23092
rect 13944 23028 13970 23092
rect 14034 23028 14039 23092
rect 13515 23011 14039 23028
rect 13515 22947 13520 23011
rect 13584 22947 13610 23011
rect 13674 22947 13700 23011
rect 13764 22947 13790 23011
rect 13854 22947 13880 23011
rect 13944 22947 13970 23011
rect 14034 22947 14039 23011
rect 13515 22930 14039 22947
rect 13515 22866 13520 22930
rect 13584 22866 13610 22930
rect 13674 22866 13700 22930
rect 13764 22866 13790 22930
rect 13854 22866 13880 22930
rect 13944 22866 13970 22930
rect 14034 22866 14039 22930
rect 13515 22849 14039 22866
rect 13515 22785 13520 22849
rect 13584 22785 13610 22849
rect 13674 22785 13700 22849
rect 13764 22785 13790 22849
rect 13854 22785 13880 22849
rect 13944 22785 13970 22849
rect 14034 22785 14039 22849
rect 13515 22768 14039 22785
rect 13515 22704 13520 22768
rect 13584 22704 13610 22768
rect 13674 22704 13700 22768
rect 13764 22704 13790 22768
rect 13854 22704 13880 22768
rect 13944 22704 13970 22768
rect 14034 22704 14039 22768
rect 13515 22687 14039 22704
rect 13515 22623 13520 22687
rect 13584 22623 13610 22687
rect 13674 22623 13700 22687
rect 13764 22623 13790 22687
rect 13854 22623 13880 22687
rect 13944 22623 13970 22687
rect 14034 22623 14039 22687
rect 13515 22606 14039 22623
rect 13515 22542 13520 22606
rect 13584 22542 13610 22606
rect 13674 22542 13700 22606
rect 13764 22542 13790 22606
rect 13854 22542 13880 22606
rect 13944 22542 13970 22606
rect 14034 22542 14039 22606
rect 13515 22525 14039 22542
rect 13515 22461 13520 22525
rect 13584 22461 13610 22525
rect 13674 22461 13700 22525
rect 13764 22461 13790 22525
rect 13854 22461 13880 22525
rect 13944 22461 13970 22525
rect 14034 22461 14039 22525
rect 13515 22444 14039 22461
rect 13515 22380 13520 22444
rect 13584 22380 13610 22444
rect 13674 22380 13700 22444
rect 13764 22380 13790 22444
rect 13854 22380 13880 22444
rect 13944 22380 13970 22444
rect 14034 22380 14039 22444
rect 13515 22363 14039 22380
rect 13515 22299 13520 22363
rect 13584 22299 13610 22363
rect 13674 22299 13700 22363
rect 13764 22299 13790 22363
rect 13854 22299 13880 22363
rect 13944 22299 13970 22363
rect 14034 22299 14039 22363
rect 13515 22282 14039 22299
rect 13515 22218 13520 22282
rect 13584 22218 13610 22282
rect 13674 22218 13700 22282
rect 13764 22218 13790 22282
rect 13854 22218 13880 22282
rect 13944 22218 13970 22282
rect 14034 22218 14039 22282
rect 13515 22201 14039 22218
rect 13515 22137 13520 22201
rect 13584 22137 13610 22201
rect 13674 22137 13700 22201
rect 13764 22137 13790 22201
rect 13854 22137 13880 22201
rect 13944 22137 13970 22201
rect 14034 22137 14039 22201
rect 13515 22120 14039 22137
rect 13515 22056 13520 22120
rect 13584 22056 13610 22120
rect 13674 22056 13700 22120
rect 13764 22056 13790 22120
rect 13854 22056 13880 22120
rect 13944 22056 13970 22120
rect 14034 22056 14039 22120
rect 13515 22039 14039 22056
rect 13515 21975 13520 22039
rect 13584 21975 13610 22039
rect 13674 21975 13700 22039
rect 13764 21975 13790 22039
rect 13854 21975 13880 22039
rect 13944 21975 13970 22039
rect 14034 21975 14039 22039
rect 13515 21958 14039 21975
rect 13515 21894 13520 21958
rect 13584 21894 13610 21958
rect 13674 21894 13700 21958
rect 13764 21894 13790 21958
rect 13854 21894 13880 21958
rect 13944 21894 13970 21958
rect 14034 21894 14039 21958
rect 13515 21877 14039 21894
rect 13515 21813 13520 21877
rect 13584 21813 13610 21877
rect 13674 21813 13700 21877
rect 13764 21813 13790 21877
rect 13854 21813 13880 21877
rect 13944 21813 13970 21877
rect 14034 21813 14039 21877
rect 13515 21796 14039 21813
rect 13515 21732 13520 21796
rect 13584 21732 13610 21796
rect 13674 21732 13700 21796
rect 13764 21732 13790 21796
rect 13854 21732 13880 21796
rect 13944 21732 13970 21796
rect 14034 21732 14039 21796
rect 13515 21715 14039 21732
rect 13515 21651 13520 21715
rect 13584 21651 13610 21715
rect 13674 21651 13700 21715
rect 13764 21651 13790 21715
rect 13854 21651 13880 21715
rect 13944 21651 13970 21715
rect 14034 21651 14039 21715
rect 13515 21634 14039 21651
rect 13515 21570 13520 21634
rect 13584 21570 13610 21634
rect 13674 21570 13700 21634
rect 13764 21570 13790 21634
rect 13854 21570 13880 21634
rect 13944 21570 13970 21634
rect 14034 21570 14039 21634
rect 13515 21553 14039 21570
rect 13515 21489 13520 21553
rect 13584 21489 13610 21553
rect 13674 21489 13700 21553
rect 13764 21489 13790 21553
rect 13854 21489 13880 21553
rect 13944 21489 13970 21553
rect 14034 21489 14039 21553
rect 13515 21472 14039 21489
rect 13515 21408 13520 21472
rect 13584 21408 13610 21472
rect 13674 21408 13700 21472
rect 13764 21408 13790 21472
rect 13854 21408 13880 21472
rect 13944 21408 13970 21472
rect 14034 21408 14039 21472
rect 13515 21391 14039 21408
rect 13515 21327 13520 21391
rect 13584 21327 13610 21391
rect 13674 21327 13700 21391
rect 13764 21327 13790 21391
rect 13854 21327 13880 21391
rect 13944 21327 13970 21391
rect 14034 21327 14039 21391
rect 13515 21310 14039 21327
rect 13515 21246 13520 21310
rect 13584 21246 13610 21310
rect 13674 21246 13700 21310
rect 13764 21246 13790 21310
rect 13854 21246 13880 21310
rect 13944 21246 13970 21310
rect 14034 21246 14039 21310
rect 13515 21229 14039 21246
rect 13515 21165 13520 21229
rect 13584 21165 13610 21229
rect 13674 21165 13700 21229
rect 13764 21165 13790 21229
rect 13854 21165 13880 21229
rect 13944 21165 13970 21229
rect 14034 21165 14039 21229
rect 13515 21148 14039 21165
rect 13515 21084 13520 21148
rect 13584 21084 13610 21148
rect 13674 21084 13700 21148
rect 13764 21084 13790 21148
rect 13854 21084 13880 21148
rect 13944 21084 13970 21148
rect 14034 21084 14039 21148
rect 13515 21067 14039 21084
rect 13515 21003 13520 21067
rect 13584 21003 13610 21067
rect 13674 21003 13700 21067
rect 13764 21003 13790 21067
rect 13854 21003 13880 21067
rect 13944 21003 13970 21067
rect 14034 21003 14039 21067
rect 13515 20986 14039 21003
rect 13515 20958 13520 20986
rect 1496 20925 1596 20958
rect 1496 20922 1531 20925
rect 977 20905 1531 20922
rect 977 20841 982 20905
rect 1046 20841 1072 20905
rect 1136 20841 1162 20905
rect 1226 20841 1252 20905
rect 1316 20841 1342 20905
rect 1406 20841 1432 20905
rect 1496 20861 1531 20905
rect 1595 20861 1596 20925
rect 1496 20841 1596 20861
rect 977 20840 1596 20841
rect 1471 20828 1596 20840
rect 13420 20925 13520 20958
rect 13420 20861 13421 20925
rect 13485 20922 13520 20925
rect 13584 20922 13610 20986
rect 13674 20922 13700 20986
rect 13764 20922 13790 20986
rect 13854 20922 13880 20986
rect 13944 20922 13970 20986
rect 14034 20922 14039 20986
rect 13485 20905 14039 20922
rect 13485 20861 13520 20905
rect 13420 20841 13520 20861
rect 13584 20841 13610 20905
rect 13674 20841 13700 20905
rect 13764 20841 13790 20905
rect 13854 20841 13880 20905
rect 13944 20841 13970 20905
rect 14034 20841 14039 20905
rect 13420 20840 14039 20841
rect 13420 20828 13545 20840
rect 1311 20811 1736 20813
rect 1140 20769 1265 20802
rect 1140 20705 1141 20769
rect 1205 20705 1265 20769
rect 1140 20672 1265 20705
rect 1311 20747 1312 20811
rect 1376 20747 1401 20811
rect 1465 20747 1491 20811
rect 1555 20747 1581 20811
rect 1645 20747 1671 20811
rect 1735 20747 1736 20811
rect 1311 20695 1736 20747
rect 1311 20631 1312 20695
rect 1376 20631 1401 20695
rect 1465 20631 1491 20695
rect 1555 20631 1581 20695
rect 1645 20631 1671 20695
rect 1735 20631 1736 20695
rect 13280 20811 13705 20813
rect 13280 20747 13281 20811
rect 13345 20747 13371 20811
rect 13435 20747 13461 20811
rect 13525 20747 13551 20811
rect 13615 20747 13640 20811
rect 13704 20747 13705 20811
rect 13280 20695 13705 20747
rect 1311 20579 1736 20631
rect 1311 20515 1312 20579
rect 1376 20515 1401 20579
rect 1465 20515 1491 20579
rect 1555 20515 1581 20579
rect 1645 20515 1671 20579
rect 1735 20515 1736 20579
rect 1752 20617 1877 20650
rect 1752 20553 1812 20617
rect 1876 20553 1877 20617
rect 1752 20520 1877 20553
rect 13139 20617 13264 20650
rect 13139 20553 13140 20617
rect 13204 20553 13264 20617
rect 13139 20520 13264 20553
rect 13280 20631 13281 20695
rect 13345 20631 13371 20695
rect 13435 20631 13461 20695
rect 13525 20631 13551 20695
rect 13615 20631 13640 20695
rect 13704 20631 13705 20695
rect 13719 20809 13843 20810
rect 13719 20745 13749 20809
rect 13813 20745 13843 20809
rect 13719 20698 13843 20745
rect 13849 20802 13916 20835
rect 13849 20738 13851 20802
rect 13915 20738 13916 20802
rect 13849 20705 13916 20738
rect 13719 20634 13749 20698
rect 13813 20634 13843 20698
rect 13719 20633 13843 20634
rect 13280 20579 13705 20631
rect 1311 20513 1736 20515
rect 13280 20515 13281 20579
rect 13345 20515 13371 20579
rect 13435 20515 13461 20579
rect 13525 20515 13551 20579
rect 13615 20515 13640 20579
rect 13704 20515 13705 20579
rect 13280 20513 13705 20515
rect 1631 20491 2056 20493
rect 1464 20455 1589 20488
rect 1464 20391 1524 20455
rect 1588 20391 1589 20455
rect 1464 20358 1589 20391
rect 1631 20427 1632 20491
rect 1696 20427 1721 20491
rect 1785 20427 1811 20491
rect 1875 20427 1901 20491
rect 1965 20427 1991 20491
rect 2055 20427 2056 20491
rect 1631 20375 2056 20427
rect 1631 20311 1632 20375
rect 1696 20311 1721 20375
rect 1785 20311 1811 20375
rect 1875 20311 1901 20375
rect 1965 20311 1991 20375
rect 2055 20311 2056 20375
rect 12960 20491 13385 20493
rect 12960 20427 12961 20491
rect 13025 20427 13051 20491
rect 13115 20427 13141 20491
rect 13205 20427 13231 20491
rect 13295 20427 13320 20491
rect 13384 20427 13385 20491
rect 12960 20375 13385 20427
rect 1631 20259 2056 20311
rect 1631 20195 1632 20259
rect 1696 20195 1721 20259
rect 1785 20195 1811 20259
rect 1875 20195 1901 20259
rect 1965 20195 1991 20259
rect 2055 20195 2056 20259
rect 2077 20292 2202 20325
rect 2077 20228 2137 20292
rect 2201 20228 2202 20292
rect 2077 20195 2202 20228
rect 12814 20292 12939 20325
rect 12814 20228 12815 20292
rect 12879 20228 12939 20292
rect 12814 20195 12939 20228
rect 12960 20311 12961 20375
rect 13025 20311 13051 20375
rect 13115 20311 13141 20375
rect 13205 20311 13231 20375
rect 13295 20311 13320 20375
rect 13384 20311 13385 20375
rect 13427 20455 13552 20488
rect 13427 20391 13428 20455
rect 13492 20391 13552 20455
rect 13427 20358 13552 20391
rect 12960 20259 13385 20311
rect 12960 20195 12961 20259
rect 13025 20195 13051 20259
rect 13115 20195 13141 20259
rect 13205 20195 13231 20259
rect 13295 20195 13320 20259
rect 13384 20195 13385 20259
rect 1631 20193 2056 20195
rect 12960 20193 13385 20195
rect 1955 20167 2380 20169
rect 1792 20127 1917 20160
rect 1792 20063 1852 20127
rect 1916 20063 1917 20127
rect 1792 20030 1917 20063
rect 1955 20103 1956 20167
rect 2020 20103 2045 20167
rect 2109 20103 2135 20167
rect 2199 20103 2225 20167
rect 2289 20103 2315 20167
rect 2379 20103 2380 20167
rect 1955 20051 2380 20103
rect 12636 20167 13061 20169
rect 12636 20103 12637 20167
rect 12701 20103 12727 20167
rect 12791 20103 12817 20167
rect 12881 20103 12907 20167
rect 12971 20103 12996 20167
rect 13060 20103 13061 20167
rect 1955 19987 1956 20051
rect 2020 19987 2045 20051
rect 2109 19987 2135 20051
rect 2199 19987 2225 20051
rect 2289 19987 2315 20051
rect 2379 19987 2380 20051
rect 1955 19935 2380 19987
rect 1955 19871 1956 19935
rect 2020 19871 2045 19935
rect 2109 19871 2135 19935
rect 2199 19871 2225 19935
rect 2289 19871 2315 19935
rect 2379 19871 2380 19935
rect 2455 20056 2867 20057
rect 2455 19992 2456 20056
rect 2520 19992 2571 20056
rect 2635 19992 2686 20056
rect 2750 19992 2802 20056
rect 2866 19992 2867 20056
rect 2455 19936 2867 19992
rect 12149 20056 12561 20057
rect 12149 19992 12150 20056
rect 12214 19992 12266 20056
rect 12330 19992 12381 20056
rect 12445 19992 12496 20056
rect 12560 19992 12561 20056
rect 2455 19872 2456 19936
rect 2520 19872 2571 19936
rect 2635 19872 2686 19936
rect 2750 19872 2802 19936
rect 2866 19872 2867 19936
rect 2455 19871 2867 19872
rect 2881 19941 2971 19974
rect 2881 19877 2906 19941
rect 2970 19877 2971 19941
rect 1955 19869 2380 19871
rect 2881 19844 2971 19877
rect 12045 19941 12135 19974
rect 12045 19877 12046 19941
rect 12110 19877 12135 19941
rect 12045 19844 12135 19877
rect 12149 19936 12561 19992
rect 12149 19872 12150 19936
rect 12214 19872 12266 19936
rect 12330 19872 12381 19936
rect 12445 19872 12496 19936
rect 12560 19872 12561 19936
rect 12149 19871 12561 19872
rect 12636 20051 13061 20103
rect 12636 19987 12637 20051
rect 12701 19987 12727 20051
rect 12791 19987 12817 20051
rect 12881 19987 12907 20051
rect 12971 19987 12996 20051
rect 13060 19987 13061 20051
rect 13099 20127 13224 20160
rect 13099 20063 13100 20127
rect 13164 20063 13224 20127
rect 13099 20030 13224 20063
rect 12636 19935 13061 19987
rect 12636 19871 12637 19935
rect 12701 19871 12727 19935
rect 12791 19871 12817 19935
rect 12881 19871 12907 19935
rect 12971 19871 12996 19935
rect 13060 19871 13061 19935
rect 12636 19869 13061 19871
rect 2292 19830 3114 19832
rect 2133 19786 2258 19819
rect 2133 19722 2193 19786
rect 2257 19722 2258 19786
rect 2133 19689 2258 19722
rect 2292 19766 2293 19830
rect 2357 19766 2377 19830
rect 2441 19766 2461 19830
rect 2525 19766 2545 19830
rect 2609 19766 2629 19830
rect 2693 19766 2713 19830
rect 2777 19766 2797 19830
rect 2861 19766 2881 19830
rect 2945 19766 2965 19830
rect 3029 19766 3049 19830
rect 3113 19766 3114 19830
rect 2292 19714 3114 19766
rect 2292 19650 2293 19714
rect 2357 19650 2377 19714
rect 2441 19650 2461 19714
rect 2525 19650 2545 19714
rect 2609 19650 2629 19714
rect 2693 19650 2713 19714
rect 2777 19650 2797 19714
rect 2861 19650 2881 19714
rect 2945 19650 2965 19714
rect 3029 19650 3049 19714
rect 3113 19650 3114 19714
rect 11902 19830 12724 19832
rect 11902 19766 11903 19830
rect 11967 19766 11987 19830
rect 12051 19766 12071 19830
rect 12135 19766 12155 19830
rect 12219 19766 12239 19830
rect 12303 19766 12323 19830
rect 12387 19766 12407 19830
rect 12471 19766 12491 19830
rect 12555 19766 12575 19830
rect 12639 19766 12659 19830
rect 12723 19766 12724 19830
rect 11902 19714 12724 19766
rect 2292 19598 3114 19650
rect 2292 19534 2293 19598
rect 2357 19534 2377 19598
rect 2441 19534 2461 19598
rect 2525 19534 2545 19598
rect 2609 19534 2629 19598
rect 2693 19534 2713 19598
rect 2777 19534 2797 19598
rect 2861 19534 2881 19598
rect 2945 19534 2965 19598
rect 3029 19534 3049 19598
rect 3113 19534 3114 19598
rect 3123 19693 3247 19694
rect 3123 19629 3153 19693
rect 3217 19629 3247 19693
rect 3123 19600 3247 19629
rect 3123 19536 3153 19600
rect 3217 19536 3247 19600
rect 3123 19535 3247 19536
rect 11769 19693 11893 19694
rect 11769 19629 11799 19693
rect 11863 19629 11893 19693
rect 11769 19600 11893 19629
rect 11769 19536 11799 19600
rect 11863 19536 11893 19600
rect 11769 19535 11893 19536
rect 11902 19650 11903 19714
rect 11967 19650 11987 19714
rect 12051 19650 12071 19714
rect 12135 19650 12155 19714
rect 12219 19650 12239 19714
rect 12303 19650 12323 19714
rect 12387 19650 12407 19714
rect 12471 19650 12491 19714
rect 12555 19650 12575 19714
rect 12639 19650 12659 19714
rect 12723 19650 12724 19714
rect 12758 19786 12883 19819
rect 12758 19722 12759 19786
rect 12823 19722 12883 19786
rect 12758 19689 12883 19722
rect 11902 19598 12724 19650
rect 2292 19532 3114 19534
rect 11902 19534 11903 19598
rect 11967 19534 11987 19598
rect 12051 19534 12071 19598
rect 12135 19534 12155 19598
rect 12219 19534 12239 19598
rect 12303 19534 12323 19598
rect 12387 19534 12407 19598
rect 12471 19534 12491 19598
rect 12555 19534 12575 19598
rect 12639 19534 12659 19598
rect 12723 19534 12724 19598
rect 11902 19532 12724 19534
rect 4912 18895 7268 18934
rect 4912 17311 4938 18895
rect 7242 17311 7268 18895
rect 4912 17273 7268 17311
rect 7712 18895 10068 18934
rect 7712 17311 7738 18895
rect 10042 17311 10068 18895
rect 7712 17273 10068 17311
rect 5077 17218 7265 17231
rect 5077 17074 5099 17218
rect 7243 17074 7265 17218
rect 5077 17061 7265 17074
rect 7713 17218 9901 17231
rect 7713 17074 7735 17218
rect 9879 17074 9901 17218
rect 7713 17061 9901 17074
rect 2423 6025 3607 6053
rect 2423 5213 3607 5241
rect 11297 6024 12481 6052
rect 11297 5212 12481 5240
rect 886 4811 2072 4856
rect 886 4027 887 4811
rect 2071 4027 2072 4811
rect 886 3983 2072 4027
rect 12886 4811 14072 4856
rect 12886 4027 12887 4811
rect 14071 4027 14072 4811
rect 12886 3983 14072 4027
use sky130_ef_io__esd_ndiode_11v0_single  sky130_ef_io__minesd_vddio
timestamp 1701704242
transform 0 1 7496 -1 0 26758
box 160 -5766 1962 5766
use sky130_ef_io__esd_pdiode_11v0_single  sky130_ef_io__minesd_vssio
timestamp 1701704242
transform 0 1 7508 -1 0 29198
box 896 -5188 1566 5188
use sky130_fd_io__com_busses_esd  sky130_fd_io__com_busses_esd_0
timestamp 1701704242
transform 1 0 8 0 1 536
box 0 -142 15000 39451
<< properties >>
string GDS_END 9369002
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io__analog.gds
string GDS_START 7537944
<< end >>
