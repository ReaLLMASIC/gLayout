magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -119 -66 319 266
<< mvpmos >>
rect 0 0 200 200
<< mvpdiff >>
rect -50 0 0 200
rect 200 182 253 200
rect 200 148 211 182
rect 245 148 253 182
rect 200 114 253 148
rect 200 80 211 114
rect 245 80 253 114
rect 200 46 253 80
rect 200 12 211 46
rect 245 12 253 46
rect 200 0 253 12
<< mvpdiffc >>
rect 211 148 245 182
rect 211 80 245 114
rect 211 12 245 46
<< poly >>
rect 0 200 200 226
rect 0 -26 200 0
<< locali >>
rect 211 182 245 198
rect 211 114 245 148
rect 211 46 245 80
rect 211 -4 245 12
<< metal1 >>
rect -51 -16 -5 186
use hvDFL1sd_CDNS_5246887918589  hvDFL1sd_CDNS_5246887918589_0
timestamp 1701704242
transform 1 0 200 0 1 0
box 0 0 1 1
use hvDFM1sd_CDNS_52468879185130  hvDFM1sd_CDNS_52468879185130_0
timestamp 1701704242
transform -1 0 0 0 1 0
box -36 -36 89 236
<< labels >>
flabel comment s -28 85 -28 85 0 FreeSans 300 0 0 0 S
flabel comment s 228 97 228 97 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 85952772
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85951754
<< end >>
