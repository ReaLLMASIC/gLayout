magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -38 261 1602 582
<< pwell >>
rect 1 21 1487 203
rect 31 -17 65 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 247 47 277 177
rect 331 47 361 177
rect 415 47 445 177
rect 499 47 529 177
rect 687 47 717 177
rect 771 47 801 177
rect 855 47 885 177
rect 939 47 969 177
rect 1023 47 1053 177
rect 1107 47 1137 177
rect 1295 47 1325 177
rect 1379 47 1409 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 247 297 277 497
rect 331 297 361 497
rect 415 297 445 497
rect 499 297 529 497
rect 583 297 613 497
rect 668 297 698 497
rect 857 297 887 497
rect 941 297 971 497
rect 1025 297 1055 497
rect 1109 297 1139 497
rect 1277 297 1307 497
rect 1361 297 1391 497
<< ndiff >>
rect 27 95 79 177
rect 27 61 35 95
rect 69 61 79 95
rect 27 47 79 61
rect 109 163 163 177
rect 109 129 119 163
rect 153 129 163 163
rect 109 95 163 129
rect 109 61 119 95
rect 153 61 163 95
rect 109 47 163 61
rect 193 95 247 177
rect 193 61 203 95
rect 237 61 247 95
rect 193 47 247 61
rect 277 163 331 177
rect 277 129 287 163
rect 321 129 331 163
rect 277 95 331 129
rect 277 61 287 95
rect 321 61 331 95
rect 277 47 331 61
rect 361 95 415 177
rect 361 61 371 95
rect 405 61 415 95
rect 361 47 415 61
rect 445 163 499 177
rect 445 129 455 163
rect 489 129 499 163
rect 445 95 499 129
rect 445 61 455 95
rect 489 61 499 95
rect 445 47 499 61
rect 529 163 581 177
rect 529 129 539 163
rect 573 129 581 163
rect 529 47 581 129
rect 635 95 687 177
rect 635 61 643 95
rect 677 61 687 95
rect 635 47 687 61
rect 717 163 771 177
rect 717 129 727 163
rect 761 129 771 163
rect 717 47 771 129
rect 801 163 855 177
rect 801 129 811 163
rect 845 129 855 163
rect 801 95 855 129
rect 801 61 811 95
rect 845 61 855 95
rect 801 47 855 61
rect 885 95 939 177
rect 885 61 895 95
rect 929 61 939 95
rect 885 47 939 61
rect 969 163 1023 177
rect 969 129 979 163
rect 1013 129 1023 163
rect 969 95 1023 129
rect 969 61 979 95
rect 1013 61 1023 95
rect 969 47 1023 61
rect 1053 163 1107 177
rect 1053 129 1063 163
rect 1097 129 1107 163
rect 1053 47 1107 129
rect 1137 93 1189 177
rect 1137 59 1147 93
rect 1181 59 1189 93
rect 1137 47 1189 59
rect 1243 165 1295 177
rect 1243 131 1251 165
rect 1285 131 1295 165
rect 1243 47 1295 131
rect 1325 95 1379 177
rect 1325 61 1335 95
rect 1369 61 1379 95
rect 1325 47 1379 61
rect 1409 163 1461 177
rect 1409 129 1419 163
rect 1453 129 1461 163
rect 1409 95 1461 129
rect 1409 61 1419 95
rect 1453 61 1461 95
rect 1409 47 1461 61
<< pdiff >>
rect 27 477 79 497
rect 27 443 35 477
rect 69 443 79 477
rect 27 409 79 443
rect 27 375 35 409
rect 69 375 79 409
rect 27 297 79 375
rect 109 477 163 497
rect 109 443 119 477
rect 153 443 163 477
rect 109 409 163 443
rect 109 375 119 409
rect 153 375 163 409
rect 109 341 163 375
rect 109 307 119 341
rect 153 307 163 341
rect 109 297 163 307
rect 193 477 247 497
rect 193 443 203 477
rect 237 443 247 477
rect 193 409 247 443
rect 193 375 203 409
rect 237 375 247 409
rect 193 297 247 375
rect 277 477 331 497
rect 277 443 287 477
rect 321 443 331 477
rect 277 409 331 443
rect 277 375 287 409
rect 321 375 331 409
rect 277 341 331 375
rect 277 307 287 341
rect 321 307 331 341
rect 277 297 331 307
rect 361 477 415 497
rect 361 443 371 477
rect 405 443 415 477
rect 361 409 415 443
rect 361 375 371 409
rect 405 375 415 409
rect 361 297 415 375
rect 445 477 499 497
rect 445 443 455 477
rect 489 443 499 477
rect 445 409 499 443
rect 445 375 455 409
rect 489 375 499 409
rect 445 297 499 375
rect 529 477 583 497
rect 529 443 539 477
rect 573 443 583 477
rect 529 297 583 443
rect 613 477 668 497
rect 613 443 624 477
rect 658 443 668 477
rect 613 409 668 443
rect 613 375 624 409
rect 658 375 668 409
rect 613 297 668 375
rect 698 477 750 497
rect 698 443 708 477
rect 742 443 750 477
rect 698 297 750 443
rect 804 477 857 497
rect 804 443 812 477
rect 846 443 857 477
rect 804 297 857 443
rect 887 341 941 497
rect 887 307 897 341
rect 931 307 941 341
rect 887 297 941 307
rect 971 477 1025 497
rect 971 443 981 477
rect 1015 443 1025 477
rect 971 297 1025 443
rect 1055 409 1109 497
rect 1055 375 1065 409
rect 1099 375 1109 409
rect 1055 341 1109 375
rect 1055 307 1065 341
rect 1099 307 1109 341
rect 1055 297 1109 307
rect 1139 477 1277 497
rect 1139 443 1149 477
rect 1183 443 1233 477
rect 1267 443 1277 477
rect 1139 409 1277 443
rect 1139 375 1149 409
rect 1183 375 1233 409
rect 1267 375 1277 409
rect 1139 297 1277 375
rect 1307 409 1361 497
rect 1307 375 1317 409
rect 1351 375 1361 409
rect 1307 341 1361 375
rect 1307 307 1317 341
rect 1351 307 1361 341
rect 1307 297 1361 307
rect 1391 477 1445 497
rect 1391 443 1401 477
rect 1435 443 1445 477
rect 1391 409 1445 443
rect 1391 375 1401 409
rect 1435 375 1445 409
rect 1391 297 1445 375
<< ndiffc >>
rect 35 61 69 95
rect 119 129 153 163
rect 119 61 153 95
rect 203 61 237 95
rect 287 129 321 163
rect 287 61 321 95
rect 371 61 405 95
rect 455 129 489 163
rect 455 61 489 95
rect 539 129 573 163
rect 643 61 677 95
rect 727 129 761 163
rect 811 129 845 163
rect 811 61 845 95
rect 895 61 929 95
rect 979 129 1013 163
rect 979 61 1013 95
rect 1063 129 1097 163
rect 1147 59 1181 93
rect 1251 131 1285 165
rect 1335 61 1369 95
rect 1419 129 1453 163
rect 1419 61 1453 95
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 119 443 153 477
rect 119 375 153 409
rect 119 307 153 341
rect 203 443 237 477
rect 203 375 237 409
rect 287 443 321 477
rect 287 375 321 409
rect 287 307 321 341
rect 371 443 405 477
rect 371 375 405 409
rect 455 443 489 477
rect 455 375 489 409
rect 539 443 573 477
rect 624 443 658 477
rect 624 375 658 409
rect 708 443 742 477
rect 812 443 846 477
rect 897 307 931 341
rect 981 443 1015 477
rect 1065 375 1099 409
rect 1065 307 1099 341
rect 1149 443 1183 477
rect 1233 443 1267 477
rect 1149 375 1183 409
rect 1233 375 1267 409
rect 1317 375 1351 409
rect 1317 307 1351 341
rect 1401 443 1435 477
rect 1401 375 1435 409
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 247 497 277 523
rect 331 497 361 523
rect 415 497 445 523
rect 499 497 529 523
rect 583 497 613 523
rect 668 497 698 523
rect 857 497 887 523
rect 941 497 971 523
rect 1025 497 1055 523
rect 1109 497 1139 523
rect 1277 497 1307 523
rect 1361 497 1391 523
rect 79 265 109 297
rect 163 265 193 297
rect 247 265 277 297
rect 331 265 361 297
rect 415 265 445 297
rect 499 265 529 297
rect 583 265 613 297
rect 668 265 698 297
rect 857 265 887 297
rect 941 265 971 297
rect 79 249 369 265
rect 79 215 115 249
rect 149 215 183 249
rect 217 215 251 249
rect 285 215 319 249
rect 353 215 369 249
rect 79 199 369 215
rect 415 249 529 265
rect 415 215 469 249
rect 503 215 529 249
rect 415 199 529 215
rect 571 249 812 265
rect 857 250 971 265
rect 1025 265 1055 297
rect 1109 265 1139 297
rect 1277 265 1307 297
rect 1361 265 1391 297
rect 1025 251 1207 265
rect 571 215 587 249
rect 621 215 758 249
rect 792 215 812 249
rect 571 199 812 215
rect 855 249 971 250
rect 855 215 889 249
rect 923 231 971 249
rect 1023 249 1207 251
rect 923 215 969 231
rect 855 199 969 215
rect 79 177 109 199
rect 163 177 193 199
rect 247 177 277 199
rect 331 177 361 199
rect 415 177 445 199
rect 499 177 529 199
rect 687 177 717 199
rect 771 177 801 199
rect 855 177 885 199
rect 939 177 969 199
rect 1023 215 1089 249
rect 1123 215 1157 249
rect 1191 215 1207 249
rect 1023 199 1207 215
rect 1268 249 1409 265
rect 1268 215 1284 249
rect 1318 215 1352 249
rect 1386 215 1409 249
rect 1268 199 1409 215
rect 1023 177 1053 199
rect 1107 177 1137 199
rect 1295 177 1325 199
rect 1379 177 1409 199
rect 79 21 109 47
rect 163 21 193 47
rect 247 21 277 47
rect 331 21 361 47
rect 415 21 445 47
rect 499 21 529 47
rect 687 21 717 47
rect 771 21 801 47
rect 855 21 885 47
rect 939 21 969 47
rect 1023 21 1053 47
rect 1107 21 1137 47
rect 1295 21 1325 47
rect 1379 21 1409 47
<< polycont >>
rect 115 215 149 249
rect 183 215 217 249
rect 251 215 285 249
rect 319 215 353 249
rect 469 215 503 249
rect 587 215 621 249
rect 758 215 792 249
rect 889 215 923 249
rect 1089 215 1123 249
rect 1157 215 1191 249
rect 1284 215 1318 249
rect 1352 215 1386 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 31 477 77 527
rect 31 443 35 477
rect 69 443 77 477
rect 31 409 77 443
rect 31 375 35 409
rect 69 375 77 409
rect 31 359 77 375
rect 111 477 161 493
rect 111 443 119 477
rect 153 443 161 477
rect 111 409 161 443
rect 111 375 119 409
rect 153 375 161 409
rect 111 341 161 375
rect 195 477 245 527
rect 195 443 203 477
rect 237 443 245 477
rect 195 409 245 443
rect 195 375 203 409
rect 237 375 245 409
rect 195 359 245 375
rect 279 477 329 493
rect 279 443 287 477
rect 321 443 329 477
rect 279 409 329 443
rect 279 375 287 409
rect 321 375 329 409
rect 111 325 119 341
rect 19 307 119 325
rect 153 325 161 341
rect 279 341 329 375
rect 363 477 413 527
rect 363 443 371 477
rect 405 443 413 477
rect 363 409 413 443
rect 363 375 371 409
rect 405 375 413 409
rect 363 359 413 375
rect 447 477 497 493
rect 447 443 455 477
rect 489 443 497 477
rect 447 409 497 443
rect 531 477 581 527
rect 531 443 539 477
rect 573 443 581 477
rect 531 427 581 443
rect 615 477 666 493
rect 615 443 624 477
rect 658 443 666 477
rect 447 375 455 409
rect 489 393 497 409
rect 615 409 666 443
rect 700 477 750 527
rect 700 443 708 477
rect 742 443 750 477
rect 788 477 1445 493
rect 788 443 812 477
rect 846 443 981 477
rect 1015 443 1149 477
rect 1183 443 1233 477
rect 1267 459 1401 477
rect 1267 443 1277 459
rect 700 427 750 443
rect 1149 409 1277 443
rect 1395 443 1401 459
rect 1435 443 1445 477
rect 615 393 624 409
rect 489 375 624 393
rect 658 393 666 409
rect 812 393 1065 409
rect 658 375 1065 393
rect 1099 375 1115 409
rect 447 359 846 375
rect 1049 341 1115 375
rect 1183 375 1233 409
rect 1267 375 1277 409
rect 1149 359 1277 375
rect 1311 409 1361 425
rect 1311 375 1317 409
rect 1351 375 1361 409
rect 279 325 287 341
rect 153 307 287 325
rect 321 307 329 341
rect 881 325 897 341
rect 19 291 329 307
rect 363 307 897 325
rect 931 325 947 341
rect 931 307 1013 325
rect 363 291 1013 307
rect 1049 307 1065 341
rect 1099 325 1115 341
rect 1311 341 1361 375
rect 1395 409 1445 443
rect 1395 375 1401 409
rect 1435 375 1445 409
rect 1395 357 1445 375
rect 1311 325 1317 341
rect 1099 307 1317 325
rect 1351 307 1361 341
rect 1049 291 1361 307
rect 19 181 65 291
rect 363 257 397 291
rect 99 249 397 257
rect 99 215 115 249
rect 149 215 183 249
rect 217 215 251 249
rect 285 215 319 249
rect 353 223 397 249
rect 453 249 536 257
rect 353 215 369 223
rect 453 215 469 249
rect 503 215 536 249
rect 571 249 812 257
rect 571 215 587 249
rect 621 221 758 249
rect 621 215 638 221
rect 742 215 758 221
rect 792 215 812 249
rect 846 249 945 257
rect 846 215 889 249
rect 923 215 945 249
rect 389 181 399 187
rect 19 163 337 181
rect 19 147 119 163
rect 103 129 119 147
rect 153 145 287 163
rect 153 129 169 145
rect 35 95 69 111
rect 35 17 69 61
rect 103 95 169 129
rect 271 129 287 145
rect 321 129 337 163
rect 371 153 399 181
rect 663 181 680 187
rect 433 163 505 181
rect 433 153 455 163
rect 371 147 455 153
rect 103 61 119 95
rect 153 61 169 95
rect 103 51 169 61
rect 203 95 237 111
rect 203 17 237 61
rect 271 95 337 129
rect 439 129 455 147
rect 489 129 505 163
rect 271 61 287 95
rect 321 61 337 95
rect 271 51 337 61
rect 371 95 405 111
rect 371 17 405 61
rect 439 95 505 129
rect 439 61 455 95
rect 489 61 505 95
rect 439 51 505 61
rect 539 163 573 179
rect 638 153 680 181
rect 714 181 722 187
rect 979 181 1013 291
rect 1047 249 1207 257
rect 1047 215 1089 249
rect 1123 215 1157 249
rect 1191 215 1207 249
rect 1254 249 1456 257
rect 1254 215 1284 249
rect 1318 215 1352 249
rect 1386 215 1456 249
rect 714 163 777 181
rect 714 153 727 163
rect 638 147 727 153
rect 710 129 727 147
rect 761 129 777 163
rect 811 163 1013 181
rect 845 145 979 163
rect 845 129 861 145
rect 539 17 573 129
rect 811 95 861 129
rect 963 129 979 145
rect 1047 165 1469 181
rect 1047 163 1251 165
rect 1047 129 1063 163
rect 1097 131 1251 163
rect 1285 163 1469 165
rect 1285 145 1419 163
rect 1285 131 1301 145
rect 1097 129 1301 131
rect 1403 129 1419 145
rect 1453 129 1469 163
rect 616 61 643 95
rect 677 61 811 95
rect 845 61 861 95
rect 895 95 929 111
rect 895 17 929 61
rect 963 95 1013 129
rect 1335 95 1369 111
rect 963 61 979 95
rect 1013 93 1197 95
rect 1013 61 1147 93
rect 963 59 1147 61
rect 1181 59 1197 93
rect 963 51 1197 59
rect 1335 17 1369 61
rect 1403 95 1469 129
rect 1403 61 1419 95
rect 1453 61 1469 95
rect 1403 51 1469 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 399 153 433 187
rect 680 153 714 187
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
<< metal1 >>
rect 0 561 1564 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 0 496 1564 527
rect 387 187 445 193
rect 387 153 399 187
rect 433 184 445 187
rect 668 187 726 193
rect 668 184 680 187
rect 433 156 680 184
rect 433 153 445 156
rect 387 147 445 153
rect 668 153 680 156
rect 714 153 726 187
rect 668 147 726 153
rect 0 17 1564 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
rect 0 -48 1564 -17
<< labels >>
flabel locali s 583 221 617 255 0 FreeSans 400 0 0 0 A1
port 1 nsew signal input
flabel locali s 1049 221 1083 255 0 FreeSans 400 0 0 0 B1
port 3 nsew signal input
flabel locali s 865 221 899 255 0 FreeSans 400 0 0 0 C1
port 5 nsew signal input
flabel locali s 1316 221 1350 255 0 FreeSans 400 0 0 0 B2
port 4 nsew signal input
flabel locali s 31 221 65 255 0 FreeSans 400 0 0 0 X
port 10 nsew signal output
flabel locali s 491 221 525 255 0 FreeSans 400 0 0 0 A2
port 2 nsew signal input
flabel locali s 31 153 65 187 0 FreeSans 400 0 0 0 X
port 10 nsew signal output
flabel locali s 768 221 802 255 0 FreeSans 400 0 0 0 A1
port 1 nsew signal input
flabel pwell s 31 -17 65 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 31 527 65 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel metal1 s 31 527 65 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional abutment
flabel metal1 s 31 -17 65 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional abutment
rlabel comment s 0 0 0 0 4 a221o_4
rlabel metal1 s 0 -48 1564 48 1 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1564 592 1 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1564 544
string GDS_END 3575720
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3563530
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 39.100 0.000 
<< end >>
