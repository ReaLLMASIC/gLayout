magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< poly >>
rect -50 131 0 160
rect -50 97 -34 131
rect -50 63 0 97
rect -50 29 -34 63
rect -50 0 0 29
rect 300 131 350 160
rect 334 97 350 131
rect 300 63 350 97
rect 334 29 350 63
rect 300 0 350 29
<< polycont >>
rect -34 97 0 131
rect -34 29 0 63
rect 300 97 334 131
rect 300 29 334 63
<< npolyres >>
rect 0 0 300 160
<< locali >>
rect -34 131 0 147
rect -34 63 0 97
rect -34 13 0 29
rect 300 131 334 147
rect 300 63 334 97
rect 300 13 334 29
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_0
timestamp 1701704242
transform -1 0 16 0 1 13
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_1
timestamp 1701704242
transform 1 0 284 0 1 13
box 0 0 1 1
<< properties >>
string GDS_END 90828390
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 90827952
<< end >>
