magic
tech sky130A
timestamp 1701704242
<< pwell >>
rect -13 -13 1108 122
<< psubdiff >>
rect 0 97 1095 109
rect 0 12 12 97
rect 1083 12 1095 97
rect 0 0 1095 12
<< psubdiffcont >>
rect 12 12 1083 97
<< locali >>
rect 12 97 1083 105
rect 12 4 1083 12
<< properties >>
string GDS_END 86371002
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86364662
<< end >>
