magic
tech sky130A
timestamp 1701704242
<< pwell >>
rect -13 -13 564 156
<< psubdiff >>
rect 0 131 551 143
rect 0 12 12 131
rect 539 12 551 131
rect 0 0 551 12
<< psubdiffcont >>
rect 12 12 539 131
<< locali >>
rect 12 131 539 139
rect 12 4 539 12
<< properties >>
string GDS_END 86375352
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86371060
<< end >>
