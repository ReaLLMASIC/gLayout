magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< poly >>
rect -50 67 0 100
rect -50 33 -34 67
rect -50 0 0 33
rect 600 67 650 100
rect 634 33 650 67
rect 600 0 650 33
<< polycont >>
rect -34 33 0 67
rect 600 33 634 67
<< npolyres >>
rect 0 0 600 100
<< locali >>
rect -34 67 0 83
rect -34 17 0 33
rect 600 67 634 83
rect 600 17 634 33
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_0
timestamp 1701704242
transform -1 0 16 0 1 17
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_1
timestamp 1701704242
transform 1 0 584 0 1 17
box 0 0 1 1
<< properties >>
string GDS_END 88438212
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 88437778
<< end >>
