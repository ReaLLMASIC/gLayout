magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< metal2 >>
rect 0 6705 536 6714
rect 0 0 536 9
<< via2 >>
rect 0 9 536 6705
<< metal3 >>
rect -5 6705 541 6710
rect -5 9 0 6705
rect 536 9 541 6705
rect -5 4 541 9
<< properties >>
string GDS_END 93452604
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 93414840
<< end >>
