magic
tech sky130B
timestamp 1701704242
<< viali >>
rect 0 0 53 9341
<< metal1 >>
rect -6 9341 59 9344
rect -6 0 0 9341
rect 53 0 59 9341
rect -6 -3 59 0
<< properties >>
string GDS_END 92165588
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 92132176
<< end >>
