magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -80 2915 290 7977
rect 14636 2915 15006 7977
<< poly >>
rect 249 9450 386 9467
rect 2526 9450 2663 9467
rect 249 9434 452 9450
rect 249 9400 266 9434
rect 300 9400 334 9434
rect 368 9400 402 9434
rect 436 9400 452 9434
rect 249 9384 452 9400
rect 2460 9434 2663 9450
rect 2460 9400 2476 9434
rect 2510 9400 2544 9434
rect 2578 9400 2612 9434
rect 2646 9400 2663 9434
rect 2460 9384 2663 9400
rect 249 9367 386 9384
rect 2526 9367 2663 9384
<< polycont >>
rect 266 9400 300 9434
rect 334 9400 368 9434
rect 402 9400 436 9434
rect 2476 9400 2510 9434
rect 2544 9400 2578 9434
rect 2612 9400 2646 9434
<< locali >>
rect 250 9440 452 9450
rect 250 9434 453 9440
rect 250 9400 263 9434
rect 300 9400 334 9434
rect 369 9400 402 9434
rect 441 9400 453 9434
rect 250 9394 453 9400
rect 2459 9434 2662 9508
rect 2459 9400 2471 9434
rect 2510 9400 2543 9434
rect 2578 9400 2612 9434
rect 2649 9400 2662 9434
rect 2459 9394 2662 9400
rect 250 9384 452 9394
rect 2460 9384 2662 9394
rect 54 2982 224 7910
rect 688 3618 702 7256
rect 14252 3618 14266 7256
rect 14702 2982 14872 7910
<< viali >>
rect 263 9400 266 9434
rect 266 9400 297 9434
rect 335 9400 368 9434
rect 368 9400 369 9434
rect 407 9400 436 9434
rect 436 9400 441 9434
rect 2471 9400 2476 9434
rect 2476 9400 2505 9434
rect 2543 9400 2544 9434
rect 2544 9400 2577 9434
rect 2615 9400 2646 9434
rect 2646 9400 2649 9434
<< metal1 >>
rect 421 9512 473 9520
tri 387 9440 421 9474 se
rect 421 9448 473 9460
rect 250 9434 421 9440
rect 250 9400 263 9434
rect 297 9400 335 9434
rect 369 9400 407 9434
rect 250 9396 421 9400
rect 250 9394 473 9396
tri 417 9390 421 9394 ne
rect 421 9390 473 9394
rect 2459 9434 2662 9487
rect 2459 9400 2471 9434
rect 2505 9400 2543 9434
rect 2577 9400 2615 9434
rect 2649 9400 2662 9434
rect 2459 9357 2662 9400
rect 785 4021 1705 4028
rect 785 3969 791 4021
rect 843 3969 857 4021
rect 909 3969 1705 4021
rect 785 3957 1705 3969
rect 785 3905 791 3957
rect 843 3905 857 3957
rect 909 3905 1705 3957
rect 785 3898 1705 3905
rect 2135 3976 2141 4028
rect 2193 3976 2207 4028
rect 2259 3976 2265 4028
rect 2135 3950 2265 3976
rect 2135 3898 2141 3950
rect 2193 3898 2207 3950
rect 2259 3898 2265 3950
rect 2697 4021 2827 4028
rect 2697 3969 2703 4021
rect 2755 3969 2769 4021
rect 2821 3969 2827 4021
rect 2697 3957 2827 3969
rect 2697 3905 2703 3957
rect 2755 3905 2769 3957
rect 2821 3905 2827 3957
rect 2697 3898 2827 3905
rect 3257 3898 3757 4028
rect 3810 4021 4189 4028
rect 3810 3969 3816 4021
rect 3868 3969 3895 4021
rect 3947 3969 3974 4021
rect 4026 3969 4053 4021
rect 4105 3969 4131 4021
rect 4183 3969 4189 4021
rect 3810 3957 4189 3969
rect 3810 3905 3816 3957
rect 3868 3905 3895 3957
rect 3947 3905 3974 3957
rect 4026 3905 4053 3957
rect 4105 3905 4131 3957
rect 4183 3905 4189 3957
rect 3810 3898 4189 3905
rect 4249 3898 4681 4028
rect 4686 3898 5678 4028
rect 6103 3976 6109 4028
rect 6161 3976 6174 4028
rect 6226 3976 6239 4028
rect 6291 3976 6304 4028
rect 6356 3976 6368 4028
rect 6420 3976 6432 4028
rect 6484 3976 6496 4028
rect 6548 3976 6560 4028
rect 6612 3976 6624 4028
rect 6676 3976 6688 4028
rect 6740 3976 6752 4028
rect 6804 3976 7095 4028
rect 6103 3956 7095 3976
rect 6103 3904 6109 3956
rect 6161 3904 6174 3956
rect 6226 3904 6239 3956
rect 6291 3904 6304 3956
rect 6356 3904 6368 3956
rect 6420 3904 6432 3956
rect 6484 3904 6496 3956
rect 6548 3904 6560 3956
rect 6612 3904 6624 3956
rect 6676 3904 6688 3956
rect 6740 3904 6752 3956
rect 6804 3904 7095 3956
rect 6103 3898 7095 3904
rect 7657 3976 7663 4028
rect 7715 3976 7729 4028
rect 7781 3976 7787 4028
rect 7657 3950 7787 3976
rect 7657 3898 7663 3950
rect 7715 3898 7729 3950
rect 7781 3898 7787 3950
rect 8232 3976 8595 4028
rect 8647 3976 8660 4028
rect 8712 3976 8724 4028
rect 8776 3976 8788 4028
rect 8840 3976 9202 4028
rect 8232 3954 9202 3976
rect 8232 3902 8595 3954
rect 8647 3902 8660 3954
rect 8712 3902 8724 3954
rect 8776 3902 8788 3954
rect 8840 3902 9202 3954
rect 8232 3898 9202 3902
rect 9769 3986 10750 4028
rect 9769 3934 10220 3986
rect 10272 3934 10286 3986
rect 10338 3934 10352 3986
rect 10404 3934 10418 3986
rect 10470 3934 10483 3986
rect 10535 3934 10548 3986
rect 10600 3934 10613 3986
rect 10665 3934 10678 3986
rect 10730 3934 10750 3986
rect 9769 3898 10750 3934
rect 11193 3987 12185 4028
rect 11193 3935 11631 3987
rect 11683 3935 11696 3987
rect 11748 3935 11761 3987
rect 11813 3935 11826 3987
rect 11878 3935 11891 3987
rect 11943 3935 11956 3987
rect 12008 3935 12021 3987
rect 12073 3935 12185 3987
rect 11193 3898 12185 3935
rect 12747 3976 13053 4028
rect 13105 3976 13120 4028
rect 13172 3976 13187 4028
rect 13239 3976 13254 4028
rect 13306 3976 13321 4028
rect 13373 3976 13388 4028
rect 13440 3976 13455 4028
rect 13507 3976 14039 4028
rect 12747 3950 14039 3976
rect 12747 3898 13053 3950
rect 13105 3898 13120 3950
rect 13172 3898 13187 3950
rect 13239 3898 13254 3950
rect 13306 3898 13321 3950
rect 13373 3898 13388 3950
rect 13440 3898 13455 3950
rect 13507 3898 14039 3950
rect 441 2973 641 3074
rect 896 753 904 805
rect 956 753 968 805
rect 1020 753 1266 805
rect 1318 753 1330 805
rect 1382 753 2796 805
rect 2848 753 2860 805
rect 2912 753 5653 805
rect 5705 753 5742 805
rect 5794 753 5831 805
rect 5883 753 5920 805
rect 5972 753 6809 805
rect 6861 753 6873 805
rect 6925 753 8511 805
rect 8563 753 8575 805
rect 8627 753 9991 805
rect 10043 753 10055 805
rect 10107 753 11334 805
rect 11386 753 11398 805
rect 11450 753 12768 805
rect 12820 753 12832 805
rect 12884 753 14701 805
rect 14753 753 14765 805
rect 14817 753 14823 805
rect 300 715 352 721
tri 352 673 358 679 sw
rect 655 673 663 725
rect 715 673 727 725
rect 779 673 1570 725
rect 1622 673 1634 725
rect 1686 673 3100 725
rect 3152 673 3164 725
rect 3216 673 3875 725
rect 3927 673 3939 725
rect 3991 673 4003 725
rect 4055 673 4067 725
rect 4119 673 4131 725
rect 4183 673 7239 725
rect 7291 673 7303 725
rect 7355 673 8941 725
rect 8993 673 9005 725
rect 9057 673 10421 725
rect 10473 673 10485 725
rect 10537 673 11764 725
rect 11816 673 11828 725
rect 11880 673 13198 725
rect 13250 673 13262 725
rect 13314 673 14781 725
rect 14833 673 14845 725
rect 14897 673 14903 725
rect 352 663 358 673
rect 300 651 358 663
rect 352 645 358 651
tri 358 645 386 673 sw
rect 352 599 421 645
rect 300 593 421 599
rect 473 593 485 645
rect 537 593 1853 645
rect 1905 593 1917 645
rect 1969 593 3383 645
rect 3435 593 3447 645
rect 3499 593 7669 645
rect 7721 593 7733 645
rect 7785 593 9371 645
rect 9423 593 9435 645
rect 9487 593 10851 645
rect 10903 593 10915 645
rect 10967 593 12194 645
rect 12246 593 12258 645
rect 12310 593 13628 645
rect 13680 593 13692 645
rect 13744 593 14861 645
rect 14913 593 14925 645
rect 14977 593 14983 645
rect 487 308 573 512
rect 647 307 692 494
rect 773 316 825 525
<< via1 >>
rect 421 9460 473 9512
rect 421 9434 473 9448
rect 421 9400 441 9434
rect 441 9400 473 9434
rect 421 9396 473 9400
rect 791 3969 843 4021
rect 857 3969 909 4021
rect 791 3905 843 3957
rect 857 3905 909 3957
rect 2141 3976 2193 4028
rect 2207 3976 2259 4028
rect 2141 3898 2193 3950
rect 2207 3898 2259 3950
rect 2703 3969 2755 4021
rect 2769 3969 2821 4021
rect 2703 3905 2755 3957
rect 2769 3905 2821 3957
rect 3816 3969 3868 4021
rect 3895 3969 3947 4021
rect 3974 3969 4026 4021
rect 4053 3969 4105 4021
rect 4131 3969 4183 4021
rect 3816 3905 3868 3957
rect 3895 3905 3947 3957
rect 3974 3905 4026 3957
rect 4053 3905 4105 3957
rect 4131 3905 4183 3957
rect 6109 3976 6161 4028
rect 6174 3976 6226 4028
rect 6239 3976 6291 4028
rect 6304 3976 6356 4028
rect 6368 3976 6420 4028
rect 6432 3976 6484 4028
rect 6496 3976 6548 4028
rect 6560 3976 6612 4028
rect 6624 3976 6676 4028
rect 6688 3976 6740 4028
rect 6752 3976 6804 4028
rect 6109 3904 6161 3956
rect 6174 3904 6226 3956
rect 6239 3904 6291 3956
rect 6304 3904 6356 3956
rect 6368 3904 6420 3956
rect 6432 3904 6484 3956
rect 6496 3904 6548 3956
rect 6560 3904 6612 3956
rect 6624 3904 6676 3956
rect 6688 3904 6740 3956
rect 6752 3904 6804 3956
rect 7663 3976 7715 4028
rect 7729 3976 7781 4028
rect 7663 3898 7715 3950
rect 7729 3898 7781 3950
rect 8595 3976 8647 4028
rect 8660 3976 8712 4028
rect 8724 3976 8776 4028
rect 8788 3976 8840 4028
rect 8595 3902 8647 3954
rect 8660 3902 8712 3954
rect 8724 3902 8776 3954
rect 8788 3902 8840 3954
rect 10220 3934 10272 3986
rect 10286 3934 10338 3986
rect 10352 3934 10404 3986
rect 10418 3934 10470 3986
rect 10483 3934 10535 3986
rect 10548 3934 10600 3986
rect 10613 3934 10665 3986
rect 10678 3934 10730 3986
rect 11631 3935 11683 3987
rect 11696 3935 11748 3987
rect 11761 3935 11813 3987
rect 11826 3935 11878 3987
rect 11891 3935 11943 3987
rect 11956 3935 12008 3987
rect 12021 3935 12073 3987
rect 13053 3976 13105 4028
rect 13120 3976 13172 4028
rect 13187 3976 13239 4028
rect 13254 3976 13306 4028
rect 13321 3976 13373 4028
rect 13388 3976 13440 4028
rect 13455 3976 13507 4028
rect 13053 3898 13105 3950
rect 13120 3898 13172 3950
rect 13187 3898 13239 3950
rect 13254 3898 13306 3950
rect 13321 3898 13373 3950
rect 13388 3898 13440 3950
rect 13455 3898 13507 3950
rect 904 753 956 805
rect 968 753 1020 805
rect 1266 753 1318 805
rect 1330 753 1382 805
rect 2796 753 2848 805
rect 2860 753 2912 805
rect 5653 753 5705 805
rect 5742 753 5794 805
rect 5831 753 5883 805
rect 5920 753 5972 805
rect 6809 753 6861 805
rect 6873 753 6925 805
rect 8511 753 8563 805
rect 8575 753 8627 805
rect 9991 753 10043 805
rect 10055 753 10107 805
rect 11334 753 11386 805
rect 11398 753 11450 805
rect 12768 753 12820 805
rect 12832 753 12884 805
rect 14701 753 14753 805
rect 14765 753 14817 805
rect 300 663 352 715
rect 663 673 715 725
rect 727 673 779 725
rect 1570 673 1622 725
rect 1634 673 1686 725
rect 3100 673 3152 725
rect 3164 673 3216 725
rect 3875 673 3927 725
rect 3939 673 3991 725
rect 4003 673 4055 725
rect 4067 673 4119 725
rect 4131 673 4183 725
rect 7239 673 7291 725
rect 7303 673 7355 725
rect 8941 673 8993 725
rect 9005 673 9057 725
rect 10421 673 10473 725
rect 10485 673 10537 725
rect 11764 673 11816 725
rect 11828 673 11880 725
rect 13198 673 13250 725
rect 13262 673 13314 725
rect 14781 673 14833 725
rect 14845 673 14897 725
rect 300 599 352 651
rect 421 593 473 645
rect 485 593 537 645
rect 1853 593 1905 645
rect 1917 593 1969 645
rect 3383 593 3435 645
rect 3447 593 3499 645
rect 7669 593 7721 645
rect 7733 593 7785 645
rect 9371 593 9423 645
rect 9435 593 9487 645
rect 10851 593 10903 645
rect 10915 593 10967 645
rect 12194 593 12246 645
rect 12258 593 12310 645
rect 13628 593 13680 645
rect 13692 593 13744 645
rect 14861 593 14913 645
rect 14925 593 14977 645
<< metal2 >>
rect 321 9512 473 9520
rect 321 9460 421 9512
rect 321 9448 473 9460
rect 321 9396 421 9448
rect 321 9375 473 9396
tri 304 725 321 742 se
rect 321 725 352 9375
tri 352 9254 473 9375 nw
rect 785 4021 915 4028
rect 785 3969 791 4021
rect 843 3969 857 4021
rect 909 3969 915 4021
tri 1750 3976 1802 4028 se
rect 1802 3976 2141 4028
rect 2193 3976 2207 4028
rect 2259 3976 2265 4028
tri 1743 3969 1750 3976 se
rect 1750 3969 2265 3976
rect 785 3957 915 3969
tri 1731 3957 1743 3969 se
rect 1743 3957 2265 3969
rect 785 3905 791 3957
rect 843 3905 857 3957
rect 909 3905 915 3957
tri 1724 3950 1731 3957 se
rect 1731 3950 2265 3957
tri 715 3387 785 3457 se
rect 785 3387 915 3905
tri 1672 3898 1724 3950 se
rect 1724 3898 2141 3950
rect 2193 3898 2207 3950
rect 2259 3898 2265 3950
rect 2697 4021 2827 4028
rect 2697 3969 2703 4021
rect 2755 3969 2769 4021
rect 2821 3969 2827 4021
rect 2697 3957 2827 3969
rect 2697 3905 2703 3957
rect 2755 3905 2769 3957
rect 2821 3905 2827 3957
tri 1618 3844 1672 3898 se
rect 1672 3844 1802 3898
tri 1802 3844 1856 3898 nw
rect 584 3257 915 3387
tri 1497 3723 1618 3844 se
rect 1618 3723 1681 3844
tri 1681 3723 1802 3844 nw
tri 524 1368 584 1428 se
rect 584 1368 714 3257
tri 714 3187 784 3257 nw
tri 1464 1422 1497 1455 se
rect 1497 1422 1627 3723
tri 1627 3669 1681 3723 nw
rect 2697 3319 2827 3905
rect 3810 4021 4189 4028
rect 3810 3969 3816 4021
rect 3868 3969 3895 4021
rect 3947 3969 3974 4021
rect 4026 3969 4053 4021
rect 4105 3969 4131 4021
rect 4183 3969 4189 4021
rect 3810 3957 4189 3969
rect 3810 3905 3816 3957
rect 3868 3905 3895 3957
rect 3947 3905 3974 3957
rect 4026 3905 4053 3957
rect 4105 3905 4131 3957
rect 4183 3905 4189 3957
tri 2827 3319 2852 3344 sw
rect 2697 3290 2852 3319
tri 2697 3135 2852 3290 ne
tri 2852 3135 3036 3319 sw
tri 2852 2951 3036 3135 ne
tri 3036 2951 3220 3135 sw
tri 3036 2897 3090 2951 ne
tri 714 1368 768 1422 sw
tri 1410 1368 1464 1422 se
rect 1464 1368 1627 1422
tri 1627 1368 1714 1455 sw
tri 3003 1368 3090 1455 se
rect 3090 1368 3220 2951
tri 3220 1368 3307 1455 sw
tri 300 721 304 725 se
rect 304 721 352 725
rect 300 715 352 721
rect 300 651 352 663
rect 300 593 352 599
rect 413 1254 1026 1368
rect 413 1202 543 1254
tri 543 1220 577 1254 nw
tri 621 1220 655 1254 ne
rect 414 1200 542 1201
rect 655 1202 785 1254
tri 785 1220 819 1254 nw
tri 862 1220 896 1254 ne
rect 656 1200 784 1201
rect 896 1202 1026 1254
rect 897 1200 1025 1201
rect 1260 1254 1977 1368
rect 1260 1202 1390 1254
tri 1390 1218 1426 1254 nw
tri 1528 1218 1564 1254 ne
rect 1261 1200 1389 1201
rect 1564 1202 1694 1254
tri 1694 1218 1730 1254 nw
tri 1811 1218 1847 1254 ne
rect 1565 1200 1693 1201
rect 1847 1202 1977 1254
rect 1848 1200 1976 1201
rect 2790 1254 3507 1368
rect 2790 1202 2920 1254
tri 2920 1218 2956 1254 nw
tri 3058 1218 3094 1254 ne
rect 2791 1200 2919 1201
rect 3094 1202 3224 1254
tri 3224 1218 3260 1254 nw
tri 3341 1218 3377 1254 ne
rect 3095 1200 3223 1201
rect 3377 1202 3507 1254
rect 3378 1200 3506 1201
rect 413 900 543 1200
rect 1260 900 1390 1200
rect 2790 900 2920 1200
rect 414 899 542 900
rect 413 645 543 898
rect 656 899 784 900
rect 655 725 785 898
rect 897 899 1025 900
rect 896 805 1026 898
rect 896 753 904 805
rect 956 753 968 805
rect 1020 753 1026 805
rect 1261 899 1389 900
rect 1260 805 1390 898
rect 1260 753 1266 805
rect 1318 753 1330 805
rect 1382 753 1390 805
rect 1565 899 1693 900
rect 655 673 663 725
rect 715 673 727 725
rect 779 673 785 725
rect 1564 725 1694 898
rect 1564 673 1570 725
rect 1622 673 1634 725
rect 1686 673 1694 725
rect 1848 899 1976 900
rect 413 593 421 645
rect 473 593 485 645
rect 537 593 543 645
rect 1847 645 1977 898
rect 2791 899 2919 900
rect 2790 805 2920 898
rect 2790 753 2796 805
rect 2848 753 2860 805
rect 2912 753 2920 805
rect 3095 899 3223 900
rect 3094 725 3224 898
rect 3094 673 3100 725
rect 3152 673 3164 725
rect 3216 673 3224 725
rect 3378 899 3506 900
rect 1847 593 1853 645
rect 1905 593 1917 645
rect 1969 593 1977 645
rect 3377 645 3507 898
rect 3810 725 4189 3905
rect 5647 3976 6109 4028
rect 6161 3976 6174 4028
rect 6226 3976 6239 4028
rect 6291 3976 6304 4028
rect 6356 3976 6368 4028
rect 6420 3976 6432 4028
rect 6484 3976 6496 4028
rect 6548 3976 6560 4028
rect 6612 3976 6624 4028
rect 6676 3976 6688 4028
rect 6740 3976 6752 4028
rect 6804 3976 6810 4028
rect 5647 3956 6810 3976
rect 5647 3904 6109 3956
rect 6161 3904 6174 3956
rect 6226 3904 6239 3956
rect 6291 3904 6304 3956
rect 6356 3904 6368 3956
rect 6420 3904 6432 3956
rect 6484 3904 6496 3956
rect 6548 3904 6560 3956
rect 6612 3904 6624 3956
rect 6676 3904 6688 3956
rect 6740 3904 6752 3956
rect 6804 3904 6810 3956
rect 7657 3976 7663 4028
rect 7715 3976 7729 4028
rect 7781 3976 7787 4028
rect 7657 3950 7787 3976
rect 5647 3903 6112 3904
tri 6112 3903 6113 3904 nw
rect 5647 3899 6108 3903
tri 6108 3899 6112 3903 nw
rect 5647 3898 6107 3899
tri 6107 3898 6108 3899 nw
rect 7657 3898 7663 3950
rect 7715 3898 7729 3950
rect 7781 3898 7787 3950
rect 5647 805 5978 3898
tri 5978 3769 6107 3898 nw
tri 7477 1500 7657 1680 se
rect 7657 1500 7787 3898
tri 7463 1486 7477 1500 se
rect 7477 1486 7787 1500
rect 8589 3976 8595 4028
rect 8647 3976 8660 4028
rect 8712 3976 8724 4028
rect 8776 3976 8788 4028
rect 8840 3976 8846 4028
rect 8589 3954 8846 3976
rect 8589 3902 8595 3954
rect 8647 3902 8660 3954
rect 8712 3902 8724 3954
rect 8776 3902 8788 3954
rect 8840 3902 8846 3954
tri 7457 1480 7463 1486 se
rect 7463 1480 7787 1486
tri 7787 1480 7793 1486 sw
tri 7345 1368 7457 1480 se
rect 7457 1368 7793 1480
rect 6803 1254 7793 1368
rect 6803 1202 6933 1254
tri 6933 1218 6969 1254 nw
tri 7197 1218 7233 1254 ne
rect 6804 1200 6932 1201
rect 7233 1202 7363 1254
tri 7363 1218 7399 1254 nw
tri 7627 1218 7663 1254 ne
rect 7234 1200 7362 1201
rect 7663 1202 7793 1254
rect 7664 1200 7792 1201
tri 8505 1328 8589 1412 se
rect 8589 1368 8846 3902
rect 10214 3986 10736 4017
rect 10214 3934 10220 3986
rect 10272 3934 10286 3986
rect 10338 3934 10352 3986
rect 10404 3934 10418 3986
rect 10470 3934 10483 3986
rect 10535 3934 10548 3986
rect 10600 3934 10613 3986
rect 10665 3934 10678 3986
rect 10730 3934 10736 3986
tri 10132 1418 10214 1500 se
rect 10214 1418 10736 3934
rect 11625 3987 12079 4018
rect 11625 3935 11631 3987
rect 11683 3935 11696 3987
rect 11748 3935 11761 3987
rect 11813 3935 11826 3987
rect 11878 3935 11891 3987
rect 11943 3935 11956 3987
rect 12008 3935 12021 3987
rect 12073 3935 12079 3987
tri 11587 1530 11625 1568 se
rect 11625 1530 12079 3935
rect 13047 3976 13053 4028
rect 13105 3976 13120 4028
rect 13172 3976 13187 4028
rect 13239 3976 13254 4028
rect 13306 3976 13321 4028
rect 13373 3976 13388 4028
rect 13440 3976 13455 4028
rect 13507 3976 13513 4028
rect 13047 3950 13513 3976
rect 13047 3898 13053 3950
rect 13105 3898 13120 3950
rect 13172 3898 13187 3950
rect 13239 3898 13254 3950
rect 13306 3898 13321 3950
rect 13373 3898 13388 3950
rect 13440 3898 13455 3950
rect 13507 3898 13513 3950
tri 11557 1500 11587 1530 se
rect 11587 1500 12079 1530
tri 13017 1500 13047 1530 se
rect 13047 1500 13513 3898
tri 8846 1368 8896 1418 sw
tri 10082 1368 10132 1418 se
rect 10132 1368 10736 1418
tri 10736 1368 10868 1500 sw
tri 11425 1368 11557 1500 se
rect 11557 1474 12079 1500
tri 12079 1474 12105 1500 sw
tri 12991 1474 13017 1500 se
rect 13017 1474 13513 1500
rect 11557 1368 12105 1474
tri 12105 1368 12211 1474 sw
tri 12885 1368 12991 1474 se
rect 12991 1368 13513 1474
tri 13513 1368 13619 1474 sw
rect 8589 1328 8896 1368
tri 8896 1328 8936 1368 sw
rect 8505 1254 9495 1328
rect 8505 1202 8635 1254
tri 8635 1218 8671 1254 nw
tri 8899 1218 8935 1254 ne
rect 8506 1200 8634 1201
rect 8935 1202 9065 1254
tri 9065 1218 9101 1254 nw
tri 9329 1218 9365 1254 ne
rect 8936 1200 9064 1201
rect 9365 1202 9495 1254
rect 9366 1200 9494 1201
rect 9985 1254 10975 1368
rect 9985 1202 10115 1254
tri 10115 1218 10151 1254 nw
tri 10379 1218 10415 1254 ne
rect 9986 1200 10114 1201
rect 10415 1202 10545 1254
tri 10545 1218 10581 1254 nw
tri 10809 1218 10845 1254 ne
rect 10416 1200 10544 1201
rect 10845 1202 10975 1254
rect 10846 1200 10974 1201
rect 11328 1254 12318 1368
rect 11328 1202 11458 1254
tri 11458 1218 11494 1254 nw
tri 11722 1218 11758 1254 ne
rect 11329 1200 11457 1201
rect 11758 1202 11888 1254
tri 11888 1218 11924 1254 nw
tri 12152 1218 12188 1254 ne
rect 11759 1200 11887 1201
rect 12188 1202 12318 1254
rect 12189 1200 12317 1201
rect 12762 1254 13752 1368
rect 12762 1202 12892 1254
tri 12892 1218 12928 1254 nw
tri 13156 1218 13192 1254 ne
rect 12763 1200 12891 1201
rect 13192 1202 13322 1254
tri 13322 1218 13358 1254 nw
tri 13586 1218 13622 1254 ne
rect 13193 1200 13321 1201
rect 13622 1202 13752 1254
rect 13623 1200 13751 1201
rect 7233 900 7363 1200
rect 8935 900 9065 1200
rect 10415 900 10545 1200
rect 11758 900 11888 1200
rect 13622 900 13752 1200
rect 5647 753 5653 805
rect 5705 753 5742 805
rect 5794 753 5831 805
rect 5883 753 5920 805
rect 5972 753 5978 805
rect 6804 899 6932 900
rect 6803 805 6933 898
rect 6803 753 6809 805
rect 6861 753 6873 805
rect 6925 753 6933 805
rect 7234 899 7362 900
rect 3810 673 3875 725
rect 3927 673 3939 725
rect 3991 673 4003 725
rect 4055 673 4067 725
rect 4119 673 4131 725
rect 4183 673 4189 725
rect 7233 725 7363 898
rect 7233 673 7239 725
rect 7291 673 7303 725
rect 7355 673 7363 725
rect 7664 899 7792 900
rect 3377 593 3383 645
rect 3435 593 3447 645
rect 3499 593 3507 645
rect 7663 645 7793 898
rect 8506 899 8634 900
rect 8505 805 8635 898
rect 8505 753 8511 805
rect 8563 753 8575 805
rect 8627 753 8635 805
rect 8936 899 9064 900
rect 8935 725 9065 898
rect 8935 673 8941 725
rect 8993 673 9005 725
rect 9057 673 9065 725
rect 9366 899 9494 900
rect 7663 593 7669 645
rect 7721 593 7733 645
rect 7785 593 7793 645
rect 9365 645 9495 898
rect 9986 899 10114 900
rect 9985 805 10115 898
rect 9985 753 9991 805
rect 10043 753 10055 805
rect 10107 753 10115 805
rect 10416 899 10544 900
rect 10415 725 10545 898
rect 10415 673 10421 725
rect 10473 673 10485 725
rect 10537 673 10545 725
rect 10846 899 10974 900
rect 9365 593 9371 645
rect 9423 593 9435 645
rect 9487 593 9495 645
rect 10845 645 10975 898
rect 11329 899 11457 900
rect 11328 805 11458 898
rect 11328 753 11334 805
rect 11386 753 11398 805
rect 11450 753 11458 805
rect 11759 899 11887 900
rect 11758 725 11888 898
rect 11758 673 11764 725
rect 11816 673 11828 725
rect 11880 673 11888 725
rect 12189 899 12317 900
rect 10845 593 10851 645
rect 10903 593 10915 645
rect 10967 593 10975 645
rect 12188 645 12318 898
rect 12763 899 12891 900
rect 12762 805 12892 898
rect 12762 753 12768 805
rect 12820 753 12832 805
rect 12884 753 12892 805
rect 13193 899 13321 900
rect 13192 725 13322 898
rect 13192 673 13198 725
rect 13250 673 13262 725
rect 13314 673 13322 725
rect 13623 899 13751 900
rect 12188 593 12194 645
rect 12246 593 12258 645
rect 12310 593 12318 645
rect 13622 645 13752 898
tri 14755 805 14783 833 se
rect 14695 753 14701 805
rect 14753 753 14765 805
rect 14817 753 14823 805
tri 14835 725 14863 753 se
rect 14775 673 14781 725
rect 14833 673 14845 725
rect 14897 673 14903 725
tri 14915 645 14943 673 se
rect 13622 593 13628 645
rect 13680 593 13692 645
rect 13744 593 13752 645
rect 14855 593 14861 645
rect 14913 593 14925 645
rect 14977 593 14983 645
<< rmetal2 >>
rect 413 1201 543 1202
rect 413 1200 414 1201
rect 542 1200 543 1201
rect 655 1201 785 1202
rect 655 1200 656 1201
rect 784 1200 785 1201
rect 896 1201 1026 1202
rect 896 1200 897 1201
rect 1025 1200 1026 1201
rect 1260 1201 1390 1202
rect 1260 1200 1261 1201
rect 1389 1200 1390 1201
rect 1564 1201 1694 1202
rect 1564 1200 1565 1201
rect 1693 1200 1694 1201
rect 1847 1201 1977 1202
rect 1847 1200 1848 1201
rect 1976 1200 1977 1201
rect 2790 1201 2920 1202
rect 2790 1200 2791 1201
rect 2919 1200 2920 1201
rect 3094 1201 3224 1202
rect 3094 1200 3095 1201
rect 3223 1200 3224 1201
rect 3377 1201 3507 1202
rect 3377 1200 3378 1201
rect 3506 1200 3507 1201
rect 413 899 414 900
rect 542 899 543 900
rect 413 898 543 899
rect 655 899 656 900
rect 784 899 785 900
rect 655 898 785 899
rect 896 899 897 900
rect 1025 899 1026 900
rect 896 898 1026 899
rect 1260 899 1261 900
rect 1389 899 1390 900
rect 1260 898 1390 899
rect 1564 899 1565 900
rect 1693 899 1694 900
rect 1564 898 1694 899
rect 1847 899 1848 900
rect 1976 899 1977 900
rect 1847 898 1977 899
rect 2790 899 2791 900
rect 2919 899 2920 900
rect 2790 898 2920 899
rect 3094 899 3095 900
rect 3223 899 3224 900
rect 3094 898 3224 899
rect 3377 899 3378 900
rect 3506 899 3507 900
rect 3377 898 3507 899
rect 6803 1201 6933 1202
rect 6803 1200 6804 1201
rect 6932 1200 6933 1201
rect 7233 1201 7363 1202
rect 7233 1200 7234 1201
rect 7362 1200 7363 1201
rect 7663 1201 7793 1202
rect 7663 1200 7664 1201
rect 7792 1200 7793 1201
rect 8505 1201 8635 1202
rect 8505 1200 8506 1201
rect 8634 1200 8635 1201
rect 8935 1201 9065 1202
rect 8935 1200 8936 1201
rect 9064 1200 9065 1201
rect 9365 1201 9495 1202
rect 9365 1200 9366 1201
rect 9494 1200 9495 1201
rect 9985 1201 10115 1202
rect 9985 1200 9986 1201
rect 10114 1200 10115 1201
rect 10415 1201 10545 1202
rect 10415 1200 10416 1201
rect 10544 1200 10545 1201
rect 10845 1201 10975 1202
rect 10845 1200 10846 1201
rect 10974 1200 10975 1201
rect 11328 1201 11458 1202
rect 11328 1200 11329 1201
rect 11457 1200 11458 1201
rect 11758 1201 11888 1202
rect 11758 1200 11759 1201
rect 11887 1200 11888 1201
rect 12188 1201 12318 1202
rect 12188 1200 12189 1201
rect 12317 1200 12318 1201
rect 12762 1201 12892 1202
rect 12762 1200 12763 1201
rect 12891 1200 12892 1201
rect 13192 1201 13322 1202
rect 13192 1200 13193 1201
rect 13321 1200 13322 1201
rect 13622 1201 13752 1202
rect 13622 1200 13623 1201
rect 13751 1200 13752 1201
rect 6803 899 6804 900
rect 6932 899 6933 900
rect 6803 898 6933 899
rect 7233 899 7234 900
rect 7362 899 7363 900
rect 7233 898 7363 899
rect 7663 899 7664 900
rect 7792 899 7793 900
rect 7663 898 7793 899
rect 8505 899 8506 900
rect 8634 899 8635 900
rect 8505 898 8635 899
rect 8935 899 8936 900
rect 9064 899 9065 900
rect 8935 898 9065 899
rect 9365 899 9366 900
rect 9494 899 9495 900
rect 9365 898 9495 899
rect 9985 899 9986 900
rect 10114 899 10115 900
rect 9985 898 10115 899
rect 10415 899 10416 900
rect 10544 899 10545 900
rect 10415 898 10545 899
rect 10845 899 10846 900
rect 10974 899 10975 900
rect 10845 898 10975 899
rect 11328 899 11329 900
rect 11457 899 11458 900
rect 11328 898 11458 899
rect 11758 899 11759 900
rect 11887 899 11888 900
rect 11758 898 11888 899
rect 12188 899 12189 900
rect 12317 899 12318 900
rect 12188 898 12318 899
rect 12762 899 12763 900
rect 12891 899 12892 900
rect 12762 898 12892 899
rect 13192 899 13193 900
rect 13321 899 13322 900
rect 13192 898 13322 899
rect 13622 899 13623 900
rect 13751 899 13752 900
rect 13622 898 13752 899
use PYL1_C_CDNS_524688791850  PYL1_C_CDNS_524688791850_0
timestamp 1701704242
transform -1 0 2561 0 -1 9417
box 0 0 1 1
use PYL1_C_CDNS_524688791850  PYL1_C_CDNS_524688791850_1
timestamp 1701704242
transform 1 0 351 0 -1 9417
box 0 0 1 1
use PYres_CDNS_524688791856  PYres_CDNS_524688791856_0
timestamp 1701704242
transform 1 0 436 0 1 9367
box -50 0 2090 100
use sky130_fd_io__NFET_con_diff_wo_abt_270_analog_pad  sky130_fd_io__NFET_con_diff_wo_abt_270_analog_pad_0
timestamp 1701704242
transform -1 0 15088 0 -1 8404
box 8 427 15168 5489
use sky130_fd_io__tk_em2o_CDNS_524688791854  sky130_fd_io__tk_em2o_CDNS_524688791854_0
timestamp 1701704242
transform 0 1 896 1 0 846
box 0 0 1 1
use sky130_fd_io__tk_em2o_CDNS_524688791854  sky130_fd_io__tk_em2o_CDNS_524688791854_1
timestamp 1701704242
transform 0 1 655 1 0 846
box 0 0 1 1
use sky130_fd_io__tk_em2o_CDNS_524688791854  sky130_fd_io__tk_em2o_CDNS_524688791854_2
timestamp 1701704242
transform 0 -1 1694 1 0 846
box 0 0 1 1
use sky130_fd_io__tk_em2o_CDNS_524688791854  sky130_fd_io__tk_em2o_CDNS_524688791854_3
timestamp 1701704242
transform 0 -1 1977 1 0 846
box 0 0 1 1
use sky130_fd_io__tk_em2o_CDNS_524688791854  sky130_fd_io__tk_em2o_CDNS_524688791854_4
timestamp 1701704242
transform 0 -1 3507 1 0 846
box 0 0 1 1
use sky130_fd_io__tk_em2o_CDNS_524688791854  sky130_fd_io__tk_em2o_CDNS_524688791854_5
timestamp 1701704242
transform 0 -1 7793 1 0 846
box 0 0 1 1
use sky130_fd_io__tk_em2o_CDNS_524688791854  sky130_fd_io__tk_em2o_CDNS_524688791854_6
timestamp 1701704242
transform 0 -1 12318 1 0 846
box 0 0 1 1
use sky130_fd_io__tk_em2o_CDNS_524688791854  sky130_fd_io__tk_em2o_CDNS_524688791854_7
timestamp 1701704242
transform 0 -1 9495 1 0 846
box 0 0 1 1
use sky130_fd_io__tk_em2o_CDNS_524688791854  sky130_fd_io__tk_em2o_CDNS_524688791854_8
timestamp 1701704242
transform 0 -1 10975 1 0 846
box 0 0 1 1
use sky130_fd_io__tk_em2o_CDNS_524688791854  sky130_fd_io__tk_em2o_CDNS_524688791854_9
timestamp 1701704242
transform 0 -1 3224 1 0 846
box 0 0 1 1
use sky130_fd_io__tk_em2o_CDNS_524688791854  sky130_fd_io__tk_em2o_CDNS_524688791854_10
timestamp 1701704242
transform 0 -1 13322 1 0 846
box 0 0 1 1
use sky130_fd_io__tk_em2o_CDNS_524688791854  sky130_fd_io__tk_em2o_CDNS_524688791854_11
timestamp 1701704242
transform 0 -1 6933 1 0 846
box 0 0 1 1
use sky130_fd_io__tk_em2o_CDNS_524688791854  sky130_fd_io__tk_em2o_CDNS_524688791854_12
timestamp 1701704242
transform 0 -1 8635 1 0 846
box 0 0 1 1
use sky130_fd_io__tk_em2o_CDNS_524688791854  sky130_fd_io__tk_em2o_CDNS_524688791854_13
timestamp 1701704242
transform 0 -1 10115 1 0 846
box 0 0 1 1
use sky130_fd_io__tk_em2o_CDNS_524688791854  sky130_fd_io__tk_em2o_CDNS_524688791854_14
timestamp 1701704242
transform 0 -1 11458 1 0 846
box 0 0 1 1
use sky130_fd_io__tk_em2o_CDNS_524688791854  sky130_fd_io__tk_em2o_CDNS_524688791854_15
timestamp 1701704242
transform 0 -1 12892 1 0 846
box 0 0 1 1
use sky130_fd_io__tk_em2s_CDNS_524688791855  sky130_fd_io__tk_em2s_CDNS_524688791855_0
timestamp 1701704242
transform 0 1 413 1 0 846
box 0 0 1 1
use sky130_fd_io__tk_em2s_CDNS_524688791855  sky130_fd_io__tk_em2s_CDNS_524688791855_1
timestamp 1701704242
transform 0 -1 1390 1 0 846
box 0 0 1 1
use sky130_fd_io__tk_em2s_CDNS_524688791855  sky130_fd_io__tk_em2s_CDNS_524688791855_2
timestamp 1701704242
transform 0 -1 13752 1 0 846
box 0 0 1 1
use sky130_fd_io__tk_em2s_CDNS_524688791855  sky130_fd_io__tk_em2s_CDNS_524688791855_3
timestamp 1701704242
transform 0 -1 9065 1 0 846
box 0 0 1 1
use sky130_fd_io__tk_em2s_CDNS_524688791855  sky130_fd_io__tk_em2s_CDNS_524688791855_4
timestamp 1701704242
transform 0 -1 10545 1 0 846
box 0 0 1 1
use sky130_fd_io__tk_em2s_CDNS_524688791855  sky130_fd_io__tk_em2s_CDNS_524688791855_5
timestamp 1701704242
transform 0 -1 7363 1 0 846
box 0 0 1 1
use sky130_fd_io__tk_em2s_CDNS_524688791855  sky130_fd_io__tk_em2s_CDNS_524688791855_6
timestamp 1701704242
transform 0 -1 11888 1 0 846
box 0 0 1 1
use sky130_fd_io__tk_em2s_CDNS_524688791855  sky130_fd_io__tk_em2s_CDNS_524688791855_7
timestamp 1701704242
transform 0 -1 2920 1 0 846
box 0 0 1 1
<< labels >>
flabel comment s 531 416 531 416 0 FreeSans 200 270 0 0 m1_float
flabel comment s 673 407 673 407 0 FreeSans 200 270 0 0 m1_float
flabel comment s 808 407 808 407 0 FreeSans 200 270 0 0 m1_float
flabel comment s 2310 1270 2310 1270 0 FreeSans 440 0 0 0 res
flabel comment s 1561 9429 1561 9429 0 FreeSans 440 0 0 0 leaker
flabel comment s 1276 7506 1276 7506 0 FreeSans 440 180 0 0 condiode
flabel metal1 s 490 308 570 370 3 FreeSans 520 90 0 0 force_lo_h
port 3 nsew
flabel metal1 s 653 310 687 352 3 FreeSans 520 90 0 0 force_lovol_h
port 6 nsew
flabel metal1 s 779 316 819 388 3 FreeSans 520 90 0 0 vssio_amx
port 7 nsew
flabel metal1 s 2527 9424 2599 9476 0 FreeSans 400 180 0 0 vgnd_io
port 1 nsew
flabel metal1 s 301 9395 392 9439 0 FreeSans 400 0 0 0 tie_lo_esd
port 2 nsew
flabel metal1 s 14833 593 14937 645 0 FreeSans 400 0 0 0 tie_lo_esd
port 2 nsew
flabel metal1 s 14701 673 14857 725 0 FreeSans 400 0 0 0 pd_h<3>
port 4 nsew
flabel metal1 s 14692 753 14777 805 0 FreeSans 400 0 0 0 pd_h<2>
port 5 nsew
flabel metal1 s 441 2973 641 3074 0 FreeSans 400 0 0 0 vcc_io
port 8 nsew
<< properties >>
string GDS_END 14492172
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 14466518
string path 13.575 15.475 10.325 15.475 
<< end >>
