magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -122 -66 498 1066
<< mvpmos >>
rect 0 0 160 1000
rect 216 0 376 1000
<< mvpdiff >>
rect -50 0 0 1000
rect 376 0 426 1000
<< poly >>
rect 0 1000 160 1032
rect 0 -32 160 0
rect 216 1000 376 1032
rect 216 -32 376 0
<< locali >>
rect -45 -4 -11 946
rect 171 -4 205 946
rect 387 -4 421 946
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_0
timestamp 1701704242
transform -1 0 0 0 1 0
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_1
timestamp 1701704242
transform 1 0 376 0 1 0
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_2
timestamp 1701704242
transform 1 0 160 0 1 0
box -36 -36 92 1036
<< labels >>
flabel comment s -28 471 -28 471 0 FreeSans 300 0 0 0 S
flabel comment s 188 471 188 471 0 FreeSans 300 0 0 0 D
flabel comment s 404 471 404 471 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 85605066
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85603550
<< end >>
