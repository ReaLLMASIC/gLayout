magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -119 -66 1119 266
<< mvpmos >>
rect 0 0 120 200
rect 176 0 296 200
rect 352 0 472 200
rect 528 0 648 200
rect 704 0 824 200
rect 880 0 1000 200
<< mvpdiff >>
rect -50 0 0 200
rect 1000 0 1050 200
<< poly >>
rect 0 200 120 226
rect 0 -26 120 0
rect 176 200 296 226
rect 176 -26 296 0
rect 352 200 472 226
rect 352 -26 472 0
rect 528 200 648 226
rect 528 -26 648 0
rect 704 200 824 226
rect 704 -26 824 0
rect 880 200 1000 226
rect 880 -26 1000 0
<< metal1 >>
rect -51 -16 -5 186
rect 125 -16 171 186
rect 301 -16 347 186
rect 477 -16 523 186
rect 653 -16 699 186
rect 829 -16 875 186
rect 1005 -16 1051 186
use hvDFM1sd2_CDNS_52468879185231  hvDFM1sd2_CDNS_52468879185231_0
timestamp 1701704242
transform 1 0 824 0 1 0
box -36 -36 92 236
use hvDFM1sd2_CDNS_52468879185231  hvDFM1sd2_CDNS_52468879185231_1
timestamp 1701704242
transform 1 0 648 0 1 0
box -36 -36 92 236
use hvDFM1sd2_CDNS_52468879185231  hvDFM1sd2_CDNS_52468879185231_2
timestamp 1701704242
transform 1 0 472 0 1 0
box -36 -36 92 236
use hvDFM1sd2_CDNS_52468879185231  hvDFM1sd2_CDNS_52468879185231_3
timestamp 1701704242
transform 1 0 296 0 1 0
box -36 -36 92 236
use hvDFM1sd2_CDNS_52468879185231  hvDFM1sd2_CDNS_52468879185231_4
timestamp 1701704242
transform 1 0 120 0 1 0
box -36 -36 92 236
use hvDFM1sd_CDNS_52468879185130  hvDFM1sd_CDNS_52468879185130_0
timestamp 1701704242
transform -1 0 0 0 1 0
box -36 -36 89 236
use hvDFM1sd_CDNS_52468879185130  hvDFM1sd_CDNS_52468879185130_1
timestamp 1701704242
transform 1 0 1000 0 1 0
box -36 -36 89 236
<< labels >>
flabel comment s -28 85 -28 85 0 FreeSans 300 0 0 0 S
flabel comment s 148 85 148 85 0 FreeSans 300 0 0 0 D
flabel comment s 324 85 324 85 0 FreeSans 300 0 0 0 S
flabel comment s 500 85 500 85 0 FreeSans 300 0 0 0 D
flabel comment s 676 85 676 85 0 FreeSans 300 0 0 0 S
flabel comment s 852 85 852 85 0 FreeSans 300 0 0 0 D
flabel comment s 1028 85 1028 85 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 78424438
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 78420920
<< end >>
