magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< obsli1 >>
rect 385 1369 1913 1388
rect 190 1225 256 1291
rect 385 1263 412 1369
rect 1886 1263 1913 1369
rect 385 1251 1913 1263
rect 2042 1225 2108 1291
rect 190 1203 230 1225
rect 2068 1203 2108 1225
rect 41 1179 230 1203
rect 41 1145 60 1179
rect 94 1145 230 1179
rect 41 1107 230 1145
rect 41 1073 60 1107
rect 94 1073 230 1107
rect 41 1035 230 1073
rect 41 1001 60 1035
rect 94 1001 230 1035
rect 41 963 230 1001
rect 41 929 60 963
rect 94 929 230 963
rect 41 891 230 929
rect 41 857 60 891
rect 94 857 230 891
rect 41 819 230 857
rect 41 785 60 819
rect 94 785 230 819
rect 41 747 230 785
rect 41 713 60 747
rect 94 713 230 747
rect 41 675 230 713
rect 41 641 60 675
rect 94 641 230 675
rect 41 603 230 641
rect 41 569 60 603
rect 94 569 230 603
rect 41 531 230 569
rect 41 497 60 531
rect 94 497 230 531
rect 41 459 230 497
rect 41 425 60 459
rect 94 425 230 459
rect 41 387 230 425
rect 41 353 60 387
rect 94 353 230 387
rect 41 315 230 353
rect 41 281 60 315
rect 94 281 230 315
rect 41 243 230 281
rect 41 209 60 243
rect 94 209 230 243
rect 41 185 230 209
rect 352 185 386 1203
rect 508 185 542 1203
rect 664 185 698 1203
rect 820 185 854 1203
rect 976 185 1010 1203
rect 1132 185 1166 1203
rect 1288 185 1322 1203
rect 1444 185 1478 1203
rect 1600 185 1634 1203
rect 1756 185 1790 1203
rect 1912 185 1946 1203
rect 2068 1179 2257 1203
rect 2068 1145 2204 1179
rect 2238 1145 2257 1179
rect 2068 1107 2257 1145
rect 2068 1073 2204 1107
rect 2238 1073 2257 1107
rect 2068 1035 2257 1073
rect 2068 1001 2204 1035
rect 2238 1001 2257 1035
rect 2068 963 2257 1001
rect 2068 929 2204 963
rect 2238 929 2257 963
rect 2068 891 2257 929
rect 2068 857 2204 891
rect 2238 857 2257 891
rect 2068 819 2257 857
rect 2068 785 2204 819
rect 2238 785 2257 819
rect 2068 747 2257 785
rect 2068 713 2204 747
rect 2238 713 2257 747
rect 2068 675 2257 713
rect 2068 641 2204 675
rect 2238 641 2257 675
rect 2068 603 2257 641
rect 2068 569 2204 603
rect 2238 569 2257 603
rect 2068 531 2257 569
rect 2068 497 2204 531
rect 2238 497 2257 531
rect 2068 459 2257 497
rect 2068 425 2204 459
rect 2238 425 2257 459
rect 2068 387 2257 425
rect 2068 353 2204 387
rect 2238 353 2257 387
rect 2068 315 2257 353
rect 2068 281 2204 315
rect 2238 281 2257 315
rect 2068 243 2257 281
rect 2068 209 2204 243
rect 2238 209 2257 243
rect 2068 185 2257 209
rect 190 163 230 185
rect 2068 163 2108 185
rect 190 97 256 163
rect 385 125 1913 137
rect 385 19 412 125
rect 1886 19 1913 125
rect 2042 97 2108 163
rect 385 0 1913 19
<< obsli1c >>
rect 412 1263 1886 1369
rect 60 1145 94 1179
rect 60 1073 94 1107
rect 60 1001 94 1035
rect 60 929 94 963
rect 60 857 94 891
rect 60 785 94 819
rect 60 713 94 747
rect 60 641 94 675
rect 60 569 94 603
rect 60 497 94 531
rect 60 425 94 459
rect 60 353 94 387
rect 60 281 94 315
rect 60 209 94 243
rect 2204 1145 2238 1179
rect 2204 1073 2238 1107
rect 2204 1001 2238 1035
rect 2204 929 2238 963
rect 2204 857 2238 891
rect 2204 785 2238 819
rect 2204 713 2238 747
rect 2204 641 2238 675
rect 2204 569 2238 603
rect 2204 497 2238 531
rect 2204 425 2238 459
rect 2204 353 2238 387
rect 2204 281 2238 315
rect 2204 209 2238 243
rect 412 19 1886 125
<< metal1 >>
rect 381 1369 1917 1388
rect 381 1263 412 1369
rect 1886 1263 1917 1369
rect 381 1251 1917 1263
rect 41 1179 100 1191
rect 41 1145 60 1179
rect 94 1145 100 1179
rect 41 1107 100 1145
rect 41 1073 60 1107
rect 94 1073 100 1107
rect 41 1035 100 1073
rect 41 1001 60 1035
rect 94 1001 100 1035
rect 41 963 100 1001
rect 41 929 60 963
rect 94 929 100 963
rect 41 891 100 929
rect 41 857 60 891
rect 94 857 100 891
rect 41 819 100 857
rect 41 785 60 819
rect 94 785 100 819
rect 41 747 100 785
rect 41 713 60 747
rect 94 713 100 747
rect 41 675 100 713
rect 41 641 60 675
rect 94 641 100 675
rect 41 603 100 641
rect 41 569 60 603
rect 94 569 100 603
rect 41 531 100 569
rect 41 497 60 531
rect 94 497 100 531
rect 41 459 100 497
rect 41 425 60 459
rect 94 425 100 459
rect 41 387 100 425
rect 41 353 60 387
rect 94 353 100 387
rect 41 315 100 353
rect 41 281 60 315
rect 94 281 100 315
rect 41 243 100 281
rect 41 209 60 243
rect 94 209 100 243
rect 41 197 100 209
rect 2198 1179 2257 1191
rect 2198 1145 2204 1179
rect 2238 1145 2257 1179
rect 2198 1107 2257 1145
rect 2198 1073 2204 1107
rect 2238 1073 2257 1107
rect 2198 1035 2257 1073
rect 2198 1001 2204 1035
rect 2238 1001 2257 1035
rect 2198 963 2257 1001
rect 2198 929 2204 963
rect 2238 929 2257 963
rect 2198 891 2257 929
rect 2198 857 2204 891
rect 2238 857 2257 891
rect 2198 819 2257 857
rect 2198 785 2204 819
rect 2238 785 2257 819
rect 2198 747 2257 785
rect 2198 713 2204 747
rect 2238 713 2257 747
rect 2198 675 2257 713
rect 2198 641 2204 675
rect 2238 641 2257 675
rect 2198 603 2257 641
rect 2198 569 2204 603
rect 2238 569 2257 603
rect 2198 531 2257 569
rect 2198 497 2204 531
rect 2238 497 2257 531
rect 2198 459 2257 497
rect 2198 425 2204 459
rect 2238 425 2257 459
rect 2198 387 2257 425
rect 2198 353 2204 387
rect 2238 353 2257 387
rect 2198 315 2257 353
rect 2198 281 2204 315
rect 2238 281 2257 315
rect 2198 243 2257 281
rect 2198 209 2204 243
rect 2238 209 2257 243
rect 2198 197 2257 209
rect 381 125 1917 137
rect 381 19 412 125
rect 1886 19 1917 125
rect 381 0 1917 19
<< obsm1 >>
rect 343 197 395 1191
rect 499 197 551 1191
rect 655 197 707 1191
rect 811 197 863 1191
rect 967 197 1019 1191
rect 1123 197 1175 1191
rect 1279 197 1331 1191
rect 1435 197 1487 1191
rect 1591 197 1643 1191
rect 1747 197 1799 1191
rect 1903 197 1955 1191
<< metal2 >>
rect 14 719 2284 1191
rect 14 197 2284 669
<< labels >>
rlabel metal2 s 14 719 2284 1191 6 DRAIN
port 1 nsew
rlabel metal1 s 381 1251 1917 1388 6 GATE
port 2 nsew
rlabel metal1 s 381 0 1917 137 6 GATE
port 2 nsew
rlabel metal2 s 14 197 2284 669 6 SOURCE
port 3 nsew
rlabel metal1 s 41 197 100 1191 6 SUBSTRATE
port 4 nsew
rlabel metal1 s 2198 197 2257 1191 6 SUBSTRATE
port 4 nsew
<< properties >>
string FIXED_BBOX 14 0 2284 1388
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 8617584
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 8564248
string device primitive
<< end >>
