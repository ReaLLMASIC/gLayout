magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< pwell >>
rect -76 -26 1076 626
<< mvnmos >>
rect 0 0 120 600
rect 176 0 296 600
rect 352 0 472 600
rect 528 0 648 600
rect 704 0 824 600
rect 880 0 1000 600
<< mvndiff >>
rect -50 0 0 600
rect 1000 0 1050 600
<< poly >>
rect 0 600 120 632
rect 0 -32 120 0
rect 176 600 296 632
rect 176 -32 296 0
rect 352 600 472 632
rect 352 -32 472 0
rect 528 600 648 632
rect 528 -32 648 0
rect 704 600 824 632
rect 704 -32 824 0
rect 880 600 1000 632
rect 880 -32 1000 0
<< locali >>
rect -45 -4 -11 538
rect 131 -4 165 538
rect 307 -4 341 538
rect 483 -4 517 538
rect 659 -4 693 538
rect 835 -4 869 538
rect 1011 -4 1045 538
use DFL1sd2_CDNS_52468879185189  DFL1sd2_CDNS_52468879185189_0
timestamp 1701704242
transform 1 0 824 0 1 0
box -26 -26 82 626
use DFL1sd2_CDNS_52468879185189  DFL1sd2_CDNS_52468879185189_1
timestamp 1701704242
transform 1 0 648 0 1 0
box -26 -26 82 626
use DFL1sd2_CDNS_52468879185189  DFL1sd2_CDNS_52468879185189_2
timestamp 1701704242
transform 1 0 472 0 1 0
box -26 -26 82 626
use DFL1sd2_CDNS_52468879185189  DFL1sd2_CDNS_52468879185189_3
timestamp 1701704242
transform 1 0 296 0 1 0
box -26 -26 82 626
use DFL1sd2_CDNS_52468879185189  DFL1sd2_CDNS_52468879185189_4
timestamp 1701704242
transform 1 0 120 0 1 0
box -26 -26 82 626
use hvDFL1sd2_CDNS_52468879185120  hvDFL1sd2_CDNS_52468879185120_0
timestamp 1701704242
transform -1 0 0 0 1 0
box -26 -26 82 626
use hvDFL1sd2_CDNS_52468879185120  hvDFL1sd2_CDNS_52468879185120_1
timestamp 1701704242
transform 1 0 1000 0 1 0
box -26 -26 82 626
<< labels >>
flabel comment s -28 267 -28 267 0 FreeSans 300 0 0 0 S
flabel comment s 148 267 148 267 0 FreeSans 300 0 0 0 D
flabel comment s 324 267 324 267 0 FreeSans 300 0 0 0 S
flabel comment s 500 267 500 267 0 FreeSans 300 0 0 0 D
flabel comment s 676 267 676 267 0 FreeSans 300 0 0 0 S
flabel comment s 852 267 852 267 0 FreeSans 300 0 0 0 D
flabel comment s 1028 267 1028 267 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 85620956
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85617572
<< end >>
