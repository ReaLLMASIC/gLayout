magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -119 -66 7863 1466
<< mvpmos >>
rect 0 0 100 1400
rect 156 0 256 1400
rect 312 0 412 1400
rect 468 0 568 1400
rect 624 0 724 1400
rect 780 0 880 1400
rect 936 0 1036 1400
rect 1092 0 1192 1400
rect 1248 0 1348 1400
rect 1404 0 1504 1400
rect 1560 0 1660 1400
rect 1716 0 1816 1400
rect 1872 0 1972 1400
rect 2028 0 2128 1400
rect 2184 0 2284 1400
rect 2340 0 2440 1400
rect 2496 0 2596 1400
rect 2652 0 2752 1400
rect 2808 0 2908 1400
rect 2964 0 3064 1400
rect 3120 0 3220 1400
rect 3276 0 3376 1400
rect 3432 0 3532 1400
rect 3588 0 3688 1400
rect 3744 0 3844 1400
rect 3900 0 4000 1400
rect 4056 0 4156 1400
rect 4212 0 4312 1400
rect 4368 0 4468 1400
rect 4524 0 4624 1400
rect 4680 0 4780 1400
rect 4836 0 4936 1400
rect 4992 0 5092 1400
rect 5148 0 5248 1400
rect 5304 0 5404 1400
rect 5460 0 5560 1400
rect 5616 0 5716 1400
rect 5772 0 5872 1400
rect 5928 0 6028 1400
rect 6084 0 6184 1400
rect 6240 0 6340 1400
rect 6396 0 6496 1400
rect 6552 0 6652 1400
rect 6708 0 6808 1400
rect 6864 0 6964 1400
rect 7020 0 7120 1400
rect 7176 0 7276 1400
rect 7332 0 7432 1400
rect 7488 0 7588 1400
rect 7644 0 7744 1400
<< mvpdiff >>
rect -50 0 0 1400
rect 7744 0 7794 1400
<< poly >>
rect 0 1400 100 1426
rect 0 -26 100 0
rect 156 1400 256 1426
rect 156 -26 256 0
rect 312 1400 412 1426
rect 312 -26 412 0
rect 468 1400 568 1426
rect 468 -26 568 0
rect 624 1400 724 1426
rect 624 -26 724 0
rect 780 1400 880 1426
rect 780 -26 880 0
rect 936 1400 1036 1426
rect 936 -26 1036 0
rect 1092 1400 1192 1426
rect 1092 -26 1192 0
rect 1248 1400 1348 1426
rect 1248 -26 1348 0
rect 1404 1400 1504 1426
rect 1404 -26 1504 0
rect 1560 1400 1660 1426
rect 1560 -26 1660 0
rect 1716 1400 1816 1426
rect 1716 -26 1816 0
rect 1872 1400 1972 1426
rect 1872 -26 1972 0
rect 2028 1400 2128 1426
rect 2028 -26 2128 0
rect 2184 1400 2284 1426
rect 2184 -26 2284 0
rect 2340 1400 2440 1426
rect 2340 -26 2440 0
rect 2496 1400 2596 1426
rect 2496 -26 2596 0
rect 2652 1400 2752 1426
rect 2652 -26 2752 0
rect 2808 1400 2908 1426
rect 2808 -26 2908 0
rect 2964 1400 3064 1426
rect 2964 -26 3064 0
rect 3120 1400 3220 1426
rect 3120 -26 3220 0
rect 3276 1400 3376 1426
rect 3276 -26 3376 0
rect 3432 1400 3532 1426
rect 3432 -26 3532 0
rect 3588 1400 3688 1426
rect 3588 -26 3688 0
rect 3744 1400 3844 1426
rect 3744 -26 3844 0
rect 3900 1400 4000 1426
rect 3900 -26 4000 0
rect 4056 1400 4156 1426
rect 4056 -26 4156 0
rect 4212 1400 4312 1426
rect 4212 -26 4312 0
rect 4368 1400 4468 1426
rect 4368 -26 4468 0
rect 4524 1400 4624 1426
rect 4524 -26 4624 0
rect 4680 1400 4780 1426
rect 4680 -26 4780 0
rect 4836 1400 4936 1426
rect 4836 -26 4936 0
rect 4992 1400 5092 1426
rect 4992 -26 5092 0
rect 5148 1400 5248 1426
rect 5148 -26 5248 0
rect 5304 1400 5404 1426
rect 5304 -26 5404 0
rect 5460 1400 5560 1426
rect 5460 -26 5560 0
rect 5616 1400 5716 1426
rect 5616 -26 5716 0
rect 5772 1400 5872 1426
rect 5772 -26 5872 0
rect 5928 1400 6028 1426
rect 5928 -26 6028 0
rect 6084 1400 6184 1426
rect 6084 -26 6184 0
rect 6240 1400 6340 1426
rect 6240 -26 6340 0
rect 6396 1400 6496 1426
rect 6396 -26 6496 0
rect 6552 1400 6652 1426
rect 6552 -26 6652 0
rect 6708 1400 6808 1426
rect 6708 -26 6808 0
rect 6864 1400 6964 1426
rect 6864 -26 6964 0
rect 7020 1400 7120 1426
rect 7020 -26 7120 0
rect 7176 1400 7276 1426
rect 7176 -26 7276 0
rect 7332 1400 7432 1426
rect 7332 -26 7432 0
rect 7488 1400 7588 1426
rect 7488 -26 7588 0
rect 7644 1400 7744 1426
rect 7644 -26 7744 0
<< locali >>
rect -45 -4 -11 1354
rect 111 -4 145 1354
rect 267 -4 301 1354
rect 423 -4 457 1354
rect 579 -4 613 1354
rect 735 -4 769 1354
rect 891 -4 925 1354
rect 1047 -4 1081 1354
rect 1203 -4 1237 1354
rect 1359 -4 1393 1354
rect 1515 -4 1549 1354
rect 1671 -4 1705 1354
rect 1827 -4 1861 1354
rect 1983 -4 2017 1354
rect 2139 -4 2173 1354
rect 2295 -4 2329 1354
rect 2451 -4 2485 1354
rect 2607 -4 2641 1354
rect 2763 -4 2797 1354
rect 2919 -4 2953 1354
rect 3075 -4 3109 1354
rect 3231 -4 3265 1354
rect 3387 -4 3421 1354
rect 3543 -4 3577 1354
rect 3699 -4 3733 1354
rect 3855 -4 3889 1354
rect 4011 -4 4045 1354
rect 4167 -4 4201 1354
rect 4323 -4 4357 1354
rect 4479 -4 4513 1354
rect 4635 -4 4669 1354
rect 4791 -4 4825 1354
rect 4947 -4 4981 1354
rect 5103 -4 5137 1354
rect 5259 -4 5293 1354
rect 5415 -4 5449 1354
rect 5571 -4 5605 1354
rect 5727 -4 5761 1354
rect 5883 -4 5917 1354
rect 6039 -4 6073 1354
rect 6195 -4 6229 1354
rect 6351 -4 6385 1354
rect 6507 -4 6541 1354
rect 6663 -4 6697 1354
rect 6819 -4 6853 1354
rect 6975 -4 7009 1354
rect 7131 -4 7165 1354
rect 7287 -4 7321 1354
rect 7443 -4 7477 1354
rect 7599 -4 7633 1354
rect 7755 -4 7789 1354
use DFL1sd2_CDNS_5246887918574  DFL1sd2_CDNS_5246887918574_0
timestamp 1701704242
transform 1 0 7588 0 1 0
box -36 -36 92 1436
use DFL1sd2_CDNS_5246887918574  DFL1sd2_CDNS_5246887918574_1
timestamp 1701704242
transform 1 0 7432 0 1 0
box -36 -36 92 1436
use DFL1sd2_CDNS_5246887918574  DFL1sd2_CDNS_5246887918574_2
timestamp 1701704242
transform 1 0 7276 0 1 0
box -36 -36 92 1436
use DFL1sd2_CDNS_5246887918574  DFL1sd2_CDNS_5246887918574_3
timestamp 1701704242
transform 1 0 7120 0 1 0
box -36 -36 92 1436
use DFL1sd2_CDNS_5246887918574  DFL1sd2_CDNS_5246887918574_4
timestamp 1701704242
transform 1 0 6964 0 1 0
box -36 -36 92 1436
use DFL1sd2_CDNS_5246887918574  DFL1sd2_CDNS_5246887918574_5
timestamp 1701704242
transform 1 0 6808 0 1 0
box -36 -36 92 1436
use DFL1sd2_CDNS_5246887918574  DFL1sd2_CDNS_5246887918574_6
timestamp 1701704242
transform 1 0 6652 0 1 0
box -36 -36 92 1436
use DFL1sd2_CDNS_5246887918574  DFL1sd2_CDNS_5246887918574_7
timestamp 1701704242
transform 1 0 6496 0 1 0
box -36 -36 92 1436
use DFL1sd2_CDNS_5246887918574  DFL1sd2_CDNS_5246887918574_8
timestamp 1701704242
transform 1 0 6340 0 1 0
box -36 -36 92 1436
use DFL1sd2_CDNS_5246887918574  DFL1sd2_CDNS_5246887918574_9
timestamp 1701704242
transform 1 0 6184 0 1 0
box -36 -36 92 1436
use DFL1sd2_CDNS_5246887918574  DFL1sd2_CDNS_5246887918574_10
timestamp 1701704242
transform 1 0 6028 0 1 0
box -36 -36 92 1436
use DFL1sd2_CDNS_5246887918574  DFL1sd2_CDNS_5246887918574_11
timestamp 1701704242
transform 1 0 5872 0 1 0
box -36 -36 92 1436
use DFL1sd2_CDNS_5246887918574  DFL1sd2_CDNS_5246887918574_12
timestamp 1701704242
transform 1 0 5716 0 1 0
box -36 -36 92 1436
use DFL1sd2_CDNS_5246887918574  DFL1sd2_CDNS_5246887918574_13
timestamp 1701704242
transform 1 0 5560 0 1 0
box -36 -36 92 1436
use DFL1sd2_CDNS_5246887918574  DFL1sd2_CDNS_5246887918574_14
timestamp 1701704242
transform 1 0 5404 0 1 0
box -36 -36 92 1436
use DFL1sd2_CDNS_5246887918574  DFL1sd2_CDNS_5246887918574_15
timestamp 1701704242
transform 1 0 5248 0 1 0
box -36 -36 92 1436
use DFL1sd2_CDNS_5246887918574  DFL1sd2_CDNS_5246887918574_16
timestamp 1701704242
transform 1 0 5092 0 1 0
box -36 -36 92 1436
use DFL1sd2_CDNS_5246887918574  DFL1sd2_CDNS_5246887918574_17
timestamp 1701704242
transform 1 0 4936 0 1 0
box -36 -36 92 1436
use DFL1sd2_CDNS_5246887918574  DFL1sd2_CDNS_5246887918574_18
timestamp 1701704242
transform 1 0 4780 0 1 0
box -36 -36 92 1436
use DFL1sd2_CDNS_5246887918574  DFL1sd2_CDNS_5246887918574_19
timestamp 1701704242
transform 1 0 4624 0 1 0
box -36 -36 92 1436
use DFL1sd2_CDNS_5246887918574  DFL1sd2_CDNS_5246887918574_20
timestamp 1701704242
transform 1 0 4468 0 1 0
box -36 -36 92 1436
use DFL1sd2_CDNS_5246887918574  DFL1sd2_CDNS_5246887918574_21
timestamp 1701704242
transform 1 0 4312 0 1 0
box -36 -36 92 1436
use DFL1sd2_CDNS_5246887918574  DFL1sd2_CDNS_5246887918574_22
timestamp 1701704242
transform 1 0 4156 0 1 0
box -36 -36 92 1436
use DFL1sd2_CDNS_5246887918574  DFL1sd2_CDNS_5246887918574_23
timestamp 1701704242
transform 1 0 4000 0 1 0
box -36 -36 92 1436
use DFL1sd2_CDNS_5246887918574  DFL1sd2_CDNS_5246887918574_24
timestamp 1701704242
transform 1 0 3844 0 1 0
box -36 -36 92 1436
use DFL1sd2_CDNS_5246887918574  DFL1sd2_CDNS_5246887918574_25
timestamp 1701704242
transform 1 0 3688 0 1 0
box -36 -36 92 1436
use DFL1sd2_CDNS_5246887918574  DFL1sd2_CDNS_5246887918574_26
timestamp 1701704242
transform 1 0 3532 0 1 0
box -36 -36 92 1436
use DFL1sd2_CDNS_5246887918574  DFL1sd2_CDNS_5246887918574_27
timestamp 1701704242
transform 1 0 3376 0 1 0
box -36 -36 92 1436
use DFL1sd2_CDNS_5246887918574  DFL1sd2_CDNS_5246887918574_28
timestamp 1701704242
transform 1 0 3220 0 1 0
box -36 -36 92 1436
use DFL1sd2_CDNS_5246887918574  DFL1sd2_CDNS_5246887918574_29
timestamp 1701704242
transform 1 0 3064 0 1 0
box -36 -36 92 1436
use DFL1sd2_CDNS_5246887918574  DFL1sd2_CDNS_5246887918574_30
timestamp 1701704242
transform 1 0 2908 0 1 0
box -36 -36 92 1436
use DFL1sd2_CDNS_5246887918574  DFL1sd2_CDNS_5246887918574_31
timestamp 1701704242
transform 1 0 2752 0 1 0
box -36 -36 92 1436
use DFL1sd2_CDNS_5246887918574  DFL1sd2_CDNS_5246887918574_32
timestamp 1701704242
transform 1 0 2596 0 1 0
box -36 -36 92 1436
use DFL1sd2_CDNS_5246887918574  DFL1sd2_CDNS_5246887918574_33
timestamp 1701704242
transform 1 0 2440 0 1 0
box -36 -36 92 1436
use DFL1sd2_CDNS_5246887918574  DFL1sd2_CDNS_5246887918574_34
timestamp 1701704242
transform 1 0 2284 0 1 0
box -36 -36 92 1436
use DFL1sd2_CDNS_5246887918574  DFL1sd2_CDNS_5246887918574_35
timestamp 1701704242
transform 1 0 2128 0 1 0
box -36 -36 92 1436
use DFL1sd2_CDNS_5246887918574  DFL1sd2_CDNS_5246887918574_36
timestamp 1701704242
transform 1 0 1972 0 1 0
box -36 -36 92 1436
use DFL1sd2_CDNS_5246887918574  DFL1sd2_CDNS_5246887918574_37
timestamp 1701704242
transform 1 0 1816 0 1 0
box -36 -36 92 1436
use DFL1sd2_CDNS_5246887918574  DFL1sd2_CDNS_5246887918574_38
timestamp 1701704242
transform 1 0 1660 0 1 0
box -36 -36 92 1436
use DFL1sd2_CDNS_5246887918574  DFL1sd2_CDNS_5246887918574_39
timestamp 1701704242
transform 1 0 1504 0 1 0
box -36 -36 92 1436
use DFL1sd2_CDNS_5246887918574  DFL1sd2_CDNS_5246887918574_40
timestamp 1701704242
transform 1 0 1348 0 1 0
box -36 -36 92 1436
use DFL1sd2_CDNS_5246887918574  DFL1sd2_CDNS_5246887918574_41
timestamp 1701704242
transform 1 0 1192 0 1 0
box -36 -36 92 1436
use DFL1sd2_CDNS_5246887918574  DFL1sd2_CDNS_5246887918574_42
timestamp 1701704242
transform 1 0 1036 0 1 0
box -36 -36 92 1436
use DFL1sd2_CDNS_5246887918574  DFL1sd2_CDNS_5246887918574_43
timestamp 1701704242
transform 1 0 880 0 1 0
box -36 -36 92 1436
use DFL1sd2_CDNS_5246887918574  DFL1sd2_CDNS_5246887918574_44
timestamp 1701704242
transform 1 0 724 0 1 0
box -36 -36 92 1436
use DFL1sd2_CDNS_5246887918574  DFL1sd2_CDNS_5246887918574_45
timestamp 1701704242
transform 1 0 568 0 1 0
box -36 -36 92 1436
use DFL1sd2_CDNS_5246887918574  DFL1sd2_CDNS_5246887918574_46
timestamp 1701704242
transform 1 0 412 0 1 0
box -36 -36 92 1436
use DFL1sd2_CDNS_5246887918574  DFL1sd2_CDNS_5246887918574_47
timestamp 1701704242
transform 1 0 256 0 1 0
box -36 -36 92 1436
use DFL1sd2_CDNS_5246887918574  DFL1sd2_CDNS_5246887918574_48
timestamp 1701704242
transform 1 0 100 0 1 0
box -36 -36 92 1436
use DFL1sd_CDNS_52468879185620  DFL1sd_CDNS_52468879185620_0
timestamp 1701704242
transform -1 0 0 0 1 0
box -36 -36 89 1436
use DFL1sd_CDNS_52468879185620  DFL1sd_CDNS_52468879185620_1
timestamp 1701704242
transform 1 0 7744 0 1 0
box -36 -36 89 1436
<< labels >>
flabel comment s -28 675 -28 675 0 FreeSans 300 0 0 0 S
flabel comment s 128 675 128 675 0 FreeSans 300 0 0 0 D
flabel comment s 284 675 284 675 0 FreeSans 300 0 0 0 S
flabel comment s 440 675 440 675 0 FreeSans 300 0 0 0 D
flabel comment s 596 675 596 675 0 FreeSans 300 0 0 0 S
flabel comment s 752 675 752 675 0 FreeSans 300 0 0 0 D
flabel comment s 908 675 908 675 0 FreeSans 300 0 0 0 S
flabel comment s 1064 675 1064 675 0 FreeSans 300 0 0 0 D
flabel comment s 1220 675 1220 675 0 FreeSans 300 0 0 0 S
flabel comment s 1376 675 1376 675 0 FreeSans 300 0 0 0 D
flabel comment s 1532 675 1532 675 0 FreeSans 300 0 0 0 S
flabel comment s 1688 675 1688 675 0 FreeSans 300 0 0 0 D
flabel comment s 1844 675 1844 675 0 FreeSans 300 0 0 0 S
flabel comment s 2000 675 2000 675 0 FreeSans 300 0 0 0 D
flabel comment s 2156 675 2156 675 0 FreeSans 300 0 0 0 S
flabel comment s 2312 675 2312 675 0 FreeSans 300 0 0 0 D
flabel comment s 2468 675 2468 675 0 FreeSans 300 0 0 0 S
flabel comment s 2624 675 2624 675 0 FreeSans 300 0 0 0 D
flabel comment s 2780 675 2780 675 0 FreeSans 300 0 0 0 S
flabel comment s 2936 675 2936 675 0 FreeSans 300 0 0 0 D
flabel comment s 3092 675 3092 675 0 FreeSans 300 0 0 0 S
flabel comment s 3248 675 3248 675 0 FreeSans 300 0 0 0 D
flabel comment s 3404 675 3404 675 0 FreeSans 300 0 0 0 S
flabel comment s 3560 675 3560 675 0 FreeSans 300 0 0 0 D
flabel comment s 3716 675 3716 675 0 FreeSans 300 0 0 0 S
flabel comment s 3872 675 3872 675 0 FreeSans 300 0 0 0 D
flabel comment s 4028 675 4028 675 0 FreeSans 300 0 0 0 S
flabel comment s 4184 675 4184 675 0 FreeSans 300 0 0 0 D
flabel comment s 4340 675 4340 675 0 FreeSans 300 0 0 0 S
flabel comment s 4496 675 4496 675 0 FreeSans 300 0 0 0 D
flabel comment s 4652 675 4652 675 0 FreeSans 300 0 0 0 S
flabel comment s 4808 675 4808 675 0 FreeSans 300 0 0 0 D
flabel comment s 4964 675 4964 675 0 FreeSans 300 0 0 0 S
flabel comment s 5120 675 5120 675 0 FreeSans 300 0 0 0 D
flabel comment s 5276 675 5276 675 0 FreeSans 300 0 0 0 S
flabel comment s 5432 675 5432 675 0 FreeSans 300 0 0 0 D
flabel comment s 5588 675 5588 675 0 FreeSans 300 0 0 0 S
flabel comment s 5744 675 5744 675 0 FreeSans 300 0 0 0 D
flabel comment s 5900 675 5900 675 0 FreeSans 300 0 0 0 S
flabel comment s 6056 675 6056 675 0 FreeSans 300 0 0 0 D
flabel comment s 6212 675 6212 675 0 FreeSans 300 0 0 0 S
flabel comment s 6368 675 6368 675 0 FreeSans 300 0 0 0 D
flabel comment s 6524 675 6524 675 0 FreeSans 300 0 0 0 S
flabel comment s 6680 675 6680 675 0 FreeSans 300 0 0 0 D
flabel comment s 6836 675 6836 675 0 FreeSans 300 0 0 0 S
flabel comment s 6992 675 6992 675 0 FreeSans 300 0 0 0 D
flabel comment s 7148 675 7148 675 0 FreeSans 300 0 0 0 S
flabel comment s 7304 675 7304 675 0 FreeSans 300 0 0 0 D
flabel comment s 7460 675 7460 675 0 FreeSans 300 0 0 0 S
flabel comment s 7616 675 7616 675 0 FreeSans 300 0 0 0 D
flabel comment s 7772 675 7772 675 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 34375568
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 34350250
<< end >>
