magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< pwell >>
rect -79 -26 199 226
<< mvnmos >>
rect 0 0 120 200
<< mvndiff >>
rect -53 182 0 200
rect -53 148 -45 182
rect -11 148 0 182
rect -53 114 0 148
rect -53 80 -45 114
rect -11 80 0 114
rect -53 46 0 80
rect -53 12 -45 46
rect -11 12 0 46
rect -53 0 0 12
rect 120 182 173 200
rect 120 148 131 182
rect 165 148 173 182
rect 120 114 173 148
rect 120 80 131 114
rect 165 80 173 114
rect 120 46 173 80
rect 120 12 131 46
rect 165 12 173 46
rect 120 0 173 12
<< mvndiffc >>
rect -45 148 -11 182
rect -45 80 -11 114
rect -45 12 -11 46
rect 131 148 165 182
rect 131 80 165 114
rect 131 12 165 46
<< poly >>
rect 0 200 120 232
rect 0 -32 120 0
<< locali >>
rect -45 182 -11 198
rect -45 114 -11 148
rect -45 46 -11 80
rect -45 -4 -11 12
rect 131 182 165 198
rect 131 114 165 148
rect 131 46 165 80
rect 131 -4 165 12
use DFL1sd_CDNS_5246887918538  DFL1sd_CDNS_5246887918538_0
timestamp 1701704242
transform -1 0 0 0 1 0
box 0 0 1 1
use DFL1sd_CDNS_5246887918538  DFL1sd_CDNS_5246887918538_1
timestamp 1701704242
transform 1 0 120 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s -28 97 -28 97 0 FreeSans 300 0 0 0 S
flabel comment s 148 97 148 97 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 80609116
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 80608230
<< end >>
