magic
tech sky130B
timestamp 1701704242
<< viali >>
rect 0 0 161 377
<< metal1 >>
rect -6 377 167 380
rect -6 0 0 377
rect 161 0 167 377
rect -6 -3 167 0
<< properties >>
string GDS_END 95629312
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 95625660
<< end >>
