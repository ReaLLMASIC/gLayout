magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< pwell >>
rect -26 -26 82 626
<< ndiff >>
rect 0 522 56 600
rect 0 488 11 522
rect 45 488 56 522
rect 0 454 56 488
rect 0 420 11 454
rect 45 420 56 454
rect 0 386 56 420
rect 0 352 11 386
rect 45 352 56 386
rect 0 318 56 352
rect 0 284 11 318
rect 45 284 56 318
rect 0 250 56 284
rect 0 216 11 250
rect 45 216 56 250
rect 0 182 56 216
rect 0 148 11 182
rect 45 148 56 182
rect 0 114 56 148
rect 0 80 11 114
rect 45 80 56 114
rect 0 46 56 80
rect 0 12 11 46
rect 45 12 56 46
rect 0 0 56 12
<< ndiffc >>
rect 11 488 45 522
rect 11 420 45 454
rect 11 352 45 386
rect 11 284 45 318
rect 11 216 45 250
rect 11 148 45 182
rect 11 80 45 114
rect 11 12 45 46
<< locali >>
rect 11 534 45 538
rect 11 462 45 488
rect 11 390 45 420
rect 11 318 45 352
rect 11 250 45 284
rect 11 182 45 212
rect 11 114 45 140
rect 11 46 45 68
<< viali >>
rect 11 522 45 534
rect 11 500 45 522
rect 11 454 45 462
rect 11 428 45 454
rect 11 386 45 390
rect 11 356 45 386
rect 11 284 45 318
rect 11 216 45 246
rect 11 212 45 216
rect 11 148 45 174
rect 11 140 45 148
rect 11 80 45 102
rect 11 68 45 80
rect 11 12 45 30
rect 11 -4 45 12
<< metal1 >>
rect 5 534 51 546
rect 5 500 11 534
rect 45 500 51 534
rect 5 462 51 500
rect 5 428 11 462
rect 45 428 51 462
rect 5 390 51 428
rect 5 356 11 390
rect 45 356 51 390
rect 5 318 51 356
rect 5 284 11 318
rect 45 284 51 318
rect 5 246 51 284
rect 5 212 11 246
rect 45 212 51 246
rect 5 174 51 212
rect 5 140 11 174
rect 45 140 51 174
rect 5 102 51 140
rect 5 68 11 102
rect 45 68 51 102
rect 5 30 51 68
rect 5 -4 11 30
rect 45 -4 51 30
rect 5 -16 51 -4
<< properties >>
string GDS_END 86609242
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86607958
<< end >>
