magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -429 2590 549 2758
rect -429 102 -261 2590
rect 413 2550 549 2590
rect 413 2358 3374 2550
rect 413 102 549 2358
rect -429 -66 549 102
<< pwell >>
rect -201 2444 353 2530
rect -201 248 -115 2444
rect 267 248 353 2444
rect -201 162 353 248
<< mvpsubdiff >>
rect -175 2470 -151 2504
rect -117 2470 -82 2504
rect -48 2470 -13 2504
rect 21 2470 55 2504
rect 89 2470 123 2504
rect 157 2470 191 2504
rect 225 2470 327 2504
rect -175 2394 -141 2470
rect 293 2400 327 2436
rect -175 2326 -141 2360
rect -175 2257 -141 2292
rect -175 2188 -141 2223
rect -175 2119 -141 2154
rect -175 2050 -141 2085
rect -175 1981 -141 2016
rect -175 1912 -141 1947
rect -175 1843 -141 1878
rect -175 1774 -141 1809
rect -175 1705 -141 1740
rect -175 1636 -141 1671
rect -175 1567 -141 1602
rect -175 1498 -141 1533
rect -175 1429 -141 1464
rect -175 1360 -141 1395
rect -175 1291 -141 1326
rect -175 1222 -141 1257
rect -175 1153 -141 1188
rect -175 1084 -141 1119
rect -175 1015 -141 1050
rect -175 946 -141 981
rect -175 877 -141 912
rect -175 808 -141 843
rect -175 739 -141 774
rect -175 670 -141 705
rect -175 601 -141 636
rect -175 532 -141 567
rect -175 463 -141 498
rect -175 394 -141 429
rect -175 325 -141 360
rect 293 2330 327 2366
rect 293 2260 327 2296
rect 293 2190 327 2226
rect 293 2120 327 2156
rect 293 2051 327 2086
rect 293 1982 327 2017
rect 293 1913 327 1948
rect 293 1844 327 1879
rect 293 1775 327 1810
rect 293 1706 327 1741
rect 293 1637 327 1672
rect 293 1568 327 1603
rect 293 1499 327 1534
rect 293 1430 327 1465
rect 293 1361 327 1396
rect 293 1292 327 1327
rect 293 1223 327 1258
rect 293 1154 327 1189
rect 293 1085 327 1120
rect 293 1016 327 1051
rect 293 947 327 982
rect 293 878 327 913
rect 293 809 327 844
rect 293 740 327 775
rect 293 671 327 706
rect 293 602 327 637
rect 293 533 327 568
rect 293 464 327 499
rect 293 395 327 430
rect 293 326 327 361
rect -175 256 -141 291
rect -175 188 -53 222
rect -19 188 25 222
rect 59 188 103 222
rect 137 188 181 222
rect 215 188 259 222
rect 293 188 327 292
<< mvnsubdiff >>
rect -361 2656 -337 2690
rect -303 2656 -266 2690
rect -232 2656 -195 2690
rect -161 2656 -124 2690
rect -90 2656 -53 2690
rect -19 2656 18 2690
rect 52 2656 89 2690
rect 123 2656 160 2690
rect 194 2656 231 2690
rect 265 2656 302 2690
rect 336 2656 373 2690
rect 407 2656 530 2690
rect -361 2560 -327 2656
rect -361 2491 -327 2526
rect 513 2622 530 2656
rect 479 2616 530 2622
rect 479 2587 513 2616
rect 479 2518 513 2553
rect -361 2422 -327 2457
rect -361 2353 -327 2388
rect -361 2284 -327 2319
rect -361 2215 -327 2250
rect -361 2146 -327 2181
rect -361 2077 -327 2112
rect -361 2008 -327 2043
rect -361 1939 -327 1974
rect -361 1870 -327 1905
rect -361 1801 -327 1836
rect -361 1732 -327 1767
rect -361 1663 -327 1698
rect -361 1594 -327 1629
rect -361 1525 -327 1560
rect -361 1456 -327 1491
rect -361 1387 -327 1422
rect -361 1318 -327 1353
rect -361 1249 -327 1284
rect -361 1180 -327 1215
rect -361 1111 -327 1146
rect -361 1042 -327 1077
rect -361 973 -327 1008
rect -361 904 -327 939
rect -361 835 -327 870
rect -361 766 -327 801
rect -361 697 -327 732
rect -361 628 -327 663
rect -361 558 -327 594
rect -361 488 -327 524
rect -361 418 -327 454
rect -361 348 -327 384
rect -361 278 -327 314
rect -361 208 -327 244
rect 479 2449 513 2484
rect 479 2380 513 2415
rect 479 2312 513 2346
rect 513 2278 530 2292
rect 479 2244 530 2278
rect 513 2210 530 2244
rect 479 2176 530 2210
rect 513 2142 530 2176
rect 479 2108 530 2142
rect 513 2074 530 2108
rect 479 2040 530 2074
rect 513 2006 530 2040
rect 479 1972 530 2006
rect 513 1938 530 1972
rect 479 1904 530 1938
rect 513 1870 530 1904
rect 479 1836 530 1870
rect 513 1802 530 1836
rect 479 1768 530 1802
rect 513 1734 530 1768
rect 479 1700 530 1734
rect 513 1666 530 1700
rect 479 1632 530 1666
rect 513 1598 530 1632
rect 479 1564 530 1598
rect 513 1530 530 1564
rect 479 1496 530 1530
rect 513 1462 530 1496
rect 479 1428 530 1462
rect 513 1394 530 1428
rect 479 1360 530 1394
rect 513 1326 530 1360
rect 479 1292 530 1326
rect 513 1258 530 1292
rect 479 1224 530 1258
rect 513 1190 530 1224
rect 479 1156 530 1190
rect 513 1122 530 1156
rect 479 1088 530 1122
rect 513 1054 530 1088
rect 479 1020 530 1054
rect 513 986 530 1020
rect 479 952 530 986
rect 513 918 530 952
rect 479 884 530 918
rect 513 850 530 884
rect 479 816 530 850
rect 513 782 530 816
rect 479 748 530 782
rect 513 714 530 748
rect 479 680 530 714
rect 513 646 530 680
rect 479 612 530 646
rect 513 578 530 612
rect 479 544 530 578
rect 513 510 530 544
rect 479 476 530 510
rect 513 442 530 476
rect 479 408 530 442
rect 513 374 530 408
rect 479 340 530 374
rect 513 306 530 340
rect 479 272 530 306
rect 513 238 530 272
rect 479 204 530 238
rect -361 138 -327 174
rect -361 68 -327 104
rect 513 170 530 204
rect 479 136 530 170
rect 513 102 530 136
rect -361 0 -255 34
rect -221 0 -185 34
rect -151 0 -115 34
rect -81 0 -45 34
rect -11 0 25 34
rect 59 0 95 34
rect 129 0 165 34
rect 199 0 235 34
rect 269 0 305 34
rect 339 0 375 34
rect 409 0 445 34
rect 479 0 530 102
<< mvpsubdiffcont >>
rect -151 2470 -117 2504
rect -82 2470 -48 2504
rect -13 2470 21 2504
rect 55 2470 89 2504
rect 123 2470 157 2504
rect 191 2470 225 2504
rect -175 2360 -141 2394
rect 293 2436 327 2470
rect -175 2292 -141 2326
rect -175 2223 -141 2257
rect -175 2154 -141 2188
rect -175 2085 -141 2119
rect -175 2016 -141 2050
rect -175 1947 -141 1981
rect -175 1878 -141 1912
rect -175 1809 -141 1843
rect -175 1740 -141 1774
rect -175 1671 -141 1705
rect -175 1602 -141 1636
rect -175 1533 -141 1567
rect -175 1464 -141 1498
rect -175 1395 -141 1429
rect -175 1326 -141 1360
rect -175 1257 -141 1291
rect -175 1188 -141 1222
rect -175 1119 -141 1153
rect -175 1050 -141 1084
rect -175 981 -141 1015
rect -175 912 -141 946
rect -175 843 -141 877
rect -175 774 -141 808
rect -175 705 -141 739
rect -175 636 -141 670
rect -175 567 -141 601
rect -175 498 -141 532
rect -175 429 -141 463
rect -175 360 -141 394
rect -175 291 -141 325
rect 293 2366 327 2400
rect 293 2296 327 2330
rect 293 2226 327 2260
rect 293 2156 327 2190
rect 293 2086 327 2120
rect 293 2017 327 2051
rect 293 1948 327 1982
rect 293 1879 327 1913
rect 293 1810 327 1844
rect 293 1741 327 1775
rect 293 1672 327 1706
rect 293 1603 327 1637
rect 293 1534 327 1568
rect 293 1465 327 1499
rect 293 1396 327 1430
rect 293 1327 327 1361
rect 293 1258 327 1292
rect 293 1189 327 1223
rect 293 1120 327 1154
rect 293 1051 327 1085
rect 293 982 327 1016
rect 293 913 327 947
rect 293 844 327 878
rect 293 775 327 809
rect 293 706 327 740
rect 293 637 327 671
rect 293 568 327 602
rect 293 499 327 533
rect 293 430 327 464
rect 293 361 327 395
rect -175 222 -141 256
rect 293 292 327 326
rect -53 188 -19 222
rect 25 188 59 222
rect 103 188 137 222
rect 181 188 215 222
rect 259 188 293 222
<< mvnsubdiffcont >>
rect -337 2656 -303 2690
rect -266 2656 -232 2690
rect -195 2656 -161 2690
rect -124 2656 -90 2690
rect -53 2656 -19 2690
rect 18 2656 52 2690
rect 89 2656 123 2690
rect 160 2656 194 2690
rect 231 2656 265 2690
rect 302 2656 336 2690
rect 373 2656 407 2690
rect -361 2526 -327 2560
rect 479 2622 513 2656
rect 479 2553 513 2587
rect -361 2457 -327 2491
rect -361 2388 -327 2422
rect -361 2319 -327 2353
rect -361 2250 -327 2284
rect -361 2181 -327 2215
rect -361 2112 -327 2146
rect -361 2043 -327 2077
rect -361 1974 -327 2008
rect -361 1905 -327 1939
rect -361 1836 -327 1870
rect -361 1767 -327 1801
rect -361 1698 -327 1732
rect -361 1629 -327 1663
rect -361 1560 -327 1594
rect -361 1491 -327 1525
rect -361 1422 -327 1456
rect -361 1353 -327 1387
rect -361 1284 -327 1318
rect -361 1215 -327 1249
rect -361 1146 -327 1180
rect -361 1077 -327 1111
rect -361 1008 -327 1042
rect -361 939 -327 973
rect -361 870 -327 904
rect -361 801 -327 835
rect -361 732 -327 766
rect -361 663 -327 697
rect -361 594 -327 628
rect -361 524 -327 558
rect -361 454 -327 488
rect -361 384 -327 418
rect -361 314 -327 348
rect -361 244 -327 278
rect -361 174 -327 208
rect 479 2484 513 2518
rect 479 2415 513 2449
rect 479 2346 513 2380
rect 479 2278 513 2312
rect 479 2210 513 2244
rect 479 2142 513 2176
rect 479 2074 513 2108
rect 479 2006 513 2040
rect 479 1938 513 1972
rect 479 1870 513 1904
rect 479 1802 513 1836
rect 479 1734 513 1768
rect 479 1666 513 1700
rect 479 1598 513 1632
rect 479 1530 513 1564
rect 479 1462 513 1496
rect 479 1394 513 1428
rect 479 1326 513 1360
rect 479 1258 513 1292
rect 479 1190 513 1224
rect 479 1122 513 1156
rect 479 1054 513 1088
rect 479 986 513 1020
rect 479 918 513 952
rect 479 850 513 884
rect 479 782 513 816
rect 479 714 513 748
rect 479 646 513 680
rect 479 578 513 612
rect 479 510 513 544
rect 479 442 513 476
rect 479 374 513 408
rect 479 306 513 340
rect 479 238 513 272
rect -361 104 -327 138
rect -361 34 -327 68
rect 479 170 513 204
rect 479 102 513 136
rect -255 0 -221 34
rect -185 0 -151 34
rect -115 0 -81 34
rect -45 0 -11 34
rect 25 0 59 34
rect 95 0 129 34
rect 165 0 199 34
rect 235 0 269 34
rect 305 0 339 34
rect 375 0 409 34
rect 445 0 479 34
<< poly >>
rect -14 2422 166 2438
rect -14 2388 2 2422
rect 36 2388 116 2422
rect 150 2388 166 2422
rect -14 2372 166 2388
rect -14 304 166 320
rect -14 270 2 304
rect 36 270 116 304
rect 150 270 166 304
rect -14 254 166 270
<< polycont >>
rect 2 2388 36 2422
rect 116 2388 150 2422
rect 2 270 36 304
rect 116 270 150 304
<< locali >>
rect -361 2656 -337 2690
rect -303 2656 -266 2690
rect -232 2656 -229 2690
rect -161 2656 -146 2690
rect -90 2656 -63 2690
rect -19 2656 18 2690
rect 55 2656 89 2690
rect 123 2656 160 2690
rect 194 2656 231 2690
rect 265 2656 302 2690
rect 336 2656 373 2690
rect 407 2656 530 2690
rect -361 2652 -327 2656
rect -361 2578 -327 2618
rect -361 2504 -327 2526
rect 513 2622 530 2656
rect 479 2616 530 2622
rect 479 2587 513 2616
rect 479 2518 513 2553
rect -361 2430 -327 2457
rect -361 2356 -327 2388
rect -361 2284 -327 2319
rect -361 2215 -327 2248
rect -361 2146 -327 2174
rect -361 2077 -327 2100
rect -361 2008 -327 2026
rect -361 1939 -327 1952
rect -361 1870 -327 1878
rect -361 1801 -327 1804
rect -361 1764 -327 1767
rect -361 1690 -327 1698
rect -361 1616 -327 1629
rect -361 1542 -327 1560
rect -361 1468 -327 1491
rect -361 1394 -327 1422
rect -361 1320 -327 1353
rect -361 1249 -327 1284
rect -361 1180 -327 1212
rect -361 1111 -327 1138
rect -361 1042 -327 1064
rect -361 973 -327 990
rect -361 904 -327 916
rect -361 835 -327 842
rect -361 766 -327 769
rect -361 730 -327 732
rect -361 657 -327 663
rect -361 584 -327 594
rect -361 511 -327 524
rect -361 438 -327 454
rect -361 365 -327 384
rect -361 292 -327 314
rect -361 219 -327 244
rect -117 2470 -82 2504
rect -48 2470 -13 2504
rect 21 2470 55 2504
rect 89 2470 123 2504
rect 157 2470 191 2504
rect 225 2470 327 2504
rect -175 2431 -141 2470
rect -175 2394 -141 2397
rect -14 2388 2 2422
rect 36 2388 116 2422
rect 176 2388 214 2422
rect 293 2400 327 2436
rect -175 2358 -141 2360
rect -175 2285 -141 2292
rect -175 2212 -141 2223
rect -175 2139 -141 2154
rect -175 2066 -141 2085
rect -175 1993 -141 2016
rect -175 1920 -141 1947
rect -175 1847 -141 1878
rect -175 1774 -141 1809
rect -175 1705 -141 1740
rect -175 1636 -141 1667
rect -175 1567 -141 1594
rect -175 1498 -141 1522
rect -175 1429 -141 1450
rect -175 1360 -141 1378
rect -175 1291 -141 1306
rect -175 1222 -141 1234
rect -175 1153 -141 1162
rect -175 1084 -141 1090
rect -175 1015 -141 1018
rect -175 980 -141 981
rect -175 908 -141 912
rect -175 836 -141 843
rect -175 764 -141 774
rect -175 692 -141 705
rect -175 620 -141 636
rect -175 548 -141 567
rect -175 476 -141 498
rect -175 404 -141 429
rect -175 332 -141 360
rect 9 304 143 2388
rect 293 2330 327 2366
rect 293 2260 327 2296
rect 293 2190 327 2226
rect 293 2147 327 2156
rect 293 2075 327 2086
rect 293 2003 327 2017
rect 293 1931 327 1948
rect 293 1859 327 1879
rect 293 1787 327 1810
rect 293 1715 327 1741
rect 293 1643 327 1672
rect 293 1571 327 1603
rect 293 1499 327 1534
rect 293 1430 327 1465
rect 293 1361 327 1393
rect 293 1292 327 1321
rect 293 1223 327 1248
rect 293 1154 327 1175
rect 293 1085 327 1102
rect 293 1016 327 1029
rect 293 947 327 956
rect 293 878 327 883
rect 293 809 327 810
rect 293 771 327 775
rect 293 698 327 706
rect 293 625 327 637
rect 293 552 327 568
rect 293 479 327 499
rect 293 406 327 430
rect 293 333 327 361
rect -175 256 -141 291
rect -14 270 2 304
rect 36 270 116 304
rect 150 270 166 304
rect 293 260 327 292
rect -175 188 -137 222
rect -103 188 -59 222
rect -19 188 19 222
rect 59 188 96 222
rect 137 188 173 222
rect 215 188 259 222
rect 293 188 327 226
rect 479 2449 513 2484
rect 479 2380 513 2415
rect 479 2312 513 2346
rect 513 2246 530 2292
rect 479 2244 530 2246
rect 513 2210 530 2244
rect 479 2207 530 2210
rect 513 2142 530 2207
rect 479 2134 530 2142
rect 513 2074 530 2134
rect 479 2061 530 2074
rect 513 2006 530 2061
rect 479 1988 530 2006
rect 513 1938 530 1988
rect 479 1915 530 1938
rect 513 1870 530 1915
rect 479 1842 530 1870
rect 513 1802 530 1842
rect 479 1769 530 1802
rect 513 1734 530 1769
rect 479 1700 530 1734
rect 513 1662 530 1700
rect 479 1632 530 1662
rect 513 1589 530 1632
rect 479 1564 530 1589
rect 513 1516 530 1564
rect 479 1496 530 1516
rect 513 1443 530 1496
rect 479 1428 530 1443
rect 513 1370 530 1428
rect 479 1360 530 1370
rect 513 1296 530 1360
rect 479 1292 530 1296
rect 513 1258 530 1292
rect 479 1256 530 1258
rect 513 1190 530 1256
rect 479 1182 530 1190
rect 513 1122 530 1182
rect 479 1108 530 1122
rect 513 1054 530 1108
rect 479 1034 530 1054
rect 513 986 530 1034
rect 479 960 530 986
rect 513 918 530 960
rect 479 886 530 918
rect 513 850 530 886
rect 479 816 530 850
rect 513 778 530 816
rect 479 748 530 778
rect 513 704 530 748
rect 479 680 530 704
rect 513 630 530 680
rect 479 612 530 630
rect 513 556 530 612
rect 479 544 530 556
rect 513 482 530 544
rect 479 476 530 482
rect 513 374 530 476
rect 479 368 530 374
rect 513 306 530 368
rect 479 294 530 306
rect 2494 417 2687 430
rect 2528 383 2574 417
rect 2608 383 2653 417
rect 2494 345 2687 383
rect 2528 311 2574 345
rect 2608 311 2653 345
rect 2494 298 2687 311
rect 513 238 530 294
rect 479 220 530 238
rect -361 146 -327 174
rect -361 68 -327 104
rect 513 170 530 220
rect 479 146 530 170
rect 513 102 530 146
rect 479 72 530 102
rect 513 38 530 72
rect -361 0 -323 34
rect -289 0 -255 34
rect -213 0 -185 34
rect -137 0 -115 34
rect -61 0 -45 34
rect 15 0 25 34
rect 91 0 95 34
rect 129 0 133 34
rect 199 0 209 34
rect 269 0 285 34
rect 339 0 361 34
rect 409 0 445 34
rect 479 0 530 38
<< viali >>
rect -229 2656 -195 2690
rect -146 2656 -124 2690
rect -124 2656 -112 2690
rect -63 2656 -53 2690
rect -53 2656 -29 2690
rect 21 2656 52 2690
rect 52 2656 55 2690
rect -361 2618 -327 2652
rect -361 2560 -327 2578
rect -361 2544 -327 2560
rect -361 2491 -327 2504
rect -361 2470 -327 2491
rect -361 2422 -327 2430
rect -361 2396 -327 2422
rect -361 2353 -327 2356
rect -361 2322 -327 2353
rect -361 2250 -327 2282
rect -361 2248 -327 2250
rect -361 2181 -327 2208
rect -361 2174 -327 2181
rect -361 2112 -327 2134
rect -361 2100 -327 2112
rect -361 2043 -327 2060
rect -361 2026 -327 2043
rect -361 1974 -327 1986
rect -361 1952 -327 1974
rect -361 1905 -327 1912
rect -361 1878 -327 1905
rect -361 1836 -327 1838
rect -361 1804 -327 1836
rect -361 1732 -327 1764
rect -361 1730 -327 1732
rect -361 1663 -327 1690
rect -361 1656 -327 1663
rect -361 1594 -327 1616
rect -361 1582 -327 1594
rect -361 1525 -327 1542
rect -361 1508 -327 1525
rect -361 1456 -327 1468
rect -361 1434 -327 1456
rect -361 1387 -327 1394
rect -361 1360 -327 1387
rect -361 1318 -327 1320
rect -361 1286 -327 1318
rect -361 1215 -327 1246
rect -361 1212 -327 1215
rect -361 1146 -327 1172
rect -361 1138 -327 1146
rect -361 1077 -327 1098
rect -361 1064 -327 1077
rect -361 1008 -327 1024
rect -361 990 -327 1008
rect -361 939 -327 950
rect -361 916 -327 939
rect -361 870 -327 876
rect -361 842 -327 870
rect -361 801 -327 803
rect -361 769 -327 801
rect -361 697 -327 730
rect -361 696 -327 697
rect -361 628 -327 657
rect -361 623 -327 628
rect -361 558 -327 584
rect -361 550 -327 558
rect -361 488 -327 511
rect -361 477 -327 488
rect -361 418 -327 438
rect -361 404 -327 418
rect -361 348 -327 365
rect -361 331 -327 348
rect -361 278 -327 292
rect -361 258 -327 278
rect -361 208 -327 219
rect -361 185 -327 208
rect -175 2470 -151 2504
rect -151 2470 -141 2504
rect -175 2397 -141 2431
rect 142 2388 150 2422
rect 150 2388 176 2422
rect 214 2388 248 2422
rect -175 2326 -141 2358
rect -175 2324 -141 2326
rect -175 2257 -141 2285
rect -175 2251 -141 2257
rect -175 2188 -141 2212
rect -175 2178 -141 2188
rect -175 2119 -141 2139
rect -175 2105 -141 2119
rect -175 2050 -141 2066
rect -175 2032 -141 2050
rect -175 1981 -141 1993
rect -175 1959 -141 1981
rect -175 1912 -141 1920
rect -175 1886 -141 1912
rect -175 1843 -141 1847
rect -175 1813 -141 1843
rect -175 1740 -141 1774
rect -175 1671 -141 1701
rect -175 1667 -141 1671
rect -175 1602 -141 1628
rect -175 1594 -141 1602
rect -175 1533 -141 1556
rect -175 1522 -141 1533
rect -175 1464 -141 1484
rect -175 1450 -141 1464
rect -175 1395 -141 1412
rect -175 1378 -141 1395
rect -175 1326 -141 1340
rect -175 1306 -141 1326
rect -175 1257 -141 1268
rect -175 1234 -141 1257
rect -175 1188 -141 1196
rect -175 1162 -141 1188
rect -175 1119 -141 1124
rect -175 1090 -141 1119
rect -175 1050 -141 1052
rect -175 1018 -141 1050
rect -175 946 -141 980
rect -175 877 -141 908
rect -175 874 -141 877
rect -175 808 -141 836
rect -175 802 -141 808
rect -175 739 -141 764
rect -175 730 -141 739
rect -175 670 -141 692
rect -175 658 -141 670
rect -175 601 -141 620
rect -175 586 -141 601
rect -175 532 -141 548
rect -175 514 -141 532
rect -175 463 -141 476
rect -175 442 -141 463
rect -175 394 -141 404
rect -175 370 -141 394
rect -175 325 -141 332
rect -175 298 -141 325
rect 293 2120 327 2147
rect 293 2113 327 2120
rect 293 2051 327 2075
rect 293 2041 327 2051
rect 293 1982 327 2003
rect 293 1969 327 1982
rect 293 1913 327 1931
rect 293 1897 327 1913
rect 293 1844 327 1859
rect 293 1825 327 1844
rect 293 1775 327 1787
rect 293 1753 327 1775
rect 293 1706 327 1715
rect 293 1681 327 1706
rect 293 1637 327 1643
rect 293 1609 327 1637
rect 293 1568 327 1571
rect 293 1537 327 1568
rect 293 1465 327 1499
rect 293 1396 327 1427
rect 293 1393 327 1396
rect 293 1327 327 1355
rect 293 1321 327 1327
rect 293 1258 327 1282
rect 293 1248 327 1258
rect 293 1189 327 1209
rect 293 1175 327 1189
rect 293 1120 327 1136
rect 293 1102 327 1120
rect 293 1051 327 1063
rect 293 1029 327 1051
rect 293 982 327 990
rect 293 956 327 982
rect 293 913 327 917
rect 293 883 327 913
rect 293 810 327 844
rect 293 740 327 771
rect 293 737 327 740
rect 293 671 327 698
rect 293 664 327 671
rect 293 602 327 625
rect 293 591 327 602
rect 293 533 327 552
rect 293 518 327 533
rect 293 464 327 479
rect 293 445 327 464
rect 293 395 327 406
rect 293 372 327 395
rect 293 326 327 333
rect 293 299 327 326
rect 293 226 327 260
rect -137 188 -103 222
rect -59 188 -53 222
rect -53 188 -25 222
rect 19 188 25 222
rect 25 188 53 222
rect 96 188 103 222
rect 103 188 130 222
rect 173 188 181 222
rect 181 188 207 222
rect 479 2278 513 2280
rect 479 2246 513 2278
rect 479 2176 513 2207
rect 479 2173 513 2176
rect 479 2108 513 2134
rect 479 2100 513 2108
rect 479 2040 513 2061
rect 479 2027 513 2040
rect 479 1972 513 1988
rect 479 1954 513 1972
rect 479 1904 513 1915
rect 479 1881 513 1904
rect 479 1836 513 1842
rect 479 1808 513 1836
rect 479 1768 513 1769
rect 479 1735 513 1768
rect 479 1666 513 1696
rect 479 1662 513 1666
rect 479 1598 513 1623
rect 479 1589 513 1598
rect 479 1530 513 1550
rect 479 1516 513 1530
rect 479 1462 513 1477
rect 479 1443 513 1462
rect 479 1394 513 1404
rect 479 1370 513 1394
rect 479 1326 513 1330
rect 479 1296 513 1326
rect 479 1224 513 1256
rect 479 1222 513 1224
rect 479 1156 513 1182
rect 479 1148 513 1156
rect 479 1088 513 1108
rect 479 1074 513 1088
rect 479 1020 513 1034
rect 479 1000 513 1020
rect 479 952 513 960
rect 479 926 513 952
rect 479 884 513 886
rect 479 852 513 884
rect 479 782 513 812
rect 479 778 513 782
rect 479 714 513 738
rect 479 704 513 714
rect 479 646 513 664
rect 479 630 513 646
rect 479 578 513 590
rect 479 556 513 578
rect 479 510 513 516
rect 479 482 513 510
rect 479 408 513 442
rect 479 340 513 368
rect 479 334 513 340
rect 2494 383 2528 417
rect 2574 383 2608 417
rect 2653 383 2687 417
rect 2494 311 2528 345
rect 2574 311 2608 345
rect 2653 311 2687 345
rect 479 272 513 294
rect 479 260 513 272
rect 479 204 513 220
rect -361 138 -327 146
rect -361 112 -327 138
rect 479 186 513 204
rect 479 136 513 146
rect 479 112 513 136
rect 479 38 513 72
rect -323 0 -289 34
rect -247 0 -221 34
rect -221 0 -213 34
rect -171 0 -151 34
rect -151 0 -137 34
rect -95 0 -81 34
rect -81 0 -61 34
rect -19 0 -11 34
rect -11 0 15 34
rect 57 0 59 34
rect 59 0 91 34
rect 133 0 165 34
rect 165 0 167 34
rect 209 0 235 34
rect 235 0 243 34
rect 285 0 305 34
rect 305 0 319 34
rect 361 0 375 34
rect 375 0 395 34
<< metal1 >>
tri 17 5162 145 5290 se
rect 145 5170 573 5290
rect 145 5162 419 5170
tri 419 5162 427 5170 nw
tri 521 5162 529 5170 ne
rect 529 5162 573 5170
tri 573 5162 701 5290 sw
tri 0 5145 17 5162 se
rect 17 5145 402 5162
tri 402 5145 419 5162 nw
tri 529 5145 546 5162 ne
rect 546 5145 2556 5162
tri 546 5118 573 5145 ne
rect 573 5118 2556 5145
tri 573 5045 646 5118 ne
rect 646 5045 2556 5118
rect 2538 4903 2654 4909
tri 1894 4836 1919 4861 ne
tri 1919 4836 1944 4861 nw
rect 2590 4851 2602 4903
rect 2538 4836 2654 4851
rect 1861 4823 1977 4829
rect 1913 4771 1925 4823
rect 1861 4758 1977 4771
rect 1913 4706 1925 4758
rect 1861 4693 1977 4706
rect 1913 4641 1925 4693
rect 1861 4628 1977 4641
rect 1913 4576 1925 4628
rect 2590 4784 2602 4836
rect 2538 4769 2654 4784
rect 2590 4717 2602 4769
rect 2538 4702 2654 4717
rect 2590 4650 2602 4702
rect 2538 4636 2654 4650
rect 1861 4563 1977 4576
rect 820 4549 997 4550
rect 820 4545 1048 4549
rect 820 4493 828 4545
rect 880 4493 909 4545
rect 961 4493 990 4545
rect 1042 4493 1048 4545
rect 820 4481 1048 4493
rect 820 4429 828 4481
rect 880 4429 909 4481
rect 961 4429 990 4481
rect 1042 4429 1048 4481
rect 820 4425 1048 4429
rect 1581 4544 1697 4550
rect 1633 4492 1645 4544
rect 1581 4478 1697 4492
rect 1633 4426 1645 4478
rect 820 4415 997 4425
tri 1164 4415 1167 4418 se
rect 820 4409 999 4415
rect 820 4357 947 4409
tri 1142 4393 1164 4415 se
rect 1164 4393 1167 4415
rect 1581 4412 1697 4426
rect 820 4345 999 4357
rect 820 4293 947 4345
rect 1065 4341 1071 4393
rect 1123 4341 1192 4393
rect 1244 4341 1250 4393
rect 1633 4360 1645 4412
rect 1581 4346 1697 4360
rect 820 4285 999 4293
rect 1424 4294 1476 4300
rect 820 4073 997 4285
rect 1424 4229 1476 4242
rect 1424 4164 1476 4177
rect 1424 4099 1476 4112
rect 820 4067 1000 4073
rect 872 4015 884 4067
rect 936 4015 948 4067
rect 820 4001 1000 4015
rect 542 3995 658 4001
rect 594 3943 606 3995
rect 542 3928 658 3943
rect 594 3876 606 3928
rect 542 3862 658 3876
rect 594 3810 606 3862
rect 542 3796 658 3810
rect 594 3744 606 3796
rect 542 3730 658 3744
rect 594 3678 606 3730
rect 542 3664 658 3678
rect 594 3612 606 3664
rect 542 3598 658 3612
rect 594 3546 606 3598
rect 542 3532 658 3546
rect 594 3480 606 3532
rect 542 3466 658 3480
rect 594 3414 606 3466
rect 542 3400 658 3414
rect 594 3348 606 3400
rect 542 3334 658 3348
rect 594 3282 606 3334
rect 542 3268 658 3282
rect 594 3216 606 3268
rect 542 3202 658 3216
rect 594 3150 606 3202
rect 542 3136 658 3150
rect 594 3084 606 3136
rect 542 3070 658 3084
rect 594 3018 606 3070
rect 542 3004 658 3018
rect 594 2952 606 3004
rect 542 2938 658 2952
rect 594 2886 606 2938
tri 214 2850 239 2875 ne
tri 211 2725 239 2753 se
rect 239 2725 402 2875
rect 542 2872 658 2886
rect 594 2820 606 2872
rect 542 2806 658 2820
rect 594 2754 606 2806
rect 542 2740 658 2754
tri 182 2696 211 2725 se
rect 211 2696 402 2725
tri 402 2696 431 2725 sw
rect -367 2690 67 2696
rect -367 2656 -229 2690
rect -195 2656 -146 2690
rect -112 2656 -63 2690
rect -29 2656 21 2690
rect 55 2656 67 2690
rect -367 2652 67 2656
rect -367 2618 -361 2652
rect -327 2650 67 2652
tri 136 2650 182 2696 se
rect 182 2650 431 2696
tri 431 2650 477 2696 sw
rect 594 2688 606 2740
rect 542 2674 658 2688
rect -327 2618 -321 2650
tri -321 2625 -296 2650 nw
tri 119 2633 136 2650 se
rect 136 2633 477 2650
tri 477 2633 494 2650 sw
tri 111 2625 119 2633 se
rect 119 2625 494 2633
rect -367 2578 -321 2618
tri 103 2617 111 2625 se
rect 111 2617 494 2625
tri 98 2612 103 2617 se
rect 103 2613 494 2617
rect 594 2622 606 2674
rect 542 2616 658 2622
rect 872 3949 884 4001
rect 936 3949 948 4001
rect 820 3935 1000 3949
rect 872 3883 884 3935
rect 936 3883 948 3935
rect 820 3869 1000 3883
rect 872 3817 884 3869
rect 936 3817 948 3869
rect 820 3803 1000 3817
rect 872 3751 884 3803
rect 936 3751 948 3803
rect 820 3737 1000 3751
rect 872 3685 884 3737
rect 936 3685 948 3737
rect 820 3671 1000 3685
rect 872 3619 884 3671
rect 936 3619 948 3671
rect 820 3605 1000 3619
rect 872 3553 884 3605
rect 936 3553 948 3605
rect 820 3539 1000 3553
rect 872 3487 884 3539
rect 936 3487 948 3539
rect 820 3474 1000 3487
rect 872 3422 884 3474
rect 936 3422 948 3474
rect 820 3409 1000 3422
rect 872 3357 884 3409
rect 936 3357 948 3409
rect 820 3344 1000 3357
rect 872 3292 884 3344
rect 936 3292 948 3344
rect 820 3279 1000 3292
rect 872 3227 884 3279
rect 936 3227 948 3279
rect 820 3214 1000 3227
rect 872 3162 884 3214
rect 936 3162 948 3214
rect 820 3149 1000 3162
rect 872 3097 884 3149
rect 936 3097 948 3149
rect 820 3084 1000 3097
rect 872 3032 884 3084
rect 936 3032 948 3084
rect 820 3019 1000 3032
rect 872 2967 884 3019
rect 936 2967 948 3019
rect 820 2954 1000 2967
rect 872 2902 884 2954
rect 936 2902 948 2954
rect 820 2889 1000 2902
rect 872 2837 884 2889
rect 936 2837 948 2889
rect 820 2824 1000 2837
rect 872 2772 884 2824
rect 936 2772 948 2824
rect 820 2759 1000 2772
rect 872 2707 884 2759
rect 936 2707 948 2759
rect 820 2694 1000 2707
rect 872 2642 884 2694
rect 936 2642 948 2694
rect 820 2636 1000 2642
rect 1424 4034 1476 4047
rect 1424 3969 1476 3982
rect 1424 3904 1476 3917
rect 1424 3839 1476 3852
rect 1424 3774 1476 3787
rect 1424 3709 1476 3722
rect 1424 3644 1476 3657
rect 1424 3579 1476 3592
rect 1424 3514 1476 3527
rect 1424 3449 1476 3462
rect 1424 3384 1476 3397
rect 1424 3319 1476 3332
rect 1424 3254 1476 3267
rect 1424 3189 1476 3202
rect 1424 3124 1476 3137
rect 1424 3059 1476 3072
rect 1424 2995 1476 3007
rect 1424 2931 1476 2943
rect 1633 4294 1645 4346
rect 1581 4280 1697 4294
rect 1633 4228 1645 4280
rect 1581 4214 1697 4228
rect 1633 4162 1645 4214
rect 1581 4148 1697 4162
rect 1633 4096 1645 4148
rect 1581 4082 1697 4096
rect 1633 4030 1645 4082
rect 1581 4016 1697 4030
rect 1633 3964 1645 4016
rect 1581 3950 1697 3964
rect 1633 3898 1645 3950
rect 1581 3884 1697 3898
rect 1633 3832 1645 3884
rect 1581 3818 1697 3832
rect 1633 3766 1645 3818
rect 1581 3752 1697 3766
rect 1633 3700 1645 3752
rect 1581 3686 1697 3700
rect 1633 3634 1645 3686
rect 1581 3620 1697 3634
rect 1633 3568 1645 3620
rect 1581 3555 1697 3568
rect 1633 3503 1645 3555
rect 1581 3490 1697 3503
rect 1633 3438 1645 3490
rect 1581 3425 1697 3438
rect 1633 3373 1645 3425
rect 1581 3360 1697 3373
rect 1633 3308 1645 3360
rect 1581 3295 1697 3308
rect 1633 3243 1645 3295
rect 1581 3230 1697 3243
rect 1633 3178 1645 3230
rect 1581 3165 1697 3178
rect 1633 3113 1645 3165
rect 1581 3100 1697 3113
rect 1633 3048 1645 3100
rect 1581 3035 1697 3048
rect 1633 2983 1645 3035
rect 1581 2970 1697 2983
rect 1633 2918 1645 2970
rect 1581 2912 1697 2918
rect 1913 4511 1925 4563
tri 2172 4550 2217 4595 se
rect 2217 4550 2236 4595
tri 2164 4542 2172 4550 se
rect 2172 4543 2236 4550
rect 2288 4543 2330 4595
rect 2382 4543 2388 4595
rect 2172 4542 2388 4543
rect 1861 4498 1977 4511
rect 1913 4446 1925 4498
rect 1861 4433 1977 4446
rect 1913 4381 1925 4433
rect 1861 4368 1977 4381
rect 1913 4316 1925 4368
rect 1861 4303 1977 4316
rect 1913 4251 1925 4303
rect 1861 4238 1977 4251
rect 1913 4186 1925 4238
rect 1861 4173 1977 4186
rect 1913 4121 1925 4173
rect 1861 4108 1977 4121
rect 1913 4056 1925 4108
rect 1861 4043 1977 4056
rect 1913 3991 1925 4043
rect 1861 3978 1977 3991
rect 1913 3926 1925 3978
rect 1861 3913 1977 3926
rect 1913 3861 1925 3913
rect 1861 3848 1977 3861
rect 1913 3796 1925 3848
rect 1861 3783 1977 3796
rect 1913 3731 1925 3783
rect 1861 3718 1977 3731
rect 1913 3666 1925 3718
rect 1861 3653 1977 3666
rect 1913 3601 1925 3653
rect 1861 3588 1977 3601
rect 1913 3536 1925 3588
rect 1861 3523 1977 3536
rect 1913 3471 1925 3523
rect 1861 3458 1977 3471
rect 1913 3406 1925 3458
rect 1861 3393 1977 3406
rect 1913 3341 1925 3393
rect 1861 3328 1977 3341
rect 1913 3276 1925 3328
rect 1861 3263 1977 3276
rect 1913 3211 1925 3263
rect 1861 3198 1977 3211
rect 1913 3146 1925 3198
rect 1861 3133 1977 3146
rect 1913 3081 1925 3133
rect 1861 3068 1977 3081
rect 1424 2867 1476 2879
rect 1424 2803 1476 2815
rect 1424 2739 1476 2751
rect 2205 4531 2388 4542
rect 2205 4520 2311 4531
rect 2205 4490 2217 4520
rect 2153 4476 2217 4490
rect 2205 4468 2217 4476
rect 2269 4479 2311 4520
rect 2363 4479 2388 4531
rect 2590 4584 2602 4636
rect 2538 4570 2654 4584
rect 3180 4763 3296 4769
rect 3232 4711 3244 4763
rect 3180 4697 3296 4711
rect 3232 4645 3244 4697
rect 3180 4631 3296 4645
rect 3232 4579 3244 4631
rect 2590 4518 2602 4570
rect 2538 4504 2654 4518
rect 2205 4455 2269 4468
rect 2205 4424 2217 4455
rect 2153 4410 2217 4424
rect 2205 4403 2217 4410
rect 2205 4390 2269 4403
rect 2205 4358 2217 4390
rect 2153 4344 2217 4358
rect 2205 4338 2217 4344
rect 2590 4452 2602 4504
rect 2538 4438 2654 4452
rect 2590 4386 2602 4438
rect 2876 4565 2992 4571
rect 2928 4513 2940 4565
rect 2876 4500 2992 4513
rect 2928 4448 2940 4500
rect 2876 4435 2992 4448
rect 2538 4380 2654 4386
tri 2671 4380 2688 4397 sw
rect 2928 4383 2940 4435
rect 2671 4372 2688 4380
tri 2688 4372 2696 4380 sw
rect 2671 4365 2802 4372
rect 2589 4359 2802 4365
rect 2205 4325 2269 4338
rect 2205 4292 2217 4325
rect 2153 4278 2217 4292
rect 2205 4273 2217 4278
tri 2564 4316 2589 4341 ne
rect 2205 4260 2269 4273
rect 2205 4226 2217 4260
rect 2153 4212 2217 4226
rect 2205 4208 2217 4212
rect 2205 4195 2269 4208
rect 2205 4160 2217 4195
rect 2153 4146 2217 4160
rect 2205 4143 2217 4146
rect 2205 4130 2269 4143
rect 2205 4094 2217 4130
rect 2153 4080 2217 4094
rect 2205 4078 2217 4080
rect 2205 4065 2269 4078
rect 2205 4028 2217 4065
rect 2153 4014 2217 4028
rect 2205 4013 2217 4014
rect 2205 4000 2269 4013
rect 2205 3962 2217 4000
rect 2153 3948 2217 3962
rect 2205 3935 2269 3948
rect 2205 3896 2217 3935
rect 2153 3883 2217 3896
rect 2153 3882 2269 3883
rect 2205 3870 2269 3882
rect 2205 3830 2217 3870
rect 2153 3818 2217 3830
rect 2153 3816 2269 3818
rect 2205 3805 2269 3816
rect 2205 3764 2217 3805
rect 2153 3753 2217 3764
rect 2153 3750 2269 3753
rect 2205 3740 2269 3750
rect 2205 3698 2217 3740
rect 2153 3688 2217 3698
rect 2153 3685 2269 3688
rect 2205 3675 2269 3685
rect 2205 3633 2217 3675
rect 2153 3623 2217 3633
rect 2153 3620 2269 3623
rect 2205 3610 2269 3620
rect 2205 3568 2217 3610
rect 2153 3558 2217 3568
rect 2153 3555 2269 3558
rect 2205 3546 2269 3555
rect 2205 3503 2217 3546
rect 2153 3494 2217 3503
rect 2153 3490 2269 3494
rect 2205 3482 2269 3490
rect 2205 3438 2217 3482
rect 2153 3430 2217 3438
rect 2153 3425 2269 3430
rect 2205 3418 2269 3425
rect 2205 3373 2217 3418
rect 2153 3366 2217 3373
rect 2153 3360 2269 3366
rect 2205 3354 2269 3360
rect 2205 3308 2217 3354
rect 2153 3302 2217 3308
rect 2153 3295 2269 3302
rect 2205 3290 2269 3295
rect 2205 3243 2217 3290
rect 2153 3238 2217 3243
rect 2153 3230 2269 3238
rect 2205 3226 2269 3230
rect 2205 3178 2217 3226
rect 2153 3174 2217 3178
rect 2153 3165 2269 3174
rect 2205 3162 2269 3165
rect 2205 3113 2217 3162
rect 2153 3110 2217 3113
rect 2153 3100 2269 3110
rect 2205 3098 2269 3100
rect 2205 3048 2217 3098
rect 2153 3046 2217 3048
rect 2153 3035 2269 3046
rect 2205 3034 2269 3035
rect 2205 2983 2217 3034
rect 2153 2982 2217 2983
rect 2153 2970 2269 2982
rect 2205 2918 2217 2970
rect 2153 2912 2269 2918
rect 2641 4307 2653 4359
rect 2705 4307 2717 4359
rect 2769 4307 2802 4359
rect 2589 4294 2802 4307
rect 2641 4242 2653 4294
rect 2705 4242 2717 4294
rect 2769 4259 2802 4294
rect 2876 4370 2992 4383
rect 2928 4318 2940 4370
rect 2876 4305 2992 4318
rect 2589 4229 2769 4242
rect 2641 4177 2653 4229
rect 2705 4177 2717 4229
rect 2589 4164 2769 4177
rect 2641 4112 2653 4164
rect 2705 4112 2717 4164
rect 2589 4099 2769 4112
rect 2641 4047 2653 4099
rect 2705 4047 2717 4099
rect 2589 4034 2769 4047
rect 2641 3982 2653 4034
rect 2705 3982 2717 4034
rect 2589 3969 2769 3982
rect 2641 3917 2653 3969
rect 2705 3917 2717 3969
rect 2589 3904 2769 3917
rect 2641 3852 2653 3904
rect 2705 3852 2717 3904
rect 2589 3839 2769 3852
rect 2641 3787 2653 3839
rect 2705 3787 2717 3839
rect 2589 3774 2769 3787
rect 2641 3722 2653 3774
rect 2705 3722 2717 3774
rect 2589 3709 2769 3722
rect 2641 3657 2653 3709
rect 2705 3657 2717 3709
rect 2589 3644 2769 3657
rect 2641 3592 2653 3644
rect 2705 3592 2717 3644
rect 2589 3579 2769 3592
rect 2641 3527 2653 3579
rect 2705 3527 2717 3579
rect 2589 3514 2769 3527
rect 2641 3462 2653 3514
rect 2705 3462 2717 3514
rect 2589 3449 2769 3462
rect 2641 3397 2653 3449
rect 2705 3397 2717 3449
rect 2589 3384 2769 3397
rect 2641 3332 2653 3384
rect 2705 3332 2717 3384
rect 2589 3319 2769 3332
rect 2641 3267 2653 3319
rect 2705 3267 2717 3319
rect 2589 3254 2769 3267
rect 2641 3202 2653 3254
rect 2705 3202 2717 3254
rect 2589 3189 2769 3202
rect 2641 3137 2653 3189
rect 2705 3137 2717 3189
rect 2589 3124 2769 3137
rect 2641 3072 2653 3124
rect 2705 3072 2717 3124
rect 2589 3059 2769 3072
rect 2641 3007 2653 3059
rect 2705 3007 2717 3059
rect 2589 2994 2769 3007
rect 1861 2690 1977 2696
rect 1424 2675 1476 2687
rect 820 2616 997 2636
tri 1894 2663 1919 2688 se
tri 1919 2663 1944 2688 sw
rect 1424 2617 1476 2623
rect 2928 4253 2940 4305
rect 2876 4240 2992 4253
rect 2928 4188 2940 4240
rect 2876 4175 2992 4188
rect 2928 4123 2940 4175
rect 2876 4110 2992 4123
rect 2928 4058 2940 4110
rect 2876 4045 2992 4058
rect 2928 3993 2940 4045
rect 2876 3980 2992 3993
rect 2928 3928 2940 3980
rect 2876 3915 2992 3928
rect 2928 3863 2940 3915
rect 2876 3850 2992 3863
rect 2928 3798 2940 3850
rect 2876 3785 2992 3798
rect 2928 3733 2940 3785
rect 2876 3720 2992 3733
rect 2928 3668 2940 3720
rect 2876 3655 2992 3668
rect 2928 3603 2940 3655
rect 2876 3590 2992 3603
rect 2928 3538 2940 3590
rect 2876 3525 2992 3538
rect 2928 3473 2940 3525
rect 2876 3460 2992 3473
rect 2928 3408 2940 3460
rect 2876 3395 2992 3408
rect 2928 3343 2940 3395
rect 2876 3330 2992 3343
rect 2876 2632 2992 2638
rect 3180 4565 3296 4579
rect 3232 4513 3244 4565
rect 3180 4499 3296 4513
rect 3232 4447 3244 4499
rect 3180 4434 3296 4447
rect 3232 4382 3244 4434
rect 3180 4369 3296 4382
rect 3232 4317 3244 4369
rect 3180 4304 3296 4317
rect 3232 4252 3244 4304
rect 3180 4239 3296 4252
rect 3232 4187 3244 4239
rect 3180 4174 3296 4187
rect 3232 4122 3244 4174
rect 3180 4109 3296 4122
rect 3232 4057 3244 4109
rect 3180 4044 3296 4057
rect 3232 3992 3244 4044
rect 3180 3979 3296 3992
rect 3232 3927 3244 3979
rect 3180 3914 3296 3927
rect 3232 3862 3244 3914
rect 3180 3849 3296 3862
rect 3232 3797 3244 3849
rect 3180 3784 3296 3797
rect 3232 3732 3244 3784
rect 3180 3719 3296 3732
rect 3232 3667 3244 3719
rect 3180 3654 3296 3667
rect 3232 3602 3244 3654
rect 3180 3589 3296 3602
rect 3232 3537 3244 3589
rect 3180 3524 3296 3537
rect 3232 3472 3244 3524
rect 3180 3459 3296 3472
rect 3232 3407 3244 3459
rect 3180 3394 3296 3407
rect 3232 3342 3244 3394
rect 3180 3329 3296 3342
rect 3232 3277 3244 3329
rect 3180 3264 3296 3277
rect 3232 3212 3244 3264
rect 3180 3199 3296 3212
rect 3232 3147 3244 3199
rect 3180 3134 3296 3147
rect 3232 3082 3244 3134
rect 3180 3069 3296 3082
rect 3232 3017 3244 3069
rect 3180 3004 3296 3017
rect 3232 2952 3244 3004
rect 3180 2939 3296 2952
rect 3232 2887 3244 2939
rect 3180 2874 3296 2887
rect 3232 2822 3244 2874
rect 3180 2809 3296 2822
rect 3232 2757 3244 2809
rect 3180 2744 3296 2757
rect 3232 2692 3244 2744
rect 3180 2679 3296 2692
rect 103 2612 268 2613
tri 268 2612 269 2613 nw
tri 345 2612 346 2613 ne
rect 346 2612 494 2613
rect 1036 2613 1236 2617
tri 1236 2613 1240 2617 sw
rect 2589 2616 2769 2622
rect 3232 2627 3244 2679
rect 3180 2621 3296 2627
tri 73 2587 98 2612 se
rect 98 2587 243 2612
tri 243 2587 268 2612 nw
tri 346 2587 371 2612 ne
rect 371 2588 494 2612
tri 494 2588 518 2612 sw
tri 1012 2588 1036 2612 se
rect 1036 2588 1240 2613
tri 1240 2588 1265 2613 sw
tri 2318 2588 2343 2613 se
rect 2343 2588 2543 2616
rect 371 2587 518 2588
tri 518 2587 519 2588 sw
tri 1011 2587 1012 2588 se
rect 1012 2587 2543 2588
tri 71 2585 73 2587 se
rect 73 2585 241 2587
tri 241 2585 243 2587 nw
tri 371 2585 373 2587 ne
rect 373 2585 2543 2587
tri 69 2583 71 2585 se
rect 71 2583 239 2585
tri 239 2583 241 2585 nw
tri 279 2583 281 2585 se
rect 281 2583 333 2585
tri 373 2583 375 2585 ne
rect -367 2544 -361 2578
rect -327 2544 -321 2578
rect -367 2504 -321 2544
tri 2 2516 69 2583 se
rect 69 2543 199 2583
tri 199 2543 239 2583 nw
tri 239 2543 279 2583 se
rect 279 2579 333 2583
rect 279 2543 281 2579
rect 69 2516 172 2543
tri 172 2516 199 2543 nw
tri 212 2516 239 2543 se
rect 239 2527 281 2543
rect 239 2516 333 2527
rect -367 2470 -361 2504
rect -327 2470 -321 2504
rect -367 2430 -321 2470
rect -367 2396 -361 2430
rect -327 2396 -321 2430
rect -367 2356 -321 2396
rect -367 2322 -361 2356
rect -327 2322 -321 2356
rect -367 2282 -321 2322
rect -367 2248 -361 2282
rect -327 2248 -321 2282
rect -367 2208 -321 2248
rect -367 2174 -361 2208
rect -327 2174 -321 2208
rect -367 2134 -321 2174
rect -367 2100 -361 2134
rect -327 2100 -321 2134
rect -367 2060 -321 2100
rect -367 2026 -361 2060
rect -327 2026 -321 2060
rect -367 1986 -321 2026
rect -367 1952 -361 1986
rect -327 1952 -321 1986
rect -367 1912 -321 1952
rect -367 1878 -361 1912
rect -327 1878 -321 1912
rect -367 1838 -321 1878
rect -367 1804 -361 1838
rect -327 1804 -321 1838
rect -367 1764 -321 1804
rect -367 1730 -361 1764
rect -327 1730 -321 1764
rect -367 1690 -321 1730
rect -367 1656 -361 1690
rect -327 1656 -321 1690
rect -367 1616 -321 1656
rect -367 1582 -361 1616
rect -327 1582 -321 1616
rect -367 1542 -321 1582
rect -367 1508 -361 1542
rect -327 1508 -321 1542
rect -367 1468 -321 1508
rect -367 1434 -361 1468
rect -327 1434 -321 1468
rect -367 1394 -321 1434
rect -367 1360 -361 1394
rect -327 1360 -321 1394
rect -367 1320 -321 1360
rect -367 1286 -361 1320
rect -327 1286 -321 1320
rect -367 1246 -321 1286
rect -367 1212 -361 1246
rect -327 1212 -321 1246
rect -367 1172 -321 1212
rect -367 1138 -361 1172
rect -327 1138 -321 1172
rect -367 1098 -321 1138
rect -367 1064 -361 1098
rect -327 1064 -321 1098
rect -367 1024 -321 1064
rect -367 990 -361 1024
rect -327 990 -321 1024
rect -367 950 -321 990
rect -367 916 -361 950
rect -327 916 -321 950
rect -367 876 -321 916
rect -367 842 -361 876
rect -327 842 -321 876
rect -367 803 -321 842
rect -367 769 -361 803
rect -327 769 -321 803
rect -367 730 -321 769
rect -367 696 -361 730
rect -327 696 -321 730
rect -367 657 -321 696
rect -367 623 -361 657
rect -327 623 -321 657
rect -367 584 -321 623
rect -367 550 -361 584
rect -327 550 -321 584
rect -367 511 -321 550
rect -367 477 -361 511
rect -327 477 -321 511
rect -367 438 -321 477
rect -367 404 -361 438
rect -327 404 -321 438
rect -367 365 -321 404
rect -367 331 -361 365
rect -327 331 -321 365
rect -367 292 -321 331
rect -367 258 -361 292
rect -327 258 -321 292
rect -367 219 -321 258
rect -367 185 -361 219
rect -327 185 -321 219
rect -367 146 -321 185
rect -181 2504 -135 2516
rect -181 2470 -175 2504
rect -141 2470 -135 2504
rect -181 2431 -135 2470
tri -74 2440 2 2516 se
rect 2 2480 136 2516
tri 136 2480 172 2516 nw
tri 176 2480 212 2516 se
rect 212 2513 333 2516
rect 212 2480 281 2513
rect 2 2440 96 2480
tri 96 2440 136 2480 nw
tri 136 2440 176 2480 se
rect 176 2461 281 2480
rect 375 2562 2543 2585
tri 375 2468 469 2562 ne
rect 469 2468 2543 2562
tri 2634 2468 2754 2588 se
rect 2754 2468 3479 2588
rect 176 2455 333 2461
rect 176 2440 318 2455
tri 318 2440 333 2455 nw
tri 2606 2440 2634 2468 se
rect 2634 2440 2822 2468
tri 2822 2440 2850 2468 nw
rect -181 2397 -175 2431
rect -141 2397 -135 2431
tri -86 2428 -74 2440 se
rect -74 2428 84 2440
tri 84 2428 96 2440 nw
tri 124 2428 136 2440 se
rect 136 2428 306 2440
tri 306 2428 318 2440 nw
tri 346 2428 358 2440 se
rect 358 2428 2703 2440
rect -181 2358 -135 2397
rect -181 2324 -175 2358
rect -141 2324 -135 2358
rect -181 2285 -135 2324
rect -181 2251 -175 2285
rect -141 2251 -135 2285
rect -181 2212 -135 2251
rect -181 2178 -175 2212
rect -141 2178 -135 2212
rect -181 2139 -135 2178
rect -181 2105 -175 2139
rect -141 2105 -135 2139
rect -181 2066 -135 2105
rect -181 2032 -175 2066
rect -141 2032 -135 2066
rect -181 1993 -135 2032
rect -181 1959 -175 1993
rect -141 1959 -135 1993
rect -181 1920 -135 1959
rect -181 1886 -175 1920
rect -141 1886 -135 1920
rect -181 1847 -135 1886
rect -181 1813 -175 1847
rect -141 1813 -135 1847
rect -181 1774 -135 1813
rect -181 1740 -175 1774
rect -141 1740 -135 1774
tri -87 2427 -86 2428 se
rect -86 2427 83 2428
tri 83 2427 84 2428 nw
tri 123 2427 124 2428 se
rect 124 2427 293 2428
rect -87 2422 78 2427
tri 78 2422 83 2427 nw
tri 118 2422 123 2427 se
rect 123 2422 293 2427
rect -87 2403 59 2422
tri 59 2403 78 2422 nw
tri 99 2403 118 2422 se
rect 118 2403 142 2422
rect -87 2388 44 2403
tri 44 2388 59 2403 nw
tri 84 2388 99 2403 se
rect 99 2388 142 2403
rect 176 2388 214 2422
rect 248 2415 293 2422
tri 293 2415 306 2428 nw
tri 333 2415 346 2428 se
rect 346 2415 2703 2428
rect 248 2403 281 2415
tri 281 2403 293 2415 nw
tri 321 2403 333 2415 se
rect 333 2403 2703 2415
rect 248 2388 260 2403
rect -87 2387 43 2388
tri 43 2387 44 2388 nw
tri 83 2387 84 2388 se
rect 84 2387 260 2388
rect -87 2382 38 2387
tri 38 2382 43 2387 nw
tri 78 2382 83 2387 se
rect 83 2382 260 2387
tri 260 2382 281 2403 nw
tri 300 2382 321 2403 se
rect 321 2382 2703 2403
rect -87 2176 33 2382
tri 33 2377 38 2382 nw
tri 73 2377 78 2382 se
rect 78 2377 253 2382
tri 71 2375 73 2377 se
rect 73 2375 253 2377
tri 253 2375 260 2382 nw
tri 293 2375 300 2382 se
rect 300 2375 2703 2382
rect 71 2363 241 2375
tri 241 2363 253 2375 nw
tri 281 2363 293 2375 se
rect 293 2363 2703 2375
rect 71 2332 210 2363
tri 210 2332 241 2363 nw
tri 250 2332 281 2363 se
rect 281 2332 2703 2363
rect 71 2292 170 2332
tri 170 2292 210 2332 nw
tri 210 2292 250 2332 se
rect 250 2321 2703 2332
tri 2703 2321 2822 2440 nw
rect 250 2292 380 2321
tri 380 2292 409 2321 nw
tri 1011 2296 1036 2321 ne
rect 1036 2320 2702 2321
tri 2702 2320 2703 2321 nw
rect 1036 2296 1241 2320
tri 1241 2296 1265 2320 nw
tri 2318 2296 2342 2320 ne
rect 2342 2296 2543 2320
rect 1036 2292 1237 2296
tri 1237 2292 1241 2296 nw
tri 2342 2295 2343 2296 ne
rect 2343 2292 2543 2296
tri 2543 2295 2568 2320 nw
rect 71 2280 158 2292
tri 158 2280 170 2292 nw
tri 198 2280 210 2292 se
rect 210 2280 368 2292
tri 368 2280 380 2292 nw
rect 470 2280 530 2292
rect 71 2270 148 2280
tri 148 2270 158 2280 nw
tri 188 2270 198 2280 se
rect 198 2270 358 2280
tri 358 2270 368 2280 nw
rect 71 2251 129 2270
tri 129 2251 148 2270 nw
tri 169 2251 188 2270 se
rect 188 2251 339 2270
tri 339 2251 358 2270 nw
tri 164 2246 169 2251 se
rect 169 2246 334 2251
tri 334 2246 339 2251 nw
rect 470 2246 479 2280
rect 513 2246 530 2280
tri 125 2207 164 2246 se
rect 164 2207 295 2246
tri 295 2207 334 2246 nw
rect 470 2207 530 2246
tri 119 2201 125 2207 se
rect 125 2201 264 2207
tri 33 2176 58 2201 sw
tri 94 2176 119 2201 se
rect 119 2176 264 2201
tri 264 2176 295 2207 nw
rect -87 1785 56 2176
rect 58 2175 94 2176
tri -87 1763 -65 1785 ne
rect -65 1763 56 1785
rect -181 1701 -135 1740
rect -181 1667 -175 1701
rect -141 1667 -135 1701
rect -181 1628 -135 1667
rect -181 1594 -175 1628
rect -141 1594 -135 1628
rect -181 1556 -135 1594
rect -181 1522 -175 1556
rect -141 1522 -135 1556
rect -181 1484 -135 1522
rect -181 1450 -175 1484
rect -141 1450 -135 1484
rect -181 1412 -135 1450
rect -181 1378 -175 1412
rect -141 1378 -135 1412
rect -181 1340 -135 1378
rect -181 1306 -175 1340
rect -141 1306 -135 1340
rect -181 1268 -135 1306
rect -181 1234 -175 1268
rect -141 1234 -135 1268
rect -181 1196 -135 1234
rect -181 1162 -175 1196
rect -141 1162 -135 1196
rect -181 1124 -135 1162
rect -181 1090 -175 1124
rect -141 1090 -135 1124
rect -181 1052 -135 1090
rect -181 1018 -175 1052
rect -141 1018 -135 1052
rect -181 980 -135 1018
rect -181 946 -175 980
rect -141 946 -135 980
rect -181 908 -135 946
rect -181 874 -175 908
rect -141 874 -135 908
rect -181 836 -135 874
rect -181 802 -175 836
rect -141 802 -135 836
rect -181 764 -135 802
rect -181 730 -175 764
rect -141 730 -135 764
rect -181 692 -135 730
rect -181 658 -175 692
rect -141 658 -135 692
rect -181 620 -135 658
rect -181 586 -175 620
rect -141 586 -135 620
rect -181 548 -135 586
rect -181 514 -175 548
rect -141 514 -135 548
rect -181 476 -135 514
rect -181 442 -175 476
rect -141 442 -135 476
rect -181 404 -135 442
rect -181 370 -175 404
rect -141 370 -135 404
rect -181 332 -135 370
rect -181 298 -175 332
rect -141 298 -135 332
rect -19 330 56 1763
rect 57 331 95 2175
rect 96 2173 261 2176
tri 261 2173 264 2176 nw
rect 470 2173 479 2207
rect 513 2173 530 2207
rect 96 2159 247 2173
tri 247 2159 261 2173 nw
rect 96 1785 239 2159
tri 239 2151 247 2159 nw
rect 287 2153 413 2159
rect 96 1763 217 1785
tri 217 1763 239 1785 nw
rect 287 2147 361 2153
rect 287 2113 293 2147
rect 327 2113 361 2147
rect 287 2101 361 2113
rect 287 2088 413 2101
rect 287 2075 361 2088
rect 287 2041 293 2075
rect 327 2041 361 2075
rect 287 2036 361 2041
rect 287 2022 413 2036
rect 287 2003 361 2022
rect 287 1969 293 2003
rect 327 1970 361 2003
rect 327 1969 413 1970
rect 287 1956 413 1969
rect 287 1931 361 1956
rect 287 1897 293 1931
rect 327 1904 361 1931
rect 327 1897 413 1904
rect 287 1890 413 1897
rect 287 1859 361 1890
rect 287 1825 293 1859
rect 327 1838 361 1859
rect 327 1825 413 1838
rect 287 1824 413 1825
rect 287 1787 361 1824
rect 96 395 171 1763
rect 287 1753 293 1787
rect 327 1772 361 1787
rect 327 1758 413 1772
rect 327 1753 361 1758
rect 287 1715 361 1753
rect 287 1681 293 1715
rect 327 1706 361 1715
rect 327 1692 413 1706
rect 327 1681 361 1692
rect 287 1643 361 1681
rect 287 1609 293 1643
rect 327 1640 361 1643
rect 327 1626 413 1640
rect 327 1609 361 1626
rect 287 1574 361 1609
rect 287 1571 413 1574
rect 287 1537 293 1571
rect 327 1560 413 1571
rect 327 1537 361 1560
rect 287 1508 361 1537
rect 287 1499 413 1508
rect 287 1465 293 1499
rect 327 1494 413 1499
rect 327 1465 361 1494
rect 287 1442 361 1465
rect 287 1428 413 1442
rect 287 1427 361 1428
rect 287 1393 293 1427
rect 327 1393 361 1427
rect 287 1376 361 1393
rect 287 1362 413 1376
rect 287 1355 361 1362
rect 287 1321 293 1355
rect 327 1321 361 1355
rect 287 1310 361 1321
rect 287 1296 413 1310
rect 287 1282 361 1296
rect 287 1248 293 1282
rect 327 1248 361 1282
rect 287 1244 361 1248
rect 287 1230 413 1244
rect 287 1209 361 1230
rect 287 1175 293 1209
rect 327 1178 361 1209
rect 327 1175 413 1178
rect 287 1164 413 1175
rect 287 1136 361 1164
rect 287 1102 293 1136
rect 327 1112 361 1136
rect 327 1102 413 1112
rect 287 1098 413 1102
rect 287 1063 361 1098
rect 287 1029 293 1063
rect 327 1046 361 1063
rect 327 1032 413 1046
rect 327 1029 361 1032
rect 287 990 361 1029
rect 287 956 293 990
rect 327 980 361 990
rect 327 966 413 980
rect 327 956 361 966
rect 287 917 361 956
rect 287 883 293 917
rect 327 914 361 917
rect 327 900 413 914
rect 327 883 361 900
rect 287 848 361 883
rect 287 844 413 848
rect 287 810 293 844
rect 327 834 413 844
rect 327 810 361 834
rect 287 782 361 810
rect 287 771 413 782
rect 287 737 293 771
rect 327 768 413 771
rect 327 737 361 768
rect 287 716 361 737
rect 287 702 413 716
rect 287 698 361 702
rect 287 664 293 698
rect 327 664 361 698
rect 287 650 361 664
rect 287 636 413 650
rect 287 625 361 636
rect 287 591 293 625
rect 327 591 361 625
rect 287 584 361 591
rect 287 570 413 584
rect 287 552 361 570
rect 287 518 293 552
rect 327 518 361 552
rect 287 504 413 518
rect 287 479 361 504
rect 287 445 293 479
rect 327 452 361 479
rect 327 445 413 452
rect 287 438 413 445
rect 287 406 361 438
rect 58 330 94 331
rect 96 330 217 395
rect 287 372 293 406
rect 327 386 361 406
rect 327 372 413 386
rect 287 333 361 372
rect -181 228 -135 298
rect 287 299 293 333
rect 327 320 361 333
rect 327 306 413 320
rect 327 299 361 306
rect 287 260 361 299
tri -135 228 -110 253 sw
tri 262 228 287 253 se
rect 287 228 293 260
rect -181 226 293 228
rect 327 254 361 260
rect 327 240 413 254
rect 327 226 361 240
rect -181 222 361 226
rect -181 188 -137 222
rect -103 188 -59 222
rect -25 188 19 222
rect 53 188 96 222
rect 130 188 173 222
rect 207 188 361 222
rect -181 182 413 188
rect 470 2134 530 2173
rect 470 2100 479 2134
rect 513 2100 530 2134
rect 470 2061 530 2100
rect 470 2027 479 2061
rect 513 2027 530 2061
rect 470 1988 530 2027
rect 470 1954 479 1988
rect 513 1954 530 1988
rect 470 1915 530 1954
rect 470 1881 479 1915
rect 513 1881 530 1915
rect 470 1842 530 1881
rect 470 1808 479 1842
rect 513 1808 530 1842
rect 470 1769 530 1808
rect 470 1735 479 1769
rect 513 1735 530 1769
rect 470 1696 530 1735
rect 470 1662 479 1696
rect 513 1662 530 1696
rect 470 1623 530 1662
rect 470 1589 479 1623
rect 513 1589 530 1623
rect 470 1550 530 1589
rect 470 1516 479 1550
rect 513 1516 530 1550
rect 470 1477 530 1516
rect 470 1443 479 1477
rect 513 1443 530 1477
rect 470 1404 530 1443
rect 470 1370 479 1404
rect 513 1370 530 1404
rect 470 1330 530 1370
rect 470 1296 479 1330
rect 513 1296 530 1330
rect 470 1256 530 1296
rect 470 1222 479 1256
rect 513 1222 530 1256
rect 470 1182 530 1222
rect 470 1148 479 1182
rect 513 1148 530 1182
rect 470 1108 530 1148
rect 470 1074 479 1108
rect 513 1074 530 1108
rect 470 1034 530 1074
rect 470 1000 479 1034
rect 513 1000 530 1034
rect 470 960 530 1000
rect 470 926 479 960
rect 513 926 530 960
rect 470 886 530 926
rect 470 852 479 886
rect 513 852 530 886
rect 470 812 530 852
rect 470 778 479 812
rect 513 778 530 812
rect 470 738 530 778
rect 470 704 479 738
rect 513 704 530 738
rect 470 664 530 704
rect 470 630 479 664
rect 513 630 530 664
rect 470 590 530 630
rect 470 556 479 590
rect 513 556 530 590
rect 470 516 530 556
rect 470 482 479 516
rect 513 482 530 516
rect 470 442 530 482
rect 470 408 479 442
rect 513 408 530 442
rect 470 368 530 408
rect 470 334 479 368
rect 513 334 530 368
rect 470 294 530 334
rect 470 260 479 294
rect 513 260 530 294
rect 470 220 530 260
rect 470 186 479 220
rect 513 186 530 220
tri 434 146 470 182 se
rect 470 146 530 186
rect -367 112 -361 146
rect -327 112 -321 146
tri 400 112 434 146 se
rect 434 112 479 146
rect 513 142 530 146
rect 542 2286 658 2292
rect 594 2234 606 2286
rect 542 2220 658 2234
rect 594 2168 606 2220
rect 542 2154 658 2168
rect 594 2102 606 2154
rect 542 2088 658 2102
rect 594 2036 606 2088
rect 542 2022 658 2036
rect 594 1970 606 2022
rect 542 1957 658 1970
rect 594 1905 606 1957
rect 542 1892 658 1905
rect 594 1840 606 1892
rect 542 1827 658 1840
rect 594 1775 606 1827
rect 542 1762 658 1775
rect 594 1710 606 1762
rect 542 1697 658 1710
rect 594 1645 606 1697
rect 542 1632 658 1645
rect 594 1580 606 1632
rect 542 1567 658 1580
rect 594 1515 606 1567
rect 542 1502 658 1515
rect 594 1450 606 1502
rect 542 1437 658 1450
rect 594 1385 606 1437
rect 542 1372 658 1385
rect 594 1320 606 1372
rect 542 1307 658 1320
rect 594 1255 606 1307
rect 542 1242 658 1255
rect 594 1190 606 1242
rect 542 1177 658 1190
rect 594 1125 606 1177
rect 542 1112 658 1125
rect 594 1060 606 1112
rect 542 1047 658 1060
rect 594 995 606 1047
rect 542 982 658 995
rect 594 930 606 982
rect 542 917 658 930
rect 594 865 606 917
rect 542 852 658 865
rect 594 800 606 852
rect 542 787 658 800
rect 594 735 606 787
rect 542 722 658 735
rect 594 670 606 722
rect 542 657 658 670
rect 594 605 606 657
rect 542 592 658 605
rect 594 540 606 592
rect 542 527 658 540
rect 594 475 606 527
rect 542 462 658 475
rect 594 410 606 462
rect 542 397 658 410
rect 594 345 606 397
rect 820 2286 1000 2292
rect 1036 2291 1236 2292
tri 1236 2291 1237 2292 nw
rect 872 2234 884 2286
rect 936 2234 948 2286
rect 820 2221 1000 2234
rect 872 2169 884 2221
rect 936 2169 948 2221
rect 820 2156 1000 2169
rect 872 2104 884 2156
rect 936 2104 948 2156
rect 820 2091 1000 2104
rect 872 2039 884 2091
rect 936 2039 948 2091
rect 820 2026 1000 2039
rect 872 1974 884 2026
rect 936 1974 948 2026
rect 820 1961 1000 1974
rect 872 1909 884 1961
rect 936 1909 948 1961
rect 820 1896 1000 1909
rect 872 1844 884 1896
rect 936 1844 948 1896
rect 820 1831 1000 1844
rect 872 1779 884 1831
rect 936 1779 948 1831
rect 820 1766 1000 1779
rect 872 1714 884 1766
rect 936 1714 948 1766
rect 820 1701 1000 1714
rect 872 1649 884 1701
rect 936 1649 948 1701
rect 820 1636 1000 1649
rect 872 1584 884 1636
rect 936 1584 948 1636
rect 820 1571 1000 1584
rect 872 1519 884 1571
rect 936 1519 948 1571
rect 820 1506 1000 1519
rect 872 1454 884 1506
rect 936 1454 948 1506
rect 820 1441 1000 1454
rect 872 1389 884 1441
rect 936 1389 948 1441
rect 820 1376 1000 1389
rect 1423 2286 1475 2292
rect 2589 2286 2769 2292
rect 1423 2221 1475 2234
tri 1894 2220 1919 2245 ne
tri 1919 2220 1944 2245 nw
rect 2641 2234 2653 2286
rect 2705 2234 2717 2286
rect 3180 2286 3296 2292
rect 2589 2220 2769 2234
rect 1423 2156 1475 2169
rect 1423 2091 1475 2104
rect 1423 2026 1475 2039
rect 1861 2203 1977 2209
rect 1913 2151 1925 2203
rect 1861 2138 1977 2151
rect 1913 2086 1925 2138
rect 1861 2073 1977 2086
rect 1913 2021 1925 2073
rect 1861 2008 1977 2021
rect 1423 1961 1475 1974
rect 1423 1896 1475 1909
rect 1423 1831 1475 1844
rect 1423 1766 1475 1779
rect 1423 1701 1475 1714
rect 1423 1636 1475 1649
rect 1423 1571 1475 1584
rect 1423 1506 1475 1519
rect 1423 1441 1475 1454
rect 1423 1376 1475 1389
rect 1423 1311 1475 1324
rect 1423 1246 1475 1259
rect 1423 1181 1475 1194
rect 1423 1116 1475 1129
rect 1423 1051 1475 1064
rect 1423 987 1475 999
rect 1423 923 1475 935
rect 1423 859 1475 871
rect 1423 795 1475 807
rect 1423 731 1475 743
rect 1423 667 1475 679
rect 1423 609 1475 615
rect 1581 1979 1697 1985
rect 1633 1927 1645 1979
rect 1581 1914 1697 1927
rect 1633 1862 1645 1914
rect 1581 1849 1697 1862
rect 1633 1797 1645 1849
rect 1581 1784 1697 1797
rect 1633 1732 1645 1784
rect 1581 1719 1697 1732
rect 1633 1667 1645 1719
rect 1581 1654 1697 1667
rect 1633 1602 1645 1654
rect 1581 1589 1697 1602
rect 1633 1537 1645 1589
rect 1581 1524 1697 1537
rect 1633 1472 1645 1524
rect 1581 1459 1697 1472
rect 1633 1407 1645 1459
rect 1581 1394 1697 1407
rect 1633 1342 1645 1394
rect 1581 1329 1697 1342
rect 1633 1277 1645 1329
rect 1581 1264 1697 1277
rect 1633 1212 1645 1264
rect 1581 1199 1697 1212
rect 1633 1147 1645 1199
rect 1581 1134 1697 1147
rect 1633 1082 1645 1134
rect 1581 1069 1697 1082
rect 1633 1017 1645 1069
rect 1581 1004 1697 1017
rect 1633 952 1645 1004
rect 1581 939 1697 952
rect 1633 887 1645 939
rect 1581 874 1697 887
rect 1633 822 1645 874
rect 1581 809 1697 822
tri 1100 500 1167 567 se
tri 1316 563 1320 567 sw
rect 1014 457 1167 500
rect 1184 557 1300 563
rect 1236 505 1248 557
rect 1184 488 1300 505
rect 820 358 1000 364
rect 1133 436 1184 457
rect 1236 436 1248 488
rect 1316 479 1320 563
tri 1320 479 1404 563 sw
rect 1316 457 1404 479
tri 1404 457 1426 479 sw
rect 1300 436 1350 457
rect 1133 419 1350 436
rect 1133 367 1184 419
rect 1236 367 1248 419
rect 1300 367 1350 419
rect 1581 367 1697 373
rect 1913 1956 1925 2008
rect 2641 2168 2653 2220
rect 2705 2168 2717 2220
rect 2589 2154 2769 2168
rect 2641 2102 2653 2154
rect 2705 2102 2717 2154
rect 2589 2088 2769 2102
rect 2641 2036 2653 2088
rect 2705 2036 2717 2088
rect 2589 2022 2769 2036
rect 1861 1943 1977 1956
rect 1913 1891 1925 1943
rect 1861 1878 1977 1891
rect 1913 1826 1925 1878
rect 1861 1813 1977 1826
rect 1913 1761 1925 1813
rect 1861 1748 1977 1761
rect 1913 1696 1925 1748
rect 1861 1683 1977 1696
rect 1913 1631 1925 1683
rect 1861 1618 1977 1631
rect 1913 1566 1925 1618
rect 1861 1553 1977 1566
rect 1913 1501 1925 1553
rect 1861 1488 1977 1501
rect 1913 1436 1925 1488
rect 1861 1423 1977 1436
rect 1913 1371 1925 1423
rect 1861 1358 1977 1371
rect 1913 1306 1925 1358
rect 1861 1293 1977 1306
rect 1913 1241 1925 1293
rect 1861 1228 1977 1241
rect 1913 1176 1925 1228
rect 1861 1163 1977 1176
rect 1913 1111 1925 1163
rect 1861 1098 1977 1111
rect 1913 1046 1925 1098
rect 1861 1033 1977 1046
rect 1913 981 1925 1033
rect 1861 968 1977 981
rect 1913 916 1925 968
rect 1861 903 1977 916
rect 1913 851 1925 903
rect 1861 838 1977 851
rect 1913 786 1925 838
rect 1861 773 1977 786
rect 1913 721 1925 773
rect 1861 708 1977 721
rect 542 332 658 345
rect 594 280 606 332
rect 1133 350 1350 367
rect 1133 298 1184 350
rect 1236 298 1248 350
rect 1300 298 1350 350
rect 1133 292 1350 298
tri 1133 286 1139 292 ne
rect 1139 286 1167 292
tri 1316 286 1322 292 nw
rect 542 267 658 280
rect 594 215 606 267
tri 1139 258 1167 286 ne
rect 542 202 658 215
rect 594 150 606 202
rect 542 144 658 150
rect 513 140 750 142
rect 513 128 1133 140
rect 513 112 673 128
rect -367 40 -321 112
tri 360 72 400 112 se
rect 400 76 673 112
rect 725 76 740 128
rect 792 76 807 128
rect 859 76 874 128
rect 926 76 941 128
rect 993 76 1008 128
rect 1060 76 1075 128
rect 1127 76 1133 128
rect 400 72 1133 76
tri 353 65 360 72 se
rect 360 65 479 72
tri -321 40 -296 65 sw
tri 328 40 353 65 se
rect 353 40 479 65
rect -367 38 479 40
rect 513 64 1133 72
rect 513 38 673 64
rect -367 34 673 38
rect -367 0 -323 34
rect -289 0 -247 34
rect -213 0 -171 34
rect -137 0 -95 34
rect -61 0 -19 34
rect 15 0 57 34
rect 91 0 133 34
rect 167 0 209 34
rect 243 0 285 34
rect 319 0 361 34
rect 395 12 673 34
rect 725 12 740 64
rect 792 12 807 64
rect 859 12 874 64
rect 926 12 941 64
rect 993 12 1008 64
rect 1060 12 1075 64
rect 1127 12 1133 64
rect 1350 76 1356 128
rect 1408 76 1423 128
rect 1475 76 1490 128
rect 1542 76 1557 128
rect 1609 76 1624 128
rect 1676 76 1691 128
rect 1743 76 1758 128
rect 1810 76 1816 128
rect 1350 64 1816 76
rect 2153 1990 2269 1996
rect 2205 1938 2217 1990
rect 2153 1926 2269 1938
rect 2153 1925 2217 1926
rect 2205 1874 2217 1925
rect 2205 1873 2269 1874
rect 2153 1862 2269 1873
rect 2153 1860 2217 1862
rect 2205 1810 2217 1860
rect 2205 1808 2269 1810
rect 2153 1798 2269 1808
rect 2153 1795 2217 1798
rect 2205 1746 2217 1795
rect 2205 1743 2269 1746
rect 2153 1734 2269 1743
rect 2153 1730 2217 1734
rect 2205 1682 2217 1730
rect 2205 1678 2269 1682
rect 2153 1670 2269 1678
rect 2153 1665 2217 1670
rect 2205 1618 2217 1665
rect 2205 1613 2269 1618
rect 2153 1606 2269 1613
rect 2153 1600 2217 1606
rect 2205 1554 2217 1600
rect 2205 1548 2269 1554
rect 2153 1542 2269 1548
rect 2153 1535 2217 1542
rect 2205 1490 2217 1535
rect 2205 1483 2269 1490
rect 2153 1478 2269 1483
rect 2153 1470 2217 1478
rect 2205 1426 2217 1470
rect 2205 1418 2269 1426
rect 2153 1414 2269 1418
rect 2153 1405 2217 1414
rect 2205 1362 2217 1405
rect 2205 1353 2269 1362
rect 2153 1350 2269 1353
rect 2153 1340 2217 1350
rect 2205 1298 2217 1340
rect 2205 1288 2269 1298
rect 2153 1285 2269 1288
rect 2153 1275 2217 1285
rect 2205 1233 2217 1275
rect 2205 1223 2269 1233
rect 2153 1220 2269 1223
rect 2153 1210 2217 1220
rect 2205 1168 2217 1210
rect 2205 1158 2269 1168
rect 2153 1155 2269 1158
rect 2153 1144 2217 1155
rect 2205 1103 2217 1144
rect 2205 1092 2269 1103
rect 2153 1090 2269 1092
rect 2153 1078 2217 1090
rect 2205 1038 2217 1078
rect 2205 1026 2269 1038
rect 2153 1025 2269 1026
rect 2153 1012 2217 1025
rect 2205 973 2217 1012
rect 2205 960 2269 973
rect 2153 946 2217 960
rect 2205 908 2217 946
rect 2205 895 2269 908
rect 2205 894 2217 895
rect 2153 880 2217 894
rect 2205 843 2217 880
rect 2205 830 2269 843
rect 2205 828 2217 830
rect 2153 814 2217 828
rect 2205 778 2217 814
rect 2205 765 2269 778
rect 2205 762 2217 765
rect 2153 748 2217 762
rect 2205 713 2217 748
rect 2205 700 2269 713
rect 2205 696 2217 700
rect 2153 682 2217 696
rect 2205 648 2217 682
rect 2641 1970 2653 2022
rect 2705 1970 2717 2022
rect 2589 1956 2769 1970
rect 2641 1904 2653 1956
rect 2705 1904 2717 1956
rect 2589 1890 2769 1904
rect 2641 1838 2653 1890
rect 2705 1838 2717 1890
rect 2589 1824 2769 1838
rect 2641 1772 2653 1824
rect 2705 1772 2717 1824
rect 2589 1759 2769 1772
rect 2641 1707 2653 1759
rect 2705 1707 2717 1759
rect 2589 1694 2769 1707
rect 2641 1642 2653 1694
rect 2705 1642 2717 1694
rect 2589 1629 2769 1642
rect 2641 1577 2653 1629
rect 2705 1577 2717 1629
rect 2589 1564 2769 1577
rect 2641 1512 2653 1564
rect 2705 1512 2717 1564
rect 2589 1499 2769 1512
rect 2641 1447 2653 1499
rect 2705 1447 2717 1499
rect 2589 1434 2769 1447
rect 2641 1382 2653 1434
rect 2705 1382 2717 1434
rect 2589 1369 2769 1382
rect 2641 1317 2653 1369
rect 2705 1317 2717 1369
rect 2589 1304 2769 1317
rect 2641 1252 2653 1304
rect 2705 1252 2717 1304
rect 2589 1239 2769 1252
rect 2641 1187 2653 1239
rect 2705 1187 2717 1239
rect 2589 1174 2769 1187
rect 2641 1122 2653 1174
rect 2705 1122 2717 1174
rect 2589 1109 2769 1122
rect 2641 1057 2653 1109
rect 2705 1057 2717 1109
rect 2589 1044 2769 1057
rect 2641 992 2653 1044
rect 2705 992 2717 1044
rect 2589 979 2769 992
rect 2641 927 2653 979
rect 2705 927 2717 979
rect 2589 914 2769 927
rect 2641 862 2653 914
rect 2705 862 2717 914
rect 2589 849 2769 862
rect 2641 797 2653 849
rect 2705 797 2717 849
rect 2589 784 2769 797
rect 2641 732 2653 784
rect 2705 732 2717 784
rect 2589 719 2769 732
rect 2641 667 2653 719
rect 2705 667 2717 719
rect 2589 661 2769 667
rect 2876 2270 2992 2276
rect 2876 1565 2992 1578
rect 2928 1513 2940 1565
rect 2876 1500 2992 1513
rect 2928 1448 2940 1500
rect 2876 1435 2992 1448
rect 2928 1383 2940 1435
rect 2876 1370 2992 1383
rect 2928 1318 2940 1370
rect 2876 1305 2992 1318
rect 2928 1253 2940 1305
rect 2876 1240 2992 1253
rect 2928 1188 2940 1240
rect 2876 1175 2992 1188
rect 2928 1123 2940 1175
rect 2876 1110 2992 1123
rect 2928 1058 2940 1110
rect 2876 1045 2992 1058
rect 2928 993 2940 1045
rect 2876 980 2992 993
rect 2928 928 2940 980
rect 2876 915 2992 928
rect 2928 863 2940 915
rect 2876 850 2992 863
rect 2928 798 2940 850
rect 2876 785 2992 798
rect 2928 733 2940 785
rect 2876 720 2992 733
rect 2928 668 2940 720
rect 2589 649 2602 661
rect 2876 655 2992 668
rect 2205 635 2269 648
rect 2205 630 2217 635
rect 2153 616 2217 630
rect 2205 583 2217 616
rect 2205 570 2269 583
rect 2205 564 2217 570
rect 2153 550 2217 564
rect 2205 518 2217 550
rect 2928 603 2940 655
rect 2876 590 2992 603
rect 2205 505 2269 518
rect 2205 498 2217 505
rect 2153 484 2217 498
rect 2205 453 2217 484
rect 2538 554 2654 560
rect 2590 502 2602 554
rect 2205 440 2269 453
rect 2205 432 2217 440
rect 2153 418 2217 432
rect 2205 388 2217 418
tri 2488 457 2522 491 se
rect 2538 485 2654 502
rect 2488 436 2538 457
rect 2482 433 2538 436
rect 2590 433 2602 485
rect 2928 538 2940 590
rect 2876 525 2992 538
tri 2671 457 2693 479 sw
rect 2928 473 2940 525
rect 2876 460 2992 473
rect 2654 433 2705 457
rect 2269 388 2311 429
rect 2205 377 2311 388
rect 2363 377 2388 429
rect 2205 366 2388 377
tri 2164 345 2185 366 ne
rect 2185 365 2388 366
rect 2185 345 2236 365
tri 2185 313 2217 345 ne
rect 2217 313 2236 345
rect 2288 313 2330 365
rect 2382 313 2388 365
rect 2482 417 2705 433
rect 2482 383 2494 417
rect 2528 383 2538 417
rect 2687 383 2705 417
rect 2482 365 2538 383
rect 2590 365 2602 383
rect 2654 365 2705 383
rect 2482 349 2705 365
rect 2482 345 2538 349
rect 2590 345 2602 349
rect 2654 345 2705 349
rect 2482 311 2494 345
rect 2528 311 2538 345
rect 2687 311 2705 345
rect 2928 408 2940 460
rect 2876 395 2992 408
rect 2928 343 2940 395
rect 2876 337 2992 343
rect 3232 2234 3244 2286
rect 3180 2220 3296 2234
rect 3232 2168 3244 2220
rect 3180 2154 3296 2168
rect 3232 2102 3244 2154
rect 3180 2088 3296 2102
rect 3232 2036 3244 2088
rect 3180 2022 3296 2036
rect 3232 1970 3244 2022
rect 3180 1957 3296 1970
rect 3232 1905 3244 1957
rect 3180 1892 3296 1905
rect 3232 1840 3244 1892
rect 3180 1827 3296 1840
rect 3232 1775 3244 1827
rect 3180 1762 3296 1775
rect 3232 1710 3244 1762
rect 3180 1697 3296 1710
rect 3232 1645 3244 1697
rect 3180 1632 3296 1645
rect 3232 1580 3244 1632
rect 3180 1567 3296 1580
rect 3232 1515 3244 1567
rect 3180 1502 3296 1515
rect 3232 1450 3244 1502
rect 3180 1437 3296 1450
rect 3232 1385 3244 1437
rect 3180 1372 3296 1385
rect 3232 1320 3244 1372
rect 3180 1307 3296 1320
rect 3232 1255 3244 1307
rect 3180 1242 3296 1255
rect 3232 1190 3244 1242
rect 3180 1177 3296 1190
rect 3232 1125 3244 1177
rect 3180 1112 3296 1125
rect 3232 1060 3244 1112
rect 3180 1047 3296 1060
rect 3232 995 3244 1047
rect 3180 982 3296 995
rect 3232 930 3244 982
rect 3180 917 3296 930
rect 3232 865 3244 917
rect 3180 852 3296 865
rect 3232 800 3244 852
rect 3180 787 3296 800
rect 3232 735 3244 787
rect 3180 722 3296 735
rect 3232 670 3244 722
rect 3180 657 3296 670
rect 3232 605 3244 657
rect 3180 592 3296 605
rect 3232 540 3244 592
rect 3180 527 3296 540
rect 3232 475 3244 527
rect 3180 462 3296 475
rect 3232 410 3244 462
rect 3180 397 3296 410
rect 3232 345 3244 397
rect 2482 297 2538 311
rect 2590 297 2602 311
rect 2654 297 2705 311
rect 2482 292 2705 297
tri 2488 258 2522 292 ne
rect 2538 291 2654 292
rect 2671 291 2704 292
tri 2704 291 2705 292 nw
rect 3180 332 3296 345
tri 2671 258 2704 291 nw
rect 3232 280 3244 332
rect 3180 267 3296 280
rect 3232 215 3244 267
rect 3180 202 3296 215
rect 3232 150 3244 202
rect 3180 144 3296 150
rect 1861 74 1977 80
rect 2014 76 2020 128
rect 2072 76 2087 128
rect 2139 76 2154 128
rect 2206 76 2221 128
rect 2273 76 2288 128
rect 2340 76 2355 128
rect 2407 76 2422 128
rect 2474 76 2480 128
rect 1350 12 1356 64
rect 1408 12 1423 64
rect 1475 12 1490 64
rect 1542 12 1557 64
rect 1609 12 1624 64
rect 1676 12 1691 64
rect 1743 12 1758 64
rect 1810 12 1816 64
tri 1894 47 1919 72 se
tri 1919 47 1944 72 sw
rect 2014 64 2480 76
rect 2014 12 2020 64
rect 2072 12 2087 64
rect 2139 12 2154 64
rect 2206 12 2221 64
rect 2273 12 2288 64
rect 2340 12 2355 64
rect 2407 12 2422 64
rect 2474 12 2480 64
rect 2705 76 2711 128
rect 2763 76 2778 128
rect 2830 76 2845 128
rect 2897 76 2912 128
rect 2964 76 2979 128
rect 3031 76 3046 128
rect 3098 76 3113 128
rect 3165 76 3171 128
rect 2705 64 3171 76
rect 2705 12 2711 64
rect 2763 12 2778 64
rect 2830 12 2845 64
rect 2897 12 2912 64
rect 2964 12 2979 64
rect 3031 12 3046 64
rect 3098 12 3113 64
rect 3165 12 3171 64
rect 395 0 1133 12
rect -367 -6 1133 0
<< rmetal1 >>
rect 56 2175 58 2176
rect 94 2175 96 2176
rect 56 331 57 2175
rect 95 331 96 2175
rect 56 330 58 331
rect 94 330 96 331
<< via1 >>
rect 2538 4851 2590 4903
rect 2602 4851 2654 4903
rect 1861 4771 1913 4823
rect 1925 4771 1977 4823
rect 1861 4706 1913 4758
rect 1925 4706 1977 4758
rect 1861 4641 1913 4693
rect 1925 4641 1977 4693
rect 1861 4576 1913 4628
rect 1925 4576 1977 4628
rect 2538 4784 2590 4836
rect 2602 4784 2654 4836
rect 2538 4717 2590 4769
rect 2602 4717 2654 4769
rect 2538 4650 2590 4702
rect 2602 4650 2654 4702
rect 828 4493 880 4545
rect 909 4493 961 4545
rect 990 4493 1042 4545
rect 828 4429 880 4481
rect 909 4429 961 4481
rect 990 4429 1042 4481
rect 1581 4492 1633 4544
rect 1645 4492 1697 4544
rect 1581 4426 1633 4478
rect 1645 4426 1697 4478
rect 947 4357 999 4409
rect 947 4293 999 4345
rect 1071 4341 1123 4393
rect 1192 4341 1244 4393
rect 1581 4360 1633 4412
rect 1645 4360 1697 4412
rect 1424 4242 1476 4294
rect 1424 4177 1476 4229
rect 1424 4112 1476 4164
rect 820 4015 872 4067
rect 884 4015 936 4067
rect 948 4015 1000 4067
rect 542 3943 594 3995
rect 606 3943 658 3995
rect 542 3876 594 3928
rect 606 3876 658 3928
rect 542 3810 594 3862
rect 606 3810 658 3862
rect 542 3744 594 3796
rect 606 3744 658 3796
rect 542 3678 594 3730
rect 606 3678 658 3730
rect 542 3612 594 3664
rect 606 3612 658 3664
rect 542 3546 594 3598
rect 606 3546 658 3598
rect 542 3480 594 3532
rect 606 3480 658 3532
rect 542 3414 594 3466
rect 606 3414 658 3466
rect 542 3348 594 3400
rect 606 3348 658 3400
rect 542 3282 594 3334
rect 606 3282 658 3334
rect 542 3216 594 3268
rect 606 3216 658 3268
rect 542 3150 594 3202
rect 606 3150 658 3202
rect 542 3084 594 3136
rect 606 3084 658 3136
rect 542 3018 594 3070
rect 606 3018 658 3070
rect 542 2952 594 3004
rect 606 2952 658 3004
rect 542 2886 594 2938
rect 606 2886 658 2938
rect 542 2820 594 2872
rect 606 2820 658 2872
rect 542 2754 594 2806
rect 606 2754 658 2806
rect 542 2688 594 2740
rect 606 2688 658 2740
rect 542 2622 594 2674
rect 606 2622 658 2674
rect 820 3949 872 4001
rect 884 3949 936 4001
rect 948 3949 1000 4001
rect 820 3883 872 3935
rect 884 3883 936 3935
rect 948 3883 1000 3935
rect 820 3817 872 3869
rect 884 3817 936 3869
rect 948 3817 1000 3869
rect 820 3751 872 3803
rect 884 3751 936 3803
rect 948 3751 1000 3803
rect 820 3685 872 3737
rect 884 3685 936 3737
rect 948 3685 1000 3737
rect 820 3619 872 3671
rect 884 3619 936 3671
rect 948 3619 1000 3671
rect 820 3553 872 3605
rect 884 3553 936 3605
rect 948 3553 1000 3605
rect 820 3487 872 3539
rect 884 3487 936 3539
rect 948 3487 1000 3539
rect 820 3422 872 3474
rect 884 3422 936 3474
rect 948 3422 1000 3474
rect 820 3357 872 3409
rect 884 3357 936 3409
rect 948 3357 1000 3409
rect 820 3292 872 3344
rect 884 3292 936 3344
rect 948 3292 1000 3344
rect 820 3227 872 3279
rect 884 3227 936 3279
rect 948 3227 1000 3279
rect 820 3162 872 3214
rect 884 3162 936 3214
rect 948 3162 1000 3214
rect 820 3097 872 3149
rect 884 3097 936 3149
rect 948 3097 1000 3149
rect 820 3032 872 3084
rect 884 3032 936 3084
rect 948 3032 1000 3084
rect 820 2967 872 3019
rect 884 2967 936 3019
rect 948 2967 1000 3019
rect 820 2902 872 2954
rect 884 2902 936 2954
rect 948 2902 1000 2954
rect 820 2837 872 2889
rect 884 2837 936 2889
rect 948 2837 1000 2889
rect 820 2772 872 2824
rect 884 2772 936 2824
rect 948 2772 1000 2824
rect 820 2707 872 2759
rect 884 2707 936 2759
rect 948 2707 1000 2759
rect 820 2642 872 2694
rect 884 2642 936 2694
rect 948 2642 1000 2694
rect 1424 4047 1476 4099
rect 1424 3982 1476 4034
rect 1424 3917 1476 3969
rect 1424 3852 1476 3904
rect 1424 3787 1476 3839
rect 1424 3722 1476 3774
rect 1424 3657 1476 3709
rect 1424 3592 1476 3644
rect 1424 3527 1476 3579
rect 1424 3462 1476 3514
rect 1424 3397 1476 3449
rect 1424 3332 1476 3384
rect 1424 3267 1476 3319
rect 1424 3202 1476 3254
rect 1424 3137 1476 3189
rect 1424 3072 1476 3124
rect 1424 3007 1476 3059
rect 1424 2943 1476 2995
rect 1424 2879 1476 2931
rect 1581 4294 1633 4346
rect 1645 4294 1697 4346
rect 1581 4228 1633 4280
rect 1645 4228 1697 4280
rect 1581 4162 1633 4214
rect 1645 4162 1697 4214
rect 1581 4096 1633 4148
rect 1645 4096 1697 4148
rect 1581 4030 1633 4082
rect 1645 4030 1697 4082
rect 1581 3964 1633 4016
rect 1645 3964 1697 4016
rect 1581 3898 1633 3950
rect 1645 3898 1697 3950
rect 1581 3832 1633 3884
rect 1645 3832 1697 3884
rect 1581 3766 1633 3818
rect 1645 3766 1697 3818
rect 1581 3700 1633 3752
rect 1645 3700 1697 3752
rect 1581 3634 1633 3686
rect 1645 3634 1697 3686
rect 1581 3568 1633 3620
rect 1645 3568 1697 3620
rect 1581 3503 1633 3555
rect 1645 3503 1697 3555
rect 1581 3438 1633 3490
rect 1645 3438 1697 3490
rect 1581 3373 1633 3425
rect 1645 3373 1697 3425
rect 1581 3308 1633 3360
rect 1645 3308 1697 3360
rect 1581 3243 1633 3295
rect 1645 3243 1697 3295
rect 1581 3178 1633 3230
rect 1645 3178 1697 3230
rect 1581 3113 1633 3165
rect 1645 3113 1697 3165
rect 1581 3048 1633 3100
rect 1645 3048 1697 3100
rect 1581 2983 1633 3035
rect 1645 2983 1697 3035
rect 1581 2918 1633 2970
rect 1645 2918 1697 2970
rect 1861 4511 1913 4563
rect 1925 4511 1977 4563
rect 2236 4543 2288 4595
rect 2330 4543 2382 4595
rect 1861 4446 1913 4498
rect 1925 4446 1977 4498
rect 1861 4381 1913 4433
rect 1925 4381 1977 4433
rect 1861 4316 1913 4368
rect 1925 4316 1977 4368
rect 1861 4251 1913 4303
rect 1925 4251 1977 4303
rect 1861 4186 1913 4238
rect 1925 4186 1977 4238
rect 1861 4121 1913 4173
rect 1925 4121 1977 4173
rect 1861 4056 1913 4108
rect 1925 4056 1977 4108
rect 1861 3991 1913 4043
rect 1925 3991 1977 4043
rect 1861 3926 1913 3978
rect 1925 3926 1977 3978
rect 1861 3861 1913 3913
rect 1925 3861 1977 3913
rect 1861 3796 1913 3848
rect 1925 3796 1977 3848
rect 1861 3731 1913 3783
rect 1925 3731 1977 3783
rect 1861 3666 1913 3718
rect 1925 3666 1977 3718
rect 1861 3601 1913 3653
rect 1925 3601 1977 3653
rect 1861 3536 1913 3588
rect 1925 3536 1977 3588
rect 1861 3471 1913 3523
rect 1925 3471 1977 3523
rect 1861 3406 1913 3458
rect 1925 3406 1977 3458
rect 1861 3341 1913 3393
rect 1925 3341 1977 3393
rect 1861 3276 1913 3328
rect 1925 3276 1977 3328
rect 1861 3211 1913 3263
rect 1925 3211 1977 3263
rect 1861 3146 1913 3198
rect 1925 3146 1977 3198
rect 1861 3081 1913 3133
rect 1925 3081 1977 3133
rect 1424 2815 1476 2867
rect 1424 2751 1476 2803
rect 1424 2687 1476 2739
rect 1861 2696 1977 3068
rect 2153 4490 2205 4542
rect 2153 4424 2205 4476
rect 2217 4468 2269 4520
rect 2311 4479 2363 4531
rect 2538 4584 2590 4636
rect 2602 4584 2654 4636
rect 3180 4711 3232 4763
rect 3244 4711 3296 4763
rect 3180 4645 3232 4697
rect 3244 4645 3296 4697
rect 3180 4579 3232 4631
rect 3244 4579 3296 4631
rect 2538 4518 2590 4570
rect 2602 4518 2654 4570
rect 2153 4358 2205 4410
rect 2217 4403 2269 4455
rect 2153 4292 2205 4344
rect 2217 4338 2269 4390
rect 2538 4452 2590 4504
rect 2602 4452 2654 4504
rect 2538 4386 2590 4438
rect 2602 4386 2654 4438
rect 2876 4513 2928 4565
rect 2940 4513 2992 4565
rect 2876 4448 2928 4500
rect 2940 4448 2992 4500
rect 2876 4383 2928 4435
rect 2940 4383 2992 4435
rect 2153 4226 2205 4278
rect 2217 4273 2269 4325
rect 2153 4160 2205 4212
rect 2217 4208 2269 4260
rect 2153 4094 2205 4146
rect 2217 4143 2269 4195
rect 2153 4028 2205 4080
rect 2217 4078 2269 4130
rect 2153 3962 2205 4014
rect 2217 4013 2269 4065
rect 2217 3948 2269 4000
rect 2153 3896 2205 3948
rect 2217 3883 2269 3935
rect 2153 3830 2205 3882
rect 2217 3818 2269 3870
rect 2153 3764 2205 3816
rect 2217 3753 2269 3805
rect 2153 3698 2205 3750
rect 2217 3688 2269 3740
rect 2153 3633 2205 3685
rect 2217 3623 2269 3675
rect 2153 3568 2205 3620
rect 2217 3558 2269 3610
rect 2153 3503 2205 3555
rect 2217 3494 2269 3546
rect 2153 3438 2205 3490
rect 2217 3430 2269 3482
rect 2153 3373 2205 3425
rect 2217 3366 2269 3418
rect 2153 3308 2205 3360
rect 2217 3302 2269 3354
rect 2153 3243 2205 3295
rect 2217 3238 2269 3290
rect 2153 3178 2205 3230
rect 2217 3174 2269 3226
rect 2153 3113 2205 3165
rect 2217 3110 2269 3162
rect 2153 3048 2205 3100
rect 2217 3046 2269 3098
rect 2153 2983 2205 3035
rect 2217 2982 2269 3034
rect 2153 2918 2205 2970
rect 2217 2918 2269 2970
rect 2589 4307 2641 4359
rect 2653 4307 2705 4359
rect 2717 4307 2769 4359
rect 2589 4242 2641 4294
rect 2653 4242 2705 4294
rect 2717 4242 2769 4294
rect 2876 4318 2928 4370
rect 2940 4318 2992 4370
rect 2589 4177 2641 4229
rect 2653 4177 2705 4229
rect 2717 4177 2769 4229
rect 2589 4112 2641 4164
rect 2653 4112 2705 4164
rect 2717 4112 2769 4164
rect 2589 4047 2641 4099
rect 2653 4047 2705 4099
rect 2717 4047 2769 4099
rect 2589 3982 2641 4034
rect 2653 3982 2705 4034
rect 2717 3982 2769 4034
rect 2589 3917 2641 3969
rect 2653 3917 2705 3969
rect 2717 3917 2769 3969
rect 2589 3852 2641 3904
rect 2653 3852 2705 3904
rect 2717 3852 2769 3904
rect 2589 3787 2641 3839
rect 2653 3787 2705 3839
rect 2717 3787 2769 3839
rect 2589 3722 2641 3774
rect 2653 3722 2705 3774
rect 2717 3722 2769 3774
rect 2589 3657 2641 3709
rect 2653 3657 2705 3709
rect 2717 3657 2769 3709
rect 2589 3592 2641 3644
rect 2653 3592 2705 3644
rect 2717 3592 2769 3644
rect 2589 3527 2641 3579
rect 2653 3527 2705 3579
rect 2717 3527 2769 3579
rect 2589 3462 2641 3514
rect 2653 3462 2705 3514
rect 2717 3462 2769 3514
rect 2589 3397 2641 3449
rect 2653 3397 2705 3449
rect 2717 3397 2769 3449
rect 2589 3332 2641 3384
rect 2653 3332 2705 3384
rect 2717 3332 2769 3384
rect 2589 3267 2641 3319
rect 2653 3267 2705 3319
rect 2717 3267 2769 3319
rect 2589 3202 2641 3254
rect 2653 3202 2705 3254
rect 2717 3202 2769 3254
rect 2589 3137 2641 3189
rect 2653 3137 2705 3189
rect 2717 3137 2769 3189
rect 2589 3072 2641 3124
rect 2653 3072 2705 3124
rect 2717 3072 2769 3124
rect 2589 3007 2641 3059
rect 2653 3007 2705 3059
rect 2717 3007 2769 3059
rect 1424 2623 1476 2675
rect 2589 2622 2769 2994
rect 2876 4253 2928 4305
rect 2940 4253 2992 4305
rect 2876 4188 2928 4240
rect 2940 4188 2992 4240
rect 2876 4123 2928 4175
rect 2940 4123 2992 4175
rect 2876 4058 2928 4110
rect 2940 4058 2992 4110
rect 2876 3993 2928 4045
rect 2940 3993 2992 4045
rect 2876 3928 2928 3980
rect 2940 3928 2992 3980
rect 2876 3863 2928 3915
rect 2940 3863 2992 3915
rect 2876 3798 2928 3850
rect 2940 3798 2992 3850
rect 2876 3733 2928 3785
rect 2940 3733 2992 3785
rect 2876 3668 2928 3720
rect 2940 3668 2992 3720
rect 2876 3603 2928 3655
rect 2940 3603 2992 3655
rect 2876 3538 2928 3590
rect 2940 3538 2992 3590
rect 2876 3473 2928 3525
rect 2940 3473 2992 3525
rect 2876 3408 2928 3460
rect 2940 3408 2992 3460
rect 2876 3343 2928 3395
rect 2940 3343 2992 3395
rect 2876 2638 2992 3330
rect 3180 4513 3232 4565
rect 3244 4513 3296 4565
rect 3180 4447 3232 4499
rect 3244 4447 3296 4499
rect 3180 4382 3232 4434
rect 3244 4382 3296 4434
rect 3180 4317 3232 4369
rect 3244 4317 3296 4369
rect 3180 4252 3232 4304
rect 3244 4252 3296 4304
rect 3180 4187 3232 4239
rect 3244 4187 3296 4239
rect 3180 4122 3232 4174
rect 3244 4122 3296 4174
rect 3180 4057 3232 4109
rect 3244 4057 3296 4109
rect 3180 3992 3232 4044
rect 3244 3992 3296 4044
rect 3180 3927 3232 3979
rect 3244 3927 3296 3979
rect 3180 3862 3232 3914
rect 3244 3862 3296 3914
rect 3180 3797 3232 3849
rect 3244 3797 3296 3849
rect 3180 3732 3232 3784
rect 3244 3732 3296 3784
rect 3180 3667 3232 3719
rect 3244 3667 3296 3719
rect 3180 3602 3232 3654
rect 3244 3602 3296 3654
rect 3180 3537 3232 3589
rect 3244 3537 3296 3589
rect 3180 3472 3232 3524
rect 3244 3472 3296 3524
rect 3180 3407 3232 3459
rect 3244 3407 3296 3459
rect 3180 3342 3232 3394
rect 3244 3342 3296 3394
rect 3180 3277 3232 3329
rect 3244 3277 3296 3329
rect 3180 3212 3232 3264
rect 3244 3212 3296 3264
rect 3180 3147 3232 3199
rect 3244 3147 3296 3199
rect 3180 3082 3232 3134
rect 3244 3082 3296 3134
rect 3180 3017 3232 3069
rect 3244 3017 3296 3069
rect 3180 2952 3232 3004
rect 3244 2952 3296 3004
rect 3180 2887 3232 2939
rect 3244 2887 3296 2939
rect 3180 2822 3232 2874
rect 3244 2822 3296 2874
rect 3180 2757 3232 2809
rect 3244 2757 3296 2809
rect 3180 2692 3232 2744
rect 3244 2692 3296 2744
rect 3180 2627 3232 2679
rect 3244 2627 3296 2679
rect 281 2527 333 2579
rect 281 2461 333 2513
rect 361 2101 413 2153
rect 361 2036 413 2088
rect 361 1970 413 2022
rect 361 1904 413 1956
rect 361 1838 413 1890
rect 361 1772 413 1824
rect 361 1706 413 1758
rect 361 1640 413 1692
rect 361 1574 413 1626
rect 361 1508 413 1560
rect 361 1442 413 1494
rect 361 1376 413 1428
rect 361 1310 413 1362
rect 361 1244 413 1296
rect 361 1178 413 1230
rect 361 1112 413 1164
rect 361 1046 413 1098
rect 361 980 413 1032
rect 361 914 413 966
rect 361 848 413 900
rect 361 782 413 834
rect 361 716 413 768
rect 361 650 413 702
rect 361 584 413 636
rect 361 518 413 570
rect 361 452 413 504
rect 361 386 413 438
rect 361 320 413 372
rect 361 254 413 306
rect 361 188 413 240
rect 542 2234 594 2286
rect 606 2234 658 2286
rect 542 2168 594 2220
rect 606 2168 658 2220
rect 542 2102 594 2154
rect 606 2102 658 2154
rect 542 2036 594 2088
rect 606 2036 658 2088
rect 542 1970 594 2022
rect 606 1970 658 2022
rect 542 1905 594 1957
rect 606 1905 658 1957
rect 542 1840 594 1892
rect 606 1840 658 1892
rect 542 1775 594 1827
rect 606 1775 658 1827
rect 542 1710 594 1762
rect 606 1710 658 1762
rect 542 1645 594 1697
rect 606 1645 658 1697
rect 542 1580 594 1632
rect 606 1580 658 1632
rect 542 1515 594 1567
rect 606 1515 658 1567
rect 542 1450 594 1502
rect 606 1450 658 1502
rect 542 1385 594 1437
rect 606 1385 658 1437
rect 542 1320 594 1372
rect 606 1320 658 1372
rect 542 1255 594 1307
rect 606 1255 658 1307
rect 542 1190 594 1242
rect 606 1190 658 1242
rect 542 1125 594 1177
rect 606 1125 658 1177
rect 542 1060 594 1112
rect 606 1060 658 1112
rect 542 995 594 1047
rect 606 995 658 1047
rect 542 930 594 982
rect 606 930 658 982
rect 542 865 594 917
rect 606 865 658 917
rect 542 800 594 852
rect 606 800 658 852
rect 542 735 594 787
rect 606 735 658 787
rect 542 670 594 722
rect 606 670 658 722
rect 542 605 594 657
rect 606 605 658 657
rect 542 540 594 592
rect 606 540 658 592
rect 542 475 594 527
rect 606 475 658 527
rect 542 410 594 462
rect 606 410 658 462
rect 542 345 594 397
rect 606 345 658 397
rect 820 2234 872 2286
rect 884 2234 936 2286
rect 948 2234 1000 2286
rect 820 2169 872 2221
rect 884 2169 936 2221
rect 948 2169 1000 2221
rect 820 2104 872 2156
rect 884 2104 936 2156
rect 948 2104 1000 2156
rect 820 2039 872 2091
rect 884 2039 936 2091
rect 948 2039 1000 2091
rect 820 1974 872 2026
rect 884 1974 936 2026
rect 948 1974 1000 2026
rect 820 1909 872 1961
rect 884 1909 936 1961
rect 948 1909 1000 1961
rect 820 1844 872 1896
rect 884 1844 936 1896
rect 948 1844 1000 1896
rect 820 1779 872 1831
rect 884 1779 936 1831
rect 948 1779 1000 1831
rect 820 1714 872 1766
rect 884 1714 936 1766
rect 948 1714 1000 1766
rect 820 1649 872 1701
rect 884 1649 936 1701
rect 948 1649 1000 1701
rect 820 1584 872 1636
rect 884 1584 936 1636
rect 948 1584 1000 1636
rect 820 1519 872 1571
rect 884 1519 936 1571
rect 948 1519 1000 1571
rect 820 1454 872 1506
rect 884 1454 936 1506
rect 948 1454 1000 1506
rect 820 1389 872 1441
rect 884 1389 936 1441
rect 948 1389 1000 1441
rect 820 364 1000 1376
rect 1423 2234 1475 2286
rect 1423 2169 1475 2221
rect 2589 2234 2641 2286
rect 2653 2234 2705 2286
rect 2717 2234 2769 2286
rect 1423 2104 1475 2156
rect 1423 2039 1475 2091
rect 1423 1974 1475 2026
rect 1861 2151 1913 2203
rect 1925 2151 1977 2203
rect 1861 2086 1913 2138
rect 1925 2086 1977 2138
rect 1861 2021 1913 2073
rect 1925 2021 1977 2073
rect 1423 1909 1475 1961
rect 1423 1844 1475 1896
rect 1423 1779 1475 1831
rect 1423 1714 1475 1766
rect 1423 1649 1475 1701
rect 1423 1584 1475 1636
rect 1423 1519 1475 1571
rect 1423 1454 1475 1506
rect 1423 1389 1475 1441
rect 1423 1324 1475 1376
rect 1423 1259 1475 1311
rect 1423 1194 1475 1246
rect 1423 1129 1475 1181
rect 1423 1064 1475 1116
rect 1423 999 1475 1051
rect 1423 935 1475 987
rect 1423 871 1475 923
rect 1423 807 1475 859
rect 1423 743 1475 795
rect 1423 679 1475 731
rect 1423 615 1475 667
rect 1581 1927 1633 1979
rect 1645 1927 1697 1979
rect 1581 1862 1633 1914
rect 1645 1862 1697 1914
rect 1581 1797 1633 1849
rect 1645 1797 1697 1849
rect 1581 1732 1633 1784
rect 1645 1732 1697 1784
rect 1581 1667 1633 1719
rect 1645 1667 1697 1719
rect 1581 1602 1633 1654
rect 1645 1602 1697 1654
rect 1581 1537 1633 1589
rect 1645 1537 1697 1589
rect 1581 1472 1633 1524
rect 1645 1472 1697 1524
rect 1581 1407 1633 1459
rect 1645 1407 1697 1459
rect 1581 1342 1633 1394
rect 1645 1342 1697 1394
rect 1581 1277 1633 1329
rect 1645 1277 1697 1329
rect 1581 1212 1633 1264
rect 1645 1212 1697 1264
rect 1581 1147 1633 1199
rect 1645 1147 1697 1199
rect 1581 1082 1633 1134
rect 1645 1082 1697 1134
rect 1581 1017 1633 1069
rect 1645 1017 1697 1069
rect 1581 952 1633 1004
rect 1645 952 1697 1004
rect 1581 887 1633 939
rect 1645 887 1697 939
rect 1581 822 1633 874
rect 1645 822 1697 874
rect 1184 505 1236 557
rect 1248 505 1300 557
rect 1184 436 1236 488
rect 1248 436 1300 488
rect 1184 367 1236 419
rect 1248 367 1300 419
rect 1581 373 1697 809
rect 1861 1956 1913 2008
rect 1925 1956 1977 2008
rect 2589 2168 2641 2220
rect 2653 2168 2705 2220
rect 2717 2168 2769 2220
rect 2589 2102 2641 2154
rect 2653 2102 2705 2154
rect 2717 2102 2769 2154
rect 2589 2036 2641 2088
rect 2653 2036 2705 2088
rect 2717 2036 2769 2088
rect 1861 1891 1913 1943
rect 1925 1891 1977 1943
rect 1861 1826 1913 1878
rect 1925 1826 1977 1878
rect 1861 1761 1913 1813
rect 1925 1761 1977 1813
rect 1861 1696 1913 1748
rect 1925 1696 1977 1748
rect 1861 1631 1913 1683
rect 1925 1631 1977 1683
rect 1861 1566 1913 1618
rect 1925 1566 1977 1618
rect 1861 1501 1913 1553
rect 1925 1501 1977 1553
rect 1861 1436 1913 1488
rect 1925 1436 1977 1488
rect 1861 1371 1913 1423
rect 1925 1371 1977 1423
rect 1861 1306 1913 1358
rect 1925 1306 1977 1358
rect 1861 1241 1913 1293
rect 1925 1241 1977 1293
rect 1861 1176 1913 1228
rect 1925 1176 1977 1228
rect 1861 1111 1913 1163
rect 1925 1111 1977 1163
rect 1861 1046 1913 1098
rect 1925 1046 1977 1098
rect 1861 981 1913 1033
rect 1925 981 1977 1033
rect 1861 916 1913 968
rect 1925 916 1977 968
rect 1861 851 1913 903
rect 1925 851 1977 903
rect 1861 786 1913 838
rect 1925 786 1977 838
rect 1861 721 1913 773
rect 1925 721 1977 773
rect 542 280 594 332
rect 606 280 658 332
rect 1184 298 1236 350
rect 1248 298 1300 350
rect 542 215 594 267
rect 606 215 658 267
rect 542 150 594 202
rect 606 150 658 202
rect 673 76 725 128
rect 740 76 792 128
rect 807 76 859 128
rect 874 76 926 128
rect 941 76 993 128
rect 1008 76 1060 128
rect 1075 76 1127 128
rect 673 12 725 64
rect 740 12 792 64
rect 807 12 859 64
rect 874 12 926 64
rect 941 12 993 64
rect 1008 12 1060 64
rect 1075 12 1127 64
rect 1356 76 1408 128
rect 1423 76 1475 128
rect 1490 76 1542 128
rect 1557 76 1609 128
rect 1624 76 1676 128
rect 1691 76 1743 128
rect 1758 76 1810 128
rect 1861 80 1977 708
rect 2153 1938 2205 1990
rect 2217 1938 2269 1990
rect 2153 1873 2205 1925
rect 2217 1874 2269 1926
rect 2153 1808 2205 1860
rect 2217 1810 2269 1862
rect 2153 1743 2205 1795
rect 2217 1746 2269 1798
rect 2153 1678 2205 1730
rect 2217 1682 2269 1734
rect 2153 1613 2205 1665
rect 2217 1618 2269 1670
rect 2153 1548 2205 1600
rect 2217 1554 2269 1606
rect 2153 1483 2205 1535
rect 2217 1490 2269 1542
rect 2153 1418 2205 1470
rect 2217 1426 2269 1478
rect 2153 1353 2205 1405
rect 2217 1362 2269 1414
rect 2153 1288 2205 1340
rect 2217 1298 2269 1350
rect 2153 1223 2205 1275
rect 2217 1233 2269 1285
rect 2153 1158 2205 1210
rect 2217 1168 2269 1220
rect 2153 1092 2205 1144
rect 2217 1103 2269 1155
rect 2153 1026 2205 1078
rect 2217 1038 2269 1090
rect 2153 960 2205 1012
rect 2217 973 2269 1025
rect 2153 894 2205 946
rect 2217 908 2269 960
rect 2153 828 2205 880
rect 2217 843 2269 895
rect 2153 762 2205 814
rect 2217 778 2269 830
rect 2153 696 2205 748
rect 2217 713 2269 765
rect 2153 630 2205 682
rect 2217 648 2269 700
rect 2589 1970 2641 2022
rect 2653 1970 2705 2022
rect 2717 1970 2769 2022
rect 2589 1904 2641 1956
rect 2653 1904 2705 1956
rect 2717 1904 2769 1956
rect 2589 1838 2641 1890
rect 2653 1838 2705 1890
rect 2717 1838 2769 1890
rect 2589 1772 2641 1824
rect 2653 1772 2705 1824
rect 2717 1772 2769 1824
rect 2589 1707 2641 1759
rect 2653 1707 2705 1759
rect 2717 1707 2769 1759
rect 2589 1642 2641 1694
rect 2653 1642 2705 1694
rect 2717 1642 2769 1694
rect 2589 1577 2641 1629
rect 2653 1577 2705 1629
rect 2717 1577 2769 1629
rect 2589 1512 2641 1564
rect 2653 1512 2705 1564
rect 2717 1512 2769 1564
rect 2589 1447 2641 1499
rect 2653 1447 2705 1499
rect 2717 1447 2769 1499
rect 2589 1382 2641 1434
rect 2653 1382 2705 1434
rect 2717 1382 2769 1434
rect 2589 1317 2641 1369
rect 2653 1317 2705 1369
rect 2717 1317 2769 1369
rect 2589 1252 2641 1304
rect 2653 1252 2705 1304
rect 2717 1252 2769 1304
rect 2589 1187 2641 1239
rect 2653 1187 2705 1239
rect 2717 1187 2769 1239
rect 2589 1122 2641 1174
rect 2653 1122 2705 1174
rect 2717 1122 2769 1174
rect 2589 1057 2641 1109
rect 2653 1057 2705 1109
rect 2717 1057 2769 1109
rect 2589 992 2641 1044
rect 2653 992 2705 1044
rect 2717 992 2769 1044
rect 2589 927 2641 979
rect 2653 927 2705 979
rect 2717 927 2769 979
rect 2589 862 2641 914
rect 2653 862 2705 914
rect 2717 862 2769 914
rect 2589 797 2641 849
rect 2653 797 2705 849
rect 2717 797 2769 849
rect 2589 732 2641 784
rect 2653 732 2705 784
rect 2717 732 2769 784
rect 2589 667 2641 719
rect 2653 667 2705 719
rect 2717 667 2769 719
rect 2876 1578 2992 2270
rect 2876 1513 2928 1565
rect 2940 1513 2992 1565
rect 2876 1448 2928 1500
rect 2940 1448 2992 1500
rect 2876 1383 2928 1435
rect 2940 1383 2992 1435
rect 2876 1318 2928 1370
rect 2940 1318 2992 1370
rect 2876 1253 2928 1305
rect 2940 1253 2992 1305
rect 2876 1188 2928 1240
rect 2940 1188 2992 1240
rect 2876 1123 2928 1175
rect 2940 1123 2992 1175
rect 2876 1058 2928 1110
rect 2940 1058 2992 1110
rect 2876 993 2928 1045
rect 2940 993 2992 1045
rect 2876 928 2928 980
rect 2940 928 2992 980
rect 2876 863 2928 915
rect 2940 863 2992 915
rect 2876 798 2928 850
rect 2940 798 2992 850
rect 2876 733 2928 785
rect 2940 733 2992 785
rect 2876 668 2928 720
rect 2940 668 2992 720
rect 2153 564 2205 616
rect 2217 583 2269 635
rect 2153 498 2205 550
rect 2217 518 2269 570
rect 2876 603 2928 655
rect 2940 603 2992 655
rect 2153 432 2205 484
rect 2217 453 2269 505
rect 2538 502 2590 554
rect 2602 502 2654 554
rect 2153 366 2205 418
rect 2217 388 2269 440
rect 2538 433 2590 485
rect 2602 433 2654 485
rect 2876 538 2928 590
rect 2940 538 2992 590
rect 2876 473 2928 525
rect 2940 473 2992 525
rect 2311 377 2363 429
rect 2236 313 2288 365
rect 2330 313 2382 365
rect 2538 383 2574 417
rect 2574 383 2590 417
rect 2602 383 2608 417
rect 2608 383 2653 417
rect 2653 383 2654 417
rect 2538 365 2590 383
rect 2602 365 2654 383
rect 2538 345 2590 349
rect 2602 345 2654 349
rect 2538 311 2574 345
rect 2574 311 2590 345
rect 2602 311 2608 345
rect 2608 311 2653 345
rect 2653 311 2654 345
rect 2876 408 2928 460
rect 2940 408 2992 460
rect 2876 343 2928 395
rect 2940 343 2992 395
rect 3180 2234 3232 2286
rect 3244 2234 3296 2286
rect 3180 2168 3232 2220
rect 3244 2168 3296 2220
rect 3180 2102 3232 2154
rect 3244 2102 3296 2154
rect 3180 2036 3232 2088
rect 3244 2036 3296 2088
rect 3180 1970 3232 2022
rect 3244 1970 3296 2022
rect 3180 1905 3232 1957
rect 3244 1905 3296 1957
rect 3180 1840 3232 1892
rect 3244 1840 3296 1892
rect 3180 1775 3232 1827
rect 3244 1775 3296 1827
rect 3180 1710 3232 1762
rect 3244 1710 3296 1762
rect 3180 1645 3232 1697
rect 3244 1645 3296 1697
rect 3180 1580 3232 1632
rect 3244 1580 3296 1632
rect 3180 1515 3232 1567
rect 3244 1515 3296 1567
rect 3180 1450 3232 1502
rect 3244 1450 3296 1502
rect 3180 1385 3232 1437
rect 3244 1385 3296 1437
rect 3180 1320 3232 1372
rect 3244 1320 3296 1372
rect 3180 1255 3232 1307
rect 3244 1255 3296 1307
rect 3180 1190 3232 1242
rect 3244 1190 3296 1242
rect 3180 1125 3232 1177
rect 3244 1125 3296 1177
rect 3180 1060 3232 1112
rect 3244 1060 3296 1112
rect 3180 995 3232 1047
rect 3244 995 3296 1047
rect 3180 930 3232 982
rect 3244 930 3296 982
rect 3180 865 3232 917
rect 3244 865 3296 917
rect 3180 800 3232 852
rect 3244 800 3296 852
rect 3180 735 3232 787
rect 3244 735 3296 787
rect 3180 670 3232 722
rect 3244 670 3296 722
rect 3180 605 3232 657
rect 3244 605 3296 657
rect 3180 540 3232 592
rect 3244 540 3296 592
rect 3180 475 3232 527
rect 3244 475 3296 527
rect 3180 410 3232 462
rect 3244 410 3296 462
rect 3180 345 3232 397
rect 3244 345 3296 397
rect 2538 297 2590 311
rect 2602 297 2654 311
rect 3180 280 3232 332
rect 3244 280 3296 332
rect 3180 215 3232 267
rect 3244 215 3296 267
rect 3180 150 3232 202
rect 3244 150 3296 202
rect 2020 76 2072 128
rect 2087 76 2139 128
rect 2154 76 2206 128
rect 2221 76 2273 128
rect 2288 76 2340 128
rect 2355 76 2407 128
rect 2422 76 2474 128
rect 1356 12 1408 64
rect 1423 12 1475 64
rect 1490 12 1542 64
rect 1557 12 1609 64
rect 1624 12 1676 64
rect 1691 12 1743 64
rect 1758 12 1810 64
rect 2020 12 2072 64
rect 2087 12 2139 64
rect 2154 12 2206 64
rect 2221 12 2273 64
rect 2288 12 2340 64
rect 2355 12 2407 64
rect 2422 12 2474 64
rect 2711 76 2763 128
rect 2778 76 2830 128
rect 2845 76 2897 128
rect 2912 76 2964 128
rect 2979 76 3031 128
rect 3046 76 3098 128
rect 3113 76 3165 128
rect 2711 12 2763 64
rect 2778 12 2830 64
rect 2845 12 2897 64
rect 2912 12 2964 64
rect 2979 12 3031 64
rect 3046 12 3098 64
rect 3113 12 3165 64
<< metal2 >>
tri 1928 5253 2071 5396 se
rect 2071 5253 2384 5505
tri 1571 5060 1764 5253 se
rect 1764 5060 2384 5253
rect -67 1955 253 5041
rect 281 2579 333 5041
tri 394 5009 422 5037 se
rect 422 5009 1035 5041
rect 394 4636 1035 5009
rect 1218 4945 2384 5060
tri 2574 4945 2585 4956 se
rect 2585 4945 2768 5505
rect 1218 4903 1745 4945
tri 1745 4903 1787 4945 nw
tri 2538 4909 2574 4945 se
rect 2574 4909 2768 4945
tri 2532 4903 2538 4909 se
rect 2538 4903 2768 4909
rect 1218 4851 1693 4903
tri 1693 4851 1745 4903 nw
tri 2480 4851 2532 4903 se
rect 2532 4851 2538 4903
rect 2590 4851 2602 4903
rect 2654 4851 2768 4903
rect 1218 4836 1678 4851
tri 1678 4836 1693 4851 nw
tri 2465 4836 2480 4851 se
rect 2480 4836 2768 4851
rect 1218 4823 1665 4836
tri 1665 4823 1678 4836 nw
rect 1743 4823 2040 4836
rect 1218 4774 1616 4823
tri 1616 4774 1665 4823 nw
tri 1035 4636 1036 4637 sw
rect 394 4628 1036 4636
tri 1036 4628 1044 4636 sw
rect 394 4576 1044 4628
tri 1044 4576 1096 4628 sw
rect 394 4563 1096 4576
tri 1096 4563 1109 4576 sw
rect 1218 4563 1539 4774
rect 394 4549 1109 4563
tri 1109 4549 1123 4563 sw
tri 1218 4549 1232 4563 ne
rect 1232 4549 1539 4563
rect 1743 4771 1861 4823
rect 1913 4771 1925 4823
rect 1977 4771 2040 4823
rect 1743 4758 2040 4771
rect 1743 4706 1861 4758
rect 1913 4706 1925 4758
rect 1977 4706 2040 4758
rect 1743 4693 2040 4706
rect 1743 4641 1861 4693
rect 1913 4641 1925 4693
rect 1977 4641 2040 4693
tri 2415 4786 2465 4836 se
rect 2465 4786 2538 4836
rect 2415 4784 2538 4786
rect 2590 4784 2602 4836
rect 2654 4801 2768 4836
tri 2768 4801 2769 4802 sw
rect 2654 4784 2769 4801
rect 2415 4769 2769 4784
rect 2415 4717 2538 4769
rect 2590 4717 2602 4769
rect 2654 4717 2769 4769
rect 2415 4702 2769 4717
rect 2415 4657 2538 4702
tri 2415 4656 2416 4657 ne
rect 1743 4628 2040 4641
rect 1743 4576 1861 4628
rect 1913 4576 1925 4628
rect 1977 4576 2040 4628
rect 2416 4650 2538 4657
rect 2590 4650 2602 4702
rect 2654 4650 2769 4702
rect 2416 4636 2769 4650
rect 1743 4563 2040 4576
rect 394 4545 1123 4549
rect 394 4493 828 4545
rect 880 4493 909 4545
rect 961 4493 990 4545
rect 1042 4544 1123 4545
tri 1123 4544 1128 4549 sw
tri 1232 4544 1237 4549 ne
rect 1237 4544 1539 4549
rect 1042 4493 1128 4544
rect 394 4492 1128 4493
tri 1128 4492 1180 4544 sw
tri 1237 4492 1289 4544 ne
rect 1289 4492 1539 4544
rect 394 4481 1180 4492
rect 394 4429 828 4481
rect 880 4429 909 4481
rect 961 4429 990 4481
rect 1042 4478 1180 4481
tri 1180 4478 1194 4492 sw
tri 1289 4478 1303 4492 ne
rect 1303 4478 1539 4492
rect 1042 4454 1194 4478
tri 1194 4454 1218 4478 sw
tri 1303 4454 1327 4478 ne
rect 1327 4454 1539 4478
rect 1042 4429 1218 4454
rect 394 4426 1218 4429
tri 1218 4426 1246 4454 sw
tri 1327 4426 1355 4454 ne
rect 1355 4426 1539 4454
rect 394 4425 1246 4426
tri 1246 4425 1247 4426 sw
tri 1355 4425 1356 4426 ne
rect 1356 4425 1539 4426
rect 394 4415 1247 4425
tri 1247 4415 1257 4425 sw
tri 1356 4415 1366 4425 ne
rect 1366 4415 1539 4425
rect 394 4412 1257 4415
tri 1257 4412 1260 4415 sw
tri 1366 4412 1369 4415 ne
rect 1369 4412 1539 4415
rect 394 4409 1260 4412
rect 394 4357 947 4409
rect 999 4393 1260 4409
rect 999 4357 1071 4393
rect 394 4345 1071 4357
tri 391 4293 394 4296 se
rect 394 4293 947 4345
rect 999 4341 1071 4345
rect 1123 4341 1192 4393
rect 1244 4365 1260 4393
tri 1260 4365 1307 4412 sw
tri 1369 4365 1416 4412 ne
rect 1416 4365 1539 4412
rect 1244 4360 1307 4365
tri 1307 4360 1312 4365 sw
tri 1416 4360 1421 4365 ne
rect 1421 4360 1539 4365
rect 1244 4358 1312 4360
tri 1312 4358 1314 4360 sw
tri 1421 4358 1423 4360 ne
rect 1244 4346 1314 4358
tri 1314 4346 1326 4358 sw
rect 1244 4341 1326 4346
rect 999 4305 1326 4341
tri 1326 4305 1367 4346 sw
rect 999 4293 1367 4305
rect 281 2513 333 2527
rect 281 2455 333 2461
tri 361 4263 391 4293 se
rect 391 4263 1367 4293
rect 361 4225 1367 4263
rect 361 2153 502 4225
tri 502 4195 532 4225 nw
tri 683 4195 713 4225 ne
rect 713 4195 1367 4225
tri 713 4180 728 4195 ne
rect 728 4067 1367 4195
rect 728 4015 820 4067
rect 872 4015 884 4067
rect 936 4015 948 4067
rect 1000 4015 1367 4067
rect 728 4001 1367 4015
rect 413 2101 502 2153
rect 361 2088 502 2101
rect 413 2036 502 2088
rect 361 2022 502 2036
rect 413 1970 502 2022
rect 361 1956 502 1970
rect 413 1904 502 1956
rect 361 1890 502 1904
rect 413 1838 502 1890
rect 361 1824 502 1838
rect 413 1772 502 1824
rect 361 1758 502 1772
rect 413 1706 502 1758
rect 361 1692 502 1706
rect 413 1640 502 1692
rect 361 1626 502 1640
rect 413 1574 502 1626
rect 361 1560 502 1574
rect 413 1508 502 1560
rect 361 1494 502 1508
rect 413 1442 502 1494
rect 361 1428 502 1442
rect 413 1376 502 1428
rect 361 1362 502 1376
rect 413 1310 502 1362
rect 361 1296 502 1310
rect 413 1244 502 1296
rect 361 1230 502 1244
rect 413 1178 502 1230
rect 361 1164 502 1178
rect 413 1112 502 1164
rect 361 1098 502 1112
rect 413 1046 502 1098
rect 361 1032 502 1046
rect 413 980 502 1032
rect 361 966 502 980
rect 413 914 502 966
rect 361 900 502 914
rect 413 848 502 900
rect 361 834 502 848
rect 413 782 502 834
rect 361 768 502 782
rect 413 716 502 768
rect 361 702 502 716
rect 413 650 502 702
rect 361 636 502 650
rect 413 584 502 636
rect 361 570 502 584
rect 413 518 502 570
rect 361 504 502 518
rect 413 452 502 504
rect 361 438 502 452
rect 413 386 502 438
rect 361 372 502 386
rect 413 320 502 372
rect 361 306 502 320
rect 413 254 502 306
rect 361 240 502 254
rect 413 188 502 240
rect 361 182 502 188
rect 530 3995 671 4001
rect 530 3943 542 3995
rect 594 3943 606 3995
rect 658 3943 671 3995
rect 530 3928 671 3943
rect 530 3876 542 3928
rect 594 3876 606 3928
rect 658 3876 671 3928
rect 530 3862 671 3876
rect 530 3810 542 3862
rect 594 3810 606 3862
rect 658 3810 671 3862
rect 530 3796 671 3810
rect 530 3744 542 3796
rect 594 3744 606 3796
rect 658 3744 671 3796
rect 530 3730 671 3744
rect 530 3678 542 3730
rect 594 3678 606 3730
rect 658 3678 671 3730
rect 530 3664 671 3678
rect 530 3612 542 3664
rect 594 3612 606 3664
rect 658 3612 671 3664
rect 530 3598 671 3612
rect 530 3546 542 3598
rect 594 3546 606 3598
rect 658 3546 671 3598
rect 530 3532 671 3546
rect 530 3480 542 3532
rect 594 3480 606 3532
rect 658 3480 671 3532
rect 530 3466 671 3480
rect 530 3414 542 3466
rect 594 3414 606 3466
rect 658 3414 671 3466
rect 530 3400 671 3414
rect 530 3348 542 3400
rect 594 3348 606 3400
rect 658 3348 671 3400
rect 530 3334 671 3348
rect 530 3282 542 3334
rect 594 3282 606 3334
rect 658 3282 671 3334
rect 530 3268 671 3282
rect 530 3216 542 3268
rect 594 3216 606 3268
rect 658 3216 671 3268
rect 530 3202 671 3216
rect 530 3150 542 3202
rect 594 3150 606 3202
rect 658 3150 671 3202
rect 530 3136 671 3150
rect 530 3084 542 3136
rect 594 3084 606 3136
rect 658 3084 671 3136
rect 530 3070 671 3084
rect 530 3018 542 3070
rect 594 3018 606 3070
rect 658 3018 671 3070
rect 530 3004 671 3018
rect 530 2952 542 3004
rect 594 2952 606 3004
rect 658 2952 671 3004
rect 530 2938 671 2952
rect 530 2886 542 2938
rect 594 2886 606 2938
rect 658 2886 671 2938
rect 530 2872 671 2886
rect 530 2820 542 2872
rect 594 2820 606 2872
rect 658 2820 671 2872
rect 530 2806 671 2820
rect 530 2754 542 2806
rect 594 2754 606 2806
rect 658 2754 671 2806
rect 530 2740 671 2754
rect 530 2688 542 2740
rect 594 2688 606 2740
rect 658 2688 671 2740
rect 530 2674 671 2688
rect 530 2622 542 2674
rect 594 2622 606 2674
rect 658 2622 671 2674
rect 530 2286 671 2622
rect 530 2234 542 2286
rect 594 2234 606 2286
rect 658 2234 671 2286
rect 530 2220 671 2234
rect 530 2168 542 2220
rect 594 2168 606 2220
rect 658 2168 671 2220
rect 530 2154 671 2168
rect 530 2102 542 2154
rect 594 2102 606 2154
rect 658 2102 671 2154
rect 530 2088 671 2102
rect 530 2036 542 2088
rect 594 2036 606 2088
rect 658 2036 671 2088
rect 530 2022 671 2036
rect 530 1970 542 2022
rect 594 1970 606 2022
rect 658 1970 671 2022
rect 530 1957 671 1970
rect 530 1905 542 1957
rect 594 1905 606 1957
rect 658 1905 671 1957
rect 530 1892 671 1905
rect 530 1840 542 1892
rect 594 1840 606 1892
rect 658 1840 671 1892
rect 530 1827 671 1840
rect 530 1775 542 1827
rect 594 1775 606 1827
rect 658 1775 671 1827
rect 530 1762 671 1775
rect 530 1710 542 1762
rect 594 1710 606 1762
rect 658 1710 671 1762
rect 530 1697 671 1710
rect 530 1645 542 1697
rect 594 1645 606 1697
rect 658 1645 671 1697
rect 530 1632 671 1645
rect 530 1580 542 1632
rect 594 1580 606 1632
rect 658 1580 671 1632
rect 530 1567 671 1580
rect 530 1515 542 1567
rect 594 1515 606 1567
rect 658 1515 671 1567
rect 530 1502 671 1515
rect 530 1450 542 1502
rect 594 1450 606 1502
rect 658 1450 671 1502
rect 530 1437 671 1450
rect 530 1385 542 1437
rect 594 1385 606 1437
rect 658 1385 671 1437
rect 530 1372 671 1385
rect 530 1320 542 1372
rect 594 1320 606 1372
rect 658 1320 671 1372
rect 530 1307 671 1320
rect 530 1255 542 1307
rect 594 1255 606 1307
rect 658 1255 671 1307
rect 530 1242 671 1255
rect 530 1190 542 1242
rect 594 1190 606 1242
rect 658 1190 671 1242
rect 530 1177 671 1190
rect 530 1125 542 1177
rect 594 1125 606 1177
rect 658 1125 671 1177
rect 530 1112 671 1125
rect 530 1060 542 1112
rect 594 1060 606 1112
rect 658 1060 671 1112
rect 530 1047 671 1060
rect 530 995 542 1047
rect 594 995 606 1047
rect 658 995 671 1047
rect 530 982 671 995
rect 530 930 542 982
rect 594 930 606 982
rect 658 930 671 982
rect 530 917 671 930
rect 530 865 542 917
rect 594 865 606 917
rect 658 865 671 917
rect 530 852 671 865
rect 530 800 542 852
rect 594 800 606 852
rect 658 800 671 852
rect 530 787 671 800
rect 530 735 542 787
rect 594 735 606 787
rect 658 735 671 787
rect 530 722 671 735
rect 530 670 542 722
rect 594 670 606 722
rect 658 670 671 722
rect 530 657 671 670
rect 530 605 542 657
rect 594 605 606 657
rect 658 605 671 657
rect 530 592 671 605
rect 530 540 542 592
rect 594 540 606 592
rect 658 540 671 592
rect 530 527 671 540
rect 530 475 542 527
rect 594 475 606 527
rect 658 475 671 527
rect 530 462 671 475
rect 530 410 542 462
rect 594 410 606 462
rect 658 410 671 462
rect 530 397 671 410
rect 530 345 542 397
rect 594 345 606 397
rect 658 345 671 397
rect 530 332 671 345
rect 530 280 542 332
rect 594 280 606 332
rect 658 280 671 332
rect 530 267 671 280
rect 530 215 542 267
rect 594 215 606 267
rect 658 215 671 267
rect 728 3949 820 4001
rect 872 3949 884 4001
rect 936 3949 948 4001
rect 1000 3949 1367 4001
rect 728 3935 1367 3949
rect 728 3883 820 3935
rect 872 3883 884 3935
rect 936 3883 948 3935
rect 1000 3883 1367 3935
rect 728 3869 1367 3883
rect 728 3817 820 3869
rect 872 3817 884 3869
rect 936 3817 948 3869
rect 1000 3817 1367 3869
rect 728 3803 1367 3817
rect 728 3751 820 3803
rect 872 3751 884 3803
rect 936 3751 948 3803
rect 1000 3751 1367 3803
rect 728 3737 1367 3751
rect 728 3685 820 3737
rect 872 3685 884 3737
rect 936 3685 948 3737
rect 1000 3685 1367 3737
rect 728 3671 1367 3685
rect 728 3619 820 3671
rect 872 3619 884 3671
rect 936 3619 948 3671
rect 1000 3619 1367 3671
rect 728 3605 1367 3619
rect 728 3553 820 3605
rect 872 3553 884 3605
rect 936 3553 948 3605
rect 1000 3553 1367 3605
rect 728 3539 1367 3553
rect 728 3487 820 3539
rect 872 3487 884 3539
rect 936 3487 948 3539
rect 1000 3487 1367 3539
rect 728 3474 1367 3487
rect 728 3422 820 3474
rect 872 3422 884 3474
rect 936 3422 948 3474
rect 1000 3422 1367 3474
rect 728 3409 1367 3422
rect 728 3357 820 3409
rect 872 3357 884 3409
rect 936 3357 948 3409
rect 1000 3357 1367 3409
rect 728 3344 1367 3357
rect 728 3292 820 3344
rect 872 3292 884 3344
rect 936 3292 948 3344
rect 1000 3292 1367 3344
rect 728 3279 1367 3292
rect 728 3227 820 3279
rect 872 3227 884 3279
rect 936 3227 948 3279
rect 1000 3227 1367 3279
rect 728 3214 1367 3227
rect 728 3162 820 3214
rect 872 3162 884 3214
rect 936 3162 948 3214
rect 1000 3162 1367 3214
rect 728 3149 1367 3162
rect 728 3097 820 3149
rect 872 3097 884 3149
rect 936 3097 948 3149
rect 1000 3097 1367 3149
rect 728 3084 1367 3097
rect 728 3032 820 3084
rect 872 3032 884 3084
rect 936 3032 948 3084
rect 1000 3032 1367 3084
rect 728 3019 1367 3032
rect 728 2967 820 3019
rect 872 2967 884 3019
rect 936 2967 948 3019
rect 1000 2967 1367 3019
rect 728 2954 1367 2967
rect 728 2902 820 2954
rect 872 2902 884 2954
rect 936 2902 948 2954
rect 1000 2902 1367 2954
rect 728 2889 1367 2902
rect 728 2837 820 2889
rect 872 2837 884 2889
rect 936 2837 948 2889
rect 1000 2837 1367 2889
rect 728 2824 1367 2837
rect 728 2772 820 2824
rect 872 2772 884 2824
rect 936 2772 948 2824
rect 1000 2772 1367 2824
rect 728 2759 1367 2772
rect 728 2707 820 2759
rect 872 2707 884 2759
rect 936 2707 948 2759
rect 1000 2707 1367 2759
rect 728 2694 1367 2707
rect 728 2642 820 2694
rect 872 2642 884 2694
rect 936 2642 948 2694
rect 1000 2642 1367 2694
rect 728 2286 1367 2642
rect 728 2234 820 2286
rect 872 2234 884 2286
rect 936 2234 948 2286
rect 1000 2234 1367 2286
rect 728 2221 1367 2234
rect 728 2169 820 2221
rect 872 2169 884 2221
rect 936 2169 948 2221
rect 1000 2169 1367 2221
rect 728 2156 1367 2169
rect 728 2104 820 2156
rect 872 2104 884 2156
rect 936 2104 948 2156
rect 1000 2104 1367 2156
rect 728 2091 1367 2104
rect 728 2039 820 2091
rect 872 2039 884 2091
rect 936 2039 948 2091
rect 1000 2039 1367 2091
rect 728 2026 1367 2039
rect 728 1974 820 2026
rect 872 1974 884 2026
rect 936 1974 948 2026
rect 1000 1974 1367 2026
rect 728 1961 1367 1974
rect 728 1909 820 1961
rect 872 1909 884 1961
rect 936 1909 948 1961
rect 1000 1909 1367 1961
rect 728 1896 1367 1909
rect 728 1844 820 1896
rect 872 1844 884 1896
rect 936 1844 948 1896
rect 1000 1844 1367 1896
rect 728 1831 1367 1844
rect 728 1779 820 1831
rect 872 1779 884 1831
rect 936 1779 948 1831
rect 1000 1779 1367 1831
rect 728 1766 1367 1779
rect 728 1714 820 1766
rect 872 1714 884 1766
rect 936 1714 948 1766
rect 1000 1714 1367 1766
rect 728 1701 1367 1714
rect 728 1649 820 1701
rect 872 1649 884 1701
rect 936 1649 948 1701
rect 1000 1649 1367 1701
rect 728 1636 1367 1649
rect 728 1584 820 1636
rect 872 1584 884 1636
rect 936 1584 948 1636
rect 1000 1584 1367 1636
rect 728 1571 1367 1584
rect 728 1519 820 1571
rect 872 1519 884 1571
rect 936 1519 948 1571
rect 1000 1519 1367 1571
rect 728 1506 1367 1519
rect 728 1454 820 1506
rect 872 1454 884 1506
rect 936 1454 948 1506
rect 1000 1454 1367 1506
rect 728 1441 1367 1454
rect 728 1389 820 1441
rect 872 1389 884 1441
rect 936 1389 948 1441
rect 1000 1389 1367 1441
rect 728 1376 1367 1389
rect 728 364 820 1376
rect 1000 557 1367 1376
rect 1423 4294 1539 4360
rect 1423 4242 1424 4294
rect 1476 4242 1539 4294
rect 1423 4229 1539 4242
rect 1423 4177 1424 4229
rect 1476 4177 1539 4229
rect 1423 4164 1539 4177
rect 1423 4112 1424 4164
rect 1476 4112 1539 4164
rect 1423 4099 1539 4112
rect 1423 4047 1424 4099
rect 1476 4047 1539 4099
rect 1423 4034 1539 4047
rect 1423 3982 1424 4034
rect 1476 3982 1539 4034
rect 1423 3969 1539 3982
rect 1423 3917 1424 3969
rect 1476 3917 1539 3969
rect 1423 3904 1539 3917
rect 1423 3852 1424 3904
rect 1476 3852 1539 3904
rect 1423 3839 1539 3852
rect 1423 3787 1424 3839
rect 1476 3787 1539 3839
rect 1423 3774 1539 3787
rect 1423 3722 1424 3774
rect 1476 3722 1539 3774
rect 1423 3709 1539 3722
rect 1423 3657 1424 3709
rect 1476 3657 1539 3709
rect 1423 3644 1539 3657
rect 1423 3592 1424 3644
rect 1476 3592 1539 3644
rect 1423 3579 1539 3592
rect 1423 3527 1424 3579
rect 1476 3527 1539 3579
rect 1423 3514 1539 3527
rect 1423 3462 1424 3514
rect 1476 3462 1539 3514
rect 1423 3449 1539 3462
rect 1423 3397 1424 3449
rect 1476 3397 1539 3449
rect 1423 3384 1539 3397
rect 1423 3332 1424 3384
rect 1476 3332 1539 3384
rect 1423 3319 1539 3332
rect 1423 3267 1424 3319
rect 1476 3267 1539 3319
rect 1423 3254 1539 3267
rect 1423 3202 1424 3254
rect 1476 3202 1539 3254
rect 1423 3189 1539 3202
rect 1423 3137 1424 3189
rect 1476 3137 1539 3189
rect 1423 3124 1539 3137
rect 1423 3072 1424 3124
rect 1476 3072 1539 3124
rect 1423 3059 1539 3072
rect 1423 3007 1424 3059
rect 1476 3007 1539 3059
rect 1423 2995 1539 3007
rect 1423 2943 1424 2995
rect 1476 2943 1539 2995
rect 1423 2931 1539 2943
rect 1423 2879 1424 2931
rect 1476 2879 1539 2931
rect 1423 2867 1539 2879
rect 1423 2815 1424 2867
rect 1476 2815 1539 2867
rect 1423 2803 1539 2815
rect 1423 2751 1424 2803
rect 1476 2751 1539 2803
rect 1423 2739 1539 2751
rect 1423 2687 1424 2739
rect 1476 2687 1539 2739
rect 1423 2675 1539 2687
rect 1423 2623 1424 2675
rect 1476 2623 1539 2675
rect 1423 2286 1539 2623
rect 1475 2234 1539 2286
rect 1423 2221 1539 2234
rect 1475 2169 1539 2221
rect 1423 2156 1539 2169
rect 1475 2104 1539 2156
rect 1423 2091 1539 2104
rect 1475 2039 1539 2091
rect 1423 2026 1539 2039
rect 1475 1974 1539 2026
rect 1423 1961 1539 1974
rect 1475 1909 1539 1961
rect 1423 1896 1539 1909
rect 1475 1844 1539 1896
rect 1423 1831 1539 1844
rect 1475 1779 1539 1831
rect 1423 1766 1539 1779
rect 1475 1714 1539 1766
rect 1423 1701 1539 1714
rect 1475 1649 1539 1701
rect 1423 1636 1539 1649
rect 1475 1584 1539 1636
rect 1423 1571 1539 1584
rect 1475 1519 1539 1571
rect 1423 1506 1539 1519
rect 1475 1454 1539 1506
rect 1423 1441 1539 1454
rect 1475 1389 1539 1441
rect 1423 1376 1539 1389
rect 1475 1324 1539 1376
rect 1423 1311 1539 1324
rect 1475 1259 1539 1311
rect 1423 1246 1539 1259
rect 1475 1194 1539 1246
rect 1423 1181 1539 1194
rect 1475 1129 1539 1181
rect 1423 1116 1539 1129
rect 1475 1064 1539 1116
rect 1423 1051 1539 1064
rect 1475 999 1539 1051
rect 1423 987 1539 999
rect 1475 935 1539 987
rect 1423 923 1539 935
rect 1475 871 1539 923
rect 1423 859 1539 871
rect 1475 807 1539 859
rect 1423 795 1539 807
rect 1475 743 1539 795
rect 1423 731 1539 743
rect 1475 679 1539 731
rect 1423 667 1539 679
rect 1475 615 1539 667
rect 1423 606 1539 615
rect 1567 4544 1715 4554
rect 1567 4492 1581 4544
rect 1633 4492 1645 4544
rect 1697 4492 1715 4544
rect 1567 4478 1715 4492
rect 1567 4426 1581 4478
rect 1633 4426 1645 4478
rect 1697 4426 1715 4478
rect 1567 4412 1715 4426
rect 1567 4360 1581 4412
rect 1633 4360 1645 4412
rect 1697 4360 1715 4412
rect 1567 4346 1715 4360
rect 1567 4294 1581 4346
rect 1633 4294 1645 4346
rect 1697 4294 1715 4346
rect 1567 4280 1715 4294
rect 1567 4228 1581 4280
rect 1633 4228 1645 4280
rect 1697 4228 1715 4280
rect 1567 4214 1715 4228
rect 1567 4162 1581 4214
rect 1633 4162 1645 4214
rect 1697 4162 1715 4214
rect 1567 4148 1715 4162
rect 1567 4096 1581 4148
rect 1633 4096 1645 4148
rect 1697 4096 1715 4148
rect 1567 4082 1715 4096
rect 1567 4030 1581 4082
rect 1633 4030 1645 4082
rect 1697 4030 1715 4082
rect 1567 4016 1715 4030
rect 1567 3964 1581 4016
rect 1633 3964 1645 4016
rect 1697 3964 1715 4016
rect 1567 3950 1715 3964
rect 1567 3898 1581 3950
rect 1633 3898 1645 3950
rect 1697 3898 1715 3950
rect 1567 3884 1715 3898
rect 1567 3832 1581 3884
rect 1633 3832 1645 3884
rect 1697 3832 1715 3884
rect 1567 3818 1715 3832
rect 1567 3766 1581 3818
rect 1633 3766 1645 3818
rect 1697 3766 1715 3818
rect 1567 3752 1715 3766
rect 1567 3700 1581 3752
rect 1633 3700 1645 3752
rect 1697 3700 1715 3752
rect 1567 3686 1715 3700
rect 1567 3634 1581 3686
rect 1633 3634 1645 3686
rect 1697 3634 1715 3686
rect 1567 3620 1715 3634
rect 1567 3568 1581 3620
rect 1633 3568 1645 3620
rect 1697 3568 1715 3620
rect 1567 3555 1715 3568
rect 1567 3503 1581 3555
rect 1633 3503 1645 3555
rect 1697 3503 1715 3555
rect 1567 3490 1715 3503
rect 1567 3438 1581 3490
rect 1633 3438 1645 3490
rect 1697 3438 1715 3490
rect 1567 3425 1715 3438
rect 1567 3373 1581 3425
rect 1633 3373 1645 3425
rect 1697 3373 1715 3425
rect 1567 3360 1715 3373
rect 1567 3308 1581 3360
rect 1633 3308 1645 3360
rect 1697 3308 1715 3360
rect 1567 3295 1715 3308
rect 1567 3243 1581 3295
rect 1633 3243 1645 3295
rect 1697 3243 1715 3295
rect 1567 3230 1715 3243
rect 1567 3178 1581 3230
rect 1633 3178 1645 3230
rect 1697 3178 1715 3230
rect 1567 3165 1715 3178
rect 1567 3113 1581 3165
rect 1633 3113 1645 3165
rect 1697 3113 1715 3165
rect 1567 3100 1715 3113
rect 1567 3048 1581 3100
rect 1633 3048 1645 3100
rect 1697 3048 1715 3100
rect 1567 3035 1715 3048
rect 1567 2983 1581 3035
rect 1633 2983 1645 3035
rect 1697 2983 1715 3035
rect 1567 2970 1715 2983
rect 1567 2918 1581 2970
rect 1633 2918 1645 2970
rect 1697 2918 1715 2970
rect 1567 1979 1715 2918
rect 1567 1927 1581 1979
rect 1633 1927 1645 1979
rect 1697 1927 1715 1979
rect 1567 1914 1715 1927
rect 1567 1862 1581 1914
rect 1633 1862 1645 1914
rect 1697 1862 1715 1914
rect 1567 1849 1715 1862
rect 1567 1797 1581 1849
rect 1633 1797 1645 1849
rect 1697 1797 1715 1849
rect 1567 1784 1715 1797
rect 1567 1732 1581 1784
rect 1633 1732 1645 1784
rect 1697 1732 1715 1784
rect 1567 1719 1715 1732
rect 1567 1667 1581 1719
rect 1633 1667 1645 1719
rect 1697 1667 1715 1719
rect 1567 1654 1715 1667
rect 1567 1602 1581 1654
rect 1633 1602 1645 1654
rect 1697 1602 1715 1654
rect 1567 1589 1715 1602
rect 1567 1537 1581 1589
rect 1633 1537 1645 1589
rect 1697 1537 1715 1589
rect 1567 1524 1715 1537
rect 1567 1472 1581 1524
rect 1633 1472 1645 1524
rect 1697 1472 1715 1524
rect 1567 1459 1715 1472
rect 1567 1407 1581 1459
rect 1633 1407 1645 1459
rect 1697 1407 1715 1459
rect 1567 1394 1715 1407
rect 1567 1342 1581 1394
rect 1633 1342 1645 1394
rect 1697 1342 1715 1394
rect 1567 1329 1715 1342
rect 1567 1277 1581 1329
rect 1633 1277 1645 1329
rect 1697 1277 1715 1329
rect 1567 1264 1715 1277
rect 1567 1212 1581 1264
rect 1633 1212 1645 1264
rect 1697 1212 1715 1264
rect 1567 1199 1715 1212
rect 1567 1147 1581 1199
rect 1633 1147 1645 1199
rect 1697 1147 1715 1199
rect 1567 1134 1715 1147
rect 1567 1082 1581 1134
rect 1633 1082 1645 1134
rect 1697 1082 1715 1134
rect 1567 1069 1715 1082
rect 1567 1017 1581 1069
rect 1633 1017 1645 1069
rect 1697 1017 1715 1069
rect 1567 1004 1715 1017
rect 1567 952 1581 1004
rect 1633 952 1645 1004
rect 1697 952 1715 1004
rect 1567 939 1715 952
rect 1567 887 1581 939
rect 1633 887 1645 939
rect 1697 887 1715 939
rect 1567 874 1715 887
rect 1567 822 1581 874
rect 1633 822 1645 874
rect 1697 822 1715 874
rect 1567 809 1715 822
rect 1000 505 1184 557
rect 1236 505 1248 557
rect 1300 505 1367 557
rect 1000 488 1367 505
rect 1000 436 1184 488
rect 1236 436 1248 488
rect 1300 436 1367 488
rect 1000 419 1367 436
rect 1000 367 1184 419
rect 1236 367 1248 419
rect 1300 367 1367 419
rect 1000 364 1367 367
rect 728 350 1367 364
rect 728 298 1184 350
rect 1236 298 1248 350
rect 1300 298 1367 350
rect 728 294 1367 298
tri 728 249 773 294 ne
rect 773 249 1367 294
rect 1567 373 1581 809
rect 1697 373 1715 809
tri 1367 249 1410 292 sw
tri 1542 249 1567 274 se
rect 1567 249 1715 373
rect 530 202 671 215
rect 530 150 542 202
rect 594 150 606 202
rect 658 150 671 202
tri 773 195 827 249 ne
rect 827 195 1715 249
rect 1743 4511 1861 4563
rect 1913 4511 1925 4563
rect 1977 4511 2040 4563
rect 1743 4498 2040 4511
rect 1743 4446 1861 4498
rect 1913 4446 1925 4498
rect 1977 4446 2040 4498
rect 1743 4433 2040 4446
rect 1743 4381 1861 4433
rect 1913 4381 1925 4433
rect 1977 4381 2040 4433
rect 1743 4368 2040 4381
rect 1743 4316 1861 4368
rect 1913 4316 1925 4368
rect 1977 4316 2040 4368
rect 1743 4303 2040 4316
rect 1743 4251 1861 4303
rect 1913 4251 1925 4303
rect 1977 4251 2040 4303
rect 1743 4238 2040 4251
rect 1743 4186 1861 4238
rect 1913 4186 1925 4238
rect 1977 4186 2040 4238
rect 1743 4173 2040 4186
rect 1743 4121 1861 4173
rect 1913 4121 1925 4173
rect 1977 4121 2040 4173
rect 1743 4108 2040 4121
rect 1743 4056 1861 4108
rect 1913 4056 1925 4108
rect 1977 4056 2040 4108
rect 1743 4043 2040 4056
rect 1743 3991 1861 4043
rect 1913 3991 1925 4043
rect 1977 3991 2040 4043
rect 1743 3978 2040 3991
rect 1743 3926 1861 3978
rect 1913 3926 1925 3978
rect 1977 3926 2040 3978
rect 1743 3913 2040 3926
rect 1743 3861 1861 3913
rect 1913 3861 1925 3913
rect 1977 3861 2040 3913
rect 1743 3848 2040 3861
rect 1743 3796 1861 3848
rect 1913 3796 1925 3848
rect 1977 3796 2040 3848
rect 1743 3783 2040 3796
rect 1743 3731 1861 3783
rect 1913 3731 1925 3783
rect 1977 3731 2040 3783
rect 1743 3718 2040 3731
rect 1743 3666 1861 3718
rect 1913 3666 1925 3718
rect 1977 3666 2040 3718
rect 1743 3653 2040 3666
rect 1743 3601 1861 3653
rect 1913 3601 1925 3653
rect 1977 3601 2040 3653
rect 1743 3588 2040 3601
rect 1743 3536 1861 3588
rect 1913 3536 1925 3588
rect 1977 3536 2040 3588
rect 1743 3523 2040 3536
rect 1743 3471 1861 3523
rect 1913 3471 1925 3523
rect 1977 3471 2040 3523
rect 1743 3458 2040 3471
rect 1743 3406 1861 3458
rect 1913 3406 1925 3458
rect 1977 3406 2040 3458
rect 1743 3393 2040 3406
rect 1743 3341 1861 3393
rect 1913 3341 1925 3393
rect 1977 3341 2040 3393
rect 1743 3328 2040 3341
rect 1743 3276 1861 3328
rect 1913 3276 1925 3328
rect 1977 3276 2040 3328
rect 1743 3263 2040 3276
rect 1743 3211 1861 3263
rect 1913 3211 1925 3263
rect 1977 3211 2040 3263
rect 1743 3198 2040 3211
rect 1743 3146 1861 3198
rect 1913 3146 1925 3198
rect 1977 3146 2040 3198
rect 1743 3133 2040 3146
rect 1743 3081 1861 3133
rect 1913 3081 1925 3133
rect 1977 3081 2040 3133
rect 1743 3068 2040 3081
rect 1743 2696 1861 3068
rect 1977 2696 2040 3068
rect 1743 2203 2040 2696
rect 1743 2151 1861 2203
rect 1913 2151 1925 2203
rect 1977 2151 2040 2203
rect 1743 2138 2040 2151
rect 1743 2086 1861 2138
rect 1913 2086 1925 2138
rect 1977 2086 2040 2138
rect 1743 2073 2040 2086
rect 1743 2021 1861 2073
rect 1913 2021 1925 2073
rect 1977 2021 2040 2073
rect 1743 2008 2040 2021
rect 1743 1956 1861 2008
rect 1913 1956 1925 2008
rect 1977 1956 2040 2008
rect 1743 1943 2040 1956
rect 1743 1891 1861 1943
rect 1913 1891 1925 1943
rect 1977 1891 2040 1943
rect 1743 1878 2040 1891
rect 1743 1826 1861 1878
rect 1913 1826 1925 1878
rect 1977 1826 2040 1878
rect 1743 1813 2040 1826
rect 1743 1761 1861 1813
rect 1913 1761 1925 1813
rect 1977 1761 2040 1813
rect 1743 1748 2040 1761
rect 1743 1696 1861 1748
rect 1913 1696 1925 1748
rect 1977 1696 2040 1748
rect 1743 1683 2040 1696
rect 1743 1631 1861 1683
rect 1913 1631 1925 1683
rect 1977 1631 2040 1683
rect 1743 1618 2040 1631
rect 1743 1566 1861 1618
rect 1913 1566 1925 1618
rect 1977 1566 2040 1618
rect 1743 1553 2040 1566
rect 1743 1501 1861 1553
rect 1913 1501 1925 1553
rect 1977 1501 2040 1553
rect 1743 1488 2040 1501
rect 1743 1436 1861 1488
rect 1913 1436 1925 1488
rect 1977 1436 2040 1488
rect 1743 1423 2040 1436
rect 1743 1371 1861 1423
rect 1913 1371 1925 1423
rect 1977 1371 2040 1423
rect 1743 1358 2040 1371
rect 1743 1306 1861 1358
rect 1913 1306 1925 1358
rect 1977 1306 2040 1358
rect 1743 1293 2040 1306
rect 1743 1241 1861 1293
rect 1913 1241 1925 1293
rect 1977 1241 2040 1293
rect 1743 1228 2040 1241
rect 1743 1176 1861 1228
rect 1913 1176 1925 1228
rect 1977 1176 2040 1228
rect 1743 1163 2040 1176
rect 1743 1111 1861 1163
rect 1913 1111 1925 1163
rect 1977 1111 2040 1163
rect 1743 1098 2040 1111
rect 1743 1046 1861 1098
rect 1913 1046 1925 1098
rect 1977 1046 2040 1098
rect 1743 1033 2040 1046
rect 1743 981 1861 1033
rect 1913 981 1925 1033
rect 1977 981 2040 1033
rect 1743 968 2040 981
rect 1743 916 1861 968
rect 1913 916 1925 968
rect 1977 916 2040 968
rect 1743 903 2040 916
rect 1743 851 1861 903
rect 1913 851 1925 903
rect 1977 851 2040 903
rect 1743 838 2040 851
rect 1743 786 1861 838
rect 1913 786 1925 838
rect 1977 786 2040 838
rect 1743 773 2040 786
rect 1743 721 1861 773
rect 1913 721 1925 773
rect 1977 721 2040 773
rect 1743 708 2040 721
rect 530 144 671 150
tri 671 144 689 162 sw
tri 1725 144 1743 162 se
rect 1743 144 1861 708
rect 530 137 689 144
tri 689 137 696 144 sw
tri 1718 137 1725 144 se
rect 1725 137 1861 144
rect 530 128 1861 137
rect 530 76 673 128
rect 725 76 740 128
rect 792 76 807 128
rect 859 76 874 128
rect 926 76 941 128
rect 993 76 1008 128
rect 1060 76 1075 128
rect 1127 76 1356 128
rect 1408 76 1423 128
rect 1475 76 1490 128
rect 1542 76 1557 128
rect 1609 76 1624 128
rect 1676 76 1691 128
rect 1743 76 1758 128
rect 1810 80 1861 128
rect 1977 158 2040 708
rect 2068 4595 2388 4616
rect 2068 4543 2236 4595
rect 2288 4543 2330 4595
rect 2382 4543 2388 4595
rect 2068 4542 2388 4543
rect 2068 4490 2153 4542
rect 2205 4531 2388 4542
rect 2205 4520 2311 4531
rect 2205 4490 2217 4520
rect 2068 4476 2217 4490
rect 2068 4424 2153 4476
rect 2205 4468 2217 4476
rect 2269 4479 2311 4520
rect 2363 4479 2388 4531
rect 2269 4468 2388 4479
rect 2205 4455 2388 4468
rect 2205 4424 2217 4455
rect 2068 4410 2217 4424
rect 2068 4358 2153 4410
rect 2205 4403 2217 4410
rect 2269 4403 2388 4455
rect 2205 4390 2388 4403
rect 2205 4358 2217 4390
rect 2068 4344 2217 4358
rect 2068 4292 2153 4344
rect 2205 4338 2217 4344
rect 2269 4338 2388 4390
rect 2205 4325 2388 4338
rect 2205 4292 2217 4325
rect 2068 4278 2217 4292
rect 2068 4226 2153 4278
rect 2205 4273 2217 4278
rect 2269 4273 2388 4325
rect 2205 4260 2388 4273
rect 2205 4226 2217 4260
rect 2068 4212 2217 4226
rect 2068 4160 2153 4212
rect 2205 4208 2217 4212
rect 2269 4208 2388 4260
rect 2205 4195 2388 4208
rect 2205 4160 2217 4195
rect 2068 4146 2217 4160
rect 2068 4094 2153 4146
rect 2205 4143 2217 4146
rect 2269 4143 2388 4195
rect 2205 4130 2388 4143
rect 2205 4094 2217 4130
rect 2068 4080 2217 4094
rect 2068 4028 2153 4080
rect 2205 4078 2217 4080
rect 2269 4078 2388 4130
rect 2205 4065 2388 4078
rect 2205 4028 2217 4065
rect 2068 4014 2217 4028
rect 2068 3962 2153 4014
rect 2205 4013 2217 4014
rect 2269 4013 2388 4065
rect 2205 4000 2388 4013
rect 2205 3962 2217 4000
rect 2068 3948 2217 3962
rect 2269 3948 2388 4000
rect 2068 3896 2153 3948
rect 2205 3935 2388 3948
rect 2205 3896 2217 3935
rect 2068 3883 2217 3896
rect 2269 3883 2388 3935
rect 2068 3882 2388 3883
rect 2068 3830 2153 3882
rect 2205 3870 2388 3882
rect 2205 3830 2217 3870
rect 2068 3818 2217 3830
rect 2269 3818 2388 3870
rect 2068 3816 2388 3818
rect 2068 3764 2153 3816
rect 2205 3805 2388 3816
rect 2205 3764 2217 3805
rect 2068 3753 2217 3764
rect 2269 3753 2388 3805
rect 2068 3750 2388 3753
rect 2068 3698 2153 3750
rect 2205 3740 2388 3750
rect 2205 3698 2217 3740
rect 2068 3688 2217 3698
rect 2269 3688 2388 3740
rect 2068 3685 2388 3688
rect 2068 3633 2153 3685
rect 2205 3675 2388 3685
rect 2205 3633 2217 3675
rect 2068 3623 2217 3633
rect 2269 3623 2388 3675
rect 2068 3620 2388 3623
rect 2068 3568 2153 3620
rect 2205 3610 2388 3620
rect 2205 3568 2217 3610
rect 2068 3558 2217 3568
rect 2269 3558 2388 3610
rect 2068 3555 2388 3558
rect 2068 3503 2153 3555
rect 2205 3546 2388 3555
rect 2205 3503 2217 3546
rect 2068 3494 2217 3503
rect 2269 3494 2388 3546
rect 2068 3490 2388 3494
rect 2068 3438 2153 3490
rect 2205 3482 2388 3490
rect 2205 3438 2217 3482
rect 2068 3430 2217 3438
rect 2269 3430 2388 3482
rect 2068 3425 2388 3430
rect 2068 3373 2153 3425
rect 2205 3418 2388 3425
rect 2205 3373 2217 3418
rect 2068 3366 2217 3373
rect 2269 3366 2388 3418
rect 2068 3360 2388 3366
rect 2068 3308 2153 3360
rect 2205 3354 2388 3360
rect 2205 3308 2217 3354
rect 2068 3302 2217 3308
rect 2269 3302 2388 3354
rect 2068 3295 2388 3302
rect 2068 3243 2153 3295
rect 2205 3290 2388 3295
rect 2205 3243 2217 3290
rect 2068 3238 2217 3243
rect 2269 3238 2388 3290
rect 2068 3230 2388 3238
rect 2068 3178 2153 3230
rect 2205 3226 2388 3230
rect 2205 3178 2217 3226
rect 2068 3174 2217 3178
rect 2269 3174 2388 3226
rect 2068 3165 2388 3174
rect 2068 3113 2153 3165
rect 2205 3162 2388 3165
rect 2205 3113 2217 3162
rect 2068 3110 2217 3113
rect 2269 3110 2388 3162
rect 2068 3100 2388 3110
rect 2068 3048 2153 3100
rect 2205 3098 2388 3100
rect 2205 3048 2217 3098
rect 2068 3046 2217 3048
rect 2269 3046 2388 3098
rect 2068 3035 2388 3046
rect 2068 2983 2153 3035
rect 2205 3034 2388 3035
rect 2205 2983 2217 3034
rect 2068 2982 2217 2983
rect 2269 2982 2388 3034
rect 2068 2970 2388 2982
rect 2068 2918 2153 2970
rect 2205 2918 2217 2970
rect 2269 2918 2388 2970
rect 2068 1990 2388 2918
rect 2068 1938 2153 1990
rect 2205 1938 2217 1990
rect 2269 1938 2388 1990
rect 2068 1926 2388 1938
rect 2068 1925 2217 1926
rect 2068 1873 2153 1925
rect 2205 1874 2217 1925
rect 2269 1874 2388 1926
rect 2205 1873 2388 1874
rect 2068 1862 2388 1873
rect 2068 1860 2217 1862
rect 2068 1808 2153 1860
rect 2205 1810 2217 1860
rect 2269 1810 2388 1862
rect 2205 1808 2388 1810
rect 2068 1798 2388 1808
rect 2068 1795 2217 1798
rect 2068 1743 2153 1795
rect 2205 1746 2217 1795
rect 2269 1746 2388 1798
rect 2205 1743 2388 1746
rect 2068 1734 2388 1743
rect 2068 1730 2217 1734
rect 2068 1678 2153 1730
rect 2205 1682 2217 1730
rect 2269 1682 2388 1734
rect 2205 1678 2388 1682
rect 2068 1670 2388 1678
rect 2068 1665 2217 1670
rect 2068 1613 2153 1665
rect 2205 1618 2217 1665
rect 2269 1618 2388 1670
rect 2205 1613 2388 1618
rect 2068 1606 2388 1613
rect 2068 1600 2217 1606
rect 2068 1548 2153 1600
rect 2205 1554 2217 1600
rect 2269 1554 2388 1606
rect 2205 1548 2388 1554
rect 2068 1542 2388 1548
rect 2068 1535 2217 1542
rect 2068 1483 2153 1535
rect 2205 1490 2217 1535
rect 2269 1490 2388 1542
rect 2205 1483 2388 1490
rect 2068 1478 2388 1483
rect 2068 1470 2217 1478
rect 2068 1418 2153 1470
rect 2205 1426 2217 1470
rect 2269 1426 2388 1478
rect 2205 1418 2388 1426
rect 2068 1414 2388 1418
rect 2068 1405 2217 1414
rect 2068 1353 2153 1405
rect 2205 1362 2217 1405
rect 2269 1362 2388 1414
rect 2205 1353 2388 1362
rect 2068 1350 2388 1353
rect 2068 1340 2217 1350
rect 2068 1288 2153 1340
rect 2205 1298 2217 1340
rect 2269 1298 2388 1350
rect 2205 1288 2388 1298
rect 2068 1285 2388 1288
rect 2068 1275 2217 1285
rect 2068 1223 2153 1275
rect 2205 1233 2217 1275
rect 2269 1233 2388 1285
rect 2205 1223 2388 1233
rect 2068 1220 2388 1223
rect 2068 1210 2217 1220
rect 2068 1158 2153 1210
rect 2205 1168 2217 1210
rect 2269 1168 2388 1220
rect 2205 1158 2388 1168
rect 2068 1155 2388 1158
rect 2068 1144 2217 1155
rect 2068 1092 2153 1144
rect 2205 1103 2217 1144
rect 2269 1103 2388 1155
rect 2205 1092 2388 1103
rect 2068 1090 2388 1092
rect 2068 1078 2217 1090
rect 2068 1026 2153 1078
rect 2205 1038 2217 1078
rect 2269 1038 2388 1090
rect 2205 1026 2388 1038
rect 2068 1025 2388 1026
rect 2068 1012 2217 1025
rect 2068 960 2153 1012
rect 2205 973 2217 1012
rect 2269 973 2388 1025
rect 2205 960 2388 973
rect 2068 946 2217 960
rect 2068 894 2153 946
rect 2205 908 2217 946
rect 2269 908 2388 960
rect 2205 895 2388 908
rect 2205 894 2217 895
rect 2068 880 2217 894
rect 2068 828 2153 880
rect 2205 843 2217 880
rect 2269 843 2388 895
rect 2205 830 2388 843
rect 2205 828 2217 830
rect 2068 814 2217 828
rect 2068 762 2153 814
rect 2205 778 2217 814
rect 2269 778 2388 830
rect 2205 765 2388 778
rect 2205 762 2217 765
rect 2068 748 2217 762
rect 2068 696 2153 748
rect 2205 713 2217 748
rect 2269 713 2388 765
rect 2205 700 2388 713
rect 2205 696 2217 700
rect 2068 682 2217 696
rect 2068 630 2153 682
rect 2205 648 2217 682
rect 2269 648 2388 700
rect 2205 635 2388 648
rect 2205 630 2217 635
rect 2068 616 2217 630
rect 2068 564 2153 616
rect 2205 583 2217 616
rect 2269 583 2388 635
rect 2205 570 2388 583
rect 2205 564 2217 570
rect 2068 550 2217 564
rect 2068 498 2153 550
rect 2205 518 2217 550
rect 2269 518 2388 570
rect 2205 505 2388 518
rect 2205 498 2217 505
rect 2068 484 2217 498
rect 2068 432 2153 484
rect 2205 453 2217 484
rect 2269 453 2388 505
rect 2205 440 2388 453
rect 2205 432 2217 440
rect 2068 418 2217 432
rect 2068 366 2153 418
rect 2205 388 2217 418
rect 2269 429 2388 440
rect 2269 388 2311 429
rect 2205 377 2311 388
rect 2363 377 2388 429
rect 2205 366 2388 377
rect 2068 365 2388 366
rect 2068 313 2236 365
rect 2288 313 2330 365
rect 2382 313 2388 365
rect 2068 267 2388 313
rect 2416 4584 2538 4636
rect 2590 4584 2602 4636
rect 2654 4584 2769 4636
rect 2416 4570 2769 4584
rect 2416 4518 2538 4570
rect 2590 4518 2602 4570
rect 2654 4518 2769 4570
rect 2416 4504 2769 4518
rect 2416 4452 2538 4504
rect 2590 4452 2602 4504
rect 2654 4452 2769 4504
rect 2416 4438 2769 4452
rect 2416 4386 2538 4438
rect 2590 4386 2602 4438
rect 2654 4386 2769 4438
rect 2416 4359 2769 4386
rect 2416 4307 2589 4359
rect 2641 4307 2653 4359
rect 2705 4307 2717 4359
rect 2416 4294 2769 4307
rect 2416 4242 2589 4294
rect 2641 4242 2653 4294
rect 2705 4242 2717 4294
rect 2416 4229 2769 4242
rect 2416 4177 2589 4229
rect 2641 4177 2653 4229
rect 2705 4177 2717 4229
rect 2416 4164 2769 4177
rect 2416 4112 2589 4164
rect 2641 4112 2653 4164
rect 2705 4112 2717 4164
rect 2416 4099 2769 4112
rect 2416 4047 2589 4099
rect 2641 4047 2653 4099
rect 2705 4047 2717 4099
rect 2416 4034 2769 4047
rect 2416 3982 2589 4034
rect 2641 3982 2653 4034
rect 2705 3982 2717 4034
rect 2416 3969 2769 3982
rect 2416 3917 2589 3969
rect 2641 3917 2653 3969
rect 2705 3917 2717 3969
rect 2416 3904 2769 3917
rect 2416 3852 2589 3904
rect 2641 3852 2653 3904
rect 2705 3852 2717 3904
rect 2416 3839 2769 3852
rect 2416 3787 2589 3839
rect 2641 3787 2653 3839
rect 2705 3787 2717 3839
rect 2416 3774 2769 3787
rect 2416 3722 2589 3774
rect 2641 3722 2653 3774
rect 2705 3722 2717 3774
rect 2416 3709 2769 3722
rect 2416 3657 2589 3709
rect 2641 3657 2653 3709
rect 2705 3657 2717 3709
rect 2416 3644 2769 3657
rect 2416 3592 2589 3644
rect 2641 3592 2653 3644
rect 2705 3592 2717 3644
rect 2416 3579 2769 3592
rect 2416 3527 2589 3579
rect 2641 3527 2653 3579
rect 2705 3527 2717 3579
rect 2416 3514 2769 3527
rect 2416 3462 2589 3514
rect 2641 3462 2653 3514
rect 2705 3462 2717 3514
rect 2416 3449 2769 3462
rect 2416 3397 2589 3449
rect 2641 3397 2653 3449
rect 2705 3397 2717 3449
rect 2416 3384 2769 3397
rect 2416 3332 2589 3384
rect 2641 3332 2653 3384
rect 2705 3332 2717 3384
rect 2416 3319 2769 3332
rect 2416 3267 2589 3319
rect 2641 3267 2653 3319
rect 2705 3267 2717 3319
rect 2416 3254 2769 3267
rect 2416 3202 2589 3254
rect 2641 3202 2653 3254
rect 2705 3202 2717 3254
rect 2416 3189 2769 3202
rect 2416 3137 2589 3189
rect 2641 3137 2653 3189
rect 2705 3137 2717 3189
rect 2416 3124 2769 3137
rect 2416 3072 2589 3124
rect 2641 3072 2653 3124
rect 2705 3072 2717 3124
rect 2416 3059 2769 3072
rect 2416 3007 2589 3059
rect 2641 3007 2653 3059
rect 2705 3007 2717 3059
rect 2416 2994 2769 3007
rect 2416 2622 2589 2994
rect 2416 2286 2769 2622
rect 2416 2234 2589 2286
rect 2641 2234 2653 2286
rect 2705 2234 2717 2286
rect 2416 2220 2769 2234
rect 2416 2168 2589 2220
rect 2641 2168 2653 2220
rect 2705 2168 2717 2220
rect 2416 2154 2769 2168
rect 2416 2102 2589 2154
rect 2641 2102 2653 2154
rect 2705 2102 2717 2154
rect 2416 2088 2769 2102
rect 2416 2036 2589 2088
rect 2641 2036 2653 2088
rect 2705 2036 2717 2088
rect 2416 2022 2769 2036
rect 2416 1970 2589 2022
rect 2641 1970 2653 2022
rect 2705 1970 2717 2022
rect 2416 1956 2769 1970
rect 2416 1904 2589 1956
rect 2641 1904 2653 1956
rect 2705 1904 2717 1956
rect 2416 1890 2769 1904
rect 2416 1838 2589 1890
rect 2641 1838 2653 1890
rect 2705 1838 2717 1890
rect 2416 1824 2769 1838
rect 2416 1772 2589 1824
rect 2641 1772 2653 1824
rect 2705 1772 2717 1824
rect 2416 1759 2769 1772
rect 2416 1707 2589 1759
rect 2641 1707 2653 1759
rect 2705 1707 2717 1759
rect 2416 1694 2769 1707
rect 2416 1642 2589 1694
rect 2641 1642 2653 1694
rect 2705 1642 2717 1694
rect 2416 1629 2769 1642
rect 2416 1577 2589 1629
rect 2641 1577 2653 1629
rect 2705 1577 2717 1629
rect 2416 1564 2769 1577
rect 2416 1512 2589 1564
rect 2641 1512 2653 1564
rect 2705 1512 2717 1564
rect 2416 1499 2769 1512
rect 2416 1447 2589 1499
rect 2641 1447 2653 1499
rect 2705 1447 2717 1499
rect 2416 1434 2769 1447
rect 2416 1382 2589 1434
rect 2641 1382 2653 1434
rect 2705 1382 2717 1434
rect 2416 1369 2769 1382
rect 2416 1317 2589 1369
rect 2641 1317 2653 1369
rect 2705 1317 2717 1369
rect 2416 1304 2769 1317
rect 2416 1252 2589 1304
rect 2641 1252 2653 1304
rect 2705 1252 2717 1304
rect 2416 1239 2769 1252
rect 2416 1187 2589 1239
rect 2641 1187 2653 1239
rect 2705 1187 2717 1239
rect 2416 1174 2769 1187
rect 2416 1122 2589 1174
rect 2641 1122 2653 1174
rect 2705 1122 2717 1174
rect 2416 1109 2769 1122
rect 2416 1057 2589 1109
rect 2641 1057 2653 1109
rect 2705 1057 2717 1109
rect 2416 1044 2769 1057
rect 2416 992 2589 1044
rect 2641 992 2653 1044
rect 2705 992 2717 1044
rect 2416 979 2769 992
rect 2416 927 2589 979
rect 2641 927 2653 979
rect 2705 927 2717 979
rect 2416 914 2769 927
rect 2416 862 2589 914
rect 2641 862 2653 914
rect 2705 862 2717 914
rect 2416 849 2769 862
rect 2416 797 2589 849
rect 2641 797 2653 849
rect 2705 797 2717 849
rect 2416 784 2769 797
rect 2416 732 2589 784
rect 2641 732 2653 784
rect 2705 732 2717 784
rect 2416 719 2769 732
rect 2416 667 2589 719
rect 2641 667 2653 719
rect 2705 667 2717 719
rect 2416 554 2769 667
rect 2416 502 2538 554
rect 2590 502 2602 554
rect 2654 502 2769 554
rect 2416 485 2769 502
rect 2416 433 2538 485
rect 2590 433 2602 485
rect 2654 433 2769 485
rect 2416 417 2769 433
rect 2416 365 2538 417
rect 2590 365 2602 417
rect 2654 365 2769 417
rect 2416 349 2769 365
rect 2416 297 2538 349
rect 2590 297 2602 349
rect 2654 297 2769 349
rect 2416 291 2769 297
rect 2797 4565 3117 5505
rect 3172 4945 3465 5253
tri 3172 4944 3173 4945 ne
rect 2797 4513 2876 4565
rect 2928 4513 2940 4565
rect 2992 4513 3117 4565
rect 2797 4500 3117 4513
rect 2797 4448 2876 4500
rect 2928 4448 2940 4500
rect 2992 4448 3117 4500
rect 2797 4435 3117 4448
rect 2797 4383 2876 4435
rect 2928 4383 2940 4435
rect 2992 4383 3117 4435
rect 2797 4370 3117 4383
rect 2797 4318 2876 4370
rect 2928 4318 2940 4370
rect 2992 4318 3117 4370
rect 2797 4305 3117 4318
rect 2797 4253 2876 4305
rect 2928 4253 2940 4305
rect 2992 4253 3117 4305
rect 2797 4240 3117 4253
rect 2797 4188 2876 4240
rect 2928 4188 2940 4240
rect 2992 4188 3117 4240
rect 2797 4175 3117 4188
rect 2797 4123 2876 4175
rect 2928 4123 2940 4175
rect 2992 4123 3117 4175
rect 2797 4110 3117 4123
rect 2797 4058 2876 4110
rect 2928 4058 2940 4110
rect 2992 4058 3117 4110
rect 2797 4045 3117 4058
rect 2797 3993 2876 4045
rect 2928 3993 2940 4045
rect 2992 3993 3117 4045
rect 2797 3980 3117 3993
rect 2797 3928 2876 3980
rect 2928 3928 2940 3980
rect 2992 3928 3117 3980
rect 2797 3915 3117 3928
rect 2797 3863 2876 3915
rect 2928 3863 2940 3915
rect 2992 3863 3117 3915
rect 2797 3850 3117 3863
rect 2797 3798 2876 3850
rect 2928 3798 2940 3850
rect 2992 3798 3117 3850
rect 2797 3785 3117 3798
rect 2797 3733 2876 3785
rect 2928 3733 2940 3785
rect 2992 3733 3117 3785
rect 2797 3720 3117 3733
rect 2797 3668 2876 3720
rect 2928 3668 2940 3720
rect 2992 3668 3117 3720
rect 2797 3655 3117 3668
rect 2797 3603 2876 3655
rect 2928 3603 2940 3655
rect 2992 3603 3117 3655
rect 2797 3590 3117 3603
rect 2797 3538 2876 3590
rect 2928 3538 2940 3590
rect 2992 3538 3117 3590
rect 2797 3525 3117 3538
rect 2797 3473 2876 3525
rect 2928 3473 2940 3525
rect 2992 3473 3117 3525
rect 2797 3460 3117 3473
rect 2797 3408 2876 3460
rect 2928 3408 2940 3460
rect 2992 3408 3117 3460
rect 2797 3395 3117 3408
rect 2797 3343 2876 3395
rect 2928 3343 2940 3395
rect 2992 3343 3117 3395
rect 2797 3330 3117 3343
rect 2797 2638 2876 3330
rect 2992 2638 3117 3330
rect 2797 2270 3117 2638
rect 2797 1578 2876 2270
rect 2992 1578 3117 2270
rect 2797 1565 3117 1578
rect 2797 1513 2876 1565
rect 2928 1513 2940 1565
rect 2992 1513 3117 1565
rect 2797 1500 3117 1513
rect 2797 1448 2876 1500
rect 2928 1448 2940 1500
rect 2992 1448 3117 1500
rect 2797 1435 3117 1448
rect 2797 1383 2876 1435
rect 2928 1383 2940 1435
rect 2992 1383 3117 1435
rect 2797 1370 3117 1383
rect 2797 1318 2876 1370
rect 2928 1318 2940 1370
rect 2992 1318 3117 1370
rect 2797 1305 3117 1318
rect 2797 1253 2876 1305
rect 2928 1253 2940 1305
rect 2992 1253 3117 1305
rect 2797 1240 3117 1253
rect 2797 1188 2876 1240
rect 2928 1188 2940 1240
rect 2992 1188 3117 1240
rect 2797 1175 3117 1188
rect 2797 1123 2876 1175
rect 2928 1123 2940 1175
rect 2992 1123 3117 1175
rect 2797 1110 3117 1123
rect 2797 1058 2876 1110
rect 2928 1058 2940 1110
rect 2992 1058 3117 1110
rect 2797 1045 3117 1058
rect 2797 993 2876 1045
rect 2928 993 2940 1045
rect 2992 993 3117 1045
rect 2797 980 3117 993
rect 2797 928 2876 980
rect 2928 928 2940 980
rect 2992 928 3117 980
rect 2797 915 3117 928
rect 2797 863 2876 915
rect 2928 863 2940 915
rect 2992 863 3117 915
rect 2797 850 3117 863
rect 2797 798 2876 850
rect 2928 798 2940 850
rect 2992 798 3117 850
rect 2797 785 3117 798
rect 2797 733 2876 785
rect 2928 733 2940 785
rect 2992 733 3117 785
rect 2797 720 3117 733
rect 2797 668 2876 720
rect 2928 668 2940 720
rect 2992 668 3117 720
rect 2797 655 3117 668
rect 2797 603 2876 655
rect 2928 603 2940 655
rect 2992 603 3117 655
rect 2797 590 3117 603
rect 2797 538 2876 590
rect 2928 538 2940 590
rect 2992 538 3117 590
rect 2797 525 3117 538
rect 2797 473 2876 525
rect 2928 473 2940 525
rect 2992 473 3117 525
rect 2797 460 3117 473
rect 2797 408 2876 460
rect 2928 408 2940 460
rect 2992 408 3117 460
rect 2797 395 3117 408
rect 2797 343 2876 395
rect 2928 343 2940 395
rect 2992 343 3117 395
tri 2388 267 2395 274 sw
tri 2790 267 2797 274 se
rect 2797 267 3117 343
rect 2068 249 2395 267
tri 2395 249 2413 267 sw
tri 2772 249 2790 267 se
rect 2790 249 3117 267
rect 2068 195 3117 249
rect 3173 4763 3465 4945
rect 3173 4711 3180 4763
rect 3232 4711 3244 4763
rect 3296 4711 3465 4763
rect 3173 4697 3465 4711
rect 3173 4645 3180 4697
rect 3232 4645 3244 4697
rect 3296 4645 3465 4697
rect 3173 4631 3465 4645
rect 3173 4579 3180 4631
rect 3232 4579 3244 4631
rect 3296 4579 3465 4631
rect 3173 4565 3465 4579
rect 3173 4513 3180 4565
rect 3232 4513 3244 4565
rect 3296 4513 3465 4565
rect 3173 4499 3465 4513
rect 3173 4447 3180 4499
rect 3232 4447 3244 4499
rect 3296 4447 3465 4499
rect 3173 4434 3465 4447
rect 3173 4382 3180 4434
rect 3232 4382 3244 4434
rect 3296 4382 3465 4434
rect 3173 4369 3465 4382
rect 3173 4317 3180 4369
rect 3232 4317 3244 4369
rect 3296 4317 3465 4369
rect 3173 4304 3465 4317
rect 3173 4252 3180 4304
rect 3232 4252 3244 4304
rect 3296 4252 3465 4304
rect 3173 4239 3465 4252
rect 3173 4187 3180 4239
rect 3232 4187 3244 4239
rect 3296 4187 3465 4239
rect 3173 4174 3465 4187
rect 3173 4122 3180 4174
rect 3232 4122 3244 4174
rect 3296 4122 3465 4174
rect 3173 4109 3465 4122
rect 3173 4057 3180 4109
rect 3232 4057 3244 4109
rect 3296 4057 3465 4109
rect 3173 4044 3465 4057
rect 3173 3992 3180 4044
rect 3232 3992 3244 4044
rect 3296 3992 3465 4044
rect 3173 3979 3465 3992
rect 3173 3927 3180 3979
rect 3232 3927 3244 3979
rect 3296 3927 3465 3979
rect 3173 3914 3465 3927
rect 3173 3862 3180 3914
rect 3232 3862 3244 3914
rect 3296 3862 3465 3914
rect 3173 3849 3465 3862
rect 3173 3797 3180 3849
rect 3232 3797 3244 3849
rect 3296 3797 3465 3849
rect 3173 3784 3465 3797
rect 3173 3732 3180 3784
rect 3232 3732 3244 3784
rect 3296 3732 3465 3784
rect 3173 3719 3465 3732
rect 3173 3667 3180 3719
rect 3232 3667 3244 3719
rect 3296 3667 3465 3719
rect 3173 3654 3465 3667
rect 3173 3602 3180 3654
rect 3232 3602 3244 3654
rect 3296 3602 3465 3654
rect 3173 3589 3465 3602
rect 3173 3537 3180 3589
rect 3232 3537 3244 3589
rect 3296 3537 3465 3589
rect 3173 3524 3465 3537
rect 3173 3472 3180 3524
rect 3232 3472 3244 3524
rect 3296 3472 3465 3524
rect 3173 3459 3465 3472
rect 3173 3407 3180 3459
rect 3232 3407 3244 3459
rect 3296 3407 3465 3459
rect 3173 3394 3465 3407
rect 3173 3342 3180 3394
rect 3232 3342 3244 3394
rect 3296 3342 3465 3394
rect 3173 3329 3465 3342
rect 3173 3277 3180 3329
rect 3232 3277 3244 3329
rect 3296 3277 3465 3329
rect 3173 3264 3465 3277
rect 3173 3212 3180 3264
rect 3232 3212 3244 3264
rect 3296 3212 3465 3264
rect 3173 3199 3465 3212
rect 3173 3147 3180 3199
rect 3232 3147 3244 3199
rect 3296 3147 3465 3199
rect 3173 3134 3465 3147
rect 3173 3082 3180 3134
rect 3232 3082 3244 3134
rect 3296 3082 3465 3134
rect 3173 3069 3465 3082
rect 3173 3017 3180 3069
rect 3232 3017 3244 3069
rect 3296 3017 3465 3069
rect 3173 3004 3465 3017
rect 3173 2952 3180 3004
rect 3232 2952 3244 3004
rect 3296 2952 3465 3004
rect 3173 2939 3465 2952
rect 3173 2887 3180 2939
rect 3232 2887 3244 2939
rect 3296 2887 3465 2939
rect 3173 2874 3465 2887
rect 3173 2822 3180 2874
rect 3232 2822 3244 2874
rect 3296 2822 3465 2874
rect 3173 2809 3465 2822
rect 3173 2757 3180 2809
rect 3232 2757 3244 2809
rect 3296 2757 3465 2809
rect 3173 2744 3465 2757
rect 3173 2692 3180 2744
rect 3232 2692 3244 2744
rect 3296 2692 3465 2744
rect 3173 2679 3465 2692
rect 3173 2627 3180 2679
rect 3232 2627 3244 2679
rect 3296 2627 3465 2679
rect 3173 2286 3465 2627
rect 3173 2234 3180 2286
rect 3232 2234 3244 2286
rect 3296 2234 3465 2286
rect 3173 2220 3465 2234
rect 3173 2168 3180 2220
rect 3232 2168 3244 2220
rect 3296 2168 3465 2220
rect 3173 2154 3465 2168
rect 3173 2102 3180 2154
rect 3232 2102 3244 2154
rect 3296 2102 3465 2154
rect 3173 2088 3465 2102
rect 3173 2036 3180 2088
rect 3232 2036 3244 2088
rect 3296 2036 3465 2088
rect 3173 2022 3465 2036
rect 3173 1970 3180 2022
rect 3232 1970 3244 2022
rect 3296 1970 3465 2022
rect 3173 1957 3465 1970
rect 3173 1905 3180 1957
rect 3232 1905 3244 1957
rect 3296 1905 3465 1957
rect 3173 1892 3465 1905
rect 3173 1840 3180 1892
rect 3232 1840 3244 1892
rect 3296 1840 3465 1892
rect 3173 1827 3465 1840
rect 3173 1775 3180 1827
rect 3232 1775 3244 1827
rect 3296 1775 3465 1827
rect 3173 1762 3465 1775
rect 3173 1710 3180 1762
rect 3232 1710 3244 1762
rect 3296 1710 3465 1762
rect 3173 1697 3465 1710
rect 3173 1645 3180 1697
rect 3232 1645 3244 1697
rect 3296 1645 3465 1697
rect 3173 1632 3465 1645
rect 3173 1580 3180 1632
rect 3232 1580 3244 1632
rect 3296 1580 3465 1632
rect 3173 1567 3465 1580
rect 3173 1515 3180 1567
rect 3232 1515 3244 1567
rect 3296 1515 3465 1567
rect 3173 1502 3465 1515
rect 3173 1450 3180 1502
rect 3232 1450 3244 1502
rect 3296 1450 3465 1502
rect 3173 1437 3465 1450
rect 3173 1385 3180 1437
rect 3232 1385 3244 1437
rect 3296 1385 3465 1437
rect 3173 1372 3465 1385
rect 3173 1320 3180 1372
rect 3232 1320 3244 1372
rect 3296 1320 3465 1372
rect 3173 1307 3465 1320
rect 3173 1255 3180 1307
rect 3232 1255 3244 1307
rect 3296 1255 3465 1307
rect 3173 1242 3465 1255
rect 3173 1190 3180 1242
rect 3232 1190 3244 1242
rect 3296 1190 3465 1242
rect 3173 1177 3465 1190
rect 3173 1125 3180 1177
rect 3232 1125 3244 1177
rect 3296 1125 3465 1177
rect 3173 1112 3465 1125
rect 3173 1060 3180 1112
rect 3232 1060 3244 1112
rect 3296 1060 3465 1112
rect 3173 1047 3465 1060
rect 3173 995 3180 1047
rect 3232 995 3244 1047
rect 3296 995 3465 1047
rect 3173 982 3465 995
rect 3173 930 3180 982
rect 3232 930 3244 982
rect 3296 930 3465 982
rect 3173 917 3465 930
rect 3173 865 3180 917
rect 3232 865 3244 917
rect 3296 865 3465 917
rect 3173 852 3465 865
rect 3173 800 3180 852
rect 3232 800 3244 852
rect 3296 800 3465 852
rect 3173 787 3465 800
rect 3173 735 3180 787
rect 3232 735 3244 787
rect 3296 735 3465 787
rect 3173 722 3465 735
rect 3173 670 3180 722
rect 3232 670 3244 722
rect 3296 670 3465 722
rect 3173 657 3465 670
rect 3173 605 3180 657
rect 3232 605 3244 657
rect 3296 605 3465 657
rect 3173 592 3465 605
rect 3173 540 3180 592
rect 3232 540 3244 592
rect 3296 540 3465 592
rect 3173 527 3465 540
rect 3173 475 3180 527
rect 3232 475 3244 527
rect 3296 475 3465 527
rect 3173 462 3465 475
rect 3173 410 3180 462
rect 3232 410 3244 462
rect 3296 410 3465 462
rect 3173 397 3465 410
rect 3173 345 3180 397
rect 3232 345 3244 397
rect 3296 345 3465 397
rect 3173 332 3465 345
rect 3173 280 3180 332
rect 3232 280 3244 332
rect 3296 280 3465 332
rect 3173 267 3465 280
rect 3173 215 3180 267
rect 3232 215 3244 267
rect 3296 215 3465 267
tri 3164 202 3173 211 se
rect 3173 202 3465 215
tri 3157 195 3164 202 se
rect 3164 195 3180 202
tri 3145 183 3157 195 se
rect 3157 183 3180 195
tri 2040 158 2065 183 sw
tri 3120 158 3145 183 se
rect 3145 158 3180 183
rect 1977 150 3180 158
rect 3232 150 3244 202
rect 3296 150 3465 202
rect 1977 128 3465 150
rect 1977 80 2020 128
rect 1810 76 2020 80
rect 2072 76 2087 128
rect 2139 76 2154 128
rect 2206 76 2221 128
rect 2273 76 2288 128
rect 2340 76 2355 128
rect 2407 76 2422 128
rect 2474 76 2711 128
rect 2763 76 2778 128
rect 2830 76 2845 128
rect 2897 76 2912 128
rect 2964 76 2979 128
rect 3031 76 3046 128
rect 3098 76 3113 128
rect 3165 76 3465 128
rect 530 64 3465 76
rect 530 12 673 64
rect 725 12 740 64
rect 792 12 807 64
rect 859 12 874 64
rect 926 12 941 64
rect 993 12 1008 64
rect 1060 12 1075 64
rect 1127 12 1356 64
rect 1408 12 1423 64
rect 1475 12 1490 64
rect 1542 12 1557 64
rect 1609 12 1624 64
rect 1676 12 1691 64
rect 1743 12 1758 64
rect 1810 12 2020 64
rect 2072 12 2087 64
rect 2139 12 2154 64
rect 2206 12 2221 64
rect 2273 12 2288 64
rect 2340 12 2355 64
rect 2407 12 2422 64
rect 2474 12 2711 64
rect 2763 12 2778 64
rect 2830 12 2845 64
rect 2897 12 2912 64
rect 2964 12 2979 64
rect 3031 12 3046 64
rect 3098 12 3113 64
rect 3165 12 3465 64
rect 530 0 3465 12
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1701704242
transform 1 0 142 0 -1 2422
box 0 0 1 1
use L1M1_CDNS_52468879185945  L1M1_CDNS_52468879185945_0
timestamp 1701704242
transform 0 1 177 -1 0 2241
box -12 -6 1846 40
use nfet_CDNS_524688791851289  nfet_CDNS_524688791851289_0
timestamp 1701704242
transform 1 0 -14 0 1 346
box -79 -26 259 2026
use s8_esd_res250only_small  s8_esd_res250only_small_0
timestamp 1701704242
transform 0 -1 403 -1 0 5145
box 0 0 2270 404
use s8_esd_signal_5_sym_hv_local_5term  s8_esd_signal_5_sym_hv_local_5term_0
timestamp 1701704242
transform -1 0 3374 0 1 2550
box 0 0 1591 2424
use s8_esd_signal_5_sym_hv_local_5term  s8_esd_signal_5_sym_hv_local_5term_1
timestamp 1701704242
transform -1 0 3374 0 -1 2358
box 0 0 1591 2424
use s8_esd_signal_5_sym_hv_local_5term  s8_esd_signal_5_sym_hv_local_5term_2
timestamp 1701704242
transform 1 0 464 0 -1 2358
box 0 0 1591 2424
use s8_esd_signal_5_sym_hv_local_5term  s8_esd_signal_5_sym_hv_local_5term_3
timestamp 1701704242
transform 1 0 464 0 1 2550
box 0 0 1591 2424
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851288  sky130_fd_io__sio_tk_em1s_CDNS_524688791851288_0
timestamp 1701704242
transform -1 0 148 0 1 330
box 0 0 1 1
<< labels >>
flabel comment s 1638 380 1638 380 0 FreeSans 400 0 0 0 vnb
flabel comment s 1458 671 1458 671 0 FreeSans 400 0 0 0 vcc_ioq
flabel comment s 2130 4503 2130 4503 0 FreeSans 400 0 0 0 vnb
flabel comment s 1190 350 1190 350 0 FreeSans 400 0 0 0 vgnd
flabel comment s 2606 350 2606 350 0 FreeSans 400 0 0 0 vgnd
flabel comment s 2316 350 2316 350 0 FreeSans 400 0 0 0 vnb
flabel comment s 2982 350 2982 350 0 FreeSans 400 0 0 0 vnb
flabel comment s 807 380 807 380 0 FreeSans 400 0 0 0 vnb
flabel comment s 3260 52 3260 52 0 FreeSans 400 0 0 0 vcc_io
flabel comment s 548 52 548 52 0 FreeSans 400 0 0 0 vcc_io
flabel comment s 517 4109 517 4109 0 FreeSans 400 0 0 0 vcc_io
flabel comment s 1873 37 1873 37 0 FreeSans 400 0 0 0 vcc_io
flabel comment s 1888 4800 1888 4800 0 FreeSans 400 0 0 0 vcc_io
flabel comment s -26 4898 -26 4898 0 FreeSans 400 270 0 0 vpwr_ka
flabel metal1 s 1866 5047 1994 5162 3 FreeSans 400 0 0 0 pad
port 3 nsew
flabel metal1 s 3392 2468 3479 2588 0 FreeSans 200 0 0 0 pad_sw0
port 2 nsew
flabel metal2 s 2071 5408 2384 5504 0 FreeSans 400 0 0 0 vcc_ioq
port 4 nsew
flabel metal2 s 281 5004 333 5041 0 FreeSans 400 0 0 0 ng_ctl
port 5 nsew
flabel metal2 s 2586 5409 2768 5505 0 FreeSans 400 0 0 0 vgnd
port 6 nsew
flabel metal2 s 3173 5159 3465 5253 0 FreeSans 400 0 0 0 vcc_io
port 7 nsew
flabel metal2 s 715 4945 1035 5041 0 FreeSans 400 0 0 0 vgnd
port 6 nsew
<< properties >>
string GDS_END 86349172
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86240334
string path 62.000 1.750 50.350 1.750 
<< end >>
