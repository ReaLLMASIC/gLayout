magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< poly >>
rect -50 50 0 66
rect -50 16 -34 50
rect -50 0 0 16
rect 3736 50 3786 66
rect 3770 16 3786 50
rect 3736 0 3786 16
<< polycont >>
rect -34 16 0 50
rect 3736 16 3770 50
<< npolyres >>
rect 0 0 3736 66
<< locali >>
rect -34 50 0 66
rect -34 0 0 16
rect 3736 50 3770 66
rect 3736 0 3770 16
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_0
timestamp 1701704242
transform -1 0 16 0 1 0
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_1
timestamp 1701704242
transform 1 0 3720 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 80365180
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 80364746
<< end >>
