magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< dnwell >>
rect 7815 7803 12903 8364
rect 3717 6372 12903 7803
rect 3717 991 12253 6372
<< nwell >>
rect -625 13614 1361 14286
rect -625 13477 443 13614
rect -631 11917 443 13477
rect 11807 12009 12701 13485
rect 13109 11947 14756 14833
rect 7727 8117 13038 8459
rect 7727 7883 7926 8117
rect 3637 7472 7926 7883
rect 3637 6646 3997 7472
rect 4729 6646 4897 7472
rect 5589 6646 5757 7472
rect 6599 6646 6767 7472
rect 7602 6646 7770 7472
rect 12645 6646 13038 8117
rect 3637 6478 13038 6646
rect 3637 1023 3997 6478
rect 12046 6218 13038 6478
rect 12046 1023 12419 6218
rect 3637 681 12419 1023
<< pwell >>
rect 3053 14588 5147 14674
rect 3053 11922 3139 14588
rect 5061 11922 5147 14588
rect 5384 14281 9291 14367
rect 5384 12499 5470 14281
rect 8671 14048 8857 14281
rect 5718 13808 5904 13926
rect 9205 13772 9291 14281
rect 8981 13654 9291 13772
rect 9205 12692 9291 13654
rect 8973 12499 9291 12692
rect 5384 12413 9291 12499
rect 11660 13546 12851 13632
rect 3053 11836 5147 11922
rect 11660 11947 11746 13546
rect 12765 11947 12851 13546
rect 11660 11861 12851 11947
rect 8173 7971 12407 8057
rect 4082 7326 4648 7412
rect 4082 6917 4168 7326
rect 4562 6917 4648 7326
rect 4082 6831 4648 6917
rect 4962 7326 5528 7412
rect 4962 6917 5048 7326
rect 5442 6917 5528 7326
rect 4962 6831 5528 6917
rect 5824 7326 6390 7412
rect 5824 6917 5910 7326
rect 6304 6917 6390 7326
rect 5824 6831 6390 6917
rect 6954 7326 7520 7412
rect 6954 6917 7040 7326
rect 7434 6917 7520 7326
rect 6954 6831 7520 6917
rect 8173 6706 12407 6792
rect 11897 1917 11985 5738
<< ndiff >>
rect 8697 14124 8831 14140
rect 8697 14090 8709 14124
rect 8743 14090 8785 14124
rect 8819 14090 8831 14124
rect 8697 14074 8831 14090
rect 5744 13884 5878 13900
rect 5744 13850 5756 13884
rect 5790 13850 5832 13884
rect 5866 13850 5878 13884
rect 5744 13834 5878 13850
rect 9007 13730 9141 13746
rect 9007 13696 9019 13730
rect 9053 13696 9095 13730
rect 9129 13696 9141 13730
rect 9007 13680 9141 13696
rect 8999 12650 9133 12666
rect 8999 12616 9011 12650
rect 9045 12616 9087 12650
rect 9121 12616 9133 12650
rect 8999 12600 9133 12616
<< ndiffc >>
rect 8709 14090 8743 14124
rect 8785 14090 8819 14124
rect 5756 13850 5790 13884
rect 5832 13850 5866 13884
rect 9019 13696 9053 13730
rect 9095 13696 9129 13730
rect 9011 12616 9045 12650
rect 9087 12616 9121 12650
<< psubdiff >>
rect 3079 14614 3147 14648
rect 3181 14614 3215 14648
rect 3249 14614 3283 14648
rect 3317 14614 3351 14648
rect 3385 14614 3419 14648
rect 3453 14614 3487 14648
rect 3521 14614 3555 14648
rect 3589 14614 3623 14648
rect 3657 14614 3691 14648
rect 3725 14614 3759 14648
rect 3793 14614 3827 14648
rect 3861 14614 3895 14648
rect 3929 14614 3963 14648
rect 3997 14614 4031 14648
rect 4065 14614 4099 14648
rect 4133 14614 4167 14648
rect 4201 14614 4235 14648
rect 4269 14614 4303 14648
rect 4337 14614 4371 14648
rect 4405 14614 4439 14648
rect 4473 14614 4507 14648
rect 4541 14614 4575 14648
rect 4609 14614 4643 14648
rect 4677 14614 4711 14648
rect 4745 14614 4779 14648
rect 4813 14614 4847 14648
rect 4881 14614 4915 14648
rect 4949 14614 4983 14648
rect 5017 14614 5121 14648
rect 3079 14558 3113 14614
rect 5087 14580 5121 14614
rect 3079 14490 3113 14524
rect 5087 14512 5121 14546
rect 3079 14422 3113 14456
rect 3079 14354 3113 14388
rect 3079 14286 3113 14320
rect 3079 14218 3113 14252
rect 3079 14150 3113 14184
rect 3079 14082 3113 14116
rect 3079 14014 3113 14048
rect 3079 13946 3113 13980
rect 3079 13878 3113 13912
rect 3079 13810 3113 13844
rect 3079 13742 3113 13776
rect 3079 13674 3113 13708
rect 3079 13606 3113 13640
rect 3079 13538 3113 13572
rect 3079 13470 3113 13504
rect 3079 13402 3113 13436
rect 3079 13334 3113 13368
rect 3079 13266 3113 13300
rect 3079 13198 3113 13232
rect 3079 13130 3113 13164
rect 3079 13062 3113 13096
rect 3079 12994 3113 13028
rect 5087 14444 5121 14478
rect 5087 14376 5121 14410
rect 5087 14308 5121 14342
rect 5087 14240 5121 14274
rect 5087 14172 5121 14206
rect 5087 14104 5121 14138
rect 5087 14036 5121 14070
rect 5087 13968 5121 14002
rect 5087 13900 5121 13934
rect 5087 13832 5121 13866
rect 5087 13764 5121 13798
rect 5087 13696 5121 13730
rect 5087 13628 5121 13662
rect 5087 13560 5121 13594
rect 5087 13492 5121 13526
rect 5087 13424 5121 13458
rect 5087 13356 5121 13390
rect 5087 13288 5121 13322
rect 5087 13220 5121 13254
rect 5087 13152 5121 13186
rect 5087 13084 5121 13118
rect 5087 13016 5121 13050
rect 3079 12926 3113 12960
rect 5087 12948 5121 12982
rect 3079 12858 3113 12892
rect 3079 12790 3113 12824
rect 3079 12722 3113 12756
rect 3079 12576 3113 12688
rect 3079 12508 3113 12542
rect 3079 12440 3113 12474
rect 5087 12880 5121 12914
rect 5087 12812 5121 12846
rect 5087 12744 5121 12778
rect 5087 12676 5121 12710
rect 5087 12608 5121 12642
rect 5087 12540 5121 12574
rect 5087 12472 5121 12506
rect 5410 14307 5478 14341
rect 5512 14307 5546 14341
rect 5580 14307 5614 14341
rect 5648 14307 5682 14341
rect 5716 14307 5750 14341
rect 5784 14307 5818 14341
rect 5852 14307 5886 14341
rect 5920 14307 5954 14341
rect 5988 14307 6022 14341
rect 6056 14307 6090 14341
rect 6124 14307 6158 14341
rect 6192 14307 6226 14341
rect 6260 14307 6294 14341
rect 6328 14307 6362 14341
rect 6396 14307 6430 14341
rect 6464 14307 6498 14341
rect 6532 14307 6566 14341
rect 6600 14307 6634 14341
rect 6668 14307 6702 14341
rect 6736 14307 6770 14341
rect 6804 14307 6838 14341
rect 6872 14307 6906 14341
rect 6940 14307 6974 14341
rect 7008 14307 7042 14341
rect 7076 14307 7110 14341
rect 7144 14307 7178 14341
rect 7212 14307 7246 14341
rect 7280 14307 7314 14341
rect 7348 14307 7382 14341
rect 7416 14307 7450 14341
rect 7484 14307 7518 14341
rect 7552 14307 7586 14341
rect 7620 14307 7654 14341
rect 7688 14307 7722 14341
rect 7756 14307 7790 14341
rect 7824 14307 7858 14341
rect 7892 14307 7926 14341
rect 7960 14307 7994 14341
rect 8028 14307 8062 14341
rect 8096 14307 8130 14341
rect 8164 14307 8198 14341
rect 8232 14307 8266 14341
rect 8300 14307 8334 14341
rect 8368 14307 8402 14341
rect 8436 14307 8470 14341
rect 8504 14307 8538 14341
rect 8572 14307 8606 14341
rect 8640 14307 8674 14341
rect 8708 14307 8742 14341
rect 8776 14307 8810 14341
rect 8844 14307 8878 14341
rect 8912 14307 8946 14341
rect 8980 14307 9014 14341
rect 9048 14307 9082 14341
rect 9116 14307 9150 14341
rect 9184 14307 9265 14341
rect 5410 14241 5444 14307
rect 5410 14173 5444 14207
rect 9231 14273 9265 14307
rect 9231 14205 9265 14239
rect 5410 14105 5444 14139
rect 9231 14137 9265 14171
rect 5410 14037 5444 14071
rect 5410 13969 5444 14003
rect 5410 13901 5444 13935
rect 9231 14069 9265 14103
rect 9231 14001 9265 14035
rect 9231 13933 9265 13967
rect 5410 13833 5444 13867
rect 9231 13865 9265 13899
rect 5410 13765 5444 13799
rect 9231 13797 9265 13831
rect 5410 13697 5444 13731
rect 9231 13729 9265 13763
rect 5410 13629 5444 13663
rect 5410 13561 5444 13595
rect 5410 13493 5444 13527
rect 5410 13425 5444 13459
rect 5410 13357 5444 13391
rect 5410 13289 5444 13323
rect 5410 13221 5444 13255
rect 5410 13153 5444 13187
rect 5410 13085 5444 13119
rect 5410 13017 5444 13051
rect 5410 12949 5444 12983
rect 5410 12881 5444 12915
rect 5410 12813 5444 12847
rect 5410 12745 5444 12779
rect 5410 12677 5444 12711
rect 9231 13661 9265 13695
rect 9231 13593 9265 13627
rect 9231 13525 9265 13559
rect 9231 13457 9265 13491
rect 9231 13389 9265 13423
rect 9231 13321 9265 13355
rect 9231 13253 9265 13287
rect 9231 13185 9265 13219
rect 9231 13117 9265 13151
rect 9231 13049 9265 13083
rect 9231 12981 9265 13015
rect 9231 12913 9265 12947
rect 9231 12845 9265 12879
rect 9231 12777 9265 12811
rect 9231 12709 9265 12743
rect 5410 12609 5444 12643
rect 9231 12641 9265 12675
rect 5410 12541 5444 12575
rect 5410 12473 5444 12507
rect 9231 12573 9265 12607
rect 9231 12473 9265 12539
rect 5410 12439 5524 12473
rect 5558 12439 5592 12473
rect 5626 12439 5660 12473
rect 5694 12439 5728 12473
rect 5762 12439 5796 12473
rect 5830 12439 5864 12473
rect 5898 12439 5932 12473
rect 5966 12439 6000 12473
rect 6034 12439 6068 12473
rect 6102 12439 6136 12473
rect 6170 12439 6204 12473
rect 6238 12439 6272 12473
rect 6306 12439 6340 12473
rect 6374 12439 6408 12473
rect 6442 12439 6476 12473
rect 6510 12439 6544 12473
rect 6578 12439 6612 12473
rect 6646 12439 6680 12473
rect 6714 12439 6748 12473
rect 6782 12439 6816 12473
rect 6850 12439 6884 12473
rect 6918 12439 6952 12473
rect 6986 12439 7020 12473
rect 7054 12439 7088 12473
rect 7122 12439 7156 12473
rect 7190 12439 7224 12473
rect 7258 12439 7292 12473
rect 7326 12439 7360 12473
rect 7394 12439 7428 12473
rect 7462 12439 7496 12473
rect 7530 12439 7564 12473
rect 7598 12439 7632 12473
rect 7666 12439 7700 12473
rect 7734 12439 7768 12473
rect 7802 12439 7836 12473
rect 7870 12439 7939 12473
rect 7973 12439 8007 12473
rect 8041 12439 8075 12473
rect 8109 12439 8143 12473
rect 8177 12439 8211 12473
rect 8245 12439 8279 12473
rect 8313 12439 8347 12473
rect 8381 12439 8415 12473
rect 8449 12439 8483 12473
rect 8517 12439 8551 12473
rect 8585 12439 8619 12473
rect 8653 12439 8687 12473
rect 8721 12439 8755 12473
rect 8789 12439 8823 12473
rect 8857 12439 8891 12473
rect 8925 12439 8959 12473
rect 8993 12439 9027 12473
rect 9061 12439 9095 12473
rect 9129 12439 9163 12473
rect 9197 12439 9265 12473
rect 11686 13572 11771 13606
rect 11805 13572 11839 13606
rect 11873 13572 11907 13606
rect 11941 13572 11975 13606
rect 12009 13572 12043 13606
rect 12077 13572 12111 13606
rect 12145 13572 12179 13606
rect 12213 13572 12247 13606
rect 12281 13572 12315 13606
rect 12349 13572 12383 13606
rect 12417 13572 12451 13606
rect 12485 13572 12519 13606
rect 12553 13572 12587 13606
rect 12621 13572 12655 13606
rect 12689 13572 12723 13606
rect 12757 13572 12825 13606
rect 11686 13538 11720 13572
rect 11686 13470 11720 13504
rect 11686 13402 11720 13436
rect 12791 13485 12825 13572
rect 11686 13334 11720 13368
rect 11686 13266 11720 13300
rect 11686 13198 11720 13232
rect 11686 13130 11720 13164
rect 11686 13062 11720 13096
rect 11686 12994 11720 13028
rect 11686 12926 11720 12960
rect 11686 12858 11720 12892
rect 11686 12790 11720 12824
rect 11686 12722 11720 12756
rect 11686 12654 11720 12688
rect 11686 12586 11720 12620
rect 11686 12518 11720 12552
rect 11686 12450 11720 12484
rect 3079 12372 3113 12406
rect 3079 12304 3113 12338
rect 5087 12404 5121 12438
rect 5087 12336 5121 12370
rect 3079 12236 3113 12270
rect 3079 12168 3113 12202
rect 3079 12100 3113 12134
rect 3079 12032 3113 12066
rect 5087 12268 5121 12302
rect 5087 12200 5121 12234
rect 5087 12132 5121 12166
rect 5087 12064 5121 12098
rect 3079 11964 3113 11998
rect 5087 11996 5121 12030
rect 3079 11896 3113 11930
rect 5087 11896 5121 11962
rect 3079 11862 3183 11896
rect 3217 11862 3251 11896
rect 3285 11862 3319 11896
rect 3353 11862 3387 11896
rect 3421 11862 3455 11896
rect 3489 11862 3523 11896
rect 3557 11862 3591 11896
rect 3625 11862 3659 11896
rect 3693 11862 3727 11896
rect 3761 11862 3795 11896
rect 3829 11862 3863 11896
rect 3897 11862 3931 11896
rect 3965 11862 3999 11896
rect 4033 11862 4067 11896
rect 4101 11862 4135 11896
rect 4169 11862 4203 11896
rect 4237 11862 4271 11896
rect 4305 11862 4339 11896
rect 4373 11862 4407 11896
rect 4441 11862 4475 11896
rect 4509 11862 4543 11896
rect 4577 11862 4611 11896
rect 4645 11862 4679 11896
rect 4713 11862 4747 11896
rect 4781 11862 4815 11896
rect 4849 11862 4883 11896
rect 4917 11862 4951 11896
rect 4985 11862 5019 11896
rect 5053 11862 5121 11896
rect 11686 12382 11720 12416
rect 11686 12314 11720 12348
rect 11686 12246 11720 12280
rect 11686 12178 11720 12212
rect 11686 12110 11720 12144
rect 12791 13417 12825 13451
rect 12791 13349 12825 13383
rect 12791 13281 12825 13315
rect 12791 13213 12825 13247
rect 12791 13145 12825 13179
rect 12791 13077 12825 13111
rect 12791 13009 12825 13043
rect 12791 12941 12825 12975
rect 12791 12873 12825 12907
rect 12791 12805 12825 12839
rect 12791 12737 12825 12771
rect 12791 12669 12825 12703
rect 12791 12601 12825 12635
rect 12791 12533 12825 12567
rect 12791 12465 12825 12499
rect 12791 12397 12825 12431
rect 12791 12329 12825 12363
rect 12791 12261 12825 12295
rect 12791 12193 12825 12227
rect 12791 12125 12825 12159
rect 11686 12042 11720 12076
rect 11686 11921 11720 12008
rect 12791 12057 12825 12091
rect 12791 11989 12825 12023
rect 12791 11921 12825 11955
rect 11686 11887 11754 11921
rect 11788 11887 11822 11921
rect 11856 11887 11890 11921
rect 11924 11887 11958 11921
rect 11992 11887 12026 11921
rect 12060 11887 12094 11921
rect 12128 11887 12162 11921
rect 12196 11887 12230 11921
rect 12264 11887 12298 11921
rect 12332 11887 12366 11921
rect 12400 11887 12434 11921
rect 12468 11887 12502 11921
rect 12536 11887 12570 11921
rect 12604 11887 12638 11921
rect 12672 11887 12706 11921
rect 12740 11887 12825 11921
rect 8199 7997 8233 8031
rect 8267 7997 8301 8031
rect 8335 7997 8369 8031
rect 8403 7997 8437 8031
rect 8471 7997 8505 8031
rect 8539 7997 8573 8031
rect 8607 7997 8641 8031
rect 8675 7997 8709 8031
rect 8743 7997 8777 8031
rect 8811 7997 8845 8031
rect 8879 7997 8913 8031
rect 8947 7997 8981 8031
rect 9015 7997 9049 8031
rect 9083 7997 9117 8031
rect 9151 7997 9185 8031
rect 9219 7997 9253 8031
rect 9287 7997 9321 8031
rect 9355 7997 9389 8031
rect 9423 7997 9457 8031
rect 9491 7997 9525 8031
rect 9559 7997 9593 8031
rect 9627 7997 9661 8031
rect 9695 7997 9729 8031
rect 9763 7997 9797 8031
rect 9831 7997 9865 8031
rect 9899 7997 9933 8031
rect 9967 7997 10001 8031
rect 10035 7997 10069 8031
rect 10103 7997 10137 8031
rect 10171 7997 10205 8031
rect 10239 7997 10273 8031
rect 10307 7997 10341 8031
rect 10375 7997 10409 8031
rect 10443 7997 10477 8031
rect 10511 7997 10545 8031
rect 10579 7997 10613 8031
rect 10647 7997 10681 8031
rect 10715 7997 10749 8031
rect 10783 7997 10817 8031
rect 10851 7997 10885 8031
rect 10919 7997 10953 8031
rect 10987 7997 11021 8031
rect 11055 7997 11089 8031
rect 11123 7997 11157 8031
rect 11191 7997 11225 8031
rect 11259 7997 11293 8031
rect 11327 7997 11361 8031
rect 11395 7997 11429 8031
rect 11463 7997 11497 8031
rect 11531 7997 11565 8031
rect 11599 7997 11633 8031
rect 11667 7997 11701 8031
rect 11735 7997 11769 8031
rect 11803 7997 11837 8031
rect 11871 7997 11905 8031
rect 11939 7997 11973 8031
rect 12007 7997 12041 8031
rect 12075 7997 12109 8031
rect 12143 7997 12177 8031
rect 12211 7997 12245 8031
rect 12279 7997 12313 8031
rect 12347 7997 12381 8031
rect 4108 7352 4180 7386
rect 4214 7352 4248 7386
rect 4282 7352 4316 7386
rect 4350 7352 4384 7386
rect 4418 7352 4452 7386
rect 4486 7352 4520 7386
rect 4554 7352 4622 7386
rect 4108 7318 4142 7352
rect 4108 7250 4142 7284
rect 4588 7299 4622 7352
rect 4588 7231 4622 7265
rect 4108 7182 4142 7216
rect 4108 7114 4142 7148
rect 4108 7046 4142 7080
rect 4588 7163 4622 7197
rect 4588 7095 4622 7129
rect 4108 6978 4142 7012
rect 4108 6891 4142 6944
rect 4588 7027 4622 7061
rect 4588 6959 4622 6993
rect 4588 6891 4622 6925
rect 4108 6857 4176 6891
rect 4210 6857 4244 6891
rect 4278 6857 4312 6891
rect 4346 6857 4380 6891
rect 4414 6857 4448 6891
rect 4482 6857 4622 6891
rect 4988 7352 5060 7386
rect 5094 7352 5128 7386
rect 5162 7352 5196 7386
rect 5230 7352 5264 7386
rect 5298 7352 5332 7386
rect 5366 7352 5400 7386
rect 5434 7352 5502 7386
rect 4988 7318 5022 7352
rect 4988 7250 5022 7284
rect 5468 7299 5502 7352
rect 5468 7231 5502 7265
rect 4988 7182 5022 7216
rect 4988 7114 5022 7148
rect 4988 7046 5022 7080
rect 5468 7163 5502 7197
rect 5468 7095 5502 7129
rect 4988 6978 5022 7012
rect 4988 6891 5022 6944
rect 5468 7027 5502 7061
rect 5468 6959 5502 6993
rect 5468 6891 5502 6925
rect 4988 6857 5056 6891
rect 5090 6857 5124 6891
rect 5158 6857 5192 6891
rect 5226 6857 5260 6891
rect 5294 6857 5328 6891
rect 5362 6857 5502 6891
rect 5850 7352 5922 7386
rect 5956 7352 5990 7386
rect 6024 7352 6058 7386
rect 6092 7352 6126 7386
rect 6160 7352 6194 7386
rect 6228 7352 6262 7386
rect 6296 7352 6364 7386
rect 5850 7318 5884 7352
rect 5850 7250 5884 7284
rect 6330 7299 6364 7352
rect 6330 7231 6364 7265
rect 5850 7182 5884 7216
rect 5850 7114 5884 7148
rect 5850 7046 5884 7080
rect 6330 7163 6364 7197
rect 6330 7095 6364 7129
rect 5850 6978 5884 7012
rect 5850 6891 5884 6944
rect 6330 7027 6364 7061
rect 6330 6959 6364 6993
rect 6330 6891 6364 6925
rect 5850 6857 5918 6891
rect 5952 6857 5986 6891
rect 6020 6857 6054 6891
rect 6088 6857 6122 6891
rect 6156 6857 6190 6891
rect 6224 6857 6364 6891
rect 6980 7352 7052 7386
rect 7086 7352 7120 7386
rect 7154 7352 7188 7386
rect 7222 7352 7256 7386
rect 7290 7352 7324 7386
rect 7358 7352 7392 7386
rect 7426 7352 7494 7386
rect 6980 7318 7014 7352
rect 6980 7250 7014 7284
rect 7460 7299 7494 7352
rect 7460 7231 7494 7265
rect 6980 7182 7014 7216
rect 6980 7114 7014 7148
rect 6980 7046 7014 7080
rect 7460 7163 7494 7197
rect 7460 7095 7494 7129
rect 6980 6978 7014 7012
rect 6980 6891 7014 6944
rect 7460 7027 7494 7061
rect 7460 6959 7494 6993
rect 7460 6891 7494 6925
rect 6980 6857 7048 6891
rect 7082 6857 7116 6891
rect 7150 6857 7184 6891
rect 7218 6857 7252 6891
rect 7286 6857 7320 6891
rect 7354 6857 7494 6891
rect 8199 6732 8233 6766
rect 8267 6732 8301 6766
rect 8335 6732 8369 6766
rect 8403 6732 8437 6766
rect 8471 6732 8505 6766
rect 8539 6732 8573 6766
rect 8607 6732 8641 6766
rect 8675 6732 8709 6766
rect 8743 6732 8777 6766
rect 8811 6732 8845 6766
rect 8879 6732 8913 6766
rect 8947 6732 8981 6766
rect 9015 6732 9049 6766
rect 9083 6732 9117 6766
rect 9151 6732 9185 6766
rect 9219 6732 9253 6766
rect 9287 6732 9321 6766
rect 9355 6732 9389 6766
rect 9423 6732 9457 6766
rect 9491 6732 9525 6766
rect 9559 6732 9593 6766
rect 9627 6732 9661 6766
rect 9695 6732 9729 6766
rect 9763 6732 9797 6766
rect 9831 6732 9865 6766
rect 9899 6732 9933 6766
rect 9967 6732 10001 6766
rect 10035 6732 10069 6766
rect 10103 6732 10137 6766
rect 10171 6732 10205 6766
rect 10239 6732 10273 6766
rect 10307 6732 10341 6766
rect 10375 6732 10409 6766
rect 10443 6732 10477 6766
rect 10511 6732 10545 6766
rect 10579 6732 10613 6766
rect 10647 6732 10681 6766
rect 10715 6732 10749 6766
rect 10783 6732 10817 6766
rect 10851 6732 10885 6766
rect 10919 6732 10953 6766
rect 10987 6732 11021 6766
rect 11055 6732 11089 6766
rect 11123 6732 11157 6766
rect 11191 6732 11225 6766
rect 11259 6732 11293 6766
rect 11327 6732 11361 6766
rect 11395 6732 11429 6766
rect 11463 6732 11497 6766
rect 11531 6732 11565 6766
rect 11599 6732 11633 6766
rect 11667 6732 11701 6766
rect 11735 6732 11769 6766
rect 11803 6732 11837 6766
rect 11871 6732 11905 6766
rect 11939 6732 11973 6766
rect 12007 6732 12041 6766
rect 12075 6732 12109 6766
rect 12143 6732 12177 6766
rect 12211 6732 12245 6766
rect 12279 6732 12313 6766
rect 12347 6732 12381 6766
rect 11923 5678 11959 5712
rect 11923 5644 11924 5678
rect 11958 5644 11959 5678
rect 11923 5610 11959 5644
rect 11923 5576 11924 5610
rect 11958 5576 11959 5610
rect 11923 5542 11959 5576
rect 11923 5508 11924 5542
rect 11958 5508 11959 5542
rect 11923 5474 11959 5508
rect 11923 5440 11924 5474
rect 11958 5440 11959 5474
rect 11923 5406 11959 5440
rect 11923 5372 11924 5406
rect 11958 5372 11959 5406
rect 11923 5338 11959 5372
rect 11923 5304 11924 5338
rect 11958 5304 11959 5338
rect 11923 5270 11959 5304
rect 11923 5236 11924 5270
rect 11958 5236 11959 5270
rect 11923 5202 11959 5236
rect 11923 5168 11924 5202
rect 11958 5168 11959 5202
rect 11923 5134 11959 5168
rect 11923 5100 11924 5134
rect 11958 5100 11959 5134
rect 11923 5066 11959 5100
rect 11923 5032 11924 5066
rect 11958 5032 11959 5066
rect 11923 4998 11959 5032
rect 11923 4964 11924 4998
rect 11958 4964 11959 4998
rect 11923 4930 11959 4964
rect 11923 4896 11924 4930
rect 11958 4896 11959 4930
rect 11923 4862 11959 4896
rect 11923 4828 11924 4862
rect 11958 4828 11959 4862
rect 11923 4794 11959 4828
rect 11923 4760 11924 4794
rect 11958 4760 11959 4794
rect 11923 4726 11959 4760
rect 11923 4692 11924 4726
rect 11958 4692 11959 4726
rect 11923 4658 11959 4692
rect 11923 4624 11924 4658
rect 11958 4624 11959 4658
rect 11923 4590 11959 4624
rect 11923 4556 11924 4590
rect 11958 4556 11959 4590
rect 11923 4522 11959 4556
rect 11923 4488 11924 4522
rect 11958 4488 11959 4522
rect 11923 4454 11959 4488
rect 11923 4420 11924 4454
rect 11958 4420 11959 4454
rect 11923 4386 11959 4420
rect 11923 4352 11924 4386
rect 11958 4352 11959 4386
rect 11923 4318 11959 4352
rect 11923 4284 11924 4318
rect 11958 4284 11959 4318
rect 11923 4250 11959 4284
rect 11923 4216 11924 4250
rect 11958 4216 11959 4250
rect 11923 4182 11959 4216
rect 11923 4148 11924 4182
rect 11958 4148 11959 4182
rect 11923 4114 11959 4148
rect 11923 4080 11924 4114
rect 11958 4080 11959 4114
rect 11923 4046 11959 4080
rect 11923 4012 11924 4046
rect 11958 4012 11959 4046
rect 11923 3978 11959 4012
rect 11923 3944 11924 3978
rect 11958 3944 11959 3978
rect 11923 3910 11959 3944
rect 11923 3876 11924 3910
rect 11958 3876 11959 3910
rect 11923 3842 11959 3876
rect 11923 3808 11924 3842
rect 11958 3808 11959 3842
rect 11923 3774 11959 3808
rect 11923 3740 11924 3774
rect 11958 3740 11959 3774
rect 11923 3706 11959 3740
rect 11923 3672 11924 3706
rect 11958 3672 11959 3706
rect 11923 3638 11959 3672
rect 11923 3604 11924 3638
rect 11958 3604 11959 3638
rect 11923 3570 11959 3604
rect 11923 3536 11924 3570
rect 11958 3536 11959 3570
rect 11923 3502 11959 3536
rect 11923 3468 11924 3502
rect 11958 3468 11959 3502
rect 11923 3434 11959 3468
rect 11923 3400 11924 3434
rect 11958 3400 11959 3434
rect 11923 3366 11959 3400
rect 11923 3332 11924 3366
rect 11958 3332 11959 3366
rect 11923 3298 11959 3332
rect 11923 3264 11924 3298
rect 11958 3264 11959 3298
rect 11923 3230 11959 3264
rect 11923 3196 11924 3230
rect 11958 3196 11959 3230
rect 11923 3162 11959 3196
rect 11923 3128 11924 3162
rect 11958 3128 11959 3162
rect 11923 3094 11959 3128
rect 11923 3060 11924 3094
rect 11958 3060 11959 3094
rect 11923 3026 11959 3060
rect 11923 2992 11924 3026
rect 11958 2992 11959 3026
rect 11923 2958 11959 2992
rect 11923 2924 11924 2958
rect 11958 2924 11959 2958
rect 11923 2890 11959 2924
rect 11923 2856 11924 2890
rect 11958 2856 11959 2890
rect 11923 2822 11959 2856
rect 11923 2788 11924 2822
rect 11958 2788 11959 2822
rect 11923 2754 11959 2788
rect 11923 2720 11924 2754
rect 11958 2720 11959 2754
rect 11923 2686 11959 2720
rect 11923 2652 11924 2686
rect 11958 2652 11959 2686
rect 11923 2618 11959 2652
rect 11923 2584 11924 2618
rect 11958 2584 11959 2618
rect 11923 2550 11959 2584
rect 11923 2516 11924 2550
rect 11958 2516 11959 2550
rect 11923 2482 11959 2516
rect 11923 2448 11924 2482
rect 11958 2448 11959 2482
rect 11923 2414 11959 2448
rect 11923 2380 11924 2414
rect 11958 2380 11959 2414
rect 11923 2346 11959 2380
rect 11923 2312 11924 2346
rect 11958 2312 11959 2346
rect 11923 2278 11959 2312
rect 11923 2244 11924 2278
rect 11958 2244 11959 2278
rect 11923 2210 11959 2244
rect 11923 2176 11924 2210
rect 11958 2176 11959 2210
rect 11923 2142 11959 2176
rect 11923 2108 11924 2142
rect 11958 2108 11959 2142
rect 11923 2074 11959 2108
rect 11923 2040 11924 2074
rect 11958 2040 11959 2074
rect 11923 1943 11959 2040
<< nsubdiff >>
rect 13176 14732 13244 14766
rect 13278 14732 13312 14766
rect 13346 14732 13380 14766
rect 13414 14732 13448 14766
rect 13482 14732 13516 14766
rect 13550 14732 13584 14766
rect 13618 14732 13652 14766
rect 13686 14732 13720 14766
rect 13754 14732 13788 14766
rect 13822 14732 13856 14766
rect 13890 14732 13924 14766
rect 13958 14732 13992 14766
rect 14026 14732 14060 14766
rect 14094 14732 14128 14766
rect 14162 14732 14196 14766
rect 14230 14732 14264 14766
rect 14298 14732 14332 14766
rect 14366 14732 14400 14766
rect 14434 14732 14468 14766
rect 14502 14732 14536 14766
rect 14570 14732 14689 14766
rect -564 13376 -496 13410
rect -462 13376 -428 13410
rect -394 13376 -360 13410
rect -326 13376 -292 13410
rect -258 13376 -224 13410
rect -190 13376 -156 13410
rect -122 13376 -88 13410
rect -54 13376 -20 13410
rect 14 13376 48 13410
rect 82 13376 116 13410
rect 150 13376 184 13410
rect 218 13376 252 13410
rect 286 13376 320 13410
rect 354 13376 407 13410
rect -564 13298 -530 13376
rect -564 13230 -530 13264
rect -564 13162 -530 13196
rect -564 13094 -530 13128
rect -564 13026 -530 13060
rect -564 12958 -530 12992
rect -564 12890 -530 12924
rect -564 12822 -530 12856
rect -564 12754 -530 12788
rect -564 12686 -530 12720
rect -564 12618 -530 12652
rect -564 12550 -530 12584
rect -564 12482 -530 12516
rect -564 12414 -530 12448
rect -564 12346 -530 12380
rect -564 12278 -530 12312
rect -564 12210 -530 12244
rect -564 12142 -530 12176
rect 13176 14632 13210 14732
rect 14655 14698 14689 14732
rect 14655 14630 14689 14664
rect 13176 14564 13210 14598
rect 13176 14496 13210 14530
rect 14655 14562 14689 14596
rect 13176 14428 13210 14462
rect 13176 14360 13210 14394
rect 13176 14292 13210 14326
rect 13176 14224 13210 14258
rect 13176 14156 13210 14190
rect 13176 14088 13210 14122
rect 13176 14020 13210 14054
rect 13176 13952 13210 13986
rect 13176 13884 13210 13918
rect 13176 13816 13210 13850
rect 13176 13748 13210 13782
rect 13176 13680 13210 13714
rect 13176 13612 13210 13646
rect -564 12074 -530 12108
rect -564 12006 -530 12040
rect 11874 13384 11988 13418
rect 12022 13384 12056 13418
rect 12090 13384 12124 13418
rect 12158 13384 12192 13418
rect 12226 13384 12260 13418
rect 12294 13384 12328 13418
rect 12362 13384 12396 13418
rect 12430 13384 12464 13418
rect 12498 13384 12532 13418
rect 12566 13384 12634 13418
rect 11874 13350 11908 13384
rect 11874 13282 11908 13316
rect 11874 13214 11908 13248
rect 11874 13146 11908 13180
rect 11874 13078 11908 13112
rect 11874 13010 11908 13044
rect 11874 12942 11908 12976
rect 11874 12874 11908 12908
rect 11874 12806 11908 12840
rect 11874 12738 11908 12772
rect 11874 12670 11908 12704
rect 11874 12602 11908 12636
rect 11874 12534 11908 12568
rect 11874 12466 11908 12500
rect 11874 12398 11908 12432
rect 11874 12330 11908 12364
rect 11874 12262 11908 12296
rect 11874 12110 11908 12228
rect 12600 13334 12634 13384
rect 12600 13266 12634 13300
rect 12600 13198 12634 13232
rect 12600 13130 12634 13164
rect 12600 13062 12634 13096
rect 12600 12994 12634 13028
rect 12600 12926 12634 12960
rect 12600 12858 12634 12892
rect 12600 12790 12634 12824
rect 12600 12722 12634 12756
rect 12600 12654 12634 12688
rect 12600 12586 12634 12620
rect 12600 12518 12634 12552
rect 12600 12450 12634 12484
rect 12600 12382 12634 12416
rect 12600 12314 12634 12348
rect 12600 12246 12634 12280
rect 12600 12178 12634 12212
rect 12600 12110 12634 12144
rect 11874 12076 11942 12110
rect 11976 12076 12010 12110
rect 12044 12076 12078 12110
rect 12112 12076 12146 12110
rect 12180 12076 12214 12110
rect 12248 12076 12282 12110
rect 12316 12076 12350 12110
rect 12384 12076 12418 12110
rect 12452 12076 12486 12110
rect 12520 12076 12634 12110
rect 13176 13544 13210 13578
rect 13176 13476 13210 13510
rect 14655 14494 14689 14528
rect 14655 14426 14689 14460
rect 14655 14358 14689 14392
rect 14655 14290 14689 14324
rect 14655 14222 14689 14256
rect 14655 14154 14689 14188
rect 14655 14086 14689 14120
rect 14655 14018 14689 14052
rect 14655 13950 14689 13984
rect 14655 13882 14689 13916
rect 14655 13814 14689 13848
rect 14655 13746 14689 13780
rect 14655 13678 14689 13712
rect 14655 13610 14689 13644
rect 14655 13542 14689 13576
rect 14655 13474 14689 13508
rect 13176 13408 13210 13442
rect 13176 13340 13210 13374
rect 13176 13272 13210 13306
rect 14655 13406 14689 13440
rect 14655 13338 14689 13372
rect 14655 13270 14689 13304
rect 13176 13204 13210 13238
rect 13176 13136 13210 13170
rect 13176 13068 13210 13102
rect 13176 13000 13210 13034
rect 13176 12932 13210 12966
rect 13176 12864 13210 12898
rect 13176 12796 13210 12830
rect 13176 12728 13210 12762
rect 13176 12660 13210 12694
rect 13176 12592 13210 12626
rect 13176 12524 13210 12558
rect 13176 12456 13210 12490
rect 13176 12388 13210 12422
rect 13176 12320 13210 12354
rect 13176 12252 13210 12286
rect 13176 12184 13210 12218
rect 14655 13202 14689 13236
rect 14655 13134 14689 13168
rect 14655 13066 14689 13100
rect 14655 12998 14689 13032
rect 14655 12930 14689 12964
rect 14655 12862 14689 12896
rect 14655 12794 14689 12828
rect 14655 12726 14689 12760
rect 14655 12658 14689 12692
rect 14655 12590 14689 12624
rect 14655 12522 14689 12556
rect 14655 12454 14689 12488
rect 14655 12386 14689 12420
rect 14655 12318 14689 12352
rect 14655 12250 14689 12284
rect 13176 12116 13210 12150
rect 14655 12182 14689 12216
rect 13176 12048 13210 12082
rect 14655 12048 14689 12148
rect 13176 12014 13248 12048
rect 13282 12014 13316 12048
rect 13350 12014 13384 12048
rect 13418 12014 13452 12048
rect 13486 12014 13520 12048
rect 13554 12014 13588 12048
rect 13622 12014 13656 12048
rect 13690 12014 13724 12048
rect 13758 12014 13792 12048
rect 13826 12014 13860 12048
rect 13894 12014 13928 12048
rect 13962 12014 13996 12048
rect 14030 12014 14064 12048
rect 14098 12014 14132 12048
rect 14166 12014 14200 12048
rect 14234 12014 14268 12048
rect 14302 12014 14336 12048
rect 14370 12014 14404 12048
rect 14438 12014 14472 12048
rect 14506 12014 14587 12048
rect 14621 12014 14689 12048
rect 4796 7463 4830 7472
rect 4796 7395 4830 7429
rect 5656 7463 5690 7472
rect 5656 7395 5690 7429
rect 4796 7327 4830 7361
rect 4796 7259 4830 7293
rect 4796 7191 4830 7225
rect 4796 7123 4830 7157
rect 4796 7055 4830 7089
rect 4796 6987 4830 7021
rect 4796 6919 4830 6953
rect 4796 6851 4830 6885
rect 6666 7463 6700 7472
rect 6666 7395 6700 7429
rect 5656 7327 5690 7361
rect 5656 7259 5690 7293
rect 5656 7191 5690 7225
rect 5656 7123 5690 7157
rect 5656 7055 5690 7089
rect 5656 6987 5690 7021
rect 5656 6919 5690 6953
rect 4796 6783 4830 6817
rect 4796 6715 4830 6749
rect 4796 6647 4830 6681
rect 4796 6579 4830 6613
rect 5656 6851 5690 6885
rect 7669 7463 7703 7472
rect 7669 7395 7703 7429
rect 6666 7327 6700 7361
rect 6666 7259 6700 7293
rect 6666 7191 6700 7225
rect 6666 7123 6700 7157
rect 6666 7055 6700 7089
rect 6666 6987 6700 7021
rect 6666 6919 6700 6953
rect 5656 6783 5690 6817
rect 5656 6715 5690 6749
rect 5656 6647 5690 6681
rect 5656 6579 5690 6613
rect 6666 6851 6700 6885
rect 7669 7327 7703 7361
rect 7669 7259 7703 7293
rect 7669 7191 7703 7225
rect 7669 7123 7703 7157
rect 7669 7055 7703 7089
rect 7669 6987 7703 7021
rect 7669 6919 7703 6953
rect 6666 6783 6700 6817
rect 6666 6715 6700 6749
rect 6666 6647 6700 6681
rect 6666 6579 6700 6613
rect 7669 6851 7703 6885
rect 7669 6783 7703 6817
rect 7669 6715 7703 6749
rect 7669 6647 7703 6681
rect 7669 6579 7703 6613
rect 3998 6545 4032 6579
rect 4066 6545 4100 6579
rect 4134 6545 4168 6579
rect 4202 6545 4236 6579
rect 4270 6545 4304 6579
rect 4338 6545 4372 6579
rect 4406 6545 4440 6579
rect 4474 6545 4508 6579
rect 4542 6545 4576 6579
rect 4610 6545 4644 6579
rect 4678 6545 4712 6579
rect 4746 6545 4780 6579
rect 4814 6545 4848 6579
rect 4882 6545 4916 6579
rect 4950 6545 4984 6579
rect 5018 6545 5052 6579
rect 5086 6545 5120 6579
rect 5154 6545 5188 6579
rect 5222 6545 5256 6579
rect 5290 6545 5324 6579
rect 5358 6545 5392 6579
rect 5426 6545 5460 6579
rect 5494 6545 5528 6579
rect 5562 6545 5596 6579
rect 5630 6545 5664 6579
rect 5698 6545 5732 6579
rect 5766 6545 5800 6579
rect 5834 6545 5868 6579
rect 5902 6545 5936 6579
rect 5970 6545 6004 6579
rect 6038 6545 6072 6579
rect 6106 6545 6140 6579
rect 6174 6545 6208 6579
rect 6242 6545 6276 6579
rect 6310 6545 6344 6579
rect 6378 6545 6412 6579
rect 6446 6545 6480 6579
rect 6514 6545 6548 6579
rect 6582 6545 6616 6579
rect 6650 6545 6684 6579
rect 6718 6545 6752 6579
rect 6786 6545 6820 6579
rect 6854 6545 6888 6579
rect 6922 6545 6956 6579
rect 6990 6545 7024 6579
rect 7058 6545 7092 6579
rect 7126 6545 7160 6579
rect 7194 6545 7228 6579
rect 7262 6545 7296 6579
rect 7330 6545 7364 6579
rect 7398 6545 7432 6579
rect 7466 6545 7500 6579
rect 7534 6545 7568 6579
rect 7602 6545 7636 6579
rect 7670 6545 7704 6579
rect 7738 6545 7772 6579
rect 7806 6545 7840 6579
rect 7874 6545 7908 6579
rect 7942 6545 7976 6579
rect 8010 6545 8044 6579
rect 8078 6545 8112 6579
rect 8146 6545 8180 6579
rect 8214 6545 8248 6579
rect 8282 6545 8316 6579
rect 8350 6545 8384 6579
rect 8418 6545 8452 6579
rect 8486 6545 8520 6579
rect 8554 6545 8588 6579
rect 8622 6545 8656 6579
rect 8690 6545 8724 6579
rect 8758 6545 8792 6579
rect 8826 6545 8860 6579
rect 8894 6545 8928 6579
rect 8962 6545 8996 6579
rect 9030 6545 9064 6579
rect 9098 6545 9132 6579
rect 9166 6545 9200 6579
rect 9234 6545 9268 6579
rect 9302 6545 9336 6579
rect 9370 6545 9404 6579
rect 9438 6545 9472 6579
rect 9506 6545 9540 6579
rect 9574 6545 9608 6579
rect 9642 6545 9676 6579
rect 9710 6545 9744 6579
rect 9778 6545 9812 6579
rect 9846 6545 9880 6579
rect 9914 6545 9948 6579
rect 9982 6545 10016 6579
rect 10050 6545 10084 6579
rect 10118 6545 10152 6579
rect 10186 6545 10220 6579
rect 10254 6545 10288 6579
rect 10322 6545 10356 6579
rect 10390 6545 10424 6579
rect 10458 6545 10492 6579
rect 10526 6545 10560 6579
rect 10594 6545 10628 6579
rect 10662 6545 10696 6579
rect 10730 6545 10764 6579
rect 10798 6545 10832 6579
rect 10866 6545 10900 6579
rect 10934 6545 10968 6579
rect 11002 6545 11036 6579
rect 11070 6545 11104 6579
rect 11138 6545 11172 6579
rect 11206 6545 11240 6579
rect 11274 6545 11308 6579
rect 11342 6545 11376 6579
rect 11410 6545 11444 6579
rect 11478 6545 11512 6579
rect 11546 6545 11580 6579
rect 11614 6545 11648 6579
rect 11682 6545 11716 6579
rect 11750 6545 11784 6579
rect 11818 6545 11852 6579
rect 11886 6545 11920 6579
rect 11954 6545 12046 6579
<< mvnsubdiff >>
rect 7823 8219 12931 8220
rect 7823 8185 7857 8219
rect 7891 8185 7925 8219
rect 7959 8185 7993 8219
rect 8027 8185 8061 8219
rect 8095 8185 8129 8219
rect 8163 8185 8197 8219
rect 8231 8185 8265 8219
rect 8299 8185 8333 8219
rect 8367 8185 8401 8219
rect 8435 8185 8469 8219
rect 8503 8185 8537 8219
rect 8571 8185 8605 8219
rect 8639 8185 8673 8219
rect 8707 8185 8741 8219
rect 8775 8185 8809 8219
rect 8843 8185 8877 8219
rect 8911 8185 8945 8219
rect 8979 8185 9013 8219
rect 9047 8185 9081 8219
rect 9115 8185 9149 8219
rect 9183 8185 9217 8219
rect 9251 8185 9285 8219
rect 9319 8185 9353 8219
rect 9387 8185 9421 8219
rect 9455 8185 9489 8219
rect 9523 8185 9557 8219
rect 9591 8185 9625 8219
rect 9659 8185 9693 8219
rect 9727 8185 9761 8219
rect 9795 8185 9829 8219
rect 9863 8185 9897 8219
rect 9931 8185 9965 8219
rect 9999 8185 10033 8219
rect 10067 8185 10101 8219
rect 10135 8185 10169 8219
rect 10203 8185 10237 8219
rect 10271 8185 10305 8219
rect 10339 8185 10373 8219
rect 10407 8185 10441 8219
rect 10475 8185 10509 8219
rect 10543 8185 10577 8219
rect 10611 8185 10645 8219
rect 10679 8185 10713 8219
rect 10747 8185 10781 8219
rect 10815 8185 10849 8219
rect 10883 8185 10917 8219
rect 10951 8185 10985 8219
rect 11019 8185 11053 8219
rect 11087 8185 11121 8219
rect 11155 8185 11189 8219
rect 11223 8185 11257 8219
rect 11291 8185 11325 8219
rect 11359 8185 11393 8219
rect 11427 8185 11461 8219
rect 11495 8185 11529 8219
rect 11563 8185 11597 8219
rect 11631 8185 11665 8219
rect 11699 8185 11733 8219
rect 11767 8185 11801 8219
rect 11835 8185 11869 8219
rect 11903 8185 11937 8219
rect 11971 8185 12005 8219
rect 12039 8185 12073 8219
rect 12107 8185 12141 8219
rect 12175 8185 12209 8219
rect 12243 8185 12277 8219
rect 12311 8185 12345 8219
rect 12379 8185 12413 8219
rect 12447 8185 12481 8219
rect 12515 8185 12549 8219
rect 12583 8185 12617 8219
rect 12651 8185 12685 8219
rect 12719 8185 12753 8219
rect 12787 8185 12821 8219
rect 12855 8186 12931 8219
rect 12855 8185 12896 8186
rect 7823 8184 12896 8185
rect 7823 8151 7859 8184
rect 7823 8117 7824 8151
rect 7858 8117 7859 8151
rect 7823 8083 7859 8117
rect 7823 8049 7824 8083
rect 7858 8049 7859 8083
rect 7823 8015 7859 8049
rect 12895 8152 12896 8184
rect 12930 8152 12931 8186
rect 12895 8118 12931 8152
rect 12895 8084 12896 8118
rect 12930 8084 12931 8118
rect 12895 8050 12931 8084
rect 7823 7981 7824 8015
rect 7858 7981 7859 8015
rect 12895 8016 12896 8050
rect 12930 8016 12931 8050
rect 7823 7947 7859 7981
rect 7823 7913 7824 7947
rect 7858 7913 7859 7947
rect 7823 7879 7859 7913
rect 7823 7845 7824 7879
rect 7858 7845 7859 7879
rect 12895 7982 12931 8016
rect 12895 7948 12896 7982
rect 12930 7948 12931 7982
rect 12895 7914 12931 7948
rect 12895 7880 12896 7914
rect 12930 7880 12931 7914
rect 12895 7846 12931 7880
rect 7823 7811 7859 7845
rect 7823 7777 7824 7811
rect 7858 7777 7859 7811
rect 7823 7743 7859 7777
rect 7823 7709 7824 7743
rect 7858 7709 7859 7743
rect 7823 7675 7859 7709
rect 7823 7641 7824 7675
rect 7858 7641 7859 7675
rect 12895 7812 12896 7846
rect 12930 7812 12931 7846
rect 12895 7778 12931 7812
rect 12895 7744 12896 7778
rect 12930 7744 12931 7778
rect 12895 7710 12931 7744
rect 12895 7676 12896 7710
rect 12930 7676 12931 7710
rect 7823 7607 7859 7641
rect 12895 7642 12931 7676
rect 7823 7575 7824 7607
rect 3894 7574 7824 7575
rect 3894 7540 3928 7574
rect 3962 7540 3996 7574
rect 4030 7540 4064 7574
rect 4098 7540 4132 7574
rect 4166 7540 4200 7574
rect 4234 7540 4268 7574
rect 4302 7540 4336 7574
rect 4370 7540 4404 7574
rect 4438 7540 4472 7574
rect 4506 7540 4540 7574
rect 4574 7540 4608 7574
rect 4642 7540 4676 7574
rect 4710 7540 4744 7574
rect 4778 7540 4812 7574
rect 4846 7540 4880 7574
rect 4914 7540 4948 7574
rect 4982 7540 5016 7574
rect 5050 7540 5084 7574
rect 5118 7540 5152 7574
rect 5186 7540 5220 7574
rect 5254 7540 5288 7574
rect 5322 7540 5356 7574
rect 5390 7540 5424 7574
rect 5458 7540 5492 7574
rect 5526 7540 5560 7574
rect 5594 7540 5628 7574
rect 5662 7540 5696 7574
rect 5730 7540 5764 7574
rect 5798 7540 5832 7574
rect 5866 7540 5900 7574
rect 5934 7540 5968 7574
rect 6002 7540 6036 7574
rect 6070 7540 6104 7574
rect 6138 7540 6172 7574
rect 6206 7540 6240 7574
rect 6274 7540 6308 7574
rect 6342 7540 6376 7574
rect 6410 7540 6444 7574
rect 6478 7540 6512 7574
rect 6546 7540 6580 7574
rect 6614 7540 6648 7574
rect 6682 7540 6716 7574
rect 6750 7540 6784 7574
rect 6818 7540 6852 7574
rect 6886 7540 6920 7574
rect 6954 7540 6988 7574
rect 7022 7540 7056 7574
rect 7090 7540 7124 7574
rect 7158 7540 7192 7574
rect 7226 7540 7260 7574
rect 7294 7540 7328 7574
rect 7362 7540 7396 7574
rect 7430 7540 7464 7574
rect 7498 7540 7532 7574
rect 7566 7540 7600 7574
rect 7634 7540 7668 7574
rect 7702 7540 7736 7574
rect 7770 7573 7824 7574
rect 7858 7573 7859 7607
rect 7770 7540 7859 7573
rect 3894 7539 7859 7540
rect 3894 7495 3930 7539
rect 3894 7461 3895 7495
rect 3929 7461 3930 7495
rect 3894 7427 3930 7461
rect 3894 7393 3895 7427
rect 3929 7393 3930 7427
rect 3894 7359 3930 7393
rect 4796 7472 4830 7539
rect 3894 7325 3895 7359
rect 3929 7325 3930 7359
rect 3894 7291 3930 7325
rect 3894 7257 3895 7291
rect 3929 7257 3930 7291
rect 3894 7223 3930 7257
rect 3894 7189 3895 7223
rect 3929 7189 3930 7223
rect 3894 7155 3930 7189
rect 3894 7121 3895 7155
rect 3929 7121 3930 7155
rect 3894 7087 3930 7121
rect 3894 7053 3895 7087
rect 3929 7053 3930 7087
rect 3894 7019 3930 7053
rect 3894 6985 3895 7019
rect 3929 6985 3930 7019
rect 3894 6951 3930 6985
rect 3894 6917 3895 6951
rect 3929 6917 3930 6951
rect 3894 6883 3930 6917
rect 3894 6849 3895 6883
rect 3929 6849 3930 6883
rect 5656 7472 5690 7539
rect 3894 6815 3930 6849
rect 3894 6781 3895 6815
rect 3929 6781 3930 6815
rect 3894 6747 3930 6781
rect 3894 6713 3895 6747
rect 3929 6713 3930 6747
rect 3894 6679 3930 6713
rect 3894 6645 3895 6679
rect 3929 6645 3930 6679
rect 3894 6611 3930 6645
rect 3894 6577 3895 6611
rect 3929 6579 3930 6611
rect 6666 7472 6700 7539
rect 7669 7472 7703 7539
rect 12895 7608 12896 7642
rect 12930 7608 12931 7642
rect 12895 7574 12931 7608
rect 12895 7540 12896 7574
rect 12930 7540 12931 7574
rect 12895 7506 12931 7540
rect 12895 7472 12896 7506
rect 12930 7472 12931 7506
rect 12895 7438 12931 7472
rect 12895 7404 12896 7438
rect 12930 7404 12931 7438
rect 12895 7370 12931 7404
rect 12895 7336 12896 7370
rect 12930 7336 12931 7370
rect 12895 7302 12931 7336
rect 12895 7268 12896 7302
rect 12930 7268 12931 7302
rect 12895 7234 12931 7268
rect 12895 7200 12896 7234
rect 12930 7200 12931 7234
rect 12895 7166 12931 7200
rect 12895 7132 12896 7166
rect 12930 7132 12931 7166
rect 12895 7098 12931 7132
rect 12895 7064 12896 7098
rect 12930 7064 12931 7098
rect 12895 7030 12931 7064
rect 12895 6996 12896 7030
rect 12930 6996 12931 7030
rect 12895 6962 12931 6996
rect 12895 6928 12896 6962
rect 12930 6928 12931 6962
rect 12895 6894 12931 6928
rect 12895 6860 12896 6894
rect 12930 6860 12931 6894
rect 12895 6826 12931 6860
rect 12895 6792 12896 6826
rect 12930 6792 12931 6826
rect 12895 6758 12931 6792
rect 12895 6724 12896 6758
rect 12930 6724 12931 6758
rect 12895 6690 12931 6724
rect 12895 6656 12896 6690
rect 12930 6656 12931 6690
rect 12895 6622 12931 6656
rect 12895 6588 12896 6622
rect 12930 6588 12931 6622
rect 3929 6577 3964 6579
rect 3894 6545 3964 6577
rect 12895 6554 12931 6588
rect 3894 6543 3930 6545
rect 3894 6509 3895 6543
rect 3929 6509 3930 6543
rect 3894 6475 3930 6509
rect 3894 6441 3895 6475
rect 3929 6441 3930 6475
rect 3894 6407 3930 6441
rect 3894 6373 3895 6407
rect 3929 6373 3930 6407
rect 3894 6339 3930 6373
rect 12895 6520 12896 6554
rect 12930 6520 12931 6554
rect 12895 6486 12931 6520
rect 12895 6452 12896 6486
rect 12930 6452 12931 6486
rect 12895 6354 12931 6452
rect 3894 6305 3895 6339
rect 3929 6305 3930 6339
rect 3894 6271 3930 6305
rect 3894 6237 3895 6271
rect 3929 6237 3930 6271
rect 3894 6203 3930 6237
rect 3894 6169 3895 6203
rect 3929 6169 3930 6203
rect 3894 6135 3930 6169
rect 3894 6101 3895 6135
rect 3929 6101 3930 6135
rect 3894 6067 3930 6101
rect 3894 6033 3895 6067
rect 3929 6033 3930 6067
rect 3894 5999 3930 6033
rect 3894 5965 3895 5999
rect 3929 5965 3930 5999
rect 3894 5931 3930 5965
rect 3894 5897 3895 5931
rect 3929 5897 3930 5931
rect 3894 5863 3930 5897
rect 3894 5829 3895 5863
rect 3929 5829 3930 5863
rect 3894 5795 3930 5829
rect 3894 5761 3895 5795
rect 3929 5761 3930 5795
rect 3894 5727 3930 5761
rect 3894 5693 3895 5727
rect 3929 5693 3930 5727
rect 12194 6353 12931 6354
rect 12194 6320 12319 6353
rect 12194 6286 12195 6320
rect 12229 6319 12319 6320
rect 12353 6319 12387 6353
rect 12421 6319 12455 6353
rect 12489 6319 12523 6353
rect 12557 6319 12591 6353
rect 12625 6319 12659 6353
rect 12693 6319 12727 6353
rect 12761 6319 12795 6353
rect 12829 6319 12863 6353
rect 12897 6319 12931 6353
rect 12229 6318 12931 6319
rect 12229 6286 12230 6318
rect 12194 6252 12230 6286
rect 12194 6218 12195 6252
rect 12229 6218 12230 6252
rect 12194 6184 12230 6218
rect 12194 6150 12195 6184
rect 12229 6150 12230 6184
rect 12194 6116 12230 6150
rect 12194 6082 12195 6116
rect 12229 6082 12230 6116
rect 12194 6048 12230 6082
rect 12194 6014 12195 6048
rect 12229 6014 12230 6048
rect 12194 5980 12230 6014
rect 12194 5946 12195 5980
rect 12229 5946 12230 5980
rect 12194 5912 12230 5946
rect 12194 5878 12195 5912
rect 12229 5878 12230 5912
rect 12194 5844 12230 5878
rect 12194 5810 12195 5844
rect 12229 5810 12230 5844
rect 12194 5776 12230 5810
rect 12194 5742 12195 5776
rect 12229 5742 12230 5776
rect 3894 5659 3930 5693
rect 3894 5625 3895 5659
rect 3929 5625 3930 5659
rect 3894 5591 3930 5625
rect 3894 5557 3895 5591
rect 3929 5557 3930 5591
rect 3894 5523 3930 5557
rect 3894 5489 3895 5523
rect 3929 5489 3930 5523
rect 3894 5455 3930 5489
rect 3894 5421 3895 5455
rect 3929 5421 3930 5455
rect 3894 5387 3930 5421
rect 3894 5353 3895 5387
rect 3929 5353 3930 5387
rect 3894 5319 3930 5353
rect 3894 5285 3895 5319
rect 3929 5285 3930 5319
rect 3894 5251 3930 5285
rect 3894 5217 3895 5251
rect 3929 5217 3930 5251
rect 3894 5183 3930 5217
rect 3894 5149 3895 5183
rect 3929 5149 3930 5183
rect 3894 5115 3930 5149
rect 3894 5081 3895 5115
rect 3929 5081 3930 5115
rect 3894 5047 3930 5081
rect 3894 5013 3895 5047
rect 3929 5013 3930 5047
rect 3894 4979 3930 5013
rect 3894 4945 3895 4979
rect 3929 4945 3930 4979
rect 3894 4911 3930 4945
rect 3894 4877 3895 4911
rect 3929 4877 3930 4911
rect 3894 4843 3930 4877
rect 3894 4809 3895 4843
rect 3929 4809 3930 4843
rect 3894 4775 3930 4809
rect 3894 4741 3895 4775
rect 3929 4741 3930 4775
rect 3894 4707 3930 4741
rect 3894 4673 3895 4707
rect 3929 4673 3930 4707
rect 3894 4639 3930 4673
rect 3894 4605 3895 4639
rect 3929 4605 3930 4639
rect 3894 4571 3930 4605
rect 3894 4537 3895 4571
rect 3929 4537 3930 4571
rect 3894 4503 3930 4537
rect 3894 4469 3895 4503
rect 3929 4469 3930 4503
rect 3894 4435 3930 4469
rect 3894 4401 3895 4435
rect 3929 4401 3930 4435
rect 3894 4367 3930 4401
rect 3894 4333 3895 4367
rect 3929 4333 3930 4367
rect 3894 4299 3930 4333
rect 3894 4265 3895 4299
rect 3929 4265 3930 4299
rect 3894 4231 3930 4265
rect 3894 4197 3895 4231
rect 3929 4197 3930 4231
rect 3894 4163 3930 4197
rect 3894 4129 3895 4163
rect 3929 4129 3930 4163
rect 3894 4095 3930 4129
rect 3894 4061 3895 4095
rect 3929 4061 3930 4095
rect 3894 4027 3930 4061
rect 3894 3993 3895 4027
rect 3929 3993 3930 4027
rect 3894 3959 3930 3993
rect 3894 3925 3895 3959
rect 3929 3925 3930 3959
rect 3894 3891 3930 3925
rect 3894 3857 3895 3891
rect 3929 3857 3930 3891
rect 3894 3823 3930 3857
rect 3894 3789 3895 3823
rect 3929 3789 3930 3823
rect 3894 3755 3930 3789
rect 3894 3721 3895 3755
rect 3929 3721 3930 3755
rect 3894 3687 3930 3721
rect 3894 3653 3895 3687
rect 3929 3653 3930 3687
rect 3894 3619 3930 3653
rect 3894 3585 3895 3619
rect 3929 3585 3930 3619
rect 3894 3551 3930 3585
rect 3894 3517 3895 3551
rect 3929 3517 3930 3551
rect 3894 3483 3930 3517
rect 3894 3449 3895 3483
rect 3929 3449 3930 3483
rect 3894 3415 3930 3449
rect 3894 3381 3895 3415
rect 3929 3381 3930 3415
rect 3894 3347 3930 3381
rect 3894 3313 3895 3347
rect 3929 3313 3930 3347
rect 3894 3279 3930 3313
rect 3894 3245 3895 3279
rect 3929 3245 3930 3279
rect 3894 3211 3930 3245
rect 3894 3177 3895 3211
rect 3929 3177 3930 3211
rect 3894 3143 3930 3177
rect 3894 3109 3895 3143
rect 3929 3109 3930 3143
rect 3894 3075 3930 3109
rect 3894 3041 3895 3075
rect 3929 3041 3930 3075
rect 3894 3007 3930 3041
rect 3894 2973 3895 3007
rect 3929 2973 3930 3007
rect 3894 2939 3930 2973
rect 3894 2905 3895 2939
rect 3929 2905 3930 2939
rect 3894 2871 3930 2905
rect 3894 2837 3895 2871
rect 3929 2837 3930 2871
rect 3894 2803 3930 2837
rect 3894 2769 3895 2803
rect 3929 2769 3930 2803
rect 3894 2735 3930 2769
rect 3894 2701 3895 2735
rect 3929 2701 3930 2735
rect 3894 2667 3930 2701
rect 3894 2633 3895 2667
rect 3929 2633 3930 2667
rect 3894 2599 3930 2633
rect 3894 2565 3895 2599
rect 3929 2565 3930 2599
rect 3894 2531 3930 2565
rect 3894 2497 3895 2531
rect 3929 2497 3930 2531
rect 3894 2463 3930 2497
rect 3894 2429 3895 2463
rect 3929 2429 3930 2463
rect 3894 2395 3930 2429
rect 3894 2361 3895 2395
rect 3929 2361 3930 2395
rect 3894 2327 3930 2361
rect 3894 2293 3895 2327
rect 3929 2293 3930 2327
rect 3894 2259 3930 2293
rect 3894 2225 3895 2259
rect 3929 2225 3930 2259
rect 3894 2191 3930 2225
rect 3894 2157 3895 2191
rect 3929 2157 3930 2191
rect 3894 2123 3930 2157
rect 3894 2089 3895 2123
rect 3929 2089 3930 2123
rect 3894 2055 3930 2089
rect 3894 2021 3895 2055
rect 3929 2021 3930 2055
rect 3894 1987 3930 2021
rect 3894 1953 3895 1987
rect 3929 1953 3930 1987
rect 3894 1919 3930 1953
rect 12194 5708 12230 5742
rect 12194 5674 12195 5708
rect 12229 5674 12230 5708
rect 12194 5640 12230 5674
rect 12194 5606 12195 5640
rect 12229 5606 12230 5640
rect 12194 5572 12230 5606
rect 12194 5538 12195 5572
rect 12229 5538 12230 5572
rect 12194 5504 12230 5538
rect 12194 5470 12195 5504
rect 12229 5470 12230 5504
rect 12194 5436 12230 5470
rect 12194 5402 12195 5436
rect 12229 5402 12230 5436
rect 12194 5368 12230 5402
rect 12194 5334 12195 5368
rect 12229 5334 12230 5368
rect 12194 5300 12230 5334
rect 12194 5266 12195 5300
rect 12229 5266 12230 5300
rect 12194 5232 12230 5266
rect 12194 5198 12195 5232
rect 12229 5198 12230 5232
rect 12194 5164 12230 5198
rect 12194 5130 12195 5164
rect 12229 5130 12230 5164
rect 12194 5096 12230 5130
rect 12194 5062 12195 5096
rect 12229 5062 12230 5096
rect 12194 5028 12230 5062
rect 12194 4994 12195 5028
rect 12229 4994 12230 5028
rect 12194 4960 12230 4994
rect 12194 4926 12195 4960
rect 12229 4926 12230 4960
rect 12194 4892 12230 4926
rect 12194 4858 12195 4892
rect 12229 4858 12230 4892
rect 12194 4824 12230 4858
rect 12194 4790 12195 4824
rect 12229 4790 12230 4824
rect 12194 4756 12230 4790
rect 12194 4722 12195 4756
rect 12229 4722 12230 4756
rect 12194 4688 12230 4722
rect 12194 4654 12195 4688
rect 12229 4654 12230 4688
rect 12194 4620 12230 4654
rect 12194 4586 12195 4620
rect 12229 4586 12230 4620
rect 12194 4552 12230 4586
rect 12194 4518 12195 4552
rect 12229 4518 12230 4552
rect 12194 4484 12230 4518
rect 12194 4450 12195 4484
rect 12229 4450 12230 4484
rect 12194 4416 12230 4450
rect 12194 4382 12195 4416
rect 12229 4382 12230 4416
rect 12194 4348 12230 4382
rect 12194 4314 12195 4348
rect 12229 4314 12230 4348
rect 12194 4280 12230 4314
rect 12194 4246 12195 4280
rect 12229 4246 12230 4280
rect 12194 4212 12230 4246
rect 12194 4178 12195 4212
rect 12229 4178 12230 4212
rect 12194 4144 12230 4178
rect 12194 4110 12195 4144
rect 12229 4110 12230 4144
rect 12194 4076 12230 4110
rect 12194 4042 12195 4076
rect 12229 4042 12230 4076
rect 12194 4008 12230 4042
rect 12194 3974 12195 4008
rect 12229 3974 12230 4008
rect 12194 3940 12230 3974
rect 12194 3906 12195 3940
rect 12229 3906 12230 3940
rect 12194 3872 12230 3906
rect 12194 3838 12195 3872
rect 12229 3838 12230 3872
rect 12194 3804 12230 3838
rect 12194 3770 12195 3804
rect 12229 3770 12230 3804
rect 12194 3736 12230 3770
rect 12194 3702 12195 3736
rect 12229 3702 12230 3736
rect 12194 3668 12230 3702
rect 12194 3634 12195 3668
rect 12229 3634 12230 3668
rect 12194 3600 12230 3634
rect 12194 3566 12195 3600
rect 12229 3566 12230 3600
rect 12194 3532 12230 3566
rect 12194 3498 12195 3532
rect 12229 3498 12230 3532
rect 12194 3464 12230 3498
rect 12194 3430 12195 3464
rect 12229 3430 12230 3464
rect 12194 3396 12230 3430
rect 12194 3362 12195 3396
rect 12229 3362 12230 3396
rect 12194 3328 12230 3362
rect 12194 3294 12195 3328
rect 12229 3294 12230 3328
rect 12194 3260 12230 3294
rect 12194 3226 12195 3260
rect 12229 3226 12230 3260
rect 12194 3192 12230 3226
rect 12194 3158 12195 3192
rect 12229 3158 12230 3192
rect 12194 3124 12230 3158
rect 12194 3090 12195 3124
rect 12229 3090 12230 3124
rect 12194 3056 12230 3090
rect 12194 3022 12195 3056
rect 12229 3022 12230 3056
rect 12194 2988 12230 3022
rect 12194 2954 12195 2988
rect 12229 2954 12230 2988
rect 12194 2920 12230 2954
rect 12194 2886 12195 2920
rect 12229 2886 12230 2920
rect 12194 2852 12230 2886
rect 12194 2818 12195 2852
rect 12229 2818 12230 2852
rect 12194 2784 12230 2818
rect 12194 2750 12195 2784
rect 12229 2750 12230 2784
rect 12194 2716 12230 2750
rect 12194 2682 12195 2716
rect 12229 2682 12230 2716
rect 12194 2648 12230 2682
rect 12194 2614 12195 2648
rect 12229 2614 12230 2648
rect 12194 2580 12230 2614
rect 12194 2546 12195 2580
rect 12229 2546 12230 2580
rect 12194 2512 12230 2546
rect 12194 2478 12195 2512
rect 12229 2478 12230 2512
rect 12194 2444 12230 2478
rect 12194 2410 12195 2444
rect 12229 2410 12230 2444
rect 12194 2376 12230 2410
rect 12194 2342 12195 2376
rect 12229 2342 12230 2376
rect 12194 2308 12230 2342
rect 12194 2274 12195 2308
rect 12229 2274 12230 2308
rect 12194 2240 12230 2274
rect 12194 2206 12195 2240
rect 12229 2206 12230 2240
rect 12194 2172 12230 2206
rect 12194 2138 12195 2172
rect 12229 2138 12230 2172
rect 12194 2104 12230 2138
rect 12194 2070 12195 2104
rect 12229 2070 12230 2104
rect 12194 2036 12230 2070
rect 12194 2002 12195 2036
rect 12229 2002 12230 2036
rect 12194 1968 12230 2002
rect 3894 1885 3895 1919
rect 3929 1885 3930 1919
rect 3894 1851 3930 1885
rect 3894 1817 3895 1851
rect 3929 1817 3930 1851
rect 3894 1783 3930 1817
rect 3894 1749 3895 1783
rect 3929 1749 3930 1783
rect 3894 1715 3930 1749
rect 3894 1681 3895 1715
rect 3929 1681 3930 1715
rect 3894 1647 3930 1681
rect 3894 1613 3895 1647
rect 3929 1613 3930 1647
rect 3894 1579 3930 1613
rect 3894 1545 3895 1579
rect 3929 1545 3930 1579
rect 3894 1511 3930 1545
rect 3894 1477 3895 1511
rect 3929 1477 3930 1511
rect 3894 1443 3930 1477
rect 3894 1409 3895 1443
rect 3929 1409 3930 1443
rect 3894 1375 3930 1409
rect 3894 1341 3895 1375
rect 3929 1341 3930 1375
rect 3894 1307 3930 1341
rect 3894 1273 3895 1307
rect 3929 1273 3930 1307
rect 3894 1239 3930 1273
rect 3894 1205 3895 1239
rect 3929 1205 3930 1239
rect 3894 1171 3930 1205
rect 3894 1137 3895 1171
rect 3929 1137 3930 1171
rect 3894 1103 3930 1137
rect 3894 1069 3895 1103
rect 3929 1069 3930 1103
rect 3894 1035 3930 1069
rect 3894 1001 3895 1035
rect 3929 1001 3930 1035
rect 3894 967 3930 1001
rect 3894 933 3895 967
rect 3929 933 3930 967
rect 3894 899 3930 933
rect 3894 865 3895 899
rect 3929 867 3930 899
rect 12194 1934 12195 1968
rect 12229 1934 12230 1968
rect 12194 1900 12230 1934
rect 12194 1866 12195 1900
rect 12229 1866 12230 1900
rect 12194 1832 12230 1866
rect 12194 1798 12195 1832
rect 12229 1798 12230 1832
rect 12194 1764 12230 1798
rect 12194 1730 12195 1764
rect 12229 1730 12230 1764
rect 12194 1696 12230 1730
rect 12194 1662 12195 1696
rect 12229 1662 12230 1696
rect 12194 1628 12230 1662
rect 12194 1594 12195 1628
rect 12229 1594 12230 1628
rect 12194 1560 12230 1594
rect 12194 1526 12195 1560
rect 12229 1526 12230 1560
rect 12194 1492 12230 1526
rect 12194 1458 12195 1492
rect 12229 1458 12230 1492
rect 12194 1424 12230 1458
rect 12194 1390 12195 1424
rect 12229 1390 12230 1424
rect 12194 1356 12230 1390
rect 12194 1322 12195 1356
rect 12229 1322 12230 1356
rect 12194 1288 12230 1322
rect 12194 1254 12195 1288
rect 12229 1254 12230 1288
rect 12194 1220 12230 1254
rect 12194 1186 12195 1220
rect 12229 1186 12230 1220
rect 12194 1051 12230 1186
rect 12194 1017 12195 1051
rect 12229 1017 12230 1051
rect 12194 983 12230 1017
rect 12194 949 12195 983
rect 12229 949 12230 983
rect 12194 867 12230 949
rect 3929 866 12230 867
rect 3929 865 4002 866
rect 3894 832 4002 865
rect 4036 832 4070 866
rect 4104 832 4138 866
rect 4172 832 4206 866
rect 4240 832 4274 866
rect 4308 832 4342 866
rect 4376 832 4410 866
rect 4444 832 4478 866
rect 4512 832 4546 866
rect 4580 832 4614 866
rect 4648 832 4682 866
rect 4716 832 4750 866
rect 4784 832 4818 866
rect 4852 832 4886 866
rect 4920 832 4954 866
rect 4988 832 5022 866
rect 5056 832 5090 866
rect 5124 832 5158 866
rect 5192 832 5226 866
rect 5260 832 5294 866
rect 5328 832 5362 866
rect 5396 832 5430 866
rect 5464 832 5498 866
rect 5532 832 5566 866
rect 5600 832 5634 866
rect 5668 832 5702 866
rect 5736 832 5770 866
rect 5804 832 5838 866
rect 5872 832 5906 866
rect 5940 832 5974 866
rect 6008 832 6042 866
rect 6076 832 6110 866
rect 6144 832 6178 866
rect 6212 832 6246 866
rect 6280 832 6314 866
rect 6348 832 6382 866
rect 6416 832 6450 866
rect 6484 832 6518 866
rect 6552 832 6586 866
rect 6620 832 6654 866
rect 6688 832 6722 866
rect 6756 832 6790 866
rect 6824 832 6858 866
rect 6892 832 6926 866
rect 6960 832 6994 866
rect 7028 832 7062 866
rect 7096 832 7130 866
rect 7164 832 7198 866
rect 7232 832 7266 866
rect 7300 832 7334 866
rect 7368 832 7402 866
rect 7436 832 7470 866
rect 7504 832 7538 866
rect 7572 832 7606 866
rect 7640 832 7674 866
rect 7708 832 7742 866
rect 7776 832 7810 866
rect 7844 832 7878 866
rect 7912 832 7946 866
rect 7980 832 8014 866
rect 8048 832 8082 866
rect 8116 832 8150 866
rect 8184 832 8218 866
rect 8252 832 8286 866
rect 8320 832 8354 866
rect 8388 832 8422 866
rect 8456 832 8490 866
rect 8524 832 8558 866
rect 8592 832 8626 866
rect 8660 832 8694 866
rect 8728 832 8762 866
rect 8796 832 8830 866
rect 8864 832 8898 866
rect 8932 832 8966 866
rect 9000 832 9034 866
rect 9068 832 9102 866
rect 9136 832 9170 866
rect 9204 832 9238 866
rect 9272 832 9306 866
rect 9340 832 9374 866
rect 9408 832 9442 866
rect 9476 832 9510 866
rect 9544 832 9578 866
rect 9612 832 9646 866
rect 9680 832 9714 866
rect 9748 832 9782 866
rect 9816 832 9850 866
rect 9884 832 9918 866
rect 9952 832 9986 866
rect 10020 832 10054 866
rect 10088 832 10122 866
rect 10156 832 10190 866
rect 10224 832 10258 866
rect 10292 832 10326 866
rect 10360 832 10394 866
rect 10428 832 10462 866
rect 10496 832 10530 866
rect 10564 832 10598 866
rect 10632 832 10666 866
rect 10700 832 10734 866
rect 10768 832 10802 866
rect 10836 832 10870 866
rect 10904 832 10938 866
rect 10972 832 11006 866
rect 11040 832 11074 866
rect 11108 832 11142 866
rect 11176 832 11210 866
rect 11244 832 11278 866
rect 11312 832 11346 866
rect 11380 832 11414 866
rect 11448 832 11482 866
rect 11516 832 11550 866
rect 11584 832 11618 866
rect 11652 832 11686 866
rect 11720 832 11754 866
rect 11788 832 11822 866
rect 11856 832 11890 866
rect 11924 832 11958 866
rect 11992 832 12026 866
rect 12060 832 12094 866
rect 12128 832 12162 866
rect 12196 832 12230 866
rect 3894 831 12230 832
<< psubdiffcont >>
rect 3147 14614 3181 14648
rect 3215 14614 3249 14648
rect 3283 14614 3317 14648
rect 3351 14614 3385 14648
rect 3419 14614 3453 14648
rect 3487 14614 3521 14648
rect 3555 14614 3589 14648
rect 3623 14614 3657 14648
rect 3691 14614 3725 14648
rect 3759 14614 3793 14648
rect 3827 14614 3861 14648
rect 3895 14614 3929 14648
rect 3963 14614 3997 14648
rect 4031 14614 4065 14648
rect 4099 14614 4133 14648
rect 4167 14614 4201 14648
rect 4235 14614 4269 14648
rect 4303 14614 4337 14648
rect 4371 14614 4405 14648
rect 4439 14614 4473 14648
rect 4507 14614 4541 14648
rect 4575 14614 4609 14648
rect 4643 14614 4677 14648
rect 4711 14614 4745 14648
rect 4779 14614 4813 14648
rect 4847 14614 4881 14648
rect 4915 14614 4949 14648
rect 4983 14614 5017 14648
rect 3079 14524 3113 14558
rect 3079 14456 3113 14490
rect 5087 14546 5121 14580
rect 5087 14478 5121 14512
rect 3079 14388 3113 14422
rect 3079 14320 3113 14354
rect 3079 14252 3113 14286
rect 3079 14184 3113 14218
rect 3079 14116 3113 14150
rect 3079 14048 3113 14082
rect 3079 13980 3113 14014
rect 3079 13912 3113 13946
rect 3079 13844 3113 13878
rect 3079 13776 3113 13810
rect 3079 13708 3113 13742
rect 3079 13640 3113 13674
rect 3079 13572 3113 13606
rect 3079 13504 3113 13538
rect 3079 13436 3113 13470
rect 3079 13368 3113 13402
rect 3079 13300 3113 13334
rect 3079 13232 3113 13266
rect 3079 13164 3113 13198
rect 3079 13096 3113 13130
rect 3079 13028 3113 13062
rect 3079 12960 3113 12994
rect 5087 14410 5121 14444
rect 5087 14342 5121 14376
rect 5087 14274 5121 14308
rect 5087 14206 5121 14240
rect 5087 14138 5121 14172
rect 5087 14070 5121 14104
rect 5087 14002 5121 14036
rect 5087 13934 5121 13968
rect 5087 13866 5121 13900
rect 5087 13798 5121 13832
rect 5087 13730 5121 13764
rect 5087 13662 5121 13696
rect 5087 13594 5121 13628
rect 5087 13526 5121 13560
rect 5087 13458 5121 13492
rect 5087 13390 5121 13424
rect 5087 13322 5121 13356
rect 5087 13254 5121 13288
rect 5087 13186 5121 13220
rect 5087 13118 5121 13152
rect 5087 13050 5121 13084
rect 3079 12892 3113 12926
rect 5087 12982 5121 13016
rect 5087 12914 5121 12948
rect 3079 12824 3113 12858
rect 3079 12756 3113 12790
rect 3079 12688 3113 12722
rect 3079 12542 3113 12576
rect 3079 12474 3113 12508
rect 3079 12406 3113 12440
rect 5087 12846 5121 12880
rect 5087 12778 5121 12812
rect 5087 12710 5121 12744
rect 5087 12642 5121 12676
rect 5087 12574 5121 12608
rect 5087 12506 5121 12540
rect 5087 12438 5121 12472
rect 5478 14307 5512 14341
rect 5546 14307 5580 14341
rect 5614 14307 5648 14341
rect 5682 14307 5716 14341
rect 5750 14307 5784 14341
rect 5818 14307 5852 14341
rect 5886 14307 5920 14341
rect 5954 14307 5988 14341
rect 6022 14307 6056 14341
rect 6090 14307 6124 14341
rect 6158 14307 6192 14341
rect 6226 14307 6260 14341
rect 6294 14307 6328 14341
rect 6362 14307 6396 14341
rect 6430 14307 6464 14341
rect 6498 14307 6532 14341
rect 6566 14307 6600 14341
rect 6634 14307 6668 14341
rect 6702 14307 6736 14341
rect 6770 14307 6804 14341
rect 6838 14307 6872 14341
rect 6906 14307 6940 14341
rect 6974 14307 7008 14341
rect 7042 14307 7076 14341
rect 7110 14307 7144 14341
rect 7178 14307 7212 14341
rect 7246 14307 7280 14341
rect 7314 14307 7348 14341
rect 7382 14307 7416 14341
rect 7450 14307 7484 14341
rect 7518 14307 7552 14341
rect 7586 14307 7620 14341
rect 7654 14307 7688 14341
rect 7722 14307 7756 14341
rect 7790 14307 7824 14341
rect 7858 14307 7892 14341
rect 7926 14307 7960 14341
rect 7994 14307 8028 14341
rect 8062 14307 8096 14341
rect 8130 14307 8164 14341
rect 8198 14307 8232 14341
rect 8266 14307 8300 14341
rect 8334 14307 8368 14341
rect 8402 14307 8436 14341
rect 8470 14307 8504 14341
rect 8538 14307 8572 14341
rect 8606 14307 8640 14341
rect 8674 14307 8708 14341
rect 8742 14307 8776 14341
rect 8810 14307 8844 14341
rect 8878 14307 8912 14341
rect 8946 14307 8980 14341
rect 9014 14307 9048 14341
rect 9082 14307 9116 14341
rect 9150 14307 9184 14341
rect 5410 14207 5444 14241
rect 5410 14139 5444 14173
rect 9231 14239 9265 14273
rect 9231 14171 9265 14205
rect 5410 14071 5444 14105
rect 9231 14103 9265 14137
rect 5410 14003 5444 14037
rect 5410 13935 5444 13969
rect 5410 13867 5444 13901
rect 9231 14035 9265 14069
rect 9231 13967 9265 14001
rect 9231 13899 9265 13933
rect 5410 13799 5444 13833
rect 5410 13731 5444 13765
rect 9231 13831 9265 13865
rect 9231 13763 9265 13797
rect 5410 13663 5444 13697
rect 9231 13695 9265 13729
rect 5410 13595 5444 13629
rect 5410 13527 5444 13561
rect 5410 13459 5444 13493
rect 5410 13391 5444 13425
rect 5410 13323 5444 13357
rect 5410 13255 5444 13289
rect 5410 13187 5444 13221
rect 5410 13119 5444 13153
rect 5410 13051 5444 13085
rect 5410 12983 5444 13017
rect 5410 12915 5444 12949
rect 5410 12847 5444 12881
rect 5410 12779 5444 12813
rect 5410 12711 5444 12745
rect 5410 12643 5444 12677
rect 9231 13627 9265 13661
rect 9231 13559 9265 13593
rect 9231 13491 9265 13525
rect 9231 13423 9265 13457
rect 9231 13355 9265 13389
rect 9231 13287 9265 13321
rect 9231 13219 9265 13253
rect 9231 13151 9265 13185
rect 9231 13083 9265 13117
rect 9231 13015 9265 13049
rect 9231 12947 9265 12981
rect 9231 12879 9265 12913
rect 9231 12811 9265 12845
rect 9231 12743 9265 12777
rect 9231 12675 9265 12709
rect 5410 12575 5444 12609
rect 9231 12607 9265 12641
rect 5410 12507 5444 12541
rect 9231 12539 9265 12573
rect 5524 12439 5558 12473
rect 5592 12439 5626 12473
rect 5660 12439 5694 12473
rect 5728 12439 5762 12473
rect 5796 12439 5830 12473
rect 5864 12439 5898 12473
rect 5932 12439 5966 12473
rect 6000 12439 6034 12473
rect 6068 12439 6102 12473
rect 6136 12439 6170 12473
rect 6204 12439 6238 12473
rect 6272 12439 6306 12473
rect 6340 12439 6374 12473
rect 6408 12439 6442 12473
rect 6476 12439 6510 12473
rect 6544 12439 6578 12473
rect 6612 12439 6646 12473
rect 6680 12439 6714 12473
rect 6748 12439 6782 12473
rect 6816 12439 6850 12473
rect 6884 12439 6918 12473
rect 6952 12439 6986 12473
rect 7020 12439 7054 12473
rect 7088 12439 7122 12473
rect 7156 12439 7190 12473
rect 7224 12439 7258 12473
rect 7292 12439 7326 12473
rect 7360 12439 7394 12473
rect 7428 12439 7462 12473
rect 7496 12439 7530 12473
rect 7564 12439 7598 12473
rect 7632 12439 7666 12473
rect 7700 12439 7734 12473
rect 7768 12439 7802 12473
rect 7836 12439 7870 12473
rect 7939 12439 7973 12473
rect 8007 12439 8041 12473
rect 8075 12439 8109 12473
rect 8143 12439 8177 12473
rect 8211 12439 8245 12473
rect 8279 12439 8313 12473
rect 8347 12439 8381 12473
rect 8415 12439 8449 12473
rect 8483 12439 8517 12473
rect 8551 12439 8585 12473
rect 8619 12439 8653 12473
rect 8687 12439 8721 12473
rect 8755 12439 8789 12473
rect 8823 12439 8857 12473
rect 8891 12439 8925 12473
rect 8959 12439 8993 12473
rect 9027 12439 9061 12473
rect 9095 12439 9129 12473
rect 9163 12439 9197 12473
rect 11771 13572 11805 13606
rect 11839 13572 11873 13606
rect 11907 13572 11941 13606
rect 11975 13572 12009 13606
rect 12043 13572 12077 13606
rect 12111 13572 12145 13606
rect 12179 13572 12213 13606
rect 12247 13572 12281 13606
rect 12315 13572 12349 13606
rect 12383 13572 12417 13606
rect 12451 13572 12485 13606
rect 12519 13572 12553 13606
rect 12587 13572 12621 13606
rect 12655 13572 12689 13606
rect 12723 13572 12757 13606
rect 11686 13504 11720 13538
rect 11686 13436 11720 13470
rect 12791 13451 12825 13485
rect 11686 13368 11720 13402
rect 11686 13300 11720 13334
rect 11686 13232 11720 13266
rect 11686 13164 11720 13198
rect 11686 13096 11720 13130
rect 11686 13028 11720 13062
rect 11686 12960 11720 12994
rect 11686 12892 11720 12926
rect 11686 12824 11720 12858
rect 11686 12756 11720 12790
rect 11686 12688 11720 12722
rect 11686 12620 11720 12654
rect 11686 12552 11720 12586
rect 11686 12484 11720 12518
rect 3079 12338 3113 12372
rect 5087 12370 5121 12404
rect 3079 12270 3113 12304
rect 3079 12202 3113 12236
rect 3079 12134 3113 12168
rect 3079 12066 3113 12100
rect 5087 12302 5121 12336
rect 5087 12234 5121 12268
rect 5087 12166 5121 12200
rect 5087 12098 5121 12132
rect 3079 11998 3113 12032
rect 3079 11930 3113 11964
rect 5087 12030 5121 12064
rect 5087 11962 5121 11996
rect 3183 11862 3217 11896
rect 3251 11862 3285 11896
rect 3319 11862 3353 11896
rect 3387 11862 3421 11896
rect 3455 11862 3489 11896
rect 3523 11862 3557 11896
rect 3591 11862 3625 11896
rect 3659 11862 3693 11896
rect 3727 11862 3761 11896
rect 3795 11862 3829 11896
rect 3863 11862 3897 11896
rect 3931 11862 3965 11896
rect 3999 11862 4033 11896
rect 4067 11862 4101 11896
rect 4135 11862 4169 11896
rect 4203 11862 4237 11896
rect 4271 11862 4305 11896
rect 4339 11862 4373 11896
rect 4407 11862 4441 11896
rect 4475 11862 4509 11896
rect 4543 11862 4577 11896
rect 4611 11862 4645 11896
rect 4679 11862 4713 11896
rect 4747 11862 4781 11896
rect 4815 11862 4849 11896
rect 4883 11862 4917 11896
rect 4951 11862 4985 11896
rect 5019 11862 5053 11896
rect 11686 12416 11720 12450
rect 11686 12348 11720 12382
rect 11686 12280 11720 12314
rect 11686 12212 11720 12246
rect 11686 12144 11720 12178
rect 11686 12076 11720 12110
rect 12791 13383 12825 13417
rect 12791 13315 12825 13349
rect 12791 13247 12825 13281
rect 12791 13179 12825 13213
rect 12791 13111 12825 13145
rect 12791 13043 12825 13077
rect 12791 12975 12825 13009
rect 12791 12907 12825 12941
rect 12791 12839 12825 12873
rect 12791 12771 12825 12805
rect 12791 12703 12825 12737
rect 12791 12635 12825 12669
rect 12791 12567 12825 12601
rect 12791 12499 12825 12533
rect 12791 12431 12825 12465
rect 12791 12363 12825 12397
rect 12791 12295 12825 12329
rect 12791 12227 12825 12261
rect 12791 12159 12825 12193
rect 12791 12091 12825 12125
rect 11686 12008 11720 12042
rect 12791 12023 12825 12057
rect 12791 11955 12825 11989
rect 11754 11887 11788 11921
rect 11822 11887 11856 11921
rect 11890 11887 11924 11921
rect 11958 11887 11992 11921
rect 12026 11887 12060 11921
rect 12094 11887 12128 11921
rect 12162 11887 12196 11921
rect 12230 11887 12264 11921
rect 12298 11887 12332 11921
rect 12366 11887 12400 11921
rect 12434 11887 12468 11921
rect 12502 11887 12536 11921
rect 12570 11887 12604 11921
rect 12638 11887 12672 11921
rect 12706 11887 12740 11921
rect 8233 7997 8267 8031
rect 8301 7997 8335 8031
rect 8369 7997 8403 8031
rect 8437 7997 8471 8031
rect 8505 7997 8539 8031
rect 8573 7997 8607 8031
rect 8641 7997 8675 8031
rect 8709 7997 8743 8031
rect 8777 7997 8811 8031
rect 8845 7997 8879 8031
rect 8913 7997 8947 8031
rect 8981 7997 9015 8031
rect 9049 7997 9083 8031
rect 9117 7997 9151 8031
rect 9185 7997 9219 8031
rect 9253 7997 9287 8031
rect 9321 7997 9355 8031
rect 9389 7997 9423 8031
rect 9457 7997 9491 8031
rect 9525 7997 9559 8031
rect 9593 7997 9627 8031
rect 9661 7997 9695 8031
rect 9729 7997 9763 8031
rect 9797 7997 9831 8031
rect 9865 7997 9899 8031
rect 9933 7997 9967 8031
rect 10001 7997 10035 8031
rect 10069 7997 10103 8031
rect 10137 7997 10171 8031
rect 10205 7997 10239 8031
rect 10273 7997 10307 8031
rect 10341 7997 10375 8031
rect 10409 7997 10443 8031
rect 10477 7997 10511 8031
rect 10545 7997 10579 8031
rect 10613 7997 10647 8031
rect 10681 7997 10715 8031
rect 10749 7997 10783 8031
rect 10817 7997 10851 8031
rect 10885 7997 10919 8031
rect 10953 7997 10987 8031
rect 11021 7997 11055 8031
rect 11089 7997 11123 8031
rect 11157 7997 11191 8031
rect 11225 7997 11259 8031
rect 11293 7997 11327 8031
rect 11361 7997 11395 8031
rect 11429 7997 11463 8031
rect 11497 7997 11531 8031
rect 11565 7997 11599 8031
rect 11633 7997 11667 8031
rect 11701 7997 11735 8031
rect 11769 7997 11803 8031
rect 11837 7997 11871 8031
rect 11905 7997 11939 8031
rect 11973 7997 12007 8031
rect 12041 7997 12075 8031
rect 12109 7997 12143 8031
rect 12177 7997 12211 8031
rect 12245 7997 12279 8031
rect 12313 7997 12347 8031
rect 4180 7352 4214 7386
rect 4248 7352 4282 7386
rect 4316 7352 4350 7386
rect 4384 7352 4418 7386
rect 4452 7352 4486 7386
rect 4520 7352 4554 7386
rect 4108 7284 4142 7318
rect 4108 7216 4142 7250
rect 4588 7265 4622 7299
rect 4108 7148 4142 7182
rect 4108 7080 4142 7114
rect 4108 7012 4142 7046
rect 4588 7197 4622 7231
rect 4588 7129 4622 7163
rect 4588 7061 4622 7095
rect 4108 6944 4142 6978
rect 4588 6993 4622 7027
rect 4588 6925 4622 6959
rect 4176 6857 4210 6891
rect 4244 6857 4278 6891
rect 4312 6857 4346 6891
rect 4380 6857 4414 6891
rect 4448 6857 4482 6891
rect 5060 7352 5094 7386
rect 5128 7352 5162 7386
rect 5196 7352 5230 7386
rect 5264 7352 5298 7386
rect 5332 7352 5366 7386
rect 5400 7352 5434 7386
rect 4988 7284 5022 7318
rect 4988 7216 5022 7250
rect 5468 7265 5502 7299
rect 4988 7148 5022 7182
rect 4988 7080 5022 7114
rect 4988 7012 5022 7046
rect 5468 7197 5502 7231
rect 5468 7129 5502 7163
rect 5468 7061 5502 7095
rect 4988 6944 5022 6978
rect 5468 6993 5502 7027
rect 5468 6925 5502 6959
rect 5056 6857 5090 6891
rect 5124 6857 5158 6891
rect 5192 6857 5226 6891
rect 5260 6857 5294 6891
rect 5328 6857 5362 6891
rect 5922 7352 5956 7386
rect 5990 7352 6024 7386
rect 6058 7352 6092 7386
rect 6126 7352 6160 7386
rect 6194 7352 6228 7386
rect 6262 7352 6296 7386
rect 5850 7284 5884 7318
rect 5850 7216 5884 7250
rect 6330 7265 6364 7299
rect 5850 7148 5884 7182
rect 5850 7080 5884 7114
rect 5850 7012 5884 7046
rect 6330 7197 6364 7231
rect 6330 7129 6364 7163
rect 6330 7061 6364 7095
rect 5850 6944 5884 6978
rect 6330 6993 6364 7027
rect 6330 6925 6364 6959
rect 5918 6857 5952 6891
rect 5986 6857 6020 6891
rect 6054 6857 6088 6891
rect 6122 6857 6156 6891
rect 6190 6857 6224 6891
rect 7052 7352 7086 7386
rect 7120 7352 7154 7386
rect 7188 7352 7222 7386
rect 7256 7352 7290 7386
rect 7324 7352 7358 7386
rect 7392 7352 7426 7386
rect 6980 7284 7014 7318
rect 6980 7216 7014 7250
rect 7460 7265 7494 7299
rect 6980 7148 7014 7182
rect 6980 7080 7014 7114
rect 6980 7012 7014 7046
rect 7460 7197 7494 7231
rect 7460 7129 7494 7163
rect 7460 7061 7494 7095
rect 6980 6944 7014 6978
rect 7460 6993 7494 7027
rect 7460 6925 7494 6959
rect 7048 6857 7082 6891
rect 7116 6857 7150 6891
rect 7184 6857 7218 6891
rect 7252 6857 7286 6891
rect 7320 6857 7354 6891
rect 8233 6732 8267 6766
rect 8301 6732 8335 6766
rect 8369 6732 8403 6766
rect 8437 6732 8471 6766
rect 8505 6732 8539 6766
rect 8573 6732 8607 6766
rect 8641 6732 8675 6766
rect 8709 6732 8743 6766
rect 8777 6732 8811 6766
rect 8845 6732 8879 6766
rect 8913 6732 8947 6766
rect 8981 6732 9015 6766
rect 9049 6732 9083 6766
rect 9117 6732 9151 6766
rect 9185 6732 9219 6766
rect 9253 6732 9287 6766
rect 9321 6732 9355 6766
rect 9389 6732 9423 6766
rect 9457 6732 9491 6766
rect 9525 6732 9559 6766
rect 9593 6732 9627 6766
rect 9661 6732 9695 6766
rect 9729 6732 9763 6766
rect 9797 6732 9831 6766
rect 9865 6732 9899 6766
rect 9933 6732 9967 6766
rect 10001 6732 10035 6766
rect 10069 6732 10103 6766
rect 10137 6732 10171 6766
rect 10205 6732 10239 6766
rect 10273 6732 10307 6766
rect 10341 6732 10375 6766
rect 10409 6732 10443 6766
rect 10477 6732 10511 6766
rect 10545 6732 10579 6766
rect 10613 6732 10647 6766
rect 10681 6732 10715 6766
rect 10749 6732 10783 6766
rect 10817 6732 10851 6766
rect 10885 6732 10919 6766
rect 10953 6732 10987 6766
rect 11021 6732 11055 6766
rect 11089 6732 11123 6766
rect 11157 6732 11191 6766
rect 11225 6732 11259 6766
rect 11293 6732 11327 6766
rect 11361 6732 11395 6766
rect 11429 6732 11463 6766
rect 11497 6732 11531 6766
rect 11565 6732 11599 6766
rect 11633 6732 11667 6766
rect 11701 6732 11735 6766
rect 11769 6732 11803 6766
rect 11837 6732 11871 6766
rect 11905 6732 11939 6766
rect 11973 6732 12007 6766
rect 12041 6732 12075 6766
rect 12109 6732 12143 6766
rect 12177 6732 12211 6766
rect 12245 6732 12279 6766
rect 12313 6732 12347 6766
rect 11924 5644 11958 5678
rect 11924 5576 11958 5610
rect 11924 5508 11958 5542
rect 11924 5440 11958 5474
rect 11924 5372 11958 5406
rect 11924 5304 11958 5338
rect 11924 5236 11958 5270
rect 11924 5168 11958 5202
rect 11924 5100 11958 5134
rect 11924 5032 11958 5066
rect 11924 4964 11958 4998
rect 11924 4896 11958 4930
rect 11924 4828 11958 4862
rect 11924 4760 11958 4794
rect 11924 4692 11958 4726
rect 11924 4624 11958 4658
rect 11924 4556 11958 4590
rect 11924 4488 11958 4522
rect 11924 4420 11958 4454
rect 11924 4352 11958 4386
rect 11924 4284 11958 4318
rect 11924 4216 11958 4250
rect 11924 4148 11958 4182
rect 11924 4080 11958 4114
rect 11924 4012 11958 4046
rect 11924 3944 11958 3978
rect 11924 3876 11958 3910
rect 11924 3808 11958 3842
rect 11924 3740 11958 3774
rect 11924 3672 11958 3706
rect 11924 3604 11958 3638
rect 11924 3536 11958 3570
rect 11924 3468 11958 3502
rect 11924 3400 11958 3434
rect 11924 3332 11958 3366
rect 11924 3264 11958 3298
rect 11924 3196 11958 3230
rect 11924 3128 11958 3162
rect 11924 3060 11958 3094
rect 11924 2992 11958 3026
rect 11924 2924 11958 2958
rect 11924 2856 11958 2890
rect 11924 2788 11958 2822
rect 11924 2720 11958 2754
rect 11924 2652 11958 2686
rect 11924 2584 11958 2618
rect 11924 2516 11958 2550
rect 11924 2448 11958 2482
rect 11924 2380 11958 2414
rect 11924 2312 11958 2346
rect 11924 2244 11958 2278
rect 11924 2176 11958 2210
rect 11924 2108 11958 2142
rect 11924 2040 11958 2074
<< nsubdiffcont >>
rect 13244 14732 13278 14766
rect 13312 14732 13346 14766
rect 13380 14732 13414 14766
rect 13448 14732 13482 14766
rect 13516 14732 13550 14766
rect 13584 14732 13618 14766
rect 13652 14732 13686 14766
rect 13720 14732 13754 14766
rect 13788 14732 13822 14766
rect 13856 14732 13890 14766
rect 13924 14732 13958 14766
rect 13992 14732 14026 14766
rect 14060 14732 14094 14766
rect 14128 14732 14162 14766
rect 14196 14732 14230 14766
rect 14264 14732 14298 14766
rect 14332 14732 14366 14766
rect 14400 14732 14434 14766
rect 14468 14732 14502 14766
rect 14536 14732 14570 14766
rect -496 13376 -462 13410
rect -428 13376 -394 13410
rect -360 13376 -326 13410
rect -292 13376 -258 13410
rect -224 13376 -190 13410
rect -156 13376 -122 13410
rect -88 13376 -54 13410
rect -20 13376 14 13410
rect 48 13376 82 13410
rect 116 13376 150 13410
rect 184 13376 218 13410
rect 252 13376 286 13410
rect 320 13376 354 13410
rect -564 13264 -530 13298
rect -564 13196 -530 13230
rect -564 13128 -530 13162
rect -564 13060 -530 13094
rect -564 12992 -530 13026
rect -564 12924 -530 12958
rect -564 12856 -530 12890
rect -564 12788 -530 12822
rect -564 12720 -530 12754
rect -564 12652 -530 12686
rect -564 12584 -530 12618
rect -564 12516 -530 12550
rect -564 12448 -530 12482
rect -564 12380 -530 12414
rect -564 12312 -530 12346
rect -564 12244 -530 12278
rect -564 12176 -530 12210
rect 13176 14598 13210 14632
rect 14655 14664 14689 14698
rect 13176 14530 13210 14564
rect 14655 14596 14689 14630
rect 14655 14528 14689 14562
rect 13176 14462 13210 14496
rect 13176 14394 13210 14428
rect 13176 14326 13210 14360
rect 13176 14258 13210 14292
rect 13176 14190 13210 14224
rect 13176 14122 13210 14156
rect 13176 14054 13210 14088
rect 13176 13986 13210 14020
rect 13176 13918 13210 13952
rect 13176 13850 13210 13884
rect 13176 13782 13210 13816
rect 13176 13714 13210 13748
rect 13176 13646 13210 13680
rect -564 12108 -530 12142
rect -564 12040 -530 12074
rect 11988 13384 12022 13418
rect 12056 13384 12090 13418
rect 12124 13384 12158 13418
rect 12192 13384 12226 13418
rect 12260 13384 12294 13418
rect 12328 13384 12362 13418
rect 12396 13384 12430 13418
rect 12464 13384 12498 13418
rect 12532 13384 12566 13418
rect 11874 13316 11908 13350
rect 11874 13248 11908 13282
rect 11874 13180 11908 13214
rect 11874 13112 11908 13146
rect 11874 13044 11908 13078
rect 11874 12976 11908 13010
rect 11874 12908 11908 12942
rect 11874 12840 11908 12874
rect 11874 12772 11908 12806
rect 11874 12704 11908 12738
rect 11874 12636 11908 12670
rect 11874 12568 11908 12602
rect 11874 12500 11908 12534
rect 11874 12432 11908 12466
rect 11874 12364 11908 12398
rect 11874 12296 11908 12330
rect 11874 12228 11908 12262
rect 12600 13300 12634 13334
rect 12600 13232 12634 13266
rect 12600 13164 12634 13198
rect 12600 13096 12634 13130
rect 12600 13028 12634 13062
rect 12600 12960 12634 12994
rect 12600 12892 12634 12926
rect 12600 12824 12634 12858
rect 12600 12756 12634 12790
rect 12600 12688 12634 12722
rect 12600 12620 12634 12654
rect 12600 12552 12634 12586
rect 12600 12484 12634 12518
rect 12600 12416 12634 12450
rect 12600 12348 12634 12382
rect 12600 12280 12634 12314
rect 12600 12212 12634 12246
rect 12600 12144 12634 12178
rect 11942 12076 11976 12110
rect 12010 12076 12044 12110
rect 12078 12076 12112 12110
rect 12146 12076 12180 12110
rect 12214 12076 12248 12110
rect 12282 12076 12316 12110
rect 12350 12076 12384 12110
rect 12418 12076 12452 12110
rect 12486 12076 12520 12110
rect 13176 13578 13210 13612
rect 13176 13510 13210 13544
rect 13176 13442 13210 13476
rect 14655 14460 14689 14494
rect 14655 14392 14689 14426
rect 14655 14324 14689 14358
rect 14655 14256 14689 14290
rect 14655 14188 14689 14222
rect 14655 14120 14689 14154
rect 14655 14052 14689 14086
rect 14655 13984 14689 14018
rect 14655 13916 14689 13950
rect 14655 13848 14689 13882
rect 14655 13780 14689 13814
rect 14655 13712 14689 13746
rect 14655 13644 14689 13678
rect 14655 13576 14689 13610
rect 14655 13508 14689 13542
rect 13176 13374 13210 13408
rect 13176 13306 13210 13340
rect 13176 13238 13210 13272
rect 14655 13440 14689 13474
rect 14655 13372 14689 13406
rect 14655 13304 14689 13338
rect 13176 13170 13210 13204
rect 13176 13102 13210 13136
rect 13176 13034 13210 13068
rect 13176 12966 13210 13000
rect 13176 12898 13210 12932
rect 13176 12830 13210 12864
rect 13176 12762 13210 12796
rect 13176 12694 13210 12728
rect 13176 12626 13210 12660
rect 13176 12558 13210 12592
rect 13176 12490 13210 12524
rect 13176 12422 13210 12456
rect 13176 12354 13210 12388
rect 13176 12286 13210 12320
rect 13176 12218 13210 12252
rect 14655 13236 14689 13270
rect 14655 13168 14689 13202
rect 14655 13100 14689 13134
rect 14655 13032 14689 13066
rect 14655 12964 14689 12998
rect 14655 12896 14689 12930
rect 14655 12828 14689 12862
rect 14655 12760 14689 12794
rect 14655 12692 14689 12726
rect 14655 12624 14689 12658
rect 14655 12556 14689 12590
rect 14655 12488 14689 12522
rect 14655 12420 14689 12454
rect 14655 12352 14689 12386
rect 14655 12284 14689 12318
rect 14655 12216 14689 12250
rect 13176 12150 13210 12184
rect 13176 12082 13210 12116
rect 14655 12148 14689 12182
rect 13248 12014 13282 12048
rect 13316 12014 13350 12048
rect 13384 12014 13418 12048
rect 13452 12014 13486 12048
rect 13520 12014 13554 12048
rect 13588 12014 13622 12048
rect 13656 12014 13690 12048
rect 13724 12014 13758 12048
rect 13792 12014 13826 12048
rect 13860 12014 13894 12048
rect 13928 12014 13962 12048
rect 13996 12014 14030 12048
rect 14064 12014 14098 12048
rect 14132 12014 14166 12048
rect 14200 12014 14234 12048
rect 14268 12014 14302 12048
rect 14336 12014 14370 12048
rect 14404 12014 14438 12048
rect 14472 12014 14506 12048
rect 14587 12014 14621 12048
rect 4796 7429 4830 7463
rect 4796 7361 4830 7395
rect 5656 7429 5690 7463
rect 4796 7293 4830 7327
rect 4796 7225 4830 7259
rect 4796 7157 4830 7191
rect 4796 7089 4830 7123
rect 4796 7021 4830 7055
rect 4796 6953 4830 6987
rect 4796 6885 4830 6919
rect 5656 7361 5690 7395
rect 6666 7429 6700 7463
rect 5656 7293 5690 7327
rect 5656 7225 5690 7259
rect 5656 7157 5690 7191
rect 5656 7089 5690 7123
rect 5656 7021 5690 7055
rect 5656 6953 5690 6987
rect 5656 6885 5690 6919
rect 4796 6817 4830 6851
rect 4796 6749 4830 6783
rect 4796 6681 4830 6715
rect 4796 6613 4830 6647
rect 6666 7361 6700 7395
rect 7669 7429 7703 7463
rect 6666 7293 6700 7327
rect 6666 7225 6700 7259
rect 6666 7157 6700 7191
rect 6666 7089 6700 7123
rect 6666 7021 6700 7055
rect 6666 6953 6700 6987
rect 6666 6885 6700 6919
rect 5656 6817 5690 6851
rect 5656 6749 5690 6783
rect 5656 6681 5690 6715
rect 5656 6613 5690 6647
rect 7669 7361 7703 7395
rect 7669 7293 7703 7327
rect 7669 7225 7703 7259
rect 7669 7157 7703 7191
rect 7669 7089 7703 7123
rect 7669 7021 7703 7055
rect 7669 6953 7703 6987
rect 7669 6885 7703 6919
rect 6666 6817 6700 6851
rect 6666 6749 6700 6783
rect 6666 6681 6700 6715
rect 6666 6613 6700 6647
rect 7669 6817 7703 6851
rect 7669 6749 7703 6783
rect 7669 6681 7703 6715
rect 7669 6613 7703 6647
rect 3997 6545 3998 6579
rect 4032 6545 4066 6579
rect 4100 6545 4134 6579
rect 4168 6545 4202 6579
rect 4236 6545 4270 6579
rect 4304 6545 4338 6579
rect 4372 6545 4406 6579
rect 4440 6545 4474 6579
rect 4508 6545 4542 6579
rect 4576 6545 4610 6579
rect 4644 6545 4678 6579
rect 4712 6545 4746 6579
rect 4780 6545 4814 6579
rect 4848 6545 4882 6579
rect 4916 6545 4950 6579
rect 4984 6545 5018 6579
rect 5052 6545 5086 6579
rect 5120 6545 5154 6579
rect 5188 6545 5222 6579
rect 5256 6545 5290 6579
rect 5324 6545 5358 6579
rect 5392 6545 5426 6579
rect 5460 6545 5494 6579
rect 5528 6545 5562 6579
rect 5596 6545 5630 6579
rect 5664 6545 5698 6579
rect 5732 6545 5766 6579
rect 5800 6545 5834 6579
rect 5868 6545 5902 6579
rect 5936 6545 5970 6579
rect 6004 6545 6038 6579
rect 6072 6545 6106 6579
rect 6140 6545 6174 6579
rect 6208 6545 6242 6579
rect 6276 6545 6310 6579
rect 6344 6545 6378 6579
rect 6412 6545 6446 6579
rect 6480 6545 6514 6579
rect 6548 6545 6582 6579
rect 6616 6545 6650 6579
rect 6684 6545 6718 6579
rect 6752 6545 6786 6579
rect 6820 6545 6854 6579
rect 6888 6545 6922 6579
rect 6956 6545 6990 6579
rect 7024 6545 7058 6579
rect 7092 6545 7126 6579
rect 7160 6545 7194 6579
rect 7228 6545 7262 6579
rect 7296 6545 7330 6579
rect 7364 6545 7398 6579
rect 7432 6545 7466 6579
rect 7500 6545 7534 6579
rect 7568 6545 7602 6579
rect 7636 6545 7670 6579
rect 7704 6545 7738 6579
rect 7772 6545 7806 6579
rect 7840 6545 7874 6579
rect 7908 6545 7942 6579
rect 7976 6545 8010 6579
rect 8044 6545 8078 6579
rect 8112 6545 8146 6579
rect 8180 6545 8214 6579
rect 8248 6545 8282 6579
rect 8316 6545 8350 6579
rect 8384 6545 8418 6579
rect 8452 6545 8486 6579
rect 8520 6545 8554 6579
rect 8588 6545 8622 6579
rect 8656 6545 8690 6579
rect 8724 6545 8758 6579
rect 8792 6545 8826 6579
rect 8860 6545 8894 6579
rect 8928 6545 8962 6579
rect 8996 6545 9030 6579
rect 9064 6545 9098 6579
rect 9132 6545 9166 6579
rect 9200 6545 9234 6579
rect 9268 6545 9302 6579
rect 9336 6545 9370 6579
rect 9404 6545 9438 6579
rect 9472 6545 9506 6579
rect 9540 6545 9574 6579
rect 9608 6545 9642 6579
rect 9676 6545 9710 6579
rect 9744 6545 9778 6579
rect 9812 6545 9846 6579
rect 9880 6545 9914 6579
rect 9948 6545 9982 6579
rect 10016 6545 10050 6579
rect 10084 6545 10118 6579
rect 10152 6545 10186 6579
rect 10220 6545 10254 6579
rect 10288 6545 10322 6579
rect 10356 6545 10390 6579
rect 10424 6545 10458 6579
rect 10492 6545 10526 6579
rect 10560 6545 10594 6579
rect 10628 6545 10662 6579
rect 10696 6545 10730 6579
rect 10764 6545 10798 6579
rect 10832 6545 10866 6579
rect 10900 6545 10934 6579
rect 10968 6545 11002 6579
rect 11036 6545 11070 6579
rect 11104 6545 11138 6579
rect 11172 6545 11206 6579
rect 11240 6545 11274 6579
rect 11308 6545 11342 6579
rect 11376 6545 11410 6579
rect 11444 6545 11478 6579
rect 11512 6545 11546 6579
rect 11580 6545 11614 6579
rect 11648 6545 11682 6579
rect 11716 6545 11750 6579
rect 11784 6545 11818 6579
rect 11852 6545 11886 6579
rect 11920 6545 11954 6579
<< mvnsubdiffcont >>
rect 7857 8185 7891 8219
rect 7925 8185 7959 8219
rect 7993 8185 8027 8219
rect 8061 8185 8095 8219
rect 8129 8185 8163 8219
rect 8197 8185 8231 8219
rect 8265 8185 8299 8219
rect 8333 8185 8367 8219
rect 8401 8185 8435 8219
rect 8469 8185 8503 8219
rect 8537 8185 8571 8219
rect 8605 8185 8639 8219
rect 8673 8185 8707 8219
rect 8741 8185 8775 8219
rect 8809 8185 8843 8219
rect 8877 8185 8911 8219
rect 8945 8185 8979 8219
rect 9013 8185 9047 8219
rect 9081 8185 9115 8219
rect 9149 8185 9183 8219
rect 9217 8185 9251 8219
rect 9285 8185 9319 8219
rect 9353 8185 9387 8219
rect 9421 8185 9455 8219
rect 9489 8185 9523 8219
rect 9557 8185 9591 8219
rect 9625 8185 9659 8219
rect 9693 8185 9727 8219
rect 9761 8185 9795 8219
rect 9829 8185 9863 8219
rect 9897 8185 9931 8219
rect 9965 8185 9999 8219
rect 10033 8185 10067 8219
rect 10101 8185 10135 8219
rect 10169 8185 10203 8219
rect 10237 8185 10271 8219
rect 10305 8185 10339 8219
rect 10373 8185 10407 8219
rect 10441 8185 10475 8219
rect 10509 8185 10543 8219
rect 10577 8185 10611 8219
rect 10645 8185 10679 8219
rect 10713 8185 10747 8219
rect 10781 8185 10815 8219
rect 10849 8185 10883 8219
rect 10917 8185 10951 8219
rect 10985 8185 11019 8219
rect 11053 8185 11087 8219
rect 11121 8185 11155 8219
rect 11189 8185 11223 8219
rect 11257 8185 11291 8219
rect 11325 8185 11359 8219
rect 11393 8185 11427 8219
rect 11461 8185 11495 8219
rect 11529 8185 11563 8219
rect 11597 8185 11631 8219
rect 11665 8185 11699 8219
rect 11733 8185 11767 8219
rect 11801 8185 11835 8219
rect 11869 8185 11903 8219
rect 11937 8185 11971 8219
rect 12005 8185 12039 8219
rect 12073 8185 12107 8219
rect 12141 8185 12175 8219
rect 12209 8185 12243 8219
rect 12277 8185 12311 8219
rect 12345 8185 12379 8219
rect 12413 8185 12447 8219
rect 12481 8185 12515 8219
rect 12549 8185 12583 8219
rect 12617 8185 12651 8219
rect 12685 8185 12719 8219
rect 12753 8185 12787 8219
rect 12821 8185 12855 8219
rect 7824 8117 7858 8151
rect 7824 8049 7858 8083
rect 12896 8152 12930 8186
rect 12896 8084 12930 8118
rect 7824 7981 7858 8015
rect 12896 8016 12930 8050
rect 7824 7913 7858 7947
rect 7824 7845 7858 7879
rect 12896 7948 12930 7982
rect 12896 7880 12930 7914
rect 7824 7777 7858 7811
rect 7824 7709 7858 7743
rect 7824 7641 7858 7675
rect 12896 7812 12930 7846
rect 12896 7744 12930 7778
rect 12896 7676 12930 7710
rect 3928 7540 3962 7574
rect 3996 7540 4030 7574
rect 4064 7540 4098 7574
rect 4132 7540 4166 7574
rect 4200 7540 4234 7574
rect 4268 7540 4302 7574
rect 4336 7540 4370 7574
rect 4404 7540 4438 7574
rect 4472 7540 4506 7574
rect 4540 7540 4574 7574
rect 4608 7540 4642 7574
rect 4676 7540 4710 7574
rect 4744 7540 4778 7574
rect 4812 7540 4846 7574
rect 4880 7540 4914 7574
rect 4948 7540 4982 7574
rect 5016 7540 5050 7574
rect 5084 7540 5118 7574
rect 5152 7540 5186 7574
rect 5220 7540 5254 7574
rect 5288 7540 5322 7574
rect 5356 7540 5390 7574
rect 5424 7540 5458 7574
rect 5492 7540 5526 7574
rect 5560 7540 5594 7574
rect 5628 7540 5662 7574
rect 5696 7540 5730 7574
rect 5764 7540 5798 7574
rect 5832 7540 5866 7574
rect 5900 7540 5934 7574
rect 5968 7540 6002 7574
rect 6036 7540 6070 7574
rect 6104 7540 6138 7574
rect 6172 7540 6206 7574
rect 6240 7540 6274 7574
rect 6308 7540 6342 7574
rect 6376 7540 6410 7574
rect 6444 7540 6478 7574
rect 6512 7540 6546 7574
rect 6580 7540 6614 7574
rect 6648 7540 6682 7574
rect 6716 7540 6750 7574
rect 6784 7540 6818 7574
rect 6852 7540 6886 7574
rect 6920 7540 6954 7574
rect 6988 7540 7022 7574
rect 7056 7540 7090 7574
rect 7124 7540 7158 7574
rect 7192 7540 7226 7574
rect 7260 7540 7294 7574
rect 7328 7540 7362 7574
rect 7396 7540 7430 7574
rect 7464 7540 7498 7574
rect 7532 7540 7566 7574
rect 7600 7540 7634 7574
rect 7668 7540 7702 7574
rect 7736 7540 7770 7574
rect 7824 7573 7858 7607
rect 3895 7461 3929 7495
rect 3895 7393 3929 7427
rect 3895 7325 3929 7359
rect 3895 7257 3929 7291
rect 3895 7189 3929 7223
rect 3895 7121 3929 7155
rect 3895 7053 3929 7087
rect 3895 6985 3929 7019
rect 3895 6917 3929 6951
rect 3895 6849 3929 6883
rect 3895 6781 3929 6815
rect 3895 6713 3929 6747
rect 3895 6645 3929 6679
rect 3895 6577 3929 6611
rect 12896 7608 12930 7642
rect 12896 7540 12930 7574
rect 12896 7472 12930 7506
rect 12896 7404 12930 7438
rect 12896 7336 12930 7370
rect 12896 7268 12930 7302
rect 12896 7200 12930 7234
rect 12896 7132 12930 7166
rect 12896 7064 12930 7098
rect 12896 6996 12930 7030
rect 12896 6928 12930 6962
rect 12896 6860 12930 6894
rect 12896 6792 12930 6826
rect 12896 6724 12930 6758
rect 12896 6656 12930 6690
rect 12896 6588 12930 6622
rect 3964 6545 3997 6579
rect 3895 6509 3929 6543
rect 3895 6441 3929 6475
rect 3895 6373 3929 6407
rect 12896 6520 12930 6554
rect 12896 6452 12930 6486
rect 3895 6305 3929 6339
rect 3895 6237 3929 6271
rect 3895 6169 3929 6203
rect 3895 6101 3929 6135
rect 3895 6033 3929 6067
rect 3895 5965 3929 5999
rect 3895 5897 3929 5931
rect 3895 5829 3929 5863
rect 3895 5761 3929 5795
rect 3895 5693 3929 5727
rect 12195 6286 12229 6320
rect 12319 6319 12353 6353
rect 12387 6319 12421 6353
rect 12455 6319 12489 6353
rect 12523 6319 12557 6353
rect 12591 6319 12625 6353
rect 12659 6319 12693 6353
rect 12727 6319 12761 6353
rect 12795 6319 12829 6353
rect 12863 6319 12897 6353
rect 12195 6218 12229 6252
rect 12195 6150 12229 6184
rect 12195 6082 12229 6116
rect 12195 6014 12229 6048
rect 12195 5946 12229 5980
rect 12195 5878 12229 5912
rect 12195 5810 12229 5844
rect 12195 5742 12229 5776
rect 3895 5625 3929 5659
rect 3895 5557 3929 5591
rect 3895 5489 3929 5523
rect 3895 5421 3929 5455
rect 3895 5353 3929 5387
rect 3895 5285 3929 5319
rect 3895 5217 3929 5251
rect 3895 5149 3929 5183
rect 3895 5081 3929 5115
rect 3895 5013 3929 5047
rect 3895 4945 3929 4979
rect 3895 4877 3929 4911
rect 3895 4809 3929 4843
rect 3895 4741 3929 4775
rect 3895 4673 3929 4707
rect 3895 4605 3929 4639
rect 3895 4537 3929 4571
rect 3895 4469 3929 4503
rect 3895 4401 3929 4435
rect 3895 4333 3929 4367
rect 3895 4265 3929 4299
rect 3895 4197 3929 4231
rect 3895 4129 3929 4163
rect 3895 4061 3929 4095
rect 3895 3993 3929 4027
rect 3895 3925 3929 3959
rect 3895 3857 3929 3891
rect 3895 3789 3929 3823
rect 3895 3721 3929 3755
rect 3895 3653 3929 3687
rect 3895 3585 3929 3619
rect 3895 3517 3929 3551
rect 3895 3449 3929 3483
rect 3895 3381 3929 3415
rect 3895 3313 3929 3347
rect 3895 3245 3929 3279
rect 3895 3177 3929 3211
rect 3895 3109 3929 3143
rect 3895 3041 3929 3075
rect 3895 2973 3929 3007
rect 3895 2905 3929 2939
rect 3895 2837 3929 2871
rect 3895 2769 3929 2803
rect 3895 2701 3929 2735
rect 3895 2633 3929 2667
rect 3895 2565 3929 2599
rect 3895 2497 3929 2531
rect 3895 2429 3929 2463
rect 3895 2361 3929 2395
rect 3895 2293 3929 2327
rect 3895 2225 3929 2259
rect 3895 2157 3929 2191
rect 3895 2089 3929 2123
rect 3895 2021 3929 2055
rect 3895 1953 3929 1987
rect 12195 5674 12229 5708
rect 12195 5606 12229 5640
rect 12195 5538 12229 5572
rect 12195 5470 12229 5504
rect 12195 5402 12229 5436
rect 12195 5334 12229 5368
rect 12195 5266 12229 5300
rect 12195 5198 12229 5232
rect 12195 5130 12229 5164
rect 12195 5062 12229 5096
rect 12195 4994 12229 5028
rect 12195 4926 12229 4960
rect 12195 4858 12229 4892
rect 12195 4790 12229 4824
rect 12195 4722 12229 4756
rect 12195 4654 12229 4688
rect 12195 4586 12229 4620
rect 12195 4518 12229 4552
rect 12195 4450 12229 4484
rect 12195 4382 12229 4416
rect 12195 4314 12229 4348
rect 12195 4246 12229 4280
rect 12195 4178 12229 4212
rect 12195 4110 12229 4144
rect 12195 4042 12229 4076
rect 12195 3974 12229 4008
rect 12195 3906 12229 3940
rect 12195 3838 12229 3872
rect 12195 3770 12229 3804
rect 12195 3702 12229 3736
rect 12195 3634 12229 3668
rect 12195 3566 12229 3600
rect 12195 3498 12229 3532
rect 12195 3430 12229 3464
rect 12195 3362 12229 3396
rect 12195 3294 12229 3328
rect 12195 3226 12229 3260
rect 12195 3158 12229 3192
rect 12195 3090 12229 3124
rect 12195 3022 12229 3056
rect 12195 2954 12229 2988
rect 12195 2886 12229 2920
rect 12195 2818 12229 2852
rect 12195 2750 12229 2784
rect 12195 2682 12229 2716
rect 12195 2614 12229 2648
rect 12195 2546 12229 2580
rect 12195 2478 12229 2512
rect 12195 2410 12229 2444
rect 12195 2342 12229 2376
rect 12195 2274 12229 2308
rect 12195 2206 12229 2240
rect 12195 2138 12229 2172
rect 12195 2070 12229 2104
rect 12195 2002 12229 2036
rect 3895 1885 3929 1919
rect 3895 1817 3929 1851
rect 3895 1749 3929 1783
rect 3895 1681 3929 1715
rect 3895 1613 3929 1647
rect 3895 1545 3929 1579
rect 3895 1477 3929 1511
rect 3895 1409 3929 1443
rect 3895 1341 3929 1375
rect 3895 1273 3929 1307
rect 3895 1205 3929 1239
rect 3895 1137 3929 1171
rect 3895 1069 3929 1103
rect 3895 1001 3929 1035
rect 3895 933 3929 967
rect 3895 865 3929 899
rect 12195 1934 12229 1968
rect 12195 1866 12229 1900
rect 12195 1798 12229 1832
rect 12195 1730 12229 1764
rect 12195 1662 12229 1696
rect 12195 1594 12229 1628
rect 12195 1526 12229 1560
rect 12195 1458 12229 1492
rect 12195 1390 12229 1424
rect 12195 1322 12229 1356
rect 12195 1254 12229 1288
rect 12195 1186 12229 1220
rect 12195 1017 12229 1051
rect 12195 949 12229 983
rect 4002 832 4036 866
rect 4070 832 4104 866
rect 4138 832 4172 866
rect 4206 832 4240 866
rect 4274 832 4308 866
rect 4342 832 4376 866
rect 4410 832 4444 866
rect 4478 832 4512 866
rect 4546 832 4580 866
rect 4614 832 4648 866
rect 4682 832 4716 866
rect 4750 832 4784 866
rect 4818 832 4852 866
rect 4886 832 4920 866
rect 4954 832 4988 866
rect 5022 832 5056 866
rect 5090 832 5124 866
rect 5158 832 5192 866
rect 5226 832 5260 866
rect 5294 832 5328 866
rect 5362 832 5396 866
rect 5430 832 5464 866
rect 5498 832 5532 866
rect 5566 832 5600 866
rect 5634 832 5668 866
rect 5702 832 5736 866
rect 5770 832 5804 866
rect 5838 832 5872 866
rect 5906 832 5940 866
rect 5974 832 6008 866
rect 6042 832 6076 866
rect 6110 832 6144 866
rect 6178 832 6212 866
rect 6246 832 6280 866
rect 6314 832 6348 866
rect 6382 832 6416 866
rect 6450 832 6484 866
rect 6518 832 6552 866
rect 6586 832 6620 866
rect 6654 832 6688 866
rect 6722 832 6756 866
rect 6790 832 6824 866
rect 6858 832 6892 866
rect 6926 832 6960 866
rect 6994 832 7028 866
rect 7062 832 7096 866
rect 7130 832 7164 866
rect 7198 832 7232 866
rect 7266 832 7300 866
rect 7334 832 7368 866
rect 7402 832 7436 866
rect 7470 832 7504 866
rect 7538 832 7572 866
rect 7606 832 7640 866
rect 7674 832 7708 866
rect 7742 832 7776 866
rect 7810 832 7844 866
rect 7878 832 7912 866
rect 7946 832 7980 866
rect 8014 832 8048 866
rect 8082 832 8116 866
rect 8150 832 8184 866
rect 8218 832 8252 866
rect 8286 832 8320 866
rect 8354 832 8388 866
rect 8422 832 8456 866
rect 8490 832 8524 866
rect 8558 832 8592 866
rect 8626 832 8660 866
rect 8694 832 8728 866
rect 8762 832 8796 866
rect 8830 832 8864 866
rect 8898 832 8932 866
rect 8966 832 9000 866
rect 9034 832 9068 866
rect 9102 832 9136 866
rect 9170 832 9204 866
rect 9238 832 9272 866
rect 9306 832 9340 866
rect 9374 832 9408 866
rect 9442 832 9476 866
rect 9510 832 9544 866
rect 9578 832 9612 866
rect 9646 832 9680 866
rect 9714 832 9748 866
rect 9782 832 9816 866
rect 9850 832 9884 866
rect 9918 832 9952 866
rect 9986 832 10020 866
rect 10054 832 10088 866
rect 10122 832 10156 866
rect 10190 832 10224 866
rect 10258 832 10292 866
rect 10326 832 10360 866
rect 10394 832 10428 866
rect 10462 832 10496 866
rect 10530 832 10564 866
rect 10598 832 10632 866
rect 10666 832 10700 866
rect 10734 832 10768 866
rect 10802 832 10836 866
rect 10870 832 10904 866
rect 10938 832 10972 866
rect 11006 832 11040 866
rect 11074 832 11108 866
rect 11142 832 11176 866
rect 11210 832 11244 866
rect 11278 832 11312 866
rect 11346 832 11380 866
rect 11414 832 11448 866
rect 11482 832 11516 866
rect 11550 832 11584 866
rect 11618 832 11652 866
rect 11686 832 11720 866
rect 11754 832 11788 866
rect 11822 832 11856 866
rect 11890 832 11924 866
rect 11958 832 11992 866
rect 12026 832 12060 866
rect 12094 832 12128 866
rect 12162 832 12196 866
<< poly >>
rect 3265 14532 3445 14554
rect 3265 14498 3302 14532
rect 3336 14498 3370 14532
rect 3404 14498 3445 14532
rect 3265 14476 3445 14498
rect 3501 14532 3681 14554
rect 3501 14498 3538 14532
rect 3572 14498 3606 14532
rect 3640 14498 3681 14532
rect 3501 14476 3681 14498
rect 3737 14532 3917 14554
rect 3737 14498 3774 14532
rect 3808 14498 3842 14532
rect 3876 14498 3917 14532
rect 3737 14476 3917 14498
rect 3973 14532 4153 14554
rect 3973 14498 4010 14532
rect 4044 14498 4078 14532
rect 4112 14498 4153 14532
rect 3973 14476 4153 14498
rect -464 13602 -264 13618
rect -464 13568 -448 13602
rect -414 13568 -314 13602
rect -280 13568 -264 13602
rect -464 13552 -264 13568
rect -208 13602 1784 13618
rect -208 13568 -192 13602
rect -158 13568 -123 13602
rect -89 13568 -54 13602
rect -20 13568 15 13602
rect 49 13568 84 13602
rect 118 13568 153 13602
rect 187 13568 222 13602
rect 256 13568 291 13602
rect 325 13568 360 13602
rect 394 13568 429 13602
rect 463 13568 498 13602
rect 532 13568 567 13602
rect 601 13568 636 13602
rect 670 13568 705 13602
rect 739 13568 774 13602
rect 808 13568 843 13602
rect 877 13568 912 13602
rect 946 13568 981 13602
rect 1015 13568 1050 13602
rect 1084 13568 1119 13602
rect 1153 13568 1188 13602
rect 1222 13568 1257 13602
rect 1291 13568 1326 13602
rect 1360 13568 1394 13602
rect 1428 13568 1462 13602
rect 1496 13568 1530 13602
rect 1564 13568 1598 13602
rect 1632 13568 1666 13602
rect 1700 13568 1734 13602
rect 1768 13568 1784 13602
rect -208 13552 1784 13568
rect 1840 13602 2040 13618
rect 1840 13568 1856 13602
rect 1890 13568 1990 13602
rect 2024 13568 2040 13602
rect 1840 13552 2040 13568
rect 13769 14583 13969 14605
rect 13769 14549 13818 14583
rect 13852 14549 13886 14583
rect 13920 14549 13969 14583
rect 13769 14527 13969 14549
rect 14025 14583 14225 14605
rect 14025 14549 14074 14583
rect 14108 14549 14142 14583
rect 14176 14549 14225 14583
rect 14025 14527 14225 14549
rect 4454 12965 4654 12987
rect 4454 12931 4503 12965
rect 4537 12931 4571 12965
rect 4605 12931 4654 12965
rect 4454 12909 4654 12931
rect 4710 12965 4910 12987
rect 4710 12931 4759 12965
rect 4793 12931 4827 12965
rect 4861 12931 4910 12965
rect 4710 12909 4910 12931
rect 3265 12390 3445 12412
rect 3265 12356 3302 12390
rect 3336 12356 3370 12390
rect 3404 12356 3445 12390
rect 3265 12334 3445 12356
rect 3501 12390 3681 12412
rect 3501 12356 3538 12390
rect 3572 12356 3606 12390
rect 3640 12356 3681 12390
rect 3501 12334 3681 12356
rect 3737 12390 3917 12412
rect 3737 12356 3774 12390
rect 3808 12356 3842 12390
rect 3876 12356 3917 12390
rect 3737 12334 3917 12356
rect 3973 12390 4153 12412
rect 3973 12356 4010 12390
rect 4044 12356 4078 12390
rect 4112 12356 4153 12390
rect 3973 12334 4153 12356
rect -376 12042 -176 12148
rect -376 12008 -327 12042
rect -293 12008 -259 12042
rect -225 12008 -176 12042
rect -376 11988 -176 12008
rect -120 12042 80 12149
rect 254 12058 354 12147
rect -120 12008 -71 12042
rect -37 12008 -3 12042
rect 31 12008 80 12042
rect -120 11988 80 12008
rect 235 12042 369 12058
rect 235 12008 251 12042
rect 285 12008 319 12042
rect 353 12008 369 12042
rect 235 11992 369 12008
rect 4421 12015 4621 12056
rect 4421 11981 4464 12015
rect 4498 11981 4532 12015
rect 4566 11981 4621 12015
rect 4421 11959 4621 11981
rect 4677 12015 4877 12052
rect 4677 11981 4720 12015
rect 4754 11981 4788 12015
rect 4822 11981 4877 12015
rect 4677 11959 4877 11981
rect 12015 12195 12215 12217
rect 12015 12161 12064 12195
rect 12098 12161 12132 12195
rect 12166 12161 12215 12195
rect 12015 12139 12215 12161
rect 12271 12195 12471 12217
rect 12271 12161 12320 12195
rect 12354 12161 12388 12195
rect 12422 12161 12471 12195
rect 12271 12139 12471 12161
rect 13513 13369 13713 13463
rect 13513 13335 13558 13369
rect 13592 13335 13626 13369
rect 13660 13335 13713 13369
rect 13513 13254 13713 13335
rect 13769 13369 13969 13463
rect 13769 13335 13814 13369
rect 13848 13335 13882 13369
rect 13916 13335 13969 13369
rect 13769 13254 13969 13335
rect 14025 13369 14225 13463
rect 14025 13335 14070 13369
rect 14104 13335 14138 13369
rect 14172 13335 14225 13369
rect 14025 13254 14225 13335
rect 14281 13369 14481 13463
rect 14281 13335 14326 13369
rect 14360 13335 14394 13369
rect 14428 13335 14481 13369
rect 14281 13254 14481 13335
rect 13769 12168 13969 12190
rect 13769 12134 13818 12168
rect 13852 12134 13886 12168
rect 13920 12134 13969 12168
rect 13769 12112 13969 12134
rect 14025 12168 14225 12190
rect 14025 12134 14074 12168
rect 14108 12134 14142 12168
rect 14176 12134 14225 12168
rect 14025 12112 14225 12134
rect 8084 7804 8161 7845
rect 8084 7770 8105 7804
rect 8139 7770 8161 7804
rect 8084 7736 8161 7770
rect 8084 7702 8105 7736
rect 8139 7702 8161 7736
rect 8084 7665 8161 7702
rect 10225 7804 10303 7845
rect 10225 7770 10247 7804
rect 10281 7770 10303 7804
rect 10225 7736 10303 7770
rect 10225 7702 10247 7736
rect 10281 7702 10303 7736
rect 10225 7665 10303 7702
rect 10401 7804 10479 7845
rect 10401 7770 10423 7804
rect 10457 7770 10479 7804
rect 10401 7736 10479 7770
rect 10401 7702 10423 7736
rect 10457 7702 10479 7736
rect 10401 7665 10479 7702
rect 12543 7804 12621 7845
rect 12543 7770 12565 7804
rect 12599 7770 12621 7804
rect 12543 7736 12621 7770
rect 12543 7702 12565 7736
rect 12599 7702 12621 7736
rect 12543 7665 12621 7702
rect 8084 7568 8161 7609
rect 4460 7177 4538 7221
rect 4460 7143 4482 7177
rect 4516 7143 4538 7177
rect 4460 7109 4538 7143
rect 4460 7075 4482 7109
rect 4516 7075 4538 7109
rect 4460 7041 4538 7075
rect 5343 7177 5421 7221
rect 5343 7143 5365 7177
rect 5399 7143 5421 7177
rect 5343 7109 5421 7143
rect 5343 7075 5365 7109
rect 5399 7075 5421 7109
rect 5343 7041 5421 7075
rect 6201 7177 6279 7221
rect 6201 7143 6223 7177
rect 6257 7143 6279 7177
rect 6201 7109 6279 7143
rect 6201 7075 6223 7109
rect 6257 7075 6279 7109
rect 6201 7041 6279 7075
rect 8084 7534 8105 7568
rect 8139 7534 8161 7568
rect 8084 7500 8161 7534
rect 8084 7466 8105 7500
rect 8139 7466 8161 7500
rect 8084 7429 8161 7466
rect 10225 7568 10303 7609
rect 10225 7534 10247 7568
rect 10281 7534 10303 7568
rect 10225 7500 10303 7534
rect 10225 7466 10247 7500
rect 10281 7466 10303 7500
rect 10225 7429 10303 7466
rect 10401 7568 10479 7609
rect 10401 7534 10423 7568
rect 10457 7534 10479 7568
rect 10401 7500 10479 7534
rect 10401 7466 10423 7500
rect 10457 7466 10479 7500
rect 10401 7429 10479 7466
rect 12543 7568 12621 7609
rect 12543 7534 12565 7568
rect 12599 7534 12621 7568
rect 12543 7500 12621 7534
rect 12543 7466 12565 7500
rect 12599 7466 12621 7500
rect 12543 7429 12621 7466
rect 7337 7177 7415 7221
rect 7337 7143 7359 7177
rect 7393 7143 7415 7177
rect 7337 7109 7415 7143
rect 7337 7075 7359 7109
rect 7393 7075 7415 7109
rect 7337 7041 7415 7075
rect 8084 7332 8161 7373
rect 8084 7298 8105 7332
rect 8139 7298 8161 7332
rect 8084 7264 8161 7298
rect 8084 7230 8105 7264
rect 8139 7230 8161 7264
rect 8084 7193 8161 7230
rect 10225 7332 10303 7373
rect 10225 7298 10247 7332
rect 10281 7298 10303 7332
rect 10225 7264 10303 7298
rect 10225 7230 10247 7264
rect 10281 7230 10303 7264
rect 10225 7193 10303 7230
rect 10401 7332 10479 7373
rect 10401 7298 10423 7332
rect 10457 7298 10479 7332
rect 10401 7264 10479 7298
rect 10401 7230 10423 7264
rect 10457 7230 10479 7264
rect 10401 7193 10479 7230
rect 12543 7332 12621 7373
rect 12543 7298 12565 7332
rect 12599 7298 12621 7332
rect 12543 7264 12621 7298
rect 12543 7230 12565 7264
rect 12599 7230 12621 7264
rect 12543 7193 12621 7230
rect 8084 7096 8161 7137
rect 8084 7062 8105 7096
rect 8139 7062 8161 7096
rect 8084 7028 8161 7062
rect 8084 6994 8105 7028
rect 8139 6994 8161 7028
rect 8084 6957 8161 6994
rect 10225 7096 10303 7137
rect 10225 7062 10247 7096
rect 10281 7062 10303 7096
rect 10225 7028 10303 7062
rect 10225 6994 10247 7028
rect 10281 6994 10303 7028
rect 10225 6957 10303 6994
rect 10401 7096 10479 7137
rect 10401 7062 10423 7096
rect 10457 7062 10479 7096
rect 10401 7028 10479 7062
rect 10401 6994 10423 7028
rect 10457 6994 10479 7028
rect 10401 6957 10479 6994
rect 12543 7096 12621 7137
rect 12543 7062 12565 7096
rect 12599 7062 12621 7096
rect 12543 7028 12621 7062
rect 12543 6994 12565 7028
rect 12599 6994 12621 7028
rect 12543 6957 12621 6994
rect 11817 5166 11889 5275
rect 11817 5132 11839 5166
rect 11873 5132 11889 5166
rect 11817 5098 11889 5132
rect 11817 5064 11839 5098
rect 11873 5064 11889 5098
rect 11817 5030 11889 5064
rect 11817 4996 11839 5030
rect 11873 4996 11889 5030
rect 11817 4962 11889 4996
rect 11817 4928 11839 4962
rect 11873 4928 11889 4962
rect 11817 4819 11889 4928
rect 11817 3178 11889 3227
rect 11817 3144 11839 3178
rect 11873 3144 11889 3178
rect 11817 3110 11889 3144
rect 11817 3076 11839 3110
rect 11873 3076 11889 3110
rect 11817 3027 11889 3076
rect 11817 2922 11889 2971
rect 11817 2888 11839 2922
rect 11873 2888 11889 2922
rect 11817 2854 11889 2888
rect 11817 2820 11839 2854
rect 11873 2820 11889 2854
rect 11817 2771 11889 2820
<< polycont >>
rect 3302 14498 3336 14532
rect 3370 14498 3404 14532
rect 3538 14498 3572 14532
rect 3606 14498 3640 14532
rect 3774 14498 3808 14532
rect 3842 14498 3876 14532
rect 4010 14498 4044 14532
rect 4078 14498 4112 14532
rect -448 13568 -414 13602
rect -314 13568 -280 13602
rect -192 13568 -158 13602
rect -123 13568 -89 13602
rect -54 13568 -20 13602
rect 15 13568 49 13602
rect 84 13568 118 13602
rect 153 13568 187 13602
rect 222 13568 256 13602
rect 291 13568 325 13602
rect 360 13568 394 13602
rect 429 13568 463 13602
rect 498 13568 532 13602
rect 567 13568 601 13602
rect 636 13568 670 13602
rect 705 13568 739 13602
rect 774 13568 808 13602
rect 843 13568 877 13602
rect 912 13568 946 13602
rect 981 13568 1015 13602
rect 1050 13568 1084 13602
rect 1119 13568 1153 13602
rect 1188 13568 1222 13602
rect 1257 13568 1291 13602
rect 1326 13568 1360 13602
rect 1394 13568 1428 13602
rect 1462 13568 1496 13602
rect 1530 13568 1564 13602
rect 1598 13568 1632 13602
rect 1666 13568 1700 13602
rect 1734 13568 1768 13602
rect 1856 13568 1890 13602
rect 1990 13568 2024 13602
rect 13818 14549 13852 14583
rect 13886 14549 13920 14583
rect 14074 14549 14108 14583
rect 14142 14549 14176 14583
rect 4503 12931 4537 12965
rect 4571 12931 4605 12965
rect 4759 12931 4793 12965
rect 4827 12931 4861 12965
rect 3302 12356 3336 12390
rect 3370 12356 3404 12390
rect 3538 12356 3572 12390
rect 3606 12356 3640 12390
rect 3774 12356 3808 12390
rect 3842 12356 3876 12390
rect 4010 12356 4044 12390
rect 4078 12356 4112 12390
rect -327 12008 -293 12042
rect -259 12008 -225 12042
rect -71 12008 -37 12042
rect -3 12008 31 12042
rect 251 12008 285 12042
rect 319 12008 353 12042
rect 4464 11981 4498 12015
rect 4532 11981 4566 12015
rect 4720 11981 4754 12015
rect 4788 11981 4822 12015
rect 12064 12161 12098 12195
rect 12132 12161 12166 12195
rect 12320 12161 12354 12195
rect 12388 12161 12422 12195
rect 13558 13335 13592 13369
rect 13626 13335 13660 13369
rect 13814 13335 13848 13369
rect 13882 13335 13916 13369
rect 14070 13335 14104 13369
rect 14138 13335 14172 13369
rect 14326 13335 14360 13369
rect 14394 13335 14428 13369
rect 13818 12134 13852 12168
rect 13886 12134 13920 12168
rect 14074 12134 14108 12168
rect 14142 12134 14176 12168
rect 8105 7770 8139 7804
rect 8105 7702 8139 7736
rect 10247 7770 10281 7804
rect 10247 7702 10281 7736
rect 10423 7770 10457 7804
rect 10423 7702 10457 7736
rect 12565 7770 12599 7804
rect 12565 7702 12599 7736
rect 4482 7143 4516 7177
rect 4482 7075 4516 7109
rect 5365 7143 5399 7177
rect 5365 7075 5399 7109
rect 6223 7143 6257 7177
rect 6223 7075 6257 7109
rect 8105 7534 8139 7568
rect 8105 7466 8139 7500
rect 10247 7534 10281 7568
rect 10247 7466 10281 7500
rect 10423 7534 10457 7568
rect 10423 7466 10457 7500
rect 12565 7534 12599 7568
rect 12565 7466 12599 7500
rect 7359 7143 7393 7177
rect 7359 7075 7393 7109
rect 8105 7298 8139 7332
rect 8105 7230 8139 7264
rect 10247 7298 10281 7332
rect 10247 7230 10281 7264
rect 10423 7298 10457 7332
rect 10423 7230 10457 7264
rect 12565 7298 12599 7332
rect 12565 7230 12599 7264
rect 8105 7062 8139 7096
rect 8105 6994 8139 7028
rect 10247 7062 10281 7096
rect 10247 6994 10281 7028
rect 10423 7062 10457 7096
rect 10423 6994 10457 7028
rect 12565 7062 12599 7096
rect 12565 6994 12599 7028
rect 11839 5132 11873 5166
rect 11839 5064 11873 5098
rect 11839 4996 11873 5030
rect 11839 4928 11873 4962
rect 11839 3144 11873 3178
rect 11839 3076 11873 3110
rect 11839 2888 11873 2922
rect 11839 2820 11873 2854
<< locali >>
rect 13176 14732 13244 14766
rect 13284 14732 13312 14766
rect 13358 14732 13380 14766
rect 13432 14732 13448 14766
rect 13506 14732 13516 14766
rect 13580 14732 13584 14766
rect 13618 14732 13620 14766
rect 13686 14732 13694 14766
rect 13754 14732 13768 14766
rect 13822 14732 13842 14766
rect 13890 14732 13916 14766
rect 13958 14732 13990 14766
rect 14026 14732 14060 14766
rect 14098 14732 14128 14766
rect 14172 14732 14196 14766
rect 14246 14732 14264 14766
rect 14320 14732 14332 14766
rect 14394 14732 14400 14766
rect 14502 14732 14508 14766
rect 14570 14732 14583 14766
rect 14617 14732 14689 14766
rect 3079 14614 3147 14648
rect 3181 14614 3215 14648
rect 3249 14614 3283 14648
rect 3317 14614 3351 14648
rect 3385 14614 3419 14648
rect 3453 14614 3487 14648
rect 3521 14614 3555 14648
rect 3589 14614 3623 14648
rect 3657 14614 3691 14648
rect 3725 14614 3759 14648
rect 3793 14614 3827 14648
rect 3861 14614 3895 14648
rect 3929 14614 3963 14648
rect 3997 14614 4031 14648
rect 4065 14614 4099 14648
rect 4133 14614 4167 14648
rect 4201 14614 4235 14648
rect 4269 14614 4303 14648
rect 4337 14614 4371 14648
rect 4405 14614 4439 14648
rect 4473 14614 4507 14648
rect 4541 14614 4575 14648
rect 4609 14614 4643 14648
rect 4677 14614 4711 14648
rect 4745 14614 4779 14648
rect 4813 14614 4847 14648
rect 4881 14614 4915 14648
rect 4949 14614 4983 14648
rect 5017 14614 5121 14648
rect 3079 14558 3113 14614
rect 5087 14580 5121 14614
rect 3105 14518 3113 14524
rect 3071 14490 3113 14518
rect 3286 14498 3300 14532
rect 3336 14498 3370 14532
rect 3406 14498 3420 14532
rect 3522 14498 3538 14532
rect 3575 14498 3606 14532
rect 3647 14498 3656 14532
rect 3758 14498 3772 14532
rect 3808 14498 3842 14532
rect 3878 14498 3892 14532
rect 3994 14498 4008 14532
rect 4044 14498 4078 14532
rect 4114 14498 4128 14532
rect 5087 14512 5121 14546
rect 3071 14476 3079 14490
rect 3105 14442 3113 14456
rect 3071 14422 3113 14442
rect 3071 14400 3079 14422
rect 3105 14366 3113 14388
rect 3071 14354 3113 14366
rect 3071 14324 3079 14354
rect 3105 14290 3113 14320
rect 3071 14286 3113 14290
rect 3071 14252 3079 14286
rect 3071 14248 3113 14252
rect 3105 14218 3113 14248
rect 3071 14184 3079 14214
rect 3071 14172 3113 14184
rect -253 14083 -219 14124
rect 259 14086 293 14124
rect 771 14086 805 14124
rect 1283 14086 1317 14124
rect 1795 14086 1829 14124
rect 3105 14150 3113 14172
rect 3071 14116 3079 14138
rect 3071 14096 3113 14116
rect 3105 14082 3113 14096
rect -253 14008 -219 14049
rect 3071 14048 3079 14062
rect 3071 14020 3113 14048
rect 3105 14014 3113 14020
rect -253 13932 -219 13974
rect 515 13916 549 13954
rect 1539 13912 1573 13954
rect 1539 13836 1573 13878
rect 3 13746 37 13784
rect 1027 13746 1061 13784
rect 1539 13760 1573 13802
rect 3071 13980 3079 13986
rect 3071 13946 3113 13980
rect 3071 13944 3079 13946
rect 3105 13910 3113 13912
rect 3071 13878 3113 13910
rect 3071 13868 3079 13878
rect 3105 13834 3113 13844
rect 3071 13810 3113 13834
rect 3071 13792 3079 13810
rect 3105 13758 3113 13776
rect 3071 13742 3113 13758
rect 3071 13716 3079 13742
rect -577 13602 -475 13712
rect 2051 13602 2153 13713
rect -577 13568 -448 13602
rect -414 13568 -314 13602
rect -280 13568 -264 13602
rect -208 13568 -192 13602
rect -158 13568 -123 13602
rect -89 13600 -54 13602
rect -89 13568 -56 13600
rect -20 13568 15 13602
rect 49 13600 84 13602
rect 118 13600 153 13602
rect 187 13600 222 13602
rect 256 13600 291 13602
rect 325 13600 360 13602
rect 53 13568 84 13600
rect 128 13568 153 13600
rect 203 13568 222 13600
rect 278 13568 291 13600
rect 353 13568 360 13600
rect 394 13600 429 13602
rect -22 13566 19 13568
rect 53 13566 94 13568
rect 128 13566 169 13568
rect 203 13566 244 13568
rect 278 13566 319 13568
rect 353 13566 394 13568
rect 428 13568 429 13600
rect 463 13600 498 13602
rect 532 13600 567 13602
rect 601 13600 636 13602
rect 670 13600 705 13602
rect 739 13600 774 13602
rect 463 13568 469 13600
rect 532 13568 544 13600
rect 601 13568 619 13600
rect 670 13568 694 13600
rect 739 13568 769 13600
rect 808 13568 843 13602
rect 877 13568 912 13602
rect 946 13600 981 13602
rect 1015 13600 1050 13602
rect 1084 13600 1119 13602
rect 1153 13600 1188 13602
rect 1222 13600 1257 13602
rect 1291 13600 1326 13602
rect 951 13568 981 13600
rect 1025 13568 1050 13600
rect 1099 13568 1119 13600
rect 1173 13568 1188 13600
rect 1247 13568 1257 13600
rect 1321 13568 1326 13600
rect 1360 13600 1394 13602
rect 1360 13568 1361 13600
rect 1428 13568 1462 13602
rect 1496 13568 1530 13602
rect 1564 13568 1598 13602
rect 1632 13568 1666 13602
rect 1700 13568 1734 13602
rect 1768 13568 1784 13602
rect 1840 13568 1856 13602
rect 1890 13568 1990 13602
rect 2024 13568 2153 13602
rect 3105 13682 3113 13708
rect 3071 13674 3113 13682
rect 3071 13640 3079 13674
rect 3071 13639 3113 13640
rect 3105 13606 3113 13639
rect 3071 13572 3079 13605
rect 428 13566 469 13568
rect 503 13566 544 13568
rect 578 13566 619 13568
rect 653 13566 694 13568
rect 728 13566 769 13568
rect 803 13566 843 13568
rect 877 13566 917 13568
rect 951 13566 991 13568
rect 1025 13566 1065 13568
rect 1099 13566 1139 13568
rect 1173 13566 1213 13568
rect 1247 13566 1287 13568
rect 1321 13566 1361 13568
rect 3071 13562 3113 13572
rect 3105 13538 3113 13562
rect 3071 13504 3079 13528
rect 3071 13485 3113 13504
rect 3105 13470 3113 13485
rect -564 13376 -496 13410
rect -458 13376 -428 13410
rect -382 13376 -360 13410
rect -306 13376 -292 13410
rect -230 13376 -224 13410
rect -190 13376 -156 13410
rect -122 13376 -88 13410
rect -54 13376 -20 13410
rect 14 13376 48 13410
rect 82 13376 116 13410
rect 150 13376 184 13410
rect 218 13376 252 13410
rect 286 13376 320 13410
rect 354 13376 407 13410
rect 3079 13402 3113 13436
rect -564 13335 -530 13376
rect -564 13298 -530 13301
rect -564 13260 -530 13264
rect -564 13185 -530 13196
rect -564 13110 -530 13128
rect -564 13035 -530 13060
rect -564 12960 -530 12992
rect -564 12890 -530 12924
rect -564 12822 -530 12851
rect -564 12754 -530 12776
rect -564 12686 -530 12701
rect -564 12618 -530 12625
rect -564 12583 -530 12584
rect -564 12507 -530 12516
rect -564 12431 -530 12448
rect -564 12355 -530 12380
rect -564 12279 -530 12312
rect -564 12210 -530 12244
rect -564 12142 -530 12169
rect -564 12074 -530 12108
rect 3079 13334 3113 13368
rect 3079 13266 3113 13300
rect 3079 13198 3113 13232
rect 3079 13130 3113 13164
rect 3079 13062 3113 13096
rect 3079 12994 3113 13028
rect 5087 14444 5121 14478
rect 5087 14386 5121 14410
rect 5087 14314 5121 14342
rect 13176 14632 13210 14732
rect 13176 14564 13210 14598
rect 14655 14698 14689 14732
rect 14655 14630 14689 14632
rect 13802 14549 13816 14583
rect 13852 14549 13886 14583
rect 13922 14549 13936 14583
rect 14058 14549 14072 14583
rect 14108 14549 14142 14583
rect 14178 14549 14192 14583
rect 14655 14565 14689 14596
rect 13176 14496 13210 14530
rect 13176 14428 13210 14462
rect 13176 14360 13210 14394
rect 5087 14242 5121 14274
rect 5087 14172 5121 14206
rect 5087 14104 5121 14136
rect 5087 14036 5121 14064
rect 5087 13968 5121 13992
rect 5087 13900 5121 13920
rect 5087 13832 5121 13848
rect 5087 13764 5121 13776
rect 5087 13696 5121 13704
rect 5087 13628 5121 13632
rect 5087 13593 5121 13594
rect 5087 13520 5121 13526
rect 5087 13447 5121 13458
rect 5087 13374 5121 13390
rect 5087 13301 5121 13322
rect 5087 13228 5121 13254
rect 5087 13155 5121 13186
rect 5087 13084 5121 13118
rect 5087 13016 5121 13048
rect 3079 12926 3113 12960
rect 4487 12962 4503 12965
rect 4487 12931 4501 12962
rect 4537 12931 4571 12965
rect 4605 12962 4621 12965
rect 4607 12931 4621 12962
rect 4743 12962 4759 12965
rect 4743 12931 4757 12962
rect 4793 12931 4827 12965
rect 4861 12962 4877 12965
rect 4863 12931 4877 12962
rect 5087 12948 5121 12975
rect 4535 12928 4573 12931
rect 4791 12928 4829 12931
rect 3079 12858 3113 12892
rect 3079 12790 3113 12824
rect 3079 12722 3113 12756
rect 3079 12576 3113 12688
rect 3079 12508 3113 12542
rect 3079 12440 3113 12474
rect 3079 12372 3113 12406
rect 5087 12880 5121 12902
rect 5087 12812 5121 12829
rect 5087 12744 5121 12756
rect 5087 12676 5121 12683
rect 5087 12608 5121 12610
rect 5087 12571 5121 12574
rect 5087 12498 5121 12506
rect 5410 14307 5478 14341
rect 5512 14307 5546 14341
rect 5580 14307 5614 14341
rect 5648 14307 5682 14341
rect 5716 14307 5750 14341
rect 5784 14307 5818 14341
rect 5852 14307 5886 14341
rect 5920 14307 5954 14341
rect 5988 14307 6022 14341
rect 6056 14307 6090 14341
rect 6124 14307 6158 14341
rect 6192 14307 6226 14341
rect 6260 14307 6294 14341
rect 6328 14307 6362 14341
rect 6396 14307 6430 14341
rect 6464 14307 6498 14341
rect 6532 14307 6566 14341
rect 6600 14307 6634 14341
rect 6668 14307 6702 14341
rect 6736 14307 6770 14341
rect 6804 14307 6838 14341
rect 6872 14307 6906 14341
rect 6940 14307 6974 14341
rect 7008 14307 7042 14341
rect 7076 14307 7110 14341
rect 7144 14307 7178 14341
rect 7212 14307 7246 14341
rect 7280 14307 7314 14341
rect 7348 14307 7382 14341
rect 7416 14307 7450 14341
rect 7484 14307 7518 14341
rect 7552 14307 7586 14341
rect 7620 14307 7654 14341
rect 7688 14307 7722 14341
rect 7756 14307 7790 14341
rect 7824 14307 7858 14341
rect 7892 14307 7926 14341
rect 7960 14307 7994 14341
rect 8028 14307 8062 14341
rect 8096 14307 8130 14341
rect 8164 14307 8198 14341
rect 8232 14307 8266 14341
rect 8300 14307 8334 14341
rect 8368 14307 8402 14341
rect 8436 14307 8470 14341
rect 8504 14307 8538 14341
rect 8572 14307 8606 14341
rect 8640 14307 8674 14341
rect 8708 14307 8742 14341
rect 8776 14307 8810 14341
rect 8844 14307 8878 14341
rect 8912 14307 8946 14341
rect 8980 14307 9014 14341
rect 9048 14307 9082 14341
rect 9116 14307 9150 14341
rect 9184 14307 9265 14341
rect 5410 14241 5444 14307
rect 5410 14173 5444 14207
rect 5410 14105 5444 14139
rect 9231 14273 9265 14307
rect 9231 14205 9265 14239
rect 9231 14137 9265 14171
rect 8693 14124 8835 14132
rect 8693 14090 8709 14124
rect 8749 14090 8785 14124
rect 8821 14090 8835 14124
rect 8693 14082 8835 14090
rect 5410 14037 5444 14071
rect 5410 13969 5444 14003
rect 5410 13901 5444 13935
rect 9231 14069 9265 14103
rect 9231 14001 9265 14035
rect 9231 13933 9265 13967
rect 5410 13833 5444 13867
rect 5740 13885 5882 13892
rect 5774 13884 5812 13885
rect 5846 13884 5882 13885
rect 5790 13851 5812 13884
rect 5740 13850 5756 13851
rect 5790 13850 5832 13851
rect 5866 13850 5882 13884
rect 5740 13842 5882 13850
rect 9231 13865 9265 13899
rect 5410 13765 5444 13799
rect 9231 13797 9265 13831
rect 5410 13697 5444 13731
rect 9003 13730 9145 13738
rect 9003 13696 9019 13730
rect 9053 13696 9091 13730
rect 9129 13696 9145 13730
rect 9003 13688 9145 13696
rect 9231 13729 9265 13763
rect 5410 13629 5444 13663
rect 5410 13561 5444 13595
rect 5410 13493 5444 13527
rect 5410 13425 5444 13459
rect 5410 13357 5444 13391
rect 5410 13289 5444 13323
rect 5410 13221 5444 13255
rect 5410 13153 5444 13187
rect 5410 13085 5444 13119
rect 5410 13017 5444 13051
rect 5410 12949 5444 12983
rect 5410 12881 5444 12915
rect 5410 12813 5444 12847
rect 5410 12745 5444 12779
rect 5410 12677 5444 12711
rect 9231 13661 9265 13695
rect 9231 13593 9265 13627
rect 13176 14292 13210 14326
rect 13176 14224 13210 14258
rect 13176 14156 13210 14190
rect 13176 14088 13210 14122
rect 13176 14020 13210 14054
rect 13176 13952 13210 13986
rect 13176 13884 13210 13918
rect 13176 13816 13210 13850
rect 13176 13748 13210 13782
rect 13176 13680 13210 13714
rect 13176 13612 13210 13646
rect 9231 13525 9265 13559
rect 9231 13457 9265 13491
rect 9231 13389 9265 13423
rect 9231 13321 9265 13355
rect 9231 13253 9265 13287
rect 9231 13185 9265 13219
rect 9231 13117 9265 13151
rect 9231 13049 9265 13083
rect 9231 12981 9265 13015
rect 9231 12913 9265 12947
rect 9231 12845 9265 12879
rect 9231 12777 9265 12811
rect 9231 12709 9265 12743
rect 9231 12658 9265 12675
rect 5410 12609 5444 12643
rect 8995 12650 9265 12658
rect 8995 12616 9011 12650
rect 9045 12616 9087 12650
rect 9121 12641 9265 12650
rect 9121 12616 9231 12641
rect 8995 12608 9231 12616
rect 5410 12541 5444 12575
rect 5410 12473 5444 12507
rect 9231 12573 9265 12607
rect 9231 12473 9265 12539
rect 5410 12439 5524 12473
rect 5558 12439 5592 12473
rect 5626 12439 5660 12473
rect 5694 12439 5728 12473
rect 5762 12439 5796 12473
rect 5830 12439 5864 12473
rect 5898 12439 5932 12473
rect 5966 12439 6000 12473
rect 6034 12439 6068 12473
rect 6102 12439 6136 12473
rect 6170 12439 6204 12473
rect 6238 12439 6272 12473
rect 6306 12439 6340 12473
rect 6374 12439 6408 12473
rect 6442 12439 6476 12473
rect 6510 12439 6544 12473
rect 6578 12439 6612 12473
rect 6646 12439 6680 12473
rect 6714 12439 6748 12473
rect 6782 12439 6816 12473
rect 6850 12439 6884 12473
rect 6918 12439 6952 12473
rect 6986 12439 7020 12473
rect 7054 12439 7088 12473
rect 7122 12439 7156 12473
rect 7190 12439 7224 12473
rect 7258 12439 7292 12473
rect 7326 12439 7360 12473
rect 7394 12439 7428 12473
rect 7462 12439 7496 12473
rect 7530 12439 7564 12473
rect 7598 12439 7632 12473
rect 7666 12439 7700 12473
rect 7734 12439 7768 12473
rect 7802 12439 7836 12473
rect 7870 12439 7939 12473
rect 7973 12439 8007 12473
rect 8041 12439 8075 12473
rect 8109 12439 8143 12473
rect 8177 12439 8211 12473
rect 8245 12439 8279 12473
rect 8313 12439 8347 12473
rect 8381 12439 8415 12473
rect 8449 12439 8483 12473
rect 8517 12439 8551 12473
rect 8585 12439 8619 12473
rect 8653 12439 8687 12473
rect 8721 12439 8755 12473
rect 8789 12439 8823 12473
rect 8857 12439 8891 12473
rect 8925 12439 8959 12473
rect 8993 12439 9027 12473
rect 9061 12439 9095 12473
rect 9129 12439 9163 12473
rect 9197 12439 9265 12473
rect 11686 13572 11758 13606
rect 11805 13572 11839 13606
rect 11875 13572 11907 13606
rect 11958 13572 11975 13606
rect 12041 13572 12043 13606
rect 12077 13572 12090 13606
rect 12145 13572 12179 13606
rect 12213 13572 12247 13606
rect 12281 13572 12315 13606
rect 12349 13572 12383 13606
rect 12417 13572 12451 13606
rect 12485 13572 12519 13606
rect 12553 13572 12565 13606
rect 12621 13572 12642 13606
rect 12689 13572 12719 13606
rect 12757 13572 12825 13606
rect 11686 13538 11720 13572
rect 11686 13470 11720 13499
rect 11686 13402 11720 13426
rect 12791 13533 12825 13572
rect 12791 13485 12825 13499
rect 11686 13334 11720 13353
rect 11686 13266 11720 13280
rect 11686 13198 11720 13207
rect 11686 13130 11720 13134
rect 11686 13095 11720 13096
rect 11686 13022 11720 13028
rect 11686 12949 11720 12960
rect 11686 12875 11720 12892
rect 11686 12801 11720 12824
rect 11686 12727 11720 12756
rect 11686 12654 11720 12688
rect 11686 12586 11720 12619
rect 11686 12518 11720 12545
rect 11686 12450 11720 12471
rect 5087 12425 5121 12438
rect 3286 12356 3300 12390
rect 3336 12356 3370 12390
rect 3406 12356 3420 12390
rect 3522 12356 3536 12390
rect 3572 12356 3606 12390
rect 3642 12356 3656 12390
rect 3758 12356 3772 12390
rect 3808 12356 3842 12390
rect 3878 12356 3892 12390
rect 3994 12356 4008 12390
rect 4044 12356 4078 12390
rect 4114 12356 4128 12390
rect 3079 12304 3113 12338
rect 3079 12236 3113 12270
rect 3079 12168 3113 12202
rect 3079 12100 3113 12134
rect -564 12006 -530 12040
rect -343 12008 -329 12042
rect -293 12008 -259 12042
rect -223 12008 -73 12042
rect -37 12008 -3 12042
rect 33 12008 47 12042
rect 235 12008 249 12042
rect 285 12008 319 12042
rect 355 12008 369 12042
rect 3079 12032 3113 12066
rect 5087 12352 5121 12370
rect 5087 12279 5121 12302
rect 5087 12206 5121 12234
rect 5087 12132 5121 12166
rect 5087 12064 5121 12098
rect 3079 11964 3113 11998
rect 4448 11981 4462 12015
rect 4498 11981 4532 12015
rect 4568 11981 4582 12015
rect 4704 11981 4718 12015
rect 4754 11981 4788 12015
rect 4824 11981 4838 12015
rect 5087 11996 5121 12030
rect 3079 11896 3113 11930
rect 5087 11896 5121 11962
rect 3079 11862 3183 11896
rect 3217 11862 3251 11896
rect 3285 11862 3319 11896
rect 3353 11862 3387 11896
rect 3421 11862 3455 11896
rect 3489 11862 3523 11896
rect 3557 11862 3591 11896
rect 3625 11862 3659 11896
rect 3693 11862 3727 11896
rect 3761 11862 3795 11896
rect 3829 11862 3863 11896
rect 3897 11862 3931 11896
rect 3965 11862 3999 11896
rect 4033 11862 4067 11896
rect 4101 11862 4135 11896
rect 4169 11862 4203 11896
rect 4237 11862 4271 11896
rect 4305 11862 4339 11896
rect 4373 11862 4407 11896
rect 4441 11862 4475 11896
rect 4509 11862 4543 11896
rect 4577 11862 4611 11896
rect 4645 11862 4679 11896
rect 4713 11862 4747 11896
rect 4781 11862 4815 11896
rect 4849 11862 4883 11896
rect 4917 11862 4951 11896
rect 4985 11862 5019 11896
rect 5053 11862 5121 11896
rect 11686 12382 11720 12397
rect 11686 12314 11720 12323
rect 11868 13418 12106 13424
rect 12476 13418 12640 13424
rect 11868 13384 11880 13418
rect 11914 13384 11952 13418
rect 11986 13384 11988 13418
rect 12022 13384 12024 13418
rect 12090 13384 12124 13418
rect 12158 13384 12192 13418
rect 12226 13384 12260 13418
rect 12294 13384 12328 13418
rect 12362 13384 12396 13418
rect 12430 13384 12464 13418
rect 12498 13384 12522 13418
rect 12566 13384 12594 13418
rect 12628 13384 12640 13418
rect 11868 13378 12106 13384
rect 12476 13378 12640 13384
rect 11868 13350 11914 13378
rect 11868 13285 11874 13350
rect 11908 13285 11914 13350
rect 11868 13282 11914 13285
rect 11868 13248 11874 13282
rect 11908 13248 11914 13282
rect 11868 13247 11914 13248
rect 12594 13340 12640 13378
rect 12594 13300 12600 13340
rect 12634 13300 12640 13340
rect 12594 13268 12640 13300
rect 11868 13180 11874 13247
rect 11908 13180 11914 13247
rect 11868 13175 11914 13180
rect 11868 13112 11874 13175
rect 11908 13112 11914 13175
rect 11868 13103 11914 13112
rect 11868 13044 11874 13103
rect 11908 13044 11914 13103
rect 11868 13031 11914 13044
rect 11868 12976 11874 13031
rect 11908 12976 11914 13031
rect 11868 12959 11914 12976
rect 11868 12908 11874 12959
rect 11908 12908 11914 12959
rect 11868 12887 11914 12908
rect 11868 12840 11874 12887
rect 11908 12840 11914 12887
rect 11868 12815 11914 12840
rect 11868 12772 11874 12815
rect 11908 12772 11914 12815
rect 11868 12743 11914 12772
rect 11868 12704 11874 12743
rect 11908 12704 11914 12743
rect 11868 12671 11914 12704
rect 11868 12636 11874 12671
rect 11908 12636 11914 12671
rect 11868 12602 11914 12636
rect 11868 12565 11874 12602
rect 11908 12565 11914 12602
rect 11868 12534 11914 12565
rect 11868 12493 11874 12534
rect 11908 12493 11914 12534
rect 12226 13170 12260 13213
rect 12226 13093 12260 13136
rect 12226 13016 12260 13059
rect 12226 12939 12260 12982
rect 12226 12862 12260 12905
rect 12226 12785 12260 12828
rect 12226 12708 12260 12751
rect 12226 12631 12260 12674
rect 12226 12554 12260 12597
rect 12594 13232 12600 13268
rect 12634 13232 12640 13268
rect 12594 13198 12640 13232
rect 12594 13162 12600 13198
rect 12634 13162 12640 13198
rect 12594 13130 12640 13162
rect 12594 13090 12600 13130
rect 12634 13090 12640 13130
rect 12594 13062 12640 13090
rect 12594 13018 12600 13062
rect 12634 13018 12640 13062
rect 12594 12994 12640 13018
rect 12594 12946 12600 12994
rect 12634 12946 12640 12994
rect 12594 12926 12640 12946
rect 12594 12874 12600 12926
rect 12634 12874 12640 12926
rect 12594 12858 12640 12874
rect 12594 12802 12600 12858
rect 12634 12802 12640 12858
rect 12594 12790 12640 12802
rect 12594 12730 12600 12790
rect 12634 12730 12640 12790
rect 12594 12722 12640 12730
rect 12594 12658 12600 12722
rect 12634 12658 12640 12722
rect 12594 12654 12640 12658
rect 12594 12552 12600 12654
rect 12634 12552 12640 12654
rect 12594 12548 12640 12552
rect 11868 12466 11914 12493
rect 11868 12421 11874 12466
rect 11908 12421 11914 12466
rect 11868 12398 11914 12421
rect 11868 12349 11874 12398
rect 11908 12349 11914 12398
rect 11868 12330 11914 12349
rect 11868 12277 11874 12330
rect 11908 12277 11914 12330
rect 11868 12265 11914 12277
rect 12594 12484 12600 12548
rect 12634 12484 12640 12548
rect 12594 12476 12640 12484
rect 12594 12416 12600 12476
rect 12634 12416 12640 12476
rect 12594 12404 12640 12416
rect 12594 12348 12600 12404
rect 12634 12348 12640 12404
rect 12594 12332 12640 12348
rect 12594 12280 12600 12332
rect 12634 12280 12640 12332
rect 11686 12246 11720 12249
rect 11686 12178 11720 12212
rect 11686 12110 11720 12144
rect 11686 12042 11720 12076
rect 11874 12262 11908 12265
rect 11874 12116 11908 12228
rect 12594 12260 12640 12280
rect 12594 12212 12600 12260
rect 12634 12212 12640 12260
rect 12048 12193 12064 12195
rect 12048 12161 12062 12193
rect 12098 12161 12132 12195
rect 12166 12193 12182 12195
rect 12168 12161 12182 12193
rect 12304 12193 12320 12195
rect 12304 12161 12318 12193
rect 12354 12161 12388 12195
rect 12422 12193 12438 12195
rect 12424 12161 12438 12193
rect 12594 12188 12640 12212
rect 12096 12159 12134 12161
rect 12352 12159 12390 12161
rect 12594 12144 12600 12188
rect 12634 12144 12640 12188
rect 12594 12116 12640 12144
rect 11874 12110 12600 12116
rect 11874 12076 11886 12110
rect 11920 12076 11942 12110
rect 11992 12076 12010 12110
rect 12064 12076 12078 12110
rect 12136 12076 12146 12110
rect 12208 12076 12214 12110
rect 12280 12076 12282 12110
rect 12316 12076 12318 12110
rect 12384 12076 12390 12110
rect 12452 12076 12462 12110
rect 12520 12082 12600 12110
rect 12634 12082 12640 12116
rect 12520 12076 12640 12082
rect 11874 12070 12640 12076
rect 12791 13417 12825 13426
rect 12791 13349 12825 13353
rect 12791 13314 12825 13315
rect 12791 13241 12825 13247
rect 12791 13168 12825 13179
rect 12791 13095 12825 13111
rect 12791 13022 12825 13043
rect 12791 12949 12825 12975
rect 12791 12876 12825 12907
rect 12791 12805 12825 12839
rect 12791 12737 12825 12769
rect 12791 12669 12825 12696
rect 12791 12601 12825 12623
rect 12791 12533 12825 12549
rect 12791 12465 12825 12475
rect 12791 12397 12825 12401
rect 12791 12361 12825 12363
rect 12791 12287 12825 12295
rect 12791 12213 12825 12227
rect 12791 12139 12825 12159
rect 11686 11921 11720 12008
rect 12791 12057 12825 12091
rect 12791 11989 12825 12023
rect 13176 13544 13210 13578
rect 13176 13476 13210 13510
rect 13176 13408 13210 13442
rect 13176 13340 13210 13374
rect 14655 14494 14689 14528
rect 14655 14426 14689 14450
rect 14655 14358 14689 14378
rect 14655 14290 14689 14306
rect 14655 14222 14689 14234
rect 14655 14154 14689 14162
rect 14655 14086 14689 14090
rect 14655 13980 14689 13984
rect 14655 13908 14689 13916
rect 14655 13836 14689 13848
rect 14655 13764 14689 13780
rect 14655 13692 14689 13712
rect 14655 13620 14689 13644
rect 14655 13548 14689 13576
rect 14655 13476 14689 13508
rect 14655 13406 14689 13440
rect 13542 13335 13556 13369
rect 13592 13335 13626 13369
rect 13662 13335 13676 13369
rect 13798 13335 13812 13369
rect 13848 13335 13882 13369
rect 13918 13335 14068 13369
rect 14104 13335 14138 13369
rect 14174 13335 14188 13369
rect 14310 13335 14324 13369
rect 14360 13335 14394 13369
rect 14430 13335 14444 13369
rect 14655 13338 14689 13370
rect 13176 13272 13210 13306
rect 13176 13204 13210 13238
rect 13176 13136 13210 13170
rect 13176 13068 13210 13102
rect 13176 13000 13210 13034
rect 13176 12932 13210 12966
rect 13176 12864 13210 12898
rect 13176 12796 13210 12830
rect 13176 12728 13210 12762
rect 13176 12660 13210 12694
rect 13176 12592 13210 12626
rect 13176 12524 13210 12558
rect 13176 12456 13210 12490
rect 13176 12388 13210 12422
rect 13176 12320 13210 12354
rect 13176 12252 13210 12286
rect 13176 12184 13210 12218
rect 14655 13270 14689 13298
rect 14655 13202 14689 13226
rect 14655 13134 14689 13154
rect 14655 13066 14689 13082
rect 14655 12998 14689 13010
rect 14655 12930 14689 12938
rect 14655 12862 14689 12866
rect 14655 12827 14689 12828
rect 14655 12754 14689 12760
rect 14655 12681 14689 12692
rect 14655 12608 14689 12624
rect 14655 12535 14689 12556
rect 14655 12462 14689 12488
rect 14655 12389 14689 12420
rect 14655 12318 14689 12352
rect 14655 12250 14689 12282
rect 14655 12182 14689 12209
rect 13176 12116 13210 12150
rect 13802 12134 13816 12168
rect 13852 12134 13886 12168
rect 13922 12134 13936 12168
rect 14058 12134 14072 12168
rect 14108 12134 14142 12168
rect 14178 12134 14192 12168
rect 13176 12048 13210 12082
rect 14655 12097 14689 12136
rect 14655 12048 14689 12063
rect 13176 12014 13248 12048
rect 13282 12014 13316 12048
rect 13350 12014 13384 12048
rect 13418 12014 13452 12048
rect 13486 12014 13520 12048
rect 13554 12014 13588 12048
rect 13622 12014 13656 12048
rect 13690 12014 13724 12048
rect 13758 12014 13792 12048
rect 13826 12014 13860 12048
rect 13894 12014 13928 12048
rect 13962 12014 13996 12048
rect 14030 12014 14064 12048
rect 14098 12014 14132 12048
rect 14166 12014 14200 12048
rect 14234 12014 14268 12048
rect 14302 12014 14336 12048
rect 14370 12014 14404 12048
rect 14438 12014 14472 12048
rect 14506 12014 14587 12048
rect 14621 12014 14689 12048
rect 12791 11921 12825 11955
rect 11686 11887 11754 11921
rect 11788 11887 11822 11921
rect 11856 11887 11890 11921
rect 11924 11887 11958 11921
rect 11992 11887 12026 11921
rect 12060 11887 12094 11921
rect 12128 11887 12162 11921
rect 12196 11887 12230 11921
rect 12264 11887 12298 11921
rect 12332 11887 12366 11921
rect 12400 11887 12434 11921
rect 12468 11887 12502 11921
rect 12536 11887 12570 11921
rect 12604 11887 12638 11921
rect 12672 11887 12706 11921
rect 12740 11887 12825 11921
rect 7823 8219 12931 8220
rect 7823 8185 7857 8219
rect 7891 8185 7925 8219
rect 7959 8185 7993 8219
rect 8027 8185 8061 8219
rect 8095 8185 8129 8219
rect 8163 8185 8197 8219
rect 8231 8185 8265 8219
rect 8299 8185 8333 8219
rect 8367 8185 8401 8219
rect 8435 8185 8469 8219
rect 8503 8185 8537 8219
rect 8571 8185 8605 8219
rect 8639 8185 8673 8219
rect 8707 8185 8741 8219
rect 8775 8185 8809 8219
rect 8843 8185 8877 8219
rect 8911 8185 8945 8219
rect 8979 8185 9013 8219
rect 9047 8185 9081 8219
rect 9115 8185 9149 8219
rect 9183 8185 9217 8219
rect 9251 8185 9285 8219
rect 9319 8185 9353 8219
rect 9387 8185 9421 8219
rect 9455 8185 9489 8219
rect 9523 8185 9557 8219
rect 9591 8185 9625 8219
rect 9659 8185 9693 8219
rect 9727 8185 9761 8219
rect 9795 8185 9829 8219
rect 9863 8185 9897 8219
rect 9931 8185 9965 8219
rect 9999 8185 10033 8219
rect 10067 8185 10101 8219
rect 10135 8185 10169 8219
rect 10203 8185 10237 8219
rect 10271 8185 10305 8219
rect 10339 8185 10373 8219
rect 10407 8185 10441 8219
rect 10475 8185 10509 8219
rect 10543 8185 10577 8219
rect 10611 8185 10645 8219
rect 10679 8185 10713 8219
rect 10747 8185 10781 8219
rect 10815 8185 10849 8219
rect 10883 8185 10917 8219
rect 10951 8185 10985 8219
rect 11019 8185 11053 8219
rect 11087 8185 11121 8219
rect 11155 8185 11189 8219
rect 11223 8185 11257 8219
rect 11291 8185 11325 8219
rect 11359 8185 11393 8219
rect 11427 8185 11461 8219
rect 11495 8185 11529 8219
rect 11563 8185 11597 8219
rect 11631 8185 11665 8219
rect 11699 8185 11733 8219
rect 11767 8185 11801 8219
rect 11835 8185 11869 8219
rect 11903 8185 11937 8219
rect 11971 8185 12005 8219
rect 12039 8185 12073 8219
rect 12107 8185 12141 8219
rect 12175 8185 12209 8219
rect 12243 8185 12277 8219
rect 12311 8185 12345 8219
rect 12379 8185 12413 8219
rect 12447 8185 12481 8219
rect 12515 8185 12549 8219
rect 12583 8185 12617 8219
rect 12651 8185 12685 8219
rect 12719 8185 12753 8219
rect 12787 8185 12821 8219
rect 12855 8186 12931 8219
rect 12855 8185 12896 8186
rect 7823 8184 12896 8185
rect 7823 8151 7859 8184
rect 7823 8117 7824 8151
rect 7858 8117 7859 8151
rect 7823 8083 7859 8117
rect 7823 8049 7824 8083
rect 7858 8049 7859 8083
rect 7823 8015 7859 8049
rect 12895 8152 12896 8184
rect 12930 8152 12931 8186
rect 12895 8118 12931 8152
rect 12895 8084 12896 8118
rect 12930 8084 12931 8118
rect 12895 8050 12931 8084
rect 7823 7981 7824 8015
rect 7858 7981 7859 8015
rect 7823 7947 7859 7981
rect 7823 7913 7824 7947
rect 7858 7913 7859 7947
rect 7823 7879 7859 7913
rect 7823 7845 7824 7879
rect 7858 7845 7859 7879
rect 7823 7811 7859 7845
rect 7823 7777 7824 7811
rect 7858 7777 7859 7811
rect 7823 7743 7859 7777
rect 7823 7709 7824 7743
rect 7858 7709 7859 7743
rect 7823 7675 7859 7709
rect 7823 7641 7824 7675
rect 7858 7641 7859 7675
rect 7823 7607 7859 7641
rect 7823 7575 7824 7607
rect 3894 7574 7824 7575
rect 3894 7540 3901 7574
rect 3962 7540 3974 7574
rect 4030 7540 4047 7574
rect 4098 7540 4120 7574
rect 4166 7540 4193 7574
rect 4234 7540 4266 7574
rect 4302 7540 4336 7574
rect 4373 7540 4404 7574
rect 4446 7540 4472 7574
rect 4519 7540 4540 7574
rect 4592 7540 4608 7574
rect 4665 7540 4676 7574
rect 4738 7540 4744 7574
rect 4811 7540 4812 7574
rect 4846 7540 4850 7574
rect 4914 7540 4923 7574
rect 4982 7540 4996 7574
rect 5050 7540 5069 7574
rect 5118 7540 5142 7574
rect 5186 7540 5215 7574
rect 5254 7540 5288 7574
rect 5322 7540 5356 7574
rect 5395 7540 5424 7574
rect 5468 7540 5492 7574
rect 5541 7540 5560 7574
rect 5614 7540 5628 7574
rect 5687 7540 5696 7574
rect 5760 7540 5764 7574
rect 5798 7540 5799 7574
rect 5866 7540 5872 7574
rect 5934 7540 5945 7574
rect 6002 7540 6018 7574
rect 6070 7540 6091 7574
rect 6138 7540 6164 7574
rect 6206 7540 6237 7574
rect 6274 7540 6308 7574
rect 6344 7540 6376 7574
rect 6417 7540 6444 7574
rect 6490 7540 6512 7574
rect 6564 7540 6580 7574
rect 6638 7540 6648 7574
rect 6712 7540 6716 7574
rect 6750 7540 6752 7574
rect 6818 7540 6826 7574
rect 6886 7540 6900 7574
rect 6954 7540 6974 7574
rect 7022 7540 7048 7574
rect 7090 7540 7122 7574
rect 7158 7540 7192 7574
rect 7230 7540 7260 7574
rect 7304 7540 7328 7574
rect 7378 7540 7396 7574
rect 7452 7540 7464 7574
rect 7526 7540 7532 7574
rect 7634 7540 7640 7574
rect 7702 7540 7714 7574
rect 7770 7573 7824 7574
rect 7858 7573 7859 7607
rect 7770 7540 7859 7573
rect 3894 7539 7859 7540
rect 7925 7999 8221 8033
rect 3894 7495 3930 7539
rect 3894 7449 3895 7495
rect 3929 7449 3930 7495
rect 3894 7427 3930 7449
rect 3894 7367 3895 7427
rect 3929 7367 3930 7427
rect 4796 7463 4830 7539
rect 4796 7395 4830 7429
rect 3894 7359 3930 7367
rect 3894 7325 3895 7359
rect 3929 7325 3930 7359
rect 3894 7319 3930 7325
rect 3894 7257 3895 7319
rect 3929 7257 3930 7319
rect 3894 7237 3930 7257
rect 3894 7189 3895 7237
rect 3929 7189 3930 7237
rect 3894 7155 3930 7189
rect 3894 7121 3895 7155
rect 3929 7121 3930 7155
rect 3894 7087 3930 7121
rect 3894 7040 3895 7087
rect 3929 7040 3930 7087
rect 3894 7019 3930 7040
rect 3894 6959 3895 7019
rect 3929 6959 3930 7019
rect 3894 6951 3930 6959
rect 3894 6917 3895 6951
rect 3929 6917 3930 6951
rect 3894 6883 3930 6917
rect 3894 6849 3895 6883
rect 3929 6849 3930 6883
rect 4108 7352 4180 7386
rect 4214 7352 4248 7386
rect 4305 7352 4316 7386
rect 4350 7352 4361 7386
rect 4418 7352 4452 7386
rect 4486 7352 4520 7386
rect 4554 7352 4622 7386
rect 4108 7318 4142 7352
rect 4108 7250 4142 7268
rect 4588 7299 4622 7352
rect 4588 7231 4622 7265
rect 4108 7182 4142 7184
rect 4108 7133 4142 7148
rect 4108 7048 4142 7080
rect 4482 7182 4516 7193
rect 4482 7110 4516 7143
rect 4482 7059 4516 7075
rect 4588 7163 4622 7197
rect 4588 7095 4622 7129
rect 4108 6978 4142 7012
rect 4108 6891 4142 6929
rect 4588 7027 4622 7061
rect 4588 6959 4622 6993
rect 4588 6891 4622 6925
rect 4108 6857 4176 6891
rect 4215 6857 4244 6891
rect 4288 6857 4312 6891
rect 4361 6857 4380 6891
rect 4434 6857 4448 6891
rect 4507 6857 4546 6891
rect 4580 6857 4622 6891
rect 5656 7463 5690 7539
rect 5656 7395 5690 7429
rect 4796 7327 4830 7361
rect 4796 7259 4830 7293
rect 4796 7191 4830 7225
rect 4796 7123 4830 7157
rect 4796 7055 4830 7089
rect 4796 6987 4830 7021
rect 4796 6919 4830 6953
rect 3894 6815 3930 6849
rect 3894 6781 3895 6815
rect 3929 6781 3930 6815
rect 3894 6747 3930 6781
rect 3894 6713 3895 6747
rect 3929 6713 3930 6747
rect 3894 6679 3930 6713
rect 3894 6645 3895 6679
rect 3929 6645 3930 6679
rect 3894 6611 3930 6645
rect 3894 6577 3895 6611
rect 3929 6579 3930 6611
rect 4796 6851 4830 6885
rect 4988 7352 5005 7386
rect 5039 7352 5060 7386
rect 5117 7352 5128 7386
rect 5195 7352 5196 7386
rect 5230 7352 5239 7386
rect 5298 7352 5317 7386
rect 5366 7352 5396 7386
rect 5434 7352 5502 7386
rect 4988 7318 5022 7352
rect 4988 7250 5022 7284
rect 4988 7182 5022 7216
rect 5468 7301 5502 7352
rect 5468 7231 5502 7265
rect 4988 7114 5022 7148
rect 4988 7046 5022 7080
rect 5365 7182 5399 7193
rect 5365 7110 5399 7143
rect 5365 7059 5399 7075
rect 5468 7163 5502 7181
rect 4988 6978 5022 7012
rect 4988 6891 5022 6944
rect 5468 7027 5502 7061
rect 5468 6959 5502 6993
rect 5468 6912 5502 6925
rect 4988 6857 5000 6891
rect 5034 6857 5056 6891
rect 5112 6857 5124 6891
rect 5190 6857 5192 6891
rect 5226 6857 5234 6891
rect 5294 6857 5312 6891
rect 5362 6857 5390 6891
rect 5424 6878 5468 6891
rect 5424 6857 5502 6878
rect 6666 7463 6700 7539
rect 6666 7395 6700 7429
rect 5656 7327 5690 7361
rect 5656 7259 5690 7293
rect 5656 7191 5690 7225
rect 5656 7123 5690 7157
rect 5656 7055 5690 7089
rect 5656 6987 5690 7021
rect 5656 6919 5690 6953
rect 4796 6783 4830 6817
rect 4796 6715 4830 6749
rect 4796 6647 4830 6681
rect 4796 6579 4830 6613
rect 5656 6851 5690 6885
rect 5850 7352 5890 7386
rect 5956 7352 5963 7386
rect 6024 7352 6036 7386
rect 6092 7352 6110 7386
rect 6160 7352 6184 7386
rect 6228 7352 6258 7386
rect 6296 7352 6364 7386
rect 5850 7318 5884 7352
rect 5850 7250 5884 7284
rect 5850 7182 5884 7216
rect 6330 7312 6364 7352
rect 6330 7238 6364 7265
rect 5850 7114 5884 7148
rect 5850 7046 5884 7080
rect 6223 7182 6257 7193
rect 6223 7110 6257 7143
rect 6223 7059 6257 7075
rect 6330 7163 6364 7197
rect 6330 7095 6364 7129
rect 5850 6978 5884 7012
rect 5850 6891 5884 6944
rect 6330 7027 6364 7061
rect 6330 6959 6364 6993
rect 6330 6891 6364 6925
rect 7669 7463 7703 7539
rect 7669 7395 7703 7429
rect 6666 7327 6700 7361
rect 6666 7259 6700 7293
rect 6666 7191 6700 7225
rect 6666 7123 6700 7157
rect 6666 7055 6700 7089
rect 6666 6987 6700 7021
rect 6666 6919 6700 6953
rect 5850 6857 5913 6891
rect 5952 6857 5986 6891
rect 6029 6857 6054 6891
rect 6106 6857 6122 6891
rect 6183 6857 6190 6891
rect 6255 6857 6340 6891
rect 5656 6783 5690 6817
rect 5656 6715 5690 6749
rect 5656 6647 5690 6681
rect 5656 6579 5690 6613
rect 6666 6851 6700 6885
rect 6980 7352 7008 7386
rect 7042 7352 7052 7386
rect 7086 7352 7090 7386
rect 7154 7352 7172 7386
rect 7222 7352 7254 7386
rect 7290 7352 7324 7386
rect 7358 7352 7392 7386
rect 7426 7352 7494 7386
rect 6980 7318 7014 7352
rect 6980 7250 7014 7284
rect 6980 7182 7014 7216
rect 7460 7302 7494 7352
rect 7460 7231 7494 7265
rect 6980 7114 7014 7148
rect 6980 7046 7014 7080
rect 7359 7179 7393 7193
rect 7359 7109 7393 7143
rect 7359 7059 7393 7073
rect 7460 7163 7494 7184
rect 7460 7095 7494 7099
rect 6980 6994 7014 7012
rect 6980 6891 7014 6944
rect 7460 7048 7494 7061
rect 7460 6963 7494 6993
rect 7460 6891 7494 6925
rect 6980 6857 7048 6891
rect 7086 6857 7116 6891
rect 7168 6857 7184 6891
rect 7250 6857 7252 6891
rect 7286 6857 7298 6891
rect 7354 6857 7379 6891
rect 7413 6857 7494 6891
rect 7669 7327 7703 7361
rect 7669 7259 7703 7293
rect 7669 7191 7703 7225
rect 7669 7123 7703 7157
rect 7669 7055 7703 7089
rect 7669 6987 7703 7021
rect 7669 6919 7703 6953
rect 6666 6783 6700 6817
rect 6666 6715 6700 6749
rect 6666 6647 6700 6681
rect 6666 6579 6700 6613
rect 7669 6851 7703 6885
rect 7669 6783 7703 6817
rect 7669 6715 7703 6749
rect 7925 6766 7959 7999
rect 8199 7997 8221 7999
rect 8267 7997 8294 8031
rect 8335 7997 8367 8031
rect 8403 7997 8437 8031
rect 8474 7997 8505 8031
rect 8547 7997 8573 8031
rect 8620 7997 8641 8031
rect 8693 7997 8709 8031
rect 8766 7997 8777 8031
rect 8839 7997 8845 8031
rect 8912 7997 8913 8031
rect 8947 7997 8951 8031
rect 9015 7997 9024 8031
rect 9083 7997 9097 8031
rect 9151 7997 9170 8031
rect 9219 7997 9243 8031
rect 9287 7997 9316 8031
rect 9355 7997 9389 8031
rect 9423 7997 9457 8031
rect 9496 7997 9525 8031
rect 9569 7997 9593 8031
rect 9642 7997 9661 8031
rect 9715 7997 9729 8031
rect 9788 7997 9797 8031
rect 9861 7997 9865 8031
rect 9899 7997 9900 8031
rect 9967 7997 9973 8031
rect 10035 7997 10046 8031
rect 10103 7997 10119 8031
rect 10171 7997 10192 8031
rect 10239 7997 10265 8031
rect 10307 7997 10338 8031
rect 10375 7997 10409 8031
rect 10445 7997 10477 8031
rect 10518 7997 10545 8031
rect 10591 7997 10613 8031
rect 10664 7997 10681 8031
rect 10737 7997 10749 8031
rect 10810 7997 10817 8031
rect 10883 7997 10885 8031
rect 10919 7997 10922 8031
rect 10987 7997 10995 8031
rect 11055 7997 11068 8031
rect 11123 7997 11141 8031
rect 11191 7997 11214 8031
rect 11259 7997 11286 8031
rect 11327 7997 11358 8031
rect 11395 7997 11429 8031
rect 11464 7997 11497 8031
rect 11536 7997 11565 8031
rect 11608 7997 11633 8031
rect 11680 7997 11701 8031
rect 11752 7997 11769 8031
rect 11824 7997 11837 8031
rect 11896 7997 11905 8031
rect 11968 7997 11973 8031
rect 12040 7997 12041 8031
rect 12075 7997 12078 8031
rect 12143 7997 12150 8031
rect 12211 7997 12222 8031
rect 12279 7997 12294 8031
rect 12347 7997 12724 8031
rect 8105 7806 8139 7820
rect 8105 7736 8139 7770
rect 8105 7686 8139 7700
rect 10247 7806 10281 7820
rect 10247 7736 10281 7770
rect 10247 7686 10281 7700
rect 10423 7806 10457 7820
rect 10423 7736 10457 7770
rect 10423 7686 10457 7700
rect 12565 7806 12599 7820
rect 12565 7736 12599 7770
rect 12565 7686 12599 7700
rect 8105 7570 8139 7584
rect 8105 7500 8139 7534
rect 8105 7450 8139 7464
rect 10247 7570 10281 7584
rect 10247 7500 10281 7534
rect 10247 7450 10281 7464
rect 10423 7570 10457 7584
rect 10423 7500 10457 7534
rect 10423 7450 10457 7464
rect 12565 7570 12599 7584
rect 12565 7500 12599 7534
rect 12565 7450 12599 7464
rect 8105 7338 8139 7348
rect 8105 7266 8139 7298
rect 8105 7214 8139 7230
rect 10247 7334 10281 7348
rect 10247 7264 10281 7298
rect 10247 7214 10281 7228
rect 10423 7334 10457 7348
rect 10423 7264 10457 7298
rect 10423 7214 10457 7228
rect 12565 7334 12599 7348
rect 12565 7264 12599 7298
rect 12565 7214 12599 7228
rect 8105 7098 8139 7112
rect 8105 7028 8139 7062
rect 8105 6978 8139 6992
rect 10247 7098 10281 7112
rect 10247 7028 10281 7062
rect 10247 6978 10281 6992
rect 10423 7098 10457 7112
rect 10423 7028 10457 7062
rect 10423 6978 10457 6992
rect 12565 7098 12599 7112
rect 12565 7028 12599 7062
rect 12565 6978 12599 6992
rect 12690 6766 12724 7997
rect 7925 6732 8233 6766
rect 8267 6732 8301 6766
rect 8335 6732 8369 6766
rect 8403 6732 8437 6766
rect 8471 6732 8505 6766
rect 8539 6732 8573 6766
rect 8607 6732 8641 6766
rect 8675 6732 8709 6766
rect 8743 6732 8777 6766
rect 8811 6732 8845 6766
rect 8879 6732 8913 6766
rect 8947 6732 8981 6766
rect 9015 6732 9049 6766
rect 9083 6732 9117 6766
rect 9151 6732 9185 6766
rect 9219 6732 9253 6766
rect 9287 6732 9321 6766
rect 9355 6732 9389 6766
rect 9423 6732 9457 6766
rect 9491 6732 9525 6766
rect 9559 6732 9593 6766
rect 9627 6732 9661 6766
rect 9695 6732 9729 6766
rect 9763 6732 9797 6766
rect 9831 6732 9865 6766
rect 9899 6732 9933 6766
rect 9967 6732 10001 6766
rect 10035 6732 10069 6766
rect 10103 6732 10137 6766
rect 10171 6732 10205 6766
rect 10239 6732 10273 6766
rect 10307 6732 10341 6766
rect 10375 6732 10409 6766
rect 10443 6732 10477 6766
rect 10511 6732 10545 6766
rect 10579 6732 10613 6766
rect 10647 6732 10681 6766
rect 10715 6732 10749 6766
rect 10783 6732 10817 6766
rect 10851 6732 10885 6766
rect 10919 6732 10953 6766
rect 10987 6732 11021 6766
rect 11055 6732 11089 6766
rect 11123 6732 11157 6766
rect 11191 6732 11225 6766
rect 11259 6732 11293 6766
rect 11327 6732 11361 6766
rect 11395 6732 11429 6766
rect 11463 6732 11497 6766
rect 11531 6732 11565 6766
rect 11599 6732 11633 6766
rect 11667 6732 11701 6766
rect 11735 6732 11769 6766
rect 11803 6732 11837 6766
rect 11871 6732 11905 6766
rect 11939 6732 11973 6766
rect 12007 6732 12041 6766
rect 12075 6732 12109 6766
rect 12143 6732 12177 6766
rect 12211 6732 12245 6766
rect 12279 6732 12313 6766
rect 12347 6732 12724 6766
rect 12895 8016 12896 8050
rect 12930 8016 12931 8050
rect 12895 7982 12931 8016
rect 12895 7948 12896 7982
rect 12930 7948 12931 7982
rect 12895 7914 12931 7948
rect 12895 7880 12896 7914
rect 12930 7880 12931 7914
rect 12895 7846 12931 7880
rect 12895 7812 12896 7846
rect 12930 7812 12931 7846
rect 12895 7778 12931 7812
rect 12895 7744 12896 7778
rect 12930 7744 12931 7778
rect 12895 7710 12931 7744
rect 12895 7676 12896 7710
rect 12930 7676 12931 7710
rect 12895 7642 12931 7676
rect 12895 7608 12896 7642
rect 12930 7608 12931 7642
rect 12895 7574 12931 7608
rect 12895 7540 12896 7574
rect 12930 7540 12931 7574
rect 12895 7506 12931 7540
rect 12895 7472 12896 7506
rect 12930 7472 12931 7506
rect 12895 7438 12931 7472
rect 12895 7404 12896 7438
rect 12930 7404 12931 7438
rect 12895 7370 12931 7404
rect 12895 7336 12896 7370
rect 12930 7336 12931 7370
rect 12895 7302 12931 7336
rect 12895 7268 12896 7302
rect 12930 7268 12931 7302
rect 12895 7234 12931 7268
rect 12895 7200 12896 7234
rect 12930 7200 12931 7234
rect 12895 7166 12931 7200
rect 12895 7132 12896 7166
rect 12930 7132 12931 7166
rect 12895 7098 12931 7132
rect 12895 7064 12896 7098
rect 12930 7064 12931 7098
rect 12895 7030 12931 7064
rect 12895 6996 12896 7030
rect 12930 6996 12931 7030
rect 12895 6962 12931 6996
rect 12895 6928 12896 6962
rect 12930 6928 12931 6962
rect 12895 6894 12931 6928
rect 12895 6860 12896 6894
rect 12930 6860 12931 6894
rect 12895 6826 12931 6860
rect 12895 6792 12896 6826
rect 12930 6792 12931 6826
rect 12895 6758 12931 6792
rect 7669 6647 7703 6681
rect 7669 6579 7703 6613
rect 12895 6724 12896 6758
rect 12930 6724 12931 6758
rect 12895 6690 12931 6724
rect 12895 6656 12896 6690
rect 12930 6656 12931 6690
rect 12895 6622 12931 6656
rect 12895 6588 12896 6622
rect 12930 6588 12931 6622
rect 3929 6577 3964 6579
rect 3894 6545 3964 6577
rect 3998 6545 4032 6579
rect 4066 6545 4100 6579
rect 4134 6545 4168 6579
rect 4202 6545 4236 6579
rect 4270 6545 4304 6579
rect 4338 6545 4372 6579
rect 4406 6545 4440 6579
rect 4474 6545 4508 6579
rect 4542 6545 4576 6579
rect 4610 6545 4644 6579
rect 4678 6545 4712 6579
rect 4746 6545 4780 6579
rect 4814 6545 4848 6579
rect 4882 6545 4916 6579
rect 4950 6545 4984 6579
rect 5018 6545 5052 6579
rect 5086 6545 5120 6579
rect 5154 6545 5188 6579
rect 5222 6545 5256 6579
rect 5290 6545 5324 6579
rect 5358 6545 5392 6579
rect 5426 6545 5460 6579
rect 5494 6545 5528 6579
rect 5562 6545 5596 6579
rect 5630 6545 5664 6579
rect 5698 6545 5732 6579
rect 5766 6545 5800 6579
rect 5834 6545 5868 6579
rect 5902 6545 5936 6579
rect 5970 6545 6004 6579
rect 6038 6545 6072 6579
rect 6106 6545 6140 6579
rect 6174 6545 6208 6579
rect 6242 6545 6276 6579
rect 6310 6545 6344 6579
rect 6378 6545 6412 6579
rect 6446 6545 6480 6579
rect 6514 6545 6548 6579
rect 6582 6545 6616 6579
rect 6650 6545 6684 6579
rect 6718 6545 6752 6579
rect 6786 6545 6820 6579
rect 6854 6545 6888 6579
rect 6922 6545 6956 6579
rect 6990 6545 7024 6579
rect 7058 6545 7092 6579
rect 7126 6545 7160 6579
rect 7194 6545 7228 6579
rect 7262 6545 7296 6579
rect 7330 6545 7364 6579
rect 7398 6545 7432 6579
rect 7466 6545 7500 6579
rect 7534 6545 7568 6579
rect 7602 6545 7636 6579
rect 7670 6545 7704 6579
rect 7738 6545 7772 6579
rect 7806 6545 7840 6579
rect 7874 6545 7908 6579
rect 7942 6545 7976 6579
rect 8010 6545 8044 6579
rect 8078 6545 8112 6579
rect 8146 6545 8180 6579
rect 8214 6545 8248 6579
rect 8282 6545 8316 6579
rect 8350 6545 8384 6579
rect 8418 6545 8452 6579
rect 8486 6545 8520 6579
rect 8554 6545 8588 6579
rect 8622 6545 8656 6579
rect 8690 6545 8724 6579
rect 8758 6545 8792 6579
rect 8826 6545 8860 6579
rect 8894 6545 8928 6579
rect 8962 6545 8996 6579
rect 9030 6545 9064 6579
rect 9098 6545 9132 6579
rect 9166 6545 9200 6579
rect 9234 6545 9268 6579
rect 9302 6545 9336 6579
rect 9370 6545 9404 6579
rect 9438 6545 9472 6579
rect 9506 6545 9540 6579
rect 9574 6545 9608 6579
rect 9642 6545 9676 6579
rect 9710 6545 9744 6579
rect 9778 6545 9812 6579
rect 9846 6545 9880 6579
rect 9914 6545 9948 6579
rect 9982 6545 10016 6579
rect 10050 6545 10084 6579
rect 10118 6545 10152 6579
rect 10186 6545 10220 6579
rect 10254 6545 10288 6579
rect 10322 6545 10356 6579
rect 10390 6545 10424 6579
rect 10458 6545 10492 6579
rect 10526 6545 10560 6579
rect 10594 6545 10628 6579
rect 10662 6545 10696 6579
rect 10730 6545 10764 6579
rect 10798 6545 10832 6579
rect 10866 6545 10900 6579
rect 10934 6545 10968 6579
rect 11002 6545 11036 6579
rect 11070 6545 11104 6579
rect 11138 6545 11172 6579
rect 11206 6545 11240 6579
rect 11274 6545 11308 6579
rect 11342 6545 11376 6579
rect 11410 6545 11444 6579
rect 11478 6545 11512 6579
rect 11546 6545 11580 6579
rect 11614 6545 11648 6579
rect 11682 6545 11716 6579
rect 11750 6545 11784 6579
rect 11818 6545 11852 6579
rect 11886 6545 11920 6579
rect 11954 6545 12046 6579
rect 12895 6554 12931 6588
rect 3894 6543 3930 6545
rect 3894 6509 3895 6543
rect 3929 6509 3930 6543
rect 3894 6475 3930 6509
rect 3894 6441 3895 6475
rect 3929 6441 3930 6475
rect 3894 6407 3930 6441
rect 3894 6373 3895 6407
rect 3929 6373 3930 6407
rect 3894 6339 3930 6373
rect 12895 6520 12896 6554
rect 12930 6520 12931 6554
rect 12895 6486 12931 6520
rect 12895 6452 12896 6486
rect 12930 6452 12931 6486
rect 12895 6354 12931 6452
rect 3894 6305 3895 6339
rect 3929 6305 3930 6339
rect 3894 6271 3930 6305
rect 3894 6237 3895 6271
rect 3929 6237 3930 6271
rect 3894 6203 3930 6237
rect 3894 6169 3895 6203
rect 3929 6169 3930 6203
rect 3894 6135 3930 6169
rect 3894 6101 3895 6135
rect 3929 6101 3930 6135
rect 3894 6067 3930 6101
rect 3894 6033 3895 6067
rect 3929 6033 3930 6067
rect 3894 5999 3930 6033
rect 3894 5965 3895 5999
rect 3929 5965 3930 5999
rect 3894 5931 3930 5965
rect 3894 5897 3895 5931
rect 3929 5897 3930 5931
rect 3894 5863 3930 5897
rect 3894 5829 3895 5863
rect 3929 5829 3930 5863
rect 3894 5795 3930 5829
rect 3894 5761 3895 5795
rect 3929 5761 3930 5795
rect 3894 5727 3930 5761
rect 3894 5693 3895 5727
rect 3929 5693 3930 5727
rect 12194 6353 12931 6354
rect 12194 6320 12319 6353
rect 12194 6286 12195 6320
rect 12229 6319 12319 6320
rect 12353 6319 12387 6353
rect 12421 6319 12455 6353
rect 12489 6319 12523 6353
rect 12557 6319 12591 6353
rect 12625 6319 12659 6353
rect 12693 6319 12727 6353
rect 12761 6319 12795 6353
rect 12829 6319 12863 6353
rect 12897 6319 12931 6353
rect 12229 6318 12931 6319
rect 12229 6286 12230 6318
rect 12194 6252 12230 6286
rect 12194 6218 12195 6252
rect 12229 6218 12230 6252
rect 12194 6184 12230 6218
rect 12194 6150 12195 6184
rect 12229 6150 12230 6184
rect 12194 6116 12230 6150
rect 12194 6082 12195 6116
rect 12229 6082 12230 6116
rect 12194 6048 12230 6082
rect 12194 6014 12195 6048
rect 12229 6014 12230 6048
rect 12194 5980 12230 6014
rect 12194 5946 12195 5980
rect 12229 5946 12230 5980
rect 12194 5912 12230 5946
rect 12194 5878 12195 5912
rect 12229 5878 12230 5912
rect 12194 5844 12230 5878
rect 12194 5810 12195 5844
rect 12229 5810 12230 5844
rect 12194 5776 12230 5810
rect 12194 5742 12195 5776
rect 12229 5742 12230 5776
rect 3894 5659 3930 5693
rect 3894 5625 3895 5659
rect 3929 5625 3930 5659
rect 3894 5591 3930 5625
rect 3894 5557 3895 5591
rect 3929 5557 3930 5591
rect 3894 5523 3930 5557
rect 3894 5489 3895 5523
rect 3929 5489 3930 5523
rect 3894 5455 3930 5489
rect 3894 5421 3895 5455
rect 3929 5421 3930 5455
rect 3894 5387 3930 5421
rect 3894 5353 3895 5387
rect 3929 5353 3930 5387
rect 3894 5319 3930 5353
rect 3894 5285 3895 5319
rect 3929 5285 3930 5319
rect 3894 5251 3930 5285
rect 3894 5217 3895 5251
rect 3929 5217 3930 5251
rect 3894 5183 3930 5217
rect 3894 5149 3895 5183
rect 3929 5149 3930 5183
rect 11923 5678 11959 5712
rect 11923 5644 11924 5678
rect 11958 5644 11959 5678
rect 11923 5610 11959 5644
rect 11923 5576 11924 5610
rect 11958 5576 11959 5610
rect 11923 5542 11959 5576
rect 11923 5508 11924 5542
rect 11958 5508 11959 5542
rect 11923 5474 11959 5508
rect 11923 5440 11924 5474
rect 11958 5440 11959 5474
rect 11923 5406 11959 5440
rect 11923 5372 11924 5406
rect 11958 5372 11959 5406
rect 11923 5338 11959 5372
rect 11923 5304 11924 5338
rect 11958 5304 11959 5338
rect 11923 5270 11959 5304
rect 11923 5236 11924 5270
rect 11958 5236 11959 5270
rect 11923 5202 11959 5236
rect 3894 5115 3930 5149
rect 3894 5081 3895 5115
rect 3929 5081 3930 5115
rect 3894 5047 3930 5081
rect 3894 5013 3895 5047
rect 3929 5013 3930 5047
rect 3894 4979 3930 5013
rect 3894 4945 3895 4979
rect 3929 4945 3930 4979
rect 3894 4911 3930 4945
rect 11839 5166 11873 5182
rect 11839 5103 11873 5132
rect 11923 5168 11924 5202
rect 11958 5168 11959 5202
rect 11923 5134 11959 5168
rect 11839 5098 11841 5103
rect 11873 5064 11875 5069
rect 11839 5030 11875 5064
rect 11923 5100 11924 5134
rect 11958 5100 11959 5134
rect 11923 5066 11959 5100
rect 11923 5032 11924 5066
rect 11958 5032 11959 5066
rect 11923 4998 11959 5032
rect 11839 4962 11873 4996
rect 11839 4912 11873 4928
rect 11923 4964 11924 4998
rect 11958 4964 11959 4998
rect 11923 4930 11959 4964
rect 3894 4877 3895 4911
rect 3929 4877 3930 4911
rect 3894 4843 3930 4877
rect 3894 4809 3895 4843
rect 3929 4809 3930 4843
rect 3894 4775 3930 4809
rect 3894 4741 3895 4775
rect 3929 4741 3930 4775
rect 3894 4707 3930 4741
rect 3894 4673 3895 4707
rect 3929 4673 3930 4707
rect 3894 4639 3930 4673
rect 3894 4605 3895 4639
rect 3929 4605 3930 4639
rect 3894 4571 3930 4605
rect 3894 4537 3895 4571
rect 3929 4537 3930 4571
rect 3894 4503 3930 4537
rect 3894 4469 3895 4503
rect 3929 4469 3930 4503
rect 3894 4435 3930 4469
rect 3894 4401 3895 4435
rect 3929 4401 3930 4435
rect 3894 4367 3930 4401
rect 3894 4333 3895 4367
rect 3929 4333 3930 4367
rect 3894 4299 3930 4333
rect 3894 4265 3895 4299
rect 3929 4265 3930 4299
rect 3894 4231 3930 4265
rect 3894 4197 3895 4231
rect 3929 4197 3930 4231
rect 3894 4163 3930 4197
rect 3894 4129 3895 4163
rect 3929 4129 3930 4163
rect 3894 4095 3930 4129
rect 3894 4061 3895 4095
rect 3929 4061 3930 4095
rect 3894 4027 3930 4061
rect 3894 3993 3895 4027
rect 3929 3993 3930 4027
rect 3894 3959 3930 3993
rect 3894 3925 3895 3959
rect 3929 3925 3930 3959
rect 3894 3891 3930 3925
rect 3894 3857 3895 3891
rect 3929 3857 3930 3891
rect 3894 3823 3930 3857
rect 3894 3789 3895 3823
rect 3929 3789 3930 3823
rect 3894 3755 3930 3789
rect 3894 3721 3895 3755
rect 3929 3721 3930 3755
rect 3894 3687 3930 3721
rect 3894 3653 3895 3687
rect 3929 3653 3930 3687
rect 3894 3619 3930 3653
rect 3894 3585 3895 3619
rect 3929 3585 3930 3619
rect 3894 3551 3930 3585
rect 3894 3517 3895 3551
rect 3929 3517 3930 3551
rect 3894 3483 3930 3517
rect 3894 3449 3895 3483
rect 3929 3449 3930 3483
rect 3894 3415 3930 3449
rect 3894 3381 3895 3415
rect 3929 3381 3930 3415
rect 3894 3347 3930 3381
rect 3894 3313 3895 3347
rect 3929 3313 3930 3347
rect 3894 3279 3930 3313
rect 3894 3245 3895 3279
rect 3929 3245 3930 3279
rect 3894 3211 3930 3245
rect 3894 3177 3895 3211
rect 3929 3177 3930 3211
rect 11923 4896 11924 4930
rect 11958 4896 11959 4930
rect 11923 4862 11959 4896
rect 11923 4828 11924 4862
rect 11958 4828 11959 4862
rect 11923 4794 11959 4828
rect 11923 4760 11924 4794
rect 11958 4760 11959 4794
rect 11923 4726 11959 4760
rect 11923 4692 11924 4726
rect 11958 4692 11959 4726
rect 11923 4658 11959 4692
rect 11923 4624 11924 4658
rect 11958 4624 11959 4658
rect 11923 4590 11959 4624
rect 11923 4556 11924 4590
rect 11958 4556 11959 4590
rect 11923 4522 11959 4556
rect 11923 4488 11924 4522
rect 11958 4488 11959 4522
rect 11923 4454 11959 4488
rect 11923 4420 11924 4454
rect 11958 4420 11959 4454
rect 11923 4386 11959 4420
rect 11923 4352 11924 4386
rect 11958 4352 11959 4386
rect 11923 4318 11959 4352
rect 11923 4284 11924 4318
rect 11958 4284 11959 4318
rect 11923 4250 11959 4284
rect 11923 4216 11924 4250
rect 11958 4216 11959 4250
rect 11923 4182 11959 4216
rect 11923 4148 11924 4182
rect 11958 4148 11959 4182
rect 11923 4114 11959 4148
rect 11923 4080 11924 4114
rect 11958 4080 11959 4114
rect 11923 4046 11959 4080
rect 11923 4012 11924 4046
rect 11958 4012 11959 4046
rect 11923 3978 11959 4012
rect 11923 3944 11924 3978
rect 11958 3944 11959 3978
rect 11923 3910 11959 3944
rect 11923 3876 11924 3910
rect 11958 3876 11959 3910
rect 11923 3842 11959 3876
rect 11923 3808 11924 3842
rect 11958 3808 11959 3842
rect 11923 3774 11959 3808
rect 11923 3740 11924 3774
rect 11958 3740 11959 3774
rect 11923 3706 11959 3740
rect 11923 3672 11924 3706
rect 11958 3672 11959 3706
rect 11923 3638 11959 3672
rect 11923 3604 11924 3638
rect 11958 3604 11959 3638
rect 11923 3570 11959 3604
rect 11923 3536 11924 3570
rect 11958 3536 11959 3570
rect 11923 3502 11959 3536
rect 11923 3468 11924 3502
rect 11958 3468 11959 3502
rect 11923 3434 11959 3468
rect 11923 3400 11924 3434
rect 11958 3400 11959 3434
rect 11923 3366 11959 3400
rect 11923 3332 11924 3366
rect 11958 3332 11959 3366
rect 11923 3298 11959 3332
rect 11923 3264 11924 3298
rect 11958 3264 11959 3298
rect 11923 3230 11959 3264
rect 11923 3196 11924 3230
rect 11958 3196 11959 3230
rect 3894 3143 3930 3177
rect 3894 3109 3895 3143
rect 3929 3109 3930 3143
rect 3894 3075 3930 3109
rect 3894 3041 3895 3075
rect 3929 3041 3930 3075
rect 11839 3180 11873 3194
rect 11839 3110 11873 3144
rect 11839 3060 11873 3074
rect 11923 3162 11959 3196
rect 11923 3128 11924 3162
rect 11958 3128 11959 3162
rect 11923 3094 11959 3128
rect 11923 3060 11924 3094
rect 11958 3060 11959 3094
rect 3894 3007 3930 3041
rect 3894 2973 3895 3007
rect 3929 2973 3930 3007
rect 3894 2939 3930 2973
rect 3894 2905 3895 2939
rect 3929 2905 3930 2939
rect 11923 3026 11959 3060
rect 11923 2992 11924 3026
rect 11958 2992 11959 3026
rect 11923 2958 11959 2992
rect 3894 2871 3930 2905
rect 3894 2837 3895 2871
rect 3929 2837 3930 2871
rect 3894 2803 3930 2837
rect 11839 2924 11873 2938
rect 11839 2854 11873 2888
rect 11839 2804 11873 2818
rect 11923 2924 11924 2958
rect 11958 2924 11959 2958
rect 11923 2890 11959 2924
rect 11923 2856 11924 2890
rect 11958 2856 11959 2890
rect 11923 2822 11959 2856
rect 3894 2769 3895 2803
rect 3929 2769 3930 2803
rect 3894 2735 3930 2769
rect 3894 2701 3895 2735
rect 3929 2701 3930 2735
rect 3894 2667 3930 2701
rect 3894 2633 3895 2667
rect 3929 2633 3930 2667
rect 3894 2599 3930 2633
rect 3894 2565 3895 2599
rect 3929 2565 3930 2599
rect 3894 2531 3930 2565
rect 3894 2497 3895 2531
rect 3929 2497 3930 2531
rect 3894 2463 3930 2497
rect 3894 2429 3895 2463
rect 3929 2429 3930 2463
rect 3894 2395 3930 2429
rect 3894 2361 3895 2395
rect 3929 2361 3930 2395
rect 3894 2327 3930 2361
rect 3894 2293 3895 2327
rect 3929 2293 3930 2327
rect 3894 2259 3930 2293
rect 3894 2225 3895 2259
rect 3929 2225 3930 2259
rect 3894 2191 3930 2225
rect 3894 2157 3895 2191
rect 3929 2157 3930 2191
rect 3894 2123 3930 2157
rect 3894 2089 3895 2123
rect 3929 2089 3930 2123
rect 3894 2055 3930 2089
rect 3894 2021 3895 2055
rect 3929 2021 3930 2055
rect 3894 1987 3930 2021
rect 3894 1953 3895 1987
rect 3929 1953 3930 1987
rect 3894 1919 3930 1953
rect 11923 2788 11924 2822
rect 11958 2788 11959 2822
rect 11923 2754 11959 2788
rect 11923 2720 11924 2754
rect 11958 2720 11959 2754
rect 11923 2686 11959 2720
rect 11923 2652 11924 2686
rect 11958 2652 11959 2686
rect 11923 2618 11959 2652
rect 11923 2584 11924 2618
rect 11958 2584 11959 2618
rect 11923 2550 11959 2584
rect 11923 2516 11924 2550
rect 11958 2516 11959 2550
rect 11923 2482 11959 2516
rect 11923 2448 11924 2482
rect 11958 2448 11959 2482
rect 11923 2414 11959 2448
rect 11923 2380 11924 2414
rect 11958 2380 11959 2414
rect 11923 2346 11959 2380
rect 11923 2312 11924 2346
rect 11958 2312 11959 2346
rect 11923 2278 11959 2312
rect 11923 2244 11924 2278
rect 11958 2244 11959 2278
rect 11923 2210 11959 2244
rect 11923 2176 11924 2210
rect 11958 2176 11959 2210
rect 11923 2142 11959 2176
rect 11923 2108 11924 2142
rect 11958 2108 11959 2142
rect 11923 2074 11959 2108
rect 11923 2040 11924 2074
rect 11958 2040 11959 2074
rect 11923 1943 11959 2040
rect 12194 5708 12230 5742
rect 12194 5674 12195 5708
rect 12229 5674 12230 5708
rect 12194 5640 12230 5674
rect 12194 5606 12195 5640
rect 12229 5606 12230 5640
rect 12194 5572 12230 5606
rect 12194 5538 12195 5572
rect 12229 5538 12230 5572
rect 12194 5504 12230 5538
rect 12194 5470 12195 5504
rect 12229 5470 12230 5504
rect 12194 5436 12230 5470
rect 12194 5402 12195 5436
rect 12229 5402 12230 5436
rect 12194 5368 12230 5402
rect 12194 5334 12195 5368
rect 12229 5334 12230 5368
rect 12194 5300 12230 5334
rect 12194 5266 12195 5300
rect 12229 5266 12230 5300
rect 12194 5232 12230 5266
rect 12194 5198 12195 5232
rect 12229 5198 12230 5232
rect 12194 5164 12230 5198
rect 12194 5130 12195 5164
rect 12229 5130 12230 5164
rect 12194 5096 12230 5130
rect 12194 5062 12195 5096
rect 12229 5062 12230 5096
rect 12194 5028 12230 5062
rect 12194 4994 12195 5028
rect 12229 4994 12230 5028
rect 12194 4960 12230 4994
rect 12194 4926 12195 4960
rect 12229 4926 12230 4960
rect 12194 4892 12230 4926
rect 12194 4858 12195 4892
rect 12229 4858 12230 4892
rect 12194 4824 12230 4858
rect 12194 4790 12195 4824
rect 12229 4790 12230 4824
rect 12194 4756 12230 4790
rect 12194 4722 12195 4756
rect 12229 4722 12230 4756
rect 12194 4688 12230 4722
rect 12194 4654 12195 4688
rect 12229 4654 12230 4688
rect 12194 4620 12230 4654
rect 12194 4586 12195 4620
rect 12229 4586 12230 4620
rect 12194 4552 12230 4586
rect 12194 4518 12195 4552
rect 12229 4518 12230 4552
rect 12194 4484 12230 4518
rect 12194 4450 12195 4484
rect 12229 4450 12230 4484
rect 12194 4416 12230 4450
rect 12194 4382 12195 4416
rect 12229 4382 12230 4416
rect 12194 4348 12230 4382
rect 12194 4314 12195 4348
rect 12229 4314 12230 4348
rect 12194 4280 12230 4314
rect 12194 4246 12195 4280
rect 12229 4246 12230 4280
rect 12194 4212 12230 4246
rect 12194 4178 12195 4212
rect 12229 4178 12230 4212
rect 12194 4144 12230 4178
rect 12194 4110 12195 4144
rect 12229 4110 12230 4144
rect 12194 4076 12230 4110
rect 12194 4042 12195 4076
rect 12229 4042 12230 4076
rect 12194 4008 12230 4042
rect 12194 3974 12195 4008
rect 12229 3974 12230 4008
rect 12194 3940 12230 3974
rect 12194 3906 12195 3940
rect 12229 3906 12230 3940
rect 12194 3872 12230 3906
rect 12194 3838 12195 3872
rect 12229 3838 12230 3872
rect 12194 3804 12230 3838
rect 12194 3770 12195 3804
rect 12229 3770 12230 3804
rect 12194 3736 12230 3770
rect 12194 3702 12195 3736
rect 12229 3702 12230 3736
rect 12194 3668 12230 3702
rect 12194 3634 12195 3668
rect 12229 3634 12230 3668
rect 12194 3600 12230 3634
rect 12194 3566 12195 3600
rect 12229 3566 12230 3600
rect 12194 3532 12230 3566
rect 12194 3498 12195 3532
rect 12229 3498 12230 3532
rect 12194 3464 12230 3498
rect 12194 3430 12195 3464
rect 12229 3430 12230 3464
rect 12194 3396 12230 3430
rect 12194 3362 12195 3396
rect 12229 3362 12230 3396
rect 12194 3328 12230 3362
rect 12194 3294 12195 3328
rect 12229 3294 12230 3328
rect 12194 3260 12230 3294
rect 12194 3226 12195 3260
rect 12229 3226 12230 3260
rect 12194 3192 12230 3226
rect 12194 3158 12195 3192
rect 12229 3158 12230 3192
rect 12194 3124 12230 3158
rect 12194 3090 12195 3124
rect 12229 3090 12230 3124
rect 12194 3056 12230 3090
rect 12194 3022 12195 3056
rect 12229 3022 12230 3056
rect 12194 2988 12230 3022
rect 12194 2954 12195 2988
rect 12229 2954 12230 2988
rect 12194 2920 12230 2954
rect 12194 2886 12195 2920
rect 12229 2886 12230 2920
rect 12194 2852 12230 2886
rect 12194 2818 12195 2852
rect 12229 2818 12230 2852
rect 12194 2784 12230 2818
rect 12194 2750 12195 2784
rect 12229 2750 12230 2784
rect 12194 2716 12230 2750
rect 12194 2682 12195 2716
rect 12229 2682 12230 2716
rect 12194 2648 12230 2682
rect 12194 2614 12195 2648
rect 12229 2614 12230 2648
rect 12194 2580 12230 2614
rect 12194 2546 12195 2580
rect 12229 2546 12230 2580
rect 12194 2512 12230 2546
rect 12194 2478 12195 2512
rect 12229 2478 12230 2512
rect 12194 2444 12230 2478
rect 12194 2410 12195 2444
rect 12229 2410 12230 2444
rect 12194 2376 12230 2410
rect 12194 2342 12195 2376
rect 12229 2342 12230 2376
rect 12194 2308 12230 2342
rect 12194 2274 12195 2308
rect 12229 2274 12230 2308
rect 12194 2240 12230 2274
rect 12194 2206 12195 2240
rect 12229 2206 12230 2240
rect 12194 2172 12230 2206
rect 12194 2138 12195 2172
rect 12229 2138 12230 2172
rect 12194 2104 12230 2138
rect 12194 2070 12195 2104
rect 12229 2070 12230 2104
rect 12194 2036 12230 2070
rect 12194 2002 12195 2036
rect 12229 2002 12230 2036
rect 12194 1968 12230 2002
rect 3894 1885 3895 1919
rect 3929 1885 3930 1919
rect 3894 1851 3930 1885
rect 3894 1817 3895 1851
rect 3929 1817 3930 1851
rect 3894 1783 3930 1817
rect 3894 1749 3895 1783
rect 3929 1749 3930 1783
rect 3894 1715 3930 1749
rect 3894 1681 3895 1715
rect 3929 1681 3930 1715
rect 3894 1647 3930 1681
rect 3894 1613 3895 1647
rect 3929 1613 3930 1647
rect 3894 1579 3930 1613
rect 3894 1545 3895 1579
rect 3929 1545 3930 1579
rect 3894 1511 3930 1545
rect 3894 1477 3895 1511
rect 3929 1477 3930 1511
rect 3894 1443 3930 1477
rect 3894 1409 3895 1443
rect 3929 1409 3930 1443
rect 3894 1375 3930 1409
rect 3894 1341 3895 1375
rect 3929 1341 3930 1375
rect 3894 1307 3930 1341
rect 3894 1273 3895 1307
rect 3929 1273 3930 1307
rect 3894 1239 3930 1273
rect 3894 1205 3895 1239
rect 3929 1205 3930 1239
rect 3894 1171 3930 1205
rect 3894 1137 3895 1171
rect 3929 1137 3930 1171
rect 3894 1103 3930 1137
rect 3894 1069 3895 1103
rect 3929 1069 3930 1103
rect 3894 1035 3930 1069
rect 3894 1001 3895 1035
rect 3929 1001 3930 1035
rect 3894 967 3930 1001
rect 3894 933 3895 967
rect 3929 933 3930 967
rect 3894 899 3930 933
rect 3894 865 3895 899
rect 3929 867 3930 899
rect 12194 1934 12195 1968
rect 12229 1934 12230 1968
rect 12194 1900 12230 1934
rect 12194 1866 12195 1900
rect 12229 1866 12230 1900
rect 12194 1832 12230 1866
rect 12194 1798 12195 1832
rect 12229 1798 12230 1832
rect 12194 1764 12230 1798
rect 12194 1730 12195 1764
rect 12229 1730 12230 1764
rect 12194 1696 12230 1730
rect 12194 1662 12195 1696
rect 12229 1662 12230 1696
rect 12194 1628 12230 1662
rect 12194 1594 12195 1628
rect 12229 1594 12230 1628
rect 12194 1560 12230 1594
rect 12194 1526 12195 1560
rect 12229 1526 12230 1560
rect 12194 1492 12230 1526
rect 12194 1458 12195 1492
rect 12229 1458 12230 1492
rect 12194 1424 12230 1458
rect 12194 1390 12195 1424
rect 12229 1390 12230 1424
rect 12194 1356 12230 1390
rect 12194 1322 12195 1356
rect 12229 1322 12230 1356
rect 12194 1288 12230 1322
rect 12194 1254 12195 1288
rect 12229 1254 12230 1288
rect 12194 1220 12230 1254
rect 12194 1186 12195 1220
rect 12229 1186 12230 1220
rect 12194 1051 12230 1186
rect 12194 1017 12195 1051
rect 12229 1017 12230 1051
rect 12194 983 12230 1017
rect 12194 949 12195 983
rect 12229 949 12230 983
rect 12194 867 12230 949
rect 3929 866 12230 867
rect 3929 865 4002 866
rect 3894 832 4002 865
rect 4036 832 4070 866
rect 4104 832 4138 866
rect 4172 832 4206 866
rect 4240 832 4274 866
rect 4308 832 4342 866
rect 4376 832 4410 866
rect 4444 832 4478 866
rect 4512 832 4546 866
rect 4580 832 4614 866
rect 4648 832 4682 866
rect 4716 832 4750 866
rect 4784 832 4818 866
rect 4852 832 4886 866
rect 4920 832 4954 866
rect 4988 832 5022 866
rect 5056 832 5090 866
rect 5124 832 5158 866
rect 5192 832 5226 866
rect 5260 832 5294 866
rect 5328 832 5362 866
rect 5396 832 5430 866
rect 5464 832 5498 866
rect 5532 832 5566 866
rect 5600 832 5634 866
rect 5668 832 5702 866
rect 5736 832 5770 866
rect 5804 832 5838 866
rect 5872 832 5906 866
rect 5940 832 5974 866
rect 6008 832 6042 866
rect 6076 832 6110 866
rect 6144 832 6178 866
rect 6212 832 6246 866
rect 6280 832 6314 866
rect 6348 832 6382 866
rect 6416 832 6450 866
rect 6484 832 6518 866
rect 6552 832 6586 866
rect 6620 832 6654 866
rect 6688 832 6722 866
rect 6756 832 6790 866
rect 6824 832 6858 866
rect 6892 832 6926 866
rect 6960 832 6994 866
rect 7028 832 7062 866
rect 7096 832 7130 866
rect 7164 832 7198 866
rect 7232 832 7266 866
rect 7300 832 7334 866
rect 7368 832 7402 866
rect 7436 832 7470 866
rect 7504 832 7538 866
rect 7572 832 7606 866
rect 7640 832 7674 866
rect 7708 832 7742 866
rect 7776 832 7810 866
rect 7844 832 7878 866
rect 7912 832 7946 866
rect 7980 832 8014 866
rect 8048 832 8082 866
rect 8116 832 8150 866
rect 8184 832 8218 866
rect 8252 832 8286 866
rect 8320 832 8354 866
rect 8388 832 8422 866
rect 8456 832 8490 866
rect 8524 832 8558 866
rect 8592 832 8626 866
rect 8660 832 8694 866
rect 8728 832 8762 866
rect 8796 832 8830 866
rect 8864 832 8898 866
rect 8932 832 8966 866
rect 9000 832 9034 866
rect 9068 832 9102 866
rect 9136 832 9170 866
rect 9204 832 9238 866
rect 9272 832 9306 866
rect 9340 832 9374 866
rect 9408 832 9442 866
rect 9476 832 9510 866
rect 9544 832 9578 866
rect 9612 832 9646 866
rect 9680 832 9714 866
rect 9748 832 9782 866
rect 9816 832 9850 866
rect 9884 832 9918 866
rect 9952 832 9986 866
rect 10020 832 10054 866
rect 10088 832 10122 866
rect 10156 832 10190 866
rect 10224 832 10258 866
rect 10292 832 10326 866
rect 10360 832 10394 866
rect 10428 832 10462 866
rect 10496 832 10530 866
rect 10564 832 10598 866
rect 10632 832 10666 866
rect 10700 832 10734 866
rect 10768 832 10802 866
rect 10836 832 10870 866
rect 10904 832 10938 866
rect 10972 832 11006 866
rect 11040 832 11074 866
rect 11108 832 11142 866
rect 11176 832 11210 866
rect 11244 832 11278 866
rect 11312 832 11346 866
rect 11380 832 11414 866
rect 11448 832 11482 866
rect 11516 832 11550 866
rect 11584 832 11618 866
rect 11652 832 11686 866
rect 11720 832 11754 866
rect 11788 832 11822 866
rect 11856 832 11890 866
rect 11924 832 11958 866
rect 11992 832 12026 866
rect 12060 832 12094 866
rect 12128 832 12162 866
rect 12196 832 12230 866
rect 3894 831 12230 832
<< viali >>
rect 13250 14732 13278 14766
rect 13278 14732 13284 14766
rect 13324 14732 13346 14766
rect 13346 14732 13358 14766
rect 13398 14732 13414 14766
rect 13414 14732 13432 14766
rect 13472 14732 13482 14766
rect 13482 14732 13506 14766
rect 13546 14732 13550 14766
rect 13550 14732 13580 14766
rect 13620 14732 13652 14766
rect 13652 14732 13654 14766
rect 13694 14732 13720 14766
rect 13720 14732 13728 14766
rect 13768 14732 13788 14766
rect 13788 14732 13802 14766
rect 13842 14732 13856 14766
rect 13856 14732 13876 14766
rect 13916 14732 13924 14766
rect 13924 14732 13950 14766
rect 13990 14732 13992 14766
rect 13992 14732 14024 14766
rect 14064 14732 14094 14766
rect 14094 14732 14098 14766
rect 14138 14732 14162 14766
rect 14162 14732 14172 14766
rect 14212 14732 14230 14766
rect 14230 14732 14246 14766
rect 14286 14732 14298 14766
rect 14298 14732 14320 14766
rect 14360 14732 14366 14766
rect 14366 14732 14394 14766
rect 14434 14732 14468 14766
rect 14508 14732 14536 14766
rect 14536 14732 14542 14766
rect 14583 14732 14617 14766
rect 3071 14524 3079 14552
rect 3079 14524 3105 14552
rect 3071 14518 3105 14524
rect 3300 14498 3302 14532
rect 3302 14498 3334 14532
rect 3372 14498 3404 14532
rect 3404 14498 3406 14532
rect 3541 14498 3572 14532
rect 3572 14498 3575 14532
rect 3613 14498 3640 14532
rect 3640 14498 3647 14532
rect 3772 14498 3774 14532
rect 3774 14498 3806 14532
rect 3844 14498 3876 14532
rect 3876 14498 3878 14532
rect 4008 14498 4010 14532
rect 4010 14498 4042 14532
rect 4080 14498 4112 14532
rect 4112 14498 4114 14532
rect 3071 14456 3079 14476
rect 3079 14456 3105 14476
rect 3071 14442 3105 14456
rect 3071 14388 3079 14400
rect 3079 14388 3105 14400
rect 3071 14366 3105 14388
rect 3071 14320 3079 14324
rect 3079 14320 3105 14324
rect 3071 14290 3105 14320
rect 3071 14218 3105 14248
rect 3071 14214 3079 14218
rect 3079 14214 3105 14218
rect -253 14124 -219 14158
rect -253 14049 -219 14083
rect 259 14124 293 14158
rect 259 14052 293 14086
rect 771 14124 805 14158
rect 771 14052 805 14086
rect 1283 14124 1317 14158
rect 1283 14052 1317 14086
rect 1795 14124 1829 14158
rect 1795 14052 1829 14086
rect 3071 14150 3105 14172
rect 3071 14138 3079 14150
rect 3079 14138 3105 14150
rect 3071 14082 3105 14096
rect 3071 14062 3079 14082
rect 3079 14062 3105 14082
rect -253 13974 -219 14008
rect 3071 14014 3105 14020
rect -253 13898 -219 13932
rect 515 13954 549 13988
rect 515 13882 549 13916
rect 1539 13954 1573 13988
rect 1539 13878 1573 13912
rect 3 13784 37 13818
rect 3 13712 37 13746
rect 1027 13784 1061 13818
rect 1027 13712 1061 13746
rect 1539 13802 1573 13836
rect 1539 13726 1573 13760
rect 3071 13986 3079 14014
rect 3079 13986 3105 14014
rect 3071 13912 3079 13944
rect 3079 13912 3105 13944
rect 3071 13910 3105 13912
rect 3071 13844 3079 13868
rect 3079 13844 3105 13868
rect 3071 13834 3105 13844
rect 3071 13776 3079 13792
rect 3079 13776 3105 13792
rect 3071 13758 3105 13776
rect -56 13568 -54 13600
rect -54 13568 -22 13600
rect 19 13568 49 13600
rect 49 13568 53 13600
rect 94 13568 118 13600
rect 118 13568 128 13600
rect 169 13568 187 13600
rect 187 13568 203 13600
rect 244 13568 256 13600
rect 256 13568 278 13600
rect 319 13568 325 13600
rect 325 13568 353 13600
rect -56 13566 -22 13568
rect 19 13566 53 13568
rect 94 13566 128 13568
rect 169 13566 203 13568
rect 244 13566 278 13568
rect 319 13566 353 13568
rect 394 13566 428 13600
rect 469 13568 498 13600
rect 498 13568 503 13600
rect 544 13568 567 13600
rect 567 13568 578 13600
rect 619 13568 636 13600
rect 636 13568 653 13600
rect 694 13568 705 13600
rect 705 13568 728 13600
rect 769 13568 774 13600
rect 774 13568 803 13600
rect 843 13568 877 13600
rect 917 13568 946 13600
rect 946 13568 951 13600
rect 991 13568 1015 13600
rect 1015 13568 1025 13600
rect 1065 13568 1084 13600
rect 1084 13568 1099 13600
rect 1139 13568 1153 13600
rect 1153 13568 1173 13600
rect 1213 13568 1222 13600
rect 1222 13568 1247 13600
rect 1287 13568 1291 13600
rect 1291 13568 1321 13600
rect 1361 13568 1394 13600
rect 1394 13568 1395 13600
rect 3071 13708 3079 13716
rect 3079 13708 3105 13716
rect 3071 13682 3105 13708
rect 3071 13606 3105 13639
rect 3071 13605 3079 13606
rect 3079 13605 3105 13606
rect 469 13566 503 13568
rect 544 13566 578 13568
rect 619 13566 653 13568
rect 694 13566 728 13568
rect 769 13566 803 13568
rect 843 13566 877 13568
rect 917 13566 951 13568
rect 991 13566 1025 13568
rect 1065 13566 1099 13568
rect 1139 13566 1173 13568
rect 1213 13566 1247 13568
rect 1287 13566 1321 13568
rect 1361 13566 1395 13568
rect 3071 13538 3105 13562
rect 3071 13528 3079 13538
rect 3079 13528 3105 13538
rect 3071 13470 3105 13485
rect 3071 13451 3079 13470
rect 3079 13451 3105 13470
rect -492 13376 -462 13410
rect -462 13376 -458 13410
rect -416 13376 -394 13410
rect -394 13376 -382 13410
rect -340 13376 -326 13410
rect -326 13376 -306 13410
rect -264 13376 -258 13410
rect -258 13376 -230 13410
rect -564 13301 -530 13335
rect -564 13230 -530 13260
rect -564 13226 -530 13230
rect -564 13162 -530 13185
rect -564 13151 -530 13162
rect -564 13094 -530 13110
rect -564 13076 -530 13094
rect -564 13026 -530 13035
rect -564 13001 -530 13026
rect -564 12958 -530 12960
rect -564 12926 -530 12958
rect -564 12856 -530 12885
rect -564 12851 -530 12856
rect -564 12788 -530 12810
rect -564 12776 -530 12788
rect -564 12720 -530 12735
rect -564 12701 -530 12720
rect -564 12652 -530 12659
rect -564 12625 -530 12652
rect -564 12550 -530 12583
rect -564 12549 -530 12550
rect -564 12482 -530 12507
rect -564 12473 -530 12482
rect -564 12414 -530 12431
rect -564 12397 -530 12414
rect -564 12346 -530 12355
rect -564 12321 -530 12346
rect -564 12278 -530 12279
rect -564 12245 -530 12278
rect -564 12176 -530 12203
rect -564 12169 -530 12176
rect 5087 14376 5121 14386
rect 5087 14352 5121 14376
rect 14655 14664 14689 14666
rect 14655 14632 14689 14664
rect 13816 14549 13818 14583
rect 13818 14549 13850 14583
rect 13888 14549 13920 14583
rect 13920 14549 13922 14583
rect 14072 14549 14074 14583
rect 14074 14549 14106 14583
rect 14144 14549 14176 14583
rect 14176 14549 14178 14583
rect 14655 14562 14689 14565
rect 5087 14308 5121 14314
rect 5087 14280 5121 14308
rect 5087 14240 5121 14242
rect 5087 14208 5121 14240
rect 5087 14138 5121 14170
rect 5087 14136 5121 14138
rect 5087 14070 5121 14098
rect 5087 14064 5121 14070
rect 5087 14002 5121 14026
rect 5087 13992 5121 14002
rect 5087 13934 5121 13954
rect 5087 13920 5121 13934
rect 5087 13866 5121 13882
rect 5087 13848 5121 13866
rect 5087 13798 5121 13810
rect 5087 13776 5121 13798
rect 5087 13730 5121 13738
rect 5087 13704 5121 13730
rect 5087 13662 5121 13666
rect 5087 13632 5121 13662
rect 5087 13560 5121 13593
rect 5087 13559 5121 13560
rect 5087 13492 5121 13520
rect 5087 13486 5121 13492
rect 5087 13424 5121 13447
rect 5087 13413 5121 13424
rect 5087 13356 5121 13374
rect 5087 13340 5121 13356
rect 5087 13288 5121 13301
rect 5087 13267 5121 13288
rect 5087 13220 5121 13228
rect 5087 13194 5121 13220
rect 5087 13152 5121 13155
rect 5087 13121 5121 13152
rect 5087 13050 5121 13082
rect 5087 13048 5121 13050
rect 5087 12982 5121 13009
rect 5087 12975 5121 12982
rect 4501 12931 4503 12962
rect 4503 12931 4535 12962
rect 4573 12931 4605 12962
rect 4605 12931 4607 12962
rect 4757 12931 4759 12962
rect 4759 12931 4791 12962
rect 4829 12931 4861 12962
rect 4861 12931 4863 12962
rect 4501 12928 4535 12931
rect 4573 12928 4607 12931
rect 4757 12928 4791 12931
rect 4829 12928 4863 12931
rect 5087 12914 5121 12936
rect 5087 12902 5121 12914
rect 5087 12846 5121 12863
rect 5087 12829 5121 12846
rect 5087 12778 5121 12790
rect 5087 12756 5121 12778
rect 5087 12710 5121 12717
rect 5087 12683 5121 12710
rect 5087 12642 5121 12644
rect 5087 12610 5121 12642
rect 5087 12540 5121 12571
rect 5087 12537 5121 12540
rect 5087 12472 5121 12498
rect 5087 12464 5121 12472
rect 8715 14090 8743 14124
rect 8743 14090 8749 14124
rect 8787 14090 8819 14124
rect 8819 14090 8821 14124
rect 5740 13884 5774 13885
rect 5812 13884 5846 13885
rect 5740 13851 5756 13884
rect 5756 13851 5774 13884
rect 5812 13851 5832 13884
rect 5832 13851 5846 13884
rect 9019 13696 9053 13730
rect 9091 13696 9095 13730
rect 9095 13696 9125 13730
rect 11758 13572 11771 13606
rect 11771 13572 11792 13606
rect 11841 13572 11873 13606
rect 11873 13572 11875 13606
rect 11924 13572 11941 13606
rect 11941 13572 11958 13606
rect 12007 13572 12009 13606
rect 12009 13572 12041 13606
rect 12090 13572 12111 13606
rect 12111 13572 12124 13606
rect 12565 13572 12587 13606
rect 12587 13572 12599 13606
rect 12642 13572 12655 13606
rect 12655 13572 12676 13606
rect 12719 13572 12723 13606
rect 12723 13572 12753 13606
rect 11686 13504 11720 13533
rect 11686 13499 11720 13504
rect 11686 13436 11720 13460
rect 11686 13426 11720 13436
rect 12791 13499 12825 13533
rect 12791 13451 12825 13460
rect 12791 13426 12825 13451
rect 11686 13368 11720 13387
rect 11686 13353 11720 13368
rect 11686 13300 11720 13314
rect 11686 13280 11720 13300
rect 11686 13232 11720 13241
rect 11686 13207 11720 13232
rect 11686 13164 11720 13168
rect 11686 13134 11720 13164
rect 11686 13062 11720 13095
rect 11686 13061 11720 13062
rect 11686 12994 11720 13022
rect 11686 12988 11720 12994
rect 11686 12926 11720 12949
rect 11686 12915 11720 12926
rect 11686 12858 11720 12875
rect 11686 12841 11720 12858
rect 11686 12790 11720 12801
rect 11686 12767 11720 12790
rect 11686 12722 11720 12727
rect 11686 12693 11720 12722
rect 11686 12620 11720 12653
rect 11686 12619 11720 12620
rect 11686 12552 11720 12579
rect 11686 12545 11720 12552
rect 11686 12484 11720 12505
rect 11686 12471 11720 12484
rect 5087 12404 5121 12425
rect 5087 12391 5121 12404
rect 3300 12356 3302 12390
rect 3302 12356 3334 12390
rect 3372 12356 3404 12390
rect 3404 12356 3406 12390
rect 3536 12356 3538 12390
rect 3538 12356 3570 12390
rect 3608 12356 3640 12390
rect 3640 12356 3642 12390
rect 3772 12356 3774 12390
rect 3774 12356 3806 12390
rect 3844 12356 3876 12390
rect 3876 12356 3878 12390
rect 4008 12356 4010 12390
rect 4010 12356 4042 12390
rect 4080 12356 4112 12390
rect 4112 12356 4114 12390
rect -329 12008 -327 12042
rect -327 12008 -295 12042
rect -257 12008 -225 12042
rect -225 12008 -223 12042
rect -73 12008 -71 12042
rect -71 12008 -39 12042
rect -1 12008 31 12042
rect 31 12008 33 12042
rect 249 12008 251 12042
rect 251 12008 283 12042
rect 321 12008 353 12042
rect 353 12008 355 12042
rect 5087 12336 5121 12352
rect 5087 12318 5121 12336
rect 5087 12268 5121 12279
rect 5087 12245 5121 12268
rect 5087 12200 5121 12206
rect 5087 12172 5121 12200
rect 4462 11981 4464 12015
rect 4464 11981 4496 12015
rect 4534 11981 4566 12015
rect 4566 11981 4568 12015
rect 4718 11981 4720 12015
rect 4720 11981 4752 12015
rect 4790 11981 4822 12015
rect 4822 11981 4824 12015
rect 11686 12416 11720 12431
rect 11686 12397 11720 12416
rect 11686 12348 11720 12357
rect 11686 12323 11720 12348
rect 11686 12280 11720 12283
rect 11686 12249 11720 12280
rect 11880 13384 11914 13418
rect 11952 13384 11986 13418
rect 12024 13384 12056 13418
rect 12056 13384 12058 13418
rect 12522 13384 12532 13418
rect 12532 13384 12556 13418
rect 12594 13384 12628 13418
rect 11874 13316 11908 13319
rect 11874 13285 11908 13316
rect 12600 13334 12634 13340
rect 12600 13306 12634 13334
rect 11874 13214 11908 13247
rect 11874 13213 11908 13214
rect 11874 13146 11908 13175
rect 11874 13141 11908 13146
rect 11874 13078 11908 13103
rect 11874 13069 11908 13078
rect 11874 13010 11908 13031
rect 11874 12997 11908 13010
rect 11874 12942 11908 12959
rect 11874 12925 11908 12942
rect 11874 12874 11908 12887
rect 11874 12853 11908 12874
rect 11874 12806 11908 12815
rect 11874 12781 11908 12806
rect 11874 12738 11908 12743
rect 11874 12709 11908 12738
rect 11874 12670 11908 12671
rect 11874 12637 11908 12670
rect 11874 12568 11908 12599
rect 11874 12565 11908 12568
rect 11874 12500 11908 12527
rect 11874 12493 11908 12500
rect 12226 13213 12260 13247
rect 12226 13136 12260 13170
rect 12226 13059 12260 13093
rect 12226 12982 12260 13016
rect 12226 12905 12260 12939
rect 12226 12828 12260 12862
rect 12226 12751 12260 12785
rect 12226 12674 12260 12708
rect 12226 12597 12260 12631
rect 12226 12520 12260 12554
rect 12600 13266 12634 13268
rect 12600 13234 12634 13266
rect 12600 13164 12634 13196
rect 12600 13162 12634 13164
rect 12600 13096 12634 13124
rect 12600 13090 12634 13096
rect 12600 13028 12634 13052
rect 12600 13018 12634 13028
rect 12600 12960 12634 12980
rect 12600 12946 12634 12960
rect 12600 12892 12634 12908
rect 12600 12874 12634 12892
rect 12600 12824 12634 12836
rect 12600 12802 12634 12824
rect 12600 12756 12634 12764
rect 12600 12730 12634 12756
rect 12600 12688 12634 12692
rect 12600 12658 12634 12688
rect 12600 12586 12634 12620
rect 11874 12432 11908 12455
rect 11874 12421 11908 12432
rect 11874 12364 11908 12383
rect 11874 12349 11908 12364
rect 11874 12296 11908 12311
rect 11874 12277 11908 12296
rect 12600 12518 12634 12548
rect 12600 12514 12634 12518
rect 12600 12450 12634 12476
rect 12600 12442 12634 12450
rect 12600 12382 12634 12404
rect 12600 12370 12634 12382
rect 12600 12314 12634 12332
rect 12600 12298 12634 12314
rect 12600 12246 12634 12260
rect 12600 12226 12634 12246
rect 12062 12161 12064 12193
rect 12064 12161 12096 12193
rect 12134 12161 12166 12193
rect 12166 12161 12168 12193
rect 12318 12161 12320 12193
rect 12320 12161 12352 12193
rect 12390 12161 12422 12193
rect 12422 12161 12424 12193
rect 12062 12159 12096 12161
rect 12134 12159 12168 12161
rect 12318 12159 12352 12161
rect 12390 12159 12424 12161
rect 12600 12178 12634 12188
rect 12600 12154 12634 12178
rect 11886 12076 11920 12110
rect 11958 12076 11976 12110
rect 11976 12076 11992 12110
rect 12030 12076 12044 12110
rect 12044 12076 12064 12110
rect 12102 12076 12112 12110
rect 12112 12076 12136 12110
rect 12174 12076 12180 12110
rect 12180 12076 12208 12110
rect 12246 12076 12248 12110
rect 12248 12076 12280 12110
rect 12318 12076 12350 12110
rect 12350 12076 12352 12110
rect 12390 12076 12418 12110
rect 12418 12076 12424 12110
rect 12462 12076 12486 12110
rect 12486 12076 12496 12110
rect 12600 12082 12634 12116
rect 12791 13383 12825 13387
rect 12791 13353 12825 13383
rect 12791 13281 12825 13314
rect 12791 13280 12825 13281
rect 12791 13213 12825 13241
rect 12791 13207 12825 13213
rect 12791 13145 12825 13168
rect 12791 13134 12825 13145
rect 12791 13077 12825 13095
rect 12791 13061 12825 13077
rect 12791 13009 12825 13022
rect 12791 12988 12825 13009
rect 12791 12941 12825 12949
rect 12791 12915 12825 12941
rect 12791 12873 12825 12876
rect 12791 12842 12825 12873
rect 12791 12771 12825 12803
rect 12791 12769 12825 12771
rect 12791 12703 12825 12730
rect 12791 12696 12825 12703
rect 12791 12635 12825 12657
rect 12791 12623 12825 12635
rect 12791 12567 12825 12583
rect 12791 12549 12825 12567
rect 12791 12499 12825 12509
rect 12791 12475 12825 12499
rect 12791 12431 12825 12435
rect 12791 12401 12825 12431
rect 12791 12329 12825 12361
rect 12791 12327 12825 12329
rect 12791 12261 12825 12287
rect 12791 12253 12825 12261
rect 12791 12193 12825 12213
rect 12791 12179 12825 12193
rect 12791 12125 12825 12139
rect 12791 12105 12825 12125
rect 14655 14531 14689 14562
rect 14655 14460 14689 14484
rect 14655 14450 14689 14460
rect 14655 14392 14689 14412
rect 14655 14378 14689 14392
rect 14655 14324 14689 14340
rect 14655 14306 14689 14324
rect 14655 14256 14689 14268
rect 14655 14234 14689 14256
rect 14655 14188 14689 14196
rect 14655 14162 14689 14188
rect 14655 14120 14689 14124
rect 14655 14090 14689 14120
rect 14655 14018 14689 14052
rect 14655 13950 14689 13980
rect 14655 13946 14689 13950
rect 14655 13882 14689 13908
rect 14655 13874 14689 13882
rect 14655 13814 14689 13836
rect 14655 13802 14689 13814
rect 14655 13746 14689 13764
rect 14655 13730 14689 13746
rect 14655 13678 14689 13692
rect 14655 13658 14689 13678
rect 14655 13610 14689 13620
rect 14655 13586 14689 13610
rect 14655 13542 14689 13548
rect 14655 13514 14689 13542
rect 14655 13474 14689 13476
rect 14655 13442 14689 13474
rect 14655 13372 14689 13404
rect 14655 13370 14689 13372
rect 13556 13335 13558 13369
rect 13558 13335 13590 13369
rect 13628 13335 13660 13369
rect 13660 13335 13662 13369
rect 13812 13335 13814 13369
rect 13814 13335 13846 13369
rect 13884 13335 13916 13369
rect 13916 13335 13918 13369
rect 14068 13335 14070 13369
rect 14070 13335 14102 13369
rect 14140 13335 14172 13369
rect 14172 13335 14174 13369
rect 14324 13335 14326 13369
rect 14326 13335 14358 13369
rect 14396 13335 14428 13369
rect 14428 13335 14430 13369
rect 14655 13304 14689 13332
rect 14655 13298 14689 13304
rect 14655 13236 14689 13260
rect 14655 13226 14689 13236
rect 14655 13168 14689 13188
rect 14655 13154 14689 13168
rect 14655 13100 14689 13116
rect 14655 13082 14689 13100
rect 14655 13032 14689 13044
rect 14655 13010 14689 13032
rect 14655 12964 14689 12972
rect 14655 12938 14689 12964
rect 14655 12896 14689 12900
rect 14655 12866 14689 12896
rect 14655 12794 14689 12827
rect 14655 12793 14689 12794
rect 14655 12726 14689 12754
rect 14655 12720 14689 12726
rect 14655 12658 14689 12681
rect 14655 12647 14689 12658
rect 14655 12590 14689 12608
rect 14655 12574 14689 12590
rect 14655 12522 14689 12535
rect 14655 12501 14689 12522
rect 14655 12454 14689 12462
rect 14655 12428 14689 12454
rect 14655 12386 14689 12389
rect 14655 12355 14689 12386
rect 14655 12284 14689 12316
rect 14655 12282 14689 12284
rect 14655 12216 14689 12243
rect 14655 12209 14689 12216
rect 13816 12134 13818 12168
rect 13818 12134 13850 12168
rect 13888 12134 13920 12168
rect 13920 12134 13922 12168
rect 14072 12134 14074 12168
rect 14074 12134 14106 12168
rect 14144 12134 14176 12168
rect 14176 12134 14178 12168
rect 14655 12148 14689 12170
rect 14655 12136 14689 12148
rect 14655 12063 14689 12097
rect 3901 7540 3928 7574
rect 3928 7540 3935 7574
rect 3974 7540 3996 7574
rect 3996 7540 4008 7574
rect 4047 7540 4064 7574
rect 4064 7540 4081 7574
rect 4120 7540 4132 7574
rect 4132 7540 4154 7574
rect 4193 7540 4200 7574
rect 4200 7540 4227 7574
rect 4266 7540 4268 7574
rect 4268 7540 4300 7574
rect 4339 7540 4370 7574
rect 4370 7540 4373 7574
rect 4412 7540 4438 7574
rect 4438 7540 4446 7574
rect 4485 7540 4506 7574
rect 4506 7540 4519 7574
rect 4558 7540 4574 7574
rect 4574 7540 4592 7574
rect 4631 7540 4642 7574
rect 4642 7540 4665 7574
rect 4704 7540 4710 7574
rect 4710 7540 4738 7574
rect 4777 7540 4778 7574
rect 4778 7540 4811 7574
rect 4850 7540 4880 7574
rect 4880 7540 4884 7574
rect 4923 7540 4948 7574
rect 4948 7540 4957 7574
rect 4996 7540 5016 7574
rect 5016 7540 5030 7574
rect 5069 7540 5084 7574
rect 5084 7540 5103 7574
rect 5142 7540 5152 7574
rect 5152 7540 5176 7574
rect 5215 7540 5220 7574
rect 5220 7540 5249 7574
rect 5288 7540 5322 7574
rect 5361 7540 5390 7574
rect 5390 7540 5395 7574
rect 5434 7540 5458 7574
rect 5458 7540 5468 7574
rect 5507 7540 5526 7574
rect 5526 7540 5541 7574
rect 5580 7540 5594 7574
rect 5594 7540 5614 7574
rect 5653 7540 5662 7574
rect 5662 7540 5687 7574
rect 5726 7540 5730 7574
rect 5730 7540 5760 7574
rect 5799 7540 5832 7574
rect 5832 7540 5833 7574
rect 5872 7540 5900 7574
rect 5900 7540 5906 7574
rect 5945 7540 5968 7574
rect 5968 7540 5979 7574
rect 6018 7540 6036 7574
rect 6036 7540 6052 7574
rect 6091 7540 6104 7574
rect 6104 7540 6125 7574
rect 6164 7540 6172 7574
rect 6172 7540 6198 7574
rect 6237 7540 6240 7574
rect 6240 7540 6271 7574
rect 6310 7540 6342 7574
rect 6342 7540 6344 7574
rect 6383 7540 6410 7574
rect 6410 7540 6417 7574
rect 6456 7540 6478 7574
rect 6478 7540 6490 7574
rect 6530 7540 6546 7574
rect 6546 7540 6564 7574
rect 6604 7540 6614 7574
rect 6614 7540 6638 7574
rect 6678 7540 6682 7574
rect 6682 7540 6712 7574
rect 6752 7540 6784 7574
rect 6784 7540 6786 7574
rect 6826 7540 6852 7574
rect 6852 7540 6860 7574
rect 6900 7540 6920 7574
rect 6920 7540 6934 7574
rect 6974 7540 6988 7574
rect 6988 7540 7008 7574
rect 7048 7540 7056 7574
rect 7056 7540 7082 7574
rect 7122 7540 7124 7574
rect 7124 7540 7156 7574
rect 7196 7540 7226 7574
rect 7226 7540 7230 7574
rect 7270 7540 7294 7574
rect 7294 7540 7304 7574
rect 7344 7540 7362 7574
rect 7362 7540 7378 7574
rect 7418 7540 7430 7574
rect 7430 7540 7452 7574
rect 7492 7540 7498 7574
rect 7498 7540 7526 7574
rect 7566 7540 7600 7574
rect 7640 7540 7668 7574
rect 7668 7540 7674 7574
rect 7714 7540 7736 7574
rect 7736 7540 7748 7574
rect 3895 7461 3929 7483
rect 3895 7449 3929 7461
rect 3895 7393 3929 7401
rect 3895 7367 3929 7393
rect 3895 7291 3929 7319
rect 3895 7285 3929 7291
rect 3895 7223 3929 7237
rect 3895 7203 3929 7223
rect 3895 7121 3929 7155
rect 3895 7053 3929 7074
rect 3895 7040 3929 7053
rect 3895 6985 3929 6993
rect 3895 6959 3929 6985
rect 4180 7352 4214 7386
rect 4271 7352 4282 7386
rect 4282 7352 4305 7386
rect 4361 7352 4384 7386
rect 4384 7352 4395 7386
rect 4108 7284 4142 7302
rect 4108 7268 4142 7284
rect 4108 7216 4142 7218
rect 4108 7184 4142 7216
rect 4108 7114 4142 7133
rect 4108 7099 4142 7114
rect 4482 7177 4516 7182
rect 4482 7148 4516 7177
rect 4482 7109 4516 7110
rect 4482 7076 4516 7109
rect 4108 7046 4142 7048
rect 4108 7014 4142 7046
rect 4108 6944 4142 6963
rect 4108 6929 4142 6944
rect 4181 6857 4210 6891
rect 4210 6857 4215 6891
rect 4254 6857 4278 6891
rect 4278 6857 4288 6891
rect 4327 6857 4346 6891
rect 4346 6857 4361 6891
rect 4400 6857 4414 6891
rect 4414 6857 4434 6891
rect 4473 6857 4482 6891
rect 4482 6857 4507 6891
rect 4546 6857 4580 6891
rect 5005 7352 5039 7386
rect 5083 7352 5094 7386
rect 5094 7352 5117 7386
rect 5161 7352 5162 7386
rect 5162 7352 5195 7386
rect 5239 7352 5264 7386
rect 5264 7352 5273 7386
rect 5317 7352 5332 7386
rect 5332 7352 5351 7386
rect 5396 7352 5400 7386
rect 5400 7352 5430 7386
rect 5468 7299 5502 7301
rect 5468 7267 5502 7299
rect 5468 7197 5502 7215
rect 5365 7177 5399 7182
rect 5365 7148 5399 7177
rect 5365 7109 5399 7110
rect 5365 7076 5399 7109
rect 5468 7181 5502 7197
rect 5468 7095 5502 7129
rect 5000 6857 5034 6891
rect 5078 6857 5090 6891
rect 5090 6857 5112 6891
rect 5156 6857 5158 6891
rect 5158 6857 5190 6891
rect 5234 6857 5260 6891
rect 5260 6857 5268 6891
rect 5312 6857 5328 6891
rect 5328 6857 5346 6891
rect 5390 6857 5424 6891
rect 5468 6878 5502 6912
rect 5890 7352 5922 7386
rect 5922 7352 5924 7386
rect 5963 7352 5990 7386
rect 5990 7352 5997 7386
rect 6036 7352 6058 7386
rect 6058 7352 6070 7386
rect 6110 7352 6126 7386
rect 6126 7352 6144 7386
rect 6184 7352 6194 7386
rect 6194 7352 6218 7386
rect 6258 7352 6262 7386
rect 6262 7352 6292 7386
rect 6330 7299 6364 7312
rect 6330 7278 6364 7299
rect 6330 7231 6364 7238
rect 6330 7204 6364 7231
rect 6223 7177 6257 7182
rect 6223 7148 6257 7177
rect 6223 7109 6257 7110
rect 6223 7076 6257 7109
rect 6330 7129 6364 7163
rect 5913 6857 5918 6891
rect 5918 6857 5947 6891
rect 5995 6857 6020 6891
rect 6020 6857 6029 6891
rect 6072 6857 6088 6891
rect 6088 6857 6106 6891
rect 6149 6857 6156 6891
rect 6156 6857 6183 6891
rect 6221 6857 6224 6891
rect 6224 6857 6255 6891
rect 6340 6857 6374 6891
rect 7008 7352 7042 7386
rect 7090 7352 7120 7386
rect 7120 7352 7124 7386
rect 7172 7352 7188 7386
rect 7188 7352 7206 7386
rect 7254 7352 7256 7386
rect 7256 7352 7288 7386
rect 7460 7299 7494 7302
rect 7460 7268 7494 7299
rect 7460 7197 7494 7218
rect 7359 7177 7393 7179
rect 7359 7145 7393 7177
rect 7359 7075 7393 7107
rect 7359 7073 7393 7075
rect 7460 7184 7494 7197
rect 7460 7129 7494 7133
rect 7460 7099 7494 7129
rect 6980 6978 7014 6994
rect 6980 6960 7014 6978
rect 7460 7027 7494 7048
rect 7460 7014 7494 7027
rect 7460 6959 7494 6963
rect 7460 6929 7494 6959
rect 7052 6857 7082 6891
rect 7082 6857 7086 6891
rect 7134 6857 7150 6891
rect 7150 6857 7168 6891
rect 7216 6857 7218 6891
rect 7218 6857 7250 6891
rect 7298 6857 7320 6891
rect 7320 6857 7332 6891
rect 7379 6857 7413 6891
rect 8221 7997 8233 8031
rect 8233 7997 8255 8031
rect 8294 7997 8301 8031
rect 8301 7997 8328 8031
rect 8367 7997 8369 8031
rect 8369 7997 8401 8031
rect 8440 7997 8471 8031
rect 8471 7997 8474 8031
rect 8513 7997 8539 8031
rect 8539 7997 8547 8031
rect 8586 7997 8607 8031
rect 8607 7997 8620 8031
rect 8659 7997 8675 8031
rect 8675 7997 8693 8031
rect 8732 7997 8743 8031
rect 8743 7997 8766 8031
rect 8805 7997 8811 8031
rect 8811 7997 8839 8031
rect 8878 7997 8879 8031
rect 8879 7997 8912 8031
rect 8951 7997 8981 8031
rect 8981 7997 8985 8031
rect 9024 7997 9049 8031
rect 9049 7997 9058 8031
rect 9097 7997 9117 8031
rect 9117 7997 9131 8031
rect 9170 7997 9185 8031
rect 9185 7997 9204 8031
rect 9243 7997 9253 8031
rect 9253 7997 9277 8031
rect 9316 7997 9321 8031
rect 9321 7997 9350 8031
rect 9389 7997 9423 8031
rect 9462 7997 9491 8031
rect 9491 7997 9496 8031
rect 9535 7997 9559 8031
rect 9559 7997 9569 8031
rect 9608 7997 9627 8031
rect 9627 7997 9642 8031
rect 9681 7997 9695 8031
rect 9695 7997 9715 8031
rect 9754 7997 9763 8031
rect 9763 7997 9788 8031
rect 9827 7997 9831 8031
rect 9831 7997 9861 8031
rect 9900 7997 9933 8031
rect 9933 7997 9934 8031
rect 9973 7997 10001 8031
rect 10001 7997 10007 8031
rect 10046 7997 10069 8031
rect 10069 7997 10080 8031
rect 10119 7997 10137 8031
rect 10137 7997 10153 8031
rect 10192 7997 10205 8031
rect 10205 7997 10226 8031
rect 10265 7997 10273 8031
rect 10273 7997 10299 8031
rect 10338 7997 10341 8031
rect 10341 7997 10372 8031
rect 10411 7997 10443 8031
rect 10443 7997 10445 8031
rect 10484 7997 10511 8031
rect 10511 7997 10518 8031
rect 10557 7997 10579 8031
rect 10579 7997 10591 8031
rect 10630 7997 10647 8031
rect 10647 7997 10664 8031
rect 10703 7997 10715 8031
rect 10715 7997 10737 8031
rect 10776 7997 10783 8031
rect 10783 7997 10810 8031
rect 10849 7997 10851 8031
rect 10851 7997 10883 8031
rect 10922 7997 10953 8031
rect 10953 7997 10956 8031
rect 10995 7997 11021 8031
rect 11021 7997 11029 8031
rect 11068 7997 11089 8031
rect 11089 7997 11102 8031
rect 11141 7997 11157 8031
rect 11157 7997 11175 8031
rect 11214 7997 11225 8031
rect 11225 7997 11248 8031
rect 11286 7997 11293 8031
rect 11293 7997 11320 8031
rect 11358 7997 11361 8031
rect 11361 7997 11392 8031
rect 11430 7997 11463 8031
rect 11463 7997 11464 8031
rect 11502 7997 11531 8031
rect 11531 7997 11536 8031
rect 11574 7997 11599 8031
rect 11599 7997 11608 8031
rect 11646 7997 11667 8031
rect 11667 7997 11680 8031
rect 11718 7997 11735 8031
rect 11735 7997 11752 8031
rect 11790 7997 11803 8031
rect 11803 7997 11824 8031
rect 11862 7997 11871 8031
rect 11871 7997 11896 8031
rect 11934 7997 11939 8031
rect 11939 7997 11968 8031
rect 12006 7997 12007 8031
rect 12007 7997 12040 8031
rect 12078 7997 12109 8031
rect 12109 7997 12112 8031
rect 12150 7997 12177 8031
rect 12177 7997 12184 8031
rect 12222 7997 12245 8031
rect 12245 7997 12256 8031
rect 12294 7997 12313 8031
rect 12313 7997 12328 8031
rect 8105 7804 8139 7806
rect 8105 7772 8139 7804
rect 8105 7702 8139 7734
rect 8105 7700 8139 7702
rect 10247 7804 10281 7806
rect 10247 7772 10281 7804
rect 10247 7702 10281 7734
rect 10247 7700 10281 7702
rect 10423 7804 10457 7806
rect 10423 7772 10457 7804
rect 10423 7702 10457 7734
rect 10423 7700 10457 7702
rect 12565 7804 12599 7806
rect 12565 7772 12599 7804
rect 12565 7702 12599 7734
rect 12565 7700 12599 7702
rect 8105 7568 8139 7570
rect 8105 7536 8139 7568
rect 8105 7466 8139 7498
rect 8105 7464 8139 7466
rect 10247 7568 10281 7570
rect 10247 7536 10281 7568
rect 10247 7466 10281 7498
rect 10247 7464 10281 7466
rect 10423 7568 10457 7570
rect 10423 7536 10457 7568
rect 10423 7466 10457 7498
rect 10423 7464 10457 7466
rect 12565 7568 12599 7570
rect 12565 7536 12599 7568
rect 12565 7466 12599 7498
rect 12565 7464 12599 7466
rect 8105 7332 8139 7338
rect 8105 7304 8139 7332
rect 8105 7264 8139 7266
rect 8105 7232 8139 7264
rect 10247 7332 10281 7334
rect 10247 7300 10281 7332
rect 10247 7230 10281 7262
rect 10247 7228 10281 7230
rect 10423 7332 10457 7334
rect 10423 7300 10457 7332
rect 10423 7230 10457 7262
rect 10423 7228 10457 7230
rect 12565 7332 12599 7334
rect 12565 7300 12599 7332
rect 12565 7230 12599 7262
rect 12565 7228 12599 7230
rect 8105 7096 8139 7098
rect 8105 7064 8139 7096
rect 8105 6994 8139 7026
rect 8105 6992 8139 6994
rect 10247 7096 10281 7098
rect 10247 7064 10281 7096
rect 10247 6994 10281 7026
rect 10247 6992 10281 6994
rect 10423 7096 10457 7098
rect 10423 7064 10457 7096
rect 10423 6994 10457 7026
rect 10423 6992 10457 6994
rect 12565 7096 12599 7098
rect 12565 7064 12599 7096
rect 12565 6994 12599 7026
rect 12565 6992 12599 6994
rect 11841 5098 11875 5103
rect 11841 5069 11873 5098
rect 11873 5069 11875 5098
rect 11841 4996 11873 5030
rect 11873 4996 11875 5030
rect 11839 3178 11873 3180
rect 11839 3146 11873 3178
rect 11839 3076 11873 3108
rect 11839 3074 11873 3076
rect 11839 2922 11873 2924
rect 11839 2890 11873 2922
rect 11839 2820 11873 2852
rect 11839 2818 11873 2820
<< metal1 >>
tri 13889 14849 13897 14857 se
rect 13897 14849 13903 14857
tri 7821 14825 7829 14833 se
rect 7829 14827 7881 14833
tri 1773 14767 1831 14825 se
rect 1831 14785 7829 14825
tri 1831 14767 1849 14785 nw
tri 7802 14767 7820 14785 ne
rect 7820 14775 7829 14785
rect 7820 14767 7881 14775
tri 1772 14766 1773 14767 se
rect 1773 14766 1830 14767
tri 1830 14766 1831 14767 nw
tri 7820 14766 7821 14767 ne
rect 7821 14766 7881 14767
tri 1756 14750 1772 14766 se
rect 1772 14750 1814 14766
tri 1814 14750 1830 14766 nw
tri 7821 14758 7829 14766 ne
rect 7829 14763 7881 14766
tri 1751 14745 1756 14750 se
rect 1756 14745 1809 14750
tri 1809 14745 1814 14750 nw
tri 7662 14745 7667 14750 se
rect 7667 14745 7673 14750
tri 1738 14732 1751 14745 se
rect 1751 14732 1796 14745
tri 1796 14732 1809 14745 nw
tri 1854 14732 1867 14745 se
rect 1867 14732 7673 14745
tri 1715 14709 1738 14732 se
rect 1738 14709 1773 14732
tri 1773 14709 1796 14732 nw
tri 1831 14709 1854 14732 se
rect 1854 14709 7673 14732
tri 1714 14708 1715 14709 se
rect 1715 14708 1772 14709
tri 1772 14708 1773 14709 nw
tri 1830 14708 1831 14709 se
rect 1831 14708 7673 14709
tri 1699 14693 1714 14708 se
rect 1714 14693 1757 14708
tri 1757 14693 1772 14708 nw
tri 1815 14693 1830 14708 se
rect 1830 14705 7673 14708
rect 1830 14693 1873 14705
tri 1873 14693 1885 14705 nw
tri 7660 14698 7667 14705 ne
rect 7667 14698 7673 14705
rect 7725 14698 7737 14750
rect 7789 14698 7795 14750
rect 7829 14705 7881 14711
rect 12750 14805 13903 14849
rect 13955 14805 13967 14857
rect 14019 14805 14025 14857
rect 12750 14772 12795 14805
tri 12795 14772 12828 14805 nw
tri 1693 14687 1699 14693 se
rect 1699 14687 1751 14693
tri 1751 14687 1757 14693 nw
tri 1809 14687 1815 14693 se
rect 1815 14687 1867 14693
tri 1867 14687 1873 14693 nw
tri 12744 14687 12750 14693 se
rect 12750 14687 12794 14772
tri 12794 14771 12795 14772 nw
rect 13170 14766 13440 14775
rect 13492 14766 13504 14775
rect 13556 14766 14695 14775
rect 13170 14732 13250 14766
rect 13284 14732 13324 14766
rect 13358 14732 13398 14766
rect 13432 14732 13440 14766
rect 13580 14732 13620 14766
rect 13654 14732 13694 14766
rect 13728 14732 13768 14766
rect 13802 14732 13842 14766
rect 13876 14732 13916 14766
rect 13950 14732 13990 14766
rect 14024 14732 14064 14766
rect 14098 14732 14138 14766
rect 14172 14732 14212 14766
rect 14246 14732 14286 14766
rect 14320 14732 14360 14766
rect 14394 14732 14434 14766
rect 14468 14732 14508 14766
rect 14542 14732 14583 14766
rect 14617 14732 14695 14766
rect 13170 14723 13440 14732
rect 13492 14723 13504 14732
rect 13556 14723 14695 14732
rect 13170 14708 13216 14723
tri 13216 14708 13231 14723 nw
tri 14454 14708 14469 14723 ne
rect 14469 14708 14695 14723
tri 14469 14693 14484 14708 ne
rect 14484 14693 14695 14708
tri 14484 14691 14486 14693 ne
tri 1686 14680 1693 14687 se
rect 1693 14680 1744 14687
tri 1744 14680 1751 14687 nw
tri 1802 14680 1809 14687 se
rect 1809 14680 1860 14687
tri 1860 14680 1867 14687 nw
tri 12737 14680 12744 14687 se
rect 12744 14680 12794 14687
tri 1672 14666 1686 14680 se
rect 1686 14666 1730 14680
tri 1730 14666 1744 14680 nw
tri 1788 14666 1802 14680 se
rect 1802 14666 1846 14680
tri 1846 14666 1860 14680 nw
tri 12723 14666 12737 14680 se
rect 12737 14666 12794 14680
tri 13219 14666 13233 14680 se
rect 13233 14666 14276 14680
tri 1665 14659 1672 14666 se
rect 1672 14659 1723 14666
tri 1723 14659 1730 14666 nw
tri 1781 14659 1788 14666 se
rect 1788 14659 1839 14666
tri 1839 14659 1846 14666 nw
tri 12716 14659 12723 14666 se
rect 12723 14659 12794 14666
tri 1657 14651 1665 14659 se
rect 1665 14651 1715 14659
tri 1715 14651 1723 14659 nw
tri 1773 14651 1781 14659 se
rect 1781 14651 1812 14659
tri 1640 14634 1657 14651 se
rect 1657 14634 1698 14651
tri 1698 14634 1715 14651 nw
tri 1756 14634 1773 14651 se
rect 1773 14634 1812 14651
rect 1640 14632 1696 14634
tri 1696 14632 1698 14634 nw
tri 1754 14632 1756 14634 se
rect 1756 14632 1812 14634
tri 1812 14632 1839 14659 nw
rect 1640 14629 1693 14632
tri 1693 14629 1696 14632 nw
tri 1751 14629 1754 14632 se
rect 1754 14629 1809 14632
tri 1809 14629 1812 14632 nw
rect 1640 14468 1680 14629
tri 1680 14616 1693 14629 nw
tri 1738 14616 1751 14629 se
rect 1751 14616 1795 14629
tri 1737 14615 1738 14616 se
rect 1738 14615 1795 14616
tri 1795 14615 1809 14629 nw
rect 3139 14615 6626 14659
tri 1735 14613 1737 14615 se
rect 1737 14613 1793 14615
tri 1793 14613 1795 14615 nw
rect 3139 14614 4237 14615
tri 4237 14614 4238 14615 nw
tri 6612 14614 6613 14615 ne
rect 6613 14614 6626 14615
rect 3139 14613 4236 14614
tri 4236 14613 4237 14614 nw
tri 6613 14613 6614 14614 ne
rect 6614 14613 6626 14614
tri 1720 14598 1735 14613 se
rect 1735 14598 1778 14613
tri 1778 14598 1793 14613 nw
rect 1720 14583 1763 14598
tri 1763 14583 1778 14598 nw
rect 3139 14583 3189 14613
tri 3189 14583 3219 14613 nw
tri 3888 14583 3918 14613 ne
rect 3918 14607 4230 14613
tri 4230 14607 4236 14613 nw
tri 6614 14607 6620 14613 ne
rect 6620 14607 6626 14613
rect 6678 14607 6690 14659
rect 6742 14615 12794 14659
tri 13185 14632 13219 14666 se
rect 13219 14634 14276 14666
rect 13219 14632 13251 14634
tri 13251 14632 13253 14634 nw
tri 13684 14632 13686 14634 ne
rect 13686 14632 13796 14634
tri 13796 14632 13798 14634 nw
tri 14196 14632 14198 14634 ne
rect 14198 14632 14276 14634
tri 13168 14615 13185 14632 se
rect 13185 14615 13233 14632
rect 6742 14614 6755 14615
tri 6755 14614 6756 14615 nw
tri 13167 14614 13168 14615 se
rect 13168 14614 13233 14615
tri 13233 14614 13251 14632 nw
tri 13686 14614 13704 14632 ne
rect 13704 14614 13778 14632
tri 13778 14614 13796 14632 nw
tri 14198 14614 14216 14632 ne
rect 14216 14614 14276 14632
rect 6742 14607 6748 14614
tri 6748 14607 6755 14614 nw
tri 13160 14607 13167 14614 se
rect 13167 14607 13208 14614
rect 3918 14589 4212 14607
tri 4212 14589 4230 14607 nw
tri 13142 14589 13160 14607 se
rect 13160 14589 13208 14607
tri 13208 14589 13233 14614 nw
tri 13704 14600 13718 14614 ne
rect 3918 14583 4206 14589
tri 4206 14583 4212 14589 nw
tri 13136 14583 13142 14589 se
rect 13142 14583 13202 14589
tri 13202 14583 13208 14589 nw
rect 1720 14468 1760 14583
tri 1760 14580 1763 14583 nw
rect 3059 14558 3111 14564
rect 3059 14492 3111 14506
rect 3059 14426 3111 14440
rect 3059 14366 3071 14374
rect 3105 14366 3111 14374
rect 3059 14360 3111 14366
rect -547 14202 2091 14308
rect 3059 14294 3071 14308
rect 3105 14294 3111 14308
rect 3059 14228 3071 14242
rect 3105 14228 3111 14242
rect -547 14196 -301 14202
tri -301 14196 -295 14202 nw
tri 1959 14196 1965 14202 ne
rect 1965 14196 2045 14202
rect -547 14172 -325 14196
tri -325 14172 -301 14196 nw
tri 1965 14172 1989 14196 ne
rect 1989 14172 2045 14196
rect -547 14170 -327 14172
tri -327 14170 -325 14172 nw
tri 1989 14170 1991 14172 ne
rect 1991 14170 2045 14172
rect -547 14158 -339 14170
tri -339 14158 -327 14170 nw
rect -259 14158 -213 14170
tri -213 14158 -201 14170 sw
tri 241 14158 253 14170 se
rect 253 14158 299 14170
tri 299 14158 311 14170 sw
tri 753 14158 765 14170 se
rect 765 14158 811 14170
tri 811 14158 823 14170 sw
tri 1265 14158 1277 14170 se
rect 1277 14158 1323 14170
tri 1323 14158 1335 14170 sw
tri 1777 14158 1789 14170 se
rect 1789 14158 1835 14170
rect -547 14124 -373 14158
tri -373 14124 -339 14158 nw
rect -259 14124 -253 14158
rect -219 14128 -201 14158
tri -201 14128 -171 14158 sw
tri 211 14128 241 14158 se
rect 241 14128 259 14158
rect -219 14124 259 14128
rect 293 14128 311 14158
tri 311 14128 341 14158 sw
tri 723 14128 753 14158 se
rect 753 14128 771 14158
rect 293 14124 771 14128
rect 805 14128 823 14158
tri 823 14128 853 14158 sw
tri 1235 14128 1265 14158 se
rect 1265 14128 1283 14158
rect 805 14124 1283 14128
rect 1317 14128 1335 14158
tri 1335 14128 1365 14158 sw
tri 1747 14128 1777 14158 se
rect 1777 14128 1795 14158
rect 1317 14124 1795 14128
rect 1829 14124 1835 14158
tri 1991 14138 2023 14170 ne
rect 2023 14138 2045 14170
tri 2023 14136 2025 14138 ne
rect 2025 14136 2045 14138
tri 2025 14124 2037 14136 ne
rect 2037 14124 2045 14136
rect -547 13623 -381 14124
tri -381 14116 -373 14124 nw
rect -259 14086 1835 14124
tri 2037 14116 2045 14124 ne
rect 3059 14172 3111 14176
rect 3059 14162 3071 14172
rect 3105 14162 3111 14172
rect -259 14083 259 14086
rect -259 14049 -253 14083
rect -219 14082 259 14083
rect -219 14052 -201 14082
tri -201 14052 -171 14082 nw
tri 211 14052 241 14082 ne
rect 241 14052 259 14082
rect 293 14082 771 14086
rect 293 14052 311 14082
tri 311 14052 341 14082 nw
tri 723 14052 753 14082 ne
rect 753 14052 771 14082
rect 805 14082 1283 14086
rect 805 14052 823 14082
tri 823 14052 853 14082 nw
tri 1235 14052 1265 14082 ne
rect 1265 14052 1283 14082
rect 1317 14082 1795 14086
rect 1317 14052 1335 14082
tri 1335 14052 1365 14082 nw
tri 1747 14052 1777 14082 ne
rect 1777 14052 1795 14082
rect 1829 14052 1835 14086
rect -219 14049 -213 14052
rect -259 14008 -213 14049
tri -213 14040 -201 14052 nw
tri 241 14040 253 14052 ne
rect 253 14040 299 14052
tri 299 14040 311 14052 nw
tri 753 14040 765 14052 ne
rect 765 14040 811 14052
tri 811 14040 823 14052 nw
tri 1265 14040 1277 14052 ne
rect 1277 14040 1323 14052
tri 1323 14040 1335 14052 nw
tri 1777 14040 1789 14052 ne
rect 1789 14040 1835 14052
rect 3059 14096 3111 14110
rect -259 13974 -253 14008
rect -219 13974 -213 14008
rect 3059 14030 3111 14044
rect -259 13932 -213 13974
rect -259 13898 -253 13932
rect -219 13898 -213 13932
rect -259 13847 -213 13898
rect 509 13988 555 14000
tri 555 13988 567 14000 sw
tri 1521 13988 1533 14000 se
rect 1533 13988 1579 14000
rect 509 13954 515 13988
rect 549 13958 567 13988
tri 567 13958 597 13988 sw
tri 1491 13958 1521 13988 se
rect 1521 13958 1539 13988
rect 549 13954 1539 13958
rect 1573 13954 1579 13988
rect 509 13916 1579 13954
rect 509 13882 515 13916
rect 549 13912 1579 13916
rect 549 13882 563 13912
rect 509 13878 563 13882
tri 563 13878 597 13912 nw
tri 1491 13893 1510 13912 ne
rect 1510 13893 1539 13912
tri 1510 13891 1512 13893 ne
rect 1512 13891 1539 13893
tri 1512 13878 1525 13891 ne
rect 1525 13878 1539 13891
rect 1573 13878 1579 13912
rect 509 13870 555 13878
tri 555 13870 563 13878 nw
tri 1525 13870 1533 13878 ne
tri -213 13847 -197 13863 sw
rect -259 13836 -197 13847
tri -197 13836 -186 13847 sw
rect 1533 13836 1579 13878
rect -259 13835 -186 13836
tri -259 13818 -242 13835 ne
rect -242 13830 -186 13835
tri -186 13830 -180 13836 sw
rect -242 13818 -180 13830
tri -180 13818 -168 13830 sw
rect -3 13818 43 13830
tri 43 13818 55 13830 sw
tri 1009 13818 1021 13830 se
rect 1021 13818 1067 13830
tri -242 13784 -208 13818 ne
rect -208 13784 -168 13818
tri -168 13784 -134 13818 sw
rect -3 13784 3 13818
rect 37 13804 55 13818
tri 55 13804 69 13818 sw
tri 995 13804 1009 13818 se
rect 1009 13804 1027 13818
rect 37 13788 69 13804
tri 69 13788 85 13804 sw
tri 979 13788 995 13804 se
rect 995 13788 1027 13804
rect 37 13784 1027 13788
rect 1061 13784 1067 13818
tri -208 13773 -197 13784 ne
rect -197 13773 -134 13784
tri -134 13773 -123 13784 sw
tri -197 13760 -184 13773 ne
rect -184 13760 -123 13773
tri -184 13751 -175 13760 ne
rect -570 13572 -381 13623
rect -597 13466 -381 13572
rect -570 13451 -381 13466
tri -381 13451 -373 13459 sw
rect -570 13447 -373 13451
tri -373 13447 -369 13451 sw
rect -570 13416 -369 13447
tri -369 13416 -338 13447 sw
rect -570 13410 -218 13416
rect -570 13376 -492 13410
rect -458 13376 -416 13410
rect -382 13376 -340 13410
rect -306 13376 -264 13410
rect -230 13376 -218 13410
rect -570 13370 -218 13376
rect -570 13340 -368 13370
tri -368 13340 -338 13370 nw
rect -570 13335 -381 13340
rect -570 13301 -564 13335
rect -530 13301 -381 13335
tri -381 13327 -368 13340 nw
rect -570 13260 -381 13301
rect -570 13226 -564 13260
rect -530 13226 -381 13260
rect -570 13185 -381 13226
rect -570 13151 -564 13185
rect -530 13151 -381 13185
rect -570 13110 -381 13151
rect -570 13076 -564 13110
rect -530 13076 -381 13110
rect -570 13035 -381 13076
rect -570 13001 -564 13035
rect -530 13001 -381 13035
rect -570 12960 -381 13001
rect -570 12926 -564 12960
rect -530 12926 -381 12960
rect -570 12885 -381 12926
rect -570 12851 -564 12885
rect -530 12851 -381 12885
rect -570 12810 -381 12851
rect -570 12776 -564 12810
rect -530 12776 -381 12810
rect -570 12735 -381 12776
rect -570 12701 -564 12735
rect -530 12701 -381 12735
rect -570 12659 -381 12701
rect -570 12625 -564 12659
rect -530 12625 -381 12659
rect -570 12583 -381 12625
rect -570 12549 -564 12583
rect -530 12549 -381 12583
rect -570 12507 -381 12549
rect -570 12473 -564 12507
rect -530 12473 -381 12507
rect -570 12431 -381 12473
rect -570 12397 -564 12431
rect -530 12397 -381 12431
rect -570 12355 -381 12397
rect -570 12321 -564 12355
rect -530 12321 -381 12355
rect -570 12279 -381 12321
rect -570 12245 -564 12279
rect -530 12245 -381 12279
rect -570 12203 -381 12245
rect -570 12169 -564 12203
rect -530 12169 -381 12203
rect -570 12159 -381 12169
rect -175 12992 -123 13760
rect -3 13746 1067 13784
rect -3 13712 3 13746
rect 37 13742 1027 13746
rect 37 13712 55 13742
tri 55 13712 85 13742 nw
tri 979 13712 1009 13742 ne
rect 1009 13712 1027 13742
rect 1061 13712 1067 13746
tri -4 13639 -3 13640 se
rect -3 13639 43 13712
tri 43 13700 55 13712 nw
tri 1009 13700 1021 13712 ne
rect 1021 13700 1067 13712
rect 1533 13802 1539 13836
rect 1573 13802 1579 13836
rect 1533 13760 1579 13802
rect 1533 13726 1539 13760
rect 1573 13726 1579 13760
tri 43 13639 49 13645 sw
tri -37 13606 -4 13639 se
rect -4 13606 49 13639
tri 49 13606 82 13639 sw
rect -68 13600 1407 13606
rect -68 13566 -56 13600
rect -22 13566 19 13600
rect 53 13566 94 13600
rect 128 13566 169 13600
rect 203 13566 244 13600
rect 278 13566 319 13600
rect 353 13566 394 13600
rect 428 13566 469 13600
rect 503 13566 544 13600
rect 578 13566 619 13600
rect 653 13566 694 13600
rect 728 13566 769 13600
rect 803 13566 843 13600
rect 877 13566 917 13600
rect 951 13566 991 13600
rect 1025 13566 1065 13600
rect 1099 13566 1139 13600
rect 1173 13566 1213 13600
rect 1247 13566 1287 13600
rect 1321 13566 1361 13600
rect 1395 13566 1407 13600
rect -68 13554 1407 13566
rect 1533 13562 1579 13726
rect 3059 13964 3111 13978
rect 3059 13910 3071 13912
rect 3105 13910 3111 13912
rect 3059 13898 3111 13910
rect 3059 13834 3071 13846
rect 3105 13834 3111 13846
rect 3059 13832 3111 13834
rect 3059 13765 3071 13780
rect 3105 13765 3111 13780
rect 3059 13698 3071 13713
rect 3105 13698 3111 13713
rect 3059 13639 3111 13646
rect 3059 13631 3071 13639
rect 3105 13631 3111 13639
rect 3059 13564 3111 13579
tri 1579 13562 1580 13563 sw
tri -37 13528 -11 13554 ne
rect -11 13534 57 13554
tri 57 13534 77 13554 nw
rect 1533 13543 1580 13562
tri 1533 13534 1542 13543 ne
rect 1542 13534 1580 13543
tri 1580 13534 1608 13562 sw
rect -11 13528 51 13534
tri 51 13528 57 13534 nw
tri 1542 13528 1548 13534 ne
rect 1548 13528 1608 13534
tri 1608 13528 1614 13534 sw
tri -11 13520 -3 13528 ne
rect -3 13413 43 13528
tri 43 13520 51 13528 nw
tri 1548 13520 1556 13528 ne
rect 1556 13520 1614 13528
tri 1614 13520 1622 13528 sw
tri 1556 13497 1579 13520 ne
rect 1579 13497 1622 13520
tri 1579 13486 1590 13497 ne
rect 1590 13486 1622 13497
tri 1622 13486 1656 13520 sw
rect 3059 13497 3111 13512
tri 1590 13485 1591 13486 ne
rect 1591 13485 1656 13486
tri 1656 13485 1657 13486 sw
tri 1591 13468 1608 13485 ne
rect 1608 13468 1657 13485
tri 1657 13468 1674 13485 sw
tri 1608 13451 1625 13468 ne
rect 1625 13451 1674 13468
tri 1674 13451 1691 13468 sw
tri 1625 13447 1629 13451 ne
rect 1629 13447 1691 13451
tri 1691 13447 1695 13451 sw
tri 1629 13421 1655 13447 ne
rect 1655 13421 1695 13447
tri 1695 13421 1721 13447 sw
rect 3059 13439 3111 13445
tri 43 13413 51 13421 sw
tri 1655 13413 1663 13421 ne
rect 1663 13413 1721 13421
tri 1721 13413 1729 13421 sw
rect -3 13404 51 13413
tri 51 13404 60 13413 sw
tri 1663 13404 1672 13413 ne
rect 1672 13404 1729 13413
tri 1729 13404 1738 13413 sw
rect -3 13397 60 13404
tri -3 13387 7 13397 ne
rect 7 13387 60 13397
tri 60 13387 77 13404 sw
tri 1672 13402 1674 13404 ne
rect 1674 13402 1738 13404
tri 1738 13402 1740 13404 sw
tri 1674 13387 1689 13402 ne
rect 1689 13387 1740 13402
tri 1740 13387 1755 13402 sw
tri 7 13374 20 13387 ne
rect 20 13374 77 13387
tri 77 13374 90 13387 sw
tri 1689 13374 1702 13387 ne
rect 1702 13374 1755 13387
tri 1755 13374 1768 13387 sw
tri 20 13340 54 13374 ne
rect 54 13370 90 13374
tri 90 13370 94 13374 sw
tri 1702 13370 1706 13374 ne
rect 1706 13370 1768 13374
tri 1768 13370 1772 13374 sw
rect 54 13340 94 13370
tri 94 13340 124 13370 sw
tri 1706 13340 1736 13370 ne
rect 1736 13340 1772 13370
tri 1772 13340 1802 13370 sw
tri 3109 13340 3139 13370 se
rect 3139 13340 3185 14583
tri 3185 14579 3189 14583 nw
tri 3918 14579 3922 14583 ne
tri 54 13334 60 13340 ne
rect 60 13336 124 13340
tri 124 13336 128 13340 sw
tri 1736 13336 1740 13340 ne
rect 1740 13336 1802 13340
tri 1802 13336 1806 13340 sw
tri 3105 13336 3109 13340 se
rect 3109 13336 3185 13340
rect 60 13334 128 13336
tri 128 13334 130 13336 sw
tri 1740 13334 1742 13336 ne
rect 1742 13334 3185 13336
tri 60 13319 75 13334 ne
rect 75 13319 473 13334
tri 473 13319 488 13334 sw
tri 1742 13319 1757 13334 ne
rect 1757 13319 3185 13334
tri 75 13314 80 13319 ne
rect 80 13314 488 13319
tri 488 13314 493 13319 sw
tri 1757 13314 1762 13319 ne
rect 1762 13314 3185 13319
tri 80 13310 84 13314 ne
rect 84 13310 493 13314
tri 493 13310 497 13314 sw
tri 1762 13310 1766 13314 ne
rect 1766 13310 3185 13314
tri 84 13301 93 13310 ne
rect 93 13301 497 13310
tri 497 13301 506 13310 sw
tri 1766 13301 1775 13310 ne
rect 1775 13301 3185 13310
tri 93 13284 110 13301 ne
rect 110 13284 506 13301
tri 453 13267 470 13284 ne
rect 470 13267 506 13284
tri 506 13267 540 13301 sw
tri 1775 13290 1786 13301 ne
rect 1786 13290 3185 13301
rect 3214 14532 3496 14541
rect 3214 14498 3300 14532
rect 3334 14498 3372 14532
rect 3406 14498 3496 14532
tri 470 13247 490 13267 ne
rect 490 13247 540 13267
tri 540 13247 560 13267 sw
tri 490 13241 496 13247 ne
rect 496 13241 560 13247
tri 560 13241 566 13247 sw
tri 496 13240 497 13241 ne
rect 497 13240 566 13241
tri 566 13240 567 13241 sw
tri 497 13228 509 13240 ne
rect 509 13228 567 13240
tri 567 13228 579 13240 sw
tri 509 13194 543 13228 ne
rect 543 13194 579 13228
tri 579 13194 613 13228 sw
tri 543 13175 562 13194 ne
rect 562 13175 613 13194
tri 613 13175 632 13194 sw
tri 562 13170 567 13175 ne
rect 567 13170 632 13175
tri 632 13170 637 13175 sw
tri 567 13168 569 13170 ne
rect 569 13168 637 13170
tri 637 13168 639 13170 sw
tri 569 13155 582 13168 ne
rect 582 13155 639 13168
tri 639 13155 652 13168 sw
tri 582 13151 586 13155 ne
rect 586 13151 652 13155
tri 652 13151 656 13155 sw
rect -175 12928 -123 12940
rect -175 12864 -123 12876
rect -175 12800 -123 12812
rect -175 12735 -123 12748
rect -175 12670 -123 12683
rect -175 12605 -123 12618
rect -175 12540 -123 12553
rect -175 12475 -123 12488
rect -175 12410 -123 12423
rect -175 12345 -123 12358
rect -175 12280 -123 12293
rect -175 12215 -123 12228
tri -381 12159 -377 12163 sw
rect -570 12157 -377 12159
tri -377 12157 -375 12159 sw
rect -175 12157 -123 12163
tri 81 12159 85 12163 se
rect 85 12159 249 13151
tri 586 13121 616 13151 ne
rect 616 13134 656 13151
tri 656 13134 673 13151 sw
rect 616 13121 673 13134
tri 673 13121 686 13134 sw
tri 3201 13121 3214 13134 se
rect 3214 13121 3496 14498
rect 3529 14532 3659 14541
rect 3529 14498 3541 14532
rect 3575 14498 3613 14532
rect 3647 14498 3659 14532
rect 3529 14489 3659 14498
rect 3760 14532 3890 14541
rect 3760 14498 3772 14532
rect 3806 14498 3844 14532
rect 3878 14498 3890 14532
rect 3760 14489 3890 14498
rect 3922 14532 4204 14583
tri 4204 14581 4206 14583 nw
tri 13134 14581 13136 14583 se
rect 13136 14581 13168 14583
tri 13102 14549 13134 14581 se
rect 13134 14549 13168 14581
tri 13168 14549 13202 14583 nw
tri 13101 14548 13102 14549 se
rect 13102 14548 13167 14549
tri 13167 14548 13168 14549 nw
tri 13096 14543 13101 14548 se
rect 13101 14543 13162 14548
tri 13162 14543 13167 14548 nw
tri 13091 14538 13096 14543 se
rect 13096 14538 13150 14543
rect 3922 14498 4008 14532
rect 4042 14498 4080 14532
rect 4114 14498 4204 14532
tri 13084 14531 13091 14538 se
rect 13091 14531 13150 14538
tri 13150 14531 13162 14543 nw
tri 13072 14519 13084 14531 se
rect 13084 14519 13138 14531
tri 13138 14519 13150 14531 nw
tri 13057 14504 13072 14519 se
rect 13072 14504 13103 14519
tri 3530 14484 3535 14489 ne
rect 3535 14484 3639 14489
tri 3639 14484 3644 14489 nw
tri 3770 14484 3775 14489 ne
rect 3775 14484 3879 14489
tri 3879 14484 3884 14489 nw
tri 3535 14468 3551 14484 ne
rect 3551 14468 3610 14484
tri 3551 14455 3564 14468 ne
tri 616 13103 634 13121 ne
rect 634 13103 686 13121
tri 686 13103 704 13121 sw
tri 3183 13103 3201 13121 se
rect 3201 13103 3496 13121
tri 634 13100 637 13103 ne
rect 637 13100 704 13103
tri 704 13100 707 13103 sw
tri 3180 13100 3183 13103 se
rect 3183 13100 3496 13103
tri 637 13095 642 13100 ne
rect 642 13095 3496 13100
tri 642 13082 655 13095 ne
rect 655 13082 3496 13095
tri 655 13054 683 13082 ne
rect 683 13054 3496 13082
tri 3180 13048 3186 13054 ne
rect 3186 13048 3496 13054
tri 3186 13032 3202 13048 ne
rect 3202 13032 3496 13048
tri 3202 13031 3203 13032 ne
rect 3203 13031 3496 13032
tri 3203 13022 3212 13031 ne
rect 3212 13022 3496 13031
tri 3212 13020 3214 13022 ne
rect 3214 12428 3496 13022
tri 3562 12431 3564 12433 se
rect 3564 12431 3610 14468
tri 3610 14455 3639 14484 nw
tri 3775 14455 3804 14484 ne
tri 3610 12431 3612 12433 sw
tri 3802 12431 3804 12433 se
rect 3804 12431 3850 14484
tri 3850 14455 3879 14484 nw
tri 3850 12431 3852 12433 sw
tri 3559 12428 3562 12431 se
rect 3562 12428 3612 12431
tri 3254 12425 3257 12428 ne
rect 3257 12425 3449 12428
tri 3449 12425 3452 12428 nw
tri 3556 12425 3559 12428 se
rect 3559 12425 3612 12428
tri 3612 12425 3618 12431 sw
tri 3799 12428 3802 12431 se
rect 3802 12428 3852 12431
tri 3852 12428 3855 12431 sw
rect 3922 12428 4204 14498
rect 4659 14458 12266 14504
tri 13045 14492 13057 14504 se
rect 13057 14492 13103 14504
tri 13037 14484 13045 14492 se
rect 13045 14484 13103 14492
tri 13103 14484 13138 14519 nw
tri 13035 14482 13037 14484 se
rect 13037 14482 13101 14484
tri 13101 14482 13103 14484 nw
rect 4659 14450 4731 14458
tri 4731 14450 4739 14458 nw
tri 12186 14450 12194 14458 ne
rect 12194 14450 12266 14458
tri 13003 14450 13035 14482 se
rect 13035 14450 13069 14482
tri 13069 14450 13101 14482 nw
rect 13718 14473 13764 14614
tri 13764 14600 13778 14614 nw
tri 14216 14600 14230 14614 ne
rect 13804 14583 13941 14592
rect 13804 14549 13816 14583
rect 13850 14549 13888 14583
rect 13922 14549 13941 14583
rect 13804 14540 13941 14549
rect 13993 14540 14005 14592
rect 14057 14583 14190 14592
rect 14057 14549 14072 14583
rect 14106 14549 14144 14583
rect 14178 14549 14190 14583
rect 14057 14540 14190 14549
tri 13812 14531 13821 14540 ne
rect 13821 14531 13917 14540
tri 13917 14531 13926 14540 nw
tri 14060 14531 14069 14540 ne
rect 14069 14531 14165 14540
tri 14165 14531 14174 14540 nw
tri 13821 14506 13846 14531 ne
rect 13458 14467 13510 14473
rect 4370 12875 4449 14398
rect 4659 13559 4705 14450
tri 4705 14424 4731 14450 nw
tri 12194 14424 12220 14450 ne
rect 4915 14391 5286 14398
rect 4915 14386 5132 14391
rect 4915 14352 5087 14386
rect 5121 14352 5132 14386
rect 4915 14339 5132 14352
rect 5184 14339 5232 14391
rect 5284 14339 5286 14391
rect 4915 14326 5286 14339
rect 4915 14314 5132 14326
rect 4915 14280 5087 14314
rect 5121 14280 5132 14314
rect 4915 14274 5132 14280
rect 5184 14274 5232 14326
rect 5284 14274 5286 14326
rect 4915 14261 5286 14274
rect 4915 14242 5132 14261
rect 4915 14208 5087 14242
rect 5121 14209 5132 14242
rect 5184 14209 5232 14261
rect 5284 14209 5286 14261
rect 5121 14208 5286 14209
rect 4915 14196 5286 14208
rect 4915 14170 5132 14196
rect 4915 14136 5087 14170
rect 5121 14144 5132 14170
rect 5184 14144 5232 14196
rect 5284 14144 5286 14196
rect 5121 14136 5286 14144
rect 4915 14131 5286 14136
rect 4915 14098 5132 14131
rect 4915 14064 5087 14098
rect 5121 14079 5132 14098
rect 5184 14079 5232 14131
rect 5284 14079 5286 14131
rect 8703 14124 10371 14130
rect 8703 14090 8715 14124
rect 8749 14090 8787 14124
rect 8821 14090 10319 14124
rect 8703 14084 10319 14090
rect 5121 14066 5286 14079
rect 5121 14064 5132 14066
rect 4915 14026 5132 14064
rect 4915 13992 5087 14026
rect 5121 14014 5132 14026
rect 5184 14014 5232 14066
rect 5284 14014 5286 14066
tri 10285 14052 10317 14084 ne
rect 10317 14072 10319 14084
rect 10317 14060 10371 14072
rect 10317 14052 10319 14060
tri 10317 14050 10319 14052 ne
rect 5121 14001 5286 14014
rect 10319 14002 10371 14008
rect 5121 13992 5132 14001
rect 4915 13954 5132 13992
rect 4915 13920 5087 13954
rect 5121 13949 5132 13954
rect 5184 13949 5232 14001
rect 5284 13949 5286 14001
rect 5121 13936 5286 13949
rect 5121 13920 5132 13936
rect 4915 13884 5132 13920
rect 5184 13884 5232 13936
rect 5284 13884 5286 13936
rect 7743 13969 7795 13975
rect 7743 13905 7795 13917
tri 6614 13891 6616 13893 se
rect 6616 13891 6622 13893
rect 4915 13882 5286 13884
rect 4915 13848 5087 13882
rect 5121 13870 5286 13882
rect 5121 13848 5132 13870
rect 4915 13818 5132 13848
rect 5184 13818 5232 13870
rect 5284 13818 5286 13870
rect 5728 13885 6622 13891
rect 5728 13851 5740 13885
rect 5774 13851 5812 13885
rect 5846 13851 6622 13885
rect 5728 13845 6622 13851
tri 6612 13841 6616 13845 ne
rect 6616 13841 6622 13845
rect 6674 13841 6686 13893
rect 6738 13841 6744 13893
rect 7743 13847 7795 13853
tri 7743 13841 7749 13847 ne
rect 7749 13841 7795 13847
tri 7749 13836 7754 13841 ne
rect 7754 13836 7795 13841
tri 7754 13835 7755 13836 ne
rect 4915 13810 5286 13818
rect 4915 13798 5087 13810
rect 4915 13746 4936 13798
rect 4988 13776 5087 13798
rect 5121 13804 5286 13810
rect 5121 13776 5132 13804
rect 4988 13752 5132 13776
rect 5184 13752 5232 13804
rect 5284 13752 5286 13804
rect 4988 13746 5286 13752
rect 4915 13738 5286 13746
rect 4915 13734 5087 13738
rect 4915 13682 4936 13734
rect 4988 13704 5087 13734
rect 5121 13704 5132 13738
rect 4988 13686 5132 13704
rect 5184 13686 5232 13738
rect 5284 13686 5286 13738
rect 4988 13682 5286 13686
rect 4915 13672 5286 13682
rect 4915 13670 5132 13672
rect 4915 13618 4936 13670
rect 4988 13666 5132 13670
rect 4988 13632 5087 13666
rect 5121 13632 5132 13666
rect 4988 13620 5132 13632
rect 5184 13620 5232 13672
rect 5284 13620 5286 13672
rect 4988 13618 5286 13620
rect 4915 13606 5286 13618
rect 4915 13554 4936 13606
rect 4988 13593 5132 13606
rect 4988 13559 5087 13593
rect 5121 13559 5132 13593
rect 4988 13554 5132 13559
rect 5184 13554 5232 13606
rect 5284 13554 5286 13606
rect 4915 13542 5286 13554
rect 4915 13490 4936 13542
rect 4988 13540 5286 13542
rect 4988 13520 5132 13540
rect 4988 13490 5087 13520
rect 4915 13486 5087 13490
rect 5121 13488 5132 13520
rect 5184 13488 5232 13540
rect 5284 13488 5286 13540
rect 5121 13486 5286 13488
rect 4915 13478 5286 13486
rect 4915 13426 4936 13478
rect 4988 13474 5286 13478
rect 4988 13447 5132 13474
rect 4988 13426 5087 13447
rect 4915 13414 5087 13426
rect 4915 13362 4936 13414
rect 4988 13413 5087 13414
rect 5121 13422 5132 13447
rect 5184 13422 5232 13474
rect 5284 13422 5286 13474
rect 5121 13413 5286 13422
rect 4988 13408 5286 13413
rect 4988 13374 5132 13408
rect 4988 13362 5087 13374
rect 4915 13350 5087 13362
rect 4915 13298 4936 13350
rect 4988 13340 5087 13350
rect 5121 13356 5132 13374
rect 5184 13356 5232 13408
rect 5284 13356 5286 13408
rect 5121 13342 5286 13356
rect 5121 13340 5132 13342
rect 4988 13301 5132 13340
rect 4988 13298 5087 13301
rect 4915 13285 5087 13298
rect 4915 13233 4936 13285
rect 4988 13267 5087 13285
rect 5121 13290 5132 13301
rect 5184 13290 5232 13342
rect 5284 13290 5286 13342
rect 5121 13276 5286 13290
rect 5121 13267 5132 13276
rect 4988 13233 5132 13267
rect 4915 13228 5132 13233
rect 4915 13220 5087 13228
rect 4915 13168 4936 13220
rect 4988 13194 5087 13220
rect 5121 13224 5132 13228
rect 5184 13224 5232 13276
rect 5284 13224 5286 13276
rect 5121 13210 5286 13224
rect 5121 13194 5132 13210
rect 4988 13168 5132 13194
rect 4915 13158 5132 13168
rect 5184 13158 5232 13210
rect 5284 13158 5286 13210
rect 4915 13155 5286 13158
rect 4915 13103 4936 13155
rect 4988 13121 5087 13155
rect 5121 13144 5286 13155
rect 5121 13121 5132 13144
rect 4988 13103 5132 13121
rect 4915 13092 5132 13103
rect 5184 13092 5232 13144
rect 5284 13092 5286 13144
rect 4915 13090 5286 13092
rect 4915 13038 4936 13090
rect 4988 13082 5286 13090
rect 4988 13048 5087 13082
rect 5121 13078 5286 13082
rect 5121 13048 5132 13078
rect 4988 13038 5132 13048
rect 4915 13026 5132 13038
rect 5184 13026 5232 13078
rect 5284 13026 5286 13078
rect 4915 13012 5286 13026
rect 4915 13009 5132 13012
rect 4915 12975 5087 13009
rect 5121 12975 5132 13009
rect 4489 12962 4728 12969
rect 4780 12962 4792 12969
rect 4844 12962 4875 12969
rect 4489 12928 4501 12962
rect 4535 12928 4573 12962
rect 4607 12928 4728 12962
rect 4791 12928 4792 12962
rect 4863 12928 4875 12962
rect 4489 12917 4728 12928
rect 4780 12917 4792 12928
rect 4844 12917 4875 12928
rect 4915 12960 5132 12975
rect 5184 12960 5232 13012
rect 5284 12960 5286 13012
rect 4915 12946 5286 12960
rect 4915 12936 5132 12946
rect 4915 12902 5087 12936
rect 5121 12902 5132 12936
rect 4915 12894 5132 12902
rect 5184 12894 5232 12946
rect 5284 12894 5286 12946
tri 4449 12875 4461 12887 sw
tri 4903 12875 4915 12887 se
rect 4915 12880 5286 12894
rect 4915 12875 5132 12880
rect 4370 12863 4461 12875
tri 4461 12863 4473 12875 sw
tri 4891 12863 4903 12875 se
rect 4903 12863 5132 12875
rect 4370 12853 4473 12863
tri 4473 12853 4483 12863 sw
tri 4881 12853 4891 12863 se
rect 4891 12853 5087 12863
rect 4370 12852 5087 12853
rect 4370 12800 4384 12852
rect 4436 12800 4454 12852
rect 4506 12800 4524 12852
rect 4576 12800 4594 12852
rect 4646 12800 4664 12852
rect 4716 12800 4734 12852
rect 4786 12800 4803 12852
rect 4855 12829 5087 12852
rect 5121 12829 5132 12863
rect 4855 12828 5132 12829
rect 5184 12828 5232 12880
rect 5284 12828 5286 12880
rect 4855 12814 5286 12828
rect 4855 12800 5132 12814
rect 4370 12790 5132 12800
rect 4370 12782 5087 12790
rect 4370 12730 4384 12782
rect 4436 12730 4454 12782
rect 4506 12730 4524 12782
rect 4576 12730 4594 12782
rect 4646 12730 4664 12782
rect 4716 12730 4734 12782
rect 4786 12730 4803 12782
rect 4855 12756 5087 12782
rect 5121 12762 5132 12790
rect 5184 12762 5232 12814
rect 5284 12762 5286 12814
rect 5121 12756 5286 12762
rect 4855 12748 5286 12756
rect 4855 12730 5132 12748
rect 4370 12727 4447 12730
tri 4447 12727 4450 12730 nw
tri 4848 12727 4851 12730 ne
rect 4851 12727 4959 12730
tri 4959 12727 4962 12730 nw
tri 5047 12727 5050 12730 ne
rect 5050 12727 5132 12730
rect 4370 12717 4437 12727
tri 4437 12717 4447 12727 nw
tri 4851 12717 4861 12727 ne
rect 4861 12717 4949 12727
tri 4949 12717 4959 12727 nw
tri 5050 12717 5060 12727 ne
rect 5060 12717 5132 12727
tri 4364 12704 4370 12710 se
rect 4370 12704 4416 12717
rect 4364 12698 4416 12704
tri 4416 12696 4437 12717 nw
tri 4861 12696 4882 12717 ne
rect 4882 12692 4928 12717
tri 4928 12696 4949 12717 nw
tri 5060 12696 5081 12717 ne
rect 4364 12626 4416 12646
rect 4364 12553 4416 12574
rect 4364 12480 4416 12501
tri 3257 12394 3288 12425 ne
rect 3288 12399 3423 12425
tri 3423 12399 3449 12425 nw
tri 3530 12399 3556 12425 se
rect 3556 12399 3618 12425
tri 3618 12399 3644 12425 sw
rect 3288 12396 3420 12399
tri 3420 12396 3423 12399 nw
rect 3288 12390 3418 12396
tri 3418 12394 3420 12396 nw
rect 3288 12356 3300 12390
rect 3334 12356 3372 12390
rect 3406 12356 3418 12390
rect 3288 12347 3418 12356
rect 3524 12390 3654 12399
rect 3524 12356 3536 12390
rect 3570 12356 3608 12390
rect 3642 12356 3654 12390
rect 3524 12347 3654 12356
tri 3536 12318 3565 12347 ne
rect 3565 12318 3621 12347
tri 3621 12318 3650 12347 nw
tri 3565 12313 3570 12318 ne
tri 79 12157 81 12159 se
rect 81 12157 249 12159
rect -570 12154 -375 12157
tri -375 12154 -372 12157 sw
tri 76 12154 79 12157 se
rect 79 12154 249 12157
rect -570 12139 -372 12154
tri -372 12139 -357 12154 sw
tri 61 12139 76 12154 se
rect 76 12139 249 12154
rect -570 12129 -357 12139
tri -357 12129 -347 12139 sw
tri 51 12129 61 12139 se
rect 61 12129 249 12139
rect -570 12083 249 12129
rect 359 12139 405 12157
tri 405 12139 406 12140 sw
rect 359 12120 406 12139
tri 406 12120 425 12139 sw
tri 359 12116 363 12120 ne
rect 363 12116 425 12120
tri 425 12116 429 12120 sw
tri 363 12110 369 12116 ne
rect 369 12110 429 12116
tri 429 12110 435 12116 sw
tri 369 12083 396 12110 ne
rect 396 12083 435 12110
tri 396 12076 403 12083 ne
rect 403 12076 435 12083
tri 435 12076 469 12110 sw
tri 403 12063 416 12076 ne
rect 416 12063 469 12076
tri 469 12063 482 12076 sw
tri 416 12054 425 12063 ne
rect 425 12054 482 12063
tri 482 12054 491 12063 sw
tri 425 12048 431 12054 ne
rect 431 12048 491 12054
rect -341 12042 367 12048
rect -341 12008 -329 12042
rect -295 12008 -257 12042
rect -223 12033 -73 12042
rect -223 12008 -201 12033
rect -341 12002 -201 12008
rect -149 12008 -73 12033
rect -39 12008 -1 12042
rect 33 12008 249 12042
rect 283 12008 321 12042
rect 355 12008 367 12042
tri 431 12015 464 12048 ne
rect 464 12015 491 12048
tri 491 12015 530 12054 sw
rect -149 12002 367 12008
tri 464 12002 477 12015 ne
rect 477 12002 530 12015
tri 477 11988 491 12002 ne
rect 491 11993 530 12002
tri 530 11993 552 12015 sw
rect 491 11988 552 11993
tri 491 11981 498 11988 ne
rect 498 11981 552 11988
rect -201 11969 -149 11981
tri 498 11973 506 11981 ne
rect -201 11911 -149 11917
rect 506 11700 552 11981
rect 3570 11821 3616 12318
tri 3616 12313 3621 12318 nw
rect 3686 12130 3732 12428
tri 3796 12425 3799 12428 se
rect 3799 12425 3855 12428
tri 3855 12425 3858 12428 sw
tri 3962 12425 3965 12428 ne
rect 3965 12425 4157 12428
tri 4157 12425 4160 12428 nw
tri 3770 12399 3796 12425 se
rect 3796 12399 3858 12425
tri 3858 12399 3884 12425 sw
tri 3965 12399 3991 12425 ne
rect 3991 12399 4131 12425
tri 4131 12399 4157 12425 nw
rect 4364 12407 4416 12428
rect 3760 12390 3890 12399
tri 3991 12396 3994 12399 ne
rect 3994 12396 4128 12399
tri 4128 12396 4131 12399 nw
tri 3994 12394 3996 12396 ne
rect 3760 12356 3772 12390
rect 3806 12356 3844 12390
rect 3878 12356 3890 12390
rect 3760 12347 3890 12356
rect 3996 12390 4126 12396
tri 4126 12394 4128 12396 nw
rect 3996 12356 4008 12390
rect 4042 12356 4080 12390
rect 4114 12356 4126 12390
rect 3996 12347 4126 12356
tri 3770 12318 3799 12347 ne
rect 3799 12318 3855 12347
tri 3855 12318 3884 12347 nw
rect 4364 12334 4416 12355
tri 3799 12313 3804 12318 ne
rect 3804 12245 3850 12318
tri 3850 12313 3855 12318 nw
rect 4364 12261 4416 12282
tri 3850 12245 3862 12257 sw
rect 3804 12243 3862 12245
tri 3862 12243 3864 12245 sw
rect 3804 12237 3864 12243
tri 3864 12237 3870 12243 sw
tri 4053 12237 4059 12243 se
rect 4059 12237 4065 12243
tri 3804 12226 3815 12237 ne
rect 3815 12226 4065 12237
tri 3815 12213 3828 12226 ne
rect 3828 12213 4065 12226
tri 3828 12206 3835 12213 ne
rect 3835 12206 4065 12213
tri 3835 12191 3850 12206 ne
rect 3850 12191 4065 12206
rect 4117 12191 4129 12243
rect 4181 12191 4187 12243
rect 4364 12188 4416 12209
rect 5081 12683 5087 12717
rect 5121 12696 5132 12717
rect 5184 12696 5232 12748
rect 5284 12696 5286 12748
rect 5121 12683 5286 12696
rect 5081 12682 5286 12683
rect 5081 12644 5132 12682
rect 5081 12610 5087 12644
rect 5121 12630 5132 12644
rect 5184 12630 5232 12682
rect 5284 12630 5286 12682
rect 5121 12616 5286 12630
rect 5121 12610 5132 12616
rect 5081 12571 5132 12610
rect 5081 12537 5087 12571
rect 5121 12564 5132 12571
rect 5184 12564 5232 12616
rect 5284 12564 5286 12616
rect 5121 12550 5286 12564
rect 5121 12537 5132 12550
rect 5081 12498 5132 12537
rect 5184 12498 5232 12550
rect 5284 12498 5286 12550
rect 5081 12464 5087 12498
rect 5121 12484 5286 12498
rect 5121 12464 5132 12484
rect 5081 12432 5132 12464
rect 5184 12432 5232 12484
rect 5284 12432 5286 12484
rect 5081 12425 5286 12432
rect 5081 12391 5087 12425
rect 5121 12418 5286 12425
rect 5121 12391 5132 12418
rect 5081 12366 5132 12391
rect 5184 12366 5232 12418
rect 5284 12366 5286 12418
rect 5081 12352 5286 12366
rect 7755 12387 7795 13836
rect 7835 13969 7887 13975
rect 7835 13905 7887 13917
rect 7835 13847 7887 13853
rect 7835 13836 7876 13847
tri 7876 13836 7887 13847 nw
rect 7835 12436 7875 13836
tri 7875 13835 7876 13836 nw
rect 9007 13687 9013 13739
rect 9065 13687 9077 13739
rect 9129 13687 9137 13739
tri 11889 13612 11892 13615 se
rect 11892 13612 11898 13615
rect 11680 13606 11898 13612
rect 11950 13606 11988 13615
rect 12040 13606 12078 13615
rect 11680 13572 11758 13606
rect 11792 13572 11841 13606
rect 11875 13572 11898 13606
rect 11958 13572 11988 13606
rect 12041 13572 12078 13606
rect 11680 13566 11898 13572
rect 11680 13563 11771 13566
tri 11771 13563 11774 13566 nw
tri 11889 13563 11892 13566 ne
rect 11892 13563 11898 13566
rect 11950 13563 11988 13572
rect 12040 13563 12078 13572
rect 12130 13563 12136 13615
rect 11680 13548 11756 13563
tri 11756 13548 11771 13563 nw
rect 11680 13533 11741 13548
tri 11741 13533 11756 13548 nw
rect 11680 13499 11686 13533
rect 11720 13499 11726 13533
tri 11726 13518 11741 13533 nw
rect 11680 13460 11726 13499
rect 11680 13426 11686 13460
rect 11720 13426 11726 13460
rect 11680 13387 11726 13426
rect 11680 13353 11686 13387
rect 11720 13353 11726 13387
rect 11680 13314 11726 13353
rect 11680 13280 11686 13314
rect 11720 13280 11726 13314
rect 11680 13241 11726 13280
rect 11680 13207 11686 13241
rect 11720 13207 11726 13241
rect 11680 13168 11726 13207
rect 11680 13134 11686 13168
rect 11720 13134 11726 13168
rect 11680 13095 11726 13134
rect 11680 13061 11686 13095
rect 11720 13061 11726 13095
rect 11680 13022 11726 13061
rect 11680 12988 11686 13022
rect 11720 12988 11726 13022
rect 11680 12949 11726 12988
rect 11680 12915 11686 12949
rect 11720 12915 11726 12949
rect 11680 12875 11726 12915
rect 11680 12841 11686 12875
rect 11720 12841 11726 12875
rect 11680 12801 11726 12841
rect 11680 12767 11686 12801
rect 11720 12767 11726 12801
rect 11680 12727 11726 12767
rect 11680 12693 11686 12727
rect 11720 12693 11726 12727
rect 11680 12653 11726 12693
rect 11680 12619 11686 12653
rect 11720 12619 11726 12653
rect 11680 12579 11726 12619
rect 11680 12545 11686 12579
rect 11720 12545 11726 12579
rect 11680 12505 11726 12545
rect 11680 12471 11686 12505
rect 11720 12471 11726 12505
tri 7835 12431 7840 12436 ne
rect 7840 12431 7875 12436
tri 7875 12431 7898 12454 sw
rect 11680 12431 11726 12471
tri 7840 12409 7862 12431 ne
rect 7862 12409 7898 12431
tri 7898 12409 7920 12431 sw
tri 9300 12409 9312 12421 se
rect 9312 12409 9318 12421
tri 7862 12397 7874 12409 ne
rect 7874 12397 9318 12409
tri 7874 12396 7875 12397 ne
rect 7875 12396 9318 12397
tri 7875 12390 7881 12396 ne
rect 7881 12390 9318 12396
tri 7795 12387 7798 12390 sw
tri 7881 12387 7884 12390 ne
rect 7884 12387 9318 12390
rect 7755 12383 7798 12387
tri 7798 12383 7802 12387 sw
tri 7884 12383 7888 12387 ne
rect 7888 12383 9318 12387
rect 7755 12372 7802 12383
tri 7755 12357 7770 12372 ne
rect 7770 12370 7802 12372
tri 7802 12370 7815 12383 sw
tri 7888 12370 7901 12383 ne
rect 7901 12370 9318 12383
rect 7770 12357 7815 12370
tri 7815 12357 7828 12370 sw
tri 7901 12369 7902 12370 ne
rect 7902 12369 9318 12370
rect 9370 12369 9382 12421
rect 9434 12369 9440 12421
rect 11680 12397 11686 12431
rect 11720 12397 11726 12431
tri 10853 12369 10854 12370 se
rect 10854 12369 11108 12370
tri 10841 12357 10853 12369 se
rect 10853 12357 11108 12369
rect 5081 12318 5087 12352
rect 5121 12318 5132 12352
rect 5081 12300 5132 12318
rect 5184 12300 5232 12352
rect 5284 12300 5286 12352
tri 7770 12350 7777 12357 ne
rect 7777 12350 7828 12357
tri 7828 12350 7835 12357 sw
tri 10834 12350 10841 12357 se
rect 10841 12350 11108 12357
tri 7777 12347 7780 12350 ne
rect 7780 12347 7835 12350
tri 7835 12347 7838 12350 sw
tri 10831 12347 10834 12350 se
rect 10834 12347 11108 12350
tri 7780 12329 7798 12347 ne
rect 7798 12329 7838 12347
tri 7838 12329 7856 12347 sw
tri 10813 12329 10831 12347 se
rect 10831 12329 11108 12347
tri 7798 12323 7804 12329 ne
rect 7804 12323 9444 12329
tri 10807 12323 10813 12329 se
rect 10813 12323 11108 12329
tri 7804 12313 7814 12323 ne
rect 7814 12313 9392 12323
tri 7814 12311 7816 12313 ne
rect 7816 12311 9392 12313
rect 5081 12286 5286 12300
tri 7816 12289 7838 12311 ne
rect 7838 12289 9392 12311
rect 5081 12279 5132 12286
rect 5081 12245 5087 12279
rect 5121 12245 5132 12279
rect 5081 12234 5132 12245
rect 5184 12234 5232 12286
rect 5284 12234 5286 12286
rect 5081 12220 5286 12234
rect 5081 12206 5132 12220
rect 4983 12189 5035 12195
tri 3732 12130 3734 12132 sw
rect 4364 12130 4416 12136
tri 4625 12130 4626 12131 se
rect 4626 12130 4672 12145
rect 3686 12119 3734 12130
tri 3734 12119 3745 12130 sw
tri 4614 12119 4625 12130 se
rect 4625 12119 4672 12130
rect 3686 12117 3745 12119
tri 3745 12117 3747 12119 sw
tri 4612 12117 4614 12119 se
rect 4614 12117 4672 12119
rect 3686 12116 3747 12117
tri 3747 12116 3748 12117 sw
tri 4611 12116 4612 12117 se
rect 4612 12116 4672 12117
rect 3686 12112 3748 12116
tri 3748 12112 3752 12116 sw
tri 4607 12112 4611 12116 se
rect 4611 12112 4672 12116
tri 3686 12110 3688 12112 ne
rect 3688 12110 3752 12112
tri 3752 12110 3754 12112 sw
tri 4605 12110 4607 12112 se
rect 4607 12110 4672 12112
tri 3688 12097 3701 12110 ne
rect 3701 12097 3754 12110
tri 3754 12097 3767 12110 sw
tri 4592 12097 4605 12110 se
rect 4605 12097 4672 12110
tri 3701 12076 3722 12097 ne
rect 3722 12076 4672 12097
tri 3722 12067 3731 12076 ne
rect 3731 12067 4672 12076
rect 5081 12172 5087 12206
rect 5121 12172 5132 12206
rect 5081 12168 5132 12172
rect 5184 12168 5232 12220
rect 5284 12168 5286 12220
tri 10795 12311 10807 12323 se
rect 10807 12318 11108 12323
rect 11160 12318 11172 12370
rect 11224 12318 11230 12370
rect 11680 12357 11726 12397
rect 11680 12323 11686 12357
rect 11720 12323 11726 12357
rect 10807 12311 10869 12318
tri 10869 12311 10876 12318 nw
tri 10780 12296 10795 12311 se
rect 10795 12296 10854 12311
tri 10854 12296 10869 12311 nw
tri 10767 12283 10780 12296 se
rect 10780 12283 10841 12296
tri 10841 12283 10854 12296 nw
rect 11680 12283 11726 12323
rect 9392 12259 9444 12271
tri 10733 12249 10767 12283 se
rect 10767 12249 10807 12283
tri 10807 12249 10841 12283 nw
rect 11680 12249 11686 12283
rect 11720 12249 11726 12283
rect 11868 13418 12106 13424
rect 11868 13384 11880 13418
rect 11914 13384 11952 13418
rect 11986 13384 12024 13418
rect 12058 13384 12106 13418
rect 11868 13378 12106 13384
rect 11868 13353 12020 13378
tri 12020 13353 12045 13378 nw
rect 11868 13319 12010 13353
tri 12010 13343 12020 13353 nw
rect 11868 13285 11874 13319
rect 11908 13285 12010 13319
rect 11868 13247 12010 13285
rect 11868 13213 11874 13247
rect 11908 13213 12010 13247
rect 11868 13175 12010 13213
rect 11868 13141 11874 13175
rect 11908 13141 12010 13175
rect 11868 13103 12010 13141
rect 11868 13069 11874 13103
rect 11908 13069 12010 13103
rect 11868 13031 12010 13069
rect 11868 12997 11874 13031
rect 11908 12997 12010 13031
rect 11868 12959 12010 12997
rect 11868 12925 11874 12959
rect 11908 12925 12010 12959
rect 11868 12887 12010 12925
rect 11868 12853 11874 12887
rect 11908 12853 12010 12887
rect 11868 12815 12010 12853
rect 11868 12781 11874 12815
rect 11908 12781 12010 12815
rect 11868 12743 12010 12781
rect 11868 12709 11874 12743
rect 11908 12709 12010 12743
rect 11868 12671 12010 12709
rect 11868 12637 11874 12671
rect 11908 12637 12010 12671
rect 11868 12599 12010 12637
rect 11868 12565 11874 12599
rect 11908 12565 12010 12599
rect 11868 12527 12010 12565
rect 11868 12493 11874 12527
rect 11908 12493 12010 12527
rect 12220 13247 12266 14450
tri 12969 14416 13003 14450 se
rect 13003 14416 13035 14450
tri 13035 14416 13069 14450 nw
tri 12965 14412 12969 14416 se
rect 12969 14412 13031 14416
tri 13031 14412 13035 14416 nw
tri 12931 14378 12965 14412 se
rect 12965 14378 12997 14412
tri 12997 14378 13031 14412 nw
rect 13458 14390 13510 14415
tri 12903 14350 12931 14378 se
rect 12931 14350 12969 14378
tri 12969 14350 12997 14378 nw
tri 12893 14340 12903 14350 se
rect 12903 14340 12959 14350
tri 12959 14340 12969 14350 nw
tri 12859 14306 12893 14340 se
rect 12893 14306 12925 14340
tri 12925 14306 12959 14340 nw
rect 13458 14312 13510 14338
tri 12837 14284 12859 14306 se
rect 12859 14284 12903 14306
tri 12903 14284 12925 14306 nw
tri 12821 14268 12837 14284 se
rect 12837 14268 12887 14284
tri 12887 14268 12903 14284 nw
tri 12787 14234 12821 14268 se
rect 12821 14234 12853 14268
tri 12853 14234 12887 14268 nw
rect 13458 14234 13510 14260
tri 12771 14218 12787 14234 se
rect 12787 14218 12837 14234
tri 12837 14218 12853 14234 nw
tri 12749 14196 12771 14218 se
rect 12771 14196 12815 14218
tri 12815 14196 12837 14218 nw
tri 12715 14162 12749 14196 se
rect 12749 14162 12781 14196
tri 12781 14162 12815 14196 nw
tri 12705 14152 12715 14162 se
rect 12715 14152 12771 14162
tri 12771 14152 12781 14162 nw
rect 13458 14156 13510 14182
tri 12677 14124 12705 14152 se
rect 12705 14124 12743 14152
tri 12743 14124 12771 14152 nw
tri 12643 14090 12677 14124 se
rect 12677 14090 12709 14124
tri 12709 14090 12743 14124 nw
tri 12639 14086 12643 14090 se
rect 12643 14086 12705 14090
tri 12705 14086 12709 14090 nw
tri 12605 14052 12639 14086 se
rect 12639 14052 12671 14086
tri 12671 14052 12705 14086 nw
tri 12573 14020 12605 14052 se
rect 12605 14020 12639 14052
tri 12639 14020 12671 14052 nw
tri 12571 14018 12573 14020 se
rect 12573 14018 12637 14020
tri 12637 14018 12639 14020 nw
tri 12533 13980 12571 14018 se
rect 12571 13980 12599 14018
tri 12599 13980 12637 14018 nw
tri 12507 13954 12533 13980 se
rect 12533 13954 12573 13980
tri 12573 13954 12599 13980 nw
tri 12499 13946 12507 13954 se
rect 12507 13946 12565 13954
tri 12565 13946 12573 13954 nw
rect 12220 13213 12226 13247
rect 12260 13213 12266 13247
rect 12220 13170 12266 13213
rect 12220 13136 12226 13170
rect 12260 13136 12266 13170
rect 12220 13093 12266 13136
rect 12220 13059 12226 13093
rect 12260 13059 12266 13093
rect 12220 13016 12266 13059
rect 12220 12982 12226 13016
rect 12260 12982 12266 13016
rect 12220 12939 12266 12982
rect 12220 12905 12226 12939
rect 12260 12905 12266 12939
rect 12220 12862 12266 12905
rect 12220 12828 12226 12862
rect 12260 12828 12266 12862
rect 12220 12785 12266 12828
rect 12220 12751 12226 12785
rect 12260 12751 12266 12785
rect 12220 12708 12266 12751
rect 12220 12674 12226 12708
rect 12260 12674 12266 12708
rect 12220 12631 12266 12674
rect 12220 12597 12226 12631
rect 12260 12597 12266 12631
rect 12220 12554 12266 12597
rect 12220 12520 12226 12554
rect 12260 12520 12266 12554
rect 12220 12508 12266 12520
tri 12476 13923 12499 13946 se
rect 12499 13923 12542 13946
tri 12542 13923 12565 13946 nw
rect 12476 13908 12527 13923
tri 12527 13908 12542 13923 nw
rect 12476 13426 12522 13908
tri 12522 13903 12527 13908 nw
rect 12553 13563 12559 13615
rect 12611 13606 12648 13615
rect 12700 13612 12706 13615
tri 12706 13612 12709 13615 sw
rect 12700 13606 12831 13612
rect 12611 13572 12642 13606
rect 12700 13572 12719 13606
rect 12753 13572 12831 13606
rect 12611 13563 12648 13572
rect 12700 13563 12831 13572
tri 12740 13548 12755 13563 ne
rect 12755 13548 12831 13563
tri 12755 13533 12770 13548 ne
rect 12770 13533 12831 13548
tri 12770 13518 12785 13533 ne
rect 12785 13499 12791 13533
rect 12825 13499 12831 13533
rect 12785 13460 12831 13499
tri 12522 13426 12555 13459 sw
rect 12785 13426 12791 13460
rect 12825 13426 12831 13460
rect 12476 13424 12555 13426
tri 12555 13424 12557 13426 sw
rect 12476 13418 12640 13424
rect 12476 13384 12522 13418
rect 12556 13384 12594 13418
rect 12628 13384 12640 13418
rect 12476 13340 12640 13384
rect 12476 13306 12600 13340
rect 12634 13306 12640 13340
rect 12476 13268 12640 13306
rect 12476 13234 12600 13268
rect 12634 13234 12640 13268
rect 12476 13196 12640 13234
rect 12476 13162 12600 13196
rect 12634 13162 12640 13196
rect 12476 13124 12640 13162
rect 12476 13090 12600 13124
rect 12634 13090 12640 13124
rect 12476 13052 12640 13090
rect 12476 13018 12600 13052
rect 12634 13018 12640 13052
rect 12476 12980 12640 13018
rect 12476 12946 12600 12980
rect 12634 12946 12640 12980
rect 12476 12908 12640 12946
rect 12476 12874 12600 12908
rect 12634 12874 12640 12908
rect 12476 12836 12640 12874
rect 12476 12802 12600 12836
rect 12634 12802 12640 12836
rect 12476 12764 12640 12802
rect 12476 12730 12600 12764
rect 12634 12730 12640 12764
rect 12476 12692 12640 12730
rect 12476 12658 12600 12692
rect 12634 12658 12640 12692
rect 12476 12620 12640 12658
rect 12476 12586 12600 12620
rect 12634 12586 12640 12620
rect 12476 12548 12640 12586
rect 12476 12514 12600 12548
rect 12634 12514 12640 12548
rect 11868 12455 12010 12493
rect 11868 12421 11874 12455
rect 11908 12442 12010 12455
rect 12476 12476 12640 12514
tri 12010 12442 12018 12450 sw
tri 12468 12442 12476 12450 se
rect 12476 12442 12600 12476
rect 12634 12442 12640 12476
rect 11908 12435 12018 12442
tri 12018 12435 12025 12442 sw
tri 12461 12435 12468 12442 se
rect 12468 12435 12640 12442
rect 11908 12421 12025 12435
rect 11868 12415 12025 12421
tri 12025 12415 12045 12435 sw
tri 12441 12415 12461 12435 se
rect 12461 12415 12640 12435
rect 11868 12404 12640 12415
rect 11868 12383 12600 12404
rect 11868 12349 11874 12383
rect 11908 12370 12600 12383
rect 12634 12370 12640 12404
rect 11908 12349 12640 12370
rect 11868 12332 12640 12349
rect 11868 12311 12600 12332
rect 11868 12277 11874 12311
rect 11908 12298 12600 12311
rect 12634 12298 12640 12332
rect 11908 12277 12640 12298
rect 11868 12265 12640 12277
tri 12440 12260 12445 12265 ne
rect 12445 12260 12640 12265
tri 10721 12237 10733 12249 se
rect 10733 12237 10795 12249
tri 10795 12237 10807 12249 nw
tri 10717 12233 10721 12237 se
rect 10721 12233 10791 12237
tri 10791 12233 10795 12237 nw
tri 10710 12226 10717 12233 se
rect 10717 12226 10784 12233
tri 10784 12226 10791 12233 nw
rect 10958 12232 11010 12238
rect 11680 12237 11726 12249
tri 12445 12237 12468 12260 ne
rect 12468 12237 12600 12260
tri 12468 12233 12472 12237 ne
rect 12472 12233 12600 12237
tri 10706 12222 10710 12226 se
rect 10710 12222 10780 12226
tri 10780 12222 10784 12226 nw
tri 10697 12213 10706 12222 se
rect 10706 12213 10771 12222
tri 10771 12213 10780 12222 nw
rect 9392 12201 9444 12207
tri 10685 12201 10697 12213 se
rect 10697 12201 10757 12213
tri 10683 12199 10685 12201 se
rect 10685 12199 10757 12201
tri 10757 12199 10771 12213 nw
tri 10677 12193 10683 12199 se
rect 10683 12193 10751 12199
tri 10751 12193 10757 12199 nw
rect 5081 12160 5286 12168
tri 10644 12160 10677 12193 se
rect 10677 12160 10717 12193
tri 10643 12159 10644 12160 se
rect 10644 12159 10717 12160
tri 10717 12159 10751 12193 nw
tri 11010 12226 11017 12233 sw
tri 12472 12229 12476 12233 ne
rect 12476 12226 12600 12233
rect 12634 12226 12640 12260
rect 11010 12213 11017 12226
tri 11017 12213 11030 12226 sw
rect 11010 12199 11030 12213
tri 11030 12199 11044 12213 sw
rect 11010 12193 12436 12199
rect 11010 12180 12062 12193
rect 10958 12168 12062 12180
tri 10638 12154 10643 12159 se
rect 10643 12154 10712 12159
tri 10712 12154 10717 12159 nw
tri 10637 12153 10638 12154 se
rect 10638 12153 10711 12154
tri 10711 12153 10712 12154 nw
tri 10636 12152 10637 12153 se
rect 10637 12152 10706 12153
tri 5035 12148 5039 12152 sw
tri 10632 12148 10636 12152 se
rect 10636 12148 10706 12152
tri 10706 12148 10711 12153 nw
rect 5035 12139 5039 12148
tri 5039 12139 5048 12148 sw
tri 10623 12139 10632 12148 se
rect 10632 12139 10697 12148
tri 10697 12139 10706 12148 nw
rect 5035 12137 5048 12139
rect 4983 12131 5048 12137
tri 5048 12131 5056 12139 sw
tri 10615 12131 10623 12139 se
rect 10623 12131 10677 12139
rect 4983 12125 5056 12131
rect 5035 12119 5056 12125
tri 5056 12119 5068 12131 sw
tri 10603 12119 10615 12131 se
rect 10615 12119 10677 12131
tri 10677 12119 10697 12139 nw
rect 5035 12116 10674 12119
tri 10674 12116 10677 12119 nw
rect 11010 12159 12062 12168
rect 12096 12159 12134 12193
rect 12168 12159 12318 12193
rect 12352 12159 12390 12193
rect 12424 12159 12436 12193
rect 11010 12153 12436 12159
rect 12476 12188 12640 12226
rect 12476 12154 12600 12188
rect 12634 12154 12640 12188
rect 11010 12139 11030 12153
tri 11030 12139 11044 12153 nw
tri 12464 12139 12476 12151 se
rect 12476 12139 12640 12154
tri 11010 12119 11030 12139 nw
tri 12444 12119 12464 12139 se
rect 12464 12119 12640 12139
tri 12441 12116 12444 12119 se
rect 12444 12116 12640 12119
rect 5035 12110 10668 12116
tri 10668 12110 10674 12116 nw
rect 10958 12110 11010 12116
rect 11874 12110 12600 12116
rect 5035 12097 10655 12110
tri 10655 12097 10668 12110 nw
rect 5035 12083 10641 12097
tri 10641 12083 10655 12097 nw
rect 5035 12076 10634 12083
tri 10634 12076 10641 12083 nw
rect 11874 12076 11886 12110
rect 11920 12076 11958 12110
rect 11992 12076 12030 12110
rect 12064 12076 12102 12110
rect 12136 12076 12174 12110
rect 12208 12076 12246 12110
rect 12280 12076 12318 12110
rect 12352 12076 12390 12110
rect 12424 12076 12462 12110
rect 12496 12082 12600 12110
rect 12634 12082 12640 12116
rect 12785 13387 12831 13426
rect 12785 13353 12791 13387
rect 12825 13353 12831 13387
rect 12785 13314 12831 13353
rect 12785 13280 12791 13314
rect 12825 13280 12831 13314
rect 12785 13241 12831 13280
rect 12785 13207 12791 13241
rect 12825 13207 12831 13241
rect 12785 13168 12831 13207
rect 12785 13134 12791 13168
rect 12825 13134 12831 13168
rect 12785 13095 12831 13134
rect 12785 13061 12791 13095
rect 12825 13061 12831 13095
rect 12785 13022 12831 13061
rect 12785 12988 12791 13022
rect 12825 12988 12831 13022
rect 12785 12949 12831 12988
rect 12785 12915 12791 12949
rect 12825 12915 12831 12949
rect 12785 12876 12831 12915
rect 12785 12842 12791 12876
rect 12825 12842 12831 12876
rect 12785 12803 12831 12842
rect 12785 12769 12791 12803
rect 12825 12769 12831 12803
rect 12785 12730 12831 12769
rect 12785 12696 12791 12730
rect 12825 12696 12831 12730
rect 12785 12657 12831 12696
rect 12785 12623 12791 12657
rect 12825 12623 12831 12657
rect 12785 12583 12831 12623
rect 12785 12549 12791 12583
rect 12825 12549 12831 12583
rect 12785 12509 12831 12549
rect 12785 12475 12791 12509
rect 12825 12475 12831 12509
rect 12785 12435 12831 12475
rect 12785 12401 12791 12435
rect 12825 12401 12831 12435
rect 12785 12361 12831 12401
rect 12785 12327 12791 12361
rect 12825 12327 12831 12361
rect 12785 12287 12831 12327
rect 12785 12253 12791 12287
rect 12825 12253 12831 12287
rect 12785 12213 12831 12253
rect 12785 12179 12791 12213
rect 12825 12179 12831 12213
rect 13458 13404 13510 14104
tri 13843 13409 13846 13412 se
rect 13846 13409 13892 14531
tri 13892 14506 13917 14531 nw
tri 14069 14506 14094 14531 ne
rect 13970 14455 14022 14473
rect 13970 14387 14022 14403
rect 13970 14319 14022 14335
rect 13970 14251 14022 14267
rect 13970 14183 14022 14199
rect 13970 14115 14022 14131
rect 13970 14047 14022 14063
rect 13970 13978 14022 13995
rect 13970 13909 14022 13926
tri 13892 13409 13895 13412 sw
tri 13510 13404 13515 13409 sw
tri 13838 13404 13843 13409 se
rect 13843 13404 13895 13409
tri 13895 13404 13900 13409 sw
rect 13458 13375 13515 13404
tri 13515 13375 13544 13404 sw
tri 13812 13378 13838 13404 se
rect 13838 13378 13900 13404
tri 13900 13378 13926 13404 sw
rect 13458 13369 13674 13375
rect 13458 13335 13556 13369
rect 13590 13335 13628 13369
rect 13662 13335 13674 13369
rect 13458 13329 13674 13335
rect 13800 13369 13930 13378
rect 13800 13335 13812 13369
rect 13846 13335 13884 13369
rect 13918 13335 13930 13369
rect 13458 13298 13513 13329
tri 13513 13298 13544 13329 nw
rect 13800 13326 13930 13335
tri 13812 13298 13840 13326 ne
rect 13840 13298 13898 13326
tri 13898 13298 13926 13326 nw
rect 13458 12206 13510 13298
tri 13510 13295 13513 13298 nw
tri 13840 13295 13843 13298 ne
rect 13843 13295 13895 13298
tri 13895 13295 13898 13298 nw
tri 13843 13292 13846 13295 ne
tri 13844 12209 13846 12211 se
rect 13846 12209 13892 13295
tri 13892 13292 13895 13295 nw
rect 13970 13233 14022 13857
tri 14086 13404 14094 13412 se
rect 14094 13409 14140 14531
tri 14140 14506 14165 14531 nw
rect 14230 14473 14276 14614
rect 14486 14666 14695 14693
rect 14486 14632 14655 14666
rect 14689 14632 14695 14666
rect 14486 14565 14695 14632
rect 14486 14531 14655 14565
rect 14689 14531 14695 14565
rect 14486 14484 14695 14531
rect 14486 14450 14655 14484
rect 14689 14450 14695 14484
rect 14486 14412 14695 14450
rect 14486 14378 14655 14412
rect 14689 14378 14695 14412
rect 14486 14340 14695 14378
rect 14486 14306 14655 14340
rect 14689 14306 14695 14340
rect 14486 14268 14695 14306
rect 14486 14234 14655 14268
rect 14689 14234 14695 14268
rect 14486 14196 14695 14234
rect 14486 14162 14655 14196
rect 14689 14162 14695 14196
rect 14486 14124 14695 14162
rect 14486 14090 14655 14124
rect 14689 14090 14695 14124
rect 14486 14052 14695 14090
rect 14486 14018 14655 14052
rect 14689 14018 14695 14052
rect 14486 13980 14695 14018
rect 14486 13946 14655 13980
rect 14689 13946 14695 13980
rect 14486 13908 14695 13946
rect 14486 13874 14655 13908
rect 14689 13874 14695 13908
rect 14486 13836 14695 13874
rect 14486 13802 14655 13836
rect 14689 13802 14695 13836
rect 14486 13764 14695 13802
rect 14486 13730 14655 13764
rect 14689 13730 14695 13764
rect 14486 13692 14695 13730
rect 14486 13658 14655 13692
rect 14689 13658 14695 13692
rect 14486 13620 14695 13658
rect 14486 13586 14655 13620
rect 14689 13586 14695 13620
rect 14486 13548 14695 13586
rect 14486 13514 14655 13548
rect 14689 13514 14695 13548
rect 14486 13476 14695 13514
rect 14486 13442 14655 13476
rect 14689 13442 14695 13476
tri 14140 13409 14143 13412 sw
rect 14094 13404 14143 13409
tri 14143 13404 14148 13409 sw
tri 14481 13404 14486 13409 se
rect 14486 13404 14695 13442
tri 14060 13378 14086 13404 se
rect 14086 13378 14148 13404
tri 14148 13378 14174 13404 sw
tri 14455 13378 14481 13404 se
rect 14481 13378 14655 13404
rect 14056 13369 14186 13378
tri 14452 13375 14455 13378 se
rect 14455 13375 14655 13378
rect 14056 13335 14068 13369
rect 14102 13335 14140 13369
rect 14174 13335 14186 13369
rect 14056 13326 14186 13335
rect 14312 13370 14655 13375
rect 14689 13370 14695 13404
rect 14312 13369 14695 13370
rect 14312 13335 14324 13369
rect 14358 13335 14396 13369
rect 14430 13335 14695 13369
rect 14312 13332 14695 13335
rect 14312 13329 14655 13332
tri 14452 13326 14455 13329 ne
rect 14455 13326 14655 13329
tri 14060 13298 14088 13326 ne
rect 14088 13298 14146 13326
tri 14146 13298 14174 13326 nw
tri 14455 13298 14483 13326 ne
rect 14483 13298 14655 13326
rect 14689 13298 14695 13332
tri 14088 13292 14094 13298 ne
rect 14094 13295 14143 13298
tri 14143 13295 14146 13298 nw
tri 14483 13295 14486 13298 ne
tri 13970 13229 13974 13233 ne
rect 13974 13109 14020 13233
tri 14020 13231 14022 13233 nw
tri 13972 12237 13974 12239 se
tri 13970 12235 13972 12237 se
rect 13972 12235 13974 12237
tri 14020 12235 14022 12237 sw
tri 13892 12209 13894 12211 sw
tri 13841 12206 13844 12209 se
rect 13844 12206 13894 12209
tri 13894 12206 13897 12209 sw
rect 13970 12206 14022 12235
tri 14092 12209 14094 12211 se
rect 14094 12209 14140 13295
tri 14140 13292 14143 13295 nw
rect 14486 13260 14695 13298
rect 14486 13226 14655 13260
rect 14689 13226 14695 13260
rect 14486 13188 14695 13226
rect 14486 13154 14655 13188
rect 14689 13154 14695 13188
rect 14486 13116 14695 13154
rect 14486 13082 14655 13116
rect 14689 13082 14695 13116
rect 14486 13044 14695 13082
rect 14486 13010 14655 13044
rect 14689 13010 14695 13044
rect 14486 12972 14695 13010
rect 14486 12938 14655 12972
rect 14689 12938 14695 12972
rect 14486 12900 14695 12938
rect 14486 12866 14655 12900
rect 14689 12866 14695 12900
rect 14486 12827 14695 12866
rect 14486 12793 14655 12827
rect 14689 12793 14695 12827
rect 14486 12754 14695 12793
rect 14486 12720 14655 12754
rect 14689 12720 14695 12754
rect 14486 12681 14695 12720
rect 14486 12647 14655 12681
rect 14689 12647 14695 12681
rect 14486 12608 14695 12647
rect 14486 12574 14655 12608
rect 14689 12574 14695 12608
rect 14486 12535 14695 12574
rect 14486 12501 14655 12535
rect 14689 12501 14695 12535
rect 14486 12462 14695 12501
rect 14486 12428 14655 12462
rect 14689 12428 14695 12462
rect 14486 12389 14695 12428
rect 14486 12355 14655 12389
rect 14689 12355 14695 12389
rect 14486 12316 14695 12355
rect 14486 12282 14655 12316
rect 14689 12282 14695 12316
rect 14486 12243 14695 12282
tri 14140 12209 14142 12211 sw
rect 14486 12209 14655 12243
rect 14689 12209 14695 12243
tri 14089 12206 14092 12209 se
rect 14092 12206 14142 12209
tri 14142 12206 14145 12209 sw
rect 12785 12139 12831 12179
rect 12785 12105 12791 12139
rect 12825 12105 12831 12139
rect 12785 12093 12831 12105
rect 13718 12097 13764 12206
tri 13812 12177 13841 12206 se
rect 13841 12177 13897 12206
tri 13897 12177 13926 12206 sw
tri 14060 12177 14089 12206 se
rect 14089 12177 14145 12206
tri 14145 12177 14174 12206 sw
rect 13804 12168 14190 12177
rect 13804 12134 13816 12168
rect 13850 12134 13888 12168
rect 13922 12134 14072 12168
rect 14106 12134 14144 12168
rect 14178 12134 14190 12168
rect 13804 12125 14190 12134
tri 13764 12097 13791 12124 sw
tri 14203 12097 14230 12124 se
rect 14230 12097 14276 12206
rect 13718 12093 13791 12097
tri 13791 12093 13795 12097 sw
tri 14199 12093 14203 12097 se
rect 14203 12093 14276 12097
rect 12496 12076 12640 12082
rect 5035 12073 10628 12076
rect 4983 12070 10628 12073
tri 10628 12070 10634 12076 nw
rect 11874 12070 12640 12076
rect 13718 12090 13795 12093
tri 13795 12090 13798 12093 sw
tri 14196 12090 14199 12093 se
rect 14199 12090 14276 12093
rect 4983 12067 10625 12070
tri 10625 12067 10628 12070 nw
tri 3731 12063 3735 12067 ne
rect 3735 12063 4672 12067
tri 3735 12051 3747 12063 ne
rect 3747 12051 4672 12063
rect 13718 12044 14276 12090
rect 14486 12170 14695 12209
rect 14486 12136 14655 12170
rect 14689 12136 14695 12170
rect 14486 12097 14695 12136
rect 14486 12063 14655 12097
rect 14689 12063 14695 12097
rect 14486 12051 14695 12063
tri 13913 12027 13930 12044 ne
rect 13930 12027 14006 12044
tri 4829 12021 4835 12027 se
rect 4835 12021 10737 12027
tri 13930 12021 13936 12027 ne
rect 13936 12021 14006 12027
rect 4450 12015 10685 12021
rect 4450 11981 4462 12015
rect 4496 11981 4534 12015
rect 4568 11981 4718 12015
rect 4752 11981 4790 12015
rect 4824 11981 10685 12015
rect 4450 11975 10685 11981
tri 10651 11947 10679 11975 ne
rect 10679 11969 10685 11975
tri 13936 12010 13947 12021 ne
rect 11196 11993 13664 11999
tri 10737 11974 10738 11975 nw
rect 10679 11957 10737 11969
rect 10679 11947 10685 11957
tri 10679 11944 10682 11947 ne
rect 10682 11944 10685 11947
rect 3850 11892 4065 11944
rect 4117 11892 4129 11944
rect 4181 11892 7280 11944
rect 7332 11892 7344 11944
rect 7396 11892 7402 11944
tri 10682 11941 10685 11944 ne
rect 8648 11897 8700 11903
rect 10685 11899 10737 11905
rect 11248 11947 13664 11993
rect 13716 11947 13728 11999
rect 13780 11947 13786 11999
rect 11248 11941 11267 11947
rect 11196 11932 11267 11941
tri 11267 11932 11282 11947 nw
rect 11196 11929 11248 11932
tri 3616 11821 3650 11855 sw
tri 8614 11821 8648 11855 se
tri 11248 11913 11267 11932 nw
tri 13928 11913 13947 11932 se
rect 13947 11913 14006 12021
tri 14006 12010 14040 12044 nw
tri 13913 11898 13928 11913 se
rect 13928 11898 14006 11913
rect 11196 11871 11248 11877
tri 12132 11871 12159 11898 se
rect 12159 11871 14006 11898
tri 12116 11855 12132 11871 se
rect 12132 11855 14006 11871
tri 8700 11852 8703 11855 sw
tri 12113 11852 12116 11855 se
rect 12116 11852 14006 11855
rect 8700 11845 8703 11852
rect 8648 11841 8703 11845
tri 8703 11841 8714 11852 sw
tri 12102 11841 12113 11852 se
rect 12113 11841 12168 11852
tri 12168 11841 12179 11852 nw
rect 8648 11833 8714 11841
rect 3570 11781 8648 11821
rect 8700 11821 8714 11833
tri 8714 11821 8734 11841 sw
tri 12082 11821 12102 11841 se
rect 8700 11781 12102 11821
rect 3570 11775 12102 11781
tri 12102 11775 12168 11841 nw
tri 552 11700 586 11734 sw
tri 4389 11700 4395 11706 se
rect 4395 11700 4401 11706
rect 506 11654 4401 11700
rect 4453 11654 4465 11706
rect 4517 11654 4523 11706
rect 10958 11672 11010 11678
tri 10924 11595 10958 11629 se
rect 10958 11608 11010 11620
tri 5617 11553 5659 11595 se
rect 5659 11556 10958 11595
rect 5659 11553 11010 11556
rect 11196 11589 11248 11595
tri 5601 11537 5617 11553 se
rect 5617 11549 11010 11553
tri 11192 11549 11196 11553 se
rect 5617 11537 5659 11549
tri 5659 11537 5671 11549 nw
tri 11180 11537 11192 11549 se
rect 11192 11537 11196 11549
tri 5583 11519 5601 11537 se
rect 5601 11519 5641 11537
tri 5641 11519 5659 11537 nw
tri 11162 11519 11180 11537 se
rect 11180 11525 11248 11537
rect 11180 11519 11196 11525
tri 5543 11479 5583 11519 se
rect 5583 11479 5601 11519
tri 5601 11479 5641 11519 nw
tri 5659 11479 5699 11519 se
rect 5699 11479 11196 11519
tri 5486 11422 5543 11479 se
rect 5543 11461 5583 11479
tri 5583 11461 5601 11479 nw
tri 5641 11461 5659 11479 se
rect 5659 11473 11196 11479
rect 5659 11467 11248 11473
rect 5659 11461 5699 11467
tri 5699 11461 5705 11467 nw
rect 5543 11422 5544 11461
tri 5544 11422 5583 11461 nw
tri 5602 11422 5641 11461 se
tri 5470 9919 5486 9935 se
rect 5486 9919 5526 11422
tri 5526 11404 5544 11422 nw
tri 5584 11404 5602 11422 se
rect 5602 11404 5641 11422
tri 5583 11403 5584 11404 se
rect 5584 11403 5641 11404
tri 5641 11403 5699 11461 nw
rect -201 9913 -149 9919
tri 5452 9901 5470 9919 se
rect 5470 9917 5526 9919
rect 5470 9901 5510 9917
tri 5510 9901 5526 9917 nw
tri 5566 11386 5583 11403 se
rect 5583 11386 5624 11403
tri 5624 11386 5641 11403 nw
tri 5428 9877 5452 9901 se
rect 5452 9899 5508 9901
tri 5508 9899 5510 9901 nw
rect 5452 9877 5486 9899
tri 5486 9877 5508 9899 nw
tri 5544 9877 5566 9899 se
rect 5566 9881 5606 11386
tri 5606 11368 5624 11386 nw
tri 10929 10634 10963 10668 nw
tri 11005 10634 11039 10668 ne
rect 10958 10550 11010 10556
rect 10958 10471 11010 10498
rect 10958 10413 11010 10419
tri 10929 10303 10962 10336 sw
tri 11006 10303 11039 10336 se
rect 9965 10257 10025 10303
rect 10929 10302 10962 10303
tri 10962 10302 10963 10303 sw
tri 11005 10302 11006 10303 se
rect 11006 10302 11039 10303
tri 10895 10268 10929 10302 ne
tri 10467 10222 10501 10256 ne
tri 10547 10222 10581 10256 nw
tri 5698 9982 5732 10016 nw
tri 10467 9901 10501 9935 se
tri 10547 9901 10581 9935 sw
rect 5566 9877 5580 9881
tri 5413 9862 5428 9877 se
rect 5428 9862 5464 9877
rect -201 9855 -149 9861
tri -149 9855 -142 9862 sw
tri 5406 9855 5413 9862 se
rect 5413 9855 5464 9862
tri 5464 9855 5486 9877 nw
tri 5522 9855 5544 9877 se
rect 5544 9855 5580 9877
tri 5580 9855 5606 9881 nw
rect -201 9849 -142 9855
rect -149 9831 -142 9849
tri -142 9831 -118 9855 sw
tri 5382 9831 5406 9855 se
rect 5406 9841 5450 9855
tri 5450 9841 5464 9855 nw
tri 5508 9841 5522 9855 se
rect 5522 9841 5566 9855
tri 5566 9841 5580 9855 nw
tri 11263 9841 11277 9855 ne
rect 11277 9841 11297 9855
rect 5406 9831 5440 9841
tri 5440 9831 5450 9841 nw
tri 5498 9831 5508 9841 se
rect 5508 9831 5546 9841
rect -149 9821 5430 9831
tri 5430 9821 5440 9831 nw
tri 5488 9821 5498 9831 se
rect 5498 9821 5546 9831
tri 5546 9821 5566 9841 nw
tri 11277 9821 11297 9841 ne
rect -149 9797 5400 9821
rect -201 9791 5400 9797
tri 5400 9791 5430 9821 nw
tri 5458 9791 5488 9821 se
rect 5488 9791 5508 9821
tri 5450 9783 5458 9791 se
rect 5458 9783 5508 9791
tri 5508 9783 5546 9821 nw
tri 5418 9751 5450 9783 se
rect 5450 9751 5476 9783
tri 5476 9751 5508 9783 nw
rect -327 9699 -321 9751
rect -269 9699 -257 9751
rect -205 9711 5436 9751
tri 5436 9711 5476 9751 nw
rect -205 9699 -199 9711
tri -199 9699 -187 9711 nw
tri 11343 9515 11377 9549 sw
tri 12235 9515 12240 9520 se
tri 5618 9391 5652 9425 se
rect 12240 8711 12246 8763
rect 12298 8711 12318 8763
rect 12370 8711 12390 8763
rect 12442 8711 12462 8763
rect 12514 8711 12534 8763
rect 12586 8711 12592 8763
rect 7478 8210 10615 8262
rect 10667 8210 10679 8262
rect 10731 8210 10737 8262
tri 6349 8132 6383 8166 se
tri 6435 8132 6469 8166 sw
tri 8607 8037 8610 8040 se
rect 8610 8037 8616 8040
rect 8209 8031 8616 8037
rect 8668 8031 8680 8040
rect 8732 8037 8738 8040
tri 8738 8037 8741 8040 sw
rect 8732 8031 12340 8037
rect 8209 7997 8221 8031
rect 8255 7997 8294 8031
rect 8328 7997 8367 8031
rect 8401 7997 8440 8031
rect 8474 7997 8513 8031
rect 8547 7997 8586 8031
rect 8766 7997 8805 8031
rect 8839 7997 8878 8031
rect 8912 7997 8951 8031
rect 8985 7997 9024 8031
rect 9058 7997 9097 8031
rect 9131 7997 9170 8031
rect 9204 7997 9243 8031
rect 9277 7997 9316 8031
rect 9350 7997 9389 8031
rect 9423 7997 9462 8031
rect 9496 7997 9535 8031
rect 9569 7997 9608 8031
rect 9642 7997 9681 8031
rect 9715 7997 9754 8031
rect 9788 7997 9827 8031
rect 9861 7997 9900 8031
rect 9934 7997 9973 8031
rect 10007 7997 10046 8031
rect 10080 7997 10119 8031
rect 10153 7997 10192 8031
rect 10226 7997 10265 8031
rect 10299 7997 10338 8031
rect 10372 7997 10411 8031
rect 10445 7997 10484 8031
rect 10518 7997 10557 8031
rect 10591 7997 10630 8031
rect 10664 7997 10703 8031
rect 10737 7997 10776 8031
rect 10810 7997 10849 8031
rect 10883 7997 10922 8031
rect 10956 7997 10995 8031
rect 11029 7997 11068 8031
rect 11102 7997 11141 8031
rect 11175 7997 11214 8031
rect 11248 7997 11286 8031
rect 11320 7997 11358 8031
rect 11392 7997 11430 8031
rect 11464 7997 11502 8031
rect 11536 7997 11574 8031
rect 11608 7997 11646 8031
rect 11680 7997 11718 8031
rect 11752 7997 11790 8031
rect 11824 7997 11862 8031
rect 11896 7997 11934 8031
rect 11968 7997 12006 8031
rect 12040 7997 12078 8031
rect 12112 7997 12150 8031
rect 12184 7997 12222 8031
rect 12256 7997 12294 8031
rect 12328 7997 12340 8031
rect 8209 7991 8616 7997
tri 8607 7988 8610 7991 ne
rect 8610 7988 8616 7991
rect 8668 7988 8680 7997
rect 8732 7991 12340 7997
rect 8732 7988 8738 7991
tri 8738 7988 8741 7991 nw
tri 8607 7896 8610 7899 se
tri 8607 7847 8610 7850 ne
rect 8610 7847 8616 7899
rect 8668 7847 8680 7899
rect 8732 7847 8738 7899
tri 8738 7896 8741 7899 sw
rect 10209 7850 10525 7896
tri 8738 7847 8741 7850 nw
rect 8096 7806 8148 7818
tri 10238 7812 10241 7815 se
rect 10241 7812 10463 7818
tri 8148 7806 8154 7812 sw
tri 10232 7806 10238 7812 se
rect 10238 7810 10463 7812
rect 10238 7806 10319 7810
rect 8096 7772 8105 7806
rect 8139 7778 8154 7806
tri 8154 7778 8182 7806 sw
tri 10204 7778 10232 7806 se
rect 10232 7778 10247 7806
rect 8139 7772 10247 7778
rect 10281 7772 10319 7806
rect 8096 7758 10319 7772
rect 10371 7806 10463 7810
tri 10463 7806 10469 7812 sw
tri 12547 7806 12553 7812 se
rect 12553 7806 12605 7818
rect 10371 7772 10423 7806
rect 10457 7778 10469 7806
tri 10469 7778 10497 7806 sw
tri 12519 7778 12547 7806 se
rect 12547 7778 12565 7806
rect 10457 7772 12565 7778
rect 12599 7772 12605 7806
rect 10371 7758 12605 7772
rect 8096 7746 12605 7758
rect 8096 7734 10319 7746
rect 8096 7700 8105 7734
rect 8139 7732 10247 7734
rect 8139 7700 8150 7732
tri 8150 7700 8182 7732 nw
tri 10204 7700 10236 7732 ne
rect 10236 7700 10247 7732
rect 10281 7700 10319 7734
rect 8096 7688 8148 7700
tri 8148 7698 8150 7700 nw
tri 10236 7698 10238 7700 ne
rect 10238 7698 10319 7700
tri 10238 7695 10241 7698 ne
rect 10241 7694 10319 7698
rect 10371 7734 12605 7746
rect 10371 7700 10423 7734
rect 10457 7732 12565 7734
rect 10457 7700 10465 7732
tri 10465 7700 10497 7732 nw
tri 12519 7700 12551 7732 ne
rect 12551 7700 12565 7732
rect 12599 7700 12605 7734
rect 10371 7694 10463 7700
tri 10463 7698 10465 7700 nw
tri 12551 7698 12553 7700 ne
rect 10241 7688 10463 7694
rect 12553 7688 12605 7700
tri 8607 7660 8610 7663 se
tri 8607 7611 8610 7614 ne
rect 8610 7611 8616 7663
rect 8668 7611 8680 7663
rect 8732 7611 8738 7663
tri 8738 7660 8741 7663 sw
rect 10209 7614 10562 7660
tri 8738 7611 8741 7614 nw
rect 3889 7574 7760 7580
rect 3889 7540 3901 7574
rect 3935 7540 3974 7574
rect 4008 7540 4047 7574
rect 4081 7540 4120 7574
rect 4154 7540 4193 7574
rect 4227 7540 4266 7574
rect 4300 7540 4339 7574
rect 4373 7540 4412 7574
rect 4446 7540 4485 7574
rect 4519 7540 4558 7574
rect 4592 7540 4631 7574
rect 4665 7540 4704 7574
rect 4738 7540 4777 7574
rect 4811 7540 4850 7574
rect 4884 7540 4923 7574
rect 4957 7540 4996 7574
rect 5030 7540 5069 7574
rect 5103 7540 5142 7574
rect 5176 7540 5215 7574
rect 5249 7540 5288 7574
rect 5322 7540 5361 7574
rect 5395 7540 5434 7574
rect 5468 7540 5507 7574
rect 5541 7540 5580 7574
rect 5614 7540 5653 7574
rect 5687 7540 5726 7574
rect 5760 7540 5799 7574
rect 5833 7540 5872 7574
rect 5906 7540 5945 7574
rect 5979 7540 6018 7574
rect 6052 7540 6091 7574
rect 6125 7540 6164 7574
rect 6198 7540 6237 7574
rect 6271 7540 6310 7574
rect 6344 7540 6383 7574
rect 6417 7540 6456 7574
rect 6490 7540 6530 7574
rect 6564 7540 6604 7574
rect 6638 7540 6678 7574
rect 6712 7540 6752 7574
rect 6786 7540 6826 7574
rect 6860 7540 6900 7574
rect 6934 7540 6974 7574
rect 7008 7540 7048 7574
rect 7082 7540 7122 7574
rect 7156 7540 7196 7574
rect 7230 7540 7270 7574
rect 7304 7540 7344 7574
rect 7378 7540 7418 7574
rect 7452 7540 7492 7574
rect 7526 7540 7566 7574
rect 7600 7540 7640 7574
rect 7674 7540 7714 7574
rect 7748 7540 7760 7574
rect 3889 7534 7760 7540
rect 8096 7570 8148 7582
tri 10238 7576 10241 7579 se
rect 10241 7576 10463 7582
tri 8148 7570 8154 7576 sw
tri 10232 7570 10238 7576 se
rect 10238 7575 10463 7576
rect 10238 7570 10319 7575
rect 8096 7536 8105 7570
rect 8139 7542 8154 7570
tri 8154 7542 8182 7570 sw
tri 10204 7542 10232 7570 se
rect 10232 7542 10247 7570
rect 8139 7536 10247 7542
rect 10281 7536 10319 7570
rect 8096 7523 10319 7536
rect 10371 7570 10463 7575
tri 10463 7570 10469 7576 sw
tri 12547 7570 12553 7576 se
rect 12553 7570 12605 7582
rect 10371 7536 10423 7570
rect 10457 7542 10469 7570
tri 10469 7542 10497 7570 sw
tri 12519 7542 12547 7570 se
rect 12547 7542 12565 7570
rect 10457 7536 12565 7542
rect 12599 7536 12605 7570
rect 10371 7523 12605 7536
rect 8096 7511 12605 7523
rect 8096 7498 10319 7511
rect 3889 7483 3935 7495
rect 3889 7449 3895 7483
rect 3929 7449 3935 7483
rect 8096 7464 8105 7498
rect 8139 7496 10247 7498
rect 8139 7464 8150 7496
tri 8150 7464 8182 7496 nw
tri 10204 7464 10236 7496 ne
rect 10236 7464 10247 7496
rect 10281 7464 10319 7498
rect 8096 7452 8148 7464
tri 8148 7462 8150 7464 nw
tri 10236 7462 10238 7464 ne
rect 10238 7462 10319 7464
tri 10238 7459 10241 7462 ne
rect 10241 7459 10319 7462
rect 10371 7498 12605 7511
rect 10371 7464 10423 7498
rect 10457 7496 12565 7498
rect 10457 7464 10465 7496
tri 10465 7464 10497 7496 nw
tri 12519 7464 12551 7496 ne
rect 12551 7464 12565 7496
rect 12599 7464 12605 7498
rect 10371 7459 10463 7464
tri 10463 7462 10465 7464 nw
tri 12551 7462 12553 7464 ne
rect 10241 7452 10463 7459
rect 12553 7452 12605 7464
rect 3889 7401 3935 7449
tri 8607 7424 8610 7427 se
rect 3889 7367 3895 7401
rect 3929 7367 3935 7401
rect 3889 7319 3935 7367
rect 3889 7285 3895 7319
rect 3929 7285 3935 7319
rect 3889 7237 3935 7285
rect 3889 7203 3895 7237
rect 3929 7203 3935 7237
rect 3889 7155 3935 7203
rect 3889 7121 3895 7155
rect 3929 7121 3935 7155
rect 3889 7074 3935 7121
rect 3889 7040 3895 7074
rect 3929 7040 3935 7074
rect 3889 6993 3935 7040
rect 3889 6959 3895 6993
rect 3929 6959 3935 6993
rect 3889 6947 3935 6959
rect 4102 7386 4407 7392
rect 4102 7352 4180 7386
rect 4214 7352 4271 7386
rect 4305 7352 4361 7386
rect 4395 7352 4407 7386
rect 4102 7346 4407 7352
rect 4993 7386 5508 7392
rect 4993 7352 5005 7386
rect 5039 7352 5083 7386
rect 5117 7352 5161 7386
rect 5195 7352 5239 7386
rect 5273 7352 5317 7386
rect 5351 7352 5396 7386
rect 5430 7352 5508 7386
rect 4993 7346 5508 7352
rect 5878 7386 6370 7392
rect 5878 7352 5890 7386
rect 5924 7352 5963 7386
rect 5997 7352 6036 7386
rect 6070 7352 6110 7386
rect 6144 7352 6184 7386
rect 6218 7352 6258 7386
rect 6292 7352 6370 7386
rect 5878 7346 6370 7352
rect 6996 7386 7300 7392
rect 6996 7352 7008 7386
rect 7042 7352 7090 7386
rect 7124 7352 7172 7386
rect 7206 7352 7254 7386
rect 7288 7352 7300 7386
rect 6996 7346 7300 7352
rect 7428 7346 7500 7392
tri 8607 7375 8610 7378 ne
rect 8610 7375 8616 7427
rect 8668 7375 8680 7427
rect 8732 7375 8738 7427
tri 8738 7424 8741 7427 sw
rect 10209 7378 10644 7424
tri 8738 7375 8741 7378 nw
rect 4102 7338 4174 7346
tri 4174 7338 4182 7346 nw
tri 5428 7338 5436 7346 ne
rect 5436 7338 5508 7346
tri 6290 7338 6298 7346 ne
rect 6298 7338 6370 7346
tri 7428 7338 7436 7346 ne
rect 7436 7338 7500 7346
rect 4102 7302 4148 7338
tri 4148 7312 4174 7338 nw
tri 5436 7312 5462 7338 ne
rect 4102 7268 4108 7302
rect 4142 7268 4148 7302
rect 5462 7301 5508 7338
tri 6298 7312 6324 7338 ne
rect 6324 7312 6370 7338
tri 7436 7320 7454 7338 ne
rect 4102 7218 4148 7268
rect 4444 7226 4523 7272
tri 4968 7267 4973 7272 se
rect 4973 7267 5126 7272
tri 4967 7266 4968 7267 se
rect 4968 7266 5126 7267
tri 4939 7238 4967 7266 se
rect 4967 7238 5126 7266
tri 4927 7226 4939 7238 se
rect 4939 7226 5126 7238
rect 5327 7226 5405 7272
rect 4102 7184 4108 7218
rect 4142 7184 4148 7218
tri 4437 7215 4448 7226 ne
rect 4448 7215 4523 7226
tri 4916 7215 4927 7226 se
rect 4927 7215 4982 7226
tri 4982 7215 4993 7226 nw
tri 5325 7215 5336 7226 ne
rect 5336 7215 5405 7226
tri 4448 7194 4469 7215 ne
rect 4469 7194 4523 7215
tri 4895 7194 4916 7215 se
rect 4916 7194 4961 7215
tri 4961 7194 4982 7215 nw
tri 5336 7194 5357 7215 ne
rect 5357 7194 5405 7215
tri 4469 7192 4471 7194 ne
rect 4102 7133 4148 7184
rect 4102 7099 4108 7133
rect 4142 7099 4148 7133
rect 4102 7064 4148 7099
rect 4471 7186 4523 7194
tri 4889 7188 4895 7194 se
rect 4895 7192 4959 7194
tri 4959 7192 4961 7194 nw
tri 5357 7192 5359 7194 ne
rect 4895 7188 4955 7192
tri 4955 7188 4959 7192 nw
tri 4883 7182 4889 7188 se
rect 4889 7182 4949 7188
tri 4949 7182 4955 7188 nw
rect 5359 7182 5405 7194
tri 4849 7148 4883 7182 se
rect 4883 7148 4915 7182
tri 4915 7148 4949 7182 nw
rect 5359 7148 5365 7182
rect 5399 7148 5405 7182
rect 4471 7122 4523 7134
tri 4830 7129 4849 7148 se
rect 4849 7129 4896 7148
tri 4896 7129 4915 7148 nw
tri 4823 7122 4830 7129 se
rect 4830 7122 4889 7129
tri 4889 7122 4896 7129 nw
tri 4811 7110 4823 7122 se
rect 4823 7110 4877 7122
tri 4877 7110 4889 7122 nw
rect 5359 7110 5405 7148
tri 4777 7076 4811 7110 se
rect 4811 7076 4843 7110
tri 4843 7076 4877 7110 nw
rect 5359 7076 5365 7110
rect 5399 7076 5405 7110
rect 5462 7267 5468 7301
rect 5502 7267 5508 7301
rect 6324 7278 6330 7312
rect 6364 7278 6370 7312
tri 7349 7302 7350 7303 se
rect 7350 7302 7402 7307
tri 5756 7268 5760 7272 se
rect 5760 7268 5984 7272
rect 5462 7215 5508 7267
tri 5754 7266 5756 7268 se
rect 5756 7266 5984 7268
tri 5726 7238 5754 7266 se
rect 5754 7238 5984 7266
tri 5714 7226 5726 7238 se
rect 5726 7226 5984 7238
rect 6184 7226 6263 7272
rect 5462 7181 5468 7215
rect 5502 7181 5508 7215
tri 5692 7204 5714 7226 se
rect 5714 7204 5758 7226
tri 5758 7204 5780 7226 nw
tri 6184 7204 6206 7226 ne
rect 6206 7204 6263 7226
tri 5676 7188 5692 7204 se
rect 5692 7194 5748 7204
tri 5748 7194 5758 7204 nw
tri 6206 7194 6216 7204 ne
rect 6216 7194 6263 7204
rect 5692 7193 5747 7194
tri 5747 7193 5748 7194 nw
tri 6216 7193 6217 7194 ne
rect 5692 7188 5742 7193
tri 5742 7188 5747 7193 nw
tri 5672 7184 5676 7188 se
rect 5676 7184 5738 7188
tri 5738 7184 5742 7188 nw
tri 5670 7182 5672 7184 se
rect 5672 7182 5736 7184
tri 5736 7182 5738 7184 nw
rect 6217 7182 6263 7194
rect 5462 7129 5508 7181
tri 5636 7148 5670 7182 se
rect 5670 7148 5702 7182
tri 5702 7148 5736 7182 nw
rect 6217 7148 6223 7182
rect 6257 7148 6263 7182
tri 5617 7129 5636 7148 se
rect 5636 7129 5683 7148
tri 5683 7129 5702 7148 nw
rect 5462 7095 5468 7129
rect 5502 7095 5508 7129
tri 5610 7122 5617 7129 se
rect 5617 7122 5676 7129
tri 5676 7122 5683 7129 nw
tri 5598 7110 5610 7122 se
rect 5610 7110 5664 7122
tri 5664 7110 5676 7122 nw
rect 6217 7110 6263 7148
rect 6324 7238 6370 7278
tri 7319 7272 7349 7302 se
rect 7349 7301 7402 7302
rect 7349 7272 7350 7301
tri 7029 7268 7033 7272 se
rect 7033 7268 7120 7272
tri 7027 7266 7029 7268 se
rect 7029 7266 7120 7268
rect 6324 7204 6330 7238
rect 6364 7204 6370 7238
tri 6993 7232 7027 7266 se
rect 7027 7232 7120 7266
tri 6989 7228 6993 7232 se
rect 6993 7228 7120 7232
tri 6987 7226 6989 7228 se
rect 6989 7226 7120 7228
rect 7321 7249 7350 7272
rect 7321 7237 7402 7249
rect 7321 7226 7350 7237
tri 6979 7218 6987 7226 se
rect 6987 7218 7045 7226
tri 7045 7218 7053 7226 nw
tri 7319 7218 7327 7226 ne
rect 7327 7218 7350 7226
rect 6324 7163 6370 7204
tri 6949 7188 6979 7218 se
rect 6979 7192 7019 7218
tri 7019 7192 7045 7218 nw
tri 7327 7195 7350 7218 ne
rect 6979 7188 7015 7192
tri 7015 7188 7019 7192 nw
tri 6945 7184 6949 7188 se
rect 6949 7184 7011 7188
tri 7011 7184 7015 7188 nw
tri 6940 7179 6945 7184 se
rect 6945 7179 7006 7184
tri 7006 7179 7011 7184 nw
rect 7350 7179 7402 7185
rect 6324 7129 6330 7163
rect 6364 7129 6370 7163
tri 6906 7145 6940 7179 se
rect 6940 7145 6972 7179
tri 6972 7145 7006 7179 nw
rect 7350 7145 7359 7179
rect 7393 7145 7402 7179
tri 6894 7133 6906 7145 se
rect 6906 7133 6960 7145
tri 6960 7133 6972 7145 nw
rect 6324 7117 6370 7129
tri 6883 7122 6894 7133 se
rect 6894 7122 6949 7133
tri 6949 7122 6960 7133 nw
tri 6878 7117 6883 7122 se
rect 6883 7117 6944 7122
tri 6944 7117 6949 7122 nw
rect 5462 7083 5508 7095
tri 5571 7083 5598 7110 se
rect 5598 7083 5637 7110
tri 5637 7083 5664 7110 nw
tri 5564 7076 5571 7083 se
rect 5571 7076 5630 7083
tri 5630 7076 5637 7083 nw
rect 6217 7076 6223 7110
rect 6257 7076 6263 7110
tri 6868 7107 6878 7117 se
rect 6878 7107 6934 7117
tri 6934 7107 6944 7117 nw
rect 7350 7107 7402 7145
tri 4774 7073 4777 7076 se
rect 4777 7073 4840 7076
tri 4840 7073 4843 7076 nw
tri 4148 7064 4154 7070 sw
rect 4471 7064 4523 7070
tri 4765 7064 4774 7073 se
rect 4774 7064 4831 7073
tri 4831 7064 4840 7073 nw
rect 5359 7064 5405 7076
tri 5561 7073 5564 7076 se
rect 5564 7073 5627 7076
tri 5627 7073 5630 7076 nw
tri 5552 7064 5561 7073 se
rect 5561 7064 5618 7073
tri 5618 7064 5627 7073 nw
rect 6217 7064 6263 7076
tri 6834 7073 6868 7107 se
rect 6868 7073 6900 7107
tri 6900 7073 6934 7107 nw
rect 7350 7073 7359 7107
rect 7393 7073 7402 7107
tri 6825 7064 6834 7073 se
rect 6834 7064 6891 7073
tri 6891 7064 6900 7073 nw
rect 4102 7061 4154 7064
tri 4154 7061 4157 7064 sw
tri 4762 7061 4765 7064 se
rect 4765 7061 4828 7064
tri 4828 7061 4831 7064 nw
tri 5549 7061 5552 7064 se
rect 5552 7061 5615 7064
tri 5615 7061 5618 7064 nw
tri 6822 7061 6825 7064 se
rect 6825 7061 6888 7064
tri 6888 7061 6891 7064 nw
rect 7350 7061 7402 7073
rect 7454 7302 7500 7338
rect 7454 7268 7460 7302
rect 7494 7268 7500 7302
rect 7454 7218 7500 7268
rect 8096 7338 8148 7350
rect 10241 7339 10463 7346
rect 8096 7304 8105 7338
rect 8139 7334 8148 7338
tri 10238 7336 10241 7339 se
rect 10241 7336 10319 7339
tri 8148 7334 8150 7336 sw
tri 10236 7334 10238 7336 se
rect 10238 7334 10319 7336
rect 8139 7304 8150 7334
rect 8096 7302 8150 7304
tri 8150 7302 8182 7334 sw
tri 10204 7302 10236 7334 se
rect 10236 7302 10247 7334
rect 8096 7300 10247 7302
rect 10281 7300 10319 7334
rect 8096 7287 10319 7300
rect 10371 7334 10463 7339
tri 10463 7334 10465 7336 sw
tri 12551 7334 12553 7336 se
rect 12553 7334 12605 7350
rect 10371 7300 10423 7334
rect 10457 7302 10465 7334
tri 10465 7302 10497 7334 sw
tri 12519 7302 12551 7334 se
rect 12551 7302 12565 7334
rect 10457 7300 12565 7302
rect 12599 7300 12605 7334
rect 10371 7287 12605 7300
rect 8096 7275 12605 7287
rect 8096 7266 10319 7275
rect 8096 7232 8105 7266
rect 8139 7262 10319 7266
rect 8139 7256 10247 7262
rect 8139 7232 8154 7256
rect 8096 7228 8154 7232
tri 8154 7228 8182 7256 nw
tri 10204 7228 10232 7256 ne
rect 10232 7228 10247 7256
rect 10281 7228 10319 7262
rect 8096 7220 8148 7228
tri 8148 7222 8154 7228 nw
tri 10232 7222 10238 7228 ne
rect 10238 7223 10319 7228
rect 10371 7262 12605 7275
rect 10371 7228 10423 7262
rect 10457 7256 12565 7262
rect 10457 7228 10469 7256
tri 10469 7228 10497 7256 nw
tri 12519 7228 12547 7256 ne
rect 12547 7228 12565 7256
rect 12599 7228 12605 7262
rect 10371 7223 10463 7228
rect 10238 7222 10463 7223
tri 10463 7222 10469 7228 nw
tri 12547 7222 12553 7228 ne
tri 10238 7220 10240 7222 ne
rect 10240 7220 10463 7222
tri 10240 7219 10241 7220 ne
rect 7454 7184 7460 7218
rect 7494 7184 7500 7218
rect 10241 7216 10463 7220
rect 12553 7216 12605 7228
tri 8607 7188 8610 7191 se
rect 7454 7133 7500 7184
tri 8607 7139 8610 7142 ne
rect 8610 7139 8616 7191
rect 8668 7139 8680 7191
rect 8732 7139 8738 7191
tri 8738 7188 8741 7191 sw
rect 10209 7142 10525 7188
tri 8738 7139 8741 7142 nw
rect 7454 7099 7460 7133
rect 7494 7099 7500 7133
rect 4102 7048 4157 7061
tri 4157 7048 4170 7061 sw
tri 4757 7056 4762 7061 se
rect 4762 7056 4823 7061
tri 4823 7056 4828 7061 nw
tri 5544 7056 5549 7061 se
rect 5549 7056 5610 7061
tri 5610 7056 5615 7061 nw
tri 6817 7056 6822 7061 se
rect 6822 7056 6883 7061
tri 6883 7056 6888 7061 nw
tri 4749 7048 4757 7056 se
rect 4757 7048 4815 7056
tri 4815 7048 4823 7056 nw
tri 5536 7048 5544 7056 se
rect 5544 7048 5602 7056
tri 5602 7048 5610 7056 nw
tri 6809 7048 6817 7056 se
rect 6817 7048 6875 7056
tri 6875 7048 6883 7056 nw
rect 7454 7048 7500 7099
rect 4102 7014 4108 7048
rect 4142 7036 4170 7048
tri 4170 7036 4182 7048 sw
tri 4737 7036 4749 7048 se
rect 4749 7036 4803 7048
tri 4803 7036 4815 7048 nw
tri 5524 7036 5536 7048 se
rect 5536 7036 5590 7048
tri 5590 7036 5602 7048 nw
tri 6797 7036 6809 7048 se
rect 6809 7036 6863 7048
tri 6863 7036 6875 7048 nw
rect 4142 7014 4781 7036
tri 4781 7014 4803 7036 nw
rect 4988 7014 5568 7036
tri 5568 7014 5590 7036 nw
rect 5983 7014 6841 7036
tri 6841 7014 6863 7036 nw
rect 4102 6994 4761 7014
tri 4761 6994 4781 7014 nw
rect 4988 6994 5548 7014
tri 5548 6994 5568 7014 nw
rect 5983 6994 6821 7014
tri 6821 6994 6841 7014 nw
rect 6973 6994 7236 7036
rect 4102 6990 4757 6994
tri 4757 6990 4761 6994 nw
rect 4988 6990 5544 6994
tri 5544 6990 5548 6994 nw
rect 5983 6990 6817 6994
tri 6817 6990 6821 6994 nw
rect 4102 6963 4596 6990
rect 4102 6929 4108 6963
rect 4142 6960 4596 6963
tri 4596 6960 4626 6990 nw
rect 4988 6960 5514 6990
tri 5514 6960 5544 6990 nw
rect 5983 6960 6390 6990
tri 6390 6960 6420 6990 nw
rect 6973 6960 6980 6994
rect 7014 6990 7236 6994
tri 7321 7014 7331 7024 sw
tri 7444 7014 7454 7024 se
rect 7454 7014 7460 7048
rect 7494 7014 7500 7048
rect 7321 6992 7331 7014
tri 7331 6992 7353 7014 sw
tri 7422 6992 7444 7014 se
rect 7444 6992 7500 7014
rect 7321 6990 7353 6992
tri 7353 6990 7355 6992 sw
tri 7420 6990 7422 6992 se
rect 7422 6990 7500 6992
rect 7014 6963 7500 6990
rect 8096 7098 8148 7110
rect 10241 7103 10463 7110
tri 10238 7099 10241 7102 se
rect 10241 7099 10319 7103
tri 8148 7098 8149 7099 sw
tri 10237 7098 10238 7099 se
rect 10238 7098 10319 7099
rect 8096 7064 8105 7098
rect 8139 7065 8149 7098
tri 8149 7065 8182 7098 sw
tri 10204 7065 10237 7098 se
rect 10237 7065 10247 7098
rect 8139 7064 10247 7065
rect 10281 7064 10319 7098
rect 8096 7051 10319 7064
rect 10371 7098 10463 7103
tri 10463 7098 10464 7099 sw
tri 12552 7098 12553 7099 se
rect 12553 7098 12605 7110
rect 10371 7064 10423 7098
rect 10457 7065 10464 7098
tri 10464 7065 10497 7098 sw
tri 12519 7065 12552 7098 se
rect 12552 7065 12565 7098
rect 10457 7064 12565 7065
rect 12599 7064 12605 7098
rect 10371 7051 12605 7064
rect 8096 7039 12605 7051
rect 8096 7026 10319 7039
rect 8096 6992 8105 7026
rect 8139 7019 10247 7026
rect 8139 6992 8155 7019
tri 8155 6992 8182 7019 nw
tri 10204 6992 10231 7019 ne
rect 10231 6992 10247 7019
rect 10281 6992 10319 7026
rect 8096 6980 8148 6992
tri 8148 6985 8155 6992 nw
tri 10231 6985 10238 6992 ne
rect 10238 6987 10319 6992
rect 10371 7026 12605 7039
rect 10371 6992 10423 7026
rect 10457 7019 12565 7026
rect 10457 6992 10470 7019
tri 10470 6992 10497 7019 nw
tri 12519 6992 12546 7019 ne
rect 12546 6992 12565 7019
rect 12599 6992 12605 7026
rect 10371 6987 10463 6992
rect 10238 6985 10463 6987
tri 10463 6985 10470 6992 nw
tri 12546 6985 12553 6992 ne
tri 10238 6982 10241 6985 ne
rect 10241 6980 10463 6985
rect 12553 6980 12605 6992
rect 7014 6960 7460 6963
rect 4142 6929 4592 6960
tri 4592 6956 4596 6960 nw
rect 4102 6891 4592 6929
rect 4102 6857 4181 6891
rect 4215 6857 4254 6891
rect 4288 6857 4327 6891
rect 4361 6857 4400 6891
rect 4434 6857 4473 6891
rect 4507 6857 4546 6891
rect 4580 6857 4592 6891
rect 4102 6851 4592 6857
rect 4988 6912 5508 6960
tri 5508 6954 5514 6960 nw
tri 5981 6929 5983 6931 se
rect 5983 6929 6386 6960
tri 6386 6956 6390 6960 nw
rect 4988 6891 5468 6912
rect 4988 6857 5000 6891
rect 5034 6857 5078 6891
rect 5112 6857 5156 6891
rect 5190 6857 5234 6891
rect 5268 6857 5312 6891
rect 5346 6857 5390 6891
rect 5424 6878 5468 6891
rect 5502 6878 5508 6912
tri 5949 6897 5981 6929 se
rect 5981 6897 6386 6929
rect 5424 6857 5508 6878
rect 4988 6851 5508 6857
rect 5839 6891 6386 6897
rect 5839 6857 5913 6891
rect 5947 6857 5995 6891
rect 6029 6857 6072 6891
rect 6106 6857 6149 6891
rect 6183 6857 6221 6891
rect 6255 6857 6340 6891
rect 6374 6857 6386 6891
rect 5839 6851 6386 6857
rect 6973 6929 7460 6960
rect 7494 6929 7500 6963
tri 8607 6952 8610 6955 se
rect 6973 6891 7500 6929
tri 8607 6903 8610 6906 ne
rect 8610 6903 8616 6955
rect 8668 6903 8680 6955
rect 8732 6903 8738 6955
tri 8738 6952 8741 6955 sw
rect 10209 6906 10550 6952
tri 8738 6903 8741 6906 nw
rect 6973 6857 7052 6891
rect 7086 6857 7134 6891
rect 7168 6857 7216 6891
rect 7250 6857 7298 6891
rect 7332 6857 7379 6891
rect 7413 6857 7500 6891
rect 6973 6851 7500 6857
rect 11102 6552 11108 6604
rect 11160 6552 11175 6604
rect 11227 6552 11656 6604
rect 11708 6552 11723 6604
rect 11775 6552 11781 6604
rect 10704 6519 10756 6525
tri 10756 6501 10780 6525 sw
rect 10756 6467 11483 6501
rect 10704 6452 11483 6467
rect 10756 6449 11483 6452
rect 11535 6449 11550 6501
rect 11602 6449 11608 6501
tri 10756 6415 10790 6449 nw
rect 10704 6394 10756 6400
rect 11208 5277 11214 5329
rect 11266 5277 11278 5329
rect 11330 5277 11342 5329
rect 11394 5277 11406 5329
rect 11458 5277 11470 5329
rect 11522 5277 11807 5329
rect 11245 5179 11807 5240
rect 11245 5127 11556 5179
rect 11608 5127 11807 5179
rect 11245 5090 11807 5127
rect 11245 5038 11556 5090
rect 11608 5038 11807 5090
rect 11245 5001 11807 5038
rect 11245 4949 11556 5001
rect 11608 4949 11807 5001
rect 11835 5109 12071 5115
rect 11835 5103 12019 5109
rect 11835 5069 11841 5103
rect 11875 5069 12019 5103
rect 11835 5057 12019 5069
rect 11835 5042 12071 5057
rect 11835 5030 12019 5042
rect 11835 4996 11841 5030
rect 11875 4996 12019 5030
rect 11835 4990 12019 4996
rect 11835 4984 12071 4990
rect 11245 4912 11807 4949
rect 11245 4860 11556 4912
rect 11608 4860 11807 4912
rect 11245 4854 11807 4860
rect 11208 4766 11214 4818
rect 11266 4766 11278 4818
rect 11330 4766 11342 4818
rect 11394 4766 11406 4818
rect 11458 4766 11470 4818
rect 11522 4766 11807 4818
rect 11208 3230 11214 3282
rect 11266 3230 11278 3282
rect 11330 3230 11342 3282
rect 11394 3230 11406 3282
rect 11458 3230 11470 3282
rect 11522 3230 11807 3282
rect 11245 3186 11882 3192
rect 11245 3134 11556 3186
rect 11608 3180 11882 3186
rect 11608 3146 11839 3180
rect 11873 3146 11882 3180
rect 11608 3134 11882 3146
rect 11245 3108 11882 3134
rect 11245 3107 11839 3108
rect 11245 3055 11556 3107
rect 11608 3074 11839 3107
rect 11873 3074 11882 3108
rect 11608 3055 11882 3074
rect 11245 3027 11882 3055
rect 11245 2975 11556 3027
rect 11608 2975 11882 3027
rect 11245 2947 11882 2975
rect 11245 2895 11556 2947
rect 11608 2924 11882 2947
rect 11608 2895 11839 2924
rect 11245 2890 11839 2895
rect 11873 2890 11882 2924
rect 11245 2867 11882 2890
rect 11245 2815 11556 2867
rect 11608 2852 11882 2867
rect 11608 2818 11839 2852
rect 11873 2818 11882 2852
rect 11608 2815 11882 2818
rect 11245 2806 11882 2815
rect 11208 2718 11214 2770
rect 11266 2718 11278 2770
rect 11330 2718 11342 2770
rect 11394 2718 11406 2770
rect 11458 2718 11470 2770
rect 11522 2718 11807 2770
<< via1 >>
rect 7829 14775 7881 14827
rect 7673 14698 7725 14750
rect 7737 14698 7789 14750
rect 7829 14711 7881 14763
rect 13903 14805 13955 14857
rect 13967 14805 14019 14857
rect 13440 14766 13492 14775
rect 13504 14766 13556 14775
rect 13440 14732 13472 14766
rect 13472 14732 13492 14766
rect 13504 14732 13506 14766
rect 13506 14732 13546 14766
rect 13546 14732 13556 14766
rect 13440 14723 13492 14732
rect 13504 14723 13556 14732
rect 6626 14607 6678 14659
rect 6690 14607 6742 14659
rect 3059 14552 3111 14558
rect 3059 14518 3071 14552
rect 3071 14518 3105 14552
rect 3105 14518 3111 14552
rect 3059 14506 3111 14518
rect 3059 14476 3111 14492
rect 3059 14442 3071 14476
rect 3071 14442 3105 14476
rect 3105 14442 3111 14476
rect 3059 14440 3111 14442
rect 3059 14400 3111 14426
rect 3059 14374 3071 14400
rect 3071 14374 3105 14400
rect 3105 14374 3111 14400
rect 3059 14324 3111 14360
rect 3059 14308 3071 14324
rect 3071 14308 3105 14324
rect 3105 14308 3111 14324
rect 3059 14290 3071 14294
rect 3071 14290 3105 14294
rect 3105 14290 3111 14294
rect 3059 14248 3111 14290
rect 3059 14242 3071 14248
rect 3071 14242 3105 14248
rect 3105 14242 3111 14248
rect 3059 14214 3071 14228
rect 3071 14214 3105 14228
rect 3105 14214 3111 14228
rect 3059 14176 3111 14214
rect 3059 14138 3071 14162
rect 3071 14138 3105 14162
rect 3105 14138 3111 14162
rect 3059 14110 3111 14138
rect 3059 14062 3071 14096
rect 3071 14062 3105 14096
rect 3105 14062 3111 14096
rect 3059 14044 3111 14062
rect 3059 14020 3111 14030
rect 3059 13986 3071 14020
rect 3071 13986 3105 14020
rect 3105 13986 3111 14020
rect 3059 13978 3111 13986
rect 3059 13944 3111 13964
rect 3059 13912 3071 13944
rect 3071 13912 3105 13944
rect 3105 13912 3111 13944
rect 3059 13868 3111 13898
rect 3059 13846 3071 13868
rect 3071 13846 3105 13868
rect 3105 13846 3111 13868
rect 3059 13792 3111 13832
rect 3059 13780 3071 13792
rect 3071 13780 3105 13792
rect 3105 13780 3111 13792
rect 3059 13758 3071 13765
rect 3071 13758 3105 13765
rect 3105 13758 3111 13765
rect 3059 13716 3111 13758
rect 3059 13713 3071 13716
rect 3071 13713 3105 13716
rect 3105 13713 3111 13716
rect 3059 13682 3071 13698
rect 3071 13682 3105 13698
rect 3105 13682 3111 13698
rect 3059 13646 3111 13682
rect 3059 13605 3071 13631
rect 3071 13605 3105 13631
rect 3105 13605 3111 13631
rect 3059 13579 3111 13605
rect 3059 13562 3111 13564
rect 3059 13528 3071 13562
rect 3071 13528 3105 13562
rect 3105 13528 3111 13562
rect 3059 13512 3111 13528
rect 3059 13485 3111 13497
rect 3059 13451 3071 13485
rect 3071 13451 3105 13485
rect 3105 13451 3111 13485
rect 3059 13445 3111 13451
rect -175 12940 -123 12992
rect -175 12876 -123 12928
rect -175 12812 -123 12864
rect -175 12748 -123 12800
rect -175 12683 -123 12735
rect -175 12618 -123 12670
rect -175 12553 -123 12605
rect -175 12488 -123 12540
rect -175 12423 -123 12475
rect -175 12358 -123 12410
rect -175 12293 -123 12345
rect -175 12228 -123 12280
rect -175 12163 -123 12215
rect 13941 14540 13993 14592
rect 14005 14540 14057 14592
rect 5132 14339 5184 14391
rect 5232 14339 5284 14391
rect 5132 14274 5184 14326
rect 5232 14274 5284 14326
rect 5132 14209 5184 14261
rect 5232 14209 5284 14261
rect 5132 14144 5184 14196
rect 5232 14144 5284 14196
rect 5132 14079 5184 14131
rect 5232 14079 5284 14131
rect 5132 14014 5184 14066
rect 5232 14014 5284 14066
rect 10319 14072 10371 14124
rect 10319 14008 10371 14060
rect 5132 13949 5184 14001
rect 5232 13949 5284 14001
rect 5132 13884 5184 13936
rect 5232 13884 5284 13936
rect 7743 13917 7795 13969
rect 5132 13818 5184 13870
rect 5232 13818 5284 13870
rect 6622 13841 6674 13893
rect 6686 13841 6738 13893
rect 7743 13853 7795 13905
rect 4936 13746 4988 13798
rect 5132 13752 5184 13804
rect 5232 13752 5284 13804
rect 4936 13682 4988 13734
rect 5132 13686 5184 13738
rect 5232 13686 5284 13738
rect 4936 13618 4988 13670
rect 5132 13620 5184 13672
rect 5232 13620 5284 13672
rect 4936 13554 4988 13606
rect 5132 13554 5184 13606
rect 5232 13554 5284 13606
rect 4936 13490 4988 13542
rect 5132 13488 5184 13540
rect 5232 13488 5284 13540
rect 4936 13426 4988 13478
rect 4936 13362 4988 13414
rect 5132 13422 5184 13474
rect 5232 13422 5284 13474
rect 4936 13298 4988 13350
rect 5132 13356 5184 13408
rect 5232 13356 5284 13408
rect 4936 13233 4988 13285
rect 5132 13290 5184 13342
rect 5232 13290 5284 13342
rect 4936 13168 4988 13220
rect 5132 13224 5184 13276
rect 5232 13224 5284 13276
rect 5132 13158 5184 13210
rect 5232 13158 5284 13210
rect 4936 13103 4988 13155
rect 5132 13092 5184 13144
rect 5232 13092 5284 13144
rect 4936 13038 4988 13090
rect 5132 13026 5184 13078
rect 5232 13026 5284 13078
rect 4728 12962 4780 12969
rect 4792 12962 4844 12969
rect 4728 12928 4757 12962
rect 4757 12928 4780 12962
rect 4792 12928 4829 12962
rect 4829 12928 4844 12962
rect 4728 12917 4780 12928
rect 4792 12917 4844 12928
rect 5132 12960 5184 13012
rect 5232 12960 5284 13012
rect 5132 12894 5184 12946
rect 5232 12894 5284 12946
rect 4384 12800 4436 12852
rect 4454 12800 4506 12852
rect 4524 12800 4576 12852
rect 4594 12800 4646 12852
rect 4664 12800 4716 12852
rect 4734 12800 4786 12852
rect 4803 12800 4855 12852
rect 5132 12828 5184 12880
rect 5232 12828 5284 12880
rect 4384 12730 4436 12782
rect 4454 12730 4506 12782
rect 4524 12730 4576 12782
rect 4594 12730 4646 12782
rect 4664 12730 4716 12782
rect 4734 12730 4786 12782
rect 4803 12730 4855 12782
rect 5132 12762 5184 12814
rect 5232 12762 5284 12814
rect 4364 12646 4416 12698
rect 4364 12574 4416 12626
rect 4364 12501 4416 12553
rect 4364 12428 4416 12480
rect -201 11981 -149 12033
rect -201 11917 -149 11969
rect 4364 12355 4416 12407
rect 4364 12282 4416 12334
rect 4065 12191 4117 12243
rect 4129 12191 4181 12243
rect 4364 12209 4416 12261
rect 5132 12696 5184 12748
rect 5232 12696 5284 12748
rect 5132 12630 5184 12682
rect 5232 12630 5284 12682
rect 5132 12564 5184 12616
rect 5232 12564 5284 12616
rect 5132 12498 5184 12550
rect 5232 12498 5284 12550
rect 5132 12432 5184 12484
rect 5232 12432 5284 12484
rect 5132 12366 5184 12418
rect 5232 12366 5284 12418
rect 7835 13917 7887 13969
rect 7835 13853 7887 13905
rect 9013 13730 9065 13739
rect 9013 13696 9019 13730
rect 9019 13696 9053 13730
rect 9053 13696 9065 13730
rect 9013 13687 9065 13696
rect 9077 13730 9129 13739
rect 9077 13696 9091 13730
rect 9091 13696 9125 13730
rect 9125 13696 9129 13730
rect 9077 13687 9129 13696
rect 11898 13606 11950 13615
rect 11988 13606 12040 13615
rect 12078 13606 12130 13615
rect 11898 13572 11924 13606
rect 11924 13572 11950 13606
rect 11988 13572 12007 13606
rect 12007 13572 12040 13606
rect 12078 13572 12090 13606
rect 12090 13572 12124 13606
rect 12124 13572 12130 13606
rect 11898 13563 11950 13572
rect 11988 13563 12040 13572
rect 12078 13563 12130 13572
rect 9318 12369 9370 12421
rect 9382 12369 9434 12421
rect 5132 12300 5184 12352
rect 5232 12300 5284 12352
rect 5132 12234 5184 12286
rect 5232 12234 5284 12286
rect 4364 12136 4416 12188
rect 4983 12137 5035 12189
rect 5132 12168 5184 12220
rect 5232 12168 5284 12220
rect 9392 12271 9444 12323
rect 11108 12318 11160 12370
rect 11172 12318 11224 12370
rect 9392 12207 9444 12259
rect 13458 14415 13510 14467
rect 13458 14338 13510 14390
rect 13458 14260 13510 14312
rect 13458 14182 13510 14234
rect 13458 14104 13510 14156
rect 12559 13606 12611 13615
rect 12648 13606 12700 13615
rect 12559 13572 12565 13606
rect 12565 13572 12599 13606
rect 12599 13572 12611 13606
rect 12648 13572 12676 13606
rect 12676 13572 12700 13606
rect 12559 13563 12611 13572
rect 12648 13563 12700 13572
rect 10958 12180 11010 12232
rect 4983 12073 5035 12125
rect 10958 12116 11010 12168
rect 13970 14403 14022 14455
rect 13970 14335 14022 14387
rect 13970 14267 14022 14319
rect 13970 14199 14022 14251
rect 13970 14131 14022 14183
rect 13970 14063 14022 14115
rect 13970 13995 14022 14047
rect 13970 13926 14022 13978
rect 13970 13857 14022 13909
rect 10685 11969 10737 12021
rect 4065 11892 4117 11944
rect 4129 11892 4181 11944
rect 7280 11892 7332 11944
rect 7344 11892 7396 11944
rect 10685 11905 10737 11957
rect 11196 11941 11248 11993
rect 13664 11947 13716 11999
rect 13728 11947 13780 11999
rect 8648 11845 8700 11897
rect 11196 11877 11248 11929
rect 8648 11781 8700 11833
rect 4401 11654 4453 11706
rect 4465 11654 4517 11706
rect 10958 11620 11010 11672
rect 10958 11556 11010 11608
rect 11196 11537 11248 11589
rect 11196 11473 11248 11525
rect -201 9861 -149 9913
rect 10958 10498 11010 10550
rect 10958 10419 11010 10471
rect -201 9797 -149 9849
rect -321 9699 -269 9751
rect -257 9699 -205 9751
rect 12246 8711 12298 8763
rect 12318 8711 12370 8763
rect 12390 8711 12442 8763
rect 12462 8711 12514 8763
rect 12534 8711 12586 8763
rect 10615 8210 10667 8262
rect 10679 8210 10731 8262
rect 8616 8031 8668 8040
rect 8680 8031 8732 8040
rect 8616 7997 8620 8031
rect 8620 7997 8659 8031
rect 8659 7997 8668 8031
rect 8680 7997 8693 8031
rect 8693 7997 8732 8031
rect 8616 7988 8668 7997
rect 8680 7988 8732 7997
rect 8616 7847 8668 7899
rect 8680 7847 8732 7899
rect 10319 7758 10371 7810
rect 10319 7694 10371 7746
rect 8616 7611 8668 7663
rect 8680 7611 8732 7663
rect 10319 7523 10371 7575
rect 10319 7459 10371 7511
rect 8616 7375 8668 7427
rect 8680 7375 8732 7427
rect 4471 7182 4523 7186
rect 4471 7148 4482 7182
rect 4482 7148 4516 7182
rect 4516 7148 4523 7182
rect 4471 7134 4523 7148
rect 4471 7110 4523 7122
rect 4471 7076 4482 7110
rect 4482 7076 4516 7110
rect 4516 7076 4523 7110
rect 7350 7249 7402 7301
rect 7350 7185 7402 7237
rect 4471 7070 4523 7076
rect 10319 7287 10371 7339
rect 10319 7223 10371 7275
rect 8616 7139 8668 7191
rect 8680 7139 8732 7191
rect 10319 7051 10371 7103
rect 10319 6987 10371 7039
rect 8616 6903 8668 6955
rect 8680 6903 8732 6955
rect 11108 6552 11160 6604
rect 11175 6552 11227 6604
rect 11656 6552 11708 6604
rect 11723 6552 11775 6604
rect 10704 6467 10756 6519
rect 10704 6400 10756 6452
rect 11483 6449 11535 6501
rect 11550 6449 11602 6501
rect 11214 5277 11266 5329
rect 11278 5277 11330 5329
rect 11342 5277 11394 5329
rect 11406 5277 11458 5329
rect 11470 5277 11522 5329
rect 11556 5127 11608 5179
rect 11556 5038 11608 5090
rect 11556 4949 11608 5001
rect 12019 5057 12071 5109
rect 12019 4990 12071 5042
rect 11556 4860 11608 4912
rect 11214 4766 11266 4818
rect 11278 4766 11330 4818
rect 11342 4766 11394 4818
rect 11406 4766 11458 4818
rect 11470 4766 11522 4818
rect 11214 3230 11266 3282
rect 11278 3230 11330 3282
rect 11342 3230 11394 3282
rect 11406 3230 11458 3282
rect 11470 3230 11522 3282
rect 11556 3134 11608 3186
rect 11556 3055 11608 3107
rect 11556 2975 11608 3027
rect 11556 2895 11608 2947
rect 11556 2815 11608 2867
rect 11214 2718 11266 2770
rect 11278 2718 11330 2770
rect 11342 2718 11394 2770
rect 11406 2718 11458 2770
rect 11470 2718 11522 2770
<< metal2 >>
rect 7829 14827 7881 14833
rect 13897 14805 13903 14857
rect 13955 14805 13967 14857
rect 14019 14805 14025 14857
tri 13939 14775 13969 14805 ne
rect 13969 14775 14025 14805
rect 7829 14763 7881 14775
rect 7667 14698 7673 14750
rect 7725 14698 7737 14750
rect 7789 14698 7795 14750
rect 7829 14705 7881 14711
tri 7829 14699 7835 14705 ne
tri 7708 14659 7747 14698 ne
rect 7747 14659 7795 14698
rect 6620 14607 6626 14659
rect 6678 14607 6690 14659
rect 6742 14607 6748 14659
tri 7747 14651 7755 14659 ne
tri 6620 14592 6635 14607 ne
rect 6635 14592 6725 14607
tri 6725 14592 6740 14607 nw
tri 6635 14573 6654 14592 ne
rect 3059 14558 3111 14564
rect 3059 14492 3111 14506
rect 3059 14426 3111 14440
rect 3059 14360 3111 14374
rect 3059 14294 3111 14308
rect 3059 14228 3111 14242
rect 3059 14162 3111 14176
rect 3059 14096 3111 14110
rect 3059 14030 3111 14044
rect 3059 13964 3111 13978
rect 3059 13898 3111 13912
rect 3059 13832 3111 13846
rect 5132 14391 5284 14397
rect 5184 14339 5232 14391
rect 5132 14326 5284 14339
rect 5184 14274 5232 14326
rect 5132 14261 5284 14274
rect 5184 14209 5232 14261
rect 5132 14196 5284 14209
rect 5184 14144 5232 14196
rect 5132 14131 5284 14144
rect 5184 14079 5232 14131
rect 5132 14066 5284 14079
rect 5184 14014 5232 14066
rect 5132 14001 5284 14014
rect 5184 13949 5232 14001
rect 5132 13936 5284 13949
rect 5184 13884 5232 13936
tri 6644 13917 6654 13927 se
rect 6654 13917 6706 14592
tri 6706 14573 6725 14592 nw
tri 7746 13978 7755 13987 se
rect 7755 13978 7795 14659
tri 7743 13975 7746 13978 se
rect 7746 13975 7795 13978
rect 7743 13969 7795 13975
tri 6706 13917 6716 13927 sw
tri 6636 13909 6644 13917 se
rect 6644 13909 6716 13917
tri 6716 13909 6724 13917 sw
tri 6632 13905 6636 13909 se
rect 6636 13905 6724 13909
tri 6724 13905 6728 13909 sw
rect 7743 13905 7795 13917
tri 6620 13893 6632 13905 se
rect 6632 13893 6728 13905
tri 6728 13893 6740 13905 sw
rect 5132 13870 5284 13884
rect 5184 13818 5232 13870
rect 6616 13841 6622 13893
rect 6674 13841 6686 13893
rect 6738 13841 6744 13893
rect 7743 13847 7795 13853
rect 7835 13978 7875 14705
tri 7875 14699 7881 14705 nw
rect 13434 14723 13440 14775
rect 13492 14723 13504 14775
rect 13556 14723 13562 14775
tri 13969 14771 13973 14775 ne
tri 13434 14699 13458 14723 ne
rect 13458 14699 13520 14723
tri 13520 14699 13544 14723 nw
rect 13458 14467 13510 14699
tri 13510 14689 13520 14699 nw
tri 13935 14592 13973 14630 se
rect 13973 14592 14025 14775
tri 14025 14592 14063 14630 sw
rect 13935 14540 13941 14592
rect 13993 14540 14005 14592
rect 14057 14540 14063 14592
rect 13458 14390 13510 14415
rect 13458 14312 13510 14338
rect 13458 14234 13510 14260
rect 13458 14156 13510 14182
rect 10319 14124 10371 14130
rect 13458 14098 13510 14104
rect 13970 14455 14022 14461
rect 13970 14387 14022 14403
rect 13970 14319 14022 14335
rect 13970 14251 14022 14267
rect 13970 14183 14022 14199
rect 13970 14115 14022 14131
rect 10319 14060 10371 14072
tri 7875 13978 7884 13987 sw
rect 7835 13975 7884 13978
tri 7884 13975 7887 13978 sw
rect 7835 13969 7887 13975
rect 7835 13905 7887 13917
rect 7835 13847 7887 13853
rect 5132 13804 5284 13818
rect 3059 13765 3111 13780
rect 3059 13698 3111 13713
rect 3059 13631 3111 13646
rect 3059 13564 3111 13579
rect 3059 13497 3111 13512
rect 3059 13439 3111 13445
rect 4922 13798 5002 13804
rect 4922 13746 4936 13798
rect 4988 13746 5002 13798
rect 4922 13734 5002 13746
rect 4922 13682 4936 13734
rect 4988 13682 5002 13734
rect 4922 13670 5002 13682
rect 4922 13618 4936 13670
rect 4988 13618 5002 13670
rect 4922 13606 5002 13618
rect 4922 13554 4936 13606
rect 4988 13554 5002 13606
rect 4922 13542 5002 13554
rect 4922 13490 4936 13542
rect 4988 13490 5002 13542
rect 4922 13478 5002 13490
rect 4922 13426 4936 13478
rect 4988 13426 5002 13478
rect 4922 13414 5002 13426
rect 4922 13362 4936 13414
rect 4988 13362 5002 13414
rect 4922 13350 5002 13362
rect 4922 13298 4936 13350
rect 4988 13298 5002 13350
rect 4922 13285 5002 13298
rect 4922 13233 4936 13285
rect 4988 13233 5002 13285
rect 4922 13220 5002 13233
rect 4922 13168 4936 13220
rect 4988 13168 5002 13220
rect 4922 13155 5002 13168
rect 4922 13103 4936 13155
rect 4988 13103 5002 13155
rect 4922 13090 5002 13103
rect 4922 13038 4936 13090
rect 4988 13038 5002 13090
rect 4922 13032 5002 13038
rect 5184 13752 5232 13804
rect 5132 13738 5284 13752
rect 5184 13686 5232 13738
tri 8771 13687 8823 13739 se
rect 8823 13687 9013 13739
rect 9065 13687 9077 13739
rect 9129 13687 9135 13739
rect 5132 13672 5284 13686
rect 5184 13620 5232 13672
tri 8749 13665 8771 13687 se
rect 8771 13665 8823 13687
tri 8823 13665 8845 13687 nw
rect 5132 13606 5284 13620
tri 8699 13615 8749 13665 se
rect 8749 13615 8773 13665
tri 8773 13615 8823 13665 nw
rect 5184 13554 5232 13606
tri 8675 13591 8699 13615 se
rect 8699 13591 8749 13615
tri 8749 13591 8773 13615 nw
rect 5132 13540 5284 13554
rect 5184 13488 5232 13540
rect 5132 13474 5284 13488
rect 5184 13422 5232 13474
rect 5132 13408 5284 13422
rect 5184 13356 5232 13408
rect 5132 13342 5284 13356
rect 5184 13290 5232 13342
rect 5132 13276 5284 13290
rect 5184 13224 5232 13276
rect 5132 13210 5284 13224
rect 5184 13158 5232 13210
rect 5132 13144 5284 13158
rect 5184 13092 5232 13144
rect 5132 13078 5284 13092
rect 5184 13026 5232 13078
rect 5132 13012 5284 13026
rect -175 12992 -123 12998
rect -175 12928 -123 12940
rect -175 12864 -123 12876
tri 4424 12969 4442 12987 sw
rect 4424 12917 4442 12969
tri 4442 12917 4494 12969 sw
rect 4722 12917 4728 12969
rect 4780 12917 4792 12969
rect 4844 12960 4922 12969
tri 4922 12960 4931 12969 sw
rect 5184 12960 5232 13012
rect 4844 12946 4931 12960
tri 4931 12946 4945 12960 sw
rect 5132 12946 5284 12960
rect 4844 12917 4945 12946
tri 4945 12917 4974 12946 sw
rect 4424 12894 4494 12917
tri 4494 12894 4517 12917 sw
tri 4900 12894 4923 12917 ne
rect 4923 12894 4974 12917
tri 4974 12894 4997 12917 sw
rect 5184 12894 5232 12946
rect 4424 12880 4517 12894
tri 4517 12880 4531 12894 sw
tri 4923 12880 4937 12894 ne
rect 4937 12880 4997 12894
tri 4997 12880 5011 12894 sw
rect 5132 12880 5284 12894
rect 4424 12854 4531 12880
tri 4531 12854 4557 12880 sw
tri 4937 12854 4963 12880 ne
rect 4963 12856 5011 12880
tri 5011 12856 5035 12880 sw
rect 4963 12854 5035 12856
rect 4424 12852 4861 12854
rect -175 12800 -123 12812
rect -175 12735 -123 12748
rect 4378 12800 4384 12852
rect 4436 12800 4454 12852
rect 4506 12800 4524 12852
rect 4576 12800 4594 12852
rect 4646 12800 4664 12852
rect 4716 12800 4734 12852
rect 4786 12800 4803 12852
rect 4855 12800 4861 12852
tri 4963 12843 4974 12854 ne
rect 4974 12843 5035 12854
tri 4974 12834 4983 12843 ne
rect 4378 12782 4861 12800
rect 4378 12730 4384 12782
rect 4436 12730 4454 12782
rect 4506 12730 4524 12782
rect 4576 12730 4594 12782
rect 4646 12730 4664 12782
rect 4716 12730 4734 12782
rect 4786 12730 4803 12782
rect 4855 12730 4861 12782
rect 4424 12725 4861 12730
rect 4424 12704 4527 12725
tri 4527 12704 4548 12725 nw
rect -175 12670 -123 12683
rect -175 12605 -123 12618
rect -175 12540 -123 12553
rect -175 12475 -123 12488
rect -175 12410 -123 12423
rect -175 12345 -123 12358
rect -175 12280 -123 12293
rect 4364 12698 4416 12704
rect 4364 12626 4416 12646
rect 4424 12696 4519 12704
tri 4519 12696 4527 12704 nw
rect 4424 12682 4505 12696
tri 4505 12682 4519 12696 nw
rect 4424 12630 4453 12682
tri 4453 12630 4505 12682 nw
rect 4424 12616 4439 12630
tri 4439 12616 4453 12630 nw
tri 4424 12601 4439 12616 nw
rect 4364 12553 4416 12574
rect 4364 12480 4416 12501
rect 4364 12407 4416 12428
rect 4364 12334 4416 12355
rect 4364 12261 4416 12282
rect -175 12215 -123 12228
tri -191 12163 -175 12179 se
rect 4059 12191 4065 12243
rect 4117 12191 4129 12243
rect 4181 12191 4187 12243
tri 4061 12189 4063 12191 ne
rect 4063 12189 4179 12191
tri 4179 12189 4181 12191 nw
tri 4063 12188 4064 12189 ne
rect 4064 12188 4178 12189
tri 4178 12188 4179 12189 nw
rect 4364 12188 4416 12209
tri -197 12157 -191 12163 se
rect -191 12157 -123 12163
tri 4064 12157 4095 12188 ne
tri -218 12136 -197 12157 se
rect -197 12136 -144 12157
tri -144 12136 -123 12157 nw
tri -229 12125 -218 12136 se
rect -218 12125 -155 12136
tri -155 12125 -144 12136 nw
tri -249 12105 -229 12125 se
rect -229 12105 -175 12125
tri -175 12105 -155 12125 nw
tri -281 12073 -249 12105 se
rect -249 12073 -207 12105
tri -207 12073 -175 12105 nw
tri -287 12067 -281 12073 se
rect -281 12067 -213 12073
tri -213 12067 -207 12073 nw
tri -315 12039 -287 12067 se
rect -287 12039 -241 12067
tri -241 12039 -213 12067 nw
tri -321 12033 -315 12039 se
rect -315 12033 -247 12039
tri -247 12033 -241 12039 nw
rect -201 12033 -149 12039
tri -323 12031 -321 12033 se
rect -321 12031 -249 12033
tri -249 12031 -247 12033 nw
tri -327 12027 -323 12031 se
rect -323 12027 -253 12031
tri -253 12027 -249 12031 nw
rect -327 9751 -275 12027
tri -275 12005 -253 12027 nw
rect -201 11969 -149 11981
tri 4086 11969 4095 11978 se
rect 4095 11969 4147 12188
tri 4147 12157 4178 12188 nw
rect 4364 12130 4416 12136
rect 4983 12189 5035 12843
rect 5184 12828 5232 12880
rect 5132 12814 5284 12828
rect 5184 12762 5232 12814
rect 5132 12748 5284 12762
rect 5184 12696 5232 12748
rect 5132 12682 5284 12696
rect 5184 12630 5232 12682
rect 5132 12616 5284 12630
rect 5184 12564 5232 12616
rect 5132 12550 5284 12564
rect 5184 12498 5232 12550
rect 5132 12484 5284 12498
rect 5184 12432 5232 12484
rect 5132 12418 5284 12432
rect 5184 12366 5232 12418
rect 5132 12352 5284 12366
rect 5184 12300 5232 12352
rect 5132 12286 5284 12300
rect 5184 12234 5232 12286
rect 5132 12220 5284 12234
rect 5184 12168 5232 12220
rect 5132 12162 5284 12168
tri 8648 13564 8675 13591 se
rect 8675 13564 8722 13591
tri 8722 13564 8749 13591 nw
rect 8648 13563 8721 13564
tri 8721 13563 8722 13564 nw
rect 4983 12125 5035 12137
rect 4983 12067 5035 12073
tri 4147 11969 4156 11978 sw
tri 4074 11957 4086 11969 se
rect 4086 11957 4156 11969
tri 4156 11957 4168 11969 sw
tri 8433 11962 8434 11963 se
tri 4061 11944 4074 11957 se
rect 4074 11944 4168 11957
tri 4168 11944 4181 11957 sw
rect -201 9913 -149 11917
rect 4059 11892 4065 11944
rect 4117 11892 4129 11944
rect 4181 11892 4187 11944
rect 7274 11892 7280 11944
rect 7332 11892 7344 11944
rect 7396 11892 7402 11944
tri 7316 11858 7350 11892 ne
rect 4395 11654 4401 11706
rect 4453 11654 4465 11706
rect 4517 11654 4523 11706
tri 4437 11620 4471 11654 ne
rect -201 9849 -149 9861
rect -201 9791 -149 9797
tri -275 9751 -247 9779 sw
rect -327 9699 -321 9751
rect -269 9699 -257 9751
rect -205 9699 -199 9751
rect 4471 7186 4523 11654
rect 7350 7301 7402 11892
rect 8648 11897 8700 13563
tri 8700 13542 8721 13563 nw
rect 9312 12369 9318 12421
rect 9370 12369 9382 12421
rect 9434 12369 9440 12421
tri 9364 12343 9390 12369 nw
rect 9392 12323 9444 12329
rect 9392 12259 9444 12271
rect 9392 12201 9444 12207
rect 8648 11833 8700 11845
tri 8614 8040 8648 8074 se
rect 8648 8040 8700 11781
tri 8700 8040 8734 8074 sw
rect 7350 7237 7402 7249
rect 7350 7179 7402 7185
rect 8610 7988 8616 8040
rect 8668 7988 8680 8040
rect 8732 7988 8738 8040
rect 8610 7899 8738 7988
rect 8610 7847 8616 7899
rect 8668 7847 8680 7899
rect 8732 7847 8738 7899
rect 8610 7663 8738 7847
rect 8610 7611 8616 7663
rect 8668 7611 8680 7663
rect 8732 7611 8738 7663
rect 8610 7427 8738 7611
rect 8610 7375 8616 7427
rect 8668 7375 8680 7427
rect 8732 7375 8738 7427
rect 8610 7191 8738 7375
rect 4471 7122 4523 7134
rect 4471 7064 4523 7070
rect 8610 7139 8616 7191
rect 8668 7139 8680 7191
rect 8732 7139 8738 7191
rect 8610 6955 8738 7139
rect 10319 7810 10371 14008
rect 13970 14047 14022 14063
rect 13970 13978 14022 13995
rect 13970 13909 14022 13926
tri 13944 13804 13970 13830 se
rect 13970 13804 14022 13857
tri 13933 13793 13944 13804 se
rect 13944 13794 14022 13804
rect 13944 13793 14021 13794
tri 14021 13793 14022 13794 nw
tri 13752 13739 13806 13793 se
rect 13806 13741 13969 13793
tri 13969 13741 14021 13793 nw
rect 13806 13739 13808 13741
tri 13734 13721 13752 13739 se
rect 13752 13721 13808 13739
tri 13808 13721 13828 13741 nw
tri 10528 13615 10558 13645 se
tri 10518 13605 10528 13615 se
rect 10528 13605 10558 13615
tri 10814 13615 10822 13623 sw
rect 10814 13605 10822 13615
tri 10822 13605 10832 13615 sw
rect 11892 13563 11898 13615
rect 11950 13563 11988 13615
rect 12040 13563 12078 13615
rect 12130 13563 12136 13615
rect 12553 13563 12559 13615
rect 12611 13563 12648 13615
rect 12700 13563 12706 13615
tri 10543 12814 10558 12829 ne
tri 10814 12814 10829 12829 nw
rect 11102 12318 11108 12370
rect 11160 12318 11172 12370
rect 11224 12318 11230 12370
rect 10958 12232 11010 12238
rect 10958 12168 11010 12180
rect 10685 12021 10737 12027
rect 10685 11957 10737 11969
tri 10651 8262 10685 8296 se
rect 10685 8262 10737 11905
rect 10958 11672 11010 12116
rect 10958 11608 11010 11620
rect 10958 10550 11010 11556
rect 10958 10471 11010 10498
rect 10958 10413 11010 10419
rect 10609 8210 10615 8262
rect 10667 8210 10679 8262
rect 10731 8210 10737 8262
tri 10651 8176 10685 8210 ne
tri 10680 8074 10685 8079 se
rect 10685 8074 10737 8210
tri 10646 8040 10680 8074 se
rect 10680 8057 10737 8074
rect 10680 8040 10713 8057
rect 10319 7746 10371 7758
rect 10319 7575 10371 7694
rect 10319 7511 10371 7523
rect 10319 7339 10371 7459
rect 10319 7275 10371 7287
rect 10319 7103 10371 7223
rect 10319 7039 10371 7051
rect 10319 6981 10371 6987
tri 10639 8033 10646 8040 se
rect 10646 8033 10713 8040
tri 10713 8033 10737 8057 nw
rect 8610 6903 8616 6955
rect 8668 6903 8680 6955
rect 8732 6903 8738 6955
rect 10639 6591 10691 8033
tri 10691 8011 10713 8033 nw
rect 11102 6604 11154 12318
tri 11154 12284 11188 12318 nw
tri 13700 11999 13734 12033 se
rect 13734 11999 13786 13721
tri 13786 13699 13808 13721 nw
rect 11196 11993 11248 11999
rect 13658 11947 13664 11999
rect 13716 11947 13728 11999
rect 13780 11947 13786 11999
rect 11196 11929 11248 11941
rect 11196 11589 11248 11877
rect 11196 11525 11248 11537
rect 11196 11467 11248 11473
rect 12240 8763 12592 9521
rect 12240 8711 12246 8763
rect 12298 8711 12318 8763
rect 12370 8711 12390 8763
rect 12442 8711 12462 8763
rect 12514 8711 12534 8763
rect 12586 8711 12592 8763
tri 11154 6604 11188 6638 sw
tri 10691 6591 10704 6604 sw
rect 10639 6582 10704 6591
tri 10704 6582 10713 6591 sw
tri 10639 6552 10669 6582 ne
rect 10669 6552 10713 6582
tri 10713 6552 10743 6582 sw
rect 11102 6552 11108 6604
rect 11160 6552 11175 6604
rect 11227 6552 11233 6604
rect 11650 6552 11656 6604
rect 11708 6552 11723 6604
rect 11775 6594 11987 6604
tri 11987 6594 11997 6604 sw
rect 11775 6552 11997 6594
tri 11997 6552 12039 6594 sw
tri 10669 6519 10702 6552 ne
rect 10702 6539 10743 6552
tri 10743 6539 10756 6552 sw
rect 10702 6519 10756 6539
tri 11965 6520 11997 6552 ne
rect 11997 6520 12039 6552
tri 12039 6520 12071 6552 sw
tri 10702 6517 10704 6519 ne
tri 11997 6501 12016 6520 ne
rect 12016 6501 12071 6520
rect 10704 6452 10756 6467
rect 11477 6449 11483 6501
rect 11535 6449 11550 6501
rect 11602 6449 11608 6501
tri 12016 6498 12019 6501 ne
tri 11522 6415 11556 6449 ne
rect 10704 6394 10756 6400
rect 11208 5329 11528 5330
rect 11208 5277 11214 5329
rect 11266 5277 11278 5329
rect 11330 5277 11342 5329
rect 11394 5277 11406 5329
rect 11458 5277 11470 5329
rect 11522 5277 11528 5329
rect 11208 4818 11528 5277
rect 11208 4766 11214 4818
rect 11266 4766 11278 4818
rect 11330 4766 11342 4818
rect 11394 4766 11406 4818
rect 11458 4766 11470 4818
rect 11522 4766 11528 4818
rect 11556 5179 11608 6449
rect 11556 5090 11608 5127
rect 11556 5001 11608 5038
rect 12019 5109 12071 6501
rect 12019 5042 12071 5057
rect 12019 4984 12071 4990
rect 11556 4912 11608 4949
rect 11208 3230 11214 3282
rect 11266 3230 11278 3282
rect 11330 3230 11342 3282
rect 11394 3230 11406 3282
rect 11458 3230 11470 3282
rect 11522 3230 11528 3282
rect 11208 2770 11528 3230
rect 11556 3186 11608 4860
rect 11556 3107 11608 3134
rect 11556 3027 11608 3055
rect 11556 2947 11608 2975
rect 11556 2867 11608 2895
rect 11556 2809 11608 2815
rect 11208 2718 11214 2770
rect 11266 2718 11278 2770
rect 11330 2718 11342 2770
rect 11394 2718 11406 2770
rect 11458 2718 11470 2770
rect 11522 2718 11528 2770
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1701704242
transform 0 1 8105 -1 0 7570
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1701704242
transform 0 1 8105 -1 0 7338
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1701704242
transform 0 1 8105 -1 0 7098
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_3
timestamp 1701704242
transform 0 1 4482 -1 0 7182
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_4
timestamp 1701704242
transform 0 1 5365 -1 0 7182
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_5
timestamp 1701704242
transform 0 1 6223 -1 0 7182
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_6
timestamp 1701704242
transform 0 1 7359 -1 0 7179
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_7
timestamp 1701704242
transform 0 1 10247 -1 0 7806
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_8
timestamp 1701704242
transform 0 1 10247 -1 0 7570
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_9
timestamp 1701704242
transform 0 1 10247 -1 0 7098
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_10
timestamp 1701704242
transform 0 1 10247 -1 0 7334
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_11
timestamp 1701704242
transform 0 1 8105 -1 0 7806
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_12
timestamp 1701704242
transform 0 1 12565 -1 0 7806
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_13
timestamp 1701704242
transform 0 1 12565 -1 0 7570
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_14
timestamp 1701704242
transform 0 1 12565 -1 0 7098
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_15
timestamp 1701704242
transform 0 1 12565 -1 0 7334
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_16
timestamp 1701704242
transform 0 1 10423 -1 0 7806
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_17
timestamp 1701704242
transform 0 1 10423 -1 0 7570
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_18
timestamp 1701704242
transform 0 1 10423 -1 0 7334
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_19
timestamp 1701704242
transform 0 1 10423 -1 0 7098
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_20
timestamp 1701704242
transform -1 0 4568 0 1 11981
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_21
timestamp 1701704242
transform -1 0 4824 0 1 11981
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_22
timestamp 1701704242
transform -1 0 12424 0 -1 12193
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_23
timestamp 1701704242
transform -1 0 4863 0 -1 12962
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_24
timestamp 1701704242
transform -1 0 4607 0 -1 12962
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_25
timestamp 1701704242
transform -1 0 14174 0 -1 13369
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_26
timestamp 1701704242
transform -1 0 14430 0 -1 13369
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_27
timestamp 1701704242
transform -1 0 13922 0 -1 14583
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_28
timestamp 1701704242
transform -1 0 14178 0 -1 12168
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_29
timestamp 1701704242
transform -1 0 13922 0 -1 12168
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_30
timestamp 1701704242
transform -1 0 14178 0 -1 14583
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_31
timestamp 1701704242
transform -1 0 13662 0 -1 13369
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_32
timestamp 1701704242
transform -1 0 13918 0 -1 13369
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_33
timestamp 1701704242
transform -1 0 355 0 -1 12042
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_34
timestamp 1701704242
transform -1 0 33 0 -1 12042
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_35
timestamp 1701704242
transform -1 0 -223 0 -1 12042
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_36
timestamp 1701704242
transform -1 0 4114 0 -1 12390
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_37
timestamp 1701704242
transform -1 0 3878 0 -1 12390
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_38
timestamp 1701704242
transform -1 0 3406 0 -1 12390
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_39
timestamp 1701704242
transform -1 0 3642 0 -1 12390
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_40
timestamp 1701704242
transform -1 0 4114 0 -1 14532
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_41
timestamp 1701704242
transform -1 0 3878 0 -1 14532
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_42
timestamp 1701704242
transform -1 0 3647 0 -1 14532
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_43
timestamp 1701704242
transform -1 0 3406 0 -1 14532
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_44
timestamp 1701704242
transform -1 0 12168 0 -1 12193
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_45
timestamp 1701704242
transform 0 -1 11873 1 0 3074
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_46
timestamp 1701704242
transform 0 -1 11873 1 0 2818
box 0 0 1 1
use nDFbentRes_CDNS_524688791851262  nDFbentRes_CDNS_524688791851262_0
timestamp 1701704242
transform -1 0 9019 0 1 13680
box -68 -1106 3474 92
use nDFbentRes_CDNS_524688791851263  nDFbentRes_CDNS_524688791851263_0
timestamp 1701704242
transform -1 0 8709 0 1 14074
box -68 -266 2912 92
use nfet_CDNS_524688791851264  nfet_CDNS_524688791851264_0
timestamp 1701704242
transform 0 -1 11791 1 0 4819
box -79 -26 535 626
use nfet_CDNS_524688791851265  nfet_CDNS_524688791851265_0
timestamp 1701704242
transform 0 -1 11791 1 0 2771
box -79 -26 535 626
use nfet_CDNS_524688791851266  nfet_CDNS_524688791851266_0
timestamp 1701704242
transform 0 -1 4428 1 0 7041
box -79 -32 259 232
use nfet_CDNS_524688791851266  nfet_CDNS_524688791851266_1
timestamp 1701704242
transform 0 -1 5311 1 0 7041
box -79 -32 259 232
use nfet_CDNS_524688791851266  nfet_CDNS_524688791851266_2
timestamp 1701704242
transform 0 -1 6169 1 0 7041
box -79 -32 259 232
use nfet_CDNS_524688791851266  nfet_CDNS_524688791851266_3
timestamp 1701704242
transform 0 -1 7305 1 0 7041
box -79 -32 259 232
use nfet_CDNS_524688791851267  nfet_CDNS_524688791851267_0
timestamp 1701704242
transform 0 -1 10193 1 0 7193
box -79 -32 259 2032
use nfet_CDNS_524688791851267  nfet_CDNS_524688791851267_1
timestamp 1701704242
transform 0 -1 12511 1 0 7193
box -79 -32 259 2032
use nfet_CDNS_524688791851267  nfet_CDNS_524688791851267_2
timestamp 1701704242
transform 1 0 3501 0 1 12444
box -79 -32 259 2032
use nfet_CDNS_524688791851268  nfet_CDNS_524688791851268_0
timestamp 1701704242
transform 0 -1 10193 1 0 7665
box -79 -32 259 2032
use nfet_CDNS_524688791851268  nfet_CDNS_524688791851268_1
timestamp 1701704242
transform 0 -1 10193 1 0 6957
box -79 -32 259 2032
use nfet_CDNS_524688791851268  nfet_CDNS_524688791851268_2
timestamp 1701704242
transform 0 -1 12511 1 0 7665
box -79 -32 259 2032
use nfet_CDNS_524688791851268  nfet_CDNS_524688791851268_3
timestamp 1701704242
transform 0 -1 12511 1 0 6957
box -79 -32 259 2032
use nfet_CDNS_524688791851268  nfet_CDNS_524688791851268_4
timestamp 1701704242
transform 1 0 3265 0 1 12444
box -79 -32 259 2032
use nfet_CDNS_524688791851268  nfet_CDNS_524688791851268_5
timestamp 1701704242
transform 1 0 3973 0 1 12444
box -79 -32 259 2032
use nfet_CDNS_524688791851269  nfet_CDNS_524688791851269_0
timestamp 1701704242
transform 0 -1 10193 1 0 7429
box -79 -32 259 2032
use nfet_CDNS_524688791851269  nfet_CDNS_524688791851269_1
timestamp 1701704242
transform 0 -1 12511 1 0 7429
box -79 -32 259 2032
use nfet_CDNS_524688791851269  nfet_CDNS_524688791851269_2
timestamp 1701704242
transform 1 0 3737 0 1 12444
box -79 -32 259 2032
use nfet_CDNS_524688791851270  nfet_CDNS_524688791851270_0
timestamp 1701704242
transform 1 0 4421 0 -1 12676
box -79 -26 535 626
use nfet_CDNS_524688791851270  nfet_CDNS_524688791851270_1
timestamp 1701704242
transform 1 0 4454 0 1 13013
box -79 -26 535 626
use pfet_CDNS_524688791851272  pfet_CDNS_524688791851272_0
timestamp 1701704242
transform 1 0 -464 0 -1 14250
box -161 -36 2665 636
use pfet_CDNS_524688791851274  pfet_CDNS_524688791851274_0
timestamp 1701704242
transform 1 0 12015 0 -1 13243
box -89 -36 545 1036
use pfet_CDNS_524688791851275  pfet_CDNS_524688791851275_0
timestamp 1701704242
transform 1 0 -376 0 1 12173
box -89 -36 545 1036
use pfet_CDNS_524688791851276  pfet_CDNS_524688791851276_0
timestamp 1701704242
transform 1 0 254 0 1 12173
box -89 -36 189 1036
use pfet_CDNS_524688791851277  pfet_CDNS_524688791851277_0
timestamp 1701704242
transform 1 0 13513 0 1 12222
box -89 -36 1057 1036
use pfet_CDNS_524688791851277  pfet_CDNS_524688791851277_1
timestamp 1701704242
transform 1 0 13513 0 1 13495
box -89 -36 1057 1036
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_0
timestamp 1701704242
transform 0 1 12304 -1 0 12211
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_1
timestamp 1701704242
transform 0 1 4743 -1 0 12981
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_2
timestamp 1701704242
transform 0 1 4487 -1 0 12981
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_3
timestamp 1701704242
transform 0 1 14054 -1 0 13385
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_4
timestamp 1701704242
transform 0 1 14310 -1 0 13385
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_5
timestamp 1701704242
transform 0 1 14058 -1 0 12184
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_6
timestamp 1701704242
transform 0 1 13802 -1 0 12184
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_7
timestamp 1701704242
transform 0 1 13798 -1 0 13385
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_8
timestamp 1701704242
transform 0 1 14058 -1 0 14599
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_9
timestamp 1701704242
transform 0 1 13802 -1 0 14599
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_10
timestamp 1701704242
transform 0 1 13542 -1 0 13385
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_11
timestamp 1701704242
transform 0 1 235 -1 0 12058
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_12
timestamp 1701704242
transform 0 1 -87 -1 0 12058
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_13
timestamp 1701704242
transform 0 1 -343 -1 0 12058
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_14
timestamp 1701704242
transform 0 1 3994 -1 0 12406
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_15
timestamp 1701704242
transform 0 1 3758 -1 0 12406
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_16
timestamp 1701704242
transform 0 1 3286 -1 0 12406
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_17
timestamp 1701704242
transform 0 1 3522 -1 0 12406
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_18
timestamp 1701704242
transform 0 1 3758 -1 0 14548
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_19
timestamp 1701704242
transform 0 1 3994 -1 0 14548
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_20
timestamp 1701704242
transform 0 1 3286 -1 0 14548
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_21
timestamp 1701704242
transform 0 1 3522 -1 0 14548
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_22
timestamp 1701704242
transform 0 1 12048 -1 0 12211
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_23
timestamp 1701704242
transform -1 0 11889 0 -1 2938
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_24
timestamp 1701704242
transform -1 0 11889 0 -1 3194
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_25
timestamp 1701704242
transform 0 1 4448 1 0 11965
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_26
timestamp 1701704242
transform 0 1 4704 1 0 11965
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_27
timestamp 1701704242
transform 1 0 8089 0 1 7450
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_28
timestamp 1701704242
transform 1 0 8089 0 1 6978
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_29
timestamp 1701704242
transform 1 0 8089 0 1 7214
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_30
timestamp 1701704242
transform 1 0 4466 0 1 7059
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_31
timestamp 1701704242
transform 1 0 5349 0 1 7059
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_32
timestamp 1701704242
transform 1 0 6207 0 1 7059
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_33
timestamp 1701704242
transform 1 0 7343 0 1 7059
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_34
timestamp 1701704242
transform 1 0 10231 0 1 7686
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_35
timestamp 1701704242
transform 1 0 10231 0 1 7450
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_36
timestamp 1701704242
transform 1 0 10231 0 1 6978
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_37
timestamp 1701704242
transform 1 0 10231 0 1 7214
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_38
timestamp 1701704242
transform 1 0 8089 0 1 7686
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_39
timestamp 1701704242
transform 1 0 12549 0 1 7686
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_40
timestamp 1701704242
transform 1 0 12549 0 1 7450
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_41
timestamp 1701704242
transform 1 0 12549 0 1 6978
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_42
timestamp 1701704242
transform 1 0 12549 0 1 7214
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_43
timestamp 1701704242
transform 1 0 10407 0 1 7450
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_44
timestamp 1701704242
transform 1 0 10407 0 1 7686
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_45
timestamp 1701704242
transform 1 0 10407 0 1 6978
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_46
timestamp 1701704242
transform 1 0 10407 0 1 7214
box 0 0 1 1
use PYL1_CDNS_52468879185309  PYL1_CDNS_52468879185309_0
timestamp 1701704242
transform -1 0 11889 0 -1 5182
box 0 0 1 1
use sky130_fd_io__sio_biasgen_res  sky130_fd_io__sio_biasgen_res_0
timestamp 1701704242
transform 1 0 2122 0 1 7963
box -71 -20 10905 2779
<< labels >>
flabel comment s 8330 6674 8330 6674 0 FreeSans 400 0 0 0 condiode
flabel comment s 7225 6737 7225 6737 0 FreeSans 400 0 0 0 condiode
flabel comment s 6223 6738 6223 6738 0 FreeSans 400 0 0 0 condiode
flabel comment s 5238 6767 5238 6767 0 FreeSans 400 0 0 0 condiode
flabel comment s 4354 6731 4354 6731 0 FreeSans 400 0 0 0 condiode
flabel comment s 7225 6450 7225 6450 0 FreeSans 400 0 0 0 condiode
flabel metal1 s -597 13466 -505 13572 3 FreeSans 520 0 0 0 vpwr
port 2 nsew
flabel metal1 s 7177 6854 7269 6960 3 FreeSans 520 0 0 0 vgnd
port 3 nsew
flabel metal1 s 5035 12731 5127 12837 3 FreeSans 520 0 0 0 vgnd
port 3 nsew
flabel metal1 s 14514 14720 14574 14766 3 FreeSans 520 0 0 0 vpwr
port 2 nsew
flabel metal1 s 9965 10257 10025 10303 3 FreeSans 520 0 0 0 vpwr
port 2 nsew
flabel metal1 s 4905 14458 5023 14504 3 FreeSans 520 0 0 0 ngate
port 4 nsew
flabel metal1 s 10964 10414 11010 10519 3 FreeSans 520 0 0 0 ie_diff_sel_n
port 5 nsew
flabel locali s 11923 5449 11959 5555 3 FreeSans 520 0 0 0 vgnd
port 3 nsew
flabel locali s 9231 12813 9265 12919 3 FreeSans 520 0 0 0 vgnd
port 3 nsew
flabel metal2 s 11208 5224 11300 5330 3 FreeSans 520 0 0 0 vgnd
port 3 nsew
flabel metal2 s 11208 3176 11300 3282 3 FreeSans 520 0 0 0 vgnd
port 3 nsew
flabel metal2 s 11102 6742 11154 6860 3 FreeSans 520 0 0 0 ie_diff_sel_h_n
port 6 nsew
<< properties >>
string GDS_END 86825752
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86621784
string path 77.125 335.975 77.125 364.100 
<< end >>
