magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< pwell >>
rect -76 -26 332 1026
<< mvnmos >>
rect 0 0 100 1000
rect 156 0 256 1000
<< mvndiff >>
rect -50 0 0 1000
rect 256 0 306 1000
<< poly >>
rect 0 1000 100 1026
rect 0 -26 100 0
rect 156 1000 256 1026
rect 156 -26 256 0
<< locali >>
rect -45 -4 -11 946
rect 111 -4 145 946
rect 267 -4 301 946
use hvDFL1sd2_CDNS_524688791858  hvDFL1sd2_CDNS_524688791858_0
timestamp 1701704242
transform 1 0 100 0 1 0
box -26 -26 82 1026
use hvDFL1sd_CDNS_5246887918592  hvDFL1sd_CDNS_5246887918592_0
timestamp 1701704242
transform -1 0 0 0 1 0
box -26 -26 79 1026
use hvDFL1sd_CDNS_5246887918592  hvDFL1sd_CDNS_5246887918592_1
timestamp 1701704242
transform 1 0 256 0 1 0
box -26 -26 79 1026
<< labels >>
flabel comment s -28 471 -28 471 0 FreeSans 300 0 0 0 S
flabel comment s 128 471 128 471 0 FreeSans 300 0 0 0 D
flabel comment s 284 471 284 471 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 96476004
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 96474616
<< end >>
