magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< metal2 >>
rect 0 465 296 474
rect 0 0 296 9
<< via2 >>
rect 0 9 296 465
<< metal3 >>
rect -5 465 301 470
rect -5 9 0 465
rect 296 9 301 465
rect -5 4 301 9
<< properties >>
string GDS_END 88079842
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 88078174
<< end >>
