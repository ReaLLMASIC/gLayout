magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -122 -66 690 366
<< mvpmos >>
rect 0 0 100 300
rect 156 0 256 300
rect 312 0 412 300
rect 468 0 568 300
<< mvpdiff >>
rect -50 0 0 300
rect 568 0 618 300
<< poly >>
rect 0 300 100 332
rect 0 -32 100 0
rect 156 300 256 332
rect 156 -32 256 0
rect 312 300 412 332
rect 312 -32 412 0
rect 468 300 568 332
rect 468 -32 568 0
<< metal1 >>
rect -51 -16 -5 258
rect 105 -16 151 258
rect 261 -16 307 258
rect 417 -16 463 258
rect 573 -16 619 258
use hvDFM1sd2_CDNS_52468879185879  hvDFM1sd2_CDNS_52468879185879_0
timestamp 1701704242
transform -1 0 0 0 1 0
box -36 -36 92 336
use hvDFM1sd2_CDNS_52468879185879  hvDFM1sd2_CDNS_52468879185879_1
timestamp 1701704242
transform 1 0 568 0 1 0
box -36 -36 92 336
use hvDFM1sd2_CDNS_52468879185879  hvDFM1sd2_CDNS_52468879185879_2
timestamp 1701704242
transform 1 0 412 0 1 0
box -36 -36 92 336
use hvDFM1sd2_CDNS_52468879185879  hvDFM1sd2_CDNS_52468879185879_3
timestamp 1701704242
transform 1 0 256 0 1 0
box -36 -36 92 336
use hvDFM1sd2_CDNS_52468879185879  hvDFM1sd2_CDNS_52468879185879_4
timestamp 1701704242
transform 1 0 100 0 1 0
box -36 -36 92 336
<< labels >>
flabel comment s -28 121 -28 121 0 FreeSans 300 0 0 0 S
flabel comment s 128 121 128 121 0 FreeSans 300 0 0 0 D
flabel comment s 284 121 284 121 0 FreeSans 300 0 0 0 S
flabel comment s 440 121 440 121 0 FreeSans 300 0 0 0 D
flabel comment s 596 121 596 121 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 7599600
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 7597078
<< end >>
