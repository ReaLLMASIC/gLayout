magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -38 261 406 582
<< pwell >>
rect 1 21 367 183
rect 29 -17 63 21
<< scnmos >>
rect 79 47 289 157
<< scpmoshvt >>
rect 79 323 289 497
<< ndiff >>
rect 27 119 79 157
rect 27 85 35 119
rect 69 85 79 119
rect 27 47 79 85
rect 289 119 341 157
rect 289 85 299 119
rect 333 85 341 119
rect 289 47 341 85
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 383 79 451
rect 27 349 35 383
rect 69 349 79 383
rect 27 323 79 349
rect 289 485 341 497
rect 289 451 299 485
rect 333 451 341 485
rect 289 383 341 451
rect 289 349 299 383
rect 333 349 341 383
rect 289 323 341 349
<< ndiffc >>
rect 35 85 69 119
rect 299 85 333 119
<< pdiffc >>
rect 35 451 69 485
rect 35 349 69 383
rect 299 451 333 485
rect 299 349 333 383
<< poly >>
rect 79 497 289 523
rect 79 297 289 323
rect 79 291 163 297
rect 21 275 163 291
rect 21 241 37 275
rect 71 241 163 275
rect 21 225 163 241
rect 205 239 347 255
rect 205 205 297 239
rect 331 205 347 239
rect 205 189 347 205
rect 205 183 289 189
rect 79 157 289 183
rect 79 21 289 47
<< polycont >>
rect 37 241 71 275
rect 297 205 331 239
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 368 561
rect 17 485 351 527
rect 17 451 35 485
rect 69 451 299 485
rect 333 451 351 485
rect 17 383 351 451
rect 17 349 35 383
rect 69 349 299 383
rect 333 349 351 383
rect 17 309 351 349
rect 17 241 37 275
rect 71 241 167 275
rect 17 171 167 241
rect 201 239 351 309
rect 201 205 297 239
rect 331 205 351 239
rect 17 119 351 171
rect 17 85 35 119
rect 69 85 299 119
rect 333 85 351 119
rect 17 17 351 85
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 368 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
<< metal1 >>
rect 0 561 368 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 368 561
rect 0 496 368 527
rect 0 17 368 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 368 17
rect 0 -48 368 -17
<< labels >>
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 1 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 4 nsew power bidirectional abutment
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 3 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 2 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 decap_4
rlabel metal1 s 0 -48 368 48 1 VGND
port 1 nsew ground bidirectional abutment
rlabel metal1 s 0 496 368 592 1 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 368 544
string GDS_END 3328444
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3325710
string LEFclass CORE SPACER
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 9.200 0.000 
<< end >>
