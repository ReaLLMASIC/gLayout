magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< nwell >>
rect 1049 336 1215 668
rect 780 236 1215 336
<< pwell >>
rect 1107 -76 1193 176
<< mvpsubdiff >>
rect 1133 126 1167 150
rect 1133 8 1167 92
rect 1133 -50 1167 -26
<< mvnsubdiff >>
rect 1115 578 1149 602
rect 1115 505 1149 544
rect 1115 432 1149 471
rect 1115 360 1149 398
rect 1115 302 1149 326
<< mvpsubdiffcont >>
rect 1133 92 1167 126
rect 1133 -26 1167 8
<< mvnsubdiffcont >>
rect 1115 544 1149 578
rect 1115 471 1149 505
rect 1115 398 1149 432
rect 1115 326 1149 360
<< poly >>
rect 888 356 988 376
rect 888 340 1093 356
rect 888 306 975 340
rect 1009 306 1043 340
rect 1077 306 1093 340
rect 888 290 1093 306
rect 119 252 531 276
rect 619 270 719 276
rect 119 218 135 252
rect 169 218 219 252
rect 253 218 302 252
rect 336 218 531 252
rect 119 150 531 218
rect 573 254 719 270
rect 573 220 589 254
rect 623 220 657 254
rect 691 220 719 254
rect 573 204 719 220
rect 619 150 719 204
rect 873 232 1007 248
rect 873 198 889 232
rect 923 198 957 232
rect 991 198 1007 232
rect 873 182 1007 198
rect 906 176 1006 182
<< polycont >>
rect 975 306 1009 340
rect 1043 306 1077 340
rect 135 218 169 252
rect 219 218 253 252
rect 302 218 336 252
rect 589 220 623 254
rect 657 220 691 254
rect 889 198 923 232
rect 957 198 991 232
<< locali >>
rect 230 640 576 674
rect 230 606 264 640
rect 542 606 576 640
rect 74 405 108 471
rect 386 270 420 606
rect 725 271 773 606
rect 807 404 843 606
rect 999 578 1149 606
rect 999 544 1115 578
rect 999 505 1149 544
rect 999 483 1115 505
rect 911 471 1115 483
rect 911 432 1149 471
rect 386 254 691 270
rect 119 218 135 252
rect 169 218 219 252
rect 253 218 302 252
rect 336 218 352 252
rect 386 220 589 254
rect 623 220 657 254
rect 386 204 691 220
rect 74 62 108 130
rect 386 36 420 204
rect 725 170 759 271
rect 807 237 855 404
rect 911 398 1115 432
rect 911 390 1149 398
rect 911 388 950 390
rect 907 384 950 388
rect 905 380 950 384
rect 902 378 949 380
rect 902 374 946 378
rect 902 370 944 374
rect 902 248 941 370
rect 1115 360 1149 390
rect 975 340 1077 356
rect 1009 306 1043 340
rect 975 290 1077 306
rect 1115 302 1149 326
rect 659 136 759 170
rect 793 182 855 237
rect 889 232 991 248
rect 923 198 957 232
rect 889 182 991 198
rect 230 2 264 36
rect 558 2 592 36
rect 230 -32 592 2
rect 659 2 696 136
rect 793 102 827 182
rect 1025 148 1077 290
rect 764 36 827 102
rect 1033 93 1077 148
rect 1017 27 1077 93
rect 659 -32 861 2
rect 1033 -54 1077 27
rect 1133 126 1167 150
rect 1133 8 1167 92
rect 1133 -50 1167 -26
use nfet_CDNS_52468879185506  nfet_CDNS_52468879185506_0
timestamp 1701704242
transform -1 0 1006 0 1 -50
box -79 -26 179 226
use nfet_CDNS_52468879185507  nfet_CDNS_52468879185507_0
timestamp 1701704242
transform 1 0 619 0 1 40
box -95 -26 179 110
use nfet_CDNS_52468879185508  nfet_CDNS_52468879185508_0
timestamp 1701704242
transform 1 0 431 0 1 40
box -79 -26 195 110
use nfet_CDNS_52468879185509  nfet_CDNS_52468879185509_0
timestamp 1701704242
transform 1 0 275 0 1 40
box -79 -26 179 110
use nfet_CDNS_52468879185510  nfet_CDNS_52468879185510_0
timestamp 1701704242
transform 1 0 119 0 1 40
box -79 -26 179 110
use pfet_CDNS_52468879185502  pfet_CDNS_52468879185502_0
timestamp 1701704242
transform 1 0 619 0 -1 602
box -154 -66 222 366
use pfet_CDNS_52468879185503  pfet_CDNS_52468879185503_0
timestamp 1701704242
transform 1 0 275 0 -1 602
box -119 -66 375 366
use pfet_CDNS_52468879185504  pfet_CDNS_52468879185504_0
timestamp 1701704242
transform -1 0 988 0 -1 602
box -119 -66 219 266
use pfet_CDNS_52468879185505  pfet_CDNS_52468879185505_0
timestamp 1701704242
transform 1 0 119 0 -1 602
box -119 -66 219 366
<< labels >>
flabel locali s 434 658 434 658 7 FreeSans 200 0 0 0 int_p
flabel locali s 433 -12 433 -12 7 FreeSans 200 0 0 0 int_n
flabel locali s 1133 66 1167 150 0 FreeSans 200 0 0 0 vgnd
port 2 nsew
flabel locali s 543 218 559 252 3 FreeSans 200 0 0 0 out
port 3 nsew
flabel locali s 1063 405 1097 471 0 FreeSans 200 0 0 0 vcc_io
port 4 nsew
flabel locali s 119 218 135 252 3 FreeSans 200 0 0 0 in
port 5 nsew
flabel locali s 74 62 108 128 3 FreeSans 200 0 0 0 vgnd
port 2 nsew
flabel locali s 74 405 108 471 3 FreeSans 200 0 0 0 vcc_io
port 4 nsew
flabel locali s 1017 27 1051 93 3 FreeSans 200 180 0 0 vgnd
port 2 nsew
<< properties >>
string GDS_END 70902954
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 70897750
string path 28.300 15.700 28.300 6.900 
<< end >>
