magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< pwell >>
rect 10 30 1366 2082
<< mvnnmos >>
tri 798 2036 818 2056 ne
tri 798 56 818 76 se
rect 818 56 998 2056
tri 998 2036 1018 2056 nw
tri 998 56 1018 76 sw
<< mvndiff >>
rect 36 2036 798 2056
tri 798 2036 818 2056 sw
rect 36 1957 818 2036
rect 36 155 176 1957
rect 278 155 818 1957
rect 36 76 818 155
rect 36 56 798 76
tri 798 56 818 76 nw
tri 998 2036 1018 2056 se
rect 1018 2036 1340 2056
rect 998 1957 1340 2036
rect 998 155 1101 1957
rect 1203 155 1340 1957
rect 998 76 1340 155
tri 998 56 1018 76 ne
rect 1018 56 1340 76
<< mvndiffc >>
rect 176 155 278 1957
rect 1101 155 1203 1957
<< poly >>
rect 778 2076 1038 2199
tri 778 2056 798 2076 ne
rect 798 2056 1018 2076
tri 1018 2056 1038 2076 nw
tri 778 36 798 56 se
rect 798 36 1018 56
tri 1018 36 1038 56 sw
rect 778 -82 1038 36
<< locali >>
rect 36 1957 283 2056
rect 36 1923 174 1957
rect 280 1923 283 1957
rect 36 1884 176 1923
rect 278 1884 283 1923
rect 36 1850 174 1884
rect 280 1850 283 1884
rect 36 1811 176 1850
rect 278 1811 283 1850
rect 36 1777 174 1811
rect 280 1777 283 1811
rect 36 1738 176 1777
rect 278 1738 283 1777
rect 36 1704 174 1738
rect 280 1704 283 1738
rect 36 1665 176 1704
rect 278 1665 283 1704
rect 36 1631 174 1665
rect 280 1631 283 1665
rect 36 1592 176 1631
rect 278 1592 283 1631
rect 36 1558 174 1592
rect 280 1558 283 1592
rect 36 1519 176 1558
rect 278 1519 283 1558
rect 36 1485 174 1519
rect 280 1485 283 1519
rect 36 1446 176 1485
rect 278 1446 283 1485
rect 36 1412 174 1446
rect 280 1412 283 1446
rect 36 1373 176 1412
rect 278 1373 283 1412
rect 36 1339 174 1373
rect 280 1339 283 1373
rect 36 1299 176 1339
rect 278 1299 283 1339
rect 36 1265 174 1299
rect 280 1265 283 1299
rect 36 1225 176 1265
rect 278 1225 283 1265
rect 36 1191 174 1225
rect 280 1191 283 1225
rect 36 1151 176 1191
rect 278 1151 283 1191
rect 36 1117 174 1151
rect 280 1117 283 1151
rect 36 1077 176 1117
rect 278 1077 283 1117
rect 36 1043 174 1077
rect 280 1043 283 1077
rect 36 1003 176 1043
rect 278 1003 283 1043
rect 36 969 174 1003
rect 280 969 283 1003
rect 36 929 176 969
rect 278 929 283 969
rect 36 895 174 929
rect 280 895 283 929
rect 36 855 176 895
rect 278 855 283 895
rect 36 821 174 855
rect 280 821 283 855
rect 36 781 176 821
rect 278 781 283 821
rect 36 747 174 781
rect 280 747 283 781
rect 36 707 176 747
rect 278 707 283 747
rect 36 673 174 707
rect 280 673 283 707
rect 36 633 176 673
rect 278 633 283 673
rect 36 599 174 633
rect 280 599 283 633
rect 36 559 176 599
rect 278 559 283 599
rect 36 525 174 559
rect 280 525 283 559
rect 36 485 176 525
rect 278 485 283 525
rect 36 451 174 485
rect 280 451 283 485
rect 36 411 176 451
rect 278 411 283 451
rect 36 377 174 411
rect 280 377 283 411
rect 36 337 176 377
rect 278 337 283 377
rect 36 303 174 337
rect 280 303 283 337
rect 36 263 176 303
rect 278 263 283 303
rect 36 229 174 263
rect 280 229 283 263
rect 36 189 176 229
rect 278 189 283 229
rect 36 155 174 189
rect 280 155 283 189
rect 36 56 283 155
rect 876 1957 1340 2056
rect 876 1923 1099 1957
rect 1205 1923 1340 1957
rect 876 1884 1101 1923
rect 1203 1884 1340 1923
rect 876 1850 1099 1884
rect 1205 1850 1340 1884
rect 876 1811 1101 1850
rect 1203 1811 1340 1850
rect 876 1777 1099 1811
rect 1205 1777 1340 1811
rect 876 1738 1101 1777
rect 1203 1738 1340 1777
rect 876 1704 1099 1738
rect 1205 1704 1340 1738
rect 876 1665 1101 1704
rect 1203 1665 1340 1704
rect 876 1631 1099 1665
rect 1205 1631 1340 1665
rect 876 1592 1101 1631
rect 1203 1592 1340 1631
rect 876 1558 1099 1592
rect 1205 1558 1340 1592
rect 876 1519 1101 1558
rect 1203 1519 1340 1558
rect 876 1485 1099 1519
rect 1205 1485 1340 1519
rect 876 1446 1101 1485
rect 1203 1446 1340 1485
rect 876 1412 1099 1446
rect 1205 1412 1340 1446
rect 876 1373 1101 1412
rect 1203 1373 1340 1412
rect 876 1339 1099 1373
rect 1205 1339 1340 1373
rect 876 1299 1101 1339
rect 1203 1299 1340 1339
rect 876 1265 1099 1299
rect 1205 1265 1340 1299
rect 876 1225 1101 1265
rect 1203 1225 1340 1265
rect 876 1191 1099 1225
rect 1205 1191 1340 1225
rect 876 1151 1101 1191
rect 1203 1151 1340 1191
rect 876 1117 1099 1151
rect 1205 1117 1340 1151
rect 876 1077 1101 1117
rect 1203 1077 1340 1117
rect 876 1043 1099 1077
rect 1205 1043 1340 1077
rect 876 1003 1101 1043
rect 1203 1003 1340 1043
rect 876 969 1099 1003
rect 1205 969 1340 1003
rect 876 929 1101 969
rect 1203 929 1340 969
rect 876 895 1099 929
rect 1205 895 1340 929
rect 876 855 1101 895
rect 1203 855 1340 895
rect 876 821 1099 855
rect 1205 821 1340 855
rect 876 781 1101 821
rect 1203 781 1340 821
rect 876 747 1099 781
rect 1205 747 1340 781
rect 876 707 1101 747
rect 1203 707 1340 747
rect 876 673 1099 707
rect 1205 673 1340 707
rect 876 633 1101 673
rect 1203 633 1340 673
rect 876 599 1099 633
rect 1205 599 1340 633
rect 876 559 1101 599
rect 1203 559 1340 599
rect 876 525 1099 559
rect 1205 525 1340 559
rect 876 485 1101 525
rect 1203 485 1340 525
rect 876 451 1099 485
rect 1205 451 1340 485
rect 876 411 1101 451
rect 1203 411 1340 451
rect 876 377 1099 411
rect 1205 377 1340 411
rect 876 337 1101 377
rect 1203 337 1340 377
rect 876 303 1099 337
rect 1205 303 1340 337
rect 876 263 1101 303
rect 1203 263 1340 303
rect 876 229 1099 263
rect 1205 229 1340 263
rect 876 189 1101 229
rect 1203 189 1340 229
rect 876 155 1099 189
rect 1205 155 1340 189
rect 876 56 1340 155
<< viali >>
rect 174 1923 176 1957
rect 176 1923 208 1957
rect 246 1923 278 1957
rect 278 1923 280 1957
rect 174 1850 176 1884
rect 176 1850 208 1884
rect 246 1850 278 1884
rect 278 1850 280 1884
rect 174 1777 176 1811
rect 176 1777 208 1811
rect 246 1777 278 1811
rect 278 1777 280 1811
rect 174 1704 176 1738
rect 176 1704 208 1738
rect 246 1704 278 1738
rect 278 1704 280 1738
rect 174 1631 176 1665
rect 176 1631 208 1665
rect 246 1631 278 1665
rect 278 1631 280 1665
rect 174 1558 176 1592
rect 176 1558 208 1592
rect 246 1558 278 1592
rect 278 1558 280 1592
rect 174 1485 176 1519
rect 176 1485 208 1519
rect 246 1485 278 1519
rect 278 1485 280 1519
rect 174 1412 176 1446
rect 176 1412 208 1446
rect 246 1412 278 1446
rect 278 1412 280 1446
rect 174 1339 176 1373
rect 176 1339 208 1373
rect 246 1339 278 1373
rect 278 1339 280 1373
rect 174 1265 176 1299
rect 176 1265 208 1299
rect 246 1265 278 1299
rect 278 1265 280 1299
rect 174 1191 176 1225
rect 176 1191 208 1225
rect 246 1191 278 1225
rect 278 1191 280 1225
rect 174 1117 176 1151
rect 176 1117 208 1151
rect 246 1117 278 1151
rect 278 1117 280 1151
rect 174 1043 176 1077
rect 176 1043 208 1077
rect 246 1043 278 1077
rect 278 1043 280 1077
rect 174 969 176 1003
rect 176 969 208 1003
rect 246 969 278 1003
rect 278 969 280 1003
rect 174 895 176 929
rect 176 895 208 929
rect 246 895 278 929
rect 278 895 280 929
rect 174 821 176 855
rect 176 821 208 855
rect 246 821 278 855
rect 278 821 280 855
rect 174 747 176 781
rect 176 747 208 781
rect 246 747 278 781
rect 278 747 280 781
rect 174 673 176 707
rect 176 673 208 707
rect 246 673 278 707
rect 278 673 280 707
rect 174 599 176 633
rect 176 599 208 633
rect 246 599 278 633
rect 278 599 280 633
rect 174 525 176 559
rect 176 525 208 559
rect 246 525 278 559
rect 278 525 280 559
rect 174 451 176 485
rect 176 451 208 485
rect 246 451 278 485
rect 278 451 280 485
rect 174 377 176 411
rect 176 377 208 411
rect 246 377 278 411
rect 278 377 280 411
rect 174 303 176 337
rect 176 303 208 337
rect 246 303 278 337
rect 278 303 280 337
rect 174 229 176 263
rect 176 229 208 263
rect 246 229 278 263
rect 278 229 280 263
rect 174 155 176 189
rect 176 155 208 189
rect 246 155 278 189
rect 278 155 280 189
rect 1099 1923 1101 1957
rect 1101 1923 1133 1957
rect 1171 1923 1203 1957
rect 1203 1923 1205 1957
rect 1099 1850 1101 1884
rect 1101 1850 1133 1884
rect 1171 1850 1203 1884
rect 1203 1850 1205 1884
rect 1099 1777 1101 1811
rect 1101 1777 1133 1811
rect 1171 1777 1203 1811
rect 1203 1777 1205 1811
rect 1099 1704 1101 1738
rect 1101 1704 1133 1738
rect 1171 1704 1203 1738
rect 1203 1704 1205 1738
rect 1099 1631 1101 1665
rect 1101 1631 1133 1665
rect 1171 1631 1203 1665
rect 1203 1631 1205 1665
rect 1099 1558 1101 1592
rect 1101 1558 1133 1592
rect 1171 1558 1203 1592
rect 1203 1558 1205 1592
rect 1099 1485 1101 1519
rect 1101 1485 1133 1519
rect 1171 1485 1203 1519
rect 1203 1485 1205 1519
rect 1099 1412 1101 1446
rect 1101 1412 1133 1446
rect 1171 1412 1203 1446
rect 1203 1412 1205 1446
rect 1099 1339 1101 1373
rect 1101 1339 1133 1373
rect 1171 1339 1203 1373
rect 1203 1339 1205 1373
rect 1099 1265 1101 1299
rect 1101 1265 1133 1299
rect 1171 1265 1203 1299
rect 1203 1265 1205 1299
rect 1099 1191 1101 1225
rect 1101 1191 1133 1225
rect 1171 1191 1203 1225
rect 1203 1191 1205 1225
rect 1099 1117 1101 1151
rect 1101 1117 1133 1151
rect 1171 1117 1203 1151
rect 1203 1117 1205 1151
rect 1099 1043 1101 1077
rect 1101 1043 1133 1077
rect 1171 1043 1203 1077
rect 1203 1043 1205 1077
rect 1099 969 1101 1003
rect 1101 969 1133 1003
rect 1171 969 1203 1003
rect 1203 969 1205 1003
rect 1099 895 1101 929
rect 1101 895 1133 929
rect 1171 895 1203 929
rect 1203 895 1205 929
rect 1099 821 1101 855
rect 1101 821 1133 855
rect 1171 821 1203 855
rect 1203 821 1205 855
rect 1099 747 1101 781
rect 1101 747 1133 781
rect 1171 747 1203 781
rect 1203 747 1205 781
rect 1099 673 1101 707
rect 1101 673 1133 707
rect 1171 673 1203 707
rect 1203 673 1205 707
rect 1099 599 1101 633
rect 1101 599 1133 633
rect 1171 599 1203 633
rect 1203 599 1205 633
rect 1099 525 1101 559
rect 1101 525 1133 559
rect 1171 525 1203 559
rect 1203 525 1205 559
rect 1099 451 1101 485
rect 1101 451 1133 485
rect 1171 451 1203 485
rect 1203 451 1205 485
rect 1099 377 1101 411
rect 1101 377 1133 411
rect 1171 377 1203 411
rect 1203 377 1205 411
rect 1099 303 1101 337
rect 1101 303 1133 337
rect 1171 303 1203 337
rect 1203 303 1205 337
rect 1099 229 1101 263
rect 1101 229 1133 263
rect 1171 229 1203 263
rect 1203 229 1205 263
rect 1099 155 1101 189
rect 1101 155 1133 189
rect 1171 155 1203 189
rect 1203 155 1205 189
<< metal1 >>
tri -14 1957 -2 1969 se
rect -2 1957 456 1969
tri 456 1957 468 1969 sw
tri 976 1957 988 1969 se
rect 988 1957 1274 1969
tri -48 1923 -14 1957 se
rect -14 1923 174 1957
rect 208 1923 246 1957
rect 280 1923 468 1957
tri 468 1923 502 1957 sw
tri 942 1923 976 1957 se
rect 976 1923 1099 1957
rect 1133 1923 1171 1957
rect 1205 1923 1274 1957
tri -49 1922 -48 1923 se
rect -48 1922 502 1923
tri 502 1922 503 1923 sw
rect -49 1884 503 1922
tri 903 1884 942 1923 se
rect 942 1884 1274 1923
rect -49 1850 174 1884
rect 208 1850 246 1884
rect 280 1850 503 1884
tri 883 1864 903 1884 se
rect 903 1864 1099 1884
rect -49 1811 503 1850
rect -49 1777 174 1811
rect 208 1777 246 1811
rect 280 1777 503 1811
rect -49 1738 503 1777
rect -49 1704 174 1738
rect 208 1704 246 1738
rect 280 1704 503 1738
rect -49 1665 503 1704
rect -49 1631 174 1665
rect 208 1631 246 1665
rect 280 1631 503 1665
rect -49 1592 503 1631
rect -49 1558 174 1592
rect 208 1558 246 1592
rect 280 1558 503 1592
rect -49 1519 503 1558
rect -49 1485 174 1519
rect 208 1485 246 1519
rect 280 1485 503 1519
rect -49 1446 503 1485
rect -49 1412 174 1446
rect 208 1412 246 1446
rect 280 1412 503 1446
rect -49 1373 503 1412
rect -49 1339 174 1373
rect 208 1339 246 1373
rect 280 1339 503 1373
rect -49 1299 503 1339
rect -49 1265 174 1299
rect 208 1265 246 1299
rect 280 1265 503 1299
rect -49 1225 503 1265
rect -49 1191 174 1225
rect 208 1191 246 1225
rect 280 1191 503 1225
rect -49 1151 503 1191
rect -49 1117 174 1151
rect 208 1117 246 1151
rect 280 1117 503 1151
rect -49 1077 503 1117
rect -49 1043 174 1077
rect 208 1043 246 1077
rect 280 1043 503 1077
rect -49 1003 503 1043
rect -49 969 174 1003
rect 208 969 246 1003
rect 280 969 503 1003
rect -49 929 503 969
rect -49 895 174 929
rect 208 895 246 929
rect 280 895 503 929
rect -49 855 503 895
rect -49 821 174 855
rect 208 821 246 855
rect 280 821 503 855
rect -49 781 503 821
rect -49 747 174 781
rect 208 747 246 781
rect 280 747 503 781
rect -49 707 503 747
rect -49 673 174 707
rect 208 673 246 707
rect 280 673 503 707
rect -49 633 503 673
rect -49 599 174 633
rect 208 599 246 633
rect 280 599 503 633
rect -49 559 503 599
rect -49 525 174 559
rect 208 525 246 559
rect 280 525 503 559
rect -49 485 503 525
rect -49 451 174 485
rect 208 451 246 485
rect 280 451 503 485
rect -49 411 503 451
rect -49 377 174 411
rect 208 377 246 411
rect 280 377 503 411
rect -49 337 503 377
rect -49 303 174 337
rect 208 303 246 337
rect 280 303 503 337
rect -49 263 503 303
rect -49 229 174 263
rect 208 229 246 263
rect 280 229 503 263
rect -49 228 503 229
rect -49 190 465 228
tri 465 190 503 228 nw
tri 876 1857 883 1864 se
rect 883 1857 1099 1864
rect 876 1850 1099 1857
rect 1133 1850 1171 1884
rect 1205 1864 1274 1884
tri 1274 1864 1379 1969 sw
rect 1205 1850 1381 1864
rect 876 1815 1381 1850
tri 1381 1815 1428 1862 sw
rect 876 1811 1428 1815
rect 876 1777 1099 1811
rect 1133 1777 1171 1811
rect 1205 1777 1428 1811
rect 876 1738 1428 1777
rect 876 1704 1099 1738
rect 1133 1704 1171 1738
rect 1205 1704 1428 1738
rect 876 1665 1428 1704
rect 876 1631 1099 1665
rect 1133 1631 1171 1665
rect 1205 1631 1428 1665
rect 876 1592 1428 1631
rect 876 1558 1099 1592
rect 1133 1558 1171 1592
rect 1205 1558 1428 1592
rect 876 1519 1428 1558
rect 876 1485 1099 1519
rect 1133 1485 1171 1519
rect 1205 1485 1428 1519
rect 876 1446 1428 1485
rect 876 1412 1099 1446
rect 1133 1412 1171 1446
rect 1205 1412 1428 1446
rect 876 1373 1428 1412
rect 876 1339 1099 1373
rect 1133 1339 1171 1373
rect 1205 1339 1428 1373
rect 876 1299 1428 1339
rect 876 1265 1099 1299
rect 1133 1265 1171 1299
rect 1205 1265 1428 1299
rect 876 1225 1428 1265
rect 876 1191 1099 1225
rect 1133 1191 1171 1225
rect 1205 1191 1428 1225
rect 876 1151 1428 1191
rect 876 1117 1099 1151
rect 1133 1117 1171 1151
rect 1205 1117 1428 1151
rect 876 1077 1428 1117
rect 876 1043 1099 1077
rect 1133 1043 1171 1077
rect 1205 1043 1428 1077
rect 876 1003 1428 1043
rect 876 969 1099 1003
rect 1133 969 1171 1003
rect 1205 969 1428 1003
rect 876 929 1428 969
rect 876 895 1099 929
rect 1133 895 1171 929
rect 1205 895 1428 929
rect 876 855 1428 895
rect 876 821 1099 855
rect 1133 821 1171 855
rect 1205 821 1428 855
rect 876 781 1428 821
rect 876 747 1099 781
rect 1133 747 1171 781
rect 1205 747 1428 781
rect 876 707 1428 747
rect 876 673 1099 707
rect 1133 673 1171 707
rect 1205 673 1428 707
rect 876 633 1428 673
rect 876 599 1099 633
rect 1133 599 1171 633
rect 1205 599 1428 633
rect 876 559 1428 599
rect 876 525 1099 559
rect 1133 525 1171 559
rect 1205 525 1428 559
rect 876 485 1428 525
rect 876 451 1099 485
rect 1133 451 1171 485
rect 1205 451 1428 485
rect 876 411 1428 451
rect 876 377 1099 411
rect 1133 377 1171 411
rect 1205 377 1428 411
rect 876 337 1428 377
rect 876 303 1099 337
rect 1133 303 1171 337
rect 1205 303 1428 337
rect 876 263 1428 303
rect 876 229 1099 263
rect 1133 229 1171 263
rect 1205 257 1428 263
rect 1205 233 1404 257
tri 1404 233 1428 257 nw
rect 1205 229 1314 233
rect 876 190 1314 229
tri -49 189 -48 190 ne
rect -48 189 464 190
tri 464 189 465 190 nw
tri 876 189 877 190 ne
rect 877 189 1314 190
tri -48 155 -14 189 ne
rect -14 155 174 189
rect 208 155 246 189
rect 280 155 430 189
tri 430 155 464 189 nw
tri 877 155 911 189 ne
rect 911 155 1099 189
rect 1133 155 1171 189
rect 1205 155 1314 189
tri -14 143 -2 155 ne
rect -2 143 418 155
tri 418 143 430 155 nw
tri 911 143 923 155 ne
rect 923 143 1314 155
tri 1314 143 1404 233 nw
<< labels >>
flabel poly s 778 -82 1038 5 0 FreeSans 48 0 0 0 g
port 2 nsew
flabel poly s 778 2107 1038 2199 0 FreeSans 48 0 0 0 g
port 2 nsew
<< properties >>
string GDS_END 94881792
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 94866986
string path 28.800 2.925 28.800 49.875 
<< end >>
