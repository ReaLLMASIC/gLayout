magic
tech sky130B
timestamp 1701704242
<< poly >>
rect 0 25 339 33
rect 0 8 8 25
rect 25 8 42 25
rect 59 8 76 25
rect 93 8 110 25
rect 127 8 144 25
rect 161 8 178 25
rect 195 8 212 25
rect 229 8 246 25
rect 263 8 280 25
rect 297 8 314 25
rect 331 8 339 25
rect 0 0 339 8
<< polycont >>
rect 8 8 25 25
rect 42 8 59 25
rect 76 8 93 25
rect 110 8 127 25
rect 144 8 161 25
rect 178 8 195 25
rect 212 8 229 25
rect 246 8 263 25
rect 280 8 297 25
rect 314 8 331 25
<< locali >>
rect 8 25 331 33
rect 25 8 42 25
rect 59 8 76 25
rect 93 8 110 25
rect 127 8 144 25
rect 161 8 178 25
rect 195 8 212 25
rect 229 8 246 25
rect 263 8 280 25
rect 297 8 314 25
rect 8 0 331 8
<< properties >>
string GDS_END 85363028
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85362192
<< end >>
