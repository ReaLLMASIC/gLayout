magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< nwell >>
rect 81 1874 2606 1910
rect 81 1142 217 1874
rect 1640 1142 2606 1248
rect 81 1112 2606 1142
<< pwell >>
rect 57 0 143 1052
rect 993 0 1079 1052
<< mvpsubdiff >>
rect 83 1002 117 1026
rect 83 931 117 968
rect 83 860 117 897
rect 83 789 117 826
rect 83 718 117 755
rect 83 647 117 684
rect 83 576 117 613
rect 83 505 117 542
rect 83 434 117 471
rect 83 364 117 400
rect 83 294 117 330
rect 83 224 117 260
rect 83 154 117 190
rect 83 84 117 120
rect 83 26 117 50
rect 1019 1002 1053 1026
rect 1019 931 1053 968
rect 1019 860 1053 897
rect 1019 789 1053 826
rect 1019 718 1053 755
rect 1019 647 1053 684
rect 1019 576 1053 613
rect 1019 505 1053 542
rect 1019 434 1053 471
rect 1019 364 1053 400
rect 1019 294 1053 330
rect 1019 224 1053 260
rect 1019 154 1053 190
rect 1019 84 1053 120
rect 1019 26 1053 50
<< mvnsubdiff >>
rect 147 1814 181 1838
rect 147 1741 181 1780
rect 147 1668 181 1707
rect 147 1596 181 1634
rect 147 1524 181 1562
rect 147 1452 181 1490
rect 147 1380 181 1418
rect 147 1308 181 1346
rect 147 1236 181 1274
rect 147 1178 181 1202
<< mvpsubdiffcont >>
rect 83 968 117 1002
rect 83 897 117 931
rect 83 826 117 860
rect 83 755 117 789
rect 83 684 117 718
rect 83 613 117 647
rect 83 542 117 576
rect 83 471 117 505
rect 83 400 117 434
rect 83 330 117 364
rect 83 260 117 294
rect 83 190 117 224
rect 83 120 117 154
rect 83 50 117 84
rect 1019 968 1053 1002
rect 1019 897 1053 931
rect 1019 826 1053 860
rect 1019 755 1053 789
rect 1019 684 1053 718
rect 1019 613 1053 647
rect 1019 542 1053 576
rect 1019 471 1053 505
rect 1019 400 1053 434
rect 1019 330 1053 364
rect 1019 260 1053 294
rect 1019 190 1053 224
rect 1019 120 1053 154
rect 1019 50 1053 84
<< mvnsubdiffcont >>
rect 147 1780 181 1814
rect 147 1707 181 1741
rect 147 1634 181 1668
rect 147 1562 181 1596
rect 147 1490 181 1524
rect 147 1418 181 1452
rect 147 1346 181 1380
rect 147 1274 181 1308
rect 147 1202 181 1236
<< poly >>
rect 331 1834 899 1906
rect 1063 1890 1265 1906
rect 1063 1856 1079 1890
rect 1113 1856 1147 1890
rect 1181 1856 1215 1890
rect 1249 1856 1265 1890
rect 1063 1834 1265 1856
rect 1321 1890 1523 1906
rect 1321 1856 1337 1890
rect 1371 1856 1405 1890
rect 1439 1856 1473 1890
rect 1507 1856 1523 1890
rect 1321 1834 1523 1856
rect 1687 1834 2487 1906
rect 1687 1216 2487 1288
rect 244 1108 730 1182
rect 244 1074 392 1108
rect 426 1074 460 1108
rect 494 1074 528 1108
rect 562 1074 596 1108
rect 630 1074 664 1108
rect 698 1074 730 1108
rect 244 1052 730 1074
rect 772 1108 906 1124
rect 772 1074 788 1108
rect 822 1074 856 1108
rect 890 1074 906 1108
rect 772 1052 906 1074
<< polycont >>
rect 1079 1856 1113 1890
rect 1147 1856 1181 1890
rect 1215 1856 1249 1890
rect 1337 1856 1371 1890
rect 1405 1856 1439 1890
rect 1473 1856 1507 1890
rect 392 1074 426 1108
rect 460 1074 494 1108
rect 528 1074 562 1108
rect 596 1074 630 1108
rect 664 1074 698 1108
rect 788 1074 822 1108
rect 856 1074 890 1108
<< locali >>
rect 147 1814 181 1838
rect 345 1825 888 1890
rect 1063 1856 1079 1890
rect 1113 1856 1147 1890
rect 1181 1856 1215 1890
rect 1249 1856 1265 1890
rect 1321 1856 1337 1890
rect 1371 1856 1405 1890
rect 1439 1856 1473 1890
rect 1507 1856 1523 1890
rect 1710 1825 2456 1890
rect 147 1741 181 1780
rect 147 1668 181 1707
rect 147 1596 181 1634
rect 147 1524 181 1562
rect 147 1452 181 1490
rect 147 1380 181 1418
rect 147 1308 181 1346
rect 147 1253 181 1274
rect 147 1181 181 1202
rect 147 1109 181 1147
rect 278 1555 336 1746
rect 1642 1555 1828 1791
rect 278 1521 286 1555
rect 320 1521 358 1555
rect 597 1521 635 1555
rect 874 1521 912 1555
rect 1756 1521 1794 1555
rect 278 1144 336 1521
rect 2498 1512 2532 1610
rect 442 1441 480 1475
rect 1494 1441 1532 1475
rect 754 1367 792 1401
rect 1012 1367 1050 1401
rect 215 1086 336 1144
rect 1276 1253 1310 1270
rect 1276 1181 1310 1219
rect 1642 1253 1676 1310
rect 1719 1266 2464 1339
rect 1642 1181 1676 1219
rect 1276 1109 1310 1147
rect 83 1002 117 1026
rect 83 931 117 968
rect 83 860 117 897
rect 215 871 257 1086
rect 376 1074 392 1108
rect 426 1074 460 1108
rect 494 1074 528 1108
rect 562 1074 596 1108
rect 630 1074 664 1108
rect 698 1074 714 1108
rect 772 1074 788 1108
rect 822 1074 856 1108
rect 890 1074 906 1108
rect 443 1023 517 1074
rect 443 989 465 1023
rect 499 989 517 1023
rect 443 951 517 989
rect 443 917 465 951
rect 499 917 517 951
rect 443 905 517 917
rect 619 1023 693 1074
rect 619 989 633 1023
rect 667 989 693 1023
rect 619 951 693 989
rect 619 917 633 951
rect 667 917 693 951
rect 619 905 693 917
rect 795 1023 869 1074
rect 795 989 817 1023
rect 851 989 869 1023
rect 795 951 869 989
rect 795 917 817 951
rect 851 917 869 951
rect 795 905 869 917
rect 1019 1002 1053 1026
rect 1019 931 1053 968
rect 233 837 271 871
rect 547 837 585 871
rect 865 837 903 871
rect 1019 860 1053 897
rect 83 789 117 826
rect 83 718 117 755
rect 83 656 117 684
rect 83 584 117 613
rect 83 505 117 542
rect 83 434 117 471
rect 83 364 117 400
rect 83 294 117 330
rect 83 224 117 260
rect 83 154 117 190
rect 83 84 117 120
rect 83 26 117 50
rect 215 22 257 837
rect 1019 789 1053 826
rect 1019 718 1053 755
rect 1019 656 1053 684
rect 375 584 409 622
rect 727 584 761 622
rect 1019 584 1053 613
rect 1019 505 1053 542
rect 1019 434 1053 471
rect 1019 364 1053 400
rect 1019 294 1053 330
rect 1019 224 1053 260
rect 1019 154 1053 190
rect 1019 84 1053 120
rect 1019 26 1053 50
<< viali >>
rect 147 1236 181 1253
rect 147 1219 181 1236
rect 147 1147 181 1181
rect 286 1521 320 1555
rect 358 1521 392 1555
rect 563 1521 597 1555
rect 635 1521 669 1555
rect 840 1521 874 1555
rect 912 1521 946 1555
rect 1722 1521 1756 1555
rect 1794 1521 1828 1555
rect 408 1441 442 1475
rect 480 1441 514 1475
rect 1460 1441 1494 1475
rect 1532 1441 1566 1475
rect 720 1367 754 1401
rect 792 1367 826 1401
rect 978 1367 1012 1401
rect 1050 1367 1084 1401
rect 147 1075 181 1109
rect 1276 1219 1310 1253
rect 1276 1147 1310 1181
rect 1642 1219 1676 1253
rect 1642 1147 1676 1181
rect 1276 1075 1310 1109
rect 465 989 499 1023
rect 465 917 499 951
rect 633 989 667 1023
rect 633 917 667 951
rect 817 989 851 1023
rect 817 917 851 951
rect 199 837 233 871
rect 271 837 305 871
rect 513 837 547 871
rect 585 837 619 871
rect 831 837 865 871
rect 903 837 937 871
rect 83 647 117 656
rect 83 622 117 647
rect 83 576 117 584
rect 83 550 117 576
rect 375 622 409 656
rect 375 550 409 584
rect 727 622 761 656
rect 727 550 761 584
rect 1019 647 1053 656
rect 1019 622 1053 647
rect 1019 576 1053 584
rect 1019 550 1053 576
<< metal1 >>
rect -528 1819 -522 1871
rect -470 1819 -458 1871
rect -406 1819 2476 1871
rect 0 1589 2606 1791
rect 274 1555 1718 1561
rect 274 1521 286 1555
rect 320 1521 358 1555
rect 392 1521 563 1555
rect 597 1521 635 1555
rect 669 1521 840 1555
rect 874 1521 912 1555
rect 946 1521 1718 1555
rect 274 1509 1718 1521
rect 1770 1509 1782 1561
rect 1834 1509 1840 1561
rect 396 1475 1578 1481
rect 396 1441 408 1475
rect 442 1441 480 1475
rect 514 1441 1460 1475
rect 1494 1441 1532 1475
rect 1566 1441 1578 1475
rect 396 1435 1578 1441
rect 2187 1415 2239 1421
rect 708 1401 1096 1407
rect 708 1367 720 1401
rect 754 1367 792 1401
rect 826 1367 978 1401
rect 1012 1367 1050 1401
rect 1084 1367 1096 1401
rect 708 1361 1096 1367
tri 2184 1361 2187 1364 se
rect 2187 1361 2239 1363
tri 2162 1339 2184 1361 se
rect 2184 1351 2239 1361
rect 2184 1339 2187 1351
tri 2239 1339 2264 1364 sw
rect 2187 1293 2239 1299
rect 0 1253 2606 1265
rect 0 1219 147 1253
rect 181 1219 1276 1253
rect 1310 1219 1642 1253
rect 1676 1219 2606 1253
rect 0 1181 2606 1219
rect 0 1147 147 1181
rect 181 1147 1276 1181
rect 1310 1147 1642 1181
rect 1676 1147 2606 1181
rect 0 1109 2606 1147
rect 0 1075 147 1109
rect 181 1075 1276 1109
rect 1310 1075 2606 1109
rect 0 1063 2606 1075
rect -528 919 -522 1035
rect -406 1023 673 1035
rect -406 989 465 1023
rect 499 989 633 1023
rect 667 989 673 1023
rect -406 951 673 989
rect -406 919 465 951
rect -528 917 465 919
rect 499 917 633 951
rect 667 917 673 951
rect -528 905 673 917
rect 811 1027 2239 1035
rect 811 1023 2187 1027
rect 811 989 817 1023
rect 851 989 2187 1023
rect 811 975 2187 989
rect 811 963 2239 975
rect 811 951 2187 963
rect 811 917 817 951
rect 851 917 2187 951
rect 811 911 2187 917
rect 811 905 2239 911
rect 187 871 1718 877
rect 187 837 199 871
rect 233 837 271 871
rect 305 837 513 871
rect 547 837 585 871
rect 619 837 831 871
rect 865 837 903 871
rect 937 837 1718 871
rect 187 825 1718 837
rect 1770 825 1782 877
rect 1834 825 1840 877
rect 0 656 2606 668
rect 0 622 83 656
rect 117 622 375 656
rect 409 622 727 656
rect 761 622 1019 656
rect 1053 622 2606 656
rect 0 584 2606 622
rect 0 550 83 584
rect 117 550 375 584
rect 409 550 727 584
rect 761 550 1019 584
rect 1053 550 2606 584
rect 0 538 2606 550
<< via1 >>
rect -522 1819 -470 1871
rect -458 1819 -406 1871
rect 1718 1555 1770 1561
rect 1718 1521 1722 1555
rect 1722 1521 1756 1555
rect 1756 1521 1770 1555
rect 1718 1509 1770 1521
rect 1782 1555 1834 1561
rect 1782 1521 1794 1555
rect 1794 1521 1828 1555
rect 1828 1521 1834 1555
rect 1782 1509 1834 1521
rect 2187 1363 2239 1415
rect 2187 1299 2239 1351
rect -522 919 -406 1035
rect 2187 975 2239 1027
rect 2187 911 2239 963
rect 1718 825 1770 877
rect 1782 825 1834 877
<< metal2 >>
rect -528 1819 -522 1871
rect -470 1819 -458 1871
rect -406 1819 -400 1871
rect -528 1035 -400 1819
rect -528 919 -522 1035
rect -406 919 -400 1035
rect 1712 1509 1718 1561
rect 1770 1509 1782 1561
rect 1834 1509 1840 1561
rect 1712 877 1840 1509
rect 2187 1415 2239 1421
rect 2187 1351 2239 1363
rect 2187 1027 2239 1299
rect 2187 963 2239 975
rect 2187 905 2239 911
rect 1712 825 1718 877
rect 1770 825 1782 877
rect 1834 825 1840 877
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1701704242
transform 0 1 727 -1 0 656
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1701704242
transform 0 1 375 -1 0 656
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1701704242
transform 0 1 83 -1 0 656
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_3
timestamp 1701704242
transform 0 1 1019 -1 0 656
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_4
timestamp 1701704242
transform -1 0 305 0 1 837
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_5
timestamp 1701704242
transform -1 0 619 0 1 837
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_6
timestamp 1701704242
transform -1 0 937 0 1 837
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_7
timestamp 1701704242
transform -1 0 1084 0 1 1367
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_8
timestamp 1701704242
transform -1 0 826 0 1 1367
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_9
timestamp 1701704242
transform -1 0 1566 0 1 1441
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_10
timestamp 1701704242
transform -1 0 514 0 1 1441
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_11
timestamp 1701704242
transform 0 -1 1676 1 0 1147
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_12
timestamp 1701704242
transform 0 -1 667 1 0 917
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_13
timestamp 1701704242
transform 0 -1 499 1 0 917
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_14
timestamp 1701704242
transform 0 -1 851 1 0 917
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_15
timestamp 1701704242
transform 1 0 286 0 1 1521
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_16
timestamp 1701704242
transform 1 0 563 0 1 1521
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_17
timestamp 1701704242
transform 1 0 1722 0 1 1521
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_18
timestamp 1701704242
transform 1 0 840 0 1 1521
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_0
timestamp 1701704242
transform 0 -1 181 -1 0 1253
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_1
timestamp 1701704242
transform 0 -1 1310 -1 0 1253
box 0 0 1 1
use L1M1_CDNS_52468879185194  L1M1_CDNS_52468879185194_0
timestamp 1701704242
transform -1 0 2464 0 1 1825
box -12 -6 766 40
use L1M1_CDNS_52468879185195  L1M1_CDNS_52468879185195_0
timestamp 1701704242
transform 1 0 346 0 1 1825
box -12 -6 550 40
use L1M1_CDNS_52468879185326  L1M1_CDNS_52468879185326_0
timestamp 1701704242
transform 1 0 1743 0 1 1299
box -12 -6 694 40
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_0
timestamp 1701704242
transform -1 0 1840 0 -1 1561
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_1
timestamp 1701704242
transform 0 -1 2239 1 0 905
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_2
timestamp 1701704242
transform 0 -1 2239 1 0 1293
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_3
timestamp 1701704242
transform 1 0 1712 0 1 825
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_4
timestamp 1701704242
transform 1 0 -528 0 1 1819
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_0
timestamp 1701704242
transform 1 0 -528 0 -1 1035
box 0 0 1 1
use nfet_CDNS_52468879185343  nfet_CDNS_52468879185343_0
timestamp 1701704242
transform 1 0 772 0 1 26
box -79 -26 199 1026
use nfet_CDNS_524688791851403  nfet_CDNS_524688791851403_0
timestamp 1701704242
transform -1 0 716 0 1 26
box -79 -26 551 1026
use pfet_CDNS_52468879185323  pfet_CDNS_52468879185323_0
timestamp 1701704242
transform -1 0 1265 0 -1 1808
box -119 -66 319 666
use pfet_CDNS_52468879185323  pfet_CDNS_52468879185323_1
timestamp 1701704242
transform 1 0 1321 0 -1 1808
box -119 -66 319 666
use pfet_CDNS_52468879185324  pfet_CDNS_52468879185324_0
timestamp 1701704242
transform -1 0 587 0 1 1208
box -119 -66 375 666
use pfet_CDNS_52468879185324  pfet_CDNS_52468879185324_1
timestamp 1701704242
transform 1 0 643 0 1 1208
box -119 -66 375 666
use pfet_CDNS_52468879185329  pfet_CDNS_52468879185329_0
timestamp 1701704242
transform -1 0 2487 0 -1 1808
box -119 -66 919 266
use pfet_CDNS_52468879185329  pfet_CDNS_52468879185329_1
timestamp 1701704242
transform 1 0 1687 0 1 1314
box -119 -66 919 266
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_0
timestamp 1701704242
transform 0 1 772 -1 0 1124
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_0
timestamp 1701704242
transform 0 -1 1523 -1 0 1906
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_1
timestamp 1701704242
transform 0 1 1063 -1 0 1906
box 0 0 1 1
use PYL1_CDNS_52468879185289  PYL1_CDNS_52468879185289_0
timestamp 1701704242
transform 0 -1 714 -1 0 1124
box 0 0 1 1
use PYL1_CDNS_52468879185317  PYL1_CDNS_52468879185317_0
timestamp 1701704242
transform 0 -1 2465 -1 0 1282
box 0 0 66 746
use PYL1_CDNS_52468879185317  PYL1_CDNS_52468879185317_1
timestamp 1701704242
transform 0 -1 2448 1 0 1840
box 0 0 66 746
use PYL1_CDNS_52468879185318  PYL1_CDNS_52468879185318_0
timestamp 1701704242
transform 0 -1 888 -1 0 1906
box 0 0 66 542
<< labels >>
flabel comment s 882 1122 882 1122 0 FreeSans 300 0 0 0 pden_h_n
flabel comment s 2512 1553 2512 1553 0 FreeSans 300 90 0 0 int_slow
flabel comment s 1146 1890 1146 1890 0 FreeSans 300 0 0 0 en_fast_n<0>
flabel comment s 1523 1886 1523 1886 0 FreeSans 300 0 0 0 en_fast_n<1>
flabel comment s 2071 1905 2071 1905 0 FreeSans 300 0 0 0 drvlo_h_n
flabel comment s 315 861 315 861 0 FreeSans 300 0 0 0 pd_h
flabel comment s 562 1547 562 1547 0 FreeSans 300 0 0 0 pd_h
flabel comment s 1162 1465 1162 1465 0 FreeSans 300 0 0 0 intnr1
flabel comment s 993 1395 993 1395 0 FreeSans 300 0 0 0 intnr0
flabel comment s 2114 1228 2114 1228 0 FreeSans 300 0 0 0 pden_h_n
flabel metal1 s 2566 1063 2606 1265 7 FreeSans 300 180 0 0 vcc_io
port 2 nsew
flabel metal1 s 0 1063 40 1265 3 FreeSans 300 180 0 0 vcc_io
port 2 nsew
flabel metal1 s 0 538 42 668 3 FreeSans 300 180 0 0 vgnd_io
port 1 nsew
flabel metal1 s 2564 538 2606 668 7 FreeSans 300 180 0 0 vgnd_io
port 1 nsew
flabel metal1 s -528 1819 -481 1871 3 FreeSans 300 180 0 0 drvlo_h_n
port 3 nsew
flabel metal1 s 1793 825 1840 877 7 FreeSans 300 180 0 0 pd_h
port 4 nsew
flabel metal1 s 2187 905 2239 954 7 FreeSans 300 180 0 0 pden_h_n
port 5 nsew
flabel metal1 s 0 1589 42 1791 3 FreeSans 300 180 0 0 vgnd_io
port 1 nsew
flabel metal1 s 2564 1589 2606 1791 7 FreeSans 300 180 0 0 vgnd_io
port 1 nsew
flabel locali s 1477 1856 1523 1890 0 FreeSans 300 180 0 0 en_fast_n<1>
port 7 nsew
flabel locali s 1101 1856 1147 1890 0 FreeSans 300 180 0 0 en_fast_n<0>
port 8 nsew
<< properties >>
string GDS_END 87858102
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 87847588
string path 4.100 46.600 4.100 28.800 
<< end >>
