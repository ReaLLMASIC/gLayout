magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -38 261 1418 582
<< pwell >>
rect 1 21 1303 203
rect 30 -17 64 21
<< scnmos >>
rect 83 47 113 177
rect 167 47 197 177
rect 251 47 281 177
rect 335 47 365 177
rect 419 47 449 177
rect 607 47 637 177
rect 691 47 721 177
rect 775 47 805 177
rect 859 47 889 177
rect 943 47 973 177
rect 1027 47 1057 177
rect 1111 47 1141 177
rect 1195 47 1225 177
<< scpmoshvt >>
rect 83 297 113 497
rect 167 297 197 497
rect 251 297 281 497
rect 335 297 365 497
rect 419 297 449 497
rect 607 297 637 497
rect 691 297 721 497
rect 775 297 805 497
rect 859 297 889 497
rect 943 297 973 497
rect 1027 297 1057 497
rect 1111 297 1141 497
rect 1195 297 1225 497
<< ndiff >>
rect 27 163 83 177
rect 27 129 39 163
rect 73 129 83 163
rect 27 95 83 129
rect 27 61 39 95
rect 73 61 83 95
rect 27 47 83 61
rect 113 95 167 177
rect 113 61 123 95
rect 157 61 167 95
rect 113 47 167 61
rect 197 163 251 177
rect 197 129 207 163
rect 241 129 251 163
rect 197 95 251 129
rect 197 61 207 95
rect 241 61 251 95
rect 197 47 251 61
rect 281 95 335 177
rect 281 61 291 95
rect 325 61 335 95
rect 281 47 335 61
rect 365 163 419 177
rect 365 129 375 163
rect 409 129 419 163
rect 365 95 419 129
rect 365 61 375 95
rect 409 61 419 95
rect 365 47 419 61
rect 449 95 607 177
rect 449 61 459 95
rect 493 61 563 95
rect 597 61 607 95
rect 449 47 607 61
rect 637 163 691 177
rect 637 129 647 163
rect 681 129 691 163
rect 637 95 691 129
rect 637 61 647 95
rect 681 61 691 95
rect 637 47 691 61
rect 721 95 775 177
rect 721 61 731 95
rect 765 61 775 95
rect 721 47 775 61
rect 805 163 859 177
rect 805 129 815 163
rect 849 129 859 163
rect 805 95 859 129
rect 805 61 815 95
rect 849 61 859 95
rect 805 47 859 61
rect 889 95 943 177
rect 889 61 899 95
rect 933 61 943 95
rect 889 47 943 61
rect 973 163 1027 177
rect 973 129 983 163
rect 1017 129 1027 163
rect 973 95 1027 129
rect 973 61 983 95
rect 1017 61 1027 95
rect 973 47 1027 61
rect 1057 95 1111 177
rect 1057 61 1067 95
rect 1101 61 1111 95
rect 1057 47 1111 61
rect 1141 163 1195 177
rect 1141 129 1151 163
rect 1185 129 1195 163
rect 1141 95 1195 129
rect 1141 61 1151 95
rect 1185 61 1195 95
rect 1141 47 1195 61
rect 1225 95 1277 177
rect 1225 61 1235 95
rect 1269 61 1277 95
rect 1225 47 1277 61
<< pdiff >>
rect 27 477 83 497
rect 27 443 39 477
rect 73 443 83 477
rect 27 409 83 443
rect 27 375 39 409
rect 73 375 83 409
rect 27 341 83 375
rect 27 307 39 341
rect 73 307 83 341
rect 27 297 83 307
rect 113 477 167 497
rect 113 443 123 477
rect 157 443 167 477
rect 113 409 167 443
rect 113 375 123 409
rect 157 375 167 409
rect 113 297 167 375
rect 197 477 251 497
rect 197 443 207 477
rect 241 443 251 477
rect 197 409 251 443
rect 197 375 207 409
rect 241 375 251 409
rect 197 297 251 375
rect 281 477 335 497
rect 281 443 291 477
rect 325 443 335 477
rect 281 297 335 443
rect 365 477 419 497
rect 365 443 375 477
rect 409 443 419 477
rect 365 409 419 443
rect 365 375 375 409
rect 409 375 419 409
rect 365 297 419 375
rect 449 477 501 497
rect 449 443 459 477
rect 493 443 501 477
rect 449 297 501 443
rect 555 477 607 497
rect 555 443 563 477
rect 597 443 607 477
rect 555 297 607 443
rect 637 409 691 497
rect 637 375 647 409
rect 681 375 691 409
rect 637 297 691 375
rect 721 477 775 497
rect 721 443 731 477
rect 765 443 775 477
rect 721 297 775 443
rect 805 409 859 497
rect 805 375 815 409
rect 849 375 859 409
rect 805 297 859 375
rect 889 477 943 497
rect 889 443 899 477
rect 933 443 943 477
rect 889 409 943 443
rect 889 375 899 409
rect 933 375 943 409
rect 889 297 943 375
rect 973 409 1027 497
rect 973 375 983 409
rect 1017 375 1027 409
rect 973 341 1027 375
rect 973 307 983 341
rect 1017 307 1027 341
rect 973 297 1027 307
rect 1057 477 1111 497
rect 1057 443 1067 477
rect 1101 443 1111 477
rect 1057 409 1111 443
rect 1057 375 1067 409
rect 1101 375 1111 409
rect 1057 297 1111 375
rect 1141 409 1195 497
rect 1141 375 1151 409
rect 1185 375 1195 409
rect 1141 341 1195 375
rect 1141 307 1151 341
rect 1185 307 1195 341
rect 1141 297 1195 307
rect 1225 477 1277 497
rect 1225 443 1235 477
rect 1269 443 1277 477
rect 1225 409 1277 443
rect 1225 375 1235 409
rect 1269 375 1277 409
rect 1225 297 1277 375
<< ndiffc >>
rect 39 129 73 163
rect 39 61 73 95
rect 123 61 157 95
rect 207 129 241 163
rect 207 61 241 95
rect 291 61 325 95
rect 375 129 409 163
rect 375 61 409 95
rect 459 61 493 95
rect 563 61 597 95
rect 647 129 681 163
rect 647 61 681 95
rect 731 61 765 95
rect 815 129 849 163
rect 815 61 849 95
rect 899 61 933 95
rect 983 129 1017 163
rect 983 61 1017 95
rect 1067 61 1101 95
rect 1151 129 1185 163
rect 1151 61 1185 95
rect 1235 61 1269 95
<< pdiffc >>
rect 39 443 73 477
rect 39 375 73 409
rect 39 307 73 341
rect 123 443 157 477
rect 123 375 157 409
rect 207 443 241 477
rect 207 375 241 409
rect 291 443 325 477
rect 375 443 409 477
rect 375 375 409 409
rect 459 443 493 477
rect 563 443 597 477
rect 647 375 681 409
rect 731 443 765 477
rect 815 375 849 409
rect 899 443 933 477
rect 899 375 933 409
rect 983 375 1017 409
rect 983 307 1017 341
rect 1067 443 1101 477
rect 1067 375 1101 409
rect 1151 375 1185 409
rect 1151 307 1185 341
rect 1235 443 1269 477
rect 1235 375 1269 409
<< poly >>
rect 83 497 113 523
rect 167 497 197 523
rect 251 497 281 523
rect 335 497 365 523
rect 419 497 449 523
rect 607 497 637 523
rect 691 497 721 523
rect 775 497 805 523
rect 859 497 889 523
rect 943 497 973 523
rect 1027 497 1057 523
rect 1111 497 1141 523
rect 1195 497 1225 523
rect 83 265 113 297
rect 22 249 113 265
rect 22 215 38 249
rect 72 215 113 249
rect 22 199 113 215
rect 83 177 113 199
rect 167 265 197 297
rect 251 265 281 297
rect 335 265 365 297
rect 419 265 449 297
rect 167 249 449 265
rect 167 215 251 249
rect 285 215 319 249
rect 353 215 387 249
rect 421 215 449 249
rect 167 199 449 215
rect 167 177 197 199
rect 251 177 281 199
rect 335 177 365 199
rect 419 177 449 199
rect 607 265 637 297
rect 691 265 721 297
rect 775 265 805 297
rect 859 265 889 297
rect 607 249 889 265
rect 607 215 623 249
rect 657 215 691 249
rect 725 215 759 249
rect 793 215 889 249
rect 607 199 889 215
rect 607 177 637 199
rect 691 177 721 199
rect 775 177 805 199
rect 859 177 889 199
rect 943 265 973 297
rect 1027 265 1057 297
rect 1111 265 1141 297
rect 1195 265 1225 297
rect 943 249 1225 265
rect 943 215 959 249
rect 993 215 1027 249
rect 1061 215 1095 249
rect 1129 215 1163 249
rect 1197 215 1225 249
rect 943 199 1225 215
rect 943 177 973 199
rect 1027 177 1057 199
rect 1111 177 1141 199
rect 1195 177 1225 199
rect 83 21 113 47
rect 167 21 197 47
rect 251 21 281 47
rect 335 21 365 47
rect 419 21 449 47
rect 607 21 637 47
rect 691 21 721 47
rect 775 21 805 47
rect 859 21 889 47
rect 943 21 973 47
rect 1027 21 1057 47
rect 1111 21 1141 47
rect 1195 21 1225 47
<< polycont >>
rect 38 215 72 249
rect 251 215 285 249
rect 319 215 353 249
rect 387 215 421 249
rect 623 215 657 249
rect 691 215 725 249
rect 759 215 793 249
rect 959 215 993 249
rect 1027 215 1061 249
rect 1095 215 1129 249
rect 1163 215 1197 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1380 561
rect 22 477 81 493
rect 22 443 39 477
rect 73 443 81 477
rect 22 409 81 443
rect 22 375 39 409
rect 73 375 81 409
rect 22 341 81 375
rect 115 477 165 527
rect 115 443 123 477
rect 157 443 165 477
rect 115 409 165 443
rect 115 375 123 409
rect 157 375 165 409
rect 115 359 165 375
rect 199 477 249 493
rect 199 443 207 477
rect 241 443 249 477
rect 199 409 249 443
rect 283 477 333 527
rect 283 443 291 477
rect 325 443 333 477
rect 283 427 333 443
rect 367 477 417 493
rect 367 443 375 477
rect 409 443 417 477
rect 199 375 207 409
rect 241 393 249 409
rect 367 409 417 443
rect 451 477 501 527
rect 451 443 459 477
rect 493 443 501 477
rect 451 427 501 443
rect 555 477 1277 493
rect 555 443 563 477
rect 597 459 731 477
rect 597 443 605 459
rect 555 427 605 443
rect 723 443 731 459
rect 765 459 899 477
rect 765 443 773 459
rect 723 427 773 443
rect 891 443 899 459
rect 933 459 1067 477
rect 933 443 941 459
rect 367 393 375 409
rect 241 375 375 393
rect 409 393 417 409
rect 639 409 689 425
rect 639 393 647 409
rect 409 375 647 393
rect 681 393 689 409
rect 807 409 857 425
rect 807 393 815 409
rect 681 375 815 393
rect 849 375 857 409
rect 199 359 857 375
rect 891 409 941 443
rect 1059 443 1067 459
rect 1101 459 1235 477
rect 1101 443 1109 459
rect 891 375 899 409
rect 933 375 941 409
rect 891 359 941 375
rect 975 409 1025 425
rect 975 375 983 409
rect 1017 375 1025 409
rect 22 307 39 341
rect 73 325 81 341
rect 975 341 1025 375
rect 1059 409 1109 443
rect 1227 443 1235 459
rect 1269 443 1277 477
rect 1059 375 1067 409
rect 1101 375 1109 409
rect 1059 359 1109 375
rect 1143 409 1193 425
rect 1143 375 1151 409
rect 1185 375 1193 409
rect 73 307 941 325
rect 22 291 941 307
rect 975 307 983 341
rect 1017 325 1025 341
rect 1143 341 1193 375
rect 1227 409 1277 443
rect 1227 375 1235 409
rect 1269 375 1277 409
rect 1227 359 1277 375
rect 1143 325 1151 341
rect 1017 307 1151 325
rect 1185 325 1193 341
rect 1311 325 1352 483
rect 1185 307 1352 325
rect 975 291 1352 307
rect 22 249 89 257
rect 22 215 38 249
rect 72 215 89 249
rect 123 181 157 291
rect 907 257 941 291
rect 207 249 538 257
rect 207 215 251 249
rect 285 215 319 249
rect 353 215 387 249
rect 421 215 538 249
rect 607 249 860 257
rect 607 215 623 249
rect 657 215 691 249
rect 725 215 759 249
rect 793 215 860 249
rect 907 249 1225 257
rect 907 215 959 249
rect 993 215 1027 249
rect 1061 215 1095 249
rect 1129 215 1163 249
rect 1197 215 1225 249
rect 1284 181 1352 291
rect 22 163 157 181
rect 22 129 39 163
rect 73 147 157 163
rect 191 163 1352 181
rect 73 129 89 147
rect 22 95 89 129
rect 191 129 207 163
rect 241 145 375 163
rect 241 129 257 145
rect 22 61 39 95
rect 73 61 89 95
rect 22 51 89 61
rect 123 95 157 111
rect 123 17 157 61
rect 191 95 257 129
rect 359 129 375 145
rect 409 145 647 163
rect 409 129 425 145
rect 191 61 207 95
rect 241 61 257 95
rect 191 51 257 61
rect 291 95 325 111
rect 291 17 325 61
rect 359 95 425 129
rect 631 129 647 145
rect 681 145 815 163
rect 681 129 697 145
rect 359 61 375 95
rect 409 61 425 95
rect 359 51 425 61
rect 459 95 597 111
rect 493 61 563 95
rect 459 17 597 61
rect 631 95 697 129
rect 799 129 815 145
rect 849 145 983 163
rect 849 129 865 145
rect 631 61 647 95
rect 681 61 697 95
rect 631 51 697 61
rect 731 95 765 111
rect 731 17 765 61
rect 799 95 865 129
rect 967 129 983 145
rect 1017 145 1151 163
rect 1017 129 1033 145
rect 799 61 815 95
rect 849 61 865 95
rect 799 51 865 61
rect 899 95 933 111
rect 899 17 933 61
rect 967 95 1033 129
rect 1135 129 1151 145
rect 1185 145 1352 163
rect 1185 129 1201 145
rect 967 61 983 95
rect 1017 61 1033 95
rect 967 51 1033 61
rect 1067 95 1101 111
rect 1067 17 1101 61
rect 1135 95 1201 129
rect 1135 61 1151 95
rect 1185 61 1201 95
rect 1135 51 1201 61
rect 1235 95 1269 111
rect 1303 63 1352 145
rect 1235 17 1269 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1380 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
<< metal1 >>
rect 0 561 1380 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1380 561
rect 0 496 1380 527
rect 0 17 1380 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1380 17
rect 0 -48 1380 -17
<< labels >>
flabel locali s 398 221 432 255 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 490 221 524 255 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 306 221 340 255 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 400 0 0 0 C_N
port 3 nsew signal input
flabel locali s 678 221 712 255 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel locali s 1317 357 1351 391 0 FreeSans 400 0 0 0 Y
port 8 nsew signal output
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 nor3b_4
rlabel metal1 s 0 -48 1380 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1380 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1380 544
string GDS_END 1123316
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1113216
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 6.900 0.000 
<< end >>
