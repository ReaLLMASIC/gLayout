magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -38 261 2430 582
<< pwell >>
rect 1 21 2391 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 267 47 297 177
rect 351 47 381 177
rect 435 47 465 177
rect 519 47 549 177
rect 603 47 633 177
rect 687 47 717 177
rect 771 47 801 177
rect 855 47 885 177
rect 939 47 969 177
rect 1023 47 1053 177
rect 1107 47 1137 177
rect 1191 47 1221 177
rect 1275 47 1305 177
rect 1359 47 1389 177
rect 1443 47 1473 177
rect 1527 47 1557 177
rect 1611 47 1641 177
rect 1695 47 1725 177
rect 1779 47 1809 177
rect 1863 47 1893 177
rect 1947 47 1977 177
rect 2031 47 2061 177
rect 2115 47 2145 177
rect 2199 47 2229 177
rect 2283 47 2313 177
<< scpmoshvt >>
rect 79 297 109 497
rect 267 297 297 497
rect 351 297 381 497
rect 435 297 465 497
rect 519 297 549 497
rect 603 297 633 497
rect 687 297 717 497
rect 771 297 801 497
rect 855 297 885 497
rect 939 297 969 497
rect 1023 297 1053 497
rect 1107 297 1137 497
rect 1191 297 1221 497
rect 1275 297 1305 497
rect 1359 297 1389 497
rect 1443 297 1473 497
rect 1527 297 1557 497
rect 1611 297 1641 497
rect 1695 297 1725 497
rect 1779 297 1809 497
rect 1863 297 1893 497
rect 1947 297 1977 497
rect 2031 297 2061 497
rect 2115 297 2145 497
rect 2199 297 2229 497
rect 2283 297 2313 497
<< ndiff >>
rect 27 165 79 177
rect 27 131 35 165
rect 69 131 79 165
rect 27 97 79 131
rect 27 63 35 97
rect 69 63 79 97
rect 27 47 79 63
rect 109 165 161 177
rect 109 131 119 165
rect 153 131 161 165
rect 109 97 161 131
rect 109 63 119 97
rect 153 63 161 97
rect 109 47 161 63
rect 215 165 267 177
rect 215 131 223 165
rect 257 131 267 165
rect 215 97 267 131
rect 215 63 223 97
rect 257 63 267 97
rect 215 47 267 63
rect 297 97 351 177
rect 297 63 307 97
rect 341 63 351 97
rect 297 47 351 63
rect 381 165 435 177
rect 381 131 391 165
rect 425 131 435 165
rect 381 97 435 131
rect 381 63 391 97
rect 425 63 435 97
rect 381 47 435 63
rect 465 97 519 177
rect 465 63 475 97
rect 509 63 519 97
rect 465 47 519 63
rect 549 165 603 177
rect 549 131 559 165
rect 593 131 603 165
rect 549 97 603 131
rect 549 63 559 97
rect 593 63 603 97
rect 549 47 603 63
rect 633 97 687 177
rect 633 63 643 97
rect 677 63 687 97
rect 633 47 687 63
rect 717 165 771 177
rect 717 131 727 165
rect 761 131 771 165
rect 717 97 771 131
rect 717 63 727 97
rect 761 63 771 97
rect 717 47 771 63
rect 801 97 855 177
rect 801 63 811 97
rect 845 63 855 97
rect 801 47 855 63
rect 885 165 939 177
rect 885 131 895 165
rect 929 131 939 165
rect 885 97 939 131
rect 885 63 895 97
rect 929 63 939 97
rect 885 47 939 63
rect 969 97 1023 177
rect 969 63 979 97
rect 1013 63 1023 97
rect 969 47 1023 63
rect 1053 165 1107 177
rect 1053 131 1063 165
rect 1097 131 1107 165
rect 1053 97 1107 131
rect 1053 63 1063 97
rect 1097 63 1107 97
rect 1053 47 1107 63
rect 1137 97 1191 177
rect 1137 63 1147 97
rect 1181 63 1191 97
rect 1137 47 1191 63
rect 1221 165 1275 177
rect 1221 131 1231 165
rect 1265 131 1275 165
rect 1221 97 1275 131
rect 1221 63 1231 97
rect 1265 63 1275 97
rect 1221 47 1275 63
rect 1305 97 1359 177
rect 1305 63 1315 97
rect 1349 63 1359 97
rect 1305 47 1359 63
rect 1389 165 1443 177
rect 1389 131 1399 165
rect 1433 131 1443 165
rect 1389 97 1443 131
rect 1389 63 1399 97
rect 1433 63 1443 97
rect 1389 47 1443 63
rect 1473 97 1527 177
rect 1473 63 1483 97
rect 1517 63 1527 97
rect 1473 47 1527 63
rect 1557 165 1611 177
rect 1557 131 1567 165
rect 1601 131 1611 165
rect 1557 97 1611 131
rect 1557 63 1567 97
rect 1601 63 1611 97
rect 1557 47 1611 63
rect 1641 97 1695 177
rect 1641 63 1651 97
rect 1685 63 1695 97
rect 1641 47 1695 63
rect 1725 165 1779 177
rect 1725 131 1735 165
rect 1769 131 1779 165
rect 1725 97 1779 131
rect 1725 63 1735 97
rect 1769 63 1779 97
rect 1725 47 1779 63
rect 1809 97 1863 177
rect 1809 63 1819 97
rect 1853 63 1863 97
rect 1809 47 1863 63
rect 1893 165 1947 177
rect 1893 131 1903 165
rect 1937 131 1947 165
rect 1893 97 1947 131
rect 1893 63 1903 97
rect 1937 63 1947 97
rect 1893 47 1947 63
rect 1977 97 2031 177
rect 1977 63 1987 97
rect 2021 63 2031 97
rect 1977 47 2031 63
rect 2061 165 2115 177
rect 2061 131 2071 165
rect 2105 131 2115 165
rect 2061 97 2115 131
rect 2061 63 2071 97
rect 2105 63 2115 97
rect 2061 47 2115 63
rect 2145 97 2199 177
rect 2145 63 2155 97
rect 2189 63 2199 97
rect 2145 47 2199 63
rect 2229 165 2283 177
rect 2229 131 2239 165
rect 2273 131 2283 165
rect 2229 97 2283 131
rect 2229 63 2239 97
rect 2273 63 2283 97
rect 2229 47 2283 63
rect 2313 97 2365 177
rect 2313 63 2323 97
rect 2357 63 2365 97
rect 2313 47 2365 63
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 417 79 451
rect 27 383 35 417
rect 69 383 79 417
rect 27 349 79 383
rect 27 315 35 349
rect 69 315 79 349
rect 27 297 79 315
rect 109 479 161 497
rect 109 445 119 479
rect 153 445 161 479
rect 109 411 161 445
rect 109 377 119 411
rect 153 377 161 411
rect 109 343 161 377
rect 109 309 119 343
rect 153 309 161 343
rect 109 297 161 309
rect 215 479 267 497
rect 215 445 223 479
rect 257 445 267 479
rect 215 411 267 445
rect 215 377 223 411
rect 257 377 267 411
rect 215 343 267 377
rect 215 309 223 343
rect 257 309 267 343
rect 215 297 267 309
rect 297 485 351 497
rect 297 451 307 485
rect 341 451 351 485
rect 297 417 351 451
rect 297 383 307 417
rect 341 383 351 417
rect 297 297 351 383
rect 381 479 435 497
rect 381 445 391 479
rect 425 445 435 479
rect 381 411 435 445
rect 381 377 391 411
rect 425 377 435 411
rect 381 343 435 377
rect 381 309 391 343
rect 425 309 435 343
rect 381 297 435 309
rect 465 485 519 497
rect 465 451 475 485
rect 509 451 519 485
rect 465 417 519 451
rect 465 383 475 417
rect 509 383 519 417
rect 465 297 519 383
rect 549 479 603 497
rect 549 445 559 479
rect 593 445 603 479
rect 549 411 603 445
rect 549 377 559 411
rect 593 377 603 411
rect 549 343 603 377
rect 549 309 559 343
rect 593 309 603 343
rect 549 297 603 309
rect 633 485 687 497
rect 633 451 643 485
rect 677 451 687 485
rect 633 417 687 451
rect 633 383 643 417
rect 677 383 687 417
rect 633 297 687 383
rect 717 479 771 497
rect 717 445 727 479
rect 761 445 771 479
rect 717 411 771 445
rect 717 377 727 411
rect 761 377 771 411
rect 717 343 771 377
rect 717 309 727 343
rect 761 309 771 343
rect 717 297 771 309
rect 801 485 855 497
rect 801 451 811 485
rect 845 451 855 485
rect 801 417 855 451
rect 801 383 811 417
rect 845 383 855 417
rect 801 297 855 383
rect 885 479 939 497
rect 885 445 895 479
rect 929 445 939 479
rect 885 411 939 445
rect 885 377 895 411
rect 929 377 939 411
rect 885 343 939 377
rect 885 309 895 343
rect 929 309 939 343
rect 885 297 939 309
rect 969 485 1023 497
rect 969 451 979 485
rect 1013 451 1023 485
rect 969 417 1023 451
rect 969 383 979 417
rect 1013 383 1023 417
rect 969 297 1023 383
rect 1053 479 1107 497
rect 1053 445 1063 479
rect 1097 445 1107 479
rect 1053 411 1107 445
rect 1053 377 1063 411
rect 1097 377 1107 411
rect 1053 343 1107 377
rect 1053 309 1063 343
rect 1097 309 1107 343
rect 1053 297 1107 309
rect 1137 485 1191 497
rect 1137 451 1147 485
rect 1181 451 1191 485
rect 1137 417 1191 451
rect 1137 383 1147 417
rect 1181 383 1191 417
rect 1137 297 1191 383
rect 1221 479 1275 497
rect 1221 445 1231 479
rect 1265 445 1275 479
rect 1221 411 1275 445
rect 1221 377 1231 411
rect 1265 377 1275 411
rect 1221 343 1275 377
rect 1221 309 1231 343
rect 1265 309 1275 343
rect 1221 297 1275 309
rect 1305 485 1359 497
rect 1305 451 1315 485
rect 1349 451 1359 485
rect 1305 417 1359 451
rect 1305 383 1315 417
rect 1349 383 1359 417
rect 1305 297 1359 383
rect 1389 479 1443 497
rect 1389 445 1399 479
rect 1433 445 1443 479
rect 1389 411 1443 445
rect 1389 377 1399 411
rect 1433 377 1443 411
rect 1389 343 1443 377
rect 1389 309 1399 343
rect 1433 309 1443 343
rect 1389 297 1443 309
rect 1473 485 1527 497
rect 1473 451 1483 485
rect 1517 451 1527 485
rect 1473 417 1527 451
rect 1473 383 1483 417
rect 1517 383 1527 417
rect 1473 297 1527 383
rect 1557 479 1611 497
rect 1557 445 1567 479
rect 1601 445 1611 479
rect 1557 411 1611 445
rect 1557 377 1567 411
rect 1601 377 1611 411
rect 1557 343 1611 377
rect 1557 309 1567 343
rect 1601 309 1611 343
rect 1557 297 1611 309
rect 1641 485 1695 497
rect 1641 451 1651 485
rect 1685 451 1695 485
rect 1641 417 1695 451
rect 1641 383 1651 417
rect 1685 383 1695 417
rect 1641 297 1695 383
rect 1725 479 1779 497
rect 1725 445 1735 479
rect 1769 445 1779 479
rect 1725 411 1779 445
rect 1725 377 1735 411
rect 1769 377 1779 411
rect 1725 343 1779 377
rect 1725 309 1735 343
rect 1769 309 1779 343
rect 1725 297 1779 309
rect 1809 485 1863 497
rect 1809 451 1819 485
rect 1853 451 1863 485
rect 1809 417 1863 451
rect 1809 383 1819 417
rect 1853 383 1863 417
rect 1809 297 1863 383
rect 1893 479 1947 497
rect 1893 445 1903 479
rect 1937 445 1947 479
rect 1893 411 1947 445
rect 1893 377 1903 411
rect 1937 377 1947 411
rect 1893 343 1947 377
rect 1893 309 1903 343
rect 1937 309 1947 343
rect 1893 297 1947 309
rect 1977 485 2031 497
rect 1977 451 1987 485
rect 2021 451 2031 485
rect 1977 417 2031 451
rect 1977 383 1987 417
rect 2021 383 2031 417
rect 1977 297 2031 383
rect 2061 479 2115 497
rect 2061 445 2071 479
rect 2105 445 2115 479
rect 2061 411 2115 445
rect 2061 377 2071 411
rect 2105 377 2115 411
rect 2061 343 2115 377
rect 2061 309 2071 343
rect 2105 309 2115 343
rect 2061 297 2115 309
rect 2145 485 2199 497
rect 2145 451 2155 485
rect 2189 451 2199 485
rect 2145 417 2199 451
rect 2145 383 2155 417
rect 2189 383 2199 417
rect 2145 297 2199 383
rect 2229 479 2283 497
rect 2229 445 2239 479
rect 2273 445 2283 479
rect 2229 411 2283 445
rect 2229 377 2239 411
rect 2273 377 2283 411
rect 2229 343 2283 377
rect 2229 309 2239 343
rect 2273 309 2283 343
rect 2229 297 2283 309
rect 2313 485 2365 497
rect 2313 451 2323 485
rect 2357 451 2365 485
rect 2313 417 2365 451
rect 2313 383 2323 417
rect 2357 383 2365 417
rect 2313 297 2365 383
<< ndiffc >>
rect 35 131 69 165
rect 35 63 69 97
rect 119 131 153 165
rect 119 63 153 97
rect 223 131 257 165
rect 223 63 257 97
rect 307 63 341 97
rect 391 131 425 165
rect 391 63 425 97
rect 475 63 509 97
rect 559 131 593 165
rect 559 63 593 97
rect 643 63 677 97
rect 727 131 761 165
rect 727 63 761 97
rect 811 63 845 97
rect 895 131 929 165
rect 895 63 929 97
rect 979 63 1013 97
rect 1063 131 1097 165
rect 1063 63 1097 97
rect 1147 63 1181 97
rect 1231 131 1265 165
rect 1231 63 1265 97
rect 1315 63 1349 97
rect 1399 131 1433 165
rect 1399 63 1433 97
rect 1483 63 1517 97
rect 1567 131 1601 165
rect 1567 63 1601 97
rect 1651 63 1685 97
rect 1735 131 1769 165
rect 1735 63 1769 97
rect 1819 63 1853 97
rect 1903 131 1937 165
rect 1903 63 1937 97
rect 1987 63 2021 97
rect 2071 131 2105 165
rect 2071 63 2105 97
rect 2155 63 2189 97
rect 2239 131 2273 165
rect 2239 63 2273 97
rect 2323 63 2357 97
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 119 445 153 479
rect 119 377 153 411
rect 119 309 153 343
rect 223 445 257 479
rect 223 377 257 411
rect 223 309 257 343
rect 307 451 341 485
rect 307 383 341 417
rect 391 445 425 479
rect 391 377 425 411
rect 391 309 425 343
rect 475 451 509 485
rect 475 383 509 417
rect 559 445 593 479
rect 559 377 593 411
rect 559 309 593 343
rect 643 451 677 485
rect 643 383 677 417
rect 727 445 761 479
rect 727 377 761 411
rect 727 309 761 343
rect 811 451 845 485
rect 811 383 845 417
rect 895 445 929 479
rect 895 377 929 411
rect 895 309 929 343
rect 979 451 1013 485
rect 979 383 1013 417
rect 1063 445 1097 479
rect 1063 377 1097 411
rect 1063 309 1097 343
rect 1147 451 1181 485
rect 1147 383 1181 417
rect 1231 445 1265 479
rect 1231 377 1265 411
rect 1231 309 1265 343
rect 1315 451 1349 485
rect 1315 383 1349 417
rect 1399 445 1433 479
rect 1399 377 1433 411
rect 1399 309 1433 343
rect 1483 451 1517 485
rect 1483 383 1517 417
rect 1567 445 1601 479
rect 1567 377 1601 411
rect 1567 309 1601 343
rect 1651 451 1685 485
rect 1651 383 1685 417
rect 1735 445 1769 479
rect 1735 377 1769 411
rect 1735 309 1769 343
rect 1819 451 1853 485
rect 1819 383 1853 417
rect 1903 445 1937 479
rect 1903 377 1937 411
rect 1903 309 1937 343
rect 1987 451 2021 485
rect 1987 383 2021 417
rect 2071 445 2105 479
rect 2071 377 2105 411
rect 2071 309 2105 343
rect 2155 451 2189 485
rect 2155 383 2189 417
rect 2239 445 2273 479
rect 2239 377 2273 411
rect 2239 309 2273 343
rect 2323 451 2357 485
rect 2323 383 2357 417
<< poly >>
rect 79 497 109 523
rect 267 497 297 523
rect 351 497 381 523
rect 435 497 465 523
rect 519 497 549 523
rect 603 497 633 523
rect 687 497 717 523
rect 771 497 801 523
rect 855 497 885 523
rect 939 497 969 523
rect 1023 497 1053 523
rect 1107 497 1137 523
rect 1191 497 1221 523
rect 1275 497 1305 523
rect 1359 497 1389 523
rect 1443 497 1473 523
rect 1527 497 1557 523
rect 1611 497 1641 523
rect 1695 497 1725 523
rect 1779 497 1809 523
rect 1863 497 1893 523
rect 1947 497 1977 523
rect 2031 497 2061 523
rect 2115 497 2145 523
rect 2199 497 2229 523
rect 2283 497 2313 523
rect 79 265 109 297
rect 22 249 109 265
rect 22 215 38 249
rect 72 215 109 249
rect 22 199 109 215
rect 79 177 109 199
rect 267 259 297 297
rect 351 259 381 297
rect 435 259 465 297
rect 267 249 465 259
rect 267 215 307 249
rect 341 215 375 249
rect 409 215 465 249
rect 267 205 465 215
rect 267 177 297 205
rect 351 177 381 205
rect 435 177 465 205
rect 519 259 549 297
rect 603 259 633 297
rect 687 259 717 297
rect 771 259 801 297
rect 855 259 885 297
rect 939 259 969 297
rect 519 249 969 259
rect 519 215 543 249
rect 577 215 611 249
rect 645 215 679 249
rect 713 215 747 249
rect 781 215 815 249
rect 849 215 883 249
rect 917 215 969 249
rect 519 205 969 215
rect 519 177 549 205
rect 603 177 633 205
rect 687 177 717 205
rect 771 177 801 205
rect 855 177 885 205
rect 939 177 969 205
rect 1023 259 1053 297
rect 1107 259 1137 297
rect 1191 259 1221 297
rect 1275 259 1305 297
rect 1359 259 1389 297
rect 1443 259 1473 297
rect 1527 259 1557 297
rect 1611 259 1641 297
rect 1695 259 1725 297
rect 1779 259 1809 297
rect 1863 259 1893 297
rect 1947 259 1977 297
rect 2031 259 2061 297
rect 2115 259 2145 297
rect 2199 259 2229 297
rect 2283 259 2313 297
rect 1023 249 2313 259
rect 1023 215 1043 249
rect 1077 215 1111 249
rect 1145 215 1179 249
rect 1213 215 1247 249
rect 1281 215 1315 249
rect 1349 215 1383 249
rect 1417 215 1451 249
rect 1485 215 1519 249
rect 1553 215 1587 249
rect 1621 215 1655 249
rect 1689 215 1723 249
rect 1757 215 1791 249
rect 1825 215 1859 249
rect 1893 215 1927 249
rect 1961 215 1995 249
rect 2029 215 2063 249
rect 2097 215 2131 249
rect 2165 215 2199 249
rect 2233 215 2313 249
rect 1023 205 2313 215
rect 1023 177 1053 205
rect 1107 177 1137 205
rect 1191 177 1221 205
rect 1275 177 1305 205
rect 1359 177 1389 205
rect 1443 177 1473 205
rect 1527 177 1557 205
rect 1611 177 1641 205
rect 1695 177 1725 205
rect 1779 177 1809 205
rect 1863 177 1893 205
rect 1947 177 1977 205
rect 2031 177 2061 205
rect 2115 177 2145 205
rect 2199 177 2229 205
rect 2283 177 2313 205
rect 79 21 109 47
rect 267 21 297 47
rect 351 21 381 47
rect 435 21 465 47
rect 519 21 549 47
rect 603 21 633 47
rect 687 21 717 47
rect 771 21 801 47
rect 855 21 885 47
rect 939 21 969 47
rect 1023 21 1053 47
rect 1107 21 1137 47
rect 1191 21 1221 47
rect 1275 21 1305 47
rect 1359 21 1389 47
rect 1443 21 1473 47
rect 1527 21 1557 47
rect 1611 21 1641 47
rect 1695 21 1725 47
rect 1779 21 1809 47
rect 1863 21 1893 47
rect 1947 21 1977 47
rect 2031 21 2061 47
rect 2115 21 2145 47
rect 2199 21 2229 47
rect 2283 21 2313 47
<< polycont >>
rect 38 215 72 249
rect 307 215 341 249
rect 375 215 409 249
rect 543 215 577 249
rect 611 215 645 249
rect 679 215 713 249
rect 747 215 781 249
rect 815 215 849 249
rect 883 215 917 249
rect 1043 215 1077 249
rect 1111 215 1145 249
rect 1179 215 1213 249
rect 1247 215 1281 249
rect 1315 215 1349 249
rect 1383 215 1417 249
rect 1451 215 1485 249
rect 1519 215 1553 249
rect 1587 215 1621 249
rect 1655 215 1689 249
rect 1723 215 1757 249
rect 1791 215 1825 249
rect 1859 215 1893 249
rect 1927 215 1961 249
rect 1995 215 2029 249
rect 2063 215 2097 249
rect 2131 215 2165 249
rect 2199 215 2233 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2392 561
rect 35 485 69 527
rect 35 417 69 451
rect 35 349 69 383
rect 35 289 69 315
rect 103 479 169 493
rect 103 445 119 479
rect 153 445 169 479
rect 103 411 169 445
rect 103 377 119 411
rect 153 377 169 411
rect 103 343 169 377
rect 103 309 119 343
rect 153 309 169 343
rect 103 289 169 309
rect 207 479 273 493
rect 207 445 223 479
rect 257 445 273 479
rect 207 411 273 445
rect 207 377 223 411
rect 257 377 273 411
rect 207 343 273 377
rect 307 485 341 527
rect 307 417 341 451
rect 307 357 341 383
rect 375 479 441 493
rect 375 445 391 479
rect 425 445 441 479
rect 375 411 441 445
rect 375 377 391 411
rect 425 377 441 411
rect 207 309 223 343
rect 257 323 273 343
rect 375 343 441 377
rect 475 485 509 527
rect 475 417 509 451
rect 475 357 509 383
rect 543 479 609 493
rect 543 445 559 479
rect 593 445 609 479
rect 543 411 609 445
rect 543 377 559 411
rect 593 377 609 411
rect 375 323 391 343
rect 257 309 391 323
rect 425 323 441 343
rect 543 343 609 377
rect 643 485 677 527
rect 643 417 677 451
rect 643 367 677 383
rect 711 479 777 493
rect 711 445 727 479
rect 761 445 777 479
rect 711 411 777 445
rect 711 377 727 411
rect 761 377 777 411
rect 425 309 509 323
rect 207 289 509 309
rect 543 309 559 343
rect 593 323 609 343
rect 711 343 777 377
rect 811 485 845 527
rect 811 417 845 451
rect 811 367 845 383
rect 879 479 945 493
rect 879 445 895 479
rect 929 445 945 479
rect 879 411 945 445
rect 879 377 895 411
rect 929 377 945 411
rect 711 323 727 343
rect 593 309 727 323
rect 761 323 777 343
rect 879 343 945 377
rect 979 485 1013 527
rect 979 417 1013 451
rect 979 367 1013 383
rect 1047 479 1113 493
rect 1047 445 1063 479
rect 1097 445 1113 479
rect 1047 411 1113 445
rect 1047 377 1063 411
rect 1097 377 1113 411
rect 879 323 895 343
rect 761 309 895 323
rect 929 323 945 343
rect 1047 343 1113 377
rect 1147 485 1181 527
rect 1147 417 1181 451
rect 1147 367 1181 383
rect 1215 479 1281 493
rect 1215 445 1231 479
rect 1265 445 1281 479
rect 1215 411 1281 445
rect 1215 377 1231 411
rect 1265 377 1281 411
rect 929 309 1013 323
rect 543 289 1013 309
rect 1047 309 1063 343
rect 1097 323 1113 343
rect 1215 343 1281 377
rect 1315 485 1349 527
rect 1315 417 1349 451
rect 1315 367 1349 383
rect 1383 479 1449 493
rect 1383 445 1399 479
rect 1433 445 1449 479
rect 1383 411 1449 445
rect 1383 377 1399 411
rect 1433 377 1449 411
rect 1215 323 1231 343
rect 1097 309 1231 323
rect 1265 323 1281 343
rect 1383 343 1449 377
rect 1483 485 1517 527
rect 1483 417 1517 451
rect 1483 367 1517 383
rect 1551 479 1617 493
rect 1551 445 1567 479
rect 1601 445 1617 479
rect 1551 411 1617 445
rect 1551 377 1567 411
rect 1601 377 1617 411
rect 1383 323 1399 343
rect 1265 309 1399 323
rect 1433 323 1449 343
rect 1551 343 1617 377
rect 1651 485 1685 527
rect 1651 417 1685 451
rect 1651 367 1685 383
rect 1719 479 1785 493
rect 1719 445 1735 479
rect 1769 445 1785 479
rect 1719 411 1785 445
rect 1719 377 1735 411
rect 1769 377 1785 411
rect 1551 323 1567 343
rect 1433 309 1567 323
rect 1601 323 1617 343
rect 1719 343 1785 377
rect 1819 485 1853 527
rect 1819 417 1853 451
rect 1819 367 1853 383
rect 1887 479 1953 493
rect 1887 445 1903 479
rect 1937 445 1953 479
rect 1887 411 1953 445
rect 1887 377 1903 411
rect 1937 377 1953 411
rect 1719 323 1735 343
rect 1601 309 1735 323
rect 1769 323 1785 343
rect 1887 343 1953 377
rect 1987 485 2021 527
rect 1987 417 2021 451
rect 1987 367 2021 383
rect 2055 479 2121 493
rect 2055 445 2071 479
rect 2105 445 2121 479
rect 2055 411 2121 445
rect 2055 377 2071 411
rect 2105 377 2121 411
rect 1887 323 1903 343
rect 1769 309 1903 323
rect 1937 323 1953 343
rect 2055 343 2121 377
rect 2155 485 2189 527
rect 2155 417 2189 451
rect 2155 367 2189 383
rect 2223 479 2289 493
rect 2223 445 2239 479
rect 2273 445 2289 479
rect 2223 411 2289 445
rect 2223 377 2239 411
rect 2273 377 2289 411
rect 2055 323 2071 343
rect 1937 309 2071 323
rect 2105 323 2121 343
rect 2223 343 2289 377
rect 2323 485 2357 527
rect 2323 417 2357 451
rect 2323 367 2357 383
rect 2223 323 2239 343
rect 2105 309 2239 323
rect 2273 323 2289 343
rect 2273 309 2375 323
rect 1047 289 2375 309
rect 122 255 169 289
rect 475 255 509 289
rect 978 255 1013 289
rect 22 249 88 255
rect 22 215 38 249
rect 72 215 88 249
rect 122 249 441 255
rect 122 215 307 249
rect 341 215 375 249
rect 409 215 441 249
rect 475 249 937 255
rect 475 215 543 249
rect 577 215 611 249
rect 645 215 679 249
rect 713 215 747 249
rect 781 215 815 249
rect 849 215 883 249
rect 917 215 937 249
rect 978 249 2290 255
rect 978 215 1043 249
rect 1077 215 1111 249
rect 1145 215 1179 249
rect 1213 215 1247 249
rect 1281 215 1315 249
rect 1349 215 1383 249
rect 1417 215 1451 249
rect 1485 215 1519 249
rect 1553 215 1587 249
rect 1621 215 1655 249
rect 1689 215 1723 249
rect 1757 215 1791 249
rect 1825 215 1859 249
rect 1893 215 1927 249
rect 1961 215 1995 249
rect 2029 215 2063 249
rect 2097 215 2131 249
rect 2165 215 2199 249
rect 2233 215 2290 249
rect 122 181 169 215
rect 475 181 509 215
rect 978 181 1013 215
rect 2324 181 2375 289
rect 35 165 69 181
rect 35 97 69 131
rect 35 17 69 63
rect 103 165 169 181
rect 103 131 119 165
rect 153 131 169 165
rect 103 97 169 131
rect 103 63 119 97
rect 153 63 169 97
rect 103 52 169 63
rect 207 165 509 181
rect 207 131 223 165
rect 257 147 391 165
rect 257 131 273 147
rect 207 97 273 131
rect 375 131 391 147
rect 425 147 509 165
rect 543 165 1013 181
rect 425 131 441 147
rect 207 63 223 97
rect 257 63 273 97
rect 207 52 273 63
rect 307 97 341 113
rect 307 17 341 63
rect 375 97 441 131
rect 543 131 559 165
rect 593 147 727 165
rect 593 131 609 147
rect 375 63 391 97
rect 425 63 441 97
rect 375 52 441 63
rect 475 97 509 113
rect 475 17 509 63
rect 543 97 609 131
rect 711 131 727 147
rect 761 147 895 165
rect 761 131 777 147
rect 543 63 559 97
rect 593 63 609 97
rect 543 52 609 63
rect 643 97 677 113
rect 643 17 677 63
rect 711 97 777 131
rect 879 131 895 147
rect 929 147 1013 165
rect 1047 165 2375 181
rect 929 131 945 147
rect 711 63 727 97
rect 761 63 777 97
rect 711 52 777 63
rect 811 97 845 113
rect 811 17 845 63
rect 879 97 945 131
rect 1047 131 1063 165
rect 1097 147 1231 165
rect 1097 131 1113 147
rect 879 63 895 97
rect 929 63 945 97
rect 879 52 945 63
rect 979 97 1013 113
rect 979 17 1013 63
rect 1047 97 1113 131
rect 1215 131 1231 147
rect 1265 147 1399 165
rect 1265 131 1281 147
rect 1047 63 1063 97
rect 1097 63 1113 97
rect 1047 52 1113 63
rect 1147 97 1181 113
rect 1047 51 1097 52
rect 1147 17 1181 63
rect 1215 97 1281 131
rect 1383 131 1399 147
rect 1433 147 1567 165
rect 1433 131 1449 147
rect 1215 63 1231 97
rect 1265 63 1281 97
rect 1215 52 1281 63
rect 1315 97 1349 113
rect 1231 51 1265 52
rect 1315 17 1349 63
rect 1383 97 1449 131
rect 1551 131 1567 147
rect 1601 147 1735 165
rect 1601 131 1617 147
rect 1383 63 1399 97
rect 1433 63 1449 97
rect 1383 52 1449 63
rect 1483 97 1517 113
rect 1399 51 1433 52
rect 1483 17 1517 63
rect 1551 97 1617 131
rect 1719 131 1735 147
rect 1769 147 1903 165
rect 1769 131 1785 147
rect 1551 63 1567 97
rect 1601 63 1617 97
rect 1551 52 1617 63
rect 1651 97 1685 113
rect 1651 17 1685 63
rect 1719 97 1785 131
rect 1887 131 1903 147
rect 1937 147 2071 165
rect 1937 131 1953 147
rect 1719 63 1735 97
rect 1769 63 1785 97
rect 1719 52 1785 63
rect 1819 97 1853 113
rect 1819 17 1853 63
rect 1887 97 1953 131
rect 2055 131 2071 147
rect 2105 147 2239 165
rect 2105 131 2121 147
rect 1887 63 1903 97
rect 1937 63 1953 97
rect 1887 52 1953 63
rect 1987 97 2021 113
rect 1987 17 2021 63
rect 2055 97 2121 131
rect 2223 131 2239 147
rect 2273 147 2375 165
rect 2273 131 2289 147
rect 2055 63 2071 97
rect 2105 63 2121 97
rect 2055 52 2121 63
rect 2155 97 2189 113
rect 2155 17 2189 63
rect 2223 97 2289 131
rect 2223 63 2239 97
rect 2273 63 2289 97
rect 2223 52 2289 63
rect 2323 97 2357 113
rect 2323 17 2357 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2392 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
<< metal1 >>
rect 0 561 2392 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2392 561
rect 0 496 2392 527
rect 0 17 2392 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2392 17
rect 0 -48 2392 -17
<< labels >>
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 2334 221 2368 255 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 2334 289 2368 323 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 bufbuf_16
rlabel metal1 s 0 -48 2392 48 1 VGND
port 2 nsew ground bidirectional abutment
rlabel metal1 s 0 496 2392 592 1 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2392 544
string GDS_END 3243022
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3224820
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 59.800 0.000 
<< end >>
