magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -51 355 483 1087
<< pwell >>
rect -11 -103 443 149
<< mvnmos >>
rect 68 -77 188 123
rect 244 -77 364 123
<< mvpmos >>
rect 68 421 188 1021
rect 244 421 364 1021
<< mvndiff >>
rect 15 111 68 123
rect 15 77 23 111
rect 57 77 68 111
rect 15 43 68 77
rect 15 9 23 43
rect 57 9 68 43
rect 15 -25 68 9
rect 15 -59 23 -25
rect 57 -59 68 -25
rect 15 -77 68 -59
rect 188 -77 244 123
rect 364 111 417 123
rect 364 77 375 111
rect 409 77 417 111
rect 364 43 417 77
rect 364 9 375 43
rect 409 9 417 43
rect 364 -25 417 9
rect 364 -59 375 -25
rect 409 -59 417 -25
rect 364 -77 417 -59
<< mvpdiff >>
rect 15 1009 68 1021
rect 15 975 23 1009
rect 57 975 68 1009
rect 15 941 68 975
rect 15 907 23 941
rect 57 907 68 941
rect 15 873 68 907
rect 15 839 23 873
rect 57 839 68 873
rect 15 805 68 839
rect 15 771 23 805
rect 57 771 68 805
rect 15 737 68 771
rect 15 703 23 737
rect 57 703 68 737
rect 15 669 68 703
rect 15 635 23 669
rect 57 635 68 669
rect 15 601 68 635
rect 15 567 23 601
rect 57 567 68 601
rect 15 533 68 567
rect 15 499 23 533
rect 57 499 68 533
rect 15 421 68 499
rect 188 1009 244 1021
rect 188 975 199 1009
rect 233 975 244 1009
rect 188 941 244 975
rect 188 907 199 941
rect 233 907 244 941
rect 188 873 244 907
rect 188 839 199 873
rect 233 839 244 873
rect 188 805 244 839
rect 188 771 199 805
rect 233 771 244 805
rect 188 737 244 771
rect 188 703 199 737
rect 233 703 244 737
rect 188 669 244 703
rect 188 635 199 669
rect 233 635 244 669
rect 188 601 244 635
rect 188 567 199 601
rect 233 567 244 601
rect 188 533 244 567
rect 188 499 199 533
rect 233 499 244 533
rect 188 421 244 499
rect 364 1009 417 1021
rect 364 975 375 1009
rect 409 975 417 1009
rect 364 941 417 975
rect 364 907 375 941
rect 409 907 417 941
rect 364 873 417 907
rect 364 839 375 873
rect 409 839 417 873
rect 364 805 417 839
rect 364 771 375 805
rect 409 771 417 805
rect 364 737 417 771
rect 364 703 375 737
rect 409 703 417 737
rect 364 669 417 703
rect 364 635 375 669
rect 409 635 417 669
rect 364 601 417 635
rect 364 567 375 601
rect 409 567 417 601
rect 364 533 417 567
rect 364 499 375 533
rect 409 499 417 533
rect 364 421 417 499
<< mvndiffc >>
rect 23 77 57 111
rect 23 9 57 43
rect 23 -59 57 -25
rect 375 77 409 111
rect 375 9 409 43
rect 375 -59 409 -25
<< mvpdiffc >>
rect 23 975 57 1009
rect 23 907 57 941
rect 23 839 57 873
rect 23 771 57 805
rect 23 703 57 737
rect 23 635 57 669
rect 23 567 57 601
rect 23 499 57 533
rect 199 975 233 1009
rect 199 907 233 941
rect 199 839 233 873
rect 199 771 233 805
rect 199 703 233 737
rect 199 635 233 669
rect 199 567 233 601
rect 199 499 233 533
rect 375 975 409 1009
rect 375 907 409 941
rect 375 839 409 873
rect 375 771 409 805
rect 375 703 409 737
rect 375 635 409 669
rect 375 567 409 601
rect 375 499 409 533
<< poly >>
rect 68 1021 188 1047
rect 244 1021 364 1047
rect 68 307 188 421
rect 68 273 104 307
rect 138 273 188 307
rect 68 239 188 273
rect 68 205 104 239
rect 138 205 188 239
rect 68 123 188 205
rect 244 300 364 421
rect 244 266 288 300
rect 322 266 364 300
rect 244 232 364 266
rect 244 198 288 232
rect 322 198 364 232
rect 244 123 364 198
rect 68 -103 188 -77
rect 244 -103 364 -77
<< polycont >>
rect 104 273 138 307
rect 104 205 138 239
rect 288 266 322 300
rect 288 198 322 232
<< locali >>
rect 23 1055 57 1095
rect 375 1055 409 1095
rect 23 1009 57 1021
rect 23 941 57 949
rect 23 873 57 907
rect 23 805 57 839
rect 23 737 57 771
rect 23 669 57 703
rect 23 601 57 635
rect 23 533 57 567
rect 23 483 57 499
rect 199 1009 233 1025
rect 199 941 233 975
rect 199 873 233 907
rect 199 805 233 839
rect 199 737 233 771
rect 199 669 233 703
rect 199 601 233 635
rect 199 533 233 567
rect 88 273 104 307
rect 138 273 154 307
rect 88 239 154 273
rect 88 205 104 239
rect 138 205 154 239
rect 199 127 233 499
rect 375 1009 409 1021
rect 375 941 409 949
rect 375 873 409 907
rect 375 805 409 839
rect 375 737 409 771
rect 375 669 409 703
rect 375 601 409 635
rect 375 533 409 567
rect 375 483 409 499
rect 272 266 288 300
rect 322 266 338 300
rect 272 232 338 266
rect 272 198 288 232
rect 322 198 338 232
rect 23 111 233 127
rect 57 77 233 111
rect 23 43 233 77
rect 57 24 233 43
rect 375 111 409 127
rect 375 43 409 77
rect 23 -25 57 9
rect 23 -75 57 -59
rect 375 -22 409 9
rect 375 -94 409 -59
rect 375 -166 409 -128
<< viali >>
rect 23 1021 57 1055
rect 23 975 57 983
rect 23 949 57 975
rect 375 1021 409 1055
rect 375 975 409 983
rect 375 949 409 975
rect 375 -25 409 -22
rect 375 -56 409 -25
rect 375 -128 409 -94
rect 375 -200 409 -166
<< metal1 >>
rect -57 1055 482 1195
rect -57 1021 23 1055
rect 57 1021 375 1055
rect 409 1021 482 1055
rect -57 983 482 1021
rect -57 949 23 983
rect 57 949 375 983
rect 409 949 482 983
rect -57 937 482 949
rect -57 -22 473 -10
rect -57 -56 375 -22
rect 409 -56 473 -22
rect -57 -94 473 -56
rect -57 -128 375 -94
rect 409 -128 473 -94
rect -57 -166 473 -128
rect -57 -200 375 -166
rect 409 -200 473 -166
rect -57 -212 473 -200
use sky130_fd_pr__model__nfet_highvoltage__example_55959141808144  sky130_fd_pr__model__nfet_highvoltage__example_55959141808144_0
timestamp 1701704242
transform -1 0 364 0 -1 123
box -1 0 0 1
use sky130_fd_pr__model__nfet_highvoltage__example_55959141808144  sky130_fd_pr__model__nfet_highvoltage__example_55959141808144_1
timestamp 1701704242
transform 1 0 68 0 -1 123
box -1 0 0 1
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808142  sky130_fd_pr__model__pfet_highvoltage__example_55959141808142_0
timestamp 1701704242
transform 1 0 68 0 -1 1021
box -1 0 297 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1701704242
transform 0 -1 57 -1 0 1055
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_1
timestamp 1701704242
transform 0 -1 409 -1 0 1055
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_0
timestamp 1701704242
transform 0 -1 409 -1 0 -22
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_0
timestamp 1701704242
transform 0 1 88 1 0 189
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_1
timestamp 1701704242
transform 0 1 272 1 0 182
box 0 0 1 1
<< properties >>
string GDS_END 68182316
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 68181128
<< end >>
