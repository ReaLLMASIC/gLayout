magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -38 261 2062 582
<< pwell >>
rect 1174 157 1356 201
rect 1659 157 2023 203
rect 1 145 824 157
rect 1028 145 2023 157
rect 1 21 2023 145
rect 29 -17 63 21
<< locali >>
rect 19 195 89 325
rect 356 157 390 337
rect 492 271 558 337
rect 616 157 650 223
rect 706 207 804 331
rect 356 123 650 157
rect 495 61 530 123
rect 1852 301 1921 479
rect 1887 164 1921 301
rect 1852 61 1921 164
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 36 393 70 493
rect 104 427 170 527
rect 36 359 169 393
rect 123 194 169 359
rect 123 161 162 194
rect 35 127 162 161
rect 204 143 249 493
rect 35 69 69 127
rect 103 17 169 93
rect 203 69 249 143
rect 287 415 342 489
rect 376 449 442 527
rect 538 449 717 483
rect 287 372 649 415
rect 287 89 321 372
rect 424 225 458 372
rect 615 337 649 372
rect 683 399 717 449
rect 751 433 785 527
rect 842 413 889 488
rect 938 438 1152 472
rect 842 399 876 413
rect 683 365 876 399
rect 615 271 654 337
rect 424 191 492 225
rect 842 173 876 365
rect 684 139 876 173
rect 910 207 958 381
rect 996 331 1084 402
rect 1118 315 1152 438
rect 1186 367 1220 527
rect 1254 427 1304 493
rect 1349 433 1526 467
rect 1118 297 1220 315
rect 1060 263 1220 297
rect 910 141 1026 207
rect 287 55 361 89
rect 395 17 461 89
rect 684 89 718 139
rect 842 107 876 139
rect 1060 107 1094 263
rect 1186 249 1220 263
rect 1128 213 1162 219
rect 1254 213 1288 427
rect 1322 249 1360 393
rect 1394 315 1458 381
rect 1128 153 1288 213
rect 1394 207 1432 315
rect 1492 281 1526 433
rect 1562 427 1623 527
rect 1693 381 1747 491
rect 1560 315 1747 381
rect 1781 325 1816 527
rect 564 55 718 89
rect 752 17 792 105
rect 842 73 912 107
rect 946 73 1094 107
rect 1144 17 1218 117
rect 1254 107 1288 153
rect 1322 141 1432 207
rect 1466 265 1526 281
rect 1713 265 1747 315
rect 1466 199 1679 265
rect 1713 199 1853 265
rect 1466 107 1500 199
rect 1713 165 1747 199
rect 1254 73 1346 107
rect 1392 73 1500 107
rect 1549 17 1623 123
rect 1677 60 1747 165
rect 1955 281 1989 527
rect 1781 17 1815 139
rect 1955 17 1989 186
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
<< metal1 >>
rect 0 561 2024 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 0 496 2024 527
rect 0 17 2024 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
rect 0 -48 2024 -17
<< obsm1 >>
rect 116 388 174 397
rect 1029 388 1087 397
rect 1312 388 1370 397
rect 116 360 1370 388
rect 116 351 174 360
rect 1029 351 1087 360
rect 1312 351 1370 360
rect 198 184 256 193
rect 937 184 995 193
rect 1314 184 1372 193
rect 198 156 1372 184
rect 198 147 256 156
rect 937 147 995 156
rect 1314 147 1372 156
<< labels >>
rlabel locali s 19 195 89 325 6 CLK
port 1 nsew clock input
rlabel locali s 492 271 558 337 6 D
port 2 nsew signal input
rlabel locali s 706 207 804 331 6 SCD
port 3 nsew signal input
rlabel locali s 495 61 530 123 6 SCE
port 4 nsew signal input
rlabel locali s 356 123 650 157 6 SCE
port 4 nsew signal input
rlabel locali s 616 157 650 223 6 SCE
port 4 nsew signal input
rlabel locali s 356 157 390 337 6 SCE
port 4 nsew signal input
rlabel metal1 s 0 -48 2024 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1 21 2023 145 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1028 145 2023 157 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1 145 824 157 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1659 157 2023 203 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1174 157 1356 201 6 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 2062 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 2024 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 1852 61 1921 164 6 Q
port 9 nsew signal output
rlabel locali s 1887 164 1921 301 6 Q
port 9 nsew signal output
rlabel locali s 1852 301 1921 479 6 Q
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 2024 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 392160
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 376362
<< end >>
