magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< nwell >>
rect 0 1331 3633 2349
<< pwell >>
rect 561 888 813 1240
rect 123 101 213 846
rect 3543 101 3633 846
rect 123 10 3633 101
<< mvnmos >>
rect 637 914 737 1214
<< mvndiff >>
rect 587 914 637 1214
rect 737 914 787 1214
<< mvpsubdiff >>
rect 149 796 187 820
rect 149 762 151 796
rect 185 762 187 796
rect 149 728 187 762
rect 149 694 151 728
rect 185 694 187 728
rect 149 660 187 694
rect 149 626 151 660
rect 185 626 187 660
rect 149 592 187 626
rect 149 558 151 592
rect 185 558 187 592
rect 149 524 187 558
rect 149 490 151 524
rect 185 490 187 524
rect 149 456 187 490
rect 149 422 151 456
rect 185 422 187 456
rect 149 388 187 422
rect 149 354 151 388
rect 185 354 187 388
rect 149 320 187 354
rect 149 286 151 320
rect 185 286 187 320
rect 149 252 187 286
rect 149 218 151 252
rect 185 218 187 252
rect 149 184 187 218
rect 3569 796 3607 820
rect 3569 762 3571 796
rect 3605 762 3607 796
rect 3569 728 3607 762
rect 3569 694 3571 728
rect 3605 694 3607 728
rect 3569 660 3607 694
rect 3569 626 3571 660
rect 3605 626 3607 660
rect 3569 592 3607 626
rect 3569 558 3571 592
rect 3605 558 3607 592
rect 3569 524 3607 558
rect 3569 490 3571 524
rect 3605 490 3607 524
rect 3569 456 3607 490
rect 3569 422 3571 456
rect 3605 422 3607 456
rect 3569 388 3607 422
rect 3569 354 3571 388
rect 3605 354 3607 388
rect 3569 320 3607 354
rect 3569 286 3571 320
rect 3605 286 3607 320
rect 3569 252 3607 286
rect 3569 218 3571 252
rect 3605 218 3607 252
rect 149 150 151 184
rect 185 150 187 184
rect 149 75 187 150
rect 3569 184 3607 218
rect 3569 150 3571 184
rect 3605 150 3607 184
rect 3569 75 3607 150
rect 149 72 3607 75
rect 149 38 193 72
rect 227 38 261 72
rect 295 38 329 72
rect 363 38 397 72
rect 431 38 465 72
rect 499 38 533 72
rect 567 38 601 72
rect 635 38 669 72
rect 703 38 737 72
rect 771 38 805 72
rect 839 38 873 72
rect 907 38 941 72
rect 975 38 1009 72
rect 1043 38 1077 72
rect 1111 38 1145 72
rect 1179 38 1213 72
rect 1247 38 1281 72
rect 1315 38 1349 72
rect 1383 38 1417 72
rect 1451 38 1485 72
rect 1519 38 1553 72
rect 1587 38 1621 72
rect 1655 38 1689 72
rect 1723 38 1757 72
rect 1791 38 1825 72
rect 1859 38 1893 72
rect 1927 38 1961 72
rect 1995 38 2029 72
rect 2063 38 2097 72
rect 2131 38 2165 72
rect 2199 38 2233 72
rect 2267 38 2301 72
rect 2335 38 2369 72
rect 2403 38 2437 72
rect 2471 38 2505 72
rect 2539 38 2573 72
rect 2607 38 2641 72
rect 2675 38 2709 72
rect 2743 38 2777 72
rect 2811 38 2845 72
rect 2879 38 2913 72
rect 2947 38 2981 72
rect 3015 38 3049 72
rect 3083 38 3117 72
rect 3151 38 3185 72
rect 3219 38 3253 72
rect 3287 38 3321 72
rect 3355 38 3389 72
rect 3423 38 3457 72
rect 3491 38 3525 72
rect 3559 38 3607 72
rect 149 36 3607 38
<< mvnsubdiff >>
rect 92 2281 3098 2283
rect 92 2247 116 2281
rect 150 2247 184 2281
rect 218 2247 252 2281
rect 286 2247 320 2281
rect 354 2247 388 2281
rect 422 2247 456 2281
rect 490 2247 524 2281
rect 558 2247 592 2281
rect 626 2247 660 2281
rect 694 2247 728 2281
rect 762 2247 796 2281
rect 830 2247 864 2281
rect 898 2247 932 2281
rect 966 2247 1000 2281
rect 1034 2247 1068 2281
rect 1102 2247 1136 2281
rect 1170 2247 1204 2281
rect 1238 2247 1272 2281
rect 1306 2247 1340 2281
rect 1374 2247 1408 2281
rect 1442 2247 1476 2281
rect 1510 2247 1544 2281
rect 1578 2247 1612 2281
rect 1646 2247 1680 2281
rect 1714 2247 1748 2281
rect 1782 2247 1816 2281
rect 1850 2247 1884 2281
rect 1918 2247 1952 2281
rect 1986 2247 2020 2281
rect 2054 2247 2088 2281
rect 2122 2247 2156 2281
rect 2190 2247 2224 2281
rect 2258 2247 2292 2281
rect 2326 2247 2360 2281
rect 2394 2247 2428 2281
rect 2462 2247 2496 2281
rect 2530 2247 2564 2281
rect 2598 2247 2632 2281
rect 2666 2247 2700 2281
rect 2734 2247 2768 2281
rect 2802 2247 2836 2281
rect 2870 2247 2904 2281
rect 2938 2247 2972 2281
rect 3006 2247 3040 2281
rect 3074 2247 3098 2281
rect 92 2245 3098 2247
rect 2608 2181 3098 2245
<< mvpsubdiffcont >>
rect 151 762 185 796
rect 151 694 185 728
rect 151 626 185 660
rect 151 558 185 592
rect 151 490 185 524
rect 151 422 185 456
rect 151 354 185 388
rect 151 286 185 320
rect 151 218 185 252
rect 3571 762 3605 796
rect 3571 694 3605 728
rect 3571 626 3605 660
rect 3571 558 3605 592
rect 3571 490 3605 524
rect 3571 422 3605 456
rect 3571 354 3605 388
rect 3571 286 3605 320
rect 3571 218 3605 252
rect 151 150 185 184
rect 3571 150 3605 184
rect 193 38 227 72
rect 261 38 295 72
rect 329 38 363 72
rect 397 38 431 72
rect 465 38 499 72
rect 533 38 567 72
rect 601 38 635 72
rect 669 38 703 72
rect 737 38 771 72
rect 805 38 839 72
rect 873 38 907 72
rect 941 38 975 72
rect 1009 38 1043 72
rect 1077 38 1111 72
rect 1145 38 1179 72
rect 1213 38 1247 72
rect 1281 38 1315 72
rect 1349 38 1383 72
rect 1417 38 1451 72
rect 1485 38 1519 72
rect 1553 38 1587 72
rect 1621 38 1655 72
rect 1689 38 1723 72
rect 1757 38 1791 72
rect 1825 38 1859 72
rect 1893 38 1927 72
rect 1961 38 1995 72
rect 2029 38 2063 72
rect 2097 38 2131 72
rect 2165 38 2199 72
rect 2233 38 2267 72
rect 2301 38 2335 72
rect 2369 38 2403 72
rect 2437 38 2471 72
rect 2505 38 2539 72
rect 2573 38 2607 72
rect 2641 38 2675 72
rect 2709 38 2743 72
rect 2777 38 2811 72
rect 2845 38 2879 72
rect 2913 38 2947 72
rect 2981 38 3015 72
rect 3049 38 3083 72
rect 3117 38 3151 72
rect 3185 38 3219 72
rect 3253 38 3287 72
rect 3321 38 3355 72
rect 3389 38 3423 72
rect 3457 38 3491 72
rect 3525 38 3559 72
<< mvnsubdiffcont >>
rect 116 2247 150 2281
rect 184 2247 218 2281
rect 252 2247 286 2281
rect 320 2247 354 2281
rect 388 2247 422 2281
rect 456 2247 490 2281
rect 524 2247 558 2281
rect 592 2247 626 2281
rect 660 2247 694 2281
rect 728 2247 762 2281
rect 796 2247 830 2281
rect 864 2247 898 2281
rect 932 2247 966 2281
rect 1000 2247 1034 2281
rect 1068 2247 1102 2281
rect 1136 2247 1170 2281
rect 1204 2247 1238 2281
rect 1272 2247 1306 2281
rect 1340 2247 1374 2281
rect 1408 2247 1442 2281
rect 1476 2247 1510 2281
rect 1544 2247 1578 2281
rect 1612 2247 1646 2281
rect 1680 2247 1714 2281
rect 1748 2247 1782 2281
rect 1816 2247 1850 2281
rect 1884 2247 1918 2281
rect 1952 2247 1986 2281
rect 2020 2247 2054 2281
rect 2088 2247 2122 2281
rect 2156 2247 2190 2281
rect 2224 2247 2258 2281
rect 2292 2247 2326 2281
rect 2360 2247 2394 2281
rect 2428 2247 2462 2281
rect 2496 2247 2530 2281
rect 2564 2247 2598 2281
rect 2632 2247 2666 2281
rect 2700 2247 2734 2281
rect 2768 2247 2802 2281
rect 2836 2247 2870 2281
rect 2904 2247 2938 2281
rect 2972 2247 3006 2281
rect 3040 2247 3074 2281
<< poly >>
rect 445 2191 579 2207
rect 445 2157 461 2191
rect 495 2157 529 2191
rect 563 2157 579 2191
rect 445 2141 579 2157
rect 462 2124 562 2141
rect 821 1912 2187 1988
rect 2280 1926 2421 1942
rect 2280 1892 2296 1926
rect 2330 1892 2364 1926
rect 2398 1892 2421 1926
rect 2280 1876 2421 1892
rect 150 1850 250 1872
rect 150 1816 184 1850
rect 218 1816 250 1850
rect 150 1782 250 1816
rect 150 1748 184 1782
rect 218 1748 250 1782
rect 150 1714 250 1748
rect 306 1850 406 1872
rect 306 1816 340 1850
rect 374 1816 406 1850
rect 618 1847 718 1872
rect 2321 1870 2421 1876
rect 2587 1870 3155 1946
rect 306 1782 406 1816
rect 306 1748 340 1782
rect 374 1748 406 1782
rect 600 1831 734 1847
rect 600 1797 616 1831
rect 650 1797 684 1831
rect 718 1797 734 1831
rect 600 1781 734 1797
rect 306 1732 406 1748
rect 150 1680 184 1714
rect 218 1690 250 1714
rect 218 1680 406 1690
rect 150 1623 406 1680
rect 483 1679 2155 1695
rect 483 1645 527 1679
rect 561 1645 595 1679
rect 629 1645 663 1679
rect 697 1645 731 1679
rect 765 1645 982 1679
rect 1016 1645 1050 1679
rect 1084 1645 1118 1679
rect 1152 1645 1186 1679
rect 1220 1645 1483 1679
rect 1517 1645 1551 1679
rect 1585 1645 2155 1679
rect 483 1623 2155 1645
rect 150 1240 380 1371
rect 620 1313 754 1329
rect 423 1296 578 1312
rect 423 1262 460 1296
rect 494 1262 528 1296
rect 562 1262 578 1296
rect 620 1279 636 1313
rect 670 1279 704 1313
rect 738 1279 754 1313
rect 620 1263 754 1279
rect 796 1296 951 1312
rect 423 1240 578 1262
rect 637 1214 737 1263
rect 796 1262 812 1296
rect 846 1262 880 1296
rect 914 1262 951 1296
rect 796 1240 951 1262
rect 1131 1100 1833 1371
rect 3197 1196 3575 1218
rect 1913 1100 3155 1172
rect 3197 1162 3217 1196
rect 3251 1162 3285 1196
rect 3319 1162 3453 1196
rect 3487 1162 3521 1196
rect 3555 1162 3575 1196
rect 3197 1142 3575 1162
rect 637 888 737 914
rect 1672 846 2240 922
rect 314 118 882 194
rect 1048 118 1616 194
rect 2296 173 2396 194
rect 2279 157 2413 173
rect 2279 123 2295 157
rect 2329 123 2363 157
rect 2397 123 2413 157
rect 2279 107 2413 123
rect 2467 172 2708 194
rect 2467 138 2491 172
rect 2525 138 2559 172
rect 2593 138 2627 172
rect 2661 138 2708 172
rect 2467 118 2708 138
rect 2874 172 3130 194
rect 2874 138 2910 172
rect 2944 138 2978 172
rect 3012 138 3046 172
rect 3080 138 3130 172
rect 2874 118 3130 138
rect 3186 172 3442 194
rect 3186 138 3222 172
rect 3256 138 3290 172
rect 3324 138 3358 172
rect 3392 138 3442 172
rect 3186 118 3442 138
<< polycont >>
rect 461 2157 495 2191
rect 529 2157 563 2191
rect 2296 1892 2330 1926
rect 2364 1892 2398 1926
rect 184 1816 218 1850
rect 184 1748 218 1782
rect 340 1816 374 1850
rect 340 1748 374 1782
rect 616 1797 650 1831
rect 684 1797 718 1831
rect 184 1680 218 1714
rect 527 1645 561 1679
rect 595 1645 629 1679
rect 663 1645 697 1679
rect 731 1645 765 1679
rect 982 1645 1016 1679
rect 1050 1645 1084 1679
rect 1118 1645 1152 1679
rect 1186 1645 1220 1679
rect 1483 1645 1517 1679
rect 1551 1645 1585 1679
rect 460 1262 494 1296
rect 528 1262 562 1296
rect 636 1279 670 1313
rect 704 1279 738 1313
rect 812 1262 846 1296
rect 880 1262 914 1296
rect 3217 1162 3251 1196
rect 3285 1162 3319 1196
rect 3453 1162 3487 1196
rect 3521 1162 3555 1196
rect 2295 123 2329 157
rect 2363 123 2397 157
rect 2491 138 2525 172
rect 2559 138 2593 172
rect 2627 138 2661 172
rect 2910 138 2944 172
rect 2978 138 3012 172
rect 3046 138 3080 172
rect 3222 138 3256 172
rect 3290 138 3324 172
rect 3358 138 3392 172
<< locali >>
rect 100 2247 116 2281
rect 150 2247 184 2281
rect 218 2247 252 2281
rect 286 2247 320 2281
rect 354 2247 388 2281
rect 422 2247 456 2281
rect 490 2247 524 2281
rect 558 2247 592 2281
rect 626 2247 660 2281
rect 694 2247 728 2281
rect 762 2247 796 2281
rect 830 2247 864 2281
rect 898 2247 932 2281
rect 966 2247 1000 2281
rect 1034 2247 1068 2281
rect 1102 2247 1136 2281
rect 1170 2247 1204 2281
rect 1238 2247 1272 2281
rect 1306 2247 1340 2281
rect 1374 2247 1408 2281
rect 1442 2247 1476 2281
rect 1510 2247 1544 2281
rect 1578 2247 1612 2281
rect 1646 2247 1680 2281
rect 1714 2247 1748 2281
rect 1782 2247 1816 2281
rect 1850 2247 1884 2281
rect 1918 2247 1952 2281
rect 1986 2247 2020 2281
rect 2054 2247 2088 2281
rect 2122 2247 2156 2281
rect 2190 2247 2224 2281
rect 2258 2247 2292 2281
rect 2326 2247 2360 2281
rect 2394 2247 2428 2281
rect 2462 2247 2496 2281
rect 2530 2247 2564 2281
rect 2598 2247 2632 2281
rect 2666 2247 2700 2281
rect 2734 2247 2768 2281
rect 2802 2247 2836 2281
rect 2870 2247 2904 2281
rect 2938 2247 2972 2281
rect 3006 2247 3040 2281
rect 3074 2247 3090 2281
rect 105 2107 139 2247
rect 339 2153 377 2187
rect 445 2157 461 2191
rect 329 2098 411 2153
rect 105 2035 139 2073
rect 261 2007 295 2045
rect 329 1906 461 2098
rect 105 1595 139 1894
rect 184 1850 218 1866
rect 184 1782 218 1816
rect 340 1850 374 1866
rect 340 1782 374 1816
rect 218 1715 256 1749
rect 184 1714 218 1715
rect 184 1664 218 1680
rect 105 1523 139 1561
rect 105 1451 139 1489
rect 215 845 295 1595
rect 340 1296 374 1748
rect 417 1595 461 1906
rect 495 1986 529 2191
rect 563 2157 579 2191
rect 729 2147 763 2247
rect 2616 2157 3090 2247
rect 729 2075 763 2113
rect 2432 1973 2466 2014
rect 495 1914 529 1952
rect 623 1902 661 1936
rect 556 1797 616 1831
rect 650 1797 684 1831
rect 718 1797 734 1831
rect 556 1764 662 1797
rect 590 1730 628 1764
rect 511 1645 527 1679
rect 561 1645 595 1679
rect 629 1645 663 1679
rect 697 1645 731 1679
rect 765 1645 781 1679
rect 417 1561 438 1595
rect 417 1523 472 1561
rect 417 1489 438 1523
rect 417 1451 472 1489
rect 417 1417 438 1451
rect 858 1545 932 1864
rect 966 1645 982 1679
rect 1016 1645 1050 1679
rect 1084 1645 1118 1679
rect 1152 1645 1186 1679
rect 1220 1645 1236 1679
rect 858 1511 870 1545
rect 904 1511 932 1545
rect 858 1473 932 1511
rect 858 1439 870 1473
rect 904 1439 932 1473
rect 417 1393 461 1417
rect 858 1393 932 1439
rect 1270 1545 1427 1864
rect 1467 1645 1483 1679
rect 1517 1645 1551 1679
rect 1585 1645 1601 1679
rect 1641 1675 2095 1965
rect 2276 1926 2398 1942
rect 2432 1939 2444 1973
rect 2478 1939 2516 1973
rect 2276 1892 2296 1926
rect 2330 1892 2364 1926
rect 2276 1876 2398 1892
rect 2276 1819 2310 1876
rect 2238 1785 2276 1819
rect 2276 1782 2310 1785
rect 2432 1859 2624 1895
rect 2432 1756 2466 1859
rect 1675 1641 1713 1675
rect 1747 1641 1785 1675
rect 1819 1641 1857 1675
rect 1891 1641 1929 1675
rect 1963 1641 2001 1675
rect 2035 1641 2073 1675
rect 2094 1595 2200 1597
rect 1270 1511 1302 1545
rect 1336 1511 1427 1545
rect 1270 1473 1427 1511
rect 1270 1439 1302 1473
rect 1336 1439 1427 1473
rect 1270 1393 1427 1439
rect 1734 1523 1768 1561
rect 1734 1451 1768 1489
rect 654 1381 688 1393
rect 688 1347 726 1381
rect 1086 1371 1120 1393
rect 1518 1371 1552 1393
rect 1950 1371 1984 1393
rect 1086 1337 1098 1371
rect 1132 1337 1170 1371
rect 1518 1337 1556 1371
rect 1912 1337 1950 1371
rect 340 1262 456 1296
rect 494 1262 528 1296
rect 562 1262 578 1296
rect 620 1279 636 1313
rect 670 1279 704 1313
rect 738 1296 754 1313
rect 1086 1296 1204 1337
rect 742 1279 754 1296
rect 670 1262 708 1279
rect 796 1262 812 1296
rect 846 1262 880 1296
rect 918 1262 930 1296
rect 1086 1262 1098 1296
rect 1132 1262 1170 1296
rect 2094 1156 2200 1417
rect 2542 1595 2576 1617
rect 2542 1523 2576 1561
rect 2542 1451 2576 1489
rect 2854 1523 2888 1561
rect 2854 1451 2888 1489
rect 3213 1523 3247 1561
rect 3213 1451 3247 1489
rect 3525 1523 3559 1561
rect 3525 1451 3559 1489
rect 2542 1156 2576 1417
rect 2698 1171 2732 1240
rect 3010 1171 3044 1240
rect 2697 1137 2735 1171
rect 2972 1137 3010 1171
rect 3201 1177 3217 1196
rect 3201 1162 3213 1177
rect 3251 1162 3285 1196
rect 3319 1162 3335 1196
rect 3247 1143 3285 1162
rect 438 997 472 1035
rect 438 925 472 963
rect 1012 845 1046 1012
rect 1868 997 1902 1035
rect 3369 941 3403 1240
rect 3437 1162 3453 1196
rect 3487 1162 3521 1196
rect 3555 1177 3571 1196
rect 3559 1162 3571 1177
rect 3487 1143 3525 1162
rect 2985 907 3403 941
rect 215 831 219 845
rect 151 796 185 812
rect 253 811 291 845
rect 325 811 363 845
rect 1012 811 1067 845
rect 1101 811 1139 845
rect 1686 833 2228 868
rect 2719 811 2728 845
rect 2762 811 2800 845
rect 151 728 185 762
rect 2719 758 2753 811
rect 2985 758 3019 907
rect 3497 857 3537 1078
rect 3297 845 3537 857
rect 3331 811 3369 845
rect 3403 811 3441 845
rect 3475 811 3537 845
rect 3297 758 3331 811
rect 3571 796 3605 812
rect 151 660 185 694
rect 3571 728 3605 762
rect 303 651 341 685
rect 581 651 619 685
rect 855 651 893 685
rect 1158 651 1196 685
rect 1471 651 1509 685
rect 1745 651 1783 685
rect 2095 651 2133 685
rect 2457 636 2495 670
rect 2863 653 2901 687
rect 3140 653 3178 687
rect 3415 653 3453 687
rect 3571 660 3605 694
rect 151 592 185 626
rect 3571 592 3605 626
rect 151 524 185 551
rect 1003 513 1037 551
rect 1315 513 1349 551
rect 1627 513 1661 551
rect 1939 513 1973 551
rect 2251 513 2285 551
rect 2563 513 2597 551
rect 3571 524 3605 551
rect 151 456 185 479
rect 151 388 185 422
rect 151 320 185 354
rect 151 252 185 286
rect 151 184 185 218
rect 3571 456 3605 479
rect 3571 388 3605 422
rect 3571 320 3605 354
rect 3571 252 3605 286
rect 425 172 459 216
rect 737 172 771 216
rect 1159 172 1193 216
rect 1471 172 1505 216
rect 2985 172 3019 216
rect 3453 172 3487 216
rect 151 88 185 150
rect 1119 138 1157 172
rect 1191 138 1229 172
rect 1263 138 1301 172
rect 1335 138 1373 172
rect 1407 138 1445 172
rect 1479 138 1517 172
rect 2279 123 2295 157
rect 2329 123 2363 157
rect 2397 123 2413 157
rect 2475 138 2491 172
rect 2525 138 2559 172
rect 2605 138 2627 172
rect 2894 138 2910 172
rect 2944 138 2978 172
rect 3012 138 3046 172
rect 3080 138 3096 172
rect 3206 138 3222 172
rect 3256 138 3290 172
rect 3324 138 3358 172
rect 3392 138 3487 172
rect 3571 184 3605 218
rect 3571 88 3605 150
rect 151 72 3605 88
rect 151 38 193 72
rect 227 38 261 72
rect 295 38 329 72
rect 363 38 397 72
rect 431 38 465 72
rect 499 38 533 72
rect 567 38 601 72
rect 635 38 669 72
rect 703 38 737 72
rect 771 38 805 72
rect 839 38 873 72
rect 907 38 941 72
rect 975 38 1009 72
rect 1043 38 1077 72
rect 1111 38 1145 72
rect 1179 38 1213 72
rect 1247 38 1281 72
rect 1315 38 1349 72
rect 1383 38 1417 72
rect 1451 38 1485 72
rect 1519 38 1553 72
rect 1587 38 1621 72
rect 1655 38 1689 72
rect 1723 38 1757 72
rect 1791 38 1825 72
rect 1859 38 1893 72
rect 1927 38 1961 72
rect 1995 38 2029 72
rect 2063 38 2097 72
rect 2131 38 2165 72
rect 2199 38 2233 72
rect 2267 38 2301 72
rect 2335 38 2369 72
rect 2403 38 2437 72
rect 2471 38 2505 72
rect 2539 38 2573 72
rect 2607 38 2641 72
rect 2675 38 2709 72
rect 2743 38 2777 72
rect 2811 38 2845 72
rect 2879 38 2913 72
rect 2947 38 2981 72
rect 3015 38 3049 72
rect 3083 38 3117 72
rect 3151 38 3185 72
rect 3219 38 3253 72
rect 3287 38 3321 72
rect 3355 38 3389 72
rect 3423 38 3457 72
rect 3491 38 3525 72
rect 3559 38 3605 72
<< viali >>
rect 305 2153 339 2187
rect 377 2153 411 2187
rect 105 2073 139 2107
rect 105 2001 139 2035
rect 261 2045 295 2079
rect 261 1973 295 2007
rect 184 1748 218 1749
rect 184 1715 218 1748
rect 256 1715 290 1749
rect 105 1561 139 1595
rect 105 1489 139 1523
rect 105 1417 139 1451
rect 729 2113 763 2147
rect 729 2041 763 2075
rect 495 1952 529 1986
rect 495 1880 529 1914
rect 589 1902 623 1936
rect 661 1902 695 1936
rect 556 1730 590 1764
rect 628 1730 662 1764
rect 438 1561 472 1595
rect 438 1489 472 1523
rect 438 1417 472 1451
rect 870 1511 904 1545
rect 870 1439 904 1473
rect 2444 1939 2478 1973
rect 2516 1939 2550 1973
rect 2204 1785 2238 1819
rect 2276 1785 2310 1819
rect 1641 1641 1675 1675
rect 1713 1641 1747 1675
rect 1785 1641 1819 1675
rect 1857 1641 1891 1675
rect 1929 1641 1963 1675
rect 2001 1641 2035 1675
rect 2073 1641 2107 1675
rect 1302 1511 1336 1545
rect 1302 1439 1336 1473
rect 1734 1561 1768 1595
rect 1734 1489 1768 1523
rect 1734 1417 1768 1451
rect 2094 1417 2200 1595
rect 654 1347 688 1381
rect 726 1347 760 1381
rect 1098 1337 1132 1371
rect 1170 1337 1204 1371
rect 1484 1337 1518 1371
rect 1556 1337 1590 1371
rect 1878 1337 1912 1371
rect 1950 1337 1984 1371
rect 456 1262 460 1296
rect 460 1262 490 1296
rect 528 1262 562 1296
rect 636 1279 670 1296
rect 708 1279 738 1296
rect 738 1279 742 1296
rect 636 1262 670 1279
rect 708 1262 742 1279
rect 812 1262 846 1296
rect 884 1262 914 1296
rect 914 1262 918 1296
rect 1098 1262 1132 1296
rect 1170 1262 1204 1296
rect 2542 1561 2576 1595
rect 2542 1489 2576 1523
rect 2542 1417 2576 1451
rect 2854 1561 2888 1595
rect 2854 1489 2888 1523
rect 2854 1417 2888 1451
rect 3213 1561 3247 1595
rect 3213 1489 3247 1523
rect 3213 1417 3247 1451
rect 3525 1561 3559 1595
rect 3525 1489 3559 1523
rect 3525 1417 3559 1451
rect 2663 1137 2697 1171
rect 2735 1137 2769 1171
rect 2938 1137 2972 1171
rect 3010 1137 3044 1171
rect 3213 1162 3217 1177
rect 3217 1162 3247 1177
rect 3285 1162 3319 1177
rect 3213 1143 3247 1162
rect 3285 1143 3319 1162
rect 438 1035 472 1069
rect 1868 1035 1902 1069
rect 438 963 472 997
rect 438 891 472 925
rect 1868 963 1902 997
rect 3453 1162 3487 1177
rect 3525 1162 3555 1177
rect 3555 1162 3559 1177
rect 3453 1143 3487 1162
rect 3525 1143 3559 1162
rect 219 811 253 845
rect 291 811 325 845
rect 363 811 397 845
rect 1067 811 1101 845
rect 1139 811 1173 845
rect 2728 811 2762 845
rect 2800 811 2834 845
rect 3297 811 3331 845
rect 3369 811 3403 845
rect 3441 811 3475 845
rect 269 651 303 685
rect 341 651 375 685
rect 547 651 581 685
rect 619 651 653 685
rect 821 651 855 685
rect 893 651 927 685
rect 1124 651 1158 685
rect 1196 651 1230 685
rect 1437 651 1471 685
rect 1509 651 1543 685
rect 1711 651 1745 685
rect 1783 651 1817 685
rect 2061 651 2095 685
rect 2133 651 2167 685
rect 2423 636 2457 670
rect 2495 636 2529 670
rect 2829 653 2863 687
rect 2901 653 2935 687
rect 3106 653 3140 687
rect 3178 653 3212 687
rect 3381 653 3415 687
rect 3453 653 3487 687
rect 151 558 185 585
rect 151 551 185 558
rect 151 490 185 513
rect 151 479 185 490
rect 1003 551 1037 585
rect 1003 479 1037 513
rect 1315 551 1349 585
rect 1315 479 1349 513
rect 1627 551 1661 585
rect 1627 479 1661 513
rect 1939 551 1973 585
rect 1939 479 1973 513
rect 2251 551 2285 585
rect 2251 479 2285 513
rect 2563 551 2597 585
rect 2563 479 2597 513
rect 3571 558 3605 585
rect 3571 551 3605 558
rect 3571 490 3605 513
rect 3571 479 3605 490
rect 1085 138 1119 172
rect 1157 138 1191 172
rect 1229 138 1263 172
rect 1301 138 1335 172
rect 1373 138 1407 172
rect 1445 138 1479 172
rect 1517 138 1551 172
rect 2571 138 2593 172
rect 2593 138 2605 172
rect 2643 138 2661 172
rect 2661 138 2677 172
<< metal1 >>
rect 0 2187 3633 2265
rect 0 2153 305 2187
rect 339 2153 377 2187
rect 411 2153 3633 2187
rect 0 2147 3633 2153
rect 0 2119 729 2147
tri 74 2113 80 2119 ne
rect 80 2113 164 2119
tri 164 2113 170 2119 nw
tri 698 2113 704 2119 ne
rect 704 2113 729 2119
rect 763 2119 3633 2147
rect 763 2113 769 2119
tri 80 2107 86 2113 ne
rect 86 2107 145 2113
tri 86 2094 99 2107 ne
rect 99 2073 105 2107
rect 139 2073 145 2107
tri 145 2094 164 2113 nw
tri 704 2094 723 2113 ne
rect 99 2035 145 2073
rect 99 2001 105 2035
rect 139 2001 145 2035
rect 99 1989 145 2001
rect 255 2079 505 2091
rect 255 2045 261 2079
rect 295 2045 505 2079
rect 255 2039 505 2045
rect 557 2039 569 2091
rect 621 2039 627 2091
rect 723 2075 769 2113
tri 769 2094 794 2119 nw
rect 723 2041 729 2075
rect 763 2041 769 2075
rect 255 2029 321 2039
tri 321 2029 331 2039 nw
rect 723 2029 769 2041
rect 829 2039 835 2091
rect 887 2039 899 2091
rect 951 2063 3633 2091
rect 951 2039 957 2063
tri 957 2039 981 2063 nw
tri 2396 2029 2402 2035 se
rect 2402 2029 3633 2035
rect 255 2007 301 2029
tri 301 2009 321 2029 nw
tri 2376 2009 2396 2029 se
rect 2396 2009 3633 2029
rect 255 1973 261 2007
rect 295 1973 301 2007
tri 2365 1998 2376 2009 se
rect 2376 2007 3633 2009
rect 2376 1998 2410 2007
tri 2410 1998 2419 2007 nw
rect 255 1961 301 1973
rect 489 1986 2391 1998
rect 489 1952 495 1986
rect 529 1979 2391 1986
tri 2391 1979 2410 1998 nw
rect 529 1973 2385 1979
tri 2385 1973 2391 1979 nw
rect 2432 1973 2595 1979
rect 2597 1978 2633 1979
rect 529 1970 2382 1973
tri 2382 1970 2385 1973 nw
rect 529 1952 537 1970
rect 489 1942 537 1952
tri 537 1942 565 1970 nw
rect 489 1914 535 1942
tri 535 1940 537 1942 nw
rect 489 1880 495 1914
rect 529 1880 535 1914
rect 577 1939 2239 1942
tri 2239 1939 2242 1942 sw
rect 2432 1939 2444 1973
rect 2478 1939 2516 1973
rect 2550 1939 2595 1973
rect 577 1936 2242 1939
rect 577 1902 589 1936
rect 623 1902 661 1936
rect 695 1933 2242 1936
tri 2242 1933 2248 1939 sw
rect 695 1927 2248 1933
tri 2248 1927 2254 1933 sw
rect 2432 1927 2595 1939
rect 2596 1928 2634 1978
rect 2597 1927 2633 1928
rect 2635 1927 2658 1979
rect 2710 1927 2722 1979
rect 2774 1927 2780 1979
rect 695 1902 2254 1927
rect 577 1899 2254 1902
tri 2254 1899 2282 1927 sw
rect 577 1896 2589 1899
rect 489 1868 535 1880
tri 2219 1868 2247 1896 ne
rect 2247 1868 2589 1896
tri 2247 1853 2262 1868 ne
rect 2262 1853 2589 1868
rect 2837 1853 2889 1899
tri 2817 1852 2818 1853 ne
rect 2818 1852 2889 1853
rect 622 1846 674 1852
tri 612 1785 622 1795 se
rect 622 1785 674 1794
tri 597 1770 612 1785 se
rect 612 1782 674 1785
rect 612 1770 622 1782
tri 433 1764 439 1770 se
rect 439 1764 622 1770
tri 424 1755 433 1764 se
rect 433 1755 556 1764
rect 172 1749 556 1755
rect 172 1715 184 1749
rect 218 1715 256 1749
rect 290 1730 556 1749
rect 590 1730 622 1764
rect 290 1724 674 1730
rect 702 1800 708 1852
rect 760 1800 772 1852
rect 824 1833 947 1852
tri 947 1833 966 1852 sw
tri 2818 1833 2837 1852 ne
rect 2837 1833 2889 1852
tri 2889 1833 2909 1853 nw
rect 824 1831 966 1833
tri 966 1831 968 1833 sw
rect 2838 1831 2888 1832
rect 824 1825 968 1831
tri 968 1825 974 1831 sw
rect 824 1819 2486 1825
rect 824 1800 2204 1819
rect 702 1785 758 1800
tri 758 1785 773 1800 nw
tri 925 1785 940 1800 ne
rect 940 1785 2204 1800
rect 2238 1785 2276 1819
rect 2310 1795 2486 1819
tri 2486 1795 2516 1825 sw
rect 2310 1785 2516 1795
rect 702 1779 752 1785
tri 752 1779 758 1785 nw
tri 940 1779 946 1785 ne
rect 946 1779 2516 1785
tri 2516 1779 2532 1795 sw
rect 2838 1794 2888 1795
tri 2823 1779 2837 1793 se
rect 2837 1779 2889 1793
rect 702 1753 748 1779
tri 748 1775 752 1779 nw
tri 946 1775 950 1779 ne
rect 950 1775 2532 1779
tri 950 1773 952 1775 ne
rect 952 1773 2532 1775
tri 2532 1773 2538 1779 sw
tri 2817 1773 2823 1779 se
rect 2823 1773 2889 1779
tri 2889 1773 2909 1793 sw
tri 2464 1753 2484 1773 ne
rect 2484 1753 3133 1773
tri 2484 1752 2485 1753 ne
rect 2485 1752 3133 1753
rect 703 1751 747 1752
tri 2485 1751 2486 1752 ne
rect 2486 1751 3133 1752
rect 290 1715 444 1724
rect 172 1709 444 1715
tri 444 1709 459 1724 nw
rect 702 1715 748 1751
tri 2486 1721 2516 1751 ne
rect 2516 1721 3133 1751
rect 703 1714 747 1715
rect 702 1681 748 1713
tri 748 1681 773 1706 sw
rect 702 1675 3633 1681
rect 702 1641 1641 1675
rect 1675 1641 1713 1675
rect 1747 1641 1785 1675
rect 1819 1641 1857 1675
rect 1891 1641 1929 1675
rect 1963 1641 2001 1675
rect 2035 1641 2073 1675
rect 2107 1641 3633 1675
rect 702 1635 3633 1641
rect 0 1595 3633 1607
rect 0 1561 105 1595
rect 139 1561 438 1595
rect 472 1561 1734 1595
rect 1768 1561 2094 1595
rect 0 1545 2094 1561
rect 0 1523 870 1545
rect 0 1489 105 1523
rect 139 1489 438 1523
rect 472 1511 870 1523
rect 904 1511 1302 1545
rect 1336 1523 2094 1545
rect 1336 1511 1734 1523
rect 472 1489 1734 1511
rect 1768 1489 2094 1523
rect 0 1473 2094 1489
rect 0 1451 870 1473
rect 0 1417 105 1451
rect 139 1417 438 1451
rect 472 1441 870 1451
rect 472 1439 648 1441
tri 648 1439 650 1441 nw
tri 764 1439 766 1441 ne
rect 766 1439 870 1441
rect 904 1439 1302 1473
rect 1336 1451 2094 1473
rect 1336 1439 1734 1451
rect 472 1427 636 1439
tri 636 1427 648 1439 nw
tri 766 1427 778 1439 ne
rect 778 1427 1734 1439
rect 472 1417 626 1427
tri 626 1417 636 1427 nw
tri 778 1417 788 1427 ne
rect 788 1417 1734 1427
rect 1768 1417 2094 1451
rect 2200 1561 2542 1595
rect 2576 1561 2854 1595
rect 2888 1561 3213 1595
rect 3247 1561 3525 1595
rect 3559 1561 3633 1595
rect 2200 1523 3633 1561
rect 2200 1489 2542 1523
rect 2576 1489 2854 1523
rect 2888 1489 3213 1523
rect 3247 1489 3525 1523
rect 3559 1489 3633 1523
rect 2200 1451 3633 1489
rect 2200 1417 2542 1451
rect 2576 1417 2854 1451
rect 2888 1417 3213 1451
rect 3247 1417 3525 1451
rect 3559 1417 3633 1451
rect 0 1405 614 1417
tri 614 1405 626 1417 nw
tri 788 1405 800 1417 ne
rect 800 1405 3633 1417
rect 642 1381 772 1387
rect 642 1347 654 1381
rect 688 1347 726 1381
rect 760 1377 772 1381
tri 772 1377 782 1387 sw
rect 760 1371 1408 1377
rect 1410 1376 1446 1377
rect 760 1347 1098 1371
rect 642 1341 1098 1347
tri 752 1337 756 1341 ne
rect 756 1337 1098 1341
rect 1132 1337 1170 1371
rect 1204 1337 1408 1371
tri 756 1331 762 1337 ne
rect 762 1331 1408 1337
rect 1409 1332 1447 1376
rect 1448 1371 1996 1377
rect 1448 1337 1484 1371
rect 1518 1337 1556 1371
rect 1590 1337 1878 1371
rect 1912 1337 1950 1371
rect 1984 1337 1996 1371
rect 1410 1331 1446 1332
rect 1448 1331 1996 1337
rect 444 1296 574 1303
rect 444 1262 456 1296
rect 490 1262 528 1296
rect 562 1262 574 1296
rect 444 1251 574 1262
rect 575 1252 576 1302
rect 612 1252 613 1302
rect 614 1251 632 1303
rect 684 1251 696 1303
rect 748 1251 754 1303
rect 800 1251 810 1303
rect 862 1251 874 1303
rect 926 1251 932 1303
rect 960 1251 966 1303
rect 1018 1251 1030 1303
rect 1082 1296 2483 1303
rect 1082 1262 1098 1296
rect 1132 1262 1170 1296
rect 1204 1262 2483 1296
rect 1082 1251 2483 1262
rect 2535 1251 2547 1303
rect 2599 1251 3633 1303
rect 499 1131 505 1183
rect 557 1131 569 1183
rect 621 1131 2658 1183
rect 2710 1131 2722 1183
rect 2774 1177 3571 1183
rect 2774 1171 3213 1177
rect 2774 1137 2938 1171
rect 2972 1137 3010 1171
rect 3044 1143 3213 1171
rect 3247 1143 3285 1177
rect 3319 1143 3453 1177
rect 3487 1143 3525 1177
rect 3559 1143 3571 1177
rect 3044 1137 3571 1143
rect 2774 1131 3571 1137
rect 0 1071 3633 1081
rect 0 1069 2713 1071
rect 0 1035 438 1069
rect 472 1035 1868 1069
rect 1902 1035 2713 1069
rect 0 1019 2713 1035
rect 2765 1019 3633 1071
rect 0 1007 3633 1019
rect 0 997 2713 1007
rect 0 963 438 997
rect 472 963 1868 997
rect 1902 963 2713 997
rect 0 955 2713 963
rect 2765 955 3633 1007
rect 0 943 3633 955
rect 0 925 2713 943
rect 0 891 438 925
rect 472 891 2713 925
rect 2765 891 3633 943
rect 0 879 3633 891
rect 207 845 538 851
tri 538 845 544 851 sw
rect 207 811 219 845
rect 253 811 291 845
rect 325 811 363 845
rect 397 811 544 845
tri 544 811 578 845 sw
rect 207 805 578 811
tri 578 805 584 811 sw
rect 207 799 584 805
tri 584 799 590 805 sw
rect 884 799 890 851
rect 942 799 954 851
rect 1006 799 1013 851
rect 1015 850 1051 851
rect 1014 800 1052 850
rect 1053 845 1189 851
rect 1053 811 1067 845
rect 1101 811 1139 845
rect 1173 811 1189 845
rect 1015 799 1051 800
rect 1053 799 1189 811
rect 1675 845 3487 851
rect 1675 811 2728 845
rect 2762 811 2800 845
rect 2834 811 3297 845
rect 3331 811 3369 845
rect 3403 811 3441 845
rect 3475 811 3487 845
rect 1675 805 3487 811
tri 516 771 544 799 ne
rect 544 771 590 799
tri 590 771 618 799 sw
tri 544 719 596 771 ne
rect 596 765 2685 771
rect 596 719 2633 765
tri 2608 694 2633 719 ne
rect 2633 701 2685 713
rect 257 685 1607 691
rect 1609 690 1645 691
rect 257 651 269 685
rect 303 651 341 685
rect 375 651 547 685
rect 581 651 619 685
rect 653 651 821 685
rect 855 651 893 685
rect 927 651 1124 685
rect 1158 651 1196 685
rect 1230 651 1437 685
rect 1471 651 1509 685
rect 1543 651 1607 685
rect 257 645 1607 651
rect 1608 646 1646 690
rect 1647 685 2179 691
rect 1647 651 1711 685
rect 1745 651 1783 685
rect 1817 651 2061 685
rect 2095 651 2133 685
rect 2167 651 2179 685
rect 1609 645 1645 646
rect 1647 645 2179 651
rect 2411 670 2483 682
rect 2411 636 2423 670
rect 2457 636 2483 670
rect 2411 630 2483 636
rect 2535 630 2547 682
rect 2599 630 2605 682
rect 2633 643 2685 649
rect 2817 687 3499 693
rect 2817 653 2829 687
rect 2863 653 2901 687
rect 2935 653 3106 687
rect 3140 653 3178 687
rect 3212 653 3381 687
rect 3415 653 3453 687
rect 3487 653 3499 687
rect 2817 647 3499 653
rect 0 591 3633 597
rect 0 585 2713 591
rect 0 551 151 585
rect 185 551 1003 585
rect 1037 551 1315 585
rect 1349 551 1627 585
rect 1661 551 1939 585
rect 1973 551 2251 585
rect 2285 551 2563 585
rect 2597 551 2713 585
rect 0 539 2713 551
rect 2765 585 3633 591
rect 2765 551 3571 585
rect 3605 551 3633 585
rect 2765 539 3633 551
rect 0 527 3633 539
rect 0 513 2713 527
rect 0 479 151 513
rect 185 479 1003 513
rect 1037 479 1315 513
rect 1349 479 1627 513
rect 1661 479 1939 513
rect 1973 479 2251 513
rect 2285 479 2563 513
rect 2597 479 2713 513
rect 0 475 2713 479
rect 2765 513 3633 527
rect 2765 479 3571 513
rect 3605 479 3633 513
rect 2765 475 3633 479
rect 0 467 3633 475
rect 378 126 890 178
rect 942 126 954 178
rect 1006 126 1013 178
rect 1014 127 1015 177
rect 1046 177 1051 178
rect 1046 127 1052 177
rect 1053 172 1604 178
rect 1053 138 1085 172
rect 1119 138 1157 172
rect 1191 138 1229 172
rect 1263 138 1301 172
rect 1335 138 1373 172
rect 1407 138 1445 172
rect 1479 138 1517 172
rect 1551 138 1604 172
rect 1046 126 1051 127
rect 1053 126 1604 138
rect 2559 172 2639 186
rect 2559 138 2571 172
rect 2605 138 2639 172
rect 2559 134 2639 138
rect 2691 134 2703 186
rect 2755 134 2763 186
rect 2559 132 2763 134
<< rmetal1 >>
rect 2595 1978 2597 1979
rect 2633 1978 2635 1979
rect 2595 1928 2596 1978
rect 2634 1928 2635 1978
rect 2595 1927 2597 1928
rect 2633 1927 2635 1928
rect 2837 1832 2889 1833
rect 2837 1831 2838 1832
rect 2888 1831 2889 1832
rect 2837 1794 2838 1795
rect 2888 1794 2889 1795
rect 2837 1793 2889 1794
rect 702 1752 748 1753
rect 702 1751 703 1752
rect 747 1751 748 1752
rect 702 1714 703 1715
rect 747 1714 748 1715
rect 702 1713 748 1714
rect 1408 1376 1410 1377
rect 1446 1376 1448 1377
rect 1408 1332 1409 1376
rect 1447 1332 1448 1376
rect 1408 1331 1410 1332
rect 1446 1331 1448 1332
rect 574 1302 576 1303
rect 574 1252 575 1302
rect 574 1251 576 1252
rect 612 1302 614 1303
rect 613 1252 614 1302
rect 612 1251 614 1252
rect 1013 850 1015 851
rect 1051 850 1053 851
rect 1013 800 1014 850
rect 1052 800 1053 850
rect 1013 799 1015 800
rect 1051 799 1053 800
rect 1607 690 1609 691
rect 1645 690 1647 691
rect 1607 646 1608 690
rect 1646 646 1647 690
rect 1607 645 1609 646
rect 1645 645 1647 646
rect 1013 177 1015 178
rect 1013 127 1014 177
rect 1013 126 1015 127
rect 1051 177 1053 178
rect 1052 127 1053 177
rect 1051 126 1053 127
<< via1 >>
rect 505 2039 557 2091
rect 569 2039 621 2091
rect 835 2039 887 2091
rect 899 2039 951 2091
rect 2658 1927 2710 1979
rect 2722 1927 2774 1979
rect 622 1794 674 1846
rect 622 1764 674 1782
rect 622 1730 628 1764
rect 628 1730 662 1764
rect 662 1730 674 1764
rect 708 1800 760 1852
rect 772 1800 824 1852
rect 632 1296 684 1303
rect 632 1262 636 1296
rect 636 1262 670 1296
rect 670 1262 684 1296
rect 632 1251 684 1262
rect 696 1296 748 1303
rect 696 1262 708 1296
rect 708 1262 742 1296
rect 742 1262 748 1296
rect 696 1251 748 1262
rect 810 1296 862 1303
rect 810 1262 812 1296
rect 812 1262 846 1296
rect 846 1262 862 1296
rect 810 1251 862 1262
rect 874 1296 926 1303
rect 874 1262 884 1296
rect 884 1262 918 1296
rect 918 1262 926 1296
rect 874 1251 926 1262
rect 966 1251 1018 1303
rect 1030 1251 1082 1303
rect 2483 1251 2535 1303
rect 2547 1251 2599 1303
rect 505 1131 557 1183
rect 569 1131 621 1183
rect 2658 1171 2710 1183
rect 2658 1137 2663 1171
rect 2663 1137 2697 1171
rect 2697 1137 2710 1171
rect 2658 1131 2710 1137
rect 2722 1171 2774 1183
rect 2722 1137 2735 1171
rect 2735 1137 2769 1171
rect 2769 1137 2774 1171
rect 2722 1131 2774 1137
rect 2713 1019 2765 1071
rect 2713 955 2765 1007
rect 2713 891 2765 943
rect 890 799 942 851
rect 954 799 1006 851
rect 2633 713 2685 765
rect 2483 670 2535 682
rect 2483 636 2495 670
rect 2495 636 2529 670
rect 2529 636 2535 670
rect 2483 630 2535 636
rect 2547 630 2599 682
rect 2633 649 2685 701
rect 2713 539 2765 591
rect 2713 475 2765 527
rect 890 126 942 178
rect 954 126 1006 178
rect 2639 172 2691 186
rect 2639 138 2643 172
rect 2643 138 2677 172
rect 2677 138 2691 172
rect 2639 134 2691 138
rect 2703 134 2755 186
<< metal2 >>
rect 499 2039 505 2091
rect 557 2039 569 2091
rect 621 2039 627 2091
rect 829 2039 835 2091
rect 887 2039 899 2091
rect 951 2039 957 2091
rect 499 1183 563 2039
tri 563 2014 588 2039 nw
tri 855 2014 880 2039 ne
tri 855 1941 880 1966 se
rect 880 1941 932 2039
tri 932 2014 957 2039 nw
rect 622 1889 932 1941
rect 622 1846 674 1889
tri 674 1864 699 1889 nw
tri 855 1864 880 1889 ne
rect 622 1782 674 1794
rect 622 1724 674 1730
rect 702 1800 708 1852
rect 760 1800 772 1852
rect 824 1800 830 1852
tri 677 1303 702 1328 se
rect 702 1303 754 1800
tri 754 1775 779 1800 nw
tri 855 1303 880 1328 se
rect 880 1303 932 1889
rect 2652 1927 2658 1979
rect 2710 1927 2722 1979
rect 2774 1927 2780 1979
rect 626 1251 632 1303
rect 684 1251 696 1303
rect 748 1251 754 1303
rect 804 1251 810 1303
rect 862 1251 874 1303
rect 926 1251 932 1303
rect 960 1251 966 1303
rect 1018 1251 1030 1303
rect 1082 1251 1088 1303
rect 2477 1251 2483 1303
rect 2535 1251 2547 1303
rect 2599 1251 2605 1303
tri 563 1183 588 1208 sw
rect 499 1131 505 1183
rect 557 1131 569 1183
rect 621 1131 627 1183
tri 935 851 960 876 se
rect 960 851 1012 1251
tri 1012 1226 1037 1251 nw
tri 2528 1226 2553 1251 ne
rect 884 799 890 851
rect 942 799 954 851
rect 1006 799 1012 851
tri 935 774 960 799 ne
tri 943 186 960 203 se
rect 960 186 1012 799
tri 2547 701 2553 707 se
rect 2553 701 2605 1251
rect 2652 1183 2704 1927
tri 2704 1902 2729 1927 nw
tri 2704 1183 2729 1208 sw
rect 2652 1131 2658 1183
rect 2710 1131 2722 1183
rect 2774 1131 2780 1183
rect 2713 1071 2765 1081
rect 2713 1007 2765 1019
rect 2713 943 2765 955
tri 2528 682 2547 701 se
rect 2547 682 2605 701
rect 2477 630 2483 682
rect 2535 630 2547 682
rect 2599 630 2605 682
rect 2633 765 2685 771
rect 2633 701 2685 713
tri 935 178 943 186 se
rect 943 178 1012 186
rect 884 126 890 178
rect 942 126 954 178
rect 1006 126 1012 178
rect 2633 186 2685 649
rect 2713 591 2765 891
rect 2713 527 2765 539
rect 2713 469 2765 475
tri 2685 186 2710 211 sw
rect 2633 134 2639 186
rect 2691 134 2703 186
rect 2755 134 2761 186
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1701704242
transform 0 -1 1902 -1 0 1069
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1701704242
transform 0 -1 529 -1 0 1986
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1701704242
transform 0 1 729 -1 0 2147
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_3
timestamp 1701704242
transform 0 1 105 -1 0 2107
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_4
timestamp 1701704242
transform -1 0 1984 0 1 1337
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_5
timestamp 1701704242
transform -1 0 562 0 1 1262
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_6
timestamp 1701704242
transform -1 0 2310 0 1 1785
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_7
timestamp 1701704242
transform -1 0 3044 0 1 1137
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_8
timestamp 1701704242
transform -1 0 2769 0 1 1137
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_9
timestamp 1701704242
transform -1 0 1590 0 1 1337
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_10
timestamp 1701704242
transform -1 0 2550 0 -1 1973
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_11
timestamp 1701704242
transform -1 0 2529 0 -1 670
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_12
timestamp 1701704242
transform 0 1 2563 1 0 479
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_13
timestamp 1701704242
transform 0 1 1315 1 0 479
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_14
timestamp 1701704242
transform 0 1 1939 1 0 479
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_15
timestamp 1701704242
transform 0 1 1627 1 0 479
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_16
timestamp 1701704242
transform 0 1 2251 1 0 479
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_17
timestamp 1701704242
transform 0 1 1003 1 0 479
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_18
timestamp 1701704242
transform 0 1 3571 1 0 479
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_19
timestamp 1701704242
transform 0 1 151 1 0 479
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_20
timestamp 1701704242
transform 0 -1 904 1 0 1439
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_21
timestamp 1701704242
transform 0 -1 1336 1 0 1439
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_22
timestamp 1701704242
transform 0 -1 295 1 0 1973
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_23
timestamp 1701704242
transform 1 0 2061 0 -1 685
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_24
timestamp 1701704242
transform 1 0 1124 0 -1 685
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_25
timestamp 1701704242
transform 1 0 1437 0 -1 685
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_26
timestamp 1701704242
transform 1 0 1067 0 -1 845
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_27
timestamp 1701704242
transform 1 0 3213 0 -1 1177
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_28
timestamp 1701704242
transform 1 0 1711 0 -1 685
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_29
timestamp 1701704242
transform 1 0 2829 0 -1 687
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_30
timestamp 1701704242
transform 1 0 3381 0 -1 687
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_31
timestamp 1701704242
transform 1 0 269 0 -1 685
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_32
timestamp 1701704242
transform 1 0 821 0 -1 685
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_33
timestamp 1701704242
transform 1 0 3453 0 -1 1177
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_34
timestamp 1701704242
transform 1 0 3106 0 -1 687
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_35
timestamp 1701704242
transform 1 0 1098 0 -1 1371
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_36
timestamp 1701704242
transform 1 0 1098 0 -1 1296
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_37
timestamp 1701704242
transform 1 0 547 0 -1 685
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_38
timestamp 1701704242
transform 1 0 2728 0 -1 845
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_39
timestamp 1701704242
transform 1 0 654 0 -1 1381
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_40
timestamp 1701704242
transform 1 0 305 0 1 2153
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_41
timestamp 1701704242
transform 1 0 812 0 1 1262
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_42
timestamp 1701704242
transform 1 0 636 0 1 1262
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_43
timestamp 1701704242
transform 1 0 589 0 1 1902
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_44
timestamp 1701704242
transform 1 0 2571 0 1 138
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_45
timestamp 1701704242
transform 1 0 184 0 1 1715
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_46
timestamp 1701704242
transform 1 0 556 0 1 1730
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_0
timestamp 1701704242
transform 0 -1 1768 -1 0 1595
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_1
timestamp 1701704242
transform 0 -1 472 -1 0 1069
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_2
timestamp 1701704242
transform 0 -1 2576 -1 0 1595
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_3
timestamp 1701704242
transform 0 -1 2888 -1 0 1595
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_4
timestamp 1701704242
transform 0 -1 3247 -1 0 1595
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_5
timestamp 1701704242
transform 0 -1 3559 -1 0 1595
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_6
timestamp 1701704242
transform -1 0 397 0 1 811
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_7
timestamp 1701704242
transform -1 0 3475 0 -1 845
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_8
timestamp 1701704242
transform 0 -1 139 1 0 1417
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_9
timestamp 1701704242
transform 0 -1 472 1 0 1417
box 0 0 1 1
use L1M1_CDNS_52468879185195  L1M1_CDNS_52468879185195_0
timestamp 1701704242
transform -1 0 3137 0 1 1859
box -12 -6 550 40
use L1M1_CDNS_52468879185195  L1M1_CDNS_52468879185195_1
timestamp 1701704242
transform -1 0 928 0 -1 172
box -12 -6 550 40
use L1M1_CDNS_52468879185195  L1M1_CDNS_52468879185195_2
timestamp 1701704242
transform 1 0 1687 0 -1 845
box -12 -6 550 40
use L1M1_CDNS_52468879185334  L1M1_CDNS_52468879185334_0
timestamp 1701704242
transform 0 1 2094 -1 0 1595
box 0 0 1 1
use L1M1_CDNS_52468879185337  L1M1_CDNS_52468879185337_0
timestamp 1701704242
transform -1 0 2107 0 1 1641
box 0 0 1 1
use L1M1_CDNS_52468879185337  L1M1_CDNS_52468879185337_1
timestamp 1701704242
transform 1 0 1085 0 -1 172
box 0 0 1 1
use L1M1_CDNS_52468879185381  L1M1_CDNS_52468879185381_0
timestamp 1701704242
transform -1 0 1800 0 -1 1175
box -12 -6 910 40
use L1M1_CDNS_52468879185382  L1M1_CDNS_52468879185382_0
timestamp 1701704242
transform -1 0 3101 0 1 2225
box -12 -6 2998 40
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_0
timestamp 1701704242
transform 0 -1 2685 -1 0 771
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_1
timestamp 1701704242
transform -1 0 2605 0 1 630
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_2
timestamp 1701704242
transform -1 0 754 0 1 1251
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_3
timestamp 1701704242
transform -1 0 2780 0 1 1927
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_4
timestamp 1701704242
transform -1 0 1088 0 1 1251
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_5
timestamp 1701704242
transform -1 0 1012 0 1 799
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_6
timestamp 1701704242
transform -1 0 957 0 1 2039
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_7
timestamp 1701704242
transform 0 1 622 1 0 1724
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_8
timestamp 1701704242
transform 0 -1 2765 1 0 469
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_9
timestamp 1701704242
transform 1 0 804 0 -1 1303
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_10
timestamp 1701704242
transform 1 0 702 0 -1 1852
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_11
timestamp 1701704242
transform 1 0 499 0 -1 2091
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_12
timestamp 1701704242
transform 1 0 884 0 -1 178
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_13
timestamp 1701704242
transform 1 0 2633 0 -1 186
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_14
timestamp 1701704242
transform 1 0 499 0 1 1131
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_15
timestamp 1701704242
transform 1 0 2477 0 1 1251
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_16
timestamp 1701704242
transform 1 0 2652 0 1 1131
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_0
timestamp 1701704242
transform 0 -1 2765 -1 0 1077
box 0 0 1 1
use nfet_CDNS_52468879185344  nfet_CDNS_52468879185344_0
timestamp 1701704242
transform -1 0 2396 0 1 220
box -79 -26 179 626
use nfet_CDNS_52468879185344  nfet_CDNS_52468879185344_1
timestamp 1701704242
transform 1 0 2608 0 1 220
box -79 -26 179 626
use nfet_CDNS_52468879185344  nfet_CDNS_52468879185344_2
timestamp 1701704242
transform 1 0 2452 0 1 220
box -79 -26 179 626
use nfet_CDNS_52468879185374  nfet_CDNS_52468879185374_0
timestamp 1701704242
transform -1 0 1857 0 -1 1074
box -79 -26 879 110
use nfet_CDNS_52468879185375  nfet_CDNS_52468879185375_0
timestamp 1701704242
transform 1 0 483 0 1 914
box -79 -26 176 326
use nfet_CDNS_52468879185390  nfet_CDNS_52468879185390_0
timestamp 1701704242
transform 1 0 1913 0 -1 1074
box -79 -26 1679 110
use nfet_CDNS_52468879185391  nfet_CDNS_52468879185391_0
timestamp 1701704242
transform -1 0 3442 0 1 220
box -79 -26 335 626
use nfet_CDNS_52468879185392  nfet_CDNS_52468879185392_0
timestamp 1701704242
transform -1 0 1616 0 1 220
box -79 -26 647 626
use nfet_CDNS_52468879185392  nfet_CDNS_52468879185392_1
timestamp 1701704242
transform -1 0 2240 0 1 220
box -79 -26 647 626
use nfet_CDNS_52468879185392  nfet_CDNS_52468879185392_2
timestamp 1701704242
transform -1 0 882 0 1 220
box -79 -26 647 626
use nfet_CDNS_52468879185393  nfet_CDNS_52468879185393_0
timestamp 1701704242
transform 1 0 637 0 1 914
box 0 0 1 1
use nfet_CDNS_52468879185394  nfet_CDNS_52468879185394_0
timestamp 1701704242
transform 1 0 791 0 1 914
box -76 -26 179 326
use nfet_CDNS_52468879185395  nfet_CDNS_52468879185395_0
timestamp 1701704242
transform 1 0 2874 0 1 220
box -79 -26 335 626
use nfet_CDNS_52468879185396  nfet_CDNS_52468879185396_0
timestamp 1701704242
transform -1 0 380 0 1 1014
box -76 -26 199 226
use pfet_CDNS_52468879185367  pfet_CDNS_52468879185367_0
timestamp 1701704242
transform -1 0 2421 0 1 1244
box -119 -66 219 666
use pfet_CDNS_52468879185397  pfet_CDNS_52468879185397_0
timestamp 1701704242
transform 1 0 3258 0 1 1244
box -119 -66 375 1066
use pfet_CDNS_52468879185398  pfet_CDNS_52468879185398_0
timestamp 1701704242
transform -1 0 406 0 1 1898
box -119 -66 219 266
use pfet_CDNS_52468879185398  pfet_CDNS_52468879185398_1
timestamp 1701704242
transform -1 0 718 0 1 1898
box -119 -66 219 266
use pfet_CDNS_52468879185398  pfet_CDNS_52468879185398_2
timestamp 1701704242
transform 1 0 150 0 1 1898
box -119 -66 219 266
use pfet_CDNS_52468879185398  pfet_CDNS_52468879185398_3
timestamp 1701704242
transform 1 0 462 0 1 1898
box -119 -66 219 266
use pfet_CDNS_52468879185399  pfet_CDNS_52468879185399_0
timestamp 1701704242
transform 1 0 483 0 1 1397
box -119 -66 927 266
use pfet_CDNS_52468879185399  pfet_CDNS_52468879185399_1
timestamp 1701704242
transform 1 0 1347 0 1 1397
box -119 -66 927 266
use pfet_CDNS_52468879185400  pfet_CDNS_52468879185400_0
timestamp 1701704242
transform 1 0 2587 0 1 1244
box -119 -66 684 666
use pfet_CDNS_52468879185401  pfet_CDNS_52468879185401_0
timestamp 1701704242
transform 1 0 150 0 1 1397
box -119 -66 372 266
use pfet_CDNS_52468879185402  pfet_CDNS_52468879185402_0
timestamp 1701704242
transform 1 0 821 0 1 2014
box -116 -66 1719 150
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_0
timestamp 1701704242
transform 1 0 2280 0 1 1876
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_0
timestamp 1701704242
transform 0 -1 578 -1 0 1312
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_1
timestamp 1701704242
transform 0 1 796 -1 0 1312
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_2
timestamp 1701704242
transform 0 1 620 -1 0 1329
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_3
timestamp 1701704242
transform 0 1 600 -1 0 1847
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_4
timestamp 1701704242
transform 0 1 3437 1 0 1146
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_5
timestamp 1701704242
transform 0 1 2279 1 0 107
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_6
timestamp 1701704242
transform 0 1 445 1 0 2141
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_7
timestamp 1701704242
transform 0 1 3201 1 0 1146
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_8
timestamp 1701704242
transform 0 -1 1601 1 0 1629
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_9
timestamp 1701704242
transform 1 0 324 0 1 1732
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_0
timestamp 1701704242
transform 0 1 2894 1 0 122
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_1
timestamp 1701704242
transform 0 1 3206 1 0 122
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_2
timestamp 1701704242
transform 0 -1 2677 1 0 122
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_3
timestamp 1701704242
transform 1 0 168 0 -1 1866
box 0 0 1 1
use PYL1_CDNS_52468879185309  PYL1_CDNS_52468879185309_0
timestamp 1701704242
transform 0 1 511 1 0 1629
box 0 0 1 1
use PYL1_CDNS_52468879185309  PYL1_CDNS_52468879185309_1
timestamp 1701704242
transform 0 -1 1236 1 0 1629
box 0 0 1 1
use PYL1_CDNS_52468879185318  PYL1_CDNS_52468879185318_0
timestamp 1701704242
transform 0 1 1686 -1 0 918
box 0 0 66 542
use PYL1_CDNS_52468879185318  PYL1_CDNS_52468879185318_1
timestamp 1701704242
transform 0 1 1062 -1 0 188
box 0 0 66 542
use PYL1_CDNS_52468879185318  PYL1_CDNS_52468879185318_2
timestamp 1701704242
transform 0 1 328 -1 0 188
box 0 0 66 542
use PYL1_CDNS_52468879185318  PYL1_CDNS_52468879185318_3
timestamp 1701704242
transform 0 1 2598 1 0 1876
box 0 0 66 542
use PYL1_CDNS_52468879185318  PYL1_CDNS_52468879185318_4
timestamp 1701704242
transform 0 -1 1820 1 0 1253
box 0 0 66 542
use PYL1_CDNS_52468879185383  PYL1_CDNS_52468879185383_0
timestamp 1701704242
transform 0 1 1966 -1 0 1172
box 0 0 66 610
use PYL1_CDNS_52468879185384  PYL1_CDNS_52468879185384_0
timestamp 1701704242
transform 0 1 825 1 0 1916
box 0 0 66 1358
use PYL1_CDNS_52468879185385  PYL1_CDNS_52468879185385_0
timestamp 1701704242
transform 0 -1 1820 1 0 1106
box 0 0 134 678
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851254  sky130_fd_io__sio_tk_em1o_CDNS_524688791851254_0
timestamp 1701704242
transform -1 0 1105 0 1 126
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851254  sky130_fd_io__sio_tk_em1o_CDNS_524688791851254_1
timestamp 1701704242
transform 1 0 522 0 1 1251
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851420  sky130_fd_io__sio_tk_em1o_CDNS_524688791851420_0
timestamp 1701704242
transform 0 -1 2889 1 0 1741
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851255  sky130_fd_io__sio_tk_em1s_CDNS_524688791851255_0
timestamp 1701704242
transform -1 0 2687 0 1 1927
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851255  sky130_fd_io__sio_tk_em1s_CDNS_524688791851255_1
timestamp 1701704242
transform -1 0 1105 0 1 799
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851295  sky130_fd_io__sio_tk_em1s_CDNS_524688791851295_0
timestamp 1701704242
transform 1 0 1356 0 1 1331
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851295  sky130_fd_io__sio_tk_em1s_CDNS_524688791851295_1
timestamp 1701704242
transform 1 0 1555 0 1 645
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851419  sky130_fd_io__sio_tk_em1s_CDNS_524688791851419_0
timestamp 1701704242
transform 0 -1 748 -1 0 1805
box 0 0 1 1
use TPL1_CDNS_52468879185386  TPL1_CDNS_52468879185386_0
timestamp 1701704242
transform 0 1 867 -1 0 1888
box -36 -36 186 730
use TPL1_CDNS_52468879185387  TPL1_CDNS_52468879185387_0
timestamp 1701704242
transform 0 1 2608 -1 0 2182
box -36 -36 254 526
<< labels >>
flabel comment s 2992 179 2992 179 0 FreeSans 300 0 0 0 n<7>
flabel comment s 3307 179 3307 179 0 FreeSans 300 0 0 0 n<8>
flabel comment s 2215 1686 2215 1686 0 FreeSans 300 180 0 0 pu_h_n
flabel comment s 2043 1291 2043 1291 0 FreeSans 300 0 0 0 nbias
flabel comment s 887 1361 887 1361 0 FreeSans 300 0 0 0 nbias
flabel comment s 776 1151 776 1151 0 FreeSans 300 270 0 0 n<3>
flabel comment s 620 1151 620 1151 0 FreeSans 300 270 0 0 n<4>
flabel comment s 1307 1934 1307 1934 0 FreeSans 300 0 0 0 n<1>
flabel comment s 1305 1800 1305 1800 0 FreeSans 300 180 0 0 n<2>
flabel comment s 2853 920 2853 920 0 FreeSans 300 0 0 0 vgnd_io
flabel comment s 611 1709 611 1709 0 FreeSans 300 90 0 0 n<2>
flabel comment s 203 1352 203 1352 0 FreeSans 300 0 0 0 drvhi_h_n
flabel comment s 429 2046 429 2046 0 FreeSans 300 0 0 0 vccio
flabel comment s 2238 1522 2238 1522 0 FreeSans 300 0 0 0 vccio
flabel comment s 1967 1990 1967 1990 0 FreeSans 300 180 0 0 pu_h_n
flabel comment s 533 190 533 190 0 FreeSans 300 0 0 0 nbias
flabel comment s 1267 190 1267 190 0 FreeSans 300 0 0 0 n<6>
flabel comment s 2341 192 2341 192 0 FreeSans 300 0 0 0 en_h_n
flabel comment s 2587 192 2587 192 0 FreeSans 300 0 0 0 drvhi_h_n
flabel comment s 1891 857 1891 857 0 FreeSans 300 0 0 0 vccio_2vtn
flabel comment s 2755 737 2755 737 0 FreeSans 300 90 0 0 vccio_2vtn
flabel comment s 1883 525 1883 525 0 FreeSans 300 0 0 0 vgnd_io
flabel comment s 3082 677 3082 677 0 FreeSans 300 0 0 0 n<8>
flabel comment s 1881 1032 1881 1032 0 FreeSans 300 270 0 0 vgnd_io
flabel comment s 1423 1201 1423 1201 0 FreeSans 300 0 0 0 bias_g
flabel comment s 2879 1108 2879 1108 0 FreeSans 300 0 0 0 vccio
flabel comment s 1283 1629 1283 1629 0 FreeSans 300 0 0 0 bias_g
flabel comment s 3336 1210 3336 1210 0 FreeSans 300 0 0 0 bias_g
flabel comment s 2353 1940 2353 1940 0 FreeSans 300 0 0 0 n<2>
flabel comment s 2891 1884 2891 1884 0 FreeSans 300 0 0 0 n<1>
flabel comment s 508 1310 508 1310 0 FreeSans 300 0 0 0 en_h
flabel comment s 671 1239 671 1239 0 FreeSans 300 0 0 0 m1 opt en_h
flabel comment s 888 1310 888 1310 0 FreeSans 300 0 0 0 drvhi_h
flabel comment s 361 1870 361 1870 0 FreeSans 300 180 0 0 en_h
flabel comment s 3136 843 3136 843 0 FreeSans 300 0 0 0 vccio_2vtn
flabel comment s 2579 791 2579 791 0 FreeSans 300 90 0 0 nbias
flabel comment s 941 668 941 668 0 FreeSans 300 0 0 0 n<6>
flabel comment s 1970 676 1970 676 0 FreeSans 300 0 0 0 m1 opt n<6>
flabel metal1 s 3593 2119 3633 2265 7 FreeSans 300 180 0 0 vcc_io
port 1 nsew
flabel metal1 s 0 2119 37 2265 6 FreeSans 300 0 0 0 vcc_io
port 1 nsew
flabel metal1 s 702 1635 744 1681 7 FreeSans 300 180 0 0 pu_h_n
port 2 nsew
flabel metal1 s 0 1405 42 1607 6 FreeSans 300 0 0 0 vcc_io
port 1 nsew
flabel metal1 s 0 879 42 1081 7 FreeSans 300 0 0 0 vgnd_io
port 3 nsew
flabel metal1 s 0 467 42 597 7 FreeSans 300 0 0 0 vgnd_io
port 3 nsew
flabel metal1 s 3593 1635 3633 1681 7 FreeSans 300 180 0 0 pu_h_n
port 2 nsew
flabel metal1 s 3593 1405 3633 1607 7 FreeSans 300 180 0 0 vcc_io
port 1 nsew
flabel metal1 s 3591 879 3633 1081 7 FreeSans 300 180 0 0 vgnd_io
port 3 nsew
flabel metal1 s 3593 2007 3633 2035 7 FreeSans 300 180 0 0 puen_h
port 4 nsew
flabel metal1 s 3593 2063 3633 2091 7 FreeSans 300 180 0 0 drvhi_h
port 6 nsew
flabel metal1 s 3593 1251 3633 1303 7 FreeSans 300 180 0 0 nbias
port 5 nsew
flabel metal1 s 3591 467 3633 597 7 FreeSans 300 180 0 0 vgnd_io
port 3 nsew
flabel locali s 340 1795 374 1866 8 FreeSans 300 0 0 0 en_h
port 8 nsew
flabel locali s 2363 123 2413 157 0 FreeSans 300 0 0 0 en_h_n
port 9 nsew
<< properties >>
string GDS_END 87807936
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 87776894
<< end >>
