magic
tech sky130B
timestamp 1701704242
<< metal1 >>
rect 0 0 3 218
rect 157 0 160 218
<< via1 >>
rect 3 0 157 218
<< metal2 >>
rect 0 0 3 218
rect 157 0 160 218
<< properties >>
string GDS_END 85878100
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85875728
<< end >>
