magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< locali >>
rect 36531 4278 36565 4316
rect 40019 4278 40053 4316
rect 40736 4278 40770 4316
rect 44224 4278 44258 4316
<< viali >>
rect 36531 4316 36565 4350
rect 36531 4244 36565 4278
rect 40019 4316 40053 4350
rect 40019 4244 40053 4278
rect 40736 4316 40770 4350
rect 40736 4244 40770 4278
rect 44224 4316 44258 4350
rect 44224 4244 44258 4278
<< metal1 >>
tri 33158 38853 33183 38878 se
rect 33183 38853 34035 38878
rect 33158 38850 34035 38853
tri 34035 38850 34063 38878 sw
rect 33158 28712 33225 38850
tri 33225 38813 33262 38850 nw
tri 33913 38785 33938 38810 se
rect 33938 38785 34038 38810
tri 34038 38785 34063 38810 nw
rect 33913 38747 34038 38785
rect 33913 35173 33980 38747
tri 34038 35328 34097 35387 sw
rect 34038 35173 34146 35328
rect 33913 35161 34146 35173
tri 33913 35136 33938 35161 ne
rect 33938 35136 34121 35161
tri 34121 35136 34146 35161 nw
tri 33913 34924 33938 34949 se
rect 33938 34924 34121 34949
tri 34121 34924 34146 34949 sw
rect 33913 34656 34146 34924
tri 33913 34631 33938 34656 ne
rect 33938 34631 34121 34656
tri 34121 34631 34146 34656 nw
tri 33913 34412 33938 34437 se
rect 33938 34412 34041 34437
tri 34041 34412 34066 34437 nw
rect 33913 34409 34038 34412
tri 34038 34409 34041 34412 nw
rect 33913 28819 33980 34409
rect 33913 28782 34038 28819
tri 33913 28755 33940 28782 ne
rect 33940 28755 34038 28782
tri 34038 28755 34063 28780 sw
tri 33158 28703 33167 28712 ne
rect 33167 28703 33225 28712
tri 33225 28703 33276 28754 sw
tri 33167 28675 33195 28703 ne
rect 33195 28675 34035 28703
tri 34035 28675 34063 28703 nw
tri 34635 28164 34699 28228 sw
rect 34635 28081 34708 28164
tri 34534 28038 34577 28081 se
rect 34577 28044 34708 28081
rect 34577 28038 34702 28044
tri 34702 28038 34708 28044 nw
rect 34534 28019 34683 28038
tri 34683 28019 34702 28038 nw
rect 39872 26910 39992 26938
tri 39992 26912 40018 26938 nw
tri 40271 26912 40297 26938 ne
rect 40297 26912 40415 26938
tri 40297 26911 40298 26912 ne
rect 40298 26910 40415 26912
rect 39872 26420 39946 26910
rect 40344 26420 40415 26910
tri 39872 26391 39901 26420 nw
tri 41044 25984 41070 26010 se
rect 40990 25866 41070 25984
tri 41044 25840 41070 25866 ne
tri 41044 21705 41070 21731 se
rect 40990 21587 41070 21705
tri 41043 21560 41070 21587 ne
tri 39847 7540 39875 7568 ne
rect 39875 7540 44708 7568
rect 44644 7445 44708 7540
rect 44644 7338 44754 7445
tri 44754 7399 44800 7445 nw
tri 44319 7314 44343 7338 ne
rect 44343 7292 44754 7338
rect 36140 5052 36211 5902
tri 36257 5244 36365 5352 sw
tri 38305 5145 38333 5173 ne
rect 38333 5145 44018 5173
tri 44018 5145 44046 5173 nw
rect 36140 4983 37857 5052
tri 37857 4983 37926 5052 sw
rect 35647 1022 35713 4755
rect 36519 4350 36577 4356
rect 36519 4316 36531 4350
rect 36565 4316 36577 4350
rect 36519 4278 36577 4316
rect 36519 4244 36531 4278
rect 36565 4244 36577 4278
rect 36519 4238 36577 4244
rect 40007 4350 40065 4356
rect 40007 4316 40019 4350
rect 40053 4316 40065 4350
rect 40007 4278 40065 4316
rect 40007 4244 40019 4278
rect 40053 4244 40065 4278
rect 40007 4238 40065 4244
rect 40724 4350 40782 4356
rect 40724 4316 40736 4350
rect 40770 4316 40782 4350
rect 40724 4278 40782 4316
rect 40724 4244 40736 4278
rect 40770 4244 40782 4278
rect 40724 4238 40782 4244
rect 44212 4350 44270 4356
rect 44212 4316 44224 4350
rect 44258 4316 44270 4350
rect 44212 4278 44270 4316
rect 44212 4244 44224 4278
rect 44258 4244 44270 4278
rect 44212 4238 44270 4244
tri 36001 3442 36029 3470 ne
rect 36029 3442 44618 3470
tri 44618 3442 44646 3470 nw
tri 44598 3422 44618 3442 nw
rect 36029 1777 43445 1780
tri 43445 1777 43448 1780 nw
tri 36004 1752 36029 1777 se
rect 36029 1752 43420 1777
tri 43420 1752 43445 1777 nw
tri 43362 1694 43420 1752 nw
tri 43572 1379 43597 1404 se
rect 43597 1379 44223 1407
tri 44223 1379 44248 1404 sw
tri 35687 996 35713 1022 ne
rect 35045 -303 36056 -301
tri 36056 -303 36058 -301 nw
tri 35019 -329 35045 -303 se
rect 35045 -329 36030 -303
tri 36030 -329 36056 -303 nw
tri 36026 -333 36030 -329 nw
<< metal2 >>
rect 40150 11958 40206 11967
rect 40150 11758 40206 11902
rect 40150 11558 40206 11702
rect 40150 11358 40206 11502
rect 40150 11293 40206 11302
rect 41082 11958 41138 11967
rect 41082 11758 41138 11902
rect 41082 11558 41138 11702
rect 41082 11358 41138 11502
rect 41082 11293 41138 11302
rect 41548 11958 41604 11967
rect 41548 11758 41604 11902
rect 41548 11558 41604 11702
rect 41548 11358 41604 11502
rect 41548 11293 41604 11302
rect 41716 11958 41772 11967
rect 41716 11758 41772 11902
rect 41716 11558 41772 11702
rect 41716 11358 41772 11502
rect 41716 11293 41772 11302
rect 43002 11958 43058 11967
rect 43002 11758 43058 11902
rect 43002 11558 43058 11702
rect 43002 11358 43058 11502
rect 43002 11293 43058 11302
rect 43393 11958 43449 11967
rect 43393 11758 43449 11902
rect 43393 11558 43449 11702
rect 43393 11358 43449 11502
rect 43393 11293 43449 11302
rect 43743 11958 43799 11967
rect 43743 11758 43799 11902
rect 43743 11558 43799 11702
rect 43743 11358 43799 11502
rect 43743 11293 43799 11302
rect 35298 6486 35354 6495
rect 35298 6286 35354 6430
rect 35298 6086 35354 6230
rect 35298 5886 35354 6030
rect 35298 5821 35354 5830
rect 37770 6486 37826 6495
rect 37770 6286 37826 6430
rect 37770 6086 37826 6230
rect 37770 5886 37826 6030
rect 37770 5821 37826 5830
rect 32854 3737 32910 3746
rect 32854 3537 32910 3681
rect 32854 3337 32910 3481
rect 32854 3137 32910 3281
rect 32854 3072 32910 3081
rect 33940 3737 33996 3746
rect 33940 3537 33996 3681
rect 33940 3337 33996 3481
rect 33940 3137 33996 3281
rect 33940 3072 33996 3081
rect 40332 3734 40388 3743
rect 40332 3534 40388 3678
rect 40332 3334 40388 3478
rect 40332 3134 40388 3278
rect 40332 3069 40388 3078
rect 44374 3734 44430 3743
rect 44374 3534 44430 3678
rect 44374 3334 44430 3478
rect 44374 3134 44430 3278
rect 44374 3069 44430 3078
<< via2 >>
rect 40150 11902 40206 11958
rect 40150 11702 40206 11758
rect 40150 11502 40206 11558
rect 40150 11302 40206 11358
rect 41082 11902 41138 11958
rect 41082 11702 41138 11758
rect 41082 11502 41138 11558
rect 41082 11302 41138 11358
rect 41548 11902 41604 11958
rect 41548 11702 41604 11758
rect 41548 11502 41604 11558
rect 41548 11302 41604 11358
rect 41716 11902 41772 11958
rect 41716 11702 41772 11758
rect 41716 11502 41772 11558
rect 41716 11302 41772 11358
rect 43002 11902 43058 11958
rect 43002 11702 43058 11758
rect 43002 11502 43058 11558
rect 43002 11302 43058 11358
rect 43393 11902 43449 11958
rect 43393 11702 43449 11758
rect 43393 11502 43449 11558
rect 43393 11302 43449 11358
rect 43743 11902 43799 11958
rect 43743 11702 43799 11758
rect 43743 11502 43799 11558
rect 43743 11302 43799 11358
rect 35298 6430 35354 6486
rect 35298 6230 35354 6286
rect 35298 6030 35354 6086
rect 35298 5830 35354 5886
rect 37770 6430 37826 6486
rect 37770 6230 37826 6286
rect 37770 6030 37826 6086
rect 37770 5830 37826 5886
rect 32854 3681 32910 3737
rect 32854 3481 32910 3537
rect 32854 3281 32910 3337
rect 32854 3081 32910 3137
rect 33940 3681 33996 3737
rect 33940 3481 33996 3537
rect 33940 3281 33996 3337
rect 33940 3081 33996 3137
rect 40332 3678 40388 3734
rect 40332 3478 40388 3534
rect 40332 3278 40388 3334
rect 40332 3078 40388 3134
rect 44374 3678 44430 3734
rect 44374 3478 44430 3534
rect 44374 3278 44430 3334
rect 44374 3078 44430 3134
<< metal3 >>
rect 40145 11958 40211 11963
rect 40145 11902 40150 11958
rect 40206 11902 40211 11958
rect 40145 11758 40211 11902
rect 40145 11702 40150 11758
rect 40206 11702 40211 11758
rect 40145 11558 40211 11702
rect 40145 11502 40150 11558
rect 40206 11502 40211 11558
rect 40145 11358 40211 11502
rect 40145 11302 40150 11358
rect 40206 11302 40211 11358
rect 40145 11297 40211 11302
rect 41077 11958 41143 11963
rect 41077 11902 41082 11958
rect 41138 11902 41143 11958
rect 41077 11758 41143 11902
rect 41077 11702 41082 11758
rect 41138 11702 41143 11758
rect 41077 11558 41143 11702
rect 41077 11502 41082 11558
rect 41138 11502 41143 11558
rect 41077 11358 41143 11502
rect 41077 11302 41082 11358
rect 41138 11302 41143 11358
rect 41077 11297 41143 11302
rect 41543 11958 41609 11963
rect 41543 11902 41548 11958
rect 41604 11902 41609 11958
rect 41543 11758 41609 11902
rect 41543 11702 41548 11758
rect 41604 11702 41609 11758
rect 41543 11558 41609 11702
rect 41543 11502 41548 11558
rect 41604 11502 41609 11558
rect 41543 11358 41609 11502
rect 41543 11302 41548 11358
rect 41604 11302 41609 11358
rect 41543 11297 41609 11302
rect 41711 11958 41777 11963
rect 41711 11902 41716 11958
rect 41772 11902 41777 11958
rect 41711 11758 41777 11902
rect 41711 11702 41716 11758
rect 41772 11702 41777 11758
rect 41711 11558 41777 11702
rect 41711 11502 41716 11558
rect 41772 11502 41777 11558
rect 41711 11358 41777 11502
rect 41711 11302 41716 11358
rect 41772 11302 41777 11358
rect 41711 11297 41777 11302
rect 42997 11958 43063 11963
rect 42997 11902 43002 11958
rect 43058 11902 43063 11958
rect 42997 11758 43063 11902
rect 42997 11702 43002 11758
rect 43058 11702 43063 11758
rect 42997 11558 43063 11702
rect 42997 11502 43002 11558
rect 43058 11502 43063 11558
rect 42997 11358 43063 11502
rect 42997 11302 43002 11358
rect 43058 11302 43063 11358
rect 42997 11297 43063 11302
rect 43388 11958 43454 11963
rect 43388 11902 43393 11958
rect 43449 11902 43454 11958
rect 43388 11758 43454 11902
rect 43388 11702 43393 11758
rect 43449 11702 43454 11758
rect 43388 11558 43454 11702
rect 43388 11502 43393 11558
rect 43449 11502 43454 11558
rect 43388 11358 43454 11502
rect 43388 11302 43393 11358
rect 43449 11302 43454 11358
rect 43388 11297 43454 11302
rect 43738 11958 43804 11963
rect 43738 11902 43743 11958
rect 43799 11902 43804 11958
rect 43738 11758 43804 11902
rect 43738 11702 43743 11758
rect 43799 11702 43804 11758
rect 43738 11558 43804 11702
rect 43738 11502 43743 11558
rect 43799 11502 43804 11558
rect 43738 11358 43804 11502
rect 43738 11302 43743 11358
rect 43799 11302 43804 11358
rect 43738 11297 43804 11302
rect 35293 6486 35359 6491
rect 35293 6430 35298 6486
rect 35354 6430 35359 6486
rect 35293 6286 35359 6430
rect 35293 6230 35298 6286
rect 35354 6230 35359 6286
rect 35293 6086 35359 6230
rect 35293 6030 35298 6086
rect 35354 6030 35359 6086
rect 35293 5886 35359 6030
rect 35293 5830 35298 5886
rect 35354 5830 35359 5886
rect 35293 5825 35359 5830
rect 37765 6486 37831 6491
rect 37765 6430 37770 6486
rect 37826 6430 37831 6486
rect 37765 6286 37831 6430
rect 37765 6230 37770 6286
rect 37826 6230 37831 6286
rect 37765 6086 37831 6230
rect 37765 6030 37770 6086
rect 37826 6030 37831 6086
rect 37765 5886 37831 6030
rect 37765 5830 37770 5886
rect 37826 5830 37831 5886
rect 37765 5825 37831 5830
rect 32849 3737 32915 3742
rect 32849 3681 32854 3737
rect 32910 3681 32915 3737
rect 32849 3537 32915 3681
rect 32849 3481 32854 3537
rect 32910 3481 32915 3537
rect 32849 3337 32915 3481
rect 32849 3281 32854 3337
rect 32910 3281 32915 3337
rect 32849 3137 32915 3281
rect 32849 3081 32854 3137
rect 32910 3081 32915 3137
rect 32849 3076 32915 3081
rect 33935 3737 34001 3742
rect 33935 3681 33940 3737
rect 33996 3681 34001 3737
rect 33935 3537 34001 3681
rect 33935 3481 33940 3537
rect 33996 3481 34001 3537
rect 33935 3337 34001 3481
rect 33935 3281 33940 3337
rect 33996 3281 34001 3337
rect 33935 3137 34001 3281
rect 33935 3081 33940 3137
rect 33996 3081 34001 3137
rect 33935 3076 34001 3081
rect 40327 3734 40393 3739
rect 40327 3678 40332 3734
rect 40388 3678 40393 3734
rect 40327 3534 40393 3678
rect 40327 3478 40332 3534
rect 40388 3478 40393 3534
rect 40327 3334 40393 3478
rect 40327 3278 40332 3334
rect 40388 3278 40393 3334
rect 40327 3134 40393 3278
rect 40327 3078 40332 3134
rect 40388 3078 40393 3134
rect 40327 3073 40393 3078
rect 44369 3734 44435 3739
rect 44369 3678 44374 3734
rect 44430 3678 44435 3734
rect 44369 3534 44435 3678
rect 44369 3478 44374 3534
rect 44430 3478 44435 3534
rect 44369 3334 44435 3478
rect 44369 3278 44374 3334
rect 44430 3278 44435 3334
rect 44369 3134 44435 3278
rect 44369 3078 44374 3134
rect 44430 3078 44435 3134
rect 44369 3073 44435 3078
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_0
timestamp 1701704242
transform 1 0 36531 0 1 4244
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_1
timestamp 1701704242
transform 1 0 40019 0 1 4244
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_2
timestamp 1701704242
transform 1 0 40736 0 1 4244
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_3
timestamp 1701704242
transform 1 0 44224 0 1 4244
box 0 0 1 1
use M2M3_CDNS_5246887918519  M2M3_CDNS_5246887918519_0
timestamp 1701704242
transform 1 0 38912 0 1 11293
box -5 0 461 674
use M2M3_CDNS_5246887918520  M2M3_CDNS_5246887918520_0
timestamp 1701704242
transform 1 0 36530 0 1 11293
box -5 0 381 674
use M2M3_CDNS_5246887918521  M2M3_CDNS_5246887918521_0
timestamp 1701704242
transform 1 0 33600 0 1 11293
box -5 0 221 674
use M2M3_CDNS_5246887918521  M2M3_CDNS_5246887918521_1
timestamp 1701704242
transform 1 0 36078 0 1 11293
box -5 0 221 674
use M2M3_CDNS_5246887918521  M2M3_CDNS_5246887918521_2
timestamp 1701704242
transform 1 0 35129 0 1 11293
box -5 0 221 674
use M2M3_CDNS_5246887918521  M2M3_CDNS_5246887918521_3
timestamp 1701704242
transform 1 0 37751 0 1 11293
box -5 0 221 674
use M2M3_CDNS_5246887918521  M2M3_CDNS_5246887918521_4
timestamp 1701704242
transform 1 0 40416 0 1 11293
box -5 0 221 674
use M2M3_CDNS_5246887918521  M2M3_CDNS_5246887918521_5
timestamp 1701704242
transform 1 0 40740 0 1 11293
box -5 0 221 674
use M2M3_CDNS_5246887918521  M2M3_CDNS_5246887918521_6
timestamp 1701704242
transform 1 0 42036 0 1 11293
box -5 0 221 674
use M2M3_CDNS_5246887918521  M2M3_CDNS_5246887918521_7
timestamp 1701704242
transform 1 0 42364 0 1 11293
box -5 0 221 674
use M2M3_CDNS_5246887918522  M2M3_CDNS_5246887918522_0
timestamp 1701704242
transform 1 0 34253 0 1 3069
box -5 0 301 674
use M2M3_CDNS_5246887918522  M2M3_CDNS_5246887918522_1
timestamp 1701704242
transform 1 0 33114 0 1 11293
box -5 0 301 674
use M2M3_CDNS_5246887918523  M2M3_CDNS_5246887918523_0
timestamp 1701704242
transform 1 0 32854 0 1 3072
box 0 0 1 1
use M2M3_CDNS_5246887918523  M2M3_CDNS_5246887918523_1
timestamp 1701704242
transform 1 0 33940 0 1 3072
box 0 0 1 1
use M2M3_CDNS_5246887918523  M2M3_CDNS_5246887918523_2
timestamp 1701704242
transform 1 0 40332 0 1 3069
box 0 0 1 1
use M2M3_CDNS_5246887918523  M2M3_CDNS_5246887918523_3
timestamp 1701704242
transform 1 0 44374 0 1 3069
box 0 0 1 1
use M2M3_CDNS_5246887918523  M2M3_CDNS_5246887918523_4
timestamp 1701704242
transform 1 0 35298 0 1 5821
box 0 0 1 1
use M2M3_CDNS_5246887918523  M2M3_CDNS_5246887918523_5
timestamp 1701704242
transform 1 0 37770 0 1 5821
box 0 0 1 1
use M2M3_CDNS_5246887918523  M2M3_CDNS_5246887918523_6
timestamp 1701704242
transform 1 0 41082 0 1 11293
box 0 0 1 1
use M2M3_CDNS_5246887918523  M2M3_CDNS_5246887918523_7
timestamp 1701704242
transform 1 0 41548 0 1 11293
box 0 0 1 1
use M2M3_CDNS_5246887918523  M2M3_CDNS_5246887918523_8
timestamp 1701704242
transform 1 0 41716 0 1 11293
box 0 0 1 1
use M2M3_CDNS_5246887918523  M2M3_CDNS_5246887918523_9
timestamp 1701704242
transform 1 0 40150 0 1 11293
box 0 0 1 1
use M2M3_CDNS_5246887918523  M2M3_CDNS_5246887918523_10
timestamp 1701704242
transform 1 0 43743 0 1 11293
box 0 0 1 1
use M2M3_CDNS_5246887918523  M2M3_CDNS_5246887918523_11
timestamp 1701704242
transform 1 0 43393 0 1 11293
box 0 0 1 1
use M2M3_CDNS_5246887918523  M2M3_CDNS_5246887918523_12
timestamp 1701704242
transform 1 0 43002 0 1 11293
box 0 0 1 1
use M2M3_CDNS_5246887918524  M2M3_CDNS_5246887918524_0
timestamp 1701704242
transform 1 0 32764 0 1 5864
box -5 0 141 674
use M2M3_CDNS_5246887918524  M2M3_CDNS_5246887918524_1
timestamp 1701704242
transform 1 0 33909 0 1 5864
box -5 0 141 674
use M2M3_CDNS_5246887918524  M2M3_CDNS_5246887918524_2
timestamp 1701704242
transform 1 0 34462 0 1 5864
box -5 0 141 674
use M2M3_CDNS_5246887918524  M2M3_CDNS_5246887918524_3
timestamp 1701704242
transform 1 0 40432 0 1 5864
box -5 0 141 674
use M2M3_CDNS_5246887918524  M2M3_CDNS_5246887918524_4
timestamp 1701704242
transform 1 0 44368 0 1 5864
box -5 0 141 674
<< properties >>
string GDS_END 78405010
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 78401718
<< end >>
