magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< locali >>
rect -17 1137 17 1153
rect -17 1087 17 1103
rect 1784 1137 1818 1153
rect 1784 1087 1818 1103
rect 21752 1137 21786 1153
rect 21752 1087 21786 1103
rect 41720 1137 41754 1153
rect 41720 1087 41754 1103
rect 61688 1137 61722 1153
rect 61688 1087 61722 1103
rect 81229 1137 81263 1153
rect 81229 1087 81263 1103
rect 1586 535 1620 551
rect 1935 517 1969 551
rect 21554 535 21588 551
rect 1586 485 1620 501
rect 21903 517 21937 551
rect 41522 535 41556 551
rect 21554 485 21588 501
rect 41871 517 41905 551
rect 61490 535 61524 551
rect 41522 485 41556 501
rect 61839 517 61873 551
rect 61490 485 61524 501
rect 1357 287 1391 303
rect 21325 287 21359 303
rect 41293 287 41327 303
rect 61261 287 61295 303
rect 1391 253 1503 287
rect 21359 253 21471 287
rect 41327 253 41439 287
rect 61295 253 61407 287
rect 1357 237 1391 253
rect 21325 237 21359 253
rect 41293 237 41327 253
rect 61261 237 61295 253
rect -17 17 17 33
rect -17 -33 17 -17
rect 1784 17 1818 33
rect 1784 -33 1818 -17
rect 21752 17 21786 33
rect 21752 -33 21786 -17
rect 41720 17 41754 33
rect 41720 -33 41754 -17
rect 61688 17 61722 33
rect 61688 -33 61722 -17
rect 81229 17 81263 33
rect 81229 -33 81263 -17
<< viali >>
rect -17 1103 17 1137
rect 1784 1103 1818 1137
rect 21752 1103 21786 1137
rect 41720 1103 41754 1137
rect 61688 1103 61722 1137
rect 81229 1103 81263 1137
rect 1586 501 1620 535
rect 21554 501 21588 535
rect 41522 501 41556 535
rect 61490 501 61524 535
rect 1357 253 1391 287
rect 21325 253 21359 287
rect 41293 253 41327 287
rect 61261 253 61295 287
rect -17 -17 17 17
rect 1784 -17 1818 17
rect 21752 -17 21786 17
rect 41720 -17 41754 17
rect 61688 -17 61722 17
rect 81229 -17 81263 17
<< metal1 >>
rect -32 1094 -26 1146
rect 26 1134 32 1146
rect 1772 1137 1830 1143
rect 1772 1134 1784 1137
rect 26 1106 1784 1134
rect 26 1094 32 1106
rect 1772 1103 1784 1106
rect 1818 1134 1830 1137
rect 21740 1137 21798 1143
rect 21740 1134 21752 1137
rect 1818 1106 21752 1134
rect 1818 1103 1830 1106
rect 1772 1097 1830 1103
rect 21740 1103 21752 1106
rect 21786 1134 21798 1137
rect 41708 1137 41766 1143
rect 41708 1134 41720 1137
rect 21786 1106 41720 1134
rect 21786 1103 21798 1106
rect 21740 1097 21798 1103
rect 41708 1103 41720 1106
rect 41754 1134 41766 1137
rect 61676 1137 61734 1143
rect 61676 1134 61688 1137
rect 41754 1106 61688 1134
rect 41754 1103 41766 1106
rect 41708 1097 41766 1103
rect 61676 1103 61688 1106
rect 61722 1134 61734 1137
rect 81214 1134 81220 1146
rect 61722 1106 81220 1134
rect 61722 1103 61734 1106
rect 61676 1097 61734 1103
rect 81214 1094 81220 1106
rect 81272 1094 81278 1146
rect 1571 492 1577 544
rect 1629 492 1635 544
rect 21539 492 21545 544
rect 21597 492 21603 544
rect 41507 492 41513 544
rect 41565 492 41571 544
rect 61475 492 61481 544
rect 61533 492 61539 544
rect 1342 244 1348 296
rect 1400 244 1406 296
rect 21310 244 21316 296
rect 21368 244 21374 296
rect 41278 244 41284 296
rect 41336 244 41342 296
rect 61246 244 61252 296
rect 61304 244 61310 296
rect -32 -26 -26 26
rect 26 14 32 26
rect 1772 17 1830 23
rect 1772 14 1784 17
rect 26 -14 1784 14
rect 26 -26 32 -14
rect 1772 -17 1784 -14
rect 1818 14 1830 17
rect 21740 17 21798 23
rect 21740 14 21752 17
rect 1818 -14 21752 14
rect 1818 -17 1830 -14
rect 1772 -23 1830 -17
rect 21740 -17 21752 -14
rect 21786 14 21798 17
rect 41708 17 41766 23
rect 41708 14 41720 17
rect 21786 -14 41720 14
rect 21786 -17 21798 -14
rect 21740 -23 21798 -17
rect 41708 -17 41720 -14
rect 41754 14 41766 17
rect 61676 17 61734 23
rect 61676 14 61688 17
rect 41754 -14 61688 14
rect 41754 -17 41766 -14
rect 41708 -23 41766 -17
rect 61676 -17 61688 -14
rect 61722 14 61734 17
rect 81214 14 81220 26
rect 61722 -14 81220 14
rect 61722 -17 61734 -14
rect 61676 -23 61734 -17
rect 81214 -26 81220 -14
rect 81272 -26 81278 26
<< via1 >>
rect -26 1137 26 1146
rect -26 1103 -17 1137
rect -17 1103 17 1137
rect 17 1103 26 1137
rect -26 1094 26 1103
rect 81220 1137 81272 1146
rect 81220 1103 81229 1137
rect 81229 1103 81263 1137
rect 81263 1103 81272 1137
rect 81220 1094 81272 1103
rect 1577 535 1629 544
rect 1577 501 1586 535
rect 1586 501 1620 535
rect 1620 501 1629 535
rect 1577 492 1629 501
rect 21545 535 21597 544
rect 21545 501 21554 535
rect 21554 501 21588 535
rect 21588 501 21597 535
rect 21545 492 21597 501
rect 41513 535 41565 544
rect 41513 501 41522 535
rect 41522 501 41556 535
rect 41556 501 41565 535
rect 41513 492 41565 501
rect 61481 535 61533 544
rect 61481 501 61490 535
rect 61490 501 61524 535
rect 61524 501 61533 535
rect 61481 492 61533 501
rect 1348 287 1400 296
rect 1348 253 1357 287
rect 1357 253 1391 287
rect 1391 253 1400 287
rect 1348 244 1400 253
rect 21316 287 21368 296
rect 21316 253 21325 287
rect 21325 253 21359 287
rect 21359 253 21368 287
rect 21316 244 21368 253
rect 41284 287 41336 296
rect 41284 253 41293 287
rect 41293 253 41327 287
rect 41327 253 41336 287
rect 41284 244 41336 253
rect 61252 287 61304 296
rect 61252 253 61261 287
rect 61261 253 61295 287
rect 61295 253 61304 287
rect 61252 244 61304 253
rect -26 17 26 26
rect -26 -17 -17 17
rect -17 -17 17 17
rect 17 -17 26 17
rect -26 -26 26 -17
rect 81220 17 81272 26
rect 81220 -17 81229 17
rect 81229 -17 81263 17
rect 81263 -17 81272 17
rect 81220 -26 81272 -17
<< metal2 >>
rect -28 1148 28 1157
rect -28 1083 28 1092
rect 81218 1148 81274 1157
rect 81218 1083 81274 1092
rect 1575 546 1631 555
rect 1575 481 1631 490
rect 21543 546 21599 555
rect 21543 481 21599 490
rect 41511 546 41567 555
rect 41511 481 41567 490
rect 61479 546 61535 555
rect 61479 481 61535 490
rect 1348 296 1400 302
rect 1348 238 1400 244
rect 21316 296 21368 302
rect 21316 238 21368 244
rect 41284 296 41336 302
rect 41284 238 41336 244
rect 61252 296 61304 302
rect 61252 238 61304 244
rect -28 28 28 37
rect -28 -37 28 -28
rect 81218 28 81274 37
rect 81218 -37 81274 -28
<< via2 >>
rect -28 1146 28 1148
rect -28 1094 -26 1146
rect -26 1094 26 1146
rect 26 1094 28 1146
rect -28 1092 28 1094
rect 81218 1146 81274 1148
rect 81218 1094 81220 1146
rect 81220 1094 81272 1146
rect 81272 1094 81274 1146
rect 81218 1092 81274 1094
rect 1575 544 1631 546
rect 1575 492 1577 544
rect 1577 492 1629 544
rect 1629 492 1631 544
rect 1575 490 1631 492
rect 21543 544 21599 546
rect 21543 492 21545 544
rect 21545 492 21597 544
rect 21597 492 21599 544
rect 21543 490 21599 492
rect 41511 544 41567 546
rect 41511 492 41513 544
rect 41513 492 41565 544
rect 41565 492 41567 544
rect 41511 490 41567 492
rect 61479 544 61535 546
rect 61479 492 61481 544
rect 61481 492 61533 544
rect 61533 492 61535 544
rect 61479 490 61535 492
rect -28 26 28 28
rect -28 -26 -26 26
rect -26 -26 26 26
rect 26 -26 28 26
rect -28 -28 28 -26
rect 81218 26 81274 28
rect 81218 -26 81220 26
rect 81220 -26 81272 26
rect 81272 -26 81274 26
rect 81218 -28 81274 -26
<< metal3 >>
rect -49 1148 49 1169
rect -49 1092 -28 1148
rect 28 1092 49 1148
rect -49 1071 49 1092
rect 81197 1148 81295 1169
rect 81197 1092 81218 1148
rect 81274 1092 81295 1148
rect 81197 1071 81295 1092
rect 1570 548 1636 551
rect 21538 548 21604 551
rect 41506 548 41572 551
rect 61474 548 61540 551
rect 0 546 81246 548
rect 0 490 1575 546
rect 1631 490 21543 546
rect 21599 490 41511 546
rect 41567 490 61479 546
rect 61535 490 81246 546
rect 0 488 81246 490
rect 1570 485 1636 488
rect 21538 485 21604 488
rect 41506 485 41572 488
rect 61474 485 61540 488
rect -49 28 49 49
rect -49 -28 -28 28
rect 28 -28 49 28
rect -49 -49 49 -28
rect 81197 28 81295 49
rect 81197 -28 81218 28
rect 81274 -28 81295 28
rect 81197 -49 81295 -28
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_0
timestamp 1701704242
transform 1 0 81213 0 1 1083
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_1
timestamp 1701704242
transform 1 0 -33 0 1 1083
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_2
timestamp 1701704242
transform 1 0 81213 0 1 -37
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_3
timestamp 1701704242
transform 1 0 -33 0 1 -37
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_4
timestamp 1701704242
transform 1 0 61474 0 1 481
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_5
timestamp 1701704242
transform 1 0 41506 0 1 481
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_6
timestamp 1701704242
transform 1 0 21538 0 1 481
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_7
timestamp 1701704242
transform 1 0 1570 0 1 481
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_0
timestamp 1701704242
transform 1 0 81217 0 1 1087
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1
timestamp 1701704242
transform 1 0 -29 0 1 1087
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_2
timestamp 1701704242
transform 1 0 81217 0 1 -33
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_3
timestamp 1701704242
transform 1 0 -29 0 1 -33
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_4
timestamp 1701704242
transform 1 0 61676 0 1 1087
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_5
timestamp 1701704242
transform 1 0 61676 0 1 -33
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_6
timestamp 1701704242
transform 1 0 61478 0 1 485
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_7
timestamp 1701704242
transform 1 0 61249 0 1 237
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_8
timestamp 1701704242
transform 1 0 41708 0 1 1087
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_9
timestamp 1701704242
transform 1 0 41708 0 1 -33
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_10
timestamp 1701704242
transform 1 0 41510 0 1 485
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_11
timestamp 1701704242
transform 1 0 41281 0 1 237
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_12
timestamp 1701704242
transform 1 0 21740 0 1 1087
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_13
timestamp 1701704242
transform 1 0 21740 0 1 -33
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_14
timestamp 1701704242
transform 1 0 21542 0 1 485
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_15
timestamp 1701704242
transform 1 0 21313 0 1 237
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_16
timestamp 1701704242
transform 1 0 1772 0 1 1087
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_17
timestamp 1701704242
transform 1 0 1772 0 1 -33
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_18
timestamp 1701704242
transform 1 0 1574 0 1 485
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_19
timestamp 1701704242
transform 1 0 1345 0 1 237
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_0
timestamp 1701704242
transform 1 0 81214 0 1 1088
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_1
timestamp 1701704242
transform 1 0 -32 0 1 1088
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_2
timestamp 1701704242
transform 1 0 81214 0 1 -32
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_3
timestamp 1701704242
transform 1 0 -32 0 1 -32
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_4
timestamp 1701704242
transform 1 0 61475 0 1 486
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_5
timestamp 1701704242
transform 1 0 61246 0 1 238
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_6
timestamp 1701704242
transform 1 0 41507 0 1 486
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_7
timestamp 1701704242
transform 1 0 41278 0 1 238
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_8
timestamp 1701704242
transform 1 0 21539 0 1 486
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_9
timestamp 1701704242
transform 1 0 21310 0 1 238
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_10
timestamp 1701704242
transform 1 0 1571 0 1 486
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_11
timestamp 1701704242
transform 1 0 1342 0 1 238
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_pand2  sky130_sram_2kbyte_1rw1r_32x512_8_pand2_0
timestamp 1701704242
transform 1 0 61278 0 1 0
box -36 -17 890 1177
use sky130_sram_2kbyte_1rw1r_32x512_8_pand2  sky130_sram_2kbyte_1rw1r_32x512_8_pand2_1
timestamp 1701704242
transform 1 0 41310 0 1 0
box -36 -17 890 1177
use sky130_sram_2kbyte_1rw1r_32x512_8_pand2  sky130_sram_2kbyte_1rw1r_32x512_8_pand2_2
timestamp 1701704242
transform 1 0 21342 0 1 0
box -36 -17 890 1177
use sky130_sram_2kbyte_1rw1r_32x512_8_pand2  sky130_sram_2kbyte_1rw1r_32x512_8_pand2_3
timestamp 1701704242
transform 1 0 1374 0 1 0
box -36 -17 890 1177
<< labels >>
rlabel metal3 s 0 488 81246 548 4 en
port 1 nsew
rlabel metal3 s 81197 -49 81295 49 4 gnd
port 2 nsew
rlabel metal3 s -49 -49 49 49 4 gnd
port 2 nsew
rlabel metal3 s 81197 1071 81295 1169 4 vdd
port 3 nsew
rlabel metal3 s -49 1071 49 1169 4 vdd
port 3 nsew
rlabel metal2 s 1360 256 1388 284 4 wmask_in_0
port 4 nsew
rlabel metal2 s 21328 256 21356 284 4 wmask_in_1
port 5 nsew
rlabel metal2 s 41296 256 41324 284 4 wmask_in_2
port 6 nsew
rlabel metal2 s 61264 256 61292 284 4 wmask_in_3
port 7 nsew
rlabel locali s 1952 534 1952 534 4 wmask_out_0
rlabel locali s 21920 534 21920 534 4 wmask_out_1
rlabel locali s 41888 534 41888 534 4 wmask_out_2
rlabel locali s 61856 534 61856 534 4 wmask_out_3
<< properties >>
string FIXED_BBOX 81213 -37 81279 0
string GDS_END 1364624
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_2kbyte_1rw1r_32x512_8.gds
string GDS_START 1357232
<< end >>
