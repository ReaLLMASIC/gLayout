magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -161 -36 2665 636
<< pmoslvt >>
rect 0 0 200 600
rect 256 0 456 600
rect 512 0 712 600
rect 768 0 968 600
rect 1024 0 1224 600
rect 1280 0 1480 600
rect 1536 0 1736 600
rect 1792 0 1992 600
rect 2048 0 2248 600
rect 2304 0 2504 600
<< pdiff >>
rect -50 0 0 600
rect 2504 0 2554 600
<< poly >>
rect 0 600 200 632
rect 0 -32 200 0
rect 256 600 456 632
rect 256 -32 456 0
rect 512 600 712 632
rect 512 -32 712 0
rect 768 600 968 632
rect 768 -32 968 0
rect 1024 600 1224 632
rect 1024 -32 1224 0
rect 1280 600 1480 632
rect 1280 -32 1480 0
rect 1536 600 1736 632
rect 1536 -32 1736 0
rect 1792 600 1992 632
rect 1792 -32 1992 0
rect 2048 600 2248 632
rect 2048 -32 2248 0
rect 2304 600 2504 632
rect 2304 -32 2504 0
<< locali >>
rect 211 -4 245 538
rect 467 -4 501 538
rect 723 -4 757 538
rect 979 -4 1013 538
rect 1235 -4 1269 538
rect 1491 -4 1525 538
rect 1747 -4 1781 538
rect 2003 -4 2037 538
rect 2259 -4 2293 538
<< metal1 >>
rect -51 -16 -5 546
rect 2509 -16 2555 546
use DFL1sd2_CDNS_5246887918535  DFL1sd2_CDNS_5246887918535_0
timestamp 1701704242
transform 1 0 2248 0 1 0
box -36 -36 92 636
use DFL1sd2_CDNS_5246887918535  DFL1sd2_CDNS_5246887918535_1
timestamp 1701704242
transform 1 0 1992 0 1 0
box -36 -36 92 636
use DFL1sd2_CDNS_5246887918535  DFL1sd2_CDNS_5246887918535_2
timestamp 1701704242
transform 1 0 1736 0 1 0
box -36 -36 92 636
use DFL1sd2_CDNS_5246887918535  DFL1sd2_CDNS_5246887918535_3
timestamp 1701704242
transform 1 0 1480 0 1 0
box -36 -36 92 636
use DFL1sd2_CDNS_5246887918535  DFL1sd2_CDNS_5246887918535_4
timestamp 1701704242
transform 1 0 1224 0 1 0
box -36 -36 92 636
use DFL1sd2_CDNS_5246887918535  DFL1sd2_CDNS_5246887918535_5
timestamp 1701704242
transform 1 0 968 0 1 0
box -36 -36 92 636
use DFL1sd2_CDNS_5246887918535  DFL1sd2_CDNS_5246887918535_6
timestamp 1701704242
transform 1 0 712 0 1 0
box -36 -36 92 636
use DFL1sd2_CDNS_5246887918535  DFL1sd2_CDNS_5246887918535_7
timestamp 1701704242
transform 1 0 456 0 1 0
box -36 -36 92 636
use DFL1sd2_CDNS_5246887918535  DFL1sd2_CDNS_5246887918535_8
timestamp 1701704242
transform 1 0 200 0 1 0
box -36 -36 92 636
use DFTPM1s_CDNS_524688791851273  DFTPM1s_CDNS_524688791851273_0
timestamp 1701704242
transform -1 0 0 0 1 0
box -36 -36 161 636
use DFTPM1s_CDNS_524688791851273  DFTPM1s_CDNS_524688791851273_1
timestamp 1701704242
transform 1 0 2504 0 1 0
box -36 -36 161 636
<< labels >>
flabel comment s -28 265 -28 265 0 FreeSans 300 0 0 0 S
flabel comment s 228 267 228 267 0 FreeSans 300 0 0 0 D
flabel comment s 484 267 484 267 0 FreeSans 300 0 0 0 S
flabel comment s 740 267 740 267 0 FreeSans 300 0 0 0 D
flabel comment s 996 267 996 267 0 FreeSans 300 0 0 0 S
flabel comment s 1252 267 1252 267 0 FreeSans 300 0 0 0 D
flabel comment s 1508 267 1508 267 0 FreeSans 300 0 0 0 S
flabel comment s 1764 267 1764 267 0 FreeSans 300 0 0 0 D
flabel comment s 2020 267 2020 267 0 FreeSans 300 0 0 0 S
flabel comment s 2276 267 2276 267 0 FreeSans 300 0 0 0 D
flabel comment s 2532 265 2532 265 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 86606554
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86601136
<< end >>
