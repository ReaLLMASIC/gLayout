magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< pwell >>
rect -79 -26 551 226
<< mvnmos >>
rect 0 0 120 200
rect 176 0 296 200
rect 352 0 472 200
<< mvndiff >>
rect -53 182 0 200
rect -53 148 -45 182
rect -11 148 0 182
rect -53 114 0 148
rect -53 80 -45 114
rect -11 80 0 114
rect -53 46 0 80
rect -53 12 -45 46
rect -11 12 0 46
rect -53 0 0 12
rect 120 182 176 200
rect 120 148 131 182
rect 165 148 176 182
rect 120 114 176 148
rect 120 80 131 114
rect 165 80 176 114
rect 120 46 176 80
rect 120 12 131 46
rect 165 12 176 46
rect 120 0 176 12
rect 296 182 352 200
rect 296 148 307 182
rect 341 148 352 182
rect 296 114 352 148
rect 296 80 307 114
rect 341 80 352 114
rect 296 46 352 80
rect 296 12 307 46
rect 341 12 352 46
rect 296 0 352 12
rect 472 182 525 200
rect 472 148 483 182
rect 517 148 525 182
rect 472 114 525 148
rect 472 80 483 114
rect 517 80 525 114
rect 472 46 525 80
rect 472 12 483 46
rect 517 12 525 46
rect 472 0 525 12
<< mvndiffc >>
rect -45 148 -11 182
rect -45 80 -11 114
rect -45 12 -11 46
rect 131 148 165 182
rect 131 80 165 114
rect 131 12 165 46
rect 307 148 341 182
rect 307 80 341 114
rect 307 12 341 46
rect 483 148 517 182
rect 483 80 517 114
rect 483 12 517 46
<< poly >>
rect 0 200 120 226
rect 176 200 296 226
rect 352 200 472 226
rect 0 -26 120 0
rect 176 -26 296 0
rect 352 -26 472 0
<< locali >>
rect -45 182 -11 198
rect -45 114 -11 148
rect -45 46 -11 80
rect -45 -4 -11 12
rect 131 182 165 198
rect 131 114 165 148
rect 131 46 165 80
rect 131 -4 165 12
rect 307 182 341 198
rect 307 114 341 148
rect 307 46 341 80
rect 307 -4 341 12
rect 483 182 517 198
rect 483 114 517 148
rect 483 46 517 80
rect 483 -4 517 12
use hvDFL1sd2_CDNS_52468879185133  hvDFL1sd2_CDNS_52468879185133_0
timestamp 1701704242
transform 1 0 296 0 1 0
box 0 0 1 1
use hvDFL1sd2_CDNS_52468879185133  hvDFL1sd2_CDNS_52468879185133_1
timestamp 1701704242
transform 1 0 120 0 1 0
box 0 0 1 1
use hvDFL1sd_CDNS_52468879185132  hvDFL1sd_CDNS_52468879185132_0
timestamp 1701704242
transform -1 0 0 0 1 0
box 0 0 1 1
use hvDFL1sd_CDNS_52468879185132  hvDFL1sd_CDNS_52468879185132_1
timestamp 1701704242
transform 1 0 472 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s -28 97 -28 97 0 FreeSans 300 0 0 0 S
flabel comment s 148 97 148 97 0 FreeSans 300 0 0 0 D
flabel comment s 324 97 324 97 0 FreeSans 300 0 0 0 S
flabel comment s 500 97 500 97 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 85575776
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85573886
<< end >>
