magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< obsli1 >>
rect 48 102 14951 39556
<< metal1 >>
rect 5660 0 5811 244
<< obsm1 >>
rect 24 300 14957 39568
rect 24 0 5604 300
rect 5867 0 14957 300
<< metal2 >>
rect 100 0 4099 115
rect 4515 0 10707 337
rect 10943 0 14940 732
<< obsm2 >>
rect 100 788 14940 38886
rect 100 393 10887 788
rect 100 171 4459 393
rect 4155 0 4459 171
rect 10763 0 10887 393
<< metal3 >>
rect 5008 0 5092 4646
rect 5200 0 7376 4044
rect 7676 0 9851 4580
<< obsm3 >>
rect 3121 4726 12066 37903
rect 3121 4044 4928 4726
rect 5172 4660 12066 4726
rect 5172 4124 7596 4660
rect 7456 4044 7596 4124
rect 9931 4044 12066 4660
<< labels >>
rlabel metal1 s 5660 0 5811 244 6 vssd
port 1 nsew ground bidirectional
rlabel metal2 s 100 0 4099 115 6 src_bdy_lvc1
port 2 nsew ground bidirectional
rlabel metal2 s 10943 0 14940 732 6 src_bdy_lvc2
port 3 nsew ground bidirectional
rlabel metal2 s 4515 0 10707 337 6 bdy2_b2b
port 4 nsew ground bidirectional
rlabel metal3 s 7676 0 9851 4580 6 drn_lvc2
port 5 nsew power bidirectional
rlabel metal3 s 5200 0 7376 4044 6 drn_lvc1
port 6 nsew power bidirectional
rlabel metal3 s 5008 0 5092 4646 6 ogc_lvc
port 7 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 15000 39600
string LEFclass PAD
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 46487740
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 43080384
<< end >>
