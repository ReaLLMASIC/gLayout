magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< nwell >>
rect 5873 927 6041 2669
<< pwell >>
rect -278 38697 6174 38783
rect -278 3492 -192 38697
rect 1804 3492 1890 38697
rect 3946 3492 4032 38697
rect 6088 3492 6174 38697
rect -278 3153 6174 3492
rect 9062 38697 15000 38783
rect 9062 3493 9148 38697
rect 10200 3493 10286 38697
rect 11398 3493 11484 38697
rect 12870 38547 13588 38697
rect 12988 38482 13470 38547
rect 9062 3153 11484 3493
rect 11398 423 11484 3153
rect 11398 359 11682 423
rect 11398 100 11800 359
rect 13186 100 13272 38482
rect 14914 431 15000 38697
rect 14776 359 15000 431
rect 14658 100 15000 359
rect 11398 14 15000 100
rect 11581 -215 14803 14
<< mvndiff >>
rect -138 3394 -80 3466
rect -138 3360 -126 3394
rect -92 3360 -80 3394
rect -138 3352 -80 3360
rect -20 3394 38 3466
rect -20 3360 -8 3394
rect 26 3360 38 3394
rect -20 3352 38 3360
rect 98 3394 156 3466
rect 98 3360 110 3394
rect 144 3360 156 3394
rect 98 3352 156 3360
rect 216 3394 274 3466
rect 216 3360 228 3394
rect 262 3360 274 3394
rect 216 3352 274 3360
rect 334 3394 392 3466
rect 334 3360 346 3394
rect 380 3360 392 3394
rect 334 3352 392 3360
rect 452 3394 510 3466
rect 452 3360 464 3394
rect 498 3360 510 3394
rect 452 3352 510 3360
rect 570 3394 628 3466
rect 570 3360 582 3394
rect 616 3360 628 3394
rect 570 3352 628 3360
rect 688 3394 746 3466
rect 688 3360 700 3394
rect 734 3360 746 3394
rect 688 3352 746 3360
rect 806 3394 864 3466
rect 806 3360 818 3394
rect 852 3360 864 3394
rect 806 3352 864 3360
rect 924 3394 982 3466
rect 924 3360 936 3394
rect 970 3360 982 3394
rect 924 3352 982 3360
rect 1042 3394 1100 3466
rect 1042 3360 1054 3394
rect 1088 3360 1100 3394
rect 1042 3352 1100 3360
rect 1160 3394 1218 3466
rect 1160 3360 1172 3394
rect 1206 3360 1218 3394
rect 1160 3352 1218 3360
rect 1278 3394 1336 3466
rect 1278 3360 1290 3394
rect 1324 3360 1336 3394
rect 1278 3352 1336 3360
rect 1396 3394 1454 3466
rect 1396 3360 1408 3394
rect 1442 3360 1454 3394
rect 1396 3352 1454 3360
rect 1514 3394 1572 3466
rect 1514 3360 1526 3394
rect 1560 3360 1572 3394
rect 1514 3352 1572 3360
rect 1632 3394 1690 3466
rect 1632 3360 1644 3394
rect 1678 3360 1690 3394
rect 1632 3352 1690 3360
rect 2004 3394 2062 3466
rect 2004 3360 2016 3394
rect 2050 3360 2062 3394
rect 2004 3352 2062 3360
rect 2122 3394 2180 3466
rect 2122 3360 2134 3394
rect 2168 3360 2180 3394
rect 2122 3352 2180 3360
rect 2240 3394 2298 3466
rect 2240 3360 2252 3394
rect 2286 3360 2298 3394
rect 2240 3352 2298 3360
rect 2358 3394 2416 3466
rect 2358 3360 2370 3394
rect 2404 3360 2416 3394
rect 2358 3352 2416 3360
rect 2476 3394 2534 3466
rect 2476 3360 2488 3394
rect 2522 3360 2534 3394
rect 2476 3352 2534 3360
rect 2594 3394 2652 3466
rect 2594 3360 2606 3394
rect 2640 3360 2652 3394
rect 2594 3352 2652 3360
rect 2712 3394 2770 3466
rect 2712 3360 2724 3394
rect 2758 3360 2770 3394
rect 2712 3352 2770 3360
rect 2830 3394 2888 3466
rect 2830 3360 2842 3394
rect 2876 3360 2888 3394
rect 2830 3352 2888 3360
rect 2948 3394 3006 3466
rect 2948 3360 2960 3394
rect 2994 3360 3006 3394
rect 2948 3352 3006 3360
rect 3066 3394 3124 3466
rect 3066 3360 3078 3394
rect 3112 3360 3124 3394
rect 3066 3352 3124 3360
rect 3184 3394 3242 3466
rect 3184 3360 3196 3394
rect 3230 3360 3242 3394
rect 3184 3352 3242 3360
rect 3302 3394 3360 3466
rect 3302 3360 3314 3394
rect 3348 3360 3360 3394
rect 3302 3352 3360 3360
rect 3420 3394 3478 3466
rect 3420 3360 3432 3394
rect 3466 3360 3478 3394
rect 3420 3352 3478 3360
rect 3538 3394 3596 3466
rect 3538 3360 3550 3394
rect 3584 3360 3596 3394
rect 3538 3352 3596 3360
rect 3656 3394 3714 3466
rect 3656 3360 3668 3394
rect 3702 3360 3714 3394
rect 3656 3352 3714 3360
rect 3774 3394 3832 3466
rect 3774 3360 3786 3394
rect 3820 3360 3832 3394
rect 3774 3352 3832 3360
rect 4146 3395 4204 3466
rect 4146 3361 4158 3395
rect 4192 3361 4204 3395
rect 4146 3353 4204 3361
rect 4264 3395 4322 3466
rect 4264 3361 4276 3395
rect 4310 3361 4322 3395
rect 4264 3353 4322 3361
rect 4382 3395 4440 3466
rect 4382 3361 4394 3395
rect 4428 3361 4440 3395
rect 4382 3353 4440 3361
rect 4500 3395 4558 3466
rect 4500 3361 4512 3395
rect 4546 3361 4558 3395
rect 4500 3353 4558 3361
rect 4618 3395 4676 3466
rect 4618 3361 4630 3395
rect 4664 3361 4676 3395
rect 4618 3353 4676 3361
rect 4736 3395 4794 3466
rect 4736 3361 4748 3395
rect 4782 3361 4794 3395
rect 4736 3353 4794 3361
rect 4854 3395 4912 3466
rect 4854 3361 4866 3395
rect 4900 3361 4912 3395
rect 4854 3353 4912 3361
rect 4972 3395 5030 3466
rect 4972 3361 4984 3395
rect 5018 3361 5030 3395
rect 4972 3353 5030 3361
rect 5090 3395 5148 3466
rect 5090 3361 5102 3395
rect 5136 3361 5148 3395
rect 5090 3353 5148 3361
rect 5208 3395 5266 3466
rect 5208 3361 5220 3395
rect 5254 3361 5266 3395
rect 5208 3353 5266 3361
rect 5326 3395 5384 3466
rect 5326 3361 5338 3395
rect 5372 3361 5384 3395
rect 5326 3353 5384 3361
rect 5444 3395 5502 3466
rect 5444 3361 5456 3395
rect 5490 3361 5502 3395
rect 5444 3353 5502 3361
rect 5562 3395 5620 3466
rect 5562 3361 5574 3395
rect 5608 3361 5620 3395
rect 5562 3353 5620 3361
rect 5680 3395 5738 3466
rect 5680 3361 5692 3395
rect 5726 3361 5738 3395
rect 5680 3353 5738 3361
rect 5798 3395 5856 3466
rect 5798 3361 5810 3395
rect 5844 3361 5856 3395
rect 5798 3353 5856 3361
rect 5916 3395 5974 3466
rect 5916 3361 5928 3395
rect 5962 3361 5974 3395
rect 5916 3353 5974 3361
rect 9202 3395 9260 3467
rect 9202 3361 9214 3395
rect 9248 3361 9260 3395
rect 9202 3353 9260 3361
rect 9320 3395 9378 3467
rect 9320 3361 9332 3395
rect 9366 3361 9378 3395
rect 9320 3353 9378 3361
rect 9438 3395 9496 3467
rect 9438 3361 9450 3395
rect 9484 3361 9496 3395
rect 9438 3353 9496 3361
rect 9556 3395 9614 3467
rect 9556 3361 9568 3395
rect 9602 3361 9614 3395
rect 9556 3353 9614 3361
rect 9674 3395 9732 3467
rect 9674 3361 9686 3395
rect 9720 3361 9732 3395
rect 9674 3353 9732 3361
rect 9792 3395 9850 3467
rect 9792 3361 9804 3395
rect 9838 3361 9850 3395
rect 9792 3353 9850 3361
rect 9910 3395 9968 3467
rect 9910 3361 9922 3395
rect 9956 3361 9968 3395
rect 9910 3353 9968 3361
rect 10028 3395 10086 3467
rect 10028 3361 10040 3395
rect 10074 3361 10086 3395
rect 10028 3353 10086 3361
rect 12896 38615 13072 38631
rect 12896 38581 12908 38615
rect 12942 38581 13026 38615
rect 13060 38581 13072 38615
rect 12896 38573 13072 38581
rect 13014 38508 13072 38573
rect 10400 3395 10458 3467
rect 10400 3361 10412 3395
rect 10446 3361 10458 3395
rect 10400 3353 10458 3361
rect 10518 3395 10576 3467
rect 10518 3361 10530 3395
rect 10564 3361 10576 3395
rect 10518 3353 10576 3361
rect 10636 3395 10694 3467
rect 10636 3361 10648 3395
rect 10682 3361 10694 3395
rect 10636 3353 10694 3361
rect 10754 3395 10812 3467
rect 10754 3361 10766 3395
rect 10800 3361 10812 3395
rect 10754 3353 10812 3361
rect 10872 3395 10930 3467
rect 10872 3361 10884 3395
rect 10918 3361 10930 3395
rect 10872 3353 10930 3361
rect 10990 3395 11048 3467
rect 10990 3361 11002 3395
rect 11036 3361 11048 3395
rect 10990 3353 11048 3361
rect 11108 3395 11166 3467
rect 11108 3361 11120 3395
rect 11154 3361 11166 3395
rect 11108 3353 11166 3361
rect 11226 3395 11284 3467
rect 11226 3361 11238 3395
rect 11272 3361 11284 3395
rect 11226 3353 11284 3361
rect 13386 38615 13562 38631
rect 13386 38581 13398 38615
rect 13432 38581 13516 38615
rect 13550 38581 13562 38615
rect 13386 38573 13562 38581
rect 13386 38508 13444 38573
rect 11598 333 11656 397
rect 11598 325 11774 333
rect 11598 291 11610 325
rect 11644 291 11724 325
rect 11758 291 11774 325
rect 11598 275 11774 291
rect 14802 333 14860 405
rect 14684 325 14860 333
rect 14684 291 14696 325
rect 14730 291 14814 325
rect 14848 291 14860 325
rect 14684 275 14860 291
<< mvndiffc >>
rect -126 3360 -92 3394
rect -8 3360 26 3394
rect 110 3360 144 3394
rect 228 3360 262 3394
rect 346 3360 380 3394
rect 464 3360 498 3394
rect 582 3360 616 3394
rect 700 3360 734 3394
rect 818 3360 852 3394
rect 936 3360 970 3394
rect 1054 3360 1088 3394
rect 1172 3360 1206 3394
rect 1290 3360 1324 3394
rect 1408 3360 1442 3394
rect 1526 3360 1560 3394
rect 1644 3360 1678 3394
rect 2016 3360 2050 3394
rect 2134 3360 2168 3394
rect 2252 3360 2286 3394
rect 2370 3360 2404 3394
rect 2488 3360 2522 3394
rect 2606 3360 2640 3394
rect 2724 3360 2758 3394
rect 2842 3360 2876 3394
rect 2960 3360 2994 3394
rect 3078 3360 3112 3394
rect 3196 3360 3230 3394
rect 3314 3360 3348 3394
rect 3432 3360 3466 3394
rect 3550 3360 3584 3394
rect 3668 3360 3702 3394
rect 3786 3360 3820 3394
rect 4158 3361 4192 3395
rect 4276 3361 4310 3395
rect 4394 3361 4428 3395
rect 4512 3361 4546 3395
rect 4630 3361 4664 3395
rect 4748 3361 4782 3395
rect 4866 3361 4900 3395
rect 4984 3361 5018 3395
rect 5102 3361 5136 3395
rect 5220 3361 5254 3395
rect 5338 3361 5372 3395
rect 5456 3361 5490 3395
rect 5574 3361 5608 3395
rect 5692 3361 5726 3395
rect 5810 3361 5844 3395
rect 5928 3361 5962 3395
rect 9214 3361 9248 3395
rect 9332 3361 9366 3395
rect 9450 3361 9484 3395
rect 9568 3361 9602 3395
rect 9686 3361 9720 3395
rect 9804 3361 9838 3395
rect 9922 3361 9956 3395
rect 10040 3361 10074 3395
rect 12908 38581 12942 38615
rect 13026 38581 13060 38615
rect 10412 3361 10446 3395
rect 10530 3361 10564 3395
rect 10648 3361 10682 3395
rect 10766 3361 10800 3395
rect 10884 3361 10918 3395
rect 11002 3361 11036 3395
rect 11120 3361 11154 3395
rect 11238 3361 11272 3395
rect 13398 38581 13432 38615
rect 13516 38581 13550 38615
rect 11610 291 11644 325
rect 11724 291 11758 325
rect 14696 291 14730 325
rect 14814 291 14848 325
<< mvpsubdiff >>
rect -252 38723 -142 38757
rect -108 38723 -74 38757
rect -40 38723 -6 38757
rect 28 38723 62 38757
rect 96 38723 130 38757
rect 164 38723 198 38757
rect 232 38723 266 38757
rect 300 38723 334 38757
rect 368 38723 402 38757
rect 436 38723 470 38757
rect 504 38723 538 38757
rect 572 38723 606 38757
rect 640 38723 674 38757
rect 708 38723 742 38757
rect 776 38723 810 38757
rect 844 38723 878 38757
rect 912 38723 946 38757
rect 980 38723 1014 38757
rect 1048 38723 1082 38757
rect 1116 38723 1150 38757
rect 1184 38723 1218 38757
rect 1252 38723 1286 38757
rect 1320 38723 1354 38757
rect 1388 38723 1422 38757
rect 1456 38723 1490 38757
rect 1524 38723 1558 38757
rect 1592 38723 1626 38757
rect 1660 38723 1694 38757
rect 1728 38723 1762 38757
rect 1796 38723 1898 38757
rect 1932 38723 1966 38757
rect 2000 38723 2034 38757
rect 2068 38723 2102 38757
rect 2136 38723 2170 38757
rect 2204 38723 2238 38757
rect 2272 38723 2306 38757
rect 2340 38723 2374 38757
rect 2408 38723 2442 38757
rect 2476 38723 2510 38757
rect 2544 38723 2578 38757
rect 2612 38723 2646 38757
rect 2680 38723 2714 38757
rect 2748 38723 2782 38757
rect 2816 38723 2850 38757
rect 2884 38723 2918 38757
rect 2952 38723 2986 38757
rect 3020 38723 3054 38757
rect 3088 38723 3122 38757
rect 3156 38723 3190 38757
rect 3224 38723 3258 38757
rect 3292 38723 3326 38757
rect 3360 38723 3394 38757
rect 3428 38723 3462 38757
rect 3496 38723 3530 38757
rect 3564 38723 3598 38757
rect 3632 38723 3666 38757
rect 3700 38723 3734 38757
rect 3768 38723 3802 38757
rect 3836 38723 3870 38757
rect 3904 38723 4074 38757
rect 4108 38723 4142 38757
rect 4176 38723 4210 38757
rect 4244 38723 4278 38757
rect 4312 38723 4346 38757
rect 4380 38723 4414 38757
rect 4448 38723 4482 38757
rect 4516 38723 4550 38757
rect 4584 38723 4618 38757
rect 4652 38723 4686 38757
rect 4720 38723 4754 38757
rect 4788 38723 4822 38757
rect 4856 38723 4890 38757
rect 4924 38723 4958 38757
rect 4992 38723 5026 38757
rect 5060 38723 5094 38757
rect 5128 38723 5162 38757
rect 5196 38723 5230 38757
rect 5264 38723 5298 38757
rect 5332 38723 5366 38757
rect 5400 38723 5434 38757
rect 5468 38723 5502 38757
rect 5536 38723 5570 38757
rect 5604 38723 5638 38757
rect 5672 38723 5706 38757
rect 5740 38723 5774 38757
rect 5808 38723 5842 38757
rect 5876 38723 5910 38757
rect 5944 38723 5978 38757
rect 6012 38723 6046 38757
rect 6080 38723 6148 38757
rect -252 38689 -218 38723
rect -252 38621 -218 38655
rect -252 38553 -218 38587
rect -252 38485 -218 38519
rect -252 38417 -218 38451
rect -252 38349 -218 38383
rect -252 38281 -218 38315
rect -252 38213 -218 38247
rect -252 38145 -218 38179
rect -252 38077 -218 38111
rect -252 38009 -218 38043
rect -252 37941 -218 37975
rect -252 37873 -218 37907
rect -252 37805 -218 37839
rect -252 37737 -218 37771
rect -252 37669 -218 37703
rect -252 37601 -218 37635
rect -252 37533 -218 37567
rect -252 37465 -218 37499
rect -252 37397 -218 37431
rect -252 37329 -218 37363
rect -252 37261 -218 37295
rect -252 37193 -218 37227
rect -252 37125 -218 37159
rect -252 37057 -218 37091
rect -252 36989 -218 37023
rect -252 36921 -218 36955
rect -252 36853 -218 36887
rect -252 36785 -218 36819
rect -252 36717 -218 36751
rect -252 36649 -218 36683
rect -252 36581 -218 36615
rect -252 36513 -218 36547
rect -252 36445 -218 36479
rect -252 36377 -218 36411
rect -252 36309 -218 36343
rect -252 36241 -218 36275
rect -252 36173 -218 36207
rect -252 36105 -218 36139
rect -252 36037 -218 36071
rect -252 35969 -218 36003
rect -252 35901 -218 35935
rect -252 35833 -218 35867
rect -252 35765 -218 35799
rect -252 35697 -218 35731
rect -252 35629 -218 35663
rect -252 35561 -218 35595
rect -252 35493 -218 35527
rect -252 35425 -218 35459
rect -252 35357 -218 35391
rect -252 35289 -218 35323
rect -252 35221 -218 35255
rect -252 35153 -218 35187
rect -252 35085 -218 35119
rect -252 35017 -218 35051
rect -252 34949 -218 34983
rect -252 34881 -218 34915
rect -252 34813 -218 34847
rect -252 34745 -218 34779
rect -252 34677 -218 34711
rect -252 34609 -218 34643
rect -252 34541 -218 34575
rect -252 34473 -218 34507
rect -252 34405 -218 34439
rect -252 34337 -218 34371
rect -252 34269 -218 34303
rect -252 34201 -218 34235
rect -252 34133 -218 34167
rect -252 34065 -218 34099
rect -252 33997 -218 34031
rect -252 33929 -218 33963
rect -252 33861 -218 33895
rect -252 33793 -218 33827
rect -252 33725 -218 33759
rect -252 33657 -218 33691
rect -252 33589 -218 33623
rect -252 33521 -218 33555
rect -252 33453 -218 33487
rect -252 33385 -218 33419
rect -252 33317 -218 33351
rect -252 33249 -218 33283
rect -252 33181 -218 33215
rect -252 33113 -218 33147
rect -252 33045 -218 33079
rect -252 32977 -218 33011
rect -252 32909 -218 32943
rect -252 32841 -218 32875
rect -252 32773 -218 32807
rect -252 32705 -218 32739
rect -252 32637 -218 32671
rect -252 32569 -218 32603
rect -252 32501 -218 32535
rect -252 32433 -218 32467
rect -252 32365 -218 32399
rect -252 32297 -218 32331
rect -252 32229 -218 32263
rect -252 32161 -218 32195
rect -252 32093 -218 32127
rect -252 32025 -218 32059
rect -252 31957 -218 31991
rect -252 31889 -218 31923
rect -252 31821 -218 31855
rect -252 31753 -218 31787
rect -252 31685 -218 31719
rect -252 31617 -218 31651
rect -252 31549 -218 31583
rect -252 31481 -218 31515
rect -252 31413 -218 31447
rect -252 31345 -218 31379
rect -252 31277 -218 31311
rect -252 31209 -218 31243
rect -252 31141 -218 31175
rect -252 31073 -218 31107
rect -252 31005 -218 31039
rect -252 30937 -218 30971
rect -252 30869 -218 30903
rect -252 30801 -218 30835
rect -252 30733 -218 30767
rect -252 30665 -218 30699
rect -252 30597 -218 30631
rect -252 30529 -218 30563
rect -252 30461 -218 30495
rect -252 30393 -218 30427
rect -252 30325 -218 30359
rect -252 30257 -218 30291
rect -252 30189 -218 30223
rect -252 30121 -218 30155
rect -252 30053 -218 30087
rect -252 29985 -218 30019
rect -252 29917 -218 29951
rect -252 29849 -218 29883
rect -252 29781 -218 29815
rect -252 29713 -218 29747
rect -252 29645 -218 29679
rect -252 29577 -218 29611
rect -252 29509 -218 29543
rect -252 29441 -218 29475
rect -252 29373 -218 29407
rect -252 29305 -218 29339
rect -252 29237 -218 29271
rect -252 29169 -218 29203
rect -252 29101 -218 29135
rect -252 29033 -218 29067
rect -252 28965 -218 28999
rect -252 28897 -218 28931
rect -252 28829 -218 28863
rect -252 28761 -218 28795
rect -252 28693 -218 28727
rect -252 28625 -218 28659
rect -252 28557 -218 28591
rect -252 28489 -218 28523
rect -252 28421 -218 28455
rect -252 28353 -218 28387
rect -252 28285 -218 28319
rect -252 28217 -218 28251
rect -252 28149 -218 28183
rect -252 28081 -218 28115
rect -252 28013 -218 28047
rect -252 27945 -218 27979
rect -252 27877 -218 27911
rect -252 27809 -218 27843
rect -252 27741 -218 27775
rect -252 27673 -218 27707
rect -252 27605 -218 27639
rect -252 27537 -218 27571
rect -252 27469 -218 27503
rect -252 27401 -218 27435
rect -252 27333 -218 27367
rect -252 27265 -218 27299
rect -252 27197 -218 27231
rect -252 27129 -218 27163
rect -252 27061 -218 27095
rect -252 26993 -218 27027
rect -252 26925 -218 26959
rect -252 26857 -218 26891
rect -252 26789 -218 26823
rect -252 26721 -218 26755
rect -252 26653 -218 26687
rect -252 26585 -218 26619
rect -252 26517 -218 26551
rect -252 26449 -218 26483
rect -252 26381 -218 26415
rect -252 26313 -218 26347
rect -252 26245 -218 26279
rect -252 26177 -218 26211
rect -252 26109 -218 26143
rect -252 26041 -218 26075
rect -252 25973 -218 26007
rect -252 25905 -218 25939
rect -252 25837 -218 25871
rect -252 25769 -218 25803
rect -252 25701 -218 25735
rect -252 25633 -218 25667
rect -252 25565 -218 25599
rect -252 25497 -218 25531
rect -252 25429 -218 25463
rect -252 25361 -218 25395
rect -252 25293 -218 25327
rect -252 25225 -218 25259
rect -252 25157 -218 25191
rect -252 25089 -218 25123
rect -252 25021 -218 25055
rect -252 24953 -218 24987
rect -252 24885 -218 24919
rect -252 24817 -218 24851
rect -252 24749 -218 24783
rect -252 24681 -218 24715
rect -252 24613 -218 24647
rect -252 24545 -218 24579
rect -252 24477 -218 24511
rect -252 24409 -218 24443
rect -252 24341 -218 24375
rect -252 24273 -218 24307
rect -252 24205 -218 24239
rect -252 24137 -218 24171
rect -252 24069 -218 24103
rect -252 24001 -218 24035
rect -252 23933 -218 23967
rect -252 23865 -218 23899
rect -252 23797 -218 23831
rect -252 23729 -218 23763
rect -252 23661 -218 23695
rect -252 23593 -218 23627
rect -252 23525 -218 23559
rect -252 23457 -218 23491
rect -252 23389 -218 23423
rect -252 23321 -218 23355
rect -252 23253 -218 23287
rect -252 23185 -218 23219
rect -252 23117 -218 23151
rect -252 23049 -218 23083
rect -252 22981 -218 23015
rect -252 22913 -218 22947
rect -252 22845 -218 22879
rect -252 22777 -218 22811
rect -252 22709 -218 22743
rect -252 22641 -218 22675
rect -252 22573 -218 22607
rect -252 22505 -218 22539
rect -252 22437 -218 22471
rect -252 22369 -218 22403
rect -252 22301 -218 22335
rect -252 22233 -218 22267
rect -252 22165 -218 22199
rect -252 22097 -218 22131
rect -252 22029 -218 22063
rect -252 21961 -218 21995
rect -252 21893 -218 21927
rect -252 21825 -218 21859
rect -252 21757 -218 21791
rect -252 21689 -218 21723
rect -252 21621 -218 21655
rect -252 21553 -218 21587
rect -252 21485 -218 21519
rect -252 21417 -218 21451
rect -252 21349 -218 21383
rect -252 21281 -218 21315
rect -252 21213 -218 21247
rect -252 21145 -218 21179
rect -252 21077 -218 21111
rect -252 21009 -218 21043
rect -252 20941 -218 20975
rect -252 20873 -218 20907
rect -252 20805 -218 20839
rect -252 20737 -218 20771
rect -252 20669 -218 20703
rect -252 20601 -218 20635
rect -252 20533 -218 20567
rect -252 20465 -218 20499
rect -252 20397 -218 20431
rect -252 20329 -218 20363
rect -252 20261 -218 20295
rect -252 20193 -218 20227
rect -252 20125 -218 20159
rect -252 20057 -218 20091
rect -252 19989 -218 20023
rect -252 19921 -218 19955
rect -252 19853 -218 19887
rect -252 19785 -218 19819
rect -252 19717 -218 19751
rect -252 19649 -218 19683
rect -252 19581 -218 19615
rect -252 19513 -218 19547
rect -252 19445 -218 19479
rect -252 19377 -218 19411
rect -252 19309 -218 19343
rect -252 19241 -218 19275
rect -252 19173 -218 19207
rect -252 19105 -218 19139
rect -252 19037 -218 19071
rect -252 18969 -218 19003
rect -252 18901 -218 18935
rect -252 18833 -218 18867
rect -252 18765 -218 18799
rect -252 18697 -218 18731
rect -252 18629 -218 18663
rect -252 18561 -218 18595
rect -252 18493 -218 18527
rect -252 18425 -218 18459
rect -252 18357 -218 18391
rect -252 18289 -218 18323
rect -252 18221 -218 18255
rect -252 18153 -218 18187
rect -252 18085 -218 18119
rect -252 18017 -218 18051
rect -252 17949 -218 17983
rect -252 17881 -218 17915
rect -252 17813 -218 17847
rect -252 17745 -218 17779
rect -252 17677 -218 17711
rect -252 17609 -218 17643
rect -252 17541 -218 17575
rect -252 17473 -218 17507
rect -252 17405 -218 17439
rect -252 17337 -218 17371
rect -252 17269 -218 17303
rect -252 17201 -218 17235
rect -252 17133 -218 17167
rect -252 17065 -218 17099
rect -252 16997 -218 17031
rect -252 16929 -218 16963
rect -252 16861 -218 16895
rect -252 16793 -218 16827
rect -252 16725 -218 16759
rect -252 16657 -218 16691
rect -252 16589 -218 16623
rect -252 16521 -218 16555
rect -252 16453 -218 16487
rect -252 16385 -218 16419
rect -252 16317 -218 16351
rect -252 16249 -218 16283
rect -252 16181 -218 16215
rect -252 16113 -218 16147
rect -252 16045 -218 16079
rect -252 15977 -218 16011
rect -252 15909 -218 15943
rect -252 15841 -218 15875
rect -252 15773 -218 15807
rect -252 15705 -218 15739
rect -252 15637 -218 15671
rect -252 15569 -218 15603
rect -252 15501 -218 15535
rect -252 15433 -218 15467
rect -252 15365 -218 15399
rect -252 15297 -218 15331
rect -252 15229 -218 15263
rect -252 15161 -218 15195
rect -252 15093 -218 15127
rect -252 15025 -218 15059
rect -252 14957 -218 14991
rect -252 14889 -218 14923
rect -252 14821 -218 14855
rect -252 14753 -218 14787
rect -252 14685 -218 14719
rect -252 14617 -218 14651
rect -252 14549 -218 14583
rect -252 14481 -218 14515
rect -252 14413 -218 14447
rect -252 14345 -218 14379
rect -252 14277 -218 14311
rect -252 14209 -218 14243
rect -252 14141 -218 14175
rect -252 14073 -218 14107
rect -252 14005 -218 14039
rect -252 13937 -218 13971
rect -252 13869 -218 13903
rect -252 13801 -218 13835
rect -252 13733 -218 13767
rect -252 13665 -218 13699
rect -252 13597 -218 13631
rect -252 13529 -218 13563
rect -252 13461 -218 13495
rect -252 13393 -218 13427
rect -252 13325 -218 13359
rect -252 13257 -218 13291
rect -252 13189 -218 13223
rect -252 13121 -218 13155
rect -252 13053 -218 13087
rect -252 12985 -218 13019
rect -252 12917 -218 12951
rect -252 12849 -218 12883
rect -252 12781 -218 12815
rect -252 12713 -218 12747
rect -252 12645 -218 12679
rect -252 12577 -218 12611
rect -252 12509 -218 12543
rect -252 12441 -218 12475
rect -252 12373 -218 12407
rect -252 12305 -218 12339
rect -252 12237 -218 12271
rect -252 12169 -218 12203
rect -252 12101 -218 12135
rect -252 12033 -218 12067
rect -252 11965 -218 11999
rect -252 11897 -218 11931
rect -252 11829 -218 11863
rect -252 11761 -218 11795
rect -252 11693 -218 11727
rect -252 11625 -218 11659
rect -252 11557 -218 11591
rect -252 11489 -218 11523
rect -252 11421 -218 11455
rect -252 11353 -218 11387
rect -252 11285 -218 11319
rect -252 11217 -218 11251
rect -252 11149 -218 11183
rect -252 11081 -218 11115
rect -252 11013 -218 11047
rect -252 10945 -218 10979
rect -252 10877 -218 10911
rect -252 10809 -218 10843
rect -252 10741 -218 10775
rect -252 10673 -218 10707
rect -252 10605 -218 10639
rect -252 10537 -218 10571
rect -252 10469 -218 10503
rect -252 10401 -218 10435
rect -252 10333 -218 10367
rect -252 10265 -218 10299
rect -252 10197 -218 10231
rect -252 10129 -218 10163
rect -252 10061 -218 10095
rect -252 9993 -218 10027
rect -252 9925 -218 9959
rect -252 9857 -218 9891
rect -252 9789 -218 9823
rect -252 9721 -218 9755
rect -252 9653 -218 9687
rect -252 9585 -218 9619
rect -252 9517 -218 9551
rect -252 9449 -218 9483
rect -252 9381 -218 9415
rect -252 9313 -218 9347
rect -252 9245 -218 9279
rect -252 9177 -218 9211
rect -252 9109 -218 9143
rect -252 9041 -218 9075
rect -252 8973 -218 9007
rect -252 8905 -218 8939
rect -252 8837 -218 8871
rect -252 8769 -218 8803
rect -252 8701 -218 8735
rect -252 8633 -218 8667
rect -252 8565 -218 8599
rect -252 8497 -218 8531
rect -252 8429 -218 8463
rect -252 8361 -218 8395
rect -252 8293 -218 8327
rect -252 8225 -218 8259
rect -252 8157 -218 8191
rect -252 8089 -218 8123
rect -252 8021 -218 8055
rect -252 7953 -218 7987
rect -252 7885 -218 7919
rect -252 7817 -218 7851
rect -252 7749 -218 7783
rect -252 7681 -218 7715
rect -252 7613 -218 7647
rect -252 7545 -218 7579
rect -252 7477 -218 7511
rect -252 7409 -218 7443
rect -252 7341 -218 7375
rect -252 7273 -218 7307
rect -252 7205 -218 7239
rect -252 7137 -218 7171
rect -252 7069 -218 7103
rect -252 7001 -218 7035
rect -252 6933 -218 6967
rect -252 6865 -218 6899
rect -252 6797 -218 6831
rect -252 6729 -218 6763
rect -252 6661 -218 6695
rect -252 6593 -218 6627
rect -252 6525 -218 6559
rect -252 6457 -218 6491
rect -252 6389 -218 6423
rect -252 6321 -218 6355
rect -252 6253 -218 6287
rect -252 6185 -218 6219
rect -252 6117 -218 6151
rect -252 6049 -218 6083
rect -252 5981 -218 6015
rect -252 5913 -218 5947
rect -252 5845 -218 5879
rect -252 5777 -218 5811
rect -252 5709 -218 5743
rect -252 5641 -218 5675
rect -252 5573 -218 5607
rect -252 5505 -218 5539
rect -252 5437 -218 5471
rect -252 5369 -218 5403
rect -252 5301 -218 5335
rect -252 5233 -218 5267
rect -252 5165 -218 5199
rect -252 5097 -218 5131
rect -252 5029 -218 5063
rect -252 4961 -218 4995
rect -252 4893 -218 4927
rect -252 4825 -218 4859
rect -252 4757 -218 4791
rect -252 4689 -218 4723
rect -252 4621 -218 4655
rect -252 4553 -218 4587
rect -252 4485 -218 4519
rect -252 4417 -218 4451
rect -252 4349 -218 4383
rect -252 4281 -218 4315
rect -252 4213 -218 4247
rect -252 4145 -218 4179
rect -252 4077 -218 4111
rect -252 4009 -218 4043
rect -252 3941 -218 3975
rect -252 3873 -218 3907
rect -252 3805 -218 3839
rect -252 3737 -218 3771
rect -252 3669 -218 3703
rect -252 3601 -218 3635
rect -252 3533 -218 3567
rect -252 3465 -218 3499
rect 1830 38641 1864 38723
rect 1830 38573 1864 38607
rect 1830 38505 1864 38539
rect 1830 38437 1864 38471
rect 1830 38369 1864 38403
rect 1830 38301 1864 38335
rect 1830 38233 1864 38267
rect 1830 38165 1864 38199
rect 1830 38097 1864 38131
rect 1830 38029 1864 38063
rect 1830 37961 1864 37995
rect 1830 37893 1864 37927
rect 1830 37825 1864 37859
rect 1830 37757 1864 37791
rect 1830 37689 1864 37723
rect 1830 37621 1864 37655
rect 1830 37553 1864 37587
rect 1830 37485 1864 37519
rect 1830 37417 1864 37451
rect 1830 37349 1864 37383
rect 1830 37281 1864 37315
rect 1830 37213 1864 37247
rect 1830 37145 1864 37179
rect 1830 37077 1864 37111
rect 1830 37009 1864 37043
rect 1830 36941 1864 36975
rect 1830 36873 1864 36907
rect 1830 36805 1864 36839
rect 1830 36737 1864 36771
rect 1830 36669 1864 36703
rect 1830 36601 1864 36635
rect 1830 36533 1864 36567
rect 1830 36465 1864 36499
rect 1830 36397 1864 36431
rect 1830 36329 1864 36363
rect 1830 36261 1864 36295
rect 1830 36193 1864 36227
rect 1830 36125 1864 36159
rect 1830 36057 1864 36091
rect 1830 35989 1864 36023
rect 1830 35921 1864 35955
rect 1830 35853 1864 35887
rect 1830 35785 1864 35819
rect 1830 35717 1864 35751
rect 1830 35649 1864 35683
rect 1830 35581 1864 35615
rect 1830 35513 1864 35547
rect 1830 35445 1864 35479
rect 1830 35377 1864 35411
rect 1830 35309 1864 35343
rect 1830 35241 1864 35275
rect 1830 35173 1864 35207
rect 1830 35105 1864 35139
rect 1830 35037 1864 35071
rect 1830 34969 1864 35003
rect 1830 34901 1864 34935
rect 1830 34833 1864 34867
rect 1830 34765 1864 34799
rect 1830 34697 1864 34731
rect 1830 34629 1864 34663
rect 1830 34561 1864 34595
rect 1830 34493 1864 34527
rect 1830 34425 1864 34459
rect 1830 34357 1864 34391
rect 1830 34289 1864 34323
rect 1830 34221 1864 34255
rect 1830 34153 1864 34187
rect 1830 34085 1864 34119
rect 1830 34017 1864 34051
rect 1830 33949 1864 33983
rect 1830 33881 1864 33915
rect 1830 33813 1864 33847
rect 1830 33745 1864 33779
rect 1830 33677 1864 33711
rect 1830 33609 1864 33643
rect 1830 33541 1864 33575
rect 1830 33473 1864 33507
rect 1830 33405 1864 33439
rect 1830 33337 1864 33371
rect 1830 33269 1864 33303
rect 1830 33201 1864 33235
rect 1830 33133 1864 33167
rect 1830 33065 1864 33099
rect 1830 32997 1864 33031
rect 1830 32929 1864 32963
rect 1830 32861 1864 32895
rect 1830 32793 1864 32827
rect 1830 32725 1864 32759
rect 1830 32657 1864 32691
rect 1830 32589 1864 32623
rect 1830 32521 1864 32555
rect 1830 32453 1864 32487
rect 1830 32385 1864 32419
rect 1830 32317 1864 32351
rect 1830 32249 1864 32283
rect 1830 32181 1864 32215
rect 1830 32113 1864 32147
rect 1830 32045 1864 32079
rect 1830 31977 1864 32011
rect 1830 31909 1864 31943
rect 1830 31841 1864 31875
rect 1830 31773 1864 31807
rect 1830 31705 1864 31739
rect 1830 31637 1864 31671
rect 1830 31569 1864 31603
rect 1830 31501 1864 31535
rect 1830 31433 1864 31467
rect 1830 31365 1864 31399
rect 1830 31297 1864 31331
rect 1830 31229 1864 31263
rect 1830 31161 1864 31195
rect 1830 31093 1864 31127
rect 1830 31025 1864 31059
rect 1830 30957 1864 30991
rect 1830 30889 1864 30923
rect 1830 30821 1864 30855
rect 1830 30753 1864 30787
rect 1830 30685 1864 30719
rect 1830 30617 1864 30651
rect 1830 30549 1864 30583
rect 1830 30481 1864 30515
rect 1830 30413 1864 30447
rect 1830 30345 1864 30379
rect 1830 30277 1864 30311
rect 1830 30209 1864 30243
rect 1830 30141 1864 30175
rect 1830 30073 1864 30107
rect 1830 30005 1864 30039
rect 1830 29937 1864 29971
rect 1830 29869 1864 29903
rect 1830 29801 1864 29835
rect 1830 29733 1864 29767
rect 1830 29665 1864 29699
rect 1830 29597 1864 29631
rect 1830 29529 1864 29563
rect 1830 29461 1864 29495
rect 1830 29393 1864 29427
rect 1830 29325 1864 29359
rect 1830 29257 1864 29291
rect 1830 29189 1864 29223
rect 1830 29121 1864 29155
rect 1830 29053 1864 29087
rect 1830 28985 1864 29019
rect 1830 28917 1864 28951
rect 1830 28849 1864 28883
rect 1830 28781 1864 28815
rect 1830 28713 1864 28747
rect 1830 28645 1864 28679
rect 1830 28577 1864 28611
rect 1830 28509 1864 28543
rect 1830 28441 1864 28475
rect 1830 28373 1864 28407
rect 1830 28305 1864 28339
rect 1830 28237 1864 28271
rect 1830 28169 1864 28203
rect 1830 28101 1864 28135
rect 1830 28033 1864 28067
rect 1830 27965 1864 27999
rect 1830 27897 1864 27931
rect 1830 27829 1864 27863
rect 1830 27761 1864 27795
rect 1830 27693 1864 27727
rect 1830 27625 1864 27659
rect 1830 27557 1864 27591
rect 1830 27489 1864 27523
rect 1830 27421 1864 27455
rect 1830 27353 1864 27387
rect 1830 27285 1864 27319
rect 1830 27217 1864 27251
rect 1830 27149 1864 27183
rect 1830 27081 1864 27115
rect 1830 27013 1864 27047
rect 1830 26945 1864 26979
rect 1830 26877 1864 26911
rect 1830 26809 1864 26843
rect 1830 26741 1864 26775
rect 1830 26673 1864 26707
rect 1830 26605 1864 26639
rect 1830 26537 1864 26571
rect 1830 26469 1864 26503
rect 1830 26401 1864 26435
rect 1830 26333 1864 26367
rect 1830 26265 1864 26299
rect 1830 26197 1864 26231
rect 1830 26129 1864 26163
rect 1830 26061 1864 26095
rect 1830 25993 1864 26027
rect 1830 25925 1864 25959
rect 1830 25857 1864 25891
rect 1830 25789 1864 25823
rect 1830 25721 1864 25755
rect 1830 25653 1864 25687
rect 1830 25585 1864 25619
rect 1830 25517 1864 25551
rect 1830 25449 1864 25483
rect 1830 25381 1864 25415
rect 1830 25313 1864 25347
rect 1830 25245 1864 25279
rect 1830 25177 1864 25211
rect 1830 25109 1864 25143
rect 1830 25041 1864 25075
rect 1830 24973 1864 25007
rect 1830 24905 1864 24939
rect 1830 24837 1864 24871
rect 1830 24769 1864 24803
rect 1830 24701 1864 24735
rect 1830 24633 1864 24667
rect 1830 24565 1864 24599
rect 1830 24497 1864 24531
rect 1830 24429 1864 24463
rect 1830 24361 1864 24395
rect 1830 24293 1864 24327
rect 1830 24225 1864 24259
rect 1830 24157 1864 24191
rect 1830 24089 1864 24123
rect 1830 24021 1864 24055
rect 1830 23953 1864 23987
rect 1830 23885 1864 23919
rect 1830 23817 1864 23851
rect 1830 23749 1864 23783
rect 1830 23681 1864 23715
rect 1830 23613 1864 23647
rect 1830 23545 1864 23579
rect 1830 23477 1864 23511
rect 1830 23409 1864 23443
rect 1830 23341 1864 23375
rect 1830 23273 1864 23307
rect 1830 23205 1864 23239
rect 1830 23137 1864 23171
rect 1830 23069 1864 23103
rect 1830 23001 1864 23035
rect 1830 22933 1864 22967
rect 1830 22865 1864 22899
rect 1830 22797 1864 22831
rect 1830 22729 1864 22763
rect 1830 22661 1864 22695
rect 1830 22593 1864 22627
rect 1830 22525 1864 22559
rect 1830 22457 1864 22491
rect 1830 22389 1864 22423
rect 1830 22321 1864 22355
rect 1830 22253 1864 22287
rect 1830 22185 1864 22219
rect 1830 22117 1864 22151
rect 1830 22049 1864 22083
rect 1830 21981 1864 22015
rect 1830 21913 1864 21947
rect 1830 21845 1864 21879
rect 1830 21777 1864 21811
rect 1830 21709 1864 21743
rect 1830 21641 1864 21675
rect 1830 21573 1864 21607
rect 1830 21505 1864 21539
rect 1830 21437 1864 21471
rect 1830 21369 1864 21403
rect 1830 21301 1864 21335
rect 1830 21233 1864 21267
rect 1830 21165 1864 21199
rect 1830 21097 1864 21131
rect 1830 21029 1864 21063
rect 1830 20961 1864 20995
rect 1830 20893 1864 20927
rect 1830 20825 1864 20859
rect 1830 20757 1864 20791
rect 1830 20689 1864 20723
rect 1830 20621 1864 20655
rect 1830 20553 1864 20587
rect 1830 20485 1864 20519
rect 1830 20417 1864 20451
rect 1830 20349 1864 20383
rect 1830 20281 1864 20315
rect 1830 20213 1864 20247
rect 1830 20145 1864 20179
rect 1830 20077 1864 20111
rect 1830 20009 1864 20043
rect 1830 19941 1864 19975
rect 1830 19873 1864 19907
rect 1830 19805 1864 19839
rect 1830 19737 1864 19771
rect 1830 19669 1864 19703
rect 1830 19601 1864 19635
rect 1830 19533 1864 19567
rect 1830 19465 1864 19499
rect 1830 19397 1864 19431
rect 1830 19329 1864 19363
rect 1830 19261 1864 19295
rect 1830 19193 1864 19227
rect 1830 19125 1864 19159
rect 1830 19057 1864 19091
rect 1830 18989 1864 19023
rect 1830 18921 1864 18955
rect 1830 18853 1864 18887
rect 1830 18785 1864 18819
rect 1830 18717 1864 18751
rect 1830 18649 1864 18683
rect 1830 18581 1864 18615
rect 1830 18513 1864 18547
rect 1830 18445 1864 18479
rect 1830 18377 1864 18411
rect 1830 18309 1864 18343
rect 1830 18241 1864 18275
rect 1830 18173 1864 18207
rect 1830 18105 1864 18139
rect 1830 18037 1864 18071
rect 1830 17969 1864 18003
rect 1830 17901 1864 17935
rect 1830 17833 1864 17867
rect 1830 17765 1864 17799
rect 1830 17697 1864 17731
rect 1830 17629 1864 17663
rect 1830 17561 1864 17595
rect 1830 17493 1864 17527
rect 1830 17425 1864 17459
rect 1830 17357 1864 17391
rect 1830 17289 1864 17323
rect 1830 17221 1864 17255
rect 1830 17153 1864 17187
rect 1830 17085 1864 17119
rect 1830 17017 1864 17051
rect 1830 16949 1864 16983
rect 1830 16881 1864 16915
rect 1830 16813 1864 16847
rect 1830 16745 1864 16779
rect 1830 16677 1864 16711
rect 1830 16609 1864 16643
rect 1830 16541 1864 16575
rect 1830 16473 1864 16507
rect 1830 16405 1864 16439
rect 1830 16337 1864 16371
rect 1830 16269 1864 16303
rect 1830 16201 1864 16235
rect 1830 16133 1864 16167
rect 1830 16065 1864 16099
rect 1830 15997 1864 16031
rect 1830 15929 1864 15963
rect 1830 15861 1864 15895
rect 1830 15793 1864 15827
rect 1830 15725 1864 15759
rect 1830 15657 1864 15691
rect 1830 15589 1864 15623
rect 1830 15521 1864 15555
rect 1830 15453 1864 15487
rect 1830 15385 1864 15419
rect 1830 15317 1864 15351
rect 1830 15249 1864 15283
rect 1830 15181 1864 15215
rect 1830 15113 1864 15147
rect 1830 15045 1864 15079
rect 1830 14977 1864 15011
rect 1830 14909 1864 14943
rect 1830 14841 1864 14875
rect 1830 14773 1864 14807
rect 1830 14705 1864 14739
rect 1830 14637 1864 14671
rect 1830 14569 1864 14603
rect 1830 14501 1864 14535
rect 1830 14433 1864 14467
rect 1830 14365 1864 14399
rect 1830 14297 1864 14331
rect 1830 14229 1864 14263
rect 1830 14161 1864 14195
rect 1830 14093 1864 14127
rect 1830 14025 1864 14059
rect 1830 13957 1864 13991
rect 1830 13889 1864 13923
rect 1830 13821 1864 13855
rect 1830 13753 1864 13787
rect 1830 13685 1864 13719
rect 1830 13617 1864 13651
rect 1830 13549 1864 13583
rect 1830 13481 1864 13515
rect 1830 13413 1864 13447
rect 1830 13345 1864 13379
rect 1830 13277 1864 13311
rect 1830 13209 1864 13243
rect 1830 13141 1864 13175
rect 1830 13073 1864 13107
rect 1830 13005 1864 13039
rect 1830 12937 1864 12971
rect 1830 12869 1864 12903
rect 1830 12801 1864 12835
rect 1830 12733 1864 12767
rect 1830 12665 1864 12699
rect 1830 12597 1864 12631
rect 1830 12529 1864 12563
rect 1830 12461 1864 12495
rect 1830 12393 1864 12427
rect 1830 12325 1864 12359
rect 1830 12257 1864 12291
rect 1830 12189 1864 12223
rect 1830 12121 1864 12155
rect 1830 12053 1864 12087
rect 1830 11985 1864 12019
rect 1830 11917 1864 11951
rect 1830 11849 1864 11883
rect 1830 11781 1864 11815
rect 1830 11713 1864 11747
rect 1830 11645 1864 11679
rect 1830 11577 1864 11611
rect 1830 11509 1864 11543
rect 1830 11441 1864 11475
rect 1830 11373 1864 11407
rect 1830 11305 1864 11339
rect 1830 11237 1864 11271
rect 1830 11169 1864 11203
rect 1830 11101 1864 11135
rect 1830 11033 1864 11067
rect 1830 10965 1864 10999
rect 1830 10897 1864 10931
rect 1830 10829 1864 10863
rect 1830 10761 1864 10795
rect 1830 10693 1864 10727
rect 1830 10625 1864 10659
rect 1830 10557 1864 10591
rect 1830 10489 1864 10523
rect 1830 10421 1864 10455
rect 1830 10353 1864 10387
rect 1830 10285 1864 10319
rect 1830 10217 1864 10251
rect 1830 10149 1864 10183
rect 1830 10081 1864 10115
rect 1830 10013 1864 10047
rect 1830 9945 1864 9979
rect 1830 9877 1864 9911
rect 1830 9809 1864 9843
rect 1830 9741 1864 9775
rect 1830 9673 1864 9707
rect 1830 9605 1864 9639
rect 1830 9537 1864 9571
rect 1830 9469 1864 9503
rect 1830 9401 1864 9435
rect 1830 9333 1864 9367
rect 1830 9265 1864 9299
rect 1830 9197 1864 9231
rect 1830 9129 1864 9163
rect 1830 9061 1864 9095
rect 1830 8993 1864 9027
rect 1830 8925 1864 8959
rect 1830 8857 1864 8891
rect 1830 8789 1864 8823
rect 1830 8721 1864 8755
rect 1830 8653 1864 8687
rect 1830 8585 1864 8619
rect 1830 8517 1864 8551
rect 1830 8449 1864 8483
rect 1830 8381 1864 8415
rect 1830 8313 1864 8347
rect 1830 8245 1864 8279
rect 1830 8177 1864 8211
rect 1830 8109 1864 8143
rect 1830 8041 1864 8075
rect 1830 7973 1864 8007
rect 1830 7905 1864 7939
rect 1830 7837 1864 7871
rect 1830 7769 1864 7803
rect 1830 7701 1864 7735
rect 1830 7633 1864 7667
rect 1830 7565 1864 7599
rect 1830 7497 1864 7531
rect 1830 7429 1864 7463
rect 1830 7361 1864 7395
rect 1830 7293 1864 7327
rect 1830 7225 1864 7259
rect 1830 7157 1864 7191
rect 1830 7089 1864 7123
rect 1830 7021 1864 7055
rect 1830 6953 1864 6987
rect 1830 6885 1864 6919
rect 1830 6817 1864 6851
rect 1830 6749 1864 6783
rect 1830 6681 1864 6715
rect 1830 6613 1864 6647
rect 1830 6545 1864 6579
rect 1830 6477 1864 6511
rect 1830 6409 1864 6443
rect 1830 6341 1864 6375
rect 1830 6273 1864 6307
rect 1830 6205 1864 6239
rect 1830 6137 1864 6171
rect 1830 6069 1864 6103
rect 1830 6001 1864 6035
rect 1830 5933 1864 5967
rect 1830 5865 1864 5899
rect 1830 5797 1864 5831
rect 1830 5729 1864 5763
rect 1830 5661 1864 5695
rect 1830 5593 1864 5627
rect 1830 5525 1864 5559
rect 1830 5457 1864 5491
rect 1830 5389 1864 5423
rect 1830 5321 1864 5355
rect 1830 5253 1864 5287
rect 1830 5185 1864 5219
rect 1830 5117 1864 5151
rect 1830 5049 1864 5083
rect 1830 4981 1864 5015
rect 1830 4913 1864 4947
rect 1830 4845 1864 4879
rect 1830 4777 1864 4811
rect 1830 4709 1864 4743
rect 1830 4641 1864 4675
rect 1830 4573 1864 4607
rect 1830 4505 1864 4539
rect 1830 4437 1864 4471
rect 1830 4369 1864 4403
rect 1830 4301 1864 4335
rect 1830 4233 1864 4267
rect 1830 4165 1864 4199
rect 1830 4097 1864 4131
rect 1830 4029 1864 4063
rect 1830 3961 1864 3995
rect 1830 3893 1864 3927
rect 1830 3825 1864 3859
rect 1830 3757 1864 3791
rect 1830 3689 1864 3723
rect 1830 3621 1864 3655
rect 1830 3553 1864 3587
rect 1830 3485 1864 3519
rect -252 3397 -218 3431
rect -252 3329 -218 3363
rect 3972 38689 4006 38723
rect 3972 38621 4006 38655
rect 3972 38553 4006 38587
rect 3972 38485 4006 38519
rect 3972 38417 4006 38451
rect 3972 38349 4006 38383
rect 3972 38281 4006 38315
rect 3972 38213 4006 38247
rect 3972 38145 4006 38179
rect 3972 38077 4006 38111
rect 3972 38009 4006 38043
rect 3972 37941 4006 37975
rect 3972 37873 4006 37907
rect 3972 37805 4006 37839
rect 3972 37737 4006 37771
rect 3972 37669 4006 37703
rect 3972 37601 4006 37635
rect 3972 37533 4006 37567
rect 3972 37465 4006 37499
rect 3972 37397 4006 37431
rect 3972 37329 4006 37363
rect 3972 37261 4006 37295
rect 3972 37193 4006 37227
rect 3972 37125 4006 37159
rect 3972 37057 4006 37091
rect 3972 36989 4006 37023
rect 3972 36921 4006 36955
rect 3972 36853 4006 36887
rect 3972 36785 4006 36819
rect 3972 36717 4006 36751
rect 3972 36649 4006 36683
rect 3972 36581 4006 36615
rect 3972 36513 4006 36547
rect 3972 36445 4006 36479
rect 3972 36377 4006 36411
rect 3972 36309 4006 36343
rect 3972 36241 4006 36275
rect 3972 36173 4006 36207
rect 3972 36105 4006 36139
rect 3972 36037 4006 36071
rect 3972 35969 4006 36003
rect 3972 35901 4006 35935
rect 3972 35833 4006 35867
rect 3972 35765 4006 35799
rect 3972 35697 4006 35731
rect 3972 35629 4006 35663
rect 3972 35561 4006 35595
rect 3972 35493 4006 35527
rect 3972 35425 4006 35459
rect 3972 35357 4006 35391
rect 3972 35289 4006 35323
rect 3972 35221 4006 35255
rect 3972 35153 4006 35187
rect 3972 35085 4006 35119
rect 3972 35017 4006 35051
rect 3972 34949 4006 34983
rect 3972 34881 4006 34915
rect 3972 34813 4006 34847
rect 3972 34745 4006 34779
rect 3972 34677 4006 34711
rect 3972 34609 4006 34643
rect 3972 34541 4006 34575
rect 3972 34473 4006 34507
rect 3972 34405 4006 34439
rect 3972 34337 4006 34371
rect 3972 34269 4006 34303
rect 3972 34201 4006 34235
rect 3972 34133 4006 34167
rect 3972 34065 4006 34099
rect 3972 33997 4006 34031
rect 3972 33929 4006 33963
rect 3972 33861 4006 33895
rect 3972 33793 4006 33827
rect 3972 33725 4006 33759
rect 3972 33657 4006 33691
rect 3972 33589 4006 33623
rect 3972 33521 4006 33555
rect 3972 33453 4006 33487
rect 3972 33385 4006 33419
rect 3972 33317 4006 33351
rect 3972 33249 4006 33283
rect 3972 33181 4006 33215
rect 3972 33113 4006 33147
rect 3972 33045 4006 33079
rect 3972 32977 4006 33011
rect 3972 32909 4006 32943
rect 3972 32841 4006 32875
rect 3972 32773 4006 32807
rect 3972 32705 4006 32739
rect 3972 32637 4006 32671
rect 3972 32569 4006 32603
rect 3972 32501 4006 32535
rect 3972 32433 4006 32467
rect 3972 32365 4006 32399
rect 3972 32297 4006 32331
rect 3972 32229 4006 32263
rect 3972 32161 4006 32195
rect 3972 32093 4006 32127
rect 3972 32025 4006 32059
rect 3972 31957 4006 31991
rect 3972 31889 4006 31923
rect 3972 31821 4006 31855
rect 3972 31753 4006 31787
rect 3972 31685 4006 31719
rect 3972 31617 4006 31651
rect 3972 31549 4006 31583
rect 3972 31481 4006 31515
rect 3972 31413 4006 31447
rect 3972 31345 4006 31379
rect 3972 31277 4006 31311
rect 3972 31209 4006 31243
rect 3972 31141 4006 31175
rect 3972 31073 4006 31107
rect 3972 31005 4006 31039
rect 3972 30937 4006 30971
rect 3972 30869 4006 30903
rect 3972 30801 4006 30835
rect 3972 30733 4006 30767
rect 3972 30665 4006 30699
rect 3972 30597 4006 30631
rect 3972 30529 4006 30563
rect 3972 30461 4006 30495
rect 3972 30393 4006 30427
rect 3972 30325 4006 30359
rect 3972 30257 4006 30291
rect 3972 30189 4006 30223
rect 3972 30121 4006 30155
rect 3972 30053 4006 30087
rect 3972 29985 4006 30019
rect 3972 29917 4006 29951
rect 3972 29849 4006 29883
rect 3972 29781 4006 29815
rect 3972 29713 4006 29747
rect 3972 29645 4006 29679
rect 3972 29577 4006 29611
rect 3972 29509 4006 29543
rect 3972 29441 4006 29475
rect 3972 29373 4006 29407
rect 3972 29305 4006 29339
rect 3972 29237 4006 29271
rect 3972 29169 4006 29203
rect 3972 29101 4006 29135
rect 3972 29033 4006 29067
rect 3972 28965 4006 28999
rect 3972 28897 4006 28931
rect 3972 28829 4006 28863
rect 3972 28761 4006 28795
rect 3972 28693 4006 28727
rect 3972 28625 4006 28659
rect 3972 28557 4006 28591
rect 3972 28489 4006 28523
rect 3972 28421 4006 28455
rect 3972 28353 4006 28387
rect 3972 28285 4006 28319
rect 3972 28217 4006 28251
rect 3972 28149 4006 28183
rect 3972 28081 4006 28115
rect 3972 28013 4006 28047
rect 3972 27945 4006 27979
rect 3972 27877 4006 27911
rect 3972 27809 4006 27843
rect 3972 27741 4006 27775
rect 3972 27673 4006 27707
rect 3972 27605 4006 27639
rect 3972 27537 4006 27571
rect 3972 27469 4006 27503
rect 3972 27401 4006 27435
rect 3972 27333 4006 27367
rect 3972 27265 4006 27299
rect 3972 27197 4006 27231
rect 3972 27129 4006 27163
rect 3972 27061 4006 27095
rect 3972 26993 4006 27027
rect 3972 26925 4006 26959
rect 3972 26857 4006 26891
rect 3972 26789 4006 26823
rect 3972 26721 4006 26755
rect 3972 26653 4006 26687
rect 3972 26585 4006 26619
rect 3972 26517 4006 26551
rect 3972 26449 4006 26483
rect 3972 26381 4006 26415
rect 3972 26313 4006 26347
rect 3972 26245 4006 26279
rect 3972 26177 4006 26211
rect 3972 26109 4006 26143
rect 3972 26041 4006 26075
rect 3972 25973 4006 26007
rect 3972 25905 4006 25939
rect 3972 25837 4006 25871
rect 3972 25769 4006 25803
rect 3972 25701 4006 25735
rect 3972 25633 4006 25667
rect 3972 25565 4006 25599
rect 3972 25497 4006 25531
rect 3972 25429 4006 25463
rect 3972 25361 4006 25395
rect 3972 25293 4006 25327
rect 3972 25225 4006 25259
rect 3972 25157 4006 25191
rect 3972 25089 4006 25123
rect 3972 25021 4006 25055
rect 3972 24953 4006 24987
rect 3972 24885 4006 24919
rect 3972 24817 4006 24851
rect 3972 24749 4006 24783
rect 3972 24681 4006 24715
rect 3972 24613 4006 24647
rect 3972 24545 4006 24579
rect 3972 24477 4006 24511
rect 3972 24409 4006 24443
rect 3972 24341 4006 24375
rect 3972 24273 4006 24307
rect 3972 24205 4006 24239
rect 3972 24137 4006 24171
rect 3972 24069 4006 24103
rect 3972 24001 4006 24035
rect 3972 23933 4006 23967
rect 3972 23865 4006 23899
rect 3972 23797 4006 23831
rect 3972 23729 4006 23763
rect 3972 23661 4006 23695
rect 3972 23593 4006 23627
rect 3972 23525 4006 23559
rect 3972 23457 4006 23491
rect 3972 23389 4006 23423
rect 3972 23321 4006 23355
rect 3972 23253 4006 23287
rect 3972 23185 4006 23219
rect 3972 23117 4006 23151
rect 3972 23049 4006 23083
rect 3972 22981 4006 23015
rect 3972 22913 4006 22947
rect 3972 22845 4006 22879
rect 3972 22777 4006 22811
rect 3972 22709 4006 22743
rect 3972 22641 4006 22675
rect 3972 22573 4006 22607
rect 3972 22505 4006 22539
rect 3972 22437 4006 22471
rect 3972 22369 4006 22403
rect 3972 22301 4006 22335
rect 3972 22233 4006 22267
rect 3972 22165 4006 22199
rect 3972 22097 4006 22131
rect 3972 22029 4006 22063
rect 3972 21961 4006 21995
rect 3972 21893 4006 21927
rect 3972 21825 4006 21859
rect 3972 21757 4006 21791
rect 3972 21689 4006 21723
rect 3972 21621 4006 21655
rect 3972 21553 4006 21587
rect 3972 21485 4006 21519
rect 3972 21417 4006 21451
rect 3972 21349 4006 21383
rect 3972 21281 4006 21315
rect 3972 21213 4006 21247
rect 3972 21145 4006 21179
rect 3972 21077 4006 21111
rect 3972 21009 4006 21043
rect 3972 20941 4006 20975
rect 3972 20873 4006 20907
rect 3972 20805 4006 20839
rect 3972 20737 4006 20771
rect 3972 20669 4006 20703
rect 3972 20601 4006 20635
rect 3972 20533 4006 20567
rect 3972 20465 4006 20499
rect 3972 20397 4006 20431
rect 3972 20329 4006 20363
rect 3972 20261 4006 20295
rect 3972 20193 4006 20227
rect 3972 20125 4006 20159
rect 3972 20057 4006 20091
rect 3972 19989 4006 20023
rect 3972 19921 4006 19955
rect 3972 19853 4006 19887
rect 3972 19785 4006 19819
rect 3972 19717 4006 19751
rect 3972 19649 4006 19683
rect 3972 19581 4006 19615
rect 3972 19513 4006 19547
rect 3972 19445 4006 19479
rect 3972 19377 4006 19411
rect 3972 19309 4006 19343
rect 3972 19241 4006 19275
rect 3972 19173 4006 19207
rect 3972 19105 4006 19139
rect 3972 19037 4006 19071
rect 3972 18969 4006 19003
rect 3972 18901 4006 18935
rect 3972 18833 4006 18867
rect 3972 18765 4006 18799
rect 3972 18697 4006 18731
rect 3972 18629 4006 18663
rect 3972 18561 4006 18595
rect 3972 18493 4006 18527
rect 3972 18425 4006 18459
rect 3972 18357 4006 18391
rect 3972 18289 4006 18323
rect 3972 18221 4006 18255
rect 3972 18153 4006 18187
rect 3972 18085 4006 18119
rect 3972 18017 4006 18051
rect 3972 17949 4006 17983
rect 3972 17881 4006 17915
rect 3972 17813 4006 17847
rect 3972 17745 4006 17779
rect 3972 17677 4006 17711
rect 3972 17609 4006 17643
rect 3972 17541 4006 17575
rect 3972 17473 4006 17507
rect 3972 17405 4006 17439
rect 3972 17337 4006 17371
rect 3972 17269 4006 17303
rect 3972 17201 4006 17235
rect 3972 17133 4006 17167
rect 3972 17065 4006 17099
rect 3972 16997 4006 17031
rect 3972 16929 4006 16963
rect 3972 16861 4006 16895
rect 3972 16793 4006 16827
rect 3972 16725 4006 16759
rect 3972 16657 4006 16691
rect 3972 16589 4006 16623
rect 3972 16521 4006 16555
rect 3972 16453 4006 16487
rect 3972 16385 4006 16419
rect 3972 16317 4006 16351
rect 3972 16249 4006 16283
rect 3972 16181 4006 16215
rect 3972 16113 4006 16147
rect 3972 16045 4006 16079
rect 3972 15977 4006 16011
rect 3972 15909 4006 15943
rect 3972 15841 4006 15875
rect 3972 15773 4006 15807
rect 3972 15705 4006 15739
rect 3972 15637 4006 15671
rect 3972 15569 4006 15603
rect 3972 15501 4006 15535
rect 3972 15433 4006 15467
rect 3972 15365 4006 15399
rect 3972 15297 4006 15331
rect 3972 15229 4006 15263
rect 3972 15161 4006 15195
rect 3972 15093 4006 15127
rect 3972 15025 4006 15059
rect 3972 14957 4006 14991
rect 3972 14889 4006 14923
rect 3972 14821 4006 14855
rect 3972 14753 4006 14787
rect 3972 14685 4006 14719
rect 3972 14617 4006 14651
rect 3972 14549 4006 14583
rect 3972 14481 4006 14515
rect 3972 14413 4006 14447
rect 3972 14345 4006 14379
rect 3972 14277 4006 14311
rect 3972 14209 4006 14243
rect 3972 14141 4006 14175
rect 3972 14073 4006 14107
rect 3972 14005 4006 14039
rect 3972 13937 4006 13971
rect 3972 13869 4006 13903
rect 3972 13801 4006 13835
rect 3972 13733 4006 13767
rect 3972 13665 4006 13699
rect 3972 13597 4006 13631
rect 3972 13529 4006 13563
rect 3972 13461 4006 13495
rect 3972 13393 4006 13427
rect 3972 13325 4006 13359
rect 3972 13257 4006 13291
rect 3972 13189 4006 13223
rect 3972 13121 4006 13155
rect 3972 13053 4006 13087
rect 3972 12985 4006 13019
rect 3972 12917 4006 12951
rect 3972 12849 4006 12883
rect 3972 12781 4006 12815
rect 3972 12713 4006 12747
rect 3972 12645 4006 12679
rect 3972 12577 4006 12611
rect 3972 12509 4006 12543
rect 3972 12441 4006 12475
rect 3972 12373 4006 12407
rect 3972 12305 4006 12339
rect 3972 12237 4006 12271
rect 3972 12169 4006 12203
rect 3972 12101 4006 12135
rect 3972 12033 4006 12067
rect 3972 11965 4006 11999
rect 3972 11897 4006 11931
rect 3972 11829 4006 11863
rect 3972 11761 4006 11795
rect 3972 11693 4006 11727
rect 3972 11625 4006 11659
rect 3972 11557 4006 11591
rect 3972 11489 4006 11523
rect 3972 11421 4006 11455
rect 3972 11353 4006 11387
rect 3972 11285 4006 11319
rect 3972 11217 4006 11251
rect 3972 11149 4006 11183
rect 3972 11081 4006 11115
rect 3972 11013 4006 11047
rect 3972 10945 4006 10979
rect 3972 10877 4006 10911
rect 3972 10809 4006 10843
rect 3972 10741 4006 10775
rect 3972 10673 4006 10707
rect 3972 10605 4006 10639
rect 3972 10537 4006 10571
rect 3972 10469 4006 10503
rect 3972 10401 4006 10435
rect 3972 10333 4006 10367
rect 3972 10265 4006 10299
rect 3972 10197 4006 10231
rect 3972 10129 4006 10163
rect 3972 10061 4006 10095
rect 3972 9993 4006 10027
rect 3972 9925 4006 9959
rect 3972 9857 4006 9891
rect 3972 9789 4006 9823
rect 3972 9721 4006 9755
rect 3972 9653 4006 9687
rect 3972 9585 4006 9619
rect 3972 9517 4006 9551
rect 3972 9449 4006 9483
rect 3972 9381 4006 9415
rect 3972 9313 4006 9347
rect 3972 9245 4006 9279
rect 3972 9177 4006 9211
rect 3972 9109 4006 9143
rect 3972 9041 4006 9075
rect 3972 8973 4006 9007
rect 3972 8905 4006 8939
rect 3972 8837 4006 8871
rect 3972 8769 4006 8803
rect 3972 8701 4006 8735
rect 3972 8633 4006 8667
rect 3972 8565 4006 8599
rect 3972 8497 4006 8531
rect 3972 8429 4006 8463
rect 3972 8361 4006 8395
rect 3972 8293 4006 8327
rect 3972 8225 4006 8259
rect 3972 8157 4006 8191
rect 3972 8089 4006 8123
rect 3972 8021 4006 8055
rect 3972 7953 4006 7987
rect 3972 7885 4006 7919
rect 3972 7817 4006 7851
rect 3972 7749 4006 7783
rect 3972 7681 4006 7715
rect 3972 7613 4006 7647
rect 3972 7545 4006 7579
rect 3972 7477 4006 7511
rect 3972 7409 4006 7443
rect 3972 7341 4006 7375
rect 3972 7273 4006 7307
rect 3972 7205 4006 7239
rect 3972 7137 4006 7171
rect 3972 7069 4006 7103
rect 3972 7001 4006 7035
rect 3972 6933 4006 6967
rect 3972 6865 4006 6899
rect 3972 6797 4006 6831
rect 3972 6729 4006 6763
rect 3972 6661 4006 6695
rect 3972 6593 4006 6627
rect 3972 6525 4006 6559
rect 3972 6457 4006 6491
rect 3972 6389 4006 6423
rect 3972 6321 4006 6355
rect 3972 6253 4006 6287
rect 3972 6185 4006 6219
rect 3972 6117 4006 6151
rect 3972 6049 4006 6083
rect 3972 5981 4006 6015
rect 3972 5913 4006 5947
rect 3972 5845 4006 5879
rect 3972 5777 4006 5811
rect 3972 5709 4006 5743
rect 3972 5641 4006 5675
rect 3972 5573 4006 5607
rect 3972 5505 4006 5539
rect 3972 5437 4006 5471
rect 3972 5369 4006 5403
rect 3972 5301 4006 5335
rect 3972 5233 4006 5267
rect 3972 5165 4006 5199
rect 3972 5097 4006 5131
rect 3972 5029 4006 5063
rect 3972 4961 4006 4995
rect 3972 4893 4006 4927
rect 3972 4825 4006 4859
rect 3972 4757 4006 4791
rect 3972 4689 4006 4723
rect 3972 4621 4006 4655
rect 3972 4553 4006 4587
rect 3972 4485 4006 4519
rect 3972 4417 4006 4451
rect 3972 4349 4006 4383
rect 3972 4281 4006 4315
rect 3972 4213 4006 4247
rect 3972 4145 4006 4179
rect 3972 4077 4006 4111
rect 3972 4009 4006 4043
rect 3972 3941 4006 3975
rect 3972 3873 4006 3907
rect 3972 3805 4006 3839
rect 3972 3737 4006 3771
rect 3972 3669 4006 3703
rect 3972 3601 4006 3635
rect 3972 3533 4006 3567
rect 1830 3417 1864 3451
rect -252 3213 -218 3295
rect 1830 3349 1864 3383
rect 3972 3465 4006 3499
rect 6114 38641 6148 38723
rect 6114 38573 6148 38607
rect 6114 38505 6148 38539
rect 6114 38437 6148 38471
rect 6114 38369 6148 38403
rect 6114 38301 6148 38335
rect 6114 38233 6148 38267
rect 6114 38165 6148 38199
rect 6114 38097 6148 38131
rect 6114 38029 6148 38063
rect 6114 37961 6148 37995
rect 6114 37893 6148 37927
rect 6114 37825 6148 37859
rect 6114 37757 6148 37791
rect 6114 37689 6148 37723
rect 6114 37621 6148 37655
rect 6114 37553 6148 37587
rect 6114 37485 6148 37519
rect 6114 37417 6148 37451
rect 6114 37349 6148 37383
rect 6114 37281 6148 37315
rect 6114 37213 6148 37247
rect 6114 37145 6148 37179
rect 6114 37077 6148 37111
rect 6114 37009 6148 37043
rect 6114 36941 6148 36975
rect 6114 36873 6148 36907
rect 6114 36805 6148 36839
rect 6114 36737 6148 36771
rect 6114 36669 6148 36703
rect 6114 36601 6148 36635
rect 6114 36533 6148 36567
rect 6114 36465 6148 36499
rect 6114 36397 6148 36431
rect 6114 36329 6148 36363
rect 6114 36261 6148 36295
rect 6114 36193 6148 36227
rect 6114 36125 6148 36159
rect 6114 36057 6148 36091
rect 6114 35989 6148 36023
rect 6114 35921 6148 35955
rect 6114 35853 6148 35887
rect 6114 35785 6148 35819
rect 6114 35717 6148 35751
rect 6114 35649 6148 35683
rect 6114 35581 6148 35615
rect 6114 35513 6148 35547
rect 6114 35445 6148 35479
rect 6114 35377 6148 35411
rect 6114 35309 6148 35343
rect 6114 35241 6148 35275
rect 6114 35173 6148 35207
rect 6114 35105 6148 35139
rect 6114 35037 6148 35071
rect 6114 34969 6148 35003
rect 6114 34901 6148 34935
rect 6114 34833 6148 34867
rect 6114 34765 6148 34799
rect 6114 34697 6148 34731
rect 6114 34629 6148 34663
rect 6114 34561 6148 34595
rect 6114 34493 6148 34527
rect 6114 34425 6148 34459
rect 6114 34357 6148 34391
rect 6114 34289 6148 34323
rect 6114 34221 6148 34255
rect 6114 34153 6148 34187
rect 6114 34085 6148 34119
rect 6114 34017 6148 34051
rect 6114 33949 6148 33983
rect 6114 33881 6148 33915
rect 6114 33813 6148 33847
rect 6114 33745 6148 33779
rect 6114 33677 6148 33711
rect 6114 33609 6148 33643
rect 6114 33541 6148 33575
rect 6114 33473 6148 33507
rect 6114 33405 6148 33439
rect 6114 33337 6148 33371
rect 6114 33269 6148 33303
rect 6114 33201 6148 33235
rect 6114 33133 6148 33167
rect 6114 33065 6148 33099
rect 6114 32997 6148 33031
rect 6114 32929 6148 32963
rect 6114 32861 6148 32895
rect 6114 32793 6148 32827
rect 6114 32725 6148 32759
rect 6114 32657 6148 32691
rect 6114 32589 6148 32623
rect 6114 32521 6148 32555
rect 6114 32453 6148 32487
rect 6114 32385 6148 32419
rect 6114 32317 6148 32351
rect 6114 32249 6148 32283
rect 6114 32181 6148 32215
rect 6114 32113 6148 32147
rect 6114 32045 6148 32079
rect 6114 31977 6148 32011
rect 6114 31909 6148 31943
rect 6114 31841 6148 31875
rect 6114 31773 6148 31807
rect 6114 31705 6148 31739
rect 6114 31637 6148 31671
rect 6114 31569 6148 31603
rect 6114 31501 6148 31535
rect 6114 31433 6148 31467
rect 6114 31365 6148 31399
rect 6114 31297 6148 31331
rect 6114 31229 6148 31263
rect 6114 31161 6148 31195
rect 6114 31093 6148 31127
rect 6114 31025 6148 31059
rect 6114 30957 6148 30991
rect 6114 30889 6148 30923
rect 6114 30821 6148 30855
rect 6114 30753 6148 30787
rect 6114 30685 6148 30719
rect 6114 30617 6148 30651
rect 6114 30549 6148 30583
rect 6114 30481 6148 30515
rect 6114 30413 6148 30447
rect 6114 30345 6148 30379
rect 6114 30277 6148 30311
rect 6114 30209 6148 30243
rect 6114 30141 6148 30175
rect 6114 30073 6148 30107
rect 6114 30005 6148 30039
rect 6114 29937 6148 29971
rect 6114 29869 6148 29903
rect 6114 29801 6148 29835
rect 6114 29733 6148 29767
rect 6114 29665 6148 29699
rect 6114 29597 6148 29631
rect 6114 29529 6148 29563
rect 6114 29461 6148 29495
rect 6114 29393 6148 29427
rect 6114 29325 6148 29359
rect 6114 29257 6148 29291
rect 6114 29189 6148 29223
rect 6114 29121 6148 29155
rect 6114 29053 6148 29087
rect 6114 28985 6148 29019
rect 6114 28917 6148 28951
rect 6114 28849 6148 28883
rect 6114 28781 6148 28815
rect 6114 28713 6148 28747
rect 6114 28645 6148 28679
rect 6114 28577 6148 28611
rect 6114 28509 6148 28543
rect 6114 28441 6148 28475
rect 6114 28373 6148 28407
rect 6114 28305 6148 28339
rect 6114 28237 6148 28271
rect 6114 28169 6148 28203
rect 6114 28101 6148 28135
rect 6114 28033 6148 28067
rect 6114 27965 6148 27999
rect 6114 27897 6148 27931
rect 6114 27829 6148 27863
rect 6114 27761 6148 27795
rect 6114 27693 6148 27727
rect 6114 27625 6148 27659
rect 6114 27557 6148 27591
rect 6114 27489 6148 27523
rect 6114 27421 6148 27455
rect 6114 27353 6148 27387
rect 6114 27285 6148 27319
rect 6114 27217 6148 27251
rect 6114 27149 6148 27183
rect 6114 27081 6148 27115
rect 6114 27013 6148 27047
rect 6114 26945 6148 26979
rect 6114 26877 6148 26911
rect 6114 26809 6148 26843
rect 6114 26741 6148 26775
rect 6114 26673 6148 26707
rect 6114 26605 6148 26639
rect 6114 26537 6148 26571
rect 6114 26469 6148 26503
rect 6114 26401 6148 26435
rect 6114 26333 6148 26367
rect 6114 26265 6148 26299
rect 6114 26197 6148 26231
rect 6114 26129 6148 26163
rect 6114 26061 6148 26095
rect 6114 25993 6148 26027
rect 6114 25925 6148 25959
rect 6114 25857 6148 25891
rect 6114 25789 6148 25823
rect 6114 25721 6148 25755
rect 6114 25653 6148 25687
rect 6114 25585 6148 25619
rect 6114 25517 6148 25551
rect 6114 25449 6148 25483
rect 6114 25381 6148 25415
rect 6114 25313 6148 25347
rect 6114 25245 6148 25279
rect 6114 25177 6148 25211
rect 6114 25109 6148 25143
rect 6114 25041 6148 25075
rect 6114 24973 6148 25007
rect 6114 24905 6148 24939
rect 6114 24837 6148 24871
rect 6114 24769 6148 24803
rect 6114 24701 6148 24735
rect 6114 24633 6148 24667
rect 6114 24565 6148 24599
rect 6114 24497 6148 24531
rect 6114 24429 6148 24463
rect 6114 24361 6148 24395
rect 6114 24293 6148 24327
rect 6114 24225 6148 24259
rect 6114 24157 6148 24191
rect 6114 24089 6148 24123
rect 6114 24021 6148 24055
rect 6114 23953 6148 23987
rect 6114 23885 6148 23919
rect 6114 23817 6148 23851
rect 6114 23749 6148 23783
rect 6114 23681 6148 23715
rect 6114 23613 6148 23647
rect 6114 23545 6148 23579
rect 6114 23477 6148 23511
rect 6114 23409 6148 23443
rect 6114 23341 6148 23375
rect 6114 23273 6148 23307
rect 6114 23205 6148 23239
rect 6114 23137 6148 23171
rect 6114 23069 6148 23103
rect 6114 23001 6148 23035
rect 6114 22933 6148 22967
rect 6114 22865 6148 22899
rect 6114 22797 6148 22831
rect 6114 22729 6148 22763
rect 6114 22661 6148 22695
rect 6114 22593 6148 22627
rect 6114 22525 6148 22559
rect 6114 22457 6148 22491
rect 6114 22389 6148 22423
rect 6114 22321 6148 22355
rect 6114 22253 6148 22287
rect 6114 22185 6148 22219
rect 6114 22117 6148 22151
rect 6114 22049 6148 22083
rect 6114 21981 6148 22015
rect 6114 21913 6148 21947
rect 6114 21845 6148 21879
rect 6114 21777 6148 21811
rect 6114 21709 6148 21743
rect 6114 21641 6148 21675
rect 6114 21573 6148 21607
rect 6114 21505 6148 21539
rect 6114 21437 6148 21471
rect 6114 21369 6148 21403
rect 6114 21301 6148 21335
rect 6114 21233 6148 21267
rect 6114 21165 6148 21199
rect 6114 21097 6148 21131
rect 6114 21029 6148 21063
rect 6114 20961 6148 20995
rect 6114 20893 6148 20927
rect 6114 20825 6148 20859
rect 6114 20757 6148 20791
rect 6114 20689 6148 20723
rect 6114 20621 6148 20655
rect 6114 20553 6148 20587
rect 6114 20485 6148 20519
rect 6114 20417 6148 20451
rect 6114 20349 6148 20383
rect 6114 20281 6148 20315
rect 6114 20213 6148 20247
rect 6114 20145 6148 20179
rect 6114 20077 6148 20111
rect 6114 20009 6148 20043
rect 6114 19941 6148 19975
rect 6114 19873 6148 19907
rect 6114 19805 6148 19839
rect 6114 19737 6148 19771
rect 6114 19669 6148 19703
rect 6114 19601 6148 19635
rect 6114 19533 6148 19567
rect 6114 19465 6148 19499
rect 6114 19397 6148 19431
rect 6114 19329 6148 19363
rect 6114 19261 6148 19295
rect 6114 19193 6148 19227
rect 6114 19125 6148 19159
rect 6114 19057 6148 19091
rect 6114 18989 6148 19023
rect 6114 18921 6148 18955
rect 6114 18853 6148 18887
rect 6114 18785 6148 18819
rect 6114 18717 6148 18751
rect 6114 18649 6148 18683
rect 6114 18581 6148 18615
rect 6114 18513 6148 18547
rect 6114 18445 6148 18479
rect 6114 18377 6148 18411
rect 6114 18309 6148 18343
rect 6114 18241 6148 18275
rect 6114 18173 6148 18207
rect 6114 18105 6148 18139
rect 6114 18037 6148 18071
rect 6114 17969 6148 18003
rect 6114 17901 6148 17935
rect 6114 17833 6148 17867
rect 6114 17765 6148 17799
rect 6114 17697 6148 17731
rect 6114 17629 6148 17663
rect 6114 17561 6148 17595
rect 6114 17493 6148 17527
rect 6114 17425 6148 17459
rect 6114 17357 6148 17391
rect 6114 17289 6148 17323
rect 6114 17221 6148 17255
rect 6114 17153 6148 17187
rect 6114 17085 6148 17119
rect 6114 17017 6148 17051
rect 6114 16949 6148 16983
rect 6114 16881 6148 16915
rect 6114 16813 6148 16847
rect 6114 16745 6148 16779
rect 6114 16677 6148 16711
rect 6114 16609 6148 16643
rect 6114 16541 6148 16575
rect 6114 16473 6148 16507
rect 6114 16405 6148 16439
rect 6114 16337 6148 16371
rect 6114 16269 6148 16303
rect 6114 16201 6148 16235
rect 6114 16133 6148 16167
rect 6114 16065 6148 16099
rect 6114 15997 6148 16031
rect 6114 15929 6148 15963
rect 6114 15861 6148 15895
rect 6114 15793 6148 15827
rect 6114 15725 6148 15759
rect 6114 15657 6148 15691
rect 6114 15589 6148 15623
rect 6114 15521 6148 15555
rect 6114 15453 6148 15487
rect 6114 15385 6148 15419
rect 6114 15317 6148 15351
rect 6114 15249 6148 15283
rect 6114 15181 6148 15215
rect 6114 15113 6148 15147
rect 6114 15045 6148 15079
rect 6114 14977 6148 15011
rect 6114 14909 6148 14943
rect 6114 14841 6148 14875
rect 6114 14773 6148 14807
rect 6114 14705 6148 14739
rect 6114 14637 6148 14671
rect 6114 14569 6148 14603
rect 6114 14501 6148 14535
rect 6114 14433 6148 14467
rect 6114 14365 6148 14399
rect 6114 14297 6148 14331
rect 6114 14229 6148 14263
rect 6114 14161 6148 14195
rect 6114 14093 6148 14127
rect 6114 14025 6148 14059
rect 6114 13957 6148 13991
rect 6114 13889 6148 13923
rect 6114 13821 6148 13855
rect 6114 13753 6148 13787
rect 6114 13685 6148 13719
rect 6114 13617 6148 13651
rect 6114 13549 6148 13583
rect 6114 13481 6148 13515
rect 6114 13413 6148 13447
rect 6114 13345 6148 13379
rect 6114 13277 6148 13311
rect 6114 13209 6148 13243
rect 6114 13141 6148 13175
rect 6114 13073 6148 13107
rect 6114 13005 6148 13039
rect 6114 12937 6148 12971
rect 6114 12869 6148 12903
rect 6114 12801 6148 12835
rect 6114 12733 6148 12767
rect 6114 12665 6148 12699
rect 6114 12597 6148 12631
rect 6114 12529 6148 12563
rect 6114 12461 6148 12495
rect 6114 12393 6148 12427
rect 6114 12325 6148 12359
rect 6114 12257 6148 12291
rect 6114 12189 6148 12223
rect 6114 12121 6148 12155
rect 6114 12053 6148 12087
rect 6114 11985 6148 12019
rect 6114 11917 6148 11951
rect 6114 11849 6148 11883
rect 6114 11781 6148 11815
rect 6114 11713 6148 11747
rect 6114 11645 6148 11679
rect 6114 11577 6148 11611
rect 6114 11509 6148 11543
rect 6114 11441 6148 11475
rect 6114 11373 6148 11407
rect 6114 11305 6148 11339
rect 6114 11237 6148 11271
rect 6114 11169 6148 11203
rect 6114 11101 6148 11135
rect 6114 11033 6148 11067
rect 6114 10965 6148 10999
rect 6114 10897 6148 10931
rect 6114 10829 6148 10863
rect 6114 10761 6148 10795
rect 6114 10693 6148 10727
rect 6114 10625 6148 10659
rect 6114 10557 6148 10591
rect 6114 10489 6148 10523
rect 6114 10421 6148 10455
rect 6114 10353 6148 10387
rect 6114 10285 6148 10319
rect 6114 10217 6148 10251
rect 6114 10149 6148 10183
rect 6114 10081 6148 10115
rect 6114 10013 6148 10047
rect 6114 9945 6148 9979
rect 6114 9877 6148 9911
rect 6114 9809 6148 9843
rect 6114 9741 6148 9775
rect 6114 9673 6148 9707
rect 6114 9605 6148 9639
rect 6114 9537 6148 9571
rect 6114 9469 6148 9503
rect 6114 9401 6148 9435
rect 6114 9333 6148 9367
rect 6114 9265 6148 9299
rect 6114 9197 6148 9231
rect 6114 9129 6148 9163
rect 6114 9061 6148 9095
rect 6114 8993 6148 9027
rect 6114 8925 6148 8959
rect 6114 8857 6148 8891
rect 6114 8789 6148 8823
rect 6114 8721 6148 8755
rect 6114 8653 6148 8687
rect 6114 8585 6148 8619
rect 6114 8517 6148 8551
rect 6114 8449 6148 8483
rect 6114 8381 6148 8415
rect 6114 8313 6148 8347
rect 6114 8245 6148 8279
rect 6114 8177 6148 8211
rect 6114 8109 6148 8143
rect 6114 8041 6148 8075
rect 6114 7973 6148 8007
rect 6114 7905 6148 7939
rect 6114 7837 6148 7871
rect 6114 7769 6148 7803
rect 6114 7701 6148 7735
rect 6114 7633 6148 7667
rect 6114 7565 6148 7599
rect 6114 7497 6148 7531
rect 6114 7429 6148 7463
rect 6114 7361 6148 7395
rect 6114 7293 6148 7327
rect 6114 7225 6148 7259
rect 6114 7157 6148 7191
rect 6114 7089 6148 7123
rect 6114 7021 6148 7055
rect 6114 6953 6148 6987
rect 6114 6885 6148 6919
rect 6114 6817 6148 6851
rect 6114 6749 6148 6783
rect 6114 6681 6148 6715
rect 6114 6613 6148 6647
rect 6114 6545 6148 6579
rect 6114 6477 6148 6511
rect 6114 6409 6148 6443
rect 6114 6341 6148 6375
rect 6114 6273 6148 6307
rect 6114 6205 6148 6239
rect 6114 6137 6148 6171
rect 6114 6069 6148 6103
rect 6114 6001 6148 6035
rect 6114 5933 6148 5967
rect 6114 5865 6148 5899
rect 6114 5797 6148 5831
rect 6114 5729 6148 5763
rect 6114 5661 6148 5695
rect 6114 5593 6148 5627
rect 6114 5525 6148 5559
rect 6114 5457 6148 5491
rect 6114 5389 6148 5423
rect 6114 5321 6148 5355
rect 6114 5253 6148 5287
rect 6114 5185 6148 5219
rect 6114 5117 6148 5151
rect 6114 5049 6148 5083
rect 6114 4981 6148 5015
rect 6114 4913 6148 4947
rect 6114 4845 6148 4879
rect 6114 4777 6148 4811
rect 6114 4709 6148 4743
rect 6114 4641 6148 4675
rect 6114 4573 6148 4607
rect 6114 4505 6148 4539
rect 6114 4437 6148 4471
rect 6114 4369 6148 4403
rect 6114 4301 6148 4335
rect 6114 4233 6148 4267
rect 6114 4165 6148 4199
rect 6114 4097 6148 4131
rect 6114 4029 6148 4063
rect 6114 3961 6148 3995
rect 6114 3893 6148 3927
rect 6114 3825 6148 3859
rect 6114 3757 6148 3791
rect 6114 3689 6148 3723
rect 6114 3621 6148 3655
rect 6114 3553 6148 3587
rect 6114 3485 6148 3519
rect 3972 3397 4006 3431
rect 1830 3281 1864 3315
rect 1830 3213 1864 3247
rect 3972 3329 4006 3363
rect 6114 3417 6148 3451
rect 3972 3213 4006 3295
rect 6114 3349 6148 3383
rect 6114 3281 6148 3315
rect 6114 3213 6148 3247
rect -252 3179 -184 3213
rect -150 3179 -116 3213
rect -82 3179 -48 3213
rect -14 3179 20 3213
rect 54 3179 88 3213
rect 122 3179 156 3213
rect 190 3179 224 3213
rect 258 3179 292 3213
rect 326 3179 360 3213
rect 394 3179 428 3213
rect 462 3179 496 3213
rect 530 3179 564 3213
rect 598 3179 632 3213
rect 666 3179 700 3213
rect 734 3179 768 3213
rect 802 3179 836 3213
rect 870 3179 904 3213
rect 938 3179 972 3213
rect 1006 3179 1040 3213
rect 1074 3179 1108 3213
rect 1142 3179 1176 3213
rect 1210 3179 1244 3213
rect 1278 3179 1312 3213
rect 1346 3179 1380 3213
rect 1414 3179 1448 3213
rect 1482 3179 1516 3213
rect 1550 3179 1584 3213
rect 1618 3179 1652 3213
rect 1686 3179 1720 3213
rect 1754 3179 1932 3213
rect 1966 3179 2000 3213
rect 2034 3179 2068 3213
rect 2102 3179 2136 3213
rect 2170 3179 2204 3213
rect 2238 3179 2272 3213
rect 2306 3179 2340 3213
rect 2374 3179 2408 3213
rect 2442 3179 2476 3213
rect 2510 3179 2544 3213
rect 2578 3179 2612 3213
rect 2646 3179 2680 3213
rect 2714 3179 2748 3213
rect 2782 3179 2816 3213
rect 2850 3179 2884 3213
rect 2918 3179 2952 3213
rect 2986 3179 3020 3213
rect 3054 3179 3088 3213
rect 3122 3179 3156 3213
rect 3190 3179 3224 3213
rect 3258 3179 3292 3213
rect 3326 3179 3360 3213
rect 3394 3179 3428 3213
rect 3462 3179 3496 3213
rect 3530 3179 3564 3213
rect 3598 3179 3632 3213
rect 3666 3179 3700 3213
rect 3734 3179 3768 3213
rect 3802 3179 3836 3213
rect 3870 3179 3904 3213
rect 3938 3179 4040 3213
rect 4074 3179 4108 3213
rect 4142 3179 4176 3213
rect 4210 3179 4244 3213
rect 4278 3179 4312 3213
rect 4346 3179 4380 3213
rect 4414 3179 4448 3213
rect 4482 3179 4516 3213
rect 4550 3179 4584 3213
rect 4618 3179 4652 3213
rect 4686 3179 4720 3213
rect 4754 3179 4788 3213
rect 4822 3179 4856 3213
rect 4890 3179 4924 3213
rect 4958 3179 4992 3213
rect 5026 3179 5060 3213
rect 5094 3179 5128 3213
rect 5162 3179 5196 3213
rect 5230 3179 5264 3213
rect 5298 3179 5332 3213
rect 5366 3179 5400 3213
rect 5434 3179 5468 3213
rect 5502 3179 5536 3213
rect 5570 3179 5604 3213
rect 5638 3179 5672 3213
rect 5706 3179 5740 3213
rect 5774 3179 5808 3213
rect 5842 3179 5876 3213
rect 5910 3179 5944 3213
rect 5978 3179 6012 3213
rect 6046 3179 6148 3213
rect 9088 38723 9206 38757
rect 9240 38723 9274 38757
rect 9308 38723 9342 38757
rect 9376 38723 9410 38757
rect 9444 38723 9478 38757
rect 9512 38723 9546 38757
rect 9580 38723 9614 38757
rect 9648 38723 9682 38757
rect 9716 38723 9750 38757
rect 9784 38723 9818 38757
rect 9852 38723 9886 38757
rect 9920 38723 9954 38757
rect 9988 38723 10022 38757
rect 10056 38723 10090 38757
rect 10124 38723 10158 38757
rect 10192 38723 10294 38757
rect 10328 38723 10362 38757
rect 10396 38723 10430 38757
rect 10464 38723 10498 38757
rect 10532 38723 10566 38757
rect 10600 38723 10634 38757
rect 10668 38723 10702 38757
rect 10736 38723 10770 38757
rect 10804 38723 10838 38757
rect 10872 38723 10906 38757
rect 10940 38723 10974 38757
rect 11008 38723 11042 38757
rect 11076 38723 11110 38757
rect 11144 38723 11178 38757
rect 11212 38723 11246 38757
rect 11280 38723 11314 38757
rect 11348 38723 11512 38757
rect 11546 38723 11580 38757
rect 11614 38723 11648 38757
rect 11682 38723 11716 38757
rect 11750 38723 11784 38757
rect 11818 38723 11852 38757
rect 11886 38723 11920 38757
rect 11954 38723 11988 38757
rect 12022 38723 12056 38757
rect 12090 38723 12124 38757
rect 12158 38723 12192 38757
rect 12226 38723 12260 38757
rect 12294 38723 12328 38757
rect 12362 38723 12396 38757
rect 12430 38723 12464 38757
rect 12498 38723 12532 38757
rect 12566 38723 12600 38757
rect 12634 38723 12668 38757
rect 12702 38723 12736 38757
rect 12770 38723 12804 38757
rect 12838 38723 12872 38757
rect 12906 38723 12940 38757
rect 12974 38723 13008 38757
rect 13042 38723 13076 38757
rect 13110 38723 13144 38757
rect 13178 38723 13280 38757
rect 13314 38723 13348 38757
rect 13382 38723 13416 38757
rect 13450 38723 13484 38757
rect 13518 38723 13552 38757
rect 13586 38723 13620 38757
rect 13654 38723 13688 38757
rect 13722 38723 13756 38757
rect 13790 38723 13824 38757
rect 13858 38723 13892 38757
rect 13926 38723 13960 38757
rect 13994 38723 14028 38757
rect 14062 38723 14096 38757
rect 14130 38723 14164 38757
rect 14198 38723 14232 38757
rect 14266 38723 14300 38757
rect 14334 38723 14368 38757
rect 14402 38723 14436 38757
rect 14470 38723 14504 38757
rect 14538 38723 14572 38757
rect 14606 38723 14640 38757
rect 14674 38723 14708 38757
rect 14742 38723 14776 38757
rect 14810 38723 14844 38757
rect 14878 38723 14974 38757
rect 9088 38689 9122 38723
rect 9088 38621 9122 38655
rect 9088 38553 9122 38587
rect 9088 38485 9122 38519
rect 9088 38417 9122 38451
rect 9088 38349 9122 38383
rect 9088 38281 9122 38315
rect 9088 38213 9122 38247
rect 9088 38145 9122 38179
rect 9088 38077 9122 38111
rect 9088 38009 9122 38043
rect 9088 37941 9122 37975
rect 9088 37873 9122 37907
rect 9088 37805 9122 37839
rect 9088 37737 9122 37771
rect 9088 37669 9122 37703
rect 9088 37601 9122 37635
rect 9088 37533 9122 37567
rect 9088 37465 9122 37499
rect 9088 37397 9122 37431
rect 9088 37329 9122 37363
rect 9088 37261 9122 37295
rect 9088 37193 9122 37227
rect 9088 37125 9122 37159
rect 9088 37057 9122 37091
rect 9088 36989 9122 37023
rect 9088 36921 9122 36955
rect 9088 36853 9122 36887
rect 9088 36785 9122 36819
rect 9088 36717 9122 36751
rect 9088 36649 9122 36683
rect 9088 36581 9122 36615
rect 9088 36513 9122 36547
rect 9088 36445 9122 36479
rect 9088 36377 9122 36411
rect 9088 36309 9122 36343
rect 9088 36241 9122 36275
rect 9088 36173 9122 36207
rect 9088 36105 9122 36139
rect 9088 36037 9122 36071
rect 9088 35969 9122 36003
rect 9088 35901 9122 35935
rect 9088 35833 9122 35867
rect 9088 35765 9122 35799
rect 9088 35697 9122 35731
rect 9088 35629 9122 35663
rect 9088 35561 9122 35595
rect 9088 35493 9122 35527
rect 9088 35425 9122 35459
rect 9088 35357 9122 35391
rect 9088 35289 9122 35323
rect 9088 35221 9122 35255
rect 9088 35153 9122 35187
rect 9088 35085 9122 35119
rect 9088 35017 9122 35051
rect 9088 34949 9122 34983
rect 9088 34881 9122 34915
rect 9088 34813 9122 34847
rect 9088 34745 9122 34779
rect 9088 34677 9122 34711
rect 9088 34609 9122 34643
rect 9088 34541 9122 34575
rect 9088 34473 9122 34507
rect 9088 34405 9122 34439
rect 9088 34337 9122 34371
rect 9088 34269 9122 34303
rect 9088 34201 9122 34235
rect 9088 34133 9122 34167
rect 9088 34065 9122 34099
rect 9088 33997 9122 34031
rect 9088 33929 9122 33963
rect 9088 33861 9122 33895
rect 9088 33793 9122 33827
rect 9088 33725 9122 33759
rect 9088 33657 9122 33691
rect 9088 33589 9122 33623
rect 9088 33521 9122 33555
rect 9088 33453 9122 33487
rect 9088 33385 9122 33419
rect 9088 33317 9122 33351
rect 9088 33249 9122 33283
rect 9088 33181 9122 33215
rect 9088 33113 9122 33147
rect 9088 33045 9122 33079
rect 9088 32977 9122 33011
rect 9088 32909 9122 32943
rect 9088 32841 9122 32875
rect 9088 32773 9122 32807
rect 9088 32705 9122 32739
rect 9088 32637 9122 32671
rect 9088 32569 9122 32603
rect 9088 32501 9122 32535
rect 9088 32433 9122 32467
rect 9088 32365 9122 32399
rect 9088 32297 9122 32331
rect 9088 32229 9122 32263
rect 9088 32161 9122 32195
rect 9088 32093 9122 32127
rect 9088 32025 9122 32059
rect 9088 31957 9122 31991
rect 9088 31889 9122 31923
rect 9088 31821 9122 31855
rect 9088 31753 9122 31787
rect 9088 31685 9122 31719
rect 9088 31617 9122 31651
rect 9088 31549 9122 31583
rect 9088 31481 9122 31515
rect 9088 31413 9122 31447
rect 9088 31345 9122 31379
rect 9088 31277 9122 31311
rect 9088 31209 9122 31243
rect 9088 31141 9122 31175
rect 9088 31073 9122 31107
rect 9088 31005 9122 31039
rect 9088 30937 9122 30971
rect 9088 30869 9122 30903
rect 9088 30801 9122 30835
rect 9088 30733 9122 30767
rect 9088 30665 9122 30699
rect 9088 30597 9122 30631
rect 9088 30529 9122 30563
rect 9088 30461 9122 30495
rect 9088 30393 9122 30427
rect 9088 30325 9122 30359
rect 9088 30257 9122 30291
rect 9088 30189 9122 30223
rect 9088 30121 9122 30155
rect 9088 30053 9122 30087
rect 9088 29985 9122 30019
rect 9088 29917 9122 29951
rect 9088 29849 9122 29883
rect 9088 29781 9122 29815
rect 9088 29713 9122 29747
rect 9088 29645 9122 29679
rect 9088 29577 9122 29611
rect 9088 29509 9122 29543
rect 9088 29441 9122 29475
rect 9088 29373 9122 29407
rect 9088 29305 9122 29339
rect 9088 29237 9122 29271
rect 9088 29169 9122 29203
rect 9088 29101 9122 29135
rect 9088 29033 9122 29067
rect 9088 28965 9122 28999
rect 9088 28897 9122 28931
rect 9088 28829 9122 28863
rect 9088 28761 9122 28795
rect 9088 28693 9122 28727
rect 9088 28625 9122 28659
rect 9088 28557 9122 28591
rect 9088 28489 9122 28523
rect 9088 28421 9122 28455
rect 9088 28353 9122 28387
rect 9088 28285 9122 28319
rect 9088 28217 9122 28251
rect 9088 28149 9122 28183
rect 9088 28081 9122 28115
rect 9088 28013 9122 28047
rect 9088 27945 9122 27979
rect 9088 27877 9122 27911
rect 9088 27809 9122 27843
rect 9088 27741 9122 27775
rect 9088 27673 9122 27707
rect 9088 27605 9122 27639
rect 9088 27537 9122 27571
rect 9088 27469 9122 27503
rect 9088 27401 9122 27435
rect 9088 27333 9122 27367
rect 9088 27265 9122 27299
rect 9088 27197 9122 27231
rect 9088 27129 9122 27163
rect 9088 27061 9122 27095
rect 9088 26993 9122 27027
rect 9088 26925 9122 26959
rect 9088 26857 9122 26891
rect 9088 26789 9122 26823
rect 9088 26721 9122 26755
rect 9088 26653 9122 26687
rect 9088 26585 9122 26619
rect 9088 26517 9122 26551
rect 9088 26449 9122 26483
rect 9088 26381 9122 26415
rect 9088 26313 9122 26347
rect 9088 26245 9122 26279
rect 9088 26177 9122 26211
rect 9088 26109 9122 26143
rect 9088 26041 9122 26075
rect 9088 25973 9122 26007
rect 9088 25905 9122 25939
rect 9088 25837 9122 25871
rect 9088 25769 9122 25803
rect 9088 25701 9122 25735
rect 9088 25633 9122 25667
rect 9088 25565 9122 25599
rect 9088 25497 9122 25531
rect 9088 25429 9122 25463
rect 9088 25361 9122 25395
rect 9088 25293 9122 25327
rect 9088 25225 9122 25259
rect 9088 25157 9122 25191
rect 9088 25089 9122 25123
rect 9088 25021 9122 25055
rect 9088 24953 9122 24987
rect 9088 24885 9122 24919
rect 9088 24817 9122 24851
rect 9088 24749 9122 24783
rect 9088 24681 9122 24715
rect 9088 24613 9122 24647
rect 9088 24545 9122 24579
rect 9088 24477 9122 24511
rect 9088 24409 9122 24443
rect 9088 24341 9122 24375
rect 9088 24273 9122 24307
rect 9088 24205 9122 24239
rect 9088 24137 9122 24171
rect 9088 24069 9122 24103
rect 9088 24001 9122 24035
rect 9088 23933 9122 23967
rect 9088 23865 9122 23899
rect 9088 23797 9122 23831
rect 9088 23729 9122 23763
rect 9088 23661 9122 23695
rect 9088 23593 9122 23627
rect 9088 23525 9122 23559
rect 9088 23457 9122 23491
rect 9088 23389 9122 23423
rect 9088 23321 9122 23355
rect 9088 23253 9122 23287
rect 9088 23185 9122 23219
rect 9088 23117 9122 23151
rect 9088 23049 9122 23083
rect 9088 22981 9122 23015
rect 9088 22913 9122 22947
rect 9088 22845 9122 22879
rect 9088 22777 9122 22811
rect 9088 22709 9122 22743
rect 9088 22641 9122 22675
rect 9088 22573 9122 22607
rect 9088 22505 9122 22539
rect 9088 22437 9122 22471
rect 9088 22369 9122 22403
rect 9088 22301 9122 22335
rect 9088 22233 9122 22267
rect 9088 22165 9122 22199
rect 9088 22097 9122 22131
rect 9088 22029 9122 22063
rect 9088 21961 9122 21995
rect 9088 21893 9122 21927
rect 9088 21825 9122 21859
rect 9088 21757 9122 21791
rect 9088 21689 9122 21723
rect 9088 21621 9122 21655
rect 9088 21553 9122 21587
rect 9088 21485 9122 21519
rect 9088 21417 9122 21451
rect 9088 21349 9122 21383
rect 9088 21281 9122 21315
rect 9088 21213 9122 21247
rect 9088 21145 9122 21179
rect 9088 21077 9122 21111
rect 9088 21009 9122 21043
rect 9088 20941 9122 20975
rect 9088 20873 9122 20907
rect 9088 20805 9122 20839
rect 9088 20737 9122 20771
rect 9088 20669 9122 20703
rect 9088 20601 9122 20635
rect 9088 20533 9122 20567
rect 9088 20465 9122 20499
rect 9088 20397 9122 20431
rect 9088 20329 9122 20363
rect 9088 20261 9122 20295
rect 9088 20193 9122 20227
rect 9088 20125 9122 20159
rect 9088 20057 9122 20091
rect 9088 19989 9122 20023
rect 9088 19921 9122 19955
rect 9088 19853 9122 19887
rect 9088 19785 9122 19819
rect 9088 19717 9122 19751
rect 9088 19649 9122 19683
rect 9088 19581 9122 19615
rect 9088 19513 9122 19547
rect 9088 19445 9122 19479
rect 9088 19377 9122 19411
rect 9088 19309 9122 19343
rect 9088 19241 9122 19275
rect 9088 19173 9122 19207
rect 9088 19105 9122 19139
rect 9088 19037 9122 19071
rect 9088 18969 9122 19003
rect 9088 18901 9122 18935
rect 9088 18833 9122 18867
rect 9088 18765 9122 18799
rect 9088 18697 9122 18731
rect 9088 18629 9122 18663
rect 9088 18561 9122 18595
rect 9088 18493 9122 18527
rect 9088 18425 9122 18459
rect 9088 18357 9122 18391
rect 9088 18289 9122 18323
rect 9088 18221 9122 18255
rect 9088 18153 9122 18187
rect 9088 18085 9122 18119
rect 9088 18017 9122 18051
rect 9088 17949 9122 17983
rect 9088 17881 9122 17915
rect 9088 17813 9122 17847
rect 9088 17745 9122 17779
rect 9088 17677 9122 17711
rect 9088 17609 9122 17643
rect 9088 17541 9122 17575
rect 9088 17473 9122 17507
rect 9088 17405 9122 17439
rect 9088 17337 9122 17371
rect 9088 17269 9122 17303
rect 9088 17201 9122 17235
rect 9088 17133 9122 17167
rect 9088 17065 9122 17099
rect 9088 16997 9122 17031
rect 9088 16929 9122 16963
rect 9088 16861 9122 16895
rect 9088 16793 9122 16827
rect 9088 16725 9122 16759
rect 9088 16657 9122 16691
rect 9088 16589 9122 16623
rect 9088 16521 9122 16555
rect 9088 16453 9122 16487
rect 9088 16385 9122 16419
rect 9088 16317 9122 16351
rect 9088 16249 9122 16283
rect 9088 16181 9122 16215
rect 9088 16113 9122 16147
rect 9088 16045 9122 16079
rect 9088 15977 9122 16011
rect 9088 15909 9122 15943
rect 9088 15841 9122 15875
rect 9088 15773 9122 15807
rect 9088 15705 9122 15739
rect 9088 15637 9122 15671
rect 9088 15569 9122 15603
rect 9088 15501 9122 15535
rect 9088 15433 9122 15467
rect 9088 15365 9122 15399
rect 9088 15297 9122 15331
rect 9088 15229 9122 15263
rect 9088 15161 9122 15195
rect 9088 15093 9122 15127
rect 9088 15025 9122 15059
rect 9088 14957 9122 14991
rect 9088 14889 9122 14923
rect 9088 14821 9122 14855
rect 9088 14753 9122 14787
rect 9088 14685 9122 14719
rect 9088 14617 9122 14651
rect 9088 14549 9122 14583
rect 9088 14481 9122 14515
rect 9088 14413 9122 14447
rect 9088 14345 9122 14379
rect 9088 14277 9122 14311
rect 9088 14209 9122 14243
rect 9088 14141 9122 14175
rect 9088 14073 9122 14107
rect 9088 14005 9122 14039
rect 9088 13937 9122 13971
rect 9088 13869 9122 13903
rect 9088 13801 9122 13835
rect 9088 13733 9122 13767
rect 9088 13665 9122 13699
rect 9088 13597 9122 13631
rect 9088 13529 9122 13563
rect 9088 13461 9122 13495
rect 9088 13393 9122 13427
rect 9088 13325 9122 13359
rect 9088 13257 9122 13291
rect 9088 13189 9122 13223
rect 9088 13121 9122 13155
rect 9088 13053 9122 13087
rect 9088 12985 9122 13019
rect 9088 12917 9122 12951
rect 9088 12849 9122 12883
rect 9088 12781 9122 12815
rect 9088 12713 9122 12747
rect 9088 12645 9122 12679
rect 9088 12577 9122 12611
rect 9088 12509 9122 12543
rect 9088 12441 9122 12475
rect 9088 12373 9122 12407
rect 9088 12305 9122 12339
rect 9088 12237 9122 12271
rect 9088 12169 9122 12203
rect 9088 12101 9122 12135
rect 9088 12033 9122 12067
rect 9088 11965 9122 11999
rect 9088 11897 9122 11931
rect 9088 11829 9122 11863
rect 9088 11761 9122 11795
rect 9088 11693 9122 11727
rect 9088 11625 9122 11659
rect 9088 11557 9122 11591
rect 9088 11489 9122 11523
rect 9088 11421 9122 11455
rect 9088 11353 9122 11387
rect 9088 11285 9122 11319
rect 9088 11217 9122 11251
rect 9088 11149 9122 11183
rect 9088 11081 9122 11115
rect 9088 11013 9122 11047
rect 9088 10945 9122 10979
rect 9088 10877 9122 10911
rect 9088 10809 9122 10843
rect 9088 10741 9122 10775
rect 9088 10673 9122 10707
rect 9088 10605 9122 10639
rect 9088 10537 9122 10571
rect 9088 10469 9122 10503
rect 9088 10401 9122 10435
rect 9088 10333 9122 10367
rect 9088 10265 9122 10299
rect 9088 10197 9122 10231
rect 9088 10129 9122 10163
rect 9088 10061 9122 10095
rect 9088 9993 9122 10027
rect 9088 9925 9122 9959
rect 9088 9857 9122 9891
rect 9088 9789 9122 9823
rect 9088 9721 9122 9755
rect 9088 9653 9122 9687
rect 9088 9585 9122 9619
rect 9088 9517 9122 9551
rect 9088 9449 9122 9483
rect 9088 9381 9122 9415
rect 9088 9313 9122 9347
rect 9088 9245 9122 9279
rect 9088 9177 9122 9211
rect 9088 9109 9122 9143
rect 9088 9041 9122 9075
rect 9088 8973 9122 9007
rect 9088 8905 9122 8939
rect 9088 8837 9122 8871
rect 9088 8769 9122 8803
rect 9088 8701 9122 8735
rect 9088 8633 9122 8667
rect 9088 8565 9122 8599
rect 9088 8497 9122 8531
rect 9088 8429 9122 8463
rect 9088 8361 9122 8395
rect 9088 8293 9122 8327
rect 9088 8225 9122 8259
rect 9088 8157 9122 8191
rect 9088 8089 9122 8123
rect 9088 8021 9122 8055
rect 9088 7953 9122 7987
rect 9088 7885 9122 7919
rect 9088 7817 9122 7851
rect 9088 7749 9122 7783
rect 9088 7681 9122 7715
rect 9088 7613 9122 7647
rect 9088 7545 9122 7579
rect 9088 7477 9122 7511
rect 9088 7409 9122 7443
rect 9088 7341 9122 7375
rect 9088 7273 9122 7307
rect 9088 7205 9122 7239
rect 9088 7137 9122 7171
rect 9088 7069 9122 7103
rect 9088 7001 9122 7035
rect 9088 6933 9122 6967
rect 9088 6865 9122 6899
rect 9088 6797 9122 6831
rect 9088 6729 9122 6763
rect 9088 6661 9122 6695
rect 9088 6593 9122 6627
rect 9088 6525 9122 6559
rect 9088 6457 9122 6491
rect 9088 6389 9122 6423
rect 9088 6321 9122 6355
rect 9088 6253 9122 6287
rect 9088 6185 9122 6219
rect 9088 6117 9122 6151
rect 9088 6049 9122 6083
rect 9088 5981 9122 6015
rect 9088 5913 9122 5947
rect 9088 5845 9122 5879
rect 9088 5777 9122 5811
rect 9088 5709 9122 5743
rect 9088 5641 9122 5675
rect 9088 5573 9122 5607
rect 9088 5505 9122 5539
rect 9088 5437 9122 5471
rect 9088 5369 9122 5403
rect 9088 5301 9122 5335
rect 9088 5233 9122 5267
rect 9088 5165 9122 5199
rect 9088 5097 9122 5131
rect 9088 5029 9122 5063
rect 9088 4961 9122 4995
rect 9088 4893 9122 4927
rect 9088 4825 9122 4859
rect 9088 4757 9122 4791
rect 9088 4689 9122 4723
rect 9088 4621 9122 4655
rect 9088 4553 9122 4587
rect 9088 4485 9122 4519
rect 9088 4417 9122 4451
rect 9088 4349 9122 4383
rect 9088 4281 9122 4315
rect 9088 4213 9122 4247
rect 9088 4145 9122 4179
rect 9088 4077 9122 4111
rect 9088 4009 9122 4043
rect 9088 3941 9122 3975
rect 9088 3873 9122 3907
rect 9088 3805 9122 3839
rect 9088 3737 9122 3771
rect 9088 3669 9122 3703
rect 9088 3601 9122 3635
rect 9088 3533 9122 3567
rect 9088 3465 9122 3499
rect 10226 38641 10260 38723
rect 10226 38573 10260 38607
rect 10226 38505 10260 38539
rect 10226 38437 10260 38471
rect 10226 38369 10260 38403
rect 10226 38301 10260 38335
rect 10226 38233 10260 38267
rect 10226 38165 10260 38199
rect 10226 38097 10260 38131
rect 10226 38029 10260 38063
rect 10226 37961 10260 37995
rect 10226 37893 10260 37927
rect 10226 37825 10260 37859
rect 10226 37757 10260 37791
rect 10226 37689 10260 37723
rect 10226 37621 10260 37655
rect 10226 37553 10260 37587
rect 10226 37485 10260 37519
rect 10226 37417 10260 37451
rect 10226 37349 10260 37383
rect 10226 37281 10260 37315
rect 10226 37213 10260 37247
rect 10226 37145 10260 37179
rect 10226 37077 10260 37111
rect 10226 37009 10260 37043
rect 10226 36941 10260 36975
rect 10226 36873 10260 36907
rect 10226 36805 10260 36839
rect 10226 36737 10260 36771
rect 10226 36669 10260 36703
rect 10226 36601 10260 36635
rect 10226 36533 10260 36567
rect 10226 36465 10260 36499
rect 10226 36397 10260 36431
rect 10226 36329 10260 36363
rect 10226 36261 10260 36295
rect 10226 36193 10260 36227
rect 10226 36125 10260 36159
rect 10226 36057 10260 36091
rect 10226 35989 10260 36023
rect 10226 35921 10260 35955
rect 10226 35853 10260 35887
rect 10226 35785 10260 35819
rect 10226 35717 10260 35751
rect 10226 35649 10260 35683
rect 10226 35581 10260 35615
rect 10226 35513 10260 35547
rect 10226 35445 10260 35479
rect 10226 35377 10260 35411
rect 10226 35309 10260 35343
rect 10226 35241 10260 35275
rect 10226 35173 10260 35207
rect 10226 35105 10260 35139
rect 10226 35037 10260 35071
rect 10226 34969 10260 35003
rect 10226 34901 10260 34935
rect 10226 34833 10260 34867
rect 10226 34765 10260 34799
rect 10226 34697 10260 34731
rect 10226 34629 10260 34663
rect 10226 34561 10260 34595
rect 10226 34493 10260 34527
rect 10226 34425 10260 34459
rect 10226 34357 10260 34391
rect 10226 34289 10260 34323
rect 10226 34221 10260 34255
rect 10226 34153 10260 34187
rect 10226 34085 10260 34119
rect 10226 34017 10260 34051
rect 10226 33949 10260 33983
rect 10226 33881 10260 33915
rect 10226 33813 10260 33847
rect 10226 33745 10260 33779
rect 10226 33677 10260 33711
rect 10226 33609 10260 33643
rect 10226 33541 10260 33575
rect 10226 33473 10260 33507
rect 10226 33405 10260 33439
rect 10226 33337 10260 33371
rect 10226 33269 10260 33303
rect 10226 33201 10260 33235
rect 10226 33133 10260 33167
rect 10226 33065 10260 33099
rect 10226 32997 10260 33031
rect 10226 32929 10260 32963
rect 10226 32861 10260 32895
rect 10226 32793 10260 32827
rect 10226 32725 10260 32759
rect 10226 32657 10260 32691
rect 10226 32589 10260 32623
rect 10226 32521 10260 32555
rect 10226 32453 10260 32487
rect 10226 32385 10260 32419
rect 10226 32317 10260 32351
rect 10226 32249 10260 32283
rect 10226 32181 10260 32215
rect 10226 32113 10260 32147
rect 10226 32045 10260 32079
rect 10226 31977 10260 32011
rect 10226 31909 10260 31943
rect 10226 31841 10260 31875
rect 10226 31773 10260 31807
rect 10226 31705 10260 31739
rect 10226 31637 10260 31671
rect 10226 31569 10260 31603
rect 10226 31501 10260 31535
rect 10226 31433 10260 31467
rect 10226 31365 10260 31399
rect 10226 31297 10260 31331
rect 10226 31229 10260 31263
rect 10226 31161 10260 31195
rect 10226 31093 10260 31127
rect 10226 31025 10260 31059
rect 10226 30957 10260 30991
rect 10226 30889 10260 30923
rect 10226 30821 10260 30855
rect 10226 30753 10260 30787
rect 10226 30685 10260 30719
rect 10226 30617 10260 30651
rect 10226 30549 10260 30583
rect 10226 30481 10260 30515
rect 10226 30413 10260 30447
rect 10226 30345 10260 30379
rect 10226 30277 10260 30311
rect 10226 30209 10260 30243
rect 10226 30141 10260 30175
rect 10226 30073 10260 30107
rect 10226 30005 10260 30039
rect 10226 29937 10260 29971
rect 10226 29869 10260 29903
rect 10226 29801 10260 29835
rect 10226 29733 10260 29767
rect 10226 29665 10260 29699
rect 10226 29597 10260 29631
rect 10226 29529 10260 29563
rect 10226 29461 10260 29495
rect 10226 29393 10260 29427
rect 10226 29325 10260 29359
rect 10226 29257 10260 29291
rect 10226 29189 10260 29223
rect 10226 29121 10260 29155
rect 10226 29053 10260 29087
rect 10226 28985 10260 29019
rect 10226 28917 10260 28951
rect 10226 28849 10260 28883
rect 10226 28781 10260 28815
rect 10226 28713 10260 28747
rect 10226 28645 10260 28679
rect 10226 28577 10260 28611
rect 10226 28509 10260 28543
rect 10226 28441 10260 28475
rect 10226 28373 10260 28407
rect 10226 28305 10260 28339
rect 10226 28237 10260 28271
rect 10226 28169 10260 28203
rect 10226 28101 10260 28135
rect 10226 28033 10260 28067
rect 10226 27965 10260 27999
rect 10226 27897 10260 27931
rect 10226 27829 10260 27863
rect 10226 27761 10260 27795
rect 10226 27693 10260 27727
rect 10226 27625 10260 27659
rect 10226 27557 10260 27591
rect 10226 27489 10260 27523
rect 10226 27421 10260 27455
rect 10226 27353 10260 27387
rect 10226 27285 10260 27319
rect 10226 27217 10260 27251
rect 10226 27149 10260 27183
rect 10226 27081 10260 27115
rect 10226 27013 10260 27047
rect 10226 26945 10260 26979
rect 10226 26877 10260 26911
rect 10226 26809 10260 26843
rect 10226 26741 10260 26775
rect 10226 26673 10260 26707
rect 10226 26605 10260 26639
rect 10226 26537 10260 26571
rect 10226 26469 10260 26503
rect 10226 26401 10260 26435
rect 10226 26333 10260 26367
rect 10226 26265 10260 26299
rect 10226 26197 10260 26231
rect 10226 26129 10260 26163
rect 10226 26061 10260 26095
rect 10226 25993 10260 26027
rect 10226 25925 10260 25959
rect 10226 25857 10260 25891
rect 10226 25789 10260 25823
rect 10226 25721 10260 25755
rect 10226 25653 10260 25687
rect 10226 25585 10260 25619
rect 10226 25517 10260 25551
rect 10226 25449 10260 25483
rect 10226 25381 10260 25415
rect 10226 25313 10260 25347
rect 10226 25245 10260 25279
rect 10226 25177 10260 25211
rect 10226 25109 10260 25143
rect 10226 25041 10260 25075
rect 10226 24973 10260 25007
rect 10226 24905 10260 24939
rect 10226 24837 10260 24871
rect 10226 24769 10260 24803
rect 10226 24701 10260 24735
rect 10226 24633 10260 24667
rect 10226 24565 10260 24599
rect 10226 24497 10260 24531
rect 10226 24429 10260 24463
rect 10226 24361 10260 24395
rect 10226 24293 10260 24327
rect 10226 24225 10260 24259
rect 10226 24157 10260 24191
rect 10226 24089 10260 24123
rect 10226 24021 10260 24055
rect 10226 23953 10260 23987
rect 10226 23885 10260 23919
rect 10226 23817 10260 23851
rect 10226 23749 10260 23783
rect 10226 23681 10260 23715
rect 10226 23613 10260 23647
rect 10226 23545 10260 23579
rect 10226 23477 10260 23511
rect 10226 23409 10260 23443
rect 10226 23341 10260 23375
rect 10226 23273 10260 23307
rect 10226 23205 10260 23239
rect 10226 23137 10260 23171
rect 10226 23069 10260 23103
rect 10226 23001 10260 23035
rect 10226 22933 10260 22967
rect 10226 22865 10260 22899
rect 10226 22797 10260 22831
rect 10226 22729 10260 22763
rect 10226 22661 10260 22695
rect 10226 22593 10260 22627
rect 10226 22525 10260 22559
rect 10226 22457 10260 22491
rect 10226 22389 10260 22423
rect 10226 22321 10260 22355
rect 10226 22253 10260 22287
rect 10226 22185 10260 22219
rect 10226 22117 10260 22151
rect 10226 22049 10260 22083
rect 10226 21981 10260 22015
rect 10226 21913 10260 21947
rect 10226 21845 10260 21879
rect 10226 21777 10260 21811
rect 10226 21709 10260 21743
rect 10226 21641 10260 21675
rect 10226 21573 10260 21607
rect 10226 21505 10260 21539
rect 10226 21437 10260 21471
rect 10226 21369 10260 21403
rect 10226 21301 10260 21335
rect 10226 21233 10260 21267
rect 10226 21165 10260 21199
rect 10226 21097 10260 21131
rect 10226 21029 10260 21063
rect 10226 20961 10260 20995
rect 10226 20893 10260 20927
rect 10226 20825 10260 20859
rect 10226 20757 10260 20791
rect 10226 20689 10260 20723
rect 10226 20621 10260 20655
rect 10226 20553 10260 20587
rect 10226 20485 10260 20519
rect 10226 20417 10260 20451
rect 10226 20349 10260 20383
rect 10226 20281 10260 20315
rect 10226 20213 10260 20247
rect 10226 20145 10260 20179
rect 10226 20077 10260 20111
rect 10226 20009 10260 20043
rect 10226 19941 10260 19975
rect 10226 19873 10260 19907
rect 10226 19805 10260 19839
rect 10226 19737 10260 19771
rect 10226 19669 10260 19703
rect 10226 19601 10260 19635
rect 10226 19533 10260 19567
rect 10226 19465 10260 19499
rect 10226 19397 10260 19431
rect 10226 19329 10260 19363
rect 10226 19261 10260 19295
rect 10226 19193 10260 19227
rect 10226 19125 10260 19159
rect 10226 19057 10260 19091
rect 10226 18989 10260 19023
rect 10226 18921 10260 18955
rect 10226 18853 10260 18887
rect 10226 18785 10260 18819
rect 10226 18717 10260 18751
rect 10226 18649 10260 18683
rect 10226 18581 10260 18615
rect 10226 18513 10260 18547
rect 10226 18445 10260 18479
rect 10226 18377 10260 18411
rect 10226 18309 10260 18343
rect 10226 18241 10260 18275
rect 10226 18173 10260 18207
rect 10226 18105 10260 18139
rect 10226 18037 10260 18071
rect 10226 17969 10260 18003
rect 10226 17901 10260 17935
rect 10226 17833 10260 17867
rect 10226 17765 10260 17799
rect 10226 17697 10260 17731
rect 10226 17629 10260 17663
rect 10226 17561 10260 17595
rect 10226 17493 10260 17527
rect 10226 17425 10260 17459
rect 10226 17357 10260 17391
rect 10226 17289 10260 17323
rect 10226 17221 10260 17255
rect 10226 17153 10260 17187
rect 10226 17085 10260 17119
rect 10226 17017 10260 17051
rect 10226 16949 10260 16983
rect 10226 16881 10260 16915
rect 10226 16813 10260 16847
rect 10226 16745 10260 16779
rect 10226 16677 10260 16711
rect 10226 16609 10260 16643
rect 10226 16541 10260 16575
rect 10226 16473 10260 16507
rect 10226 16405 10260 16439
rect 10226 16337 10260 16371
rect 10226 16269 10260 16303
rect 10226 16201 10260 16235
rect 10226 16133 10260 16167
rect 10226 16065 10260 16099
rect 10226 15997 10260 16031
rect 10226 15929 10260 15963
rect 10226 15861 10260 15895
rect 10226 15793 10260 15827
rect 10226 15725 10260 15759
rect 10226 15657 10260 15691
rect 10226 15589 10260 15623
rect 10226 15521 10260 15555
rect 10226 15453 10260 15487
rect 10226 15385 10260 15419
rect 10226 15317 10260 15351
rect 10226 15249 10260 15283
rect 10226 15181 10260 15215
rect 10226 15113 10260 15147
rect 10226 15045 10260 15079
rect 10226 14977 10260 15011
rect 10226 14909 10260 14943
rect 10226 14841 10260 14875
rect 10226 14773 10260 14807
rect 10226 14705 10260 14739
rect 10226 14637 10260 14671
rect 10226 14569 10260 14603
rect 10226 14501 10260 14535
rect 10226 14433 10260 14467
rect 10226 14365 10260 14399
rect 10226 14297 10260 14331
rect 10226 14229 10260 14263
rect 10226 14161 10260 14195
rect 10226 14093 10260 14127
rect 10226 14025 10260 14059
rect 10226 13957 10260 13991
rect 10226 13889 10260 13923
rect 10226 13821 10260 13855
rect 10226 13753 10260 13787
rect 10226 13685 10260 13719
rect 10226 13617 10260 13651
rect 10226 13549 10260 13583
rect 10226 13481 10260 13515
rect 10226 13413 10260 13447
rect 10226 13345 10260 13379
rect 10226 13277 10260 13311
rect 10226 13209 10260 13243
rect 10226 13141 10260 13175
rect 10226 13073 10260 13107
rect 10226 13005 10260 13039
rect 10226 12937 10260 12971
rect 10226 12869 10260 12903
rect 10226 12801 10260 12835
rect 10226 12733 10260 12767
rect 10226 12665 10260 12699
rect 10226 12597 10260 12631
rect 10226 12529 10260 12563
rect 10226 12461 10260 12495
rect 10226 12393 10260 12427
rect 10226 12325 10260 12359
rect 10226 12257 10260 12291
rect 10226 12189 10260 12223
rect 10226 12121 10260 12155
rect 10226 12053 10260 12087
rect 10226 11985 10260 12019
rect 10226 11917 10260 11951
rect 10226 11849 10260 11883
rect 10226 11781 10260 11815
rect 10226 11713 10260 11747
rect 10226 11645 10260 11679
rect 10226 11577 10260 11611
rect 10226 11509 10260 11543
rect 10226 11441 10260 11475
rect 10226 11373 10260 11407
rect 10226 11305 10260 11339
rect 10226 11237 10260 11271
rect 10226 11169 10260 11203
rect 10226 11101 10260 11135
rect 10226 11033 10260 11067
rect 10226 10965 10260 10999
rect 10226 10897 10260 10931
rect 10226 10829 10260 10863
rect 10226 10761 10260 10795
rect 10226 10693 10260 10727
rect 10226 10625 10260 10659
rect 10226 10557 10260 10591
rect 10226 10489 10260 10523
rect 10226 10421 10260 10455
rect 10226 10353 10260 10387
rect 10226 10285 10260 10319
rect 10226 10217 10260 10251
rect 10226 10149 10260 10183
rect 10226 10081 10260 10115
rect 10226 10013 10260 10047
rect 10226 9945 10260 9979
rect 10226 9877 10260 9911
rect 10226 9809 10260 9843
rect 10226 9741 10260 9775
rect 10226 9673 10260 9707
rect 10226 9605 10260 9639
rect 10226 9537 10260 9571
rect 10226 9469 10260 9503
rect 10226 9401 10260 9435
rect 10226 9333 10260 9367
rect 10226 9265 10260 9299
rect 10226 9197 10260 9231
rect 10226 9129 10260 9163
rect 10226 9061 10260 9095
rect 10226 8993 10260 9027
rect 10226 8925 10260 8959
rect 10226 8857 10260 8891
rect 10226 8789 10260 8823
rect 10226 8721 10260 8755
rect 10226 8653 10260 8687
rect 10226 8585 10260 8619
rect 10226 8517 10260 8551
rect 10226 8449 10260 8483
rect 10226 8381 10260 8415
rect 10226 8313 10260 8347
rect 10226 8245 10260 8279
rect 10226 8177 10260 8211
rect 10226 8109 10260 8143
rect 10226 8041 10260 8075
rect 10226 7973 10260 8007
rect 10226 7905 10260 7939
rect 10226 7837 10260 7871
rect 10226 7769 10260 7803
rect 10226 7701 10260 7735
rect 10226 7633 10260 7667
rect 10226 7565 10260 7599
rect 10226 7497 10260 7531
rect 10226 7429 10260 7463
rect 10226 7361 10260 7395
rect 10226 7293 10260 7327
rect 10226 7225 10260 7259
rect 10226 7157 10260 7191
rect 10226 7089 10260 7123
rect 10226 7021 10260 7055
rect 10226 6953 10260 6987
rect 10226 6885 10260 6919
rect 10226 6817 10260 6851
rect 10226 6749 10260 6783
rect 10226 6681 10260 6715
rect 10226 6613 10260 6647
rect 10226 6545 10260 6579
rect 10226 6477 10260 6511
rect 10226 6409 10260 6443
rect 10226 6341 10260 6375
rect 10226 6273 10260 6307
rect 10226 6205 10260 6239
rect 10226 6137 10260 6171
rect 10226 6069 10260 6103
rect 10226 6001 10260 6035
rect 10226 5933 10260 5967
rect 10226 5865 10260 5899
rect 10226 5797 10260 5831
rect 10226 5729 10260 5763
rect 10226 5661 10260 5695
rect 10226 5593 10260 5627
rect 10226 5525 10260 5559
rect 10226 5457 10260 5491
rect 10226 5389 10260 5423
rect 10226 5321 10260 5355
rect 10226 5253 10260 5287
rect 10226 5185 10260 5219
rect 10226 5117 10260 5151
rect 10226 5049 10260 5083
rect 10226 4981 10260 5015
rect 10226 4913 10260 4947
rect 10226 4845 10260 4879
rect 10226 4777 10260 4811
rect 10226 4709 10260 4743
rect 10226 4641 10260 4675
rect 10226 4573 10260 4607
rect 10226 4505 10260 4539
rect 10226 4437 10260 4471
rect 10226 4369 10260 4403
rect 10226 4301 10260 4335
rect 10226 4233 10260 4267
rect 10226 4165 10260 4199
rect 10226 4097 10260 4131
rect 10226 4029 10260 4063
rect 10226 3961 10260 3995
rect 10226 3893 10260 3927
rect 10226 3825 10260 3859
rect 10226 3757 10260 3791
rect 10226 3689 10260 3723
rect 10226 3621 10260 3655
rect 10226 3553 10260 3587
rect 10226 3485 10260 3519
rect 9088 3397 9122 3431
rect 9088 3329 9122 3363
rect 11424 38689 11458 38723
rect 11424 38621 11458 38655
rect 11424 38553 11458 38587
rect 11424 38485 11458 38519
rect 13212 38630 13246 38723
rect 14940 38689 14974 38723
rect 13212 38562 13246 38596
rect 11424 38417 11458 38451
rect 11424 38349 11458 38383
rect 11424 38281 11458 38315
rect 11424 38213 11458 38247
rect 11424 38145 11458 38179
rect 11424 38077 11458 38111
rect 11424 38009 11458 38043
rect 11424 37941 11458 37975
rect 11424 37873 11458 37907
rect 11424 37805 11458 37839
rect 11424 37737 11458 37771
rect 11424 37669 11458 37703
rect 11424 37601 11458 37635
rect 11424 37533 11458 37567
rect 11424 37465 11458 37499
rect 11424 37397 11458 37431
rect 11424 37329 11458 37363
rect 11424 37261 11458 37295
rect 11424 37193 11458 37227
rect 11424 37125 11458 37159
rect 11424 37057 11458 37091
rect 11424 36989 11458 37023
rect 11424 36921 11458 36955
rect 11424 36853 11458 36887
rect 11424 36785 11458 36819
rect 11424 36717 11458 36751
rect 11424 36649 11458 36683
rect 11424 36581 11458 36615
rect 11424 36513 11458 36547
rect 11424 36445 11458 36479
rect 11424 36377 11458 36411
rect 11424 36309 11458 36343
rect 11424 36241 11458 36275
rect 11424 36173 11458 36207
rect 11424 36105 11458 36139
rect 11424 36037 11458 36071
rect 11424 35969 11458 36003
rect 11424 35901 11458 35935
rect 11424 35833 11458 35867
rect 11424 35765 11458 35799
rect 11424 35697 11458 35731
rect 11424 35629 11458 35663
rect 11424 35561 11458 35595
rect 11424 35493 11458 35527
rect 11424 35425 11458 35459
rect 11424 35357 11458 35391
rect 11424 35289 11458 35323
rect 11424 35221 11458 35255
rect 11424 35153 11458 35187
rect 11424 35085 11458 35119
rect 11424 35017 11458 35051
rect 11424 34949 11458 34983
rect 11424 34881 11458 34915
rect 11424 34813 11458 34847
rect 11424 34745 11458 34779
rect 11424 34677 11458 34711
rect 11424 34609 11458 34643
rect 11424 34541 11458 34575
rect 11424 34473 11458 34507
rect 11424 34405 11458 34439
rect 11424 34337 11458 34371
rect 11424 34269 11458 34303
rect 11424 34201 11458 34235
rect 11424 34133 11458 34167
rect 11424 34065 11458 34099
rect 11424 33997 11458 34031
rect 11424 33929 11458 33963
rect 11424 33861 11458 33895
rect 11424 33793 11458 33827
rect 11424 33725 11458 33759
rect 11424 33657 11458 33691
rect 11424 33589 11458 33623
rect 11424 33521 11458 33555
rect 11424 33453 11458 33487
rect 11424 33385 11458 33419
rect 11424 33317 11458 33351
rect 11424 33249 11458 33283
rect 11424 33181 11458 33215
rect 11424 33113 11458 33147
rect 11424 33045 11458 33079
rect 11424 32977 11458 33011
rect 11424 32909 11458 32943
rect 11424 32841 11458 32875
rect 11424 32773 11458 32807
rect 11424 32705 11458 32739
rect 11424 32637 11458 32671
rect 11424 32569 11458 32603
rect 11424 32501 11458 32535
rect 11424 32433 11458 32467
rect 11424 32365 11458 32399
rect 11424 32297 11458 32331
rect 11424 32229 11458 32263
rect 11424 32161 11458 32195
rect 11424 32093 11458 32127
rect 11424 32025 11458 32059
rect 11424 31957 11458 31991
rect 11424 31889 11458 31923
rect 11424 31821 11458 31855
rect 11424 31753 11458 31787
rect 11424 31685 11458 31719
rect 11424 31617 11458 31651
rect 11424 31549 11458 31583
rect 11424 31481 11458 31515
rect 11424 31413 11458 31447
rect 11424 31345 11458 31379
rect 11424 31277 11458 31311
rect 11424 31209 11458 31243
rect 11424 31141 11458 31175
rect 11424 31073 11458 31107
rect 11424 31005 11458 31039
rect 11424 30937 11458 30971
rect 11424 30869 11458 30903
rect 11424 30801 11458 30835
rect 11424 30733 11458 30767
rect 11424 30665 11458 30699
rect 11424 30597 11458 30631
rect 11424 30529 11458 30563
rect 11424 30461 11458 30495
rect 11424 30393 11458 30427
rect 11424 30325 11458 30359
rect 11424 30257 11458 30291
rect 11424 30189 11458 30223
rect 11424 30121 11458 30155
rect 11424 30053 11458 30087
rect 11424 29985 11458 30019
rect 11424 29917 11458 29951
rect 11424 29849 11458 29883
rect 11424 29781 11458 29815
rect 11424 29713 11458 29747
rect 11424 29645 11458 29679
rect 11424 29577 11458 29611
rect 11424 29509 11458 29543
rect 11424 29441 11458 29475
rect 11424 29373 11458 29407
rect 11424 29305 11458 29339
rect 11424 29237 11458 29271
rect 11424 29169 11458 29203
rect 11424 29101 11458 29135
rect 11424 29033 11458 29067
rect 11424 28965 11458 28999
rect 11424 28897 11458 28931
rect 11424 28829 11458 28863
rect 11424 28761 11458 28795
rect 11424 28693 11458 28727
rect 11424 28625 11458 28659
rect 11424 28557 11458 28591
rect 11424 28489 11458 28523
rect 11424 28421 11458 28455
rect 11424 28353 11458 28387
rect 11424 28285 11458 28319
rect 11424 28217 11458 28251
rect 11424 28149 11458 28183
rect 11424 28081 11458 28115
rect 11424 28013 11458 28047
rect 11424 27945 11458 27979
rect 11424 27877 11458 27911
rect 11424 27809 11458 27843
rect 11424 27741 11458 27775
rect 11424 27673 11458 27707
rect 11424 27605 11458 27639
rect 11424 27537 11458 27571
rect 11424 27469 11458 27503
rect 11424 27401 11458 27435
rect 11424 27333 11458 27367
rect 11424 27265 11458 27299
rect 11424 27197 11458 27231
rect 11424 27129 11458 27163
rect 11424 27061 11458 27095
rect 11424 26993 11458 27027
rect 11424 26925 11458 26959
rect 11424 26857 11458 26891
rect 11424 26789 11458 26823
rect 11424 26721 11458 26755
rect 11424 26653 11458 26687
rect 11424 26585 11458 26619
rect 11424 26517 11458 26551
rect 11424 26449 11458 26483
rect 11424 26381 11458 26415
rect 11424 26313 11458 26347
rect 11424 26245 11458 26279
rect 11424 26177 11458 26211
rect 11424 26109 11458 26143
rect 11424 26041 11458 26075
rect 11424 25973 11458 26007
rect 11424 25905 11458 25939
rect 11424 25837 11458 25871
rect 11424 25769 11458 25803
rect 11424 25701 11458 25735
rect 11424 25633 11458 25667
rect 11424 25565 11458 25599
rect 11424 25497 11458 25531
rect 11424 25429 11458 25463
rect 11424 25361 11458 25395
rect 11424 25293 11458 25327
rect 11424 25225 11458 25259
rect 11424 25157 11458 25191
rect 11424 25089 11458 25123
rect 11424 25021 11458 25055
rect 11424 24953 11458 24987
rect 11424 24885 11458 24919
rect 11424 24817 11458 24851
rect 11424 24749 11458 24783
rect 11424 24681 11458 24715
rect 11424 24613 11458 24647
rect 11424 24545 11458 24579
rect 11424 24477 11458 24511
rect 11424 24409 11458 24443
rect 11424 24341 11458 24375
rect 11424 24273 11458 24307
rect 11424 24205 11458 24239
rect 11424 24137 11458 24171
rect 11424 24069 11458 24103
rect 11424 24001 11458 24035
rect 11424 23933 11458 23967
rect 11424 23865 11458 23899
rect 11424 23797 11458 23831
rect 11424 23729 11458 23763
rect 11424 23661 11458 23695
rect 11424 23593 11458 23627
rect 11424 23525 11458 23559
rect 11424 23457 11458 23491
rect 11424 23389 11458 23423
rect 11424 23321 11458 23355
rect 11424 23253 11458 23287
rect 11424 23185 11458 23219
rect 11424 23117 11458 23151
rect 11424 23049 11458 23083
rect 11424 22981 11458 23015
rect 11424 22913 11458 22947
rect 11424 22845 11458 22879
rect 11424 22777 11458 22811
rect 11424 22709 11458 22743
rect 11424 22641 11458 22675
rect 11424 22573 11458 22607
rect 11424 22505 11458 22539
rect 11424 22437 11458 22471
rect 11424 22369 11458 22403
rect 11424 22301 11458 22335
rect 11424 22233 11458 22267
rect 11424 22165 11458 22199
rect 11424 22097 11458 22131
rect 11424 22029 11458 22063
rect 11424 21961 11458 21995
rect 11424 21893 11458 21927
rect 11424 21825 11458 21859
rect 11424 21757 11458 21791
rect 11424 21689 11458 21723
rect 11424 21621 11458 21655
rect 11424 21553 11458 21587
rect 11424 21485 11458 21519
rect 11424 21417 11458 21451
rect 11424 21349 11458 21383
rect 11424 21281 11458 21315
rect 11424 21213 11458 21247
rect 11424 21145 11458 21179
rect 11424 21077 11458 21111
rect 11424 21009 11458 21043
rect 11424 20941 11458 20975
rect 11424 20873 11458 20907
rect 11424 20805 11458 20839
rect 11424 20737 11458 20771
rect 11424 20669 11458 20703
rect 11424 20601 11458 20635
rect 11424 20533 11458 20567
rect 11424 20465 11458 20499
rect 11424 20397 11458 20431
rect 11424 20329 11458 20363
rect 11424 20261 11458 20295
rect 11424 20193 11458 20227
rect 11424 20125 11458 20159
rect 11424 20057 11458 20091
rect 11424 19989 11458 20023
rect 11424 19921 11458 19955
rect 11424 19853 11458 19887
rect 11424 19785 11458 19819
rect 11424 19717 11458 19751
rect 11424 19649 11458 19683
rect 11424 19581 11458 19615
rect 11424 19513 11458 19547
rect 11424 19445 11458 19479
rect 11424 19377 11458 19411
rect 11424 19309 11458 19343
rect 11424 19241 11458 19275
rect 11424 19173 11458 19207
rect 11424 19105 11458 19139
rect 11424 19037 11458 19071
rect 11424 18969 11458 19003
rect 11424 18901 11458 18935
rect 11424 18833 11458 18867
rect 11424 18765 11458 18799
rect 11424 18697 11458 18731
rect 11424 18629 11458 18663
rect 11424 18561 11458 18595
rect 11424 18493 11458 18527
rect 11424 18425 11458 18459
rect 11424 18357 11458 18391
rect 11424 18289 11458 18323
rect 11424 18221 11458 18255
rect 11424 18153 11458 18187
rect 11424 18085 11458 18119
rect 11424 18017 11458 18051
rect 11424 17949 11458 17983
rect 11424 17881 11458 17915
rect 11424 17813 11458 17847
rect 11424 17745 11458 17779
rect 11424 17677 11458 17711
rect 11424 17609 11458 17643
rect 11424 17541 11458 17575
rect 11424 17473 11458 17507
rect 11424 17405 11458 17439
rect 11424 17337 11458 17371
rect 11424 17269 11458 17303
rect 11424 17201 11458 17235
rect 11424 17133 11458 17167
rect 11424 17065 11458 17099
rect 11424 16997 11458 17031
rect 11424 16929 11458 16963
rect 11424 16861 11458 16895
rect 11424 16793 11458 16827
rect 11424 16725 11458 16759
rect 11424 16657 11458 16691
rect 11424 16589 11458 16623
rect 11424 16521 11458 16555
rect 11424 16453 11458 16487
rect 11424 16385 11458 16419
rect 11424 16317 11458 16351
rect 11424 16249 11458 16283
rect 11424 16181 11458 16215
rect 11424 16113 11458 16147
rect 11424 16045 11458 16079
rect 11424 15977 11458 16011
rect 11424 15909 11458 15943
rect 11424 15841 11458 15875
rect 11424 15773 11458 15807
rect 11424 15705 11458 15739
rect 11424 15637 11458 15671
rect 11424 15569 11458 15603
rect 11424 15501 11458 15535
rect 11424 15433 11458 15467
rect 11424 15365 11458 15399
rect 11424 15297 11458 15331
rect 11424 15229 11458 15263
rect 11424 15161 11458 15195
rect 11424 15093 11458 15127
rect 11424 15025 11458 15059
rect 11424 14957 11458 14991
rect 11424 14889 11458 14923
rect 11424 14821 11458 14855
rect 11424 14753 11458 14787
rect 11424 14685 11458 14719
rect 11424 14617 11458 14651
rect 11424 14549 11458 14583
rect 11424 14481 11458 14515
rect 11424 14413 11458 14447
rect 11424 14345 11458 14379
rect 11424 14277 11458 14311
rect 11424 14209 11458 14243
rect 11424 14141 11458 14175
rect 11424 14073 11458 14107
rect 11424 14005 11458 14039
rect 11424 13937 11458 13971
rect 11424 13869 11458 13903
rect 11424 13801 11458 13835
rect 11424 13733 11458 13767
rect 11424 13665 11458 13699
rect 11424 13597 11458 13631
rect 11424 13529 11458 13563
rect 11424 13461 11458 13495
rect 11424 13393 11458 13427
rect 11424 13325 11458 13359
rect 11424 13257 11458 13291
rect 11424 13189 11458 13223
rect 11424 13121 11458 13155
rect 11424 13053 11458 13087
rect 11424 12985 11458 13019
rect 11424 12917 11458 12951
rect 11424 12849 11458 12883
rect 11424 12781 11458 12815
rect 11424 12713 11458 12747
rect 11424 12645 11458 12679
rect 11424 12577 11458 12611
rect 11424 12509 11458 12543
rect 11424 12441 11458 12475
rect 11424 12373 11458 12407
rect 11424 12305 11458 12339
rect 11424 12237 11458 12271
rect 11424 12169 11458 12203
rect 11424 12101 11458 12135
rect 11424 12033 11458 12067
rect 11424 11965 11458 11999
rect 11424 11897 11458 11931
rect 11424 11829 11458 11863
rect 11424 11761 11458 11795
rect 11424 11693 11458 11727
rect 11424 11625 11458 11659
rect 11424 11557 11458 11591
rect 11424 11489 11458 11523
rect 11424 11421 11458 11455
rect 11424 11353 11458 11387
rect 11424 11285 11458 11319
rect 11424 11217 11458 11251
rect 11424 11149 11458 11183
rect 11424 11081 11458 11115
rect 11424 11013 11458 11047
rect 11424 10945 11458 10979
rect 11424 10877 11458 10911
rect 11424 10809 11458 10843
rect 11424 10741 11458 10775
rect 11424 10673 11458 10707
rect 11424 10605 11458 10639
rect 11424 10537 11458 10571
rect 11424 10469 11458 10503
rect 11424 10401 11458 10435
rect 11424 10333 11458 10367
rect 11424 10265 11458 10299
rect 11424 10197 11458 10231
rect 11424 10129 11458 10163
rect 11424 10061 11458 10095
rect 11424 9993 11458 10027
rect 11424 9925 11458 9959
rect 11424 9857 11458 9891
rect 11424 9789 11458 9823
rect 11424 9721 11458 9755
rect 11424 9653 11458 9687
rect 11424 9585 11458 9619
rect 11424 9517 11458 9551
rect 11424 9449 11458 9483
rect 11424 9381 11458 9415
rect 11424 9313 11458 9347
rect 11424 9245 11458 9279
rect 11424 9177 11458 9211
rect 11424 9109 11458 9143
rect 11424 9041 11458 9075
rect 11424 8973 11458 9007
rect 11424 8905 11458 8939
rect 11424 8837 11458 8871
rect 11424 8769 11458 8803
rect 11424 8701 11458 8735
rect 11424 8633 11458 8667
rect 11424 8565 11458 8599
rect 11424 8497 11458 8531
rect 11424 8429 11458 8463
rect 11424 8361 11458 8395
rect 11424 8293 11458 8327
rect 11424 8225 11458 8259
rect 11424 8157 11458 8191
rect 11424 8089 11458 8123
rect 11424 8021 11458 8055
rect 11424 7953 11458 7987
rect 11424 7885 11458 7919
rect 11424 7817 11458 7851
rect 11424 7749 11458 7783
rect 11424 7681 11458 7715
rect 11424 7613 11458 7647
rect 11424 7545 11458 7579
rect 11424 7477 11458 7511
rect 11424 7409 11458 7443
rect 11424 7341 11458 7375
rect 11424 7273 11458 7307
rect 11424 7205 11458 7239
rect 11424 7137 11458 7171
rect 11424 7069 11458 7103
rect 11424 7001 11458 7035
rect 11424 6933 11458 6967
rect 11424 6865 11458 6899
rect 11424 6797 11458 6831
rect 11424 6729 11458 6763
rect 11424 6661 11458 6695
rect 11424 6593 11458 6627
rect 11424 6525 11458 6559
rect 11424 6457 11458 6491
rect 11424 6389 11458 6423
rect 11424 6321 11458 6355
rect 11424 6253 11458 6287
rect 11424 6185 11458 6219
rect 11424 6117 11458 6151
rect 11424 6049 11458 6083
rect 11424 5981 11458 6015
rect 11424 5913 11458 5947
rect 11424 5845 11458 5879
rect 11424 5777 11458 5811
rect 11424 5709 11458 5743
rect 11424 5641 11458 5675
rect 11424 5573 11458 5607
rect 11424 5505 11458 5539
rect 11424 5437 11458 5471
rect 11424 5369 11458 5403
rect 11424 5301 11458 5335
rect 11424 5233 11458 5267
rect 11424 5165 11458 5199
rect 11424 5097 11458 5131
rect 11424 5029 11458 5063
rect 11424 4961 11458 4995
rect 11424 4893 11458 4927
rect 11424 4825 11458 4859
rect 11424 4757 11458 4791
rect 11424 4689 11458 4723
rect 11424 4621 11458 4655
rect 11424 4553 11458 4587
rect 11424 4485 11458 4519
rect 11424 4417 11458 4451
rect 11424 4349 11458 4383
rect 11424 4281 11458 4315
rect 11424 4213 11458 4247
rect 11424 4145 11458 4179
rect 11424 4077 11458 4111
rect 11424 4009 11458 4043
rect 11424 3941 11458 3975
rect 11424 3873 11458 3907
rect 11424 3805 11458 3839
rect 11424 3737 11458 3771
rect 11424 3669 11458 3703
rect 11424 3601 11458 3635
rect 11424 3533 11458 3567
rect 10226 3417 10260 3451
rect 9088 3213 9122 3295
rect 10226 3349 10260 3383
rect 11424 3465 11458 3499
rect 11424 3397 11458 3431
rect 10226 3281 10260 3315
rect 10226 3213 10260 3247
rect 11424 3329 11458 3363
rect 11424 3213 11458 3295
rect 9088 3179 9156 3213
rect 9190 3179 9224 3213
rect 9258 3179 9292 3213
rect 9326 3179 9360 3213
rect 9394 3179 9428 3213
rect 9462 3179 9496 3213
rect 9530 3179 9564 3213
rect 9598 3179 9632 3213
rect 9666 3179 9700 3213
rect 9734 3179 9768 3213
rect 9802 3179 9836 3213
rect 9870 3179 9904 3213
rect 9938 3179 9972 3213
rect 10006 3179 10040 3213
rect 10074 3179 10108 3213
rect 10142 3179 10336 3213
rect 10370 3179 10404 3213
rect 10438 3179 10472 3213
rect 10506 3179 10540 3213
rect 10574 3179 10608 3213
rect 10642 3179 10676 3213
rect 10710 3179 10744 3213
rect 10778 3179 10812 3213
rect 10846 3179 10880 3213
rect 10914 3179 10948 3213
rect 10982 3179 11016 3213
rect 11050 3179 11084 3213
rect 11118 3179 11152 3213
rect 11186 3179 11220 3213
rect 11254 3179 11288 3213
rect 11322 3179 11356 3213
rect 11390 3205 11458 3213
rect 11390 3179 11424 3205
rect 11424 3137 11458 3171
rect 11424 3069 11458 3103
rect 11424 3001 11458 3035
rect 11424 2933 11458 2967
rect 11424 2865 11458 2899
rect 11424 2797 11458 2831
rect 11424 2729 11458 2763
rect 11424 2661 11458 2695
rect 11424 2593 11458 2627
rect 11424 2525 11458 2559
rect 11424 2457 11458 2491
rect 11424 2389 11458 2423
rect 11424 2321 11458 2355
rect 11424 2253 11458 2287
rect 11424 2185 11458 2219
rect 11424 2117 11458 2151
rect 11424 2049 11458 2083
rect 11424 1981 11458 2015
rect 11424 1913 11458 1947
rect 11424 1845 11458 1879
rect 11424 1777 11458 1811
rect 11424 1709 11458 1743
rect 11424 1641 11458 1675
rect 11424 1573 11458 1607
rect 11424 1505 11458 1539
rect 11424 1437 11458 1471
rect 11424 1369 11458 1403
rect 11424 1301 11458 1335
rect 11424 1233 11458 1267
rect 11424 1165 11458 1199
rect 11424 1097 11458 1131
rect 11424 1029 11458 1063
rect 11424 961 11458 995
rect 11424 893 11458 927
rect 11424 825 11458 859
rect 11424 757 11458 791
rect 11424 689 11458 723
rect 11424 621 11458 655
rect 11424 553 11458 587
rect 11424 485 11458 519
rect 11424 417 11458 451
rect 13212 38494 13246 38528
rect 14940 38621 14974 38655
rect 14940 38553 14974 38587
rect 13212 38426 13246 38460
rect 13212 38358 13246 38392
rect 13212 38290 13246 38324
rect 13212 38222 13246 38256
rect 13212 38154 13246 38188
rect 13212 38086 13246 38120
rect 13212 38018 13246 38052
rect 13212 37950 13246 37984
rect 13212 37882 13246 37916
rect 13212 37814 13246 37848
rect 13212 37746 13246 37780
rect 13212 37678 13246 37712
rect 13212 37610 13246 37644
rect 13212 37542 13246 37576
rect 13212 37474 13246 37508
rect 13212 37406 13246 37440
rect 13212 37338 13246 37372
rect 13212 37270 13246 37304
rect 13212 37202 13246 37236
rect 13212 37134 13246 37168
rect 13212 37066 13246 37100
rect 13212 36998 13246 37032
rect 13212 36930 13246 36964
rect 13212 36862 13246 36896
rect 13212 36794 13246 36828
rect 13212 36726 13246 36760
rect 13212 36658 13246 36692
rect 13212 36590 13246 36624
rect 13212 36522 13246 36556
rect 13212 36454 13246 36488
rect 13212 36386 13246 36420
rect 13212 36318 13246 36352
rect 13212 36250 13246 36284
rect 13212 36182 13246 36216
rect 13212 36114 13246 36148
rect 13212 36046 13246 36080
rect 13212 35978 13246 36012
rect 13212 35910 13246 35944
rect 13212 35842 13246 35876
rect 13212 35774 13246 35808
rect 13212 35706 13246 35740
rect 13212 35638 13246 35672
rect 13212 35570 13246 35604
rect 13212 35502 13246 35536
rect 13212 35434 13246 35468
rect 13212 35366 13246 35400
rect 13212 35298 13246 35332
rect 13212 35230 13246 35264
rect 13212 35162 13246 35196
rect 13212 35094 13246 35128
rect 13212 35026 13246 35060
rect 13212 34958 13246 34992
rect 13212 34890 13246 34924
rect 13212 34822 13246 34856
rect 13212 34754 13246 34788
rect 13212 34686 13246 34720
rect 13212 34618 13246 34652
rect 13212 34550 13246 34584
rect 13212 34482 13246 34516
rect 13212 34414 13246 34448
rect 13212 34346 13246 34380
rect 13212 34278 13246 34312
rect 13212 34210 13246 34244
rect 13212 34142 13246 34176
rect 13212 34074 13246 34108
rect 13212 34006 13246 34040
rect 13212 33938 13246 33972
rect 13212 33870 13246 33904
rect 13212 33802 13246 33836
rect 13212 33734 13246 33768
rect 13212 33666 13246 33700
rect 13212 33598 13246 33632
rect 13212 33530 13246 33564
rect 13212 33462 13246 33496
rect 13212 33394 13246 33428
rect 13212 33326 13246 33360
rect 13212 33258 13246 33292
rect 13212 33190 13246 33224
rect 13212 33122 13246 33156
rect 13212 33054 13246 33088
rect 13212 32986 13246 33020
rect 13212 32918 13246 32952
rect 13212 32850 13246 32884
rect 13212 32782 13246 32816
rect 13212 32714 13246 32748
rect 13212 32646 13246 32680
rect 13212 32578 13246 32612
rect 13212 32510 13246 32544
rect 13212 32442 13246 32476
rect 13212 32374 13246 32408
rect 13212 32306 13246 32340
rect 13212 32238 13246 32272
rect 13212 32170 13246 32204
rect 13212 32102 13246 32136
rect 13212 32034 13246 32068
rect 13212 31966 13246 32000
rect 13212 31898 13246 31932
rect 13212 31830 13246 31864
rect 13212 31762 13246 31796
rect 13212 31694 13246 31728
rect 13212 31626 13246 31660
rect 13212 31558 13246 31592
rect 13212 31490 13246 31524
rect 13212 31422 13246 31456
rect 13212 31354 13246 31388
rect 13212 31286 13246 31320
rect 13212 31218 13246 31252
rect 13212 31150 13246 31184
rect 13212 31082 13246 31116
rect 13212 31014 13246 31048
rect 13212 30946 13246 30980
rect 13212 30878 13246 30912
rect 13212 30810 13246 30844
rect 13212 30742 13246 30776
rect 13212 30674 13246 30708
rect 13212 30606 13246 30640
rect 13212 30538 13246 30572
rect 13212 30470 13246 30504
rect 13212 30402 13246 30436
rect 13212 30334 13246 30368
rect 13212 30266 13246 30300
rect 13212 30198 13246 30232
rect 13212 30130 13246 30164
rect 13212 30062 13246 30096
rect 13212 29994 13246 30028
rect 13212 29926 13246 29960
rect 13212 29858 13246 29892
rect 13212 29790 13246 29824
rect 13212 29722 13246 29756
rect 13212 29654 13246 29688
rect 13212 29586 13246 29620
rect 13212 29518 13246 29552
rect 13212 29450 13246 29484
rect 13212 29382 13246 29416
rect 13212 29314 13246 29348
rect 13212 29246 13246 29280
rect 13212 29178 13246 29212
rect 13212 29110 13246 29144
rect 13212 29042 13246 29076
rect 13212 28974 13246 29008
rect 13212 28906 13246 28940
rect 13212 28838 13246 28872
rect 13212 28770 13246 28804
rect 13212 28702 13246 28736
rect 13212 28634 13246 28668
rect 13212 28566 13246 28600
rect 13212 28498 13246 28532
rect 13212 28430 13246 28464
rect 13212 28362 13246 28396
rect 13212 28294 13246 28328
rect 13212 28226 13246 28260
rect 13212 28158 13246 28192
rect 13212 28090 13246 28124
rect 13212 28022 13246 28056
rect 13212 27954 13246 27988
rect 13212 27886 13246 27920
rect 13212 27818 13246 27852
rect 13212 27750 13246 27784
rect 13212 27682 13246 27716
rect 13212 27614 13246 27648
rect 13212 27546 13246 27580
rect 13212 27478 13246 27512
rect 13212 27410 13246 27444
rect 13212 27342 13246 27376
rect 13212 27274 13246 27308
rect 13212 27206 13246 27240
rect 13212 27138 13246 27172
rect 13212 27070 13246 27104
rect 13212 27002 13246 27036
rect 13212 26934 13246 26968
rect 13212 26866 13246 26900
rect 13212 26798 13246 26832
rect 13212 26730 13246 26764
rect 13212 26662 13246 26696
rect 13212 26594 13246 26628
rect 13212 26526 13246 26560
rect 13212 26458 13246 26492
rect 13212 26390 13246 26424
rect 13212 26322 13246 26356
rect 13212 26254 13246 26288
rect 13212 26186 13246 26220
rect 13212 26118 13246 26152
rect 13212 26050 13246 26084
rect 13212 25982 13246 26016
rect 13212 25914 13246 25948
rect 13212 25846 13246 25880
rect 13212 25778 13246 25812
rect 13212 25710 13246 25744
rect 13212 25642 13246 25676
rect 13212 25574 13246 25608
rect 13212 25506 13246 25540
rect 13212 25438 13246 25472
rect 13212 25370 13246 25404
rect 13212 25302 13246 25336
rect 13212 25234 13246 25268
rect 13212 25166 13246 25200
rect 13212 25098 13246 25132
rect 13212 25030 13246 25064
rect 13212 24962 13246 24996
rect 13212 24894 13246 24928
rect 13212 24826 13246 24860
rect 13212 24758 13246 24792
rect 13212 24690 13246 24724
rect 13212 24622 13246 24656
rect 13212 24554 13246 24588
rect 13212 24486 13246 24520
rect 13212 24418 13246 24452
rect 13212 24350 13246 24384
rect 13212 24282 13246 24316
rect 13212 24214 13246 24248
rect 13212 24146 13246 24180
rect 13212 24078 13246 24112
rect 13212 24010 13246 24044
rect 13212 23942 13246 23976
rect 13212 23874 13246 23908
rect 13212 23806 13246 23840
rect 13212 23738 13246 23772
rect 13212 23670 13246 23704
rect 13212 23602 13246 23636
rect 13212 23534 13246 23568
rect 13212 23466 13246 23500
rect 13212 23398 13246 23432
rect 13212 23330 13246 23364
rect 13212 23262 13246 23296
rect 13212 23194 13246 23228
rect 13212 23126 13246 23160
rect 13212 23058 13246 23092
rect 13212 22990 13246 23024
rect 13212 22922 13246 22956
rect 13212 22854 13246 22888
rect 13212 22786 13246 22820
rect 13212 22718 13246 22752
rect 13212 22650 13246 22684
rect 13212 22582 13246 22616
rect 13212 22514 13246 22548
rect 13212 22446 13246 22480
rect 13212 22378 13246 22412
rect 13212 22310 13246 22344
rect 13212 22242 13246 22276
rect 13212 22174 13246 22208
rect 13212 22106 13246 22140
rect 13212 22038 13246 22072
rect 13212 21970 13246 22004
rect 13212 21902 13246 21936
rect 13212 21834 13246 21868
rect 13212 21766 13246 21800
rect 13212 21698 13246 21732
rect 13212 21630 13246 21664
rect 13212 21562 13246 21596
rect 13212 21494 13246 21528
rect 13212 21426 13246 21460
rect 13212 21358 13246 21392
rect 13212 21290 13246 21324
rect 13212 21222 13246 21256
rect 13212 21154 13246 21188
rect 13212 21086 13246 21120
rect 13212 21018 13246 21052
rect 13212 20950 13246 20984
rect 13212 20882 13246 20916
rect 13212 20814 13246 20848
rect 13212 20746 13246 20780
rect 13212 20678 13246 20712
rect 13212 20610 13246 20644
rect 13212 20542 13246 20576
rect 13212 20474 13246 20508
rect 13212 20406 13246 20440
rect 13212 20338 13246 20372
rect 13212 20270 13246 20304
rect 13212 20202 13246 20236
rect 13212 20134 13246 20168
rect 13212 20066 13246 20100
rect 13212 19998 13246 20032
rect 13212 19930 13246 19964
rect 13212 19862 13246 19896
rect 13212 19794 13246 19828
rect 13212 19726 13246 19760
rect 13212 19658 13246 19692
rect 13212 19590 13246 19624
rect 13212 19522 13246 19556
rect 13212 19454 13246 19488
rect 13212 19386 13246 19420
rect 13212 19318 13246 19352
rect 13212 19250 13246 19284
rect 13212 19182 13246 19216
rect 13212 19114 13246 19148
rect 13212 19046 13246 19080
rect 13212 18978 13246 19012
rect 13212 18910 13246 18944
rect 13212 18842 13246 18876
rect 13212 18774 13246 18808
rect 13212 18706 13246 18740
rect 13212 18638 13246 18672
rect 13212 18570 13246 18604
rect 13212 18502 13246 18536
rect 13212 18434 13246 18468
rect 13212 18366 13246 18400
rect 13212 18298 13246 18332
rect 13212 18230 13246 18264
rect 13212 18162 13246 18196
rect 13212 18094 13246 18128
rect 13212 18026 13246 18060
rect 13212 17958 13246 17992
rect 13212 17890 13246 17924
rect 13212 17822 13246 17856
rect 13212 17754 13246 17788
rect 13212 17686 13246 17720
rect 13212 17618 13246 17652
rect 13212 17550 13246 17584
rect 13212 17482 13246 17516
rect 13212 17414 13246 17448
rect 13212 17346 13246 17380
rect 13212 17278 13246 17312
rect 13212 17210 13246 17244
rect 13212 17142 13246 17176
rect 13212 17074 13246 17108
rect 13212 17006 13246 17040
rect 13212 16938 13246 16972
rect 13212 16870 13246 16904
rect 13212 16802 13246 16836
rect 13212 16734 13246 16768
rect 13212 16666 13246 16700
rect 13212 16598 13246 16632
rect 13212 16530 13246 16564
rect 13212 16462 13246 16496
rect 13212 16394 13246 16428
rect 13212 16326 13246 16360
rect 13212 16258 13246 16292
rect 13212 16190 13246 16224
rect 13212 16122 13246 16156
rect 13212 16054 13246 16088
rect 13212 15986 13246 16020
rect 13212 15918 13246 15952
rect 13212 15850 13246 15884
rect 13212 15782 13246 15816
rect 13212 15714 13246 15748
rect 13212 15646 13246 15680
rect 13212 15578 13246 15612
rect 13212 15510 13246 15544
rect 13212 15442 13246 15476
rect 13212 15374 13246 15408
rect 13212 15306 13246 15340
rect 13212 15238 13246 15272
rect 13212 15170 13246 15204
rect 13212 15102 13246 15136
rect 13212 15034 13246 15068
rect 13212 14966 13246 15000
rect 13212 14898 13246 14932
rect 13212 14830 13246 14864
rect 13212 14762 13246 14796
rect 13212 14694 13246 14728
rect 13212 14626 13246 14660
rect 13212 14558 13246 14592
rect 13212 14490 13246 14524
rect 13212 14422 13246 14456
rect 13212 14354 13246 14388
rect 13212 14286 13246 14320
rect 13212 14218 13246 14252
rect 13212 14150 13246 14184
rect 13212 14082 13246 14116
rect 13212 14014 13246 14048
rect 13212 13946 13246 13980
rect 13212 13878 13246 13912
rect 13212 13810 13246 13844
rect 13212 13742 13246 13776
rect 13212 13674 13246 13708
rect 13212 13606 13246 13640
rect 13212 13538 13246 13572
rect 13212 13470 13246 13504
rect 13212 13402 13246 13436
rect 13212 13334 13246 13368
rect 13212 13266 13246 13300
rect 13212 13198 13246 13232
rect 13212 13130 13246 13164
rect 13212 13062 13246 13096
rect 13212 12994 13246 13028
rect 13212 12926 13246 12960
rect 13212 12858 13246 12892
rect 13212 12790 13246 12824
rect 13212 12722 13246 12756
rect 13212 12654 13246 12688
rect 13212 12586 13246 12620
rect 13212 12518 13246 12552
rect 13212 12450 13246 12484
rect 13212 12382 13246 12416
rect 13212 12314 13246 12348
rect 13212 12246 13246 12280
rect 13212 12178 13246 12212
rect 13212 12110 13246 12144
rect 13212 12042 13246 12076
rect 13212 11974 13246 12008
rect 13212 11906 13246 11940
rect 13212 11838 13246 11872
rect 13212 11770 13246 11804
rect 13212 11702 13246 11736
rect 13212 11634 13246 11668
rect 13212 11566 13246 11600
rect 13212 11498 13246 11532
rect 13212 11430 13246 11464
rect 13212 11362 13246 11396
rect 13212 11294 13246 11328
rect 13212 11226 13246 11260
rect 13212 11158 13246 11192
rect 13212 11090 13246 11124
rect 13212 11022 13246 11056
rect 13212 10954 13246 10988
rect 13212 10886 13246 10920
rect 13212 10818 13246 10852
rect 13212 10750 13246 10784
rect 13212 10682 13246 10716
rect 13212 10614 13246 10648
rect 13212 10546 13246 10580
rect 13212 10478 13246 10512
rect 13212 10410 13246 10444
rect 13212 10342 13246 10376
rect 13212 10274 13246 10308
rect 13212 10206 13246 10240
rect 13212 10138 13246 10172
rect 13212 10070 13246 10104
rect 13212 10002 13246 10036
rect 13212 9934 13246 9968
rect 13212 9866 13246 9900
rect 13212 9798 13246 9832
rect 13212 9730 13246 9764
rect 13212 9662 13246 9696
rect 13212 9594 13246 9628
rect 13212 9526 13246 9560
rect 13212 9458 13246 9492
rect 13212 9390 13246 9424
rect 13212 9322 13246 9356
rect 13212 9254 13246 9288
rect 13212 9186 13246 9220
rect 13212 9118 13246 9152
rect 13212 9050 13246 9084
rect 13212 8982 13246 9016
rect 13212 8914 13246 8948
rect 13212 8846 13246 8880
rect 13212 8778 13246 8812
rect 13212 8710 13246 8744
rect 13212 8642 13246 8676
rect 13212 8574 13246 8608
rect 13212 8506 13246 8540
rect 13212 8438 13246 8472
rect 13212 8370 13246 8404
rect 13212 8302 13246 8336
rect 13212 8234 13246 8268
rect 13212 8166 13246 8200
rect 13212 8098 13246 8132
rect 13212 8030 13246 8064
rect 13212 7962 13246 7996
rect 13212 7894 13246 7928
rect 13212 7826 13246 7860
rect 13212 7758 13246 7792
rect 13212 7690 13246 7724
rect 13212 7622 13246 7656
rect 13212 7554 13246 7588
rect 13212 7486 13246 7520
rect 13212 7418 13246 7452
rect 13212 7350 13246 7384
rect 13212 7282 13246 7316
rect 13212 7214 13246 7248
rect 13212 7146 13246 7180
rect 13212 7078 13246 7112
rect 13212 7010 13246 7044
rect 13212 6942 13246 6976
rect 13212 6874 13246 6908
rect 13212 6806 13246 6840
rect 13212 6738 13246 6772
rect 13212 6670 13246 6704
rect 13212 6602 13246 6636
rect 13212 6534 13246 6568
rect 13212 6466 13246 6500
rect 13212 6398 13246 6432
rect 13212 6330 13246 6364
rect 13212 6262 13246 6296
rect 13212 6194 13246 6228
rect 13212 6126 13246 6160
rect 13212 6058 13246 6092
rect 13212 5990 13246 6024
rect 13212 5922 13246 5956
rect 13212 5854 13246 5888
rect 13212 5786 13246 5820
rect 13212 5718 13246 5752
rect 13212 5650 13246 5684
rect 13212 5582 13246 5616
rect 13212 5514 13246 5548
rect 13212 5446 13246 5480
rect 13212 5378 13246 5412
rect 13212 5310 13246 5344
rect 13212 5242 13246 5276
rect 13212 5174 13246 5208
rect 13212 5106 13246 5140
rect 13212 5038 13246 5072
rect 13212 4970 13246 5004
rect 13212 4902 13246 4936
rect 13212 4834 13246 4868
rect 13212 4766 13246 4800
rect 13212 4698 13246 4732
rect 13212 4630 13246 4664
rect 13212 4562 13246 4596
rect 13212 4494 13246 4528
rect 13212 4426 13246 4460
rect 13212 4358 13246 4392
rect 13212 4290 13246 4324
rect 13212 4222 13246 4256
rect 13212 4154 13246 4188
rect 13212 4086 13246 4120
rect 13212 4018 13246 4052
rect 13212 3950 13246 3984
rect 13212 3882 13246 3916
rect 13212 3814 13246 3848
rect 13212 3746 13246 3780
rect 13212 3678 13246 3712
rect 13212 3610 13246 3644
rect 13212 3542 13246 3576
rect 13212 3474 13246 3508
rect 13212 3406 13246 3440
rect 13212 3338 13246 3372
rect 13212 3270 13246 3304
rect 13212 3202 13246 3236
rect 13212 3134 13246 3168
rect 13212 3066 13246 3100
rect 13212 2998 13246 3032
rect 13212 2930 13246 2964
rect 13212 2862 13246 2896
rect 13212 2794 13246 2828
rect 13212 2726 13246 2760
rect 13212 2658 13246 2692
rect 13212 2590 13246 2624
rect 13212 2522 13246 2556
rect 13212 2454 13246 2488
rect 13212 2386 13246 2420
rect 13212 2318 13246 2352
rect 13212 2250 13246 2284
rect 13212 2182 13246 2216
rect 13212 2114 13246 2148
rect 13212 2046 13246 2080
rect 13212 1978 13246 2012
rect 13212 1910 13246 1944
rect 13212 1842 13246 1876
rect 13212 1774 13246 1808
rect 13212 1706 13246 1740
rect 13212 1638 13246 1672
rect 13212 1570 13246 1604
rect 13212 1502 13246 1536
rect 13212 1434 13246 1468
rect 13212 1366 13246 1400
rect 13212 1298 13246 1332
rect 13212 1230 13246 1264
rect 13212 1162 13246 1196
rect 13212 1094 13246 1128
rect 13212 1026 13246 1060
rect 13212 958 13246 992
rect 13212 890 13246 924
rect 13212 822 13246 856
rect 13212 754 13246 788
rect 13212 686 13246 720
rect 13212 618 13246 652
rect 13212 550 13246 584
rect 13212 482 13246 516
rect 13212 414 13246 448
rect 11424 349 11458 383
rect 11424 281 11458 315
rect 14940 38485 14974 38519
rect 14940 38417 14974 38451
rect 14940 38349 14974 38383
rect 14940 38281 14974 38315
rect 14940 38213 14974 38247
rect 14940 38145 14974 38179
rect 14940 38077 14974 38111
rect 14940 38009 14974 38043
rect 14940 37941 14974 37975
rect 14940 37873 14974 37907
rect 14940 37805 14974 37839
rect 14940 37737 14974 37771
rect 14940 37669 14974 37703
rect 14940 37601 14974 37635
rect 14940 37533 14974 37567
rect 14940 37465 14974 37499
rect 14940 37397 14974 37431
rect 14940 37329 14974 37363
rect 14940 37261 14974 37295
rect 14940 37193 14974 37227
rect 14940 37125 14974 37159
rect 14940 37057 14974 37091
rect 14940 36989 14974 37023
rect 14940 36921 14974 36955
rect 14940 36853 14974 36887
rect 14940 36785 14974 36819
rect 14940 36717 14974 36751
rect 14940 36649 14974 36683
rect 14940 36581 14974 36615
rect 14940 36513 14974 36547
rect 14940 36445 14974 36479
rect 14940 36377 14974 36411
rect 14940 36309 14974 36343
rect 14940 36241 14974 36275
rect 14940 36173 14974 36207
rect 14940 36105 14974 36139
rect 14940 36037 14974 36071
rect 14940 35969 14974 36003
rect 14940 35901 14974 35935
rect 14940 35833 14974 35867
rect 14940 35765 14974 35799
rect 14940 35697 14974 35731
rect 14940 35629 14974 35663
rect 14940 35561 14974 35595
rect 14940 35493 14974 35527
rect 14940 35425 14974 35459
rect 14940 35357 14974 35391
rect 14940 35289 14974 35323
rect 14940 35221 14974 35255
rect 14940 35153 14974 35187
rect 14940 35085 14974 35119
rect 14940 35017 14974 35051
rect 14940 34949 14974 34983
rect 14940 34881 14974 34915
rect 14940 34813 14974 34847
rect 14940 34745 14974 34779
rect 14940 34677 14974 34711
rect 14940 34609 14974 34643
rect 14940 34541 14974 34575
rect 14940 34473 14974 34507
rect 14940 34405 14974 34439
rect 14940 34337 14974 34371
rect 14940 34269 14974 34303
rect 14940 34201 14974 34235
rect 14940 34133 14974 34167
rect 14940 34065 14974 34099
rect 14940 33997 14974 34031
rect 14940 33929 14974 33963
rect 14940 33861 14974 33895
rect 14940 33793 14974 33827
rect 14940 33725 14974 33759
rect 14940 33657 14974 33691
rect 14940 33589 14974 33623
rect 14940 33521 14974 33555
rect 14940 33453 14974 33487
rect 14940 33385 14974 33419
rect 14940 33317 14974 33351
rect 14940 33249 14974 33283
rect 14940 33181 14974 33215
rect 14940 33113 14974 33147
rect 14940 33045 14974 33079
rect 14940 32977 14974 33011
rect 14940 32909 14974 32943
rect 14940 32841 14974 32875
rect 14940 32773 14974 32807
rect 14940 32705 14974 32739
rect 14940 32637 14974 32671
rect 14940 32569 14974 32603
rect 14940 32501 14974 32535
rect 14940 32433 14974 32467
rect 14940 32365 14974 32399
rect 14940 32297 14974 32331
rect 14940 32229 14974 32263
rect 14940 32161 14974 32195
rect 14940 32093 14974 32127
rect 14940 32025 14974 32059
rect 14940 31957 14974 31991
rect 14940 31889 14974 31923
rect 14940 31821 14974 31855
rect 14940 31753 14974 31787
rect 14940 31685 14974 31719
rect 14940 31617 14974 31651
rect 14940 31549 14974 31583
rect 14940 31481 14974 31515
rect 14940 31413 14974 31447
rect 14940 31345 14974 31379
rect 14940 31277 14974 31311
rect 14940 31209 14974 31243
rect 14940 31141 14974 31175
rect 14940 31073 14974 31107
rect 14940 31005 14974 31039
rect 14940 30937 14974 30971
rect 14940 30869 14974 30903
rect 14940 30801 14974 30835
rect 14940 30733 14974 30767
rect 14940 30665 14974 30699
rect 14940 30597 14974 30631
rect 14940 30529 14974 30563
rect 14940 30461 14974 30495
rect 14940 30393 14974 30427
rect 14940 30325 14974 30359
rect 14940 30257 14974 30291
rect 14940 30189 14974 30223
rect 14940 30121 14974 30155
rect 14940 30053 14974 30087
rect 14940 29985 14974 30019
rect 14940 29917 14974 29951
rect 14940 29849 14974 29883
rect 14940 29781 14974 29815
rect 14940 29713 14974 29747
rect 14940 29645 14974 29679
rect 14940 29577 14974 29611
rect 14940 29509 14974 29543
rect 14940 29441 14974 29475
rect 14940 29373 14974 29407
rect 14940 29305 14974 29339
rect 14940 29237 14974 29271
rect 14940 29169 14974 29203
rect 14940 29101 14974 29135
rect 14940 29033 14974 29067
rect 14940 28965 14974 28999
rect 14940 28897 14974 28931
rect 14940 28829 14974 28863
rect 14940 28761 14974 28795
rect 14940 28693 14974 28727
rect 14940 28625 14974 28659
rect 14940 28557 14974 28591
rect 14940 28489 14974 28523
rect 14940 28421 14974 28455
rect 14940 28353 14974 28387
rect 14940 28285 14974 28319
rect 14940 28217 14974 28251
rect 14940 28149 14974 28183
rect 14940 28081 14974 28115
rect 14940 28013 14974 28047
rect 14940 27945 14974 27979
rect 14940 27877 14974 27911
rect 14940 27809 14974 27843
rect 14940 27741 14974 27775
rect 14940 27673 14974 27707
rect 14940 27605 14974 27639
rect 14940 27537 14974 27571
rect 14940 27469 14974 27503
rect 14940 27401 14974 27435
rect 14940 27333 14974 27367
rect 14940 27265 14974 27299
rect 14940 27197 14974 27231
rect 14940 27129 14974 27163
rect 14940 27061 14974 27095
rect 14940 26993 14974 27027
rect 14940 26925 14974 26959
rect 14940 26857 14974 26891
rect 14940 26789 14974 26823
rect 14940 26721 14974 26755
rect 14940 26653 14974 26687
rect 14940 26585 14974 26619
rect 14940 26517 14974 26551
rect 14940 26449 14974 26483
rect 14940 26381 14974 26415
rect 14940 26313 14974 26347
rect 14940 26245 14974 26279
rect 14940 26177 14974 26211
rect 14940 26109 14974 26143
rect 14940 26041 14974 26075
rect 14940 25973 14974 26007
rect 14940 25905 14974 25939
rect 14940 25837 14974 25871
rect 14940 25769 14974 25803
rect 14940 25701 14974 25735
rect 14940 25633 14974 25667
rect 14940 25565 14974 25599
rect 14940 25497 14974 25531
rect 14940 25429 14974 25463
rect 14940 25361 14974 25395
rect 14940 25293 14974 25327
rect 14940 25225 14974 25259
rect 14940 25157 14974 25191
rect 14940 25089 14974 25123
rect 14940 25021 14974 25055
rect 14940 24953 14974 24987
rect 14940 24885 14974 24919
rect 14940 24817 14974 24851
rect 14940 24749 14974 24783
rect 14940 24681 14974 24715
rect 14940 24613 14974 24647
rect 14940 24545 14974 24579
rect 14940 24477 14974 24511
rect 14940 24409 14974 24443
rect 14940 24341 14974 24375
rect 14940 24273 14974 24307
rect 14940 24205 14974 24239
rect 14940 24137 14974 24171
rect 14940 24069 14974 24103
rect 14940 24001 14974 24035
rect 14940 23933 14974 23967
rect 14940 23865 14974 23899
rect 14940 23797 14974 23831
rect 14940 23729 14974 23763
rect 14940 23661 14974 23695
rect 14940 23593 14974 23627
rect 14940 23525 14974 23559
rect 14940 23457 14974 23491
rect 14940 23389 14974 23423
rect 14940 23321 14974 23355
rect 14940 23253 14974 23287
rect 14940 23185 14974 23219
rect 14940 23117 14974 23151
rect 14940 23049 14974 23083
rect 14940 22981 14974 23015
rect 14940 22913 14974 22947
rect 14940 22845 14974 22879
rect 14940 22777 14974 22811
rect 14940 22709 14974 22743
rect 14940 22641 14974 22675
rect 14940 22573 14974 22607
rect 14940 22505 14974 22539
rect 14940 22437 14974 22471
rect 14940 22369 14974 22403
rect 14940 22301 14974 22335
rect 14940 22233 14974 22267
rect 14940 22165 14974 22199
rect 14940 22097 14974 22131
rect 14940 22029 14974 22063
rect 14940 21961 14974 21995
rect 14940 21893 14974 21927
rect 14940 21825 14974 21859
rect 14940 21757 14974 21791
rect 14940 21689 14974 21723
rect 14940 21621 14974 21655
rect 14940 21553 14974 21587
rect 14940 21485 14974 21519
rect 14940 21417 14974 21451
rect 14940 21349 14974 21383
rect 14940 21281 14974 21315
rect 14940 21213 14974 21247
rect 14940 21145 14974 21179
rect 14940 21077 14974 21111
rect 14940 21009 14974 21043
rect 14940 20941 14974 20975
rect 14940 20873 14974 20907
rect 14940 20805 14974 20839
rect 14940 20737 14974 20771
rect 14940 20669 14974 20703
rect 14940 20601 14974 20635
rect 14940 20533 14974 20567
rect 14940 20465 14974 20499
rect 14940 20397 14974 20431
rect 14940 20329 14974 20363
rect 14940 20261 14974 20295
rect 14940 20193 14974 20227
rect 14940 20125 14974 20159
rect 14940 20057 14974 20091
rect 14940 19989 14974 20023
rect 14940 19921 14974 19955
rect 14940 19853 14974 19887
rect 14940 19785 14974 19819
rect 14940 19717 14974 19751
rect 14940 19649 14974 19683
rect 14940 19581 14974 19615
rect 14940 19513 14974 19547
rect 14940 19445 14974 19479
rect 14940 19377 14974 19411
rect 14940 19309 14974 19343
rect 14940 19241 14974 19275
rect 14940 19173 14974 19207
rect 14940 19105 14974 19139
rect 14940 19037 14974 19071
rect 14940 18969 14974 19003
rect 14940 18901 14974 18935
rect 14940 18833 14974 18867
rect 14940 18765 14974 18799
rect 14940 18697 14974 18731
rect 14940 18629 14974 18663
rect 14940 18561 14974 18595
rect 14940 18493 14974 18527
rect 14940 18425 14974 18459
rect 14940 18357 14974 18391
rect 14940 18289 14974 18323
rect 14940 18221 14974 18255
rect 14940 18153 14974 18187
rect 14940 18085 14974 18119
rect 14940 18017 14974 18051
rect 14940 17949 14974 17983
rect 14940 17881 14974 17915
rect 14940 17813 14974 17847
rect 14940 17745 14974 17779
rect 14940 17677 14974 17711
rect 14940 17609 14974 17643
rect 14940 17541 14974 17575
rect 14940 17473 14974 17507
rect 14940 17405 14974 17439
rect 14940 17337 14974 17371
rect 14940 17269 14974 17303
rect 14940 17201 14974 17235
rect 14940 17133 14974 17167
rect 14940 17065 14974 17099
rect 14940 16997 14974 17031
rect 14940 16929 14974 16963
rect 14940 16861 14974 16895
rect 14940 16793 14974 16827
rect 14940 16725 14974 16759
rect 14940 16657 14974 16691
rect 14940 16589 14974 16623
rect 14940 16521 14974 16555
rect 14940 16453 14974 16487
rect 14940 16385 14974 16419
rect 14940 16317 14974 16351
rect 14940 16249 14974 16283
rect 14940 16181 14974 16215
rect 14940 16113 14974 16147
rect 14940 16045 14974 16079
rect 14940 15977 14974 16011
rect 14940 15909 14974 15943
rect 14940 15841 14974 15875
rect 14940 15773 14974 15807
rect 14940 15705 14974 15739
rect 14940 15637 14974 15671
rect 14940 15569 14974 15603
rect 14940 15501 14974 15535
rect 14940 15433 14974 15467
rect 14940 15365 14974 15399
rect 14940 15297 14974 15331
rect 14940 15229 14974 15263
rect 14940 15161 14974 15195
rect 14940 15093 14974 15127
rect 14940 15025 14974 15059
rect 14940 14957 14974 14991
rect 14940 14889 14974 14923
rect 14940 14821 14974 14855
rect 14940 14753 14974 14787
rect 14940 14685 14974 14719
rect 14940 14617 14974 14651
rect 14940 14549 14974 14583
rect 14940 14481 14974 14515
rect 14940 14413 14974 14447
rect 14940 14345 14974 14379
rect 14940 14277 14974 14311
rect 14940 14209 14974 14243
rect 14940 14141 14974 14175
rect 14940 14073 14974 14107
rect 14940 14005 14974 14039
rect 14940 13937 14974 13971
rect 14940 13869 14974 13903
rect 14940 13801 14974 13835
rect 14940 13733 14974 13767
rect 14940 13665 14974 13699
rect 14940 13597 14974 13631
rect 14940 13529 14974 13563
rect 14940 13461 14974 13495
rect 14940 13393 14974 13427
rect 14940 13325 14974 13359
rect 14940 13257 14974 13291
rect 14940 13189 14974 13223
rect 14940 13121 14974 13155
rect 14940 13053 14974 13087
rect 14940 12985 14974 13019
rect 14940 12917 14974 12951
rect 14940 12849 14974 12883
rect 14940 12781 14974 12815
rect 14940 12713 14974 12747
rect 14940 12645 14974 12679
rect 14940 12577 14974 12611
rect 14940 12509 14974 12543
rect 14940 12441 14974 12475
rect 14940 12373 14974 12407
rect 14940 12305 14974 12339
rect 14940 12237 14974 12271
rect 14940 12169 14974 12203
rect 14940 12101 14974 12135
rect 14940 12033 14974 12067
rect 14940 11965 14974 11999
rect 14940 11897 14974 11931
rect 14940 11829 14974 11863
rect 14940 11761 14974 11795
rect 14940 11693 14974 11727
rect 14940 11625 14974 11659
rect 14940 11557 14974 11591
rect 14940 11489 14974 11523
rect 14940 11421 14974 11455
rect 14940 11353 14974 11387
rect 14940 11285 14974 11319
rect 14940 11217 14974 11251
rect 14940 11149 14974 11183
rect 14940 11081 14974 11115
rect 14940 11013 14974 11047
rect 14940 10945 14974 10979
rect 14940 10877 14974 10911
rect 14940 10809 14974 10843
rect 14940 10741 14974 10775
rect 14940 10673 14974 10707
rect 14940 10605 14974 10639
rect 14940 10537 14974 10571
rect 14940 10469 14974 10503
rect 14940 10401 14974 10435
rect 14940 10333 14974 10367
rect 14940 10265 14974 10299
rect 14940 10197 14974 10231
rect 14940 10129 14974 10163
rect 14940 10061 14974 10095
rect 14940 9993 14974 10027
rect 14940 9925 14974 9959
rect 14940 9857 14974 9891
rect 14940 9789 14974 9823
rect 14940 9721 14974 9755
rect 14940 9653 14974 9687
rect 14940 9585 14974 9619
rect 14940 9517 14974 9551
rect 14940 9449 14974 9483
rect 14940 9381 14974 9415
rect 14940 9313 14974 9347
rect 14940 9245 14974 9279
rect 14940 9177 14974 9211
rect 14940 9109 14974 9143
rect 14940 9041 14974 9075
rect 14940 8973 14974 9007
rect 14940 8905 14974 8939
rect 14940 8837 14974 8871
rect 14940 8769 14974 8803
rect 14940 8701 14974 8735
rect 14940 8633 14974 8667
rect 14940 8565 14974 8599
rect 14940 8497 14974 8531
rect 14940 8429 14974 8463
rect 14940 8361 14974 8395
rect 14940 8293 14974 8327
rect 14940 8225 14974 8259
rect 14940 8157 14974 8191
rect 14940 8089 14974 8123
rect 14940 8021 14974 8055
rect 14940 7953 14974 7987
rect 14940 7885 14974 7919
rect 14940 7817 14974 7851
rect 14940 7749 14974 7783
rect 14940 7681 14974 7715
rect 14940 7613 14974 7647
rect 14940 7545 14974 7579
rect 14940 7477 14974 7511
rect 14940 7409 14974 7443
rect 14940 7341 14974 7375
rect 14940 7273 14974 7307
rect 14940 7205 14974 7239
rect 14940 7137 14974 7171
rect 14940 7069 14974 7103
rect 14940 7001 14974 7035
rect 14940 6933 14974 6967
rect 14940 6865 14974 6899
rect 14940 6797 14974 6831
rect 14940 6729 14974 6763
rect 14940 6661 14974 6695
rect 14940 6593 14974 6627
rect 14940 6525 14974 6559
rect 14940 6457 14974 6491
rect 14940 6389 14974 6423
rect 14940 6321 14974 6355
rect 14940 6253 14974 6287
rect 14940 6185 14974 6219
rect 14940 6117 14974 6151
rect 14940 6049 14974 6083
rect 14940 5981 14974 6015
rect 14940 5913 14974 5947
rect 14940 5845 14974 5879
rect 14940 5777 14974 5811
rect 14940 5709 14974 5743
rect 14940 5641 14974 5675
rect 14940 5573 14974 5607
rect 14940 5505 14974 5539
rect 14940 5437 14974 5471
rect 14940 5369 14974 5403
rect 14940 5301 14974 5335
rect 14940 5233 14974 5267
rect 14940 5165 14974 5199
rect 14940 5097 14974 5131
rect 14940 5029 14974 5063
rect 14940 4961 14974 4995
rect 14940 4893 14974 4927
rect 14940 4825 14974 4859
rect 14940 4757 14974 4791
rect 14940 4689 14974 4723
rect 14940 4621 14974 4655
rect 14940 4553 14974 4587
rect 14940 4485 14974 4519
rect 14940 4417 14974 4451
rect 14940 4349 14974 4383
rect 14940 4281 14974 4315
rect 14940 4213 14974 4247
rect 14940 4145 14974 4179
rect 14940 4077 14974 4111
rect 14940 4009 14974 4043
rect 14940 3941 14974 3975
rect 14940 3873 14974 3907
rect 14940 3805 14974 3839
rect 14940 3737 14974 3771
rect 14940 3669 14974 3703
rect 14940 3601 14974 3635
rect 14940 3533 14974 3567
rect 14940 3465 14974 3499
rect 14940 3397 14974 3431
rect 14940 3329 14974 3363
rect 14940 3205 14974 3295
rect 14940 3137 14974 3171
rect 14940 3069 14974 3103
rect 14940 3001 14974 3035
rect 14940 2933 14974 2967
rect 14940 2865 14974 2899
rect 14940 2797 14974 2831
rect 14940 2729 14974 2763
rect 14940 2661 14974 2695
rect 14940 2593 14974 2627
rect 14940 2525 14974 2559
rect 14940 2457 14974 2491
rect 14940 2389 14974 2423
rect 14940 2321 14974 2355
rect 14940 2253 14974 2287
rect 14940 2185 14974 2219
rect 14940 2117 14974 2151
rect 14940 2049 14974 2083
rect 14940 1981 14974 2015
rect 14940 1913 14974 1947
rect 14940 1845 14974 1879
rect 14940 1777 14974 1811
rect 14940 1709 14974 1743
rect 14940 1641 14974 1675
rect 14940 1573 14974 1607
rect 14940 1505 14974 1539
rect 14940 1437 14974 1471
rect 14940 1369 14974 1403
rect 14940 1301 14974 1335
rect 14940 1233 14974 1267
rect 14940 1165 14974 1199
rect 14940 1097 14974 1131
rect 14940 1029 14974 1063
rect 14940 961 14974 995
rect 14940 893 14974 927
rect 14940 825 14974 859
rect 14940 757 14974 791
rect 14940 689 14974 723
rect 14940 621 14974 655
rect 14940 553 14974 587
rect 14940 485 14974 519
rect 14940 417 14974 451
rect 13212 346 13246 380
rect 13212 278 13246 312
rect 11424 213 11458 247
rect 11424 145 11458 179
rect 11424 74 11458 111
rect 14940 349 14974 383
rect 14940 281 14974 315
rect 13212 210 13246 244
rect 13212 142 13246 176
rect 13212 74 13246 108
rect 14940 213 14974 247
rect 14940 145 14974 179
rect 14940 74 14974 111
rect 11424 40 11492 74
rect 11526 40 11560 74
rect 11594 40 11628 74
rect 11662 40 11696 74
rect 11730 40 11764 74
rect 11798 40 11832 74
rect 11866 40 11900 74
rect 11934 40 11968 74
rect 12002 40 12036 74
rect 12070 40 12104 74
rect 12138 40 12172 74
rect 12206 40 12240 74
rect 12274 40 12308 74
rect 12342 40 12376 74
rect 12410 40 12444 74
rect 12478 40 12512 74
rect 12546 40 12580 74
rect 12614 40 12648 74
rect 12682 40 12716 74
rect 12750 40 12784 74
rect 12818 40 12852 74
rect 12886 40 12920 74
rect 12954 40 12988 74
rect 13022 40 13056 74
rect 13090 40 13124 74
rect 13158 40 13308 74
rect 13342 40 13376 74
rect 13410 40 13444 74
rect 13478 40 13512 74
rect 13546 40 13580 74
rect 13614 40 13648 74
rect 13682 40 13716 74
rect 13750 40 13784 74
rect 13818 40 13852 74
rect 13886 40 13920 74
rect 13954 40 13988 74
rect 14022 40 14056 74
rect 14090 40 14124 74
rect 14158 40 14192 74
rect 14226 40 14260 74
rect 14294 40 14328 74
rect 14362 40 14396 74
rect 14430 40 14464 74
rect 14498 40 14532 74
rect 14566 40 14600 74
rect 14634 40 14668 74
rect 14702 40 14736 74
rect 14770 40 14804 74
rect 14838 40 14872 74
rect 14906 40 14974 74
rect 11607 -189 11631 -155
rect 11665 -189 11699 -155
rect 11733 -189 11767 -155
rect 11801 -189 11835 -155
rect 11869 -189 11903 -155
rect 11937 -189 11971 -155
rect 12005 -189 12039 -155
rect 12073 -189 12107 -155
rect 12141 -189 12175 -155
rect 12209 -189 12243 -155
rect 12277 -189 12311 -155
rect 12345 -189 12379 -155
rect 12413 -189 12447 -155
rect 12481 -189 12515 -155
rect 12549 -189 12583 -155
rect 12617 -189 12651 -155
rect 12685 -189 12719 -155
rect 12753 -189 12787 -155
rect 12821 -189 12856 -155
rect 12890 -189 12925 -155
rect 12959 -189 12994 -155
rect 13028 -189 13063 -155
rect 13097 -189 13132 -155
rect 13166 -189 13201 -155
rect 13235 -189 13270 -155
rect 13304 -189 13339 -155
rect 13373 -189 13408 -155
rect 13442 -189 13477 -155
rect 13511 -189 13546 -155
rect 13580 -189 13615 -155
rect 13649 -189 13684 -155
rect 13718 -189 13753 -155
rect 13787 -189 13822 -155
rect 13856 -189 13891 -155
rect 13925 -189 13960 -155
rect 13994 -189 14029 -155
rect 14063 -189 14098 -155
rect 14132 -189 14167 -155
rect 14201 -189 14236 -155
rect 14270 -189 14305 -155
rect 14339 -189 14374 -155
rect 14408 -189 14443 -155
rect 14477 -189 14512 -155
rect 14546 -189 14581 -155
rect 14615 -189 14650 -155
rect 14684 -189 14719 -155
rect 14753 -189 14777 -155
<< mvnsubdiff >>
rect 5940 2568 5974 2602
rect 5940 2500 5974 2534
rect 5940 2432 5974 2466
rect 5940 2364 5974 2398
rect 5940 2296 5974 2330
rect 5940 2228 5974 2262
rect 5940 2160 5974 2194
rect 5940 2092 5974 2126
rect 5940 2024 5974 2058
rect 5940 1956 5974 1990
rect 5940 1888 5974 1922
rect 5940 1820 5974 1854
rect 5940 1752 5974 1786
rect 5940 1684 5974 1718
rect 5940 1616 5974 1650
rect 5940 1548 5974 1582
rect 5940 1480 5974 1514
rect 5940 1412 5974 1446
rect 5940 1344 5974 1378
rect 5940 1276 5974 1310
rect 5940 1208 5974 1242
rect 5940 1140 5974 1174
rect 5940 1072 5974 1106
rect 5940 994 5974 1038
<< mvpsubdiffcont >>
rect -142 38723 -108 38757
rect -74 38723 -40 38757
rect -6 38723 28 38757
rect 62 38723 96 38757
rect 130 38723 164 38757
rect 198 38723 232 38757
rect 266 38723 300 38757
rect 334 38723 368 38757
rect 402 38723 436 38757
rect 470 38723 504 38757
rect 538 38723 572 38757
rect 606 38723 640 38757
rect 674 38723 708 38757
rect 742 38723 776 38757
rect 810 38723 844 38757
rect 878 38723 912 38757
rect 946 38723 980 38757
rect 1014 38723 1048 38757
rect 1082 38723 1116 38757
rect 1150 38723 1184 38757
rect 1218 38723 1252 38757
rect 1286 38723 1320 38757
rect 1354 38723 1388 38757
rect 1422 38723 1456 38757
rect 1490 38723 1524 38757
rect 1558 38723 1592 38757
rect 1626 38723 1660 38757
rect 1694 38723 1728 38757
rect 1762 38723 1796 38757
rect 1898 38723 1932 38757
rect 1966 38723 2000 38757
rect 2034 38723 2068 38757
rect 2102 38723 2136 38757
rect 2170 38723 2204 38757
rect 2238 38723 2272 38757
rect 2306 38723 2340 38757
rect 2374 38723 2408 38757
rect 2442 38723 2476 38757
rect 2510 38723 2544 38757
rect 2578 38723 2612 38757
rect 2646 38723 2680 38757
rect 2714 38723 2748 38757
rect 2782 38723 2816 38757
rect 2850 38723 2884 38757
rect 2918 38723 2952 38757
rect 2986 38723 3020 38757
rect 3054 38723 3088 38757
rect 3122 38723 3156 38757
rect 3190 38723 3224 38757
rect 3258 38723 3292 38757
rect 3326 38723 3360 38757
rect 3394 38723 3428 38757
rect 3462 38723 3496 38757
rect 3530 38723 3564 38757
rect 3598 38723 3632 38757
rect 3666 38723 3700 38757
rect 3734 38723 3768 38757
rect 3802 38723 3836 38757
rect 3870 38723 3904 38757
rect 4074 38723 4108 38757
rect 4142 38723 4176 38757
rect 4210 38723 4244 38757
rect 4278 38723 4312 38757
rect 4346 38723 4380 38757
rect 4414 38723 4448 38757
rect 4482 38723 4516 38757
rect 4550 38723 4584 38757
rect 4618 38723 4652 38757
rect 4686 38723 4720 38757
rect 4754 38723 4788 38757
rect 4822 38723 4856 38757
rect 4890 38723 4924 38757
rect 4958 38723 4992 38757
rect 5026 38723 5060 38757
rect 5094 38723 5128 38757
rect 5162 38723 5196 38757
rect 5230 38723 5264 38757
rect 5298 38723 5332 38757
rect 5366 38723 5400 38757
rect 5434 38723 5468 38757
rect 5502 38723 5536 38757
rect 5570 38723 5604 38757
rect 5638 38723 5672 38757
rect 5706 38723 5740 38757
rect 5774 38723 5808 38757
rect 5842 38723 5876 38757
rect 5910 38723 5944 38757
rect 5978 38723 6012 38757
rect 6046 38723 6080 38757
rect -252 38655 -218 38689
rect -252 38587 -218 38621
rect -252 38519 -218 38553
rect -252 38451 -218 38485
rect -252 38383 -218 38417
rect -252 38315 -218 38349
rect -252 38247 -218 38281
rect -252 38179 -218 38213
rect -252 38111 -218 38145
rect -252 38043 -218 38077
rect -252 37975 -218 38009
rect -252 37907 -218 37941
rect -252 37839 -218 37873
rect -252 37771 -218 37805
rect -252 37703 -218 37737
rect -252 37635 -218 37669
rect -252 37567 -218 37601
rect -252 37499 -218 37533
rect -252 37431 -218 37465
rect -252 37363 -218 37397
rect -252 37295 -218 37329
rect -252 37227 -218 37261
rect -252 37159 -218 37193
rect -252 37091 -218 37125
rect -252 37023 -218 37057
rect -252 36955 -218 36989
rect -252 36887 -218 36921
rect -252 36819 -218 36853
rect -252 36751 -218 36785
rect -252 36683 -218 36717
rect -252 36615 -218 36649
rect -252 36547 -218 36581
rect -252 36479 -218 36513
rect -252 36411 -218 36445
rect -252 36343 -218 36377
rect -252 36275 -218 36309
rect -252 36207 -218 36241
rect -252 36139 -218 36173
rect -252 36071 -218 36105
rect -252 36003 -218 36037
rect -252 35935 -218 35969
rect -252 35867 -218 35901
rect -252 35799 -218 35833
rect -252 35731 -218 35765
rect -252 35663 -218 35697
rect -252 35595 -218 35629
rect -252 35527 -218 35561
rect -252 35459 -218 35493
rect -252 35391 -218 35425
rect -252 35323 -218 35357
rect -252 35255 -218 35289
rect -252 35187 -218 35221
rect -252 35119 -218 35153
rect -252 35051 -218 35085
rect -252 34983 -218 35017
rect -252 34915 -218 34949
rect -252 34847 -218 34881
rect -252 34779 -218 34813
rect -252 34711 -218 34745
rect -252 34643 -218 34677
rect -252 34575 -218 34609
rect -252 34507 -218 34541
rect -252 34439 -218 34473
rect -252 34371 -218 34405
rect -252 34303 -218 34337
rect -252 34235 -218 34269
rect -252 34167 -218 34201
rect -252 34099 -218 34133
rect -252 34031 -218 34065
rect -252 33963 -218 33997
rect -252 33895 -218 33929
rect -252 33827 -218 33861
rect -252 33759 -218 33793
rect -252 33691 -218 33725
rect -252 33623 -218 33657
rect -252 33555 -218 33589
rect -252 33487 -218 33521
rect -252 33419 -218 33453
rect -252 33351 -218 33385
rect -252 33283 -218 33317
rect -252 33215 -218 33249
rect -252 33147 -218 33181
rect -252 33079 -218 33113
rect -252 33011 -218 33045
rect -252 32943 -218 32977
rect -252 32875 -218 32909
rect -252 32807 -218 32841
rect -252 32739 -218 32773
rect -252 32671 -218 32705
rect -252 32603 -218 32637
rect -252 32535 -218 32569
rect -252 32467 -218 32501
rect -252 32399 -218 32433
rect -252 32331 -218 32365
rect -252 32263 -218 32297
rect -252 32195 -218 32229
rect -252 32127 -218 32161
rect -252 32059 -218 32093
rect -252 31991 -218 32025
rect -252 31923 -218 31957
rect -252 31855 -218 31889
rect -252 31787 -218 31821
rect -252 31719 -218 31753
rect -252 31651 -218 31685
rect -252 31583 -218 31617
rect -252 31515 -218 31549
rect -252 31447 -218 31481
rect -252 31379 -218 31413
rect -252 31311 -218 31345
rect -252 31243 -218 31277
rect -252 31175 -218 31209
rect -252 31107 -218 31141
rect -252 31039 -218 31073
rect -252 30971 -218 31005
rect -252 30903 -218 30937
rect -252 30835 -218 30869
rect -252 30767 -218 30801
rect -252 30699 -218 30733
rect -252 30631 -218 30665
rect -252 30563 -218 30597
rect -252 30495 -218 30529
rect -252 30427 -218 30461
rect -252 30359 -218 30393
rect -252 30291 -218 30325
rect -252 30223 -218 30257
rect -252 30155 -218 30189
rect -252 30087 -218 30121
rect -252 30019 -218 30053
rect -252 29951 -218 29985
rect -252 29883 -218 29917
rect -252 29815 -218 29849
rect -252 29747 -218 29781
rect -252 29679 -218 29713
rect -252 29611 -218 29645
rect -252 29543 -218 29577
rect -252 29475 -218 29509
rect -252 29407 -218 29441
rect -252 29339 -218 29373
rect -252 29271 -218 29305
rect -252 29203 -218 29237
rect -252 29135 -218 29169
rect -252 29067 -218 29101
rect -252 28999 -218 29033
rect -252 28931 -218 28965
rect -252 28863 -218 28897
rect -252 28795 -218 28829
rect -252 28727 -218 28761
rect -252 28659 -218 28693
rect -252 28591 -218 28625
rect -252 28523 -218 28557
rect -252 28455 -218 28489
rect -252 28387 -218 28421
rect -252 28319 -218 28353
rect -252 28251 -218 28285
rect -252 28183 -218 28217
rect -252 28115 -218 28149
rect -252 28047 -218 28081
rect -252 27979 -218 28013
rect -252 27911 -218 27945
rect -252 27843 -218 27877
rect -252 27775 -218 27809
rect -252 27707 -218 27741
rect -252 27639 -218 27673
rect -252 27571 -218 27605
rect -252 27503 -218 27537
rect -252 27435 -218 27469
rect -252 27367 -218 27401
rect -252 27299 -218 27333
rect -252 27231 -218 27265
rect -252 27163 -218 27197
rect -252 27095 -218 27129
rect -252 27027 -218 27061
rect -252 26959 -218 26993
rect -252 26891 -218 26925
rect -252 26823 -218 26857
rect -252 26755 -218 26789
rect -252 26687 -218 26721
rect -252 26619 -218 26653
rect -252 26551 -218 26585
rect -252 26483 -218 26517
rect -252 26415 -218 26449
rect -252 26347 -218 26381
rect -252 26279 -218 26313
rect -252 26211 -218 26245
rect -252 26143 -218 26177
rect -252 26075 -218 26109
rect -252 26007 -218 26041
rect -252 25939 -218 25973
rect -252 25871 -218 25905
rect -252 25803 -218 25837
rect -252 25735 -218 25769
rect -252 25667 -218 25701
rect -252 25599 -218 25633
rect -252 25531 -218 25565
rect -252 25463 -218 25497
rect -252 25395 -218 25429
rect -252 25327 -218 25361
rect -252 25259 -218 25293
rect -252 25191 -218 25225
rect -252 25123 -218 25157
rect -252 25055 -218 25089
rect -252 24987 -218 25021
rect -252 24919 -218 24953
rect -252 24851 -218 24885
rect -252 24783 -218 24817
rect -252 24715 -218 24749
rect -252 24647 -218 24681
rect -252 24579 -218 24613
rect -252 24511 -218 24545
rect -252 24443 -218 24477
rect -252 24375 -218 24409
rect -252 24307 -218 24341
rect -252 24239 -218 24273
rect -252 24171 -218 24205
rect -252 24103 -218 24137
rect -252 24035 -218 24069
rect -252 23967 -218 24001
rect -252 23899 -218 23933
rect -252 23831 -218 23865
rect -252 23763 -218 23797
rect -252 23695 -218 23729
rect -252 23627 -218 23661
rect -252 23559 -218 23593
rect -252 23491 -218 23525
rect -252 23423 -218 23457
rect -252 23355 -218 23389
rect -252 23287 -218 23321
rect -252 23219 -218 23253
rect -252 23151 -218 23185
rect -252 23083 -218 23117
rect -252 23015 -218 23049
rect -252 22947 -218 22981
rect -252 22879 -218 22913
rect -252 22811 -218 22845
rect -252 22743 -218 22777
rect -252 22675 -218 22709
rect -252 22607 -218 22641
rect -252 22539 -218 22573
rect -252 22471 -218 22505
rect -252 22403 -218 22437
rect -252 22335 -218 22369
rect -252 22267 -218 22301
rect -252 22199 -218 22233
rect -252 22131 -218 22165
rect -252 22063 -218 22097
rect -252 21995 -218 22029
rect -252 21927 -218 21961
rect -252 21859 -218 21893
rect -252 21791 -218 21825
rect -252 21723 -218 21757
rect -252 21655 -218 21689
rect -252 21587 -218 21621
rect -252 21519 -218 21553
rect -252 21451 -218 21485
rect -252 21383 -218 21417
rect -252 21315 -218 21349
rect -252 21247 -218 21281
rect -252 21179 -218 21213
rect -252 21111 -218 21145
rect -252 21043 -218 21077
rect -252 20975 -218 21009
rect -252 20907 -218 20941
rect -252 20839 -218 20873
rect -252 20771 -218 20805
rect -252 20703 -218 20737
rect -252 20635 -218 20669
rect -252 20567 -218 20601
rect -252 20499 -218 20533
rect -252 20431 -218 20465
rect -252 20363 -218 20397
rect -252 20295 -218 20329
rect -252 20227 -218 20261
rect -252 20159 -218 20193
rect -252 20091 -218 20125
rect -252 20023 -218 20057
rect -252 19955 -218 19989
rect -252 19887 -218 19921
rect -252 19819 -218 19853
rect -252 19751 -218 19785
rect -252 19683 -218 19717
rect -252 19615 -218 19649
rect -252 19547 -218 19581
rect -252 19479 -218 19513
rect -252 19411 -218 19445
rect -252 19343 -218 19377
rect -252 19275 -218 19309
rect -252 19207 -218 19241
rect -252 19139 -218 19173
rect -252 19071 -218 19105
rect -252 19003 -218 19037
rect -252 18935 -218 18969
rect -252 18867 -218 18901
rect -252 18799 -218 18833
rect -252 18731 -218 18765
rect -252 18663 -218 18697
rect -252 18595 -218 18629
rect -252 18527 -218 18561
rect -252 18459 -218 18493
rect -252 18391 -218 18425
rect -252 18323 -218 18357
rect -252 18255 -218 18289
rect -252 18187 -218 18221
rect -252 18119 -218 18153
rect -252 18051 -218 18085
rect -252 17983 -218 18017
rect -252 17915 -218 17949
rect -252 17847 -218 17881
rect -252 17779 -218 17813
rect -252 17711 -218 17745
rect -252 17643 -218 17677
rect -252 17575 -218 17609
rect -252 17507 -218 17541
rect -252 17439 -218 17473
rect -252 17371 -218 17405
rect -252 17303 -218 17337
rect -252 17235 -218 17269
rect -252 17167 -218 17201
rect -252 17099 -218 17133
rect -252 17031 -218 17065
rect -252 16963 -218 16997
rect -252 16895 -218 16929
rect -252 16827 -218 16861
rect -252 16759 -218 16793
rect -252 16691 -218 16725
rect -252 16623 -218 16657
rect -252 16555 -218 16589
rect -252 16487 -218 16521
rect -252 16419 -218 16453
rect -252 16351 -218 16385
rect -252 16283 -218 16317
rect -252 16215 -218 16249
rect -252 16147 -218 16181
rect -252 16079 -218 16113
rect -252 16011 -218 16045
rect -252 15943 -218 15977
rect -252 15875 -218 15909
rect -252 15807 -218 15841
rect -252 15739 -218 15773
rect -252 15671 -218 15705
rect -252 15603 -218 15637
rect -252 15535 -218 15569
rect -252 15467 -218 15501
rect -252 15399 -218 15433
rect -252 15331 -218 15365
rect -252 15263 -218 15297
rect -252 15195 -218 15229
rect -252 15127 -218 15161
rect -252 15059 -218 15093
rect -252 14991 -218 15025
rect -252 14923 -218 14957
rect -252 14855 -218 14889
rect -252 14787 -218 14821
rect -252 14719 -218 14753
rect -252 14651 -218 14685
rect -252 14583 -218 14617
rect -252 14515 -218 14549
rect -252 14447 -218 14481
rect -252 14379 -218 14413
rect -252 14311 -218 14345
rect -252 14243 -218 14277
rect -252 14175 -218 14209
rect -252 14107 -218 14141
rect -252 14039 -218 14073
rect -252 13971 -218 14005
rect -252 13903 -218 13937
rect -252 13835 -218 13869
rect -252 13767 -218 13801
rect -252 13699 -218 13733
rect -252 13631 -218 13665
rect -252 13563 -218 13597
rect -252 13495 -218 13529
rect -252 13427 -218 13461
rect -252 13359 -218 13393
rect -252 13291 -218 13325
rect -252 13223 -218 13257
rect -252 13155 -218 13189
rect -252 13087 -218 13121
rect -252 13019 -218 13053
rect -252 12951 -218 12985
rect -252 12883 -218 12917
rect -252 12815 -218 12849
rect -252 12747 -218 12781
rect -252 12679 -218 12713
rect -252 12611 -218 12645
rect -252 12543 -218 12577
rect -252 12475 -218 12509
rect -252 12407 -218 12441
rect -252 12339 -218 12373
rect -252 12271 -218 12305
rect -252 12203 -218 12237
rect -252 12135 -218 12169
rect -252 12067 -218 12101
rect -252 11999 -218 12033
rect -252 11931 -218 11965
rect -252 11863 -218 11897
rect -252 11795 -218 11829
rect -252 11727 -218 11761
rect -252 11659 -218 11693
rect -252 11591 -218 11625
rect -252 11523 -218 11557
rect -252 11455 -218 11489
rect -252 11387 -218 11421
rect -252 11319 -218 11353
rect -252 11251 -218 11285
rect -252 11183 -218 11217
rect -252 11115 -218 11149
rect -252 11047 -218 11081
rect -252 10979 -218 11013
rect -252 10911 -218 10945
rect -252 10843 -218 10877
rect -252 10775 -218 10809
rect -252 10707 -218 10741
rect -252 10639 -218 10673
rect -252 10571 -218 10605
rect -252 10503 -218 10537
rect -252 10435 -218 10469
rect -252 10367 -218 10401
rect -252 10299 -218 10333
rect -252 10231 -218 10265
rect -252 10163 -218 10197
rect -252 10095 -218 10129
rect -252 10027 -218 10061
rect -252 9959 -218 9993
rect -252 9891 -218 9925
rect -252 9823 -218 9857
rect -252 9755 -218 9789
rect -252 9687 -218 9721
rect -252 9619 -218 9653
rect -252 9551 -218 9585
rect -252 9483 -218 9517
rect -252 9415 -218 9449
rect -252 9347 -218 9381
rect -252 9279 -218 9313
rect -252 9211 -218 9245
rect -252 9143 -218 9177
rect -252 9075 -218 9109
rect -252 9007 -218 9041
rect -252 8939 -218 8973
rect -252 8871 -218 8905
rect -252 8803 -218 8837
rect -252 8735 -218 8769
rect -252 8667 -218 8701
rect -252 8599 -218 8633
rect -252 8531 -218 8565
rect -252 8463 -218 8497
rect -252 8395 -218 8429
rect -252 8327 -218 8361
rect -252 8259 -218 8293
rect -252 8191 -218 8225
rect -252 8123 -218 8157
rect -252 8055 -218 8089
rect -252 7987 -218 8021
rect -252 7919 -218 7953
rect -252 7851 -218 7885
rect -252 7783 -218 7817
rect -252 7715 -218 7749
rect -252 7647 -218 7681
rect -252 7579 -218 7613
rect -252 7511 -218 7545
rect -252 7443 -218 7477
rect -252 7375 -218 7409
rect -252 7307 -218 7341
rect -252 7239 -218 7273
rect -252 7171 -218 7205
rect -252 7103 -218 7137
rect -252 7035 -218 7069
rect -252 6967 -218 7001
rect -252 6899 -218 6933
rect -252 6831 -218 6865
rect -252 6763 -218 6797
rect -252 6695 -218 6729
rect -252 6627 -218 6661
rect -252 6559 -218 6593
rect -252 6491 -218 6525
rect -252 6423 -218 6457
rect -252 6355 -218 6389
rect -252 6287 -218 6321
rect -252 6219 -218 6253
rect -252 6151 -218 6185
rect -252 6083 -218 6117
rect -252 6015 -218 6049
rect -252 5947 -218 5981
rect -252 5879 -218 5913
rect -252 5811 -218 5845
rect -252 5743 -218 5777
rect -252 5675 -218 5709
rect -252 5607 -218 5641
rect -252 5539 -218 5573
rect -252 5471 -218 5505
rect -252 5403 -218 5437
rect -252 5335 -218 5369
rect -252 5267 -218 5301
rect -252 5199 -218 5233
rect -252 5131 -218 5165
rect -252 5063 -218 5097
rect -252 4995 -218 5029
rect -252 4927 -218 4961
rect -252 4859 -218 4893
rect -252 4791 -218 4825
rect -252 4723 -218 4757
rect -252 4655 -218 4689
rect -252 4587 -218 4621
rect -252 4519 -218 4553
rect -252 4451 -218 4485
rect -252 4383 -218 4417
rect -252 4315 -218 4349
rect -252 4247 -218 4281
rect -252 4179 -218 4213
rect -252 4111 -218 4145
rect -252 4043 -218 4077
rect -252 3975 -218 4009
rect -252 3907 -218 3941
rect -252 3839 -218 3873
rect -252 3771 -218 3805
rect -252 3703 -218 3737
rect -252 3635 -218 3669
rect -252 3567 -218 3601
rect -252 3499 -218 3533
rect 1830 38607 1864 38641
rect 1830 38539 1864 38573
rect 1830 38471 1864 38505
rect 1830 38403 1864 38437
rect 1830 38335 1864 38369
rect 1830 38267 1864 38301
rect 1830 38199 1864 38233
rect 1830 38131 1864 38165
rect 1830 38063 1864 38097
rect 1830 37995 1864 38029
rect 1830 37927 1864 37961
rect 1830 37859 1864 37893
rect 1830 37791 1864 37825
rect 1830 37723 1864 37757
rect 1830 37655 1864 37689
rect 1830 37587 1864 37621
rect 1830 37519 1864 37553
rect 1830 37451 1864 37485
rect 1830 37383 1864 37417
rect 1830 37315 1864 37349
rect 1830 37247 1864 37281
rect 1830 37179 1864 37213
rect 1830 37111 1864 37145
rect 1830 37043 1864 37077
rect 1830 36975 1864 37009
rect 1830 36907 1864 36941
rect 1830 36839 1864 36873
rect 1830 36771 1864 36805
rect 1830 36703 1864 36737
rect 1830 36635 1864 36669
rect 1830 36567 1864 36601
rect 1830 36499 1864 36533
rect 1830 36431 1864 36465
rect 1830 36363 1864 36397
rect 1830 36295 1864 36329
rect 1830 36227 1864 36261
rect 1830 36159 1864 36193
rect 1830 36091 1864 36125
rect 1830 36023 1864 36057
rect 1830 35955 1864 35989
rect 1830 35887 1864 35921
rect 1830 35819 1864 35853
rect 1830 35751 1864 35785
rect 1830 35683 1864 35717
rect 1830 35615 1864 35649
rect 1830 35547 1864 35581
rect 1830 35479 1864 35513
rect 1830 35411 1864 35445
rect 1830 35343 1864 35377
rect 1830 35275 1864 35309
rect 1830 35207 1864 35241
rect 1830 35139 1864 35173
rect 1830 35071 1864 35105
rect 1830 35003 1864 35037
rect 1830 34935 1864 34969
rect 1830 34867 1864 34901
rect 1830 34799 1864 34833
rect 1830 34731 1864 34765
rect 1830 34663 1864 34697
rect 1830 34595 1864 34629
rect 1830 34527 1864 34561
rect 1830 34459 1864 34493
rect 1830 34391 1864 34425
rect 1830 34323 1864 34357
rect 1830 34255 1864 34289
rect 1830 34187 1864 34221
rect 1830 34119 1864 34153
rect 1830 34051 1864 34085
rect 1830 33983 1864 34017
rect 1830 33915 1864 33949
rect 1830 33847 1864 33881
rect 1830 33779 1864 33813
rect 1830 33711 1864 33745
rect 1830 33643 1864 33677
rect 1830 33575 1864 33609
rect 1830 33507 1864 33541
rect 1830 33439 1864 33473
rect 1830 33371 1864 33405
rect 1830 33303 1864 33337
rect 1830 33235 1864 33269
rect 1830 33167 1864 33201
rect 1830 33099 1864 33133
rect 1830 33031 1864 33065
rect 1830 32963 1864 32997
rect 1830 32895 1864 32929
rect 1830 32827 1864 32861
rect 1830 32759 1864 32793
rect 1830 32691 1864 32725
rect 1830 32623 1864 32657
rect 1830 32555 1864 32589
rect 1830 32487 1864 32521
rect 1830 32419 1864 32453
rect 1830 32351 1864 32385
rect 1830 32283 1864 32317
rect 1830 32215 1864 32249
rect 1830 32147 1864 32181
rect 1830 32079 1864 32113
rect 1830 32011 1864 32045
rect 1830 31943 1864 31977
rect 1830 31875 1864 31909
rect 1830 31807 1864 31841
rect 1830 31739 1864 31773
rect 1830 31671 1864 31705
rect 1830 31603 1864 31637
rect 1830 31535 1864 31569
rect 1830 31467 1864 31501
rect 1830 31399 1864 31433
rect 1830 31331 1864 31365
rect 1830 31263 1864 31297
rect 1830 31195 1864 31229
rect 1830 31127 1864 31161
rect 1830 31059 1864 31093
rect 1830 30991 1864 31025
rect 1830 30923 1864 30957
rect 1830 30855 1864 30889
rect 1830 30787 1864 30821
rect 1830 30719 1864 30753
rect 1830 30651 1864 30685
rect 1830 30583 1864 30617
rect 1830 30515 1864 30549
rect 1830 30447 1864 30481
rect 1830 30379 1864 30413
rect 1830 30311 1864 30345
rect 1830 30243 1864 30277
rect 1830 30175 1864 30209
rect 1830 30107 1864 30141
rect 1830 30039 1864 30073
rect 1830 29971 1864 30005
rect 1830 29903 1864 29937
rect 1830 29835 1864 29869
rect 1830 29767 1864 29801
rect 1830 29699 1864 29733
rect 1830 29631 1864 29665
rect 1830 29563 1864 29597
rect 1830 29495 1864 29529
rect 1830 29427 1864 29461
rect 1830 29359 1864 29393
rect 1830 29291 1864 29325
rect 1830 29223 1864 29257
rect 1830 29155 1864 29189
rect 1830 29087 1864 29121
rect 1830 29019 1864 29053
rect 1830 28951 1864 28985
rect 1830 28883 1864 28917
rect 1830 28815 1864 28849
rect 1830 28747 1864 28781
rect 1830 28679 1864 28713
rect 1830 28611 1864 28645
rect 1830 28543 1864 28577
rect 1830 28475 1864 28509
rect 1830 28407 1864 28441
rect 1830 28339 1864 28373
rect 1830 28271 1864 28305
rect 1830 28203 1864 28237
rect 1830 28135 1864 28169
rect 1830 28067 1864 28101
rect 1830 27999 1864 28033
rect 1830 27931 1864 27965
rect 1830 27863 1864 27897
rect 1830 27795 1864 27829
rect 1830 27727 1864 27761
rect 1830 27659 1864 27693
rect 1830 27591 1864 27625
rect 1830 27523 1864 27557
rect 1830 27455 1864 27489
rect 1830 27387 1864 27421
rect 1830 27319 1864 27353
rect 1830 27251 1864 27285
rect 1830 27183 1864 27217
rect 1830 27115 1864 27149
rect 1830 27047 1864 27081
rect 1830 26979 1864 27013
rect 1830 26911 1864 26945
rect 1830 26843 1864 26877
rect 1830 26775 1864 26809
rect 1830 26707 1864 26741
rect 1830 26639 1864 26673
rect 1830 26571 1864 26605
rect 1830 26503 1864 26537
rect 1830 26435 1864 26469
rect 1830 26367 1864 26401
rect 1830 26299 1864 26333
rect 1830 26231 1864 26265
rect 1830 26163 1864 26197
rect 1830 26095 1864 26129
rect 1830 26027 1864 26061
rect 1830 25959 1864 25993
rect 1830 25891 1864 25925
rect 1830 25823 1864 25857
rect 1830 25755 1864 25789
rect 1830 25687 1864 25721
rect 1830 25619 1864 25653
rect 1830 25551 1864 25585
rect 1830 25483 1864 25517
rect 1830 25415 1864 25449
rect 1830 25347 1864 25381
rect 1830 25279 1864 25313
rect 1830 25211 1864 25245
rect 1830 25143 1864 25177
rect 1830 25075 1864 25109
rect 1830 25007 1864 25041
rect 1830 24939 1864 24973
rect 1830 24871 1864 24905
rect 1830 24803 1864 24837
rect 1830 24735 1864 24769
rect 1830 24667 1864 24701
rect 1830 24599 1864 24633
rect 1830 24531 1864 24565
rect 1830 24463 1864 24497
rect 1830 24395 1864 24429
rect 1830 24327 1864 24361
rect 1830 24259 1864 24293
rect 1830 24191 1864 24225
rect 1830 24123 1864 24157
rect 1830 24055 1864 24089
rect 1830 23987 1864 24021
rect 1830 23919 1864 23953
rect 1830 23851 1864 23885
rect 1830 23783 1864 23817
rect 1830 23715 1864 23749
rect 1830 23647 1864 23681
rect 1830 23579 1864 23613
rect 1830 23511 1864 23545
rect 1830 23443 1864 23477
rect 1830 23375 1864 23409
rect 1830 23307 1864 23341
rect 1830 23239 1864 23273
rect 1830 23171 1864 23205
rect 1830 23103 1864 23137
rect 1830 23035 1864 23069
rect 1830 22967 1864 23001
rect 1830 22899 1864 22933
rect 1830 22831 1864 22865
rect 1830 22763 1864 22797
rect 1830 22695 1864 22729
rect 1830 22627 1864 22661
rect 1830 22559 1864 22593
rect 1830 22491 1864 22525
rect 1830 22423 1864 22457
rect 1830 22355 1864 22389
rect 1830 22287 1864 22321
rect 1830 22219 1864 22253
rect 1830 22151 1864 22185
rect 1830 22083 1864 22117
rect 1830 22015 1864 22049
rect 1830 21947 1864 21981
rect 1830 21879 1864 21913
rect 1830 21811 1864 21845
rect 1830 21743 1864 21777
rect 1830 21675 1864 21709
rect 1830 21607 1864 21641
rect 1830 21539 1864 21573
rect 1830 21471 1864 21505
rect 1830 21403 1864 21437
rect 1830 21335 1864 21369
rect 1830 21267 1864 21301
rect 1830 21199 1864 21233
rect 1830 21131 1864 21165
rect 1830 21063 1864 21097
rect 1830 20995 1864 21029
rect 1830 20927 1864 20961
rect 1830 20859 1864 20893
rect 1830 20791 1864 20825
rect 1830 20723 1864 20757
rect 1830 20655 1864 20689
rect 1830 20587 1864 20621
rect 1830 20519 1864 20553
rect 1830 20451 1864 20485
rect 1830 20383 1864 20417
rect 1830 20315 1864 20349
rect 1830 20247 1864 20281
rect 1830 20179 1864 20213
rect 1830 20111 1864 20145
rect 1830 20043 1864 20077
rect 1830 19975 1864 20009
rect 1830 19907 1864 19941
rect 1830 19839 1864 19873
rect 1830 19771 1864 19805
rect 1830 19703 1864 19737
rect 1830 19635 1864 19669
rect 1830 19567 1864 19601
rect 1830 19499 1864 19533
rect 1830 19431 1864 19465
rect 1830 19363 1864 19397
rect 1830 19295 1864 19329
rect 1830 19227 1864 19261
rect 1830 19159 1864 19193
rect 1830 19091 1864 19125
rect 1830 19023 1864 19057
rect 1830 18955 1864 18989
rect 1830 18887 1864 18921
rect 1830 18819 1864 18853
rect 1830 18751 1864 18785
rect 1830 18683 1864 18717
rect 1830 18615 1864 18649
rect 1830 18547 1864 18581
rect 1830 18479 1864 18513
rect 1830 18411 1864 18445
rect 1830 18343 1864 18377
rect 1830 18275 1864 18309
rect 1830 18207 1864 18241
rect 1830 18139 1864 18173
rect 1830 18071 1864 18105
rect 1830 18003 1864 18037
rect 1830 17935 1864 17969
rect 1830 17867 1864 17901
rect 1830 17799 1864 17833
rect 1830 17731 1864 17765
rect 1830 17663 1864 17697
rect 1830 17595 1864 17629
rect 1830 17527 1864 17561
rect 1830 17459 1864 17493
rect 1830 17391 1864 17425
rect 1830 17323 1864 17357
rect 1830 17255 1864 17289
rect 1830 17187 1864 17221
rect 1830 17119 1864 17153
rect 1830 17051 1864 17085
rect 1830 16983 1864 17017
rect 1830 16915 1864 16949
rect 1830 16847 1864 16881
rect 1830 16779 1864 16813
rect 1830 16711 1864 16745
rect 1830 16643 1864 16677
rect 1830 16575 1864 16609
rect 1830 16507 1864 16541
rect 1830 16439 1864 16473
rect 1830 16371 1864 16405
rect 1830 16303 1864 16337
rect 1830 16235 1864 16269
rect 1830 16167 1864 16201
rect 1830 16099 1864 16133
rect 1830 16031 1864 16065
rect 1830 15963 1864 15997
rect 1830 15895 1864 15929
rect 1830 15827 1864 15861
rect 1830 15759 1864 15793
rect 1830 15691 1864 15725
rect 1830 15623 1864 15657
rect 1830 15555 1864 15589
rect 1830 15487 1864 15521
rect 1830 15419 1864 15453
rect 1830 15351 1864 15385
rect 1830 15283 1864 15317
rect 1830 15215 1864 15249
rect 1830 15147 1864 15181
rect 1830 15079 1864 15113
rect 1830 15011 1864 15045
rect 1830 14943 1864 14977
rect 1830 14875 1864 14909
rect 1830 14807 1864 14841
rect 1830 14739 1864 14773
rect 1830 14671 1864 14705
rect 1830 14603 1864 14637
rect 1830 14535 1864 14569
rect 1830 14467 1864 14501
rect 1830 14399 1864 14433
rect 1830 14331 1864 14365
rect 1830 14263 1864 14297
rect 1830 14195 1864 14229
rect 1830 14127 1864 14161
rect 1830 14059 1864 14093
rect 1830 13991 1864 14025
rect 1830 13923 1864 13957
rect 1830 13855 1864 13889
rect 1830 13787 1864 13821
rect 1830 13719 1864 13753
rect 1830 13651 1864 13685
rect 1830 13583 1864 13617
rect 1830 13515 1864 13549
rect 1830 13447 1864 13481
rect 1830 13379 1864 13413
rect 1830 13311 1864 13345
rect 1830 13243 1864 13277
rect 1830 13175 1864 13209
rect 1830 13107 1864 13141
rect 1830 13039 1864 13073
rect 1830 12971 1864 13005
rect 1830 12903 1864 12937
rect 1830 12835 1864 12869
rect 1830 12767 1864 12801
rect 1830 12699 1864 12733
rect 1830 12631 1864 12665
rect 1830 12563 1864 12597
rect 1830 12495 1864 12529
rect 1830 12427 1864 12461
rect 1830 12359 1864 12393
rect 1830 12291 1864 12325
rect 1830 12223 1864 12257
rect 1830 12155 1864 12189
rect 1830 12087 1864 12121
rect 1830 12019 1864 12053
rect 1830 11951 1864 11985
rect 1830 11883 1864 11917
rect 1830 11815 1864 11849
rect 1830 11747 1864 11781
rect 1830 11679 1864 11713
rect 1830 11611 1864 11645
rect 1830 11543 1864 11577
rect 1830 11475 1864 11509
rect 1830 11407 1864 11441
rect 1830 11339 1864 11373
rect 1830 11271 1864 11305
rect 1830 11203 1864 11237
rect 1830 11135 1864 11169
rect 1830 11067 1864 11101
rect 1830 10999 1864 11033
rect 1830 10931 1864 10965
rect 1830 10863 1864 10897
rect 1830 10795 1864 10829
rect 1830 10727 1864 10761
rect 1830 10659 1864 10693
rect 1830 10591 1864 10625
rect 1830 10523 1864 10557
rect 1830 10455 1864 10489
rect 1830 10387 1864 10421
rect 1830 10319 1864 10353
rect 1830 10251 1864 10285
rect 1830 10183 1864 10217
rect 1830 10115 1864 10149
rect 1830 10047 1864 10081
rect 1830 9979 1864 10013
rect 1830 9911 1864 9945
rect 1830 9843 1864 9877
rect 1830 9775 1864 9809
rect 1830 9707 1864 9741
rect 1830 9639 1864 9673
rect 1830 9571 1864 9605
rect 1830 9503 1864 9537
rect 1830 9435 1864 9469
rect 1830 9367 1864 9401
rect 1830 9299 1864 9333
rect 1830 9231 1864 9265
rect 1830 9163 1864 9197
rect 1830 9095 1864 9129
rect 1830 9027 1864 9061
rect 1830 8959 1864 8993
rect 1830 8891 1864 8925
rect 1830 8823 1864 8857
rect 1830 8755 1864 8789
rect 1830 8687 1864 8721
rect 1830 8619 1864 8653
rect 1830 8551 1864 8585
rect 1830 8483 1864 8517
rect 1830 8415 1864 8449
rect 1830 8347 1864 8381
rect 1830 8279 1864 8313
rect 1830 8211 1864 8245
rect 1830 8143 1864 8177
rect 1830 8075 1864 8109
rect 1830 8007 1864 8041
rect 1830 7939 1864 7973
rect 1830 7871 1864 7905
rect 1830 7803 1864 7837
rect 1830 7735 1864 7769
rect 1830 7667 1864 7701
rect 1830 7599 1864 7633
rect 1830 7531 1864 7565
rect 1830 7463 1864 7497
rect 1830 7395 1864 7429
rect 1830 7327 1864 7361
rect 1830 7259 1864 7293
rect 1830 7191 1864 7225
rect 1830 7123 1864 7157
rect 1830 7055 1864 7089
rect 1830 6987 1864 7021
rect 1830 6919 1864 6953
rect 1830 6851 1864 6885
rect 1830 6783 1864 6817
rect 1830 6715 1864 6749
rect 1830 6647 1864 6681
rect 1830 6579 1864 6613
rect 1830 6511 1864 6545
rect 1830 6443 1864 6477
rect 1830 6375 1864 6409
rect 1830 6307 1864 6341
rect 1830 6239 1864 6273
rect 1830 6171 1864 6205
rect 1830 6103 1864 6137
rect 1830 6035 1864 6069
rect 1830 5967 1864 6001
rect 1830 5899 1864 5933
rect 1830 5831 1864 5865
rect 1830 5763 1864 5797
rect 1830 5695 1864 5729
rect 1830 5627 1864 5661
rect 1830 5559 1864 5593
rect 1830 5491 1864 5525
rect 1830 5423 1864 5457
rect 1830 5355 1864 5389
rect 1830 5287 1864 5321
rect 1830 5219 1864 5253
rect 1830 5151 1864 5185
rect 1830 5083 1864 5117
rect 1830 5015 1864 5049
rect 1830 4947 1864 4981
rect 1830 4879 1864 4913
rect 1830 4811 1864 4845
rect 1830 4743 1864 4777
rect 1830 4675 1864 4709
rect 1830 4607 1864 4641
rect 1830 4539 1864 4573
rect 1830 4471 1864 4505
rect 1830 4403 1864 4437
rect 1830 4335 1864 4369
rect 1830 4267 1864 4301
rect 1830 4199 1864 4233
rect 1830 4131 1864 4165
rect 1830 4063 1864 4097
rect 1830 3995 1864 4029
rect 1830 3927 1864 3961
rect 1830 3859 1864 3893
rect 1830 3791 1864 3825
rect 1830 3723 1864 3757
rect 1830 3655 1864 3689
rect 1830 3587 1864 3621
rect 1830 3519 1864 3553
rect -252 3431 -218 3465
rect -252 3363 -218 3397
rect 1830 3451 1864 3485
rect 3972 38655 4006 38689
rect 3972 38587 4006 38621
rect 3972 38519 4006 38553
rect 3972 38451 4006 38485
rect 3972 38383 4006 38417
rect 3972 38315 4006 38349
rect 3972 38247 4006 38281
rect 3972 38179 4006 38213
rect 3972 38111 4006 38145
rect 3972 38043 4006 38077
rect 3972 37975 4006 38009
rect 3972 37907 4006 37941
rect 3972 37839 4006 37873
rect 3972 37771 4006 37805
rect 3972 37703 4006 37737
rect 3972 37635 4006 37669
rect 3972 37567 4006 37601
rect 3972 37499 4006 37533
rect 3972 37431 4006 37465
rect 3972 37363 4006 37397
rect 3972 37295 4006 37329
rect 3972 37227 4006 37261
rect 3972 37159 4006 37193
rect 3972 37091 4006 37125
rect 3972 37023 4006 37057
rect 3972 36955 4006 36989
rect 3972 36887 4006 36921
rect 3972 36819 4006 36853
rect 3972 36751 4006 36785
rect 3972 36683 4006 36717
rect 3972 36615 4006 36649
rect 3972 36547 4006 36581
rect 3972 36479 4006 36513
rect 3972 36411 4006 36445
rect 3972 36343 4006 36377
rect 3972 36275 4006 36309
rect 3972 36207 4006 36241
rect 3972 36139 4006 36173
rect 3972 36071 4006 36105
rect 3972 36003 4006 36037
rect 3972 35935 4006 35969
rect 3972 35867 4006 35901
rect 3972 35799 4006 35833
rect 3972 35731 4006 35765
rect 3972 35663 4006 35697
rect 3972 35595 4006 35629
rect 3972 35527 4006 35561
rect 3972 35459 4006 35493
rect 3972 35391 4006 35425
rect 3972 35323 4006 35357
rect 3972 35255 4006 35289
rect 3972 35187 4006 35221
rect 3972 35119 4006 35153
rect 3972 35051 4006 35085
rect 3972 34983 4006 35017
rect 3972 34915 4006 34949
rect 3972 34847 4006 34881
rect 3972 34779 4006 34813
rect 3972 34711 4006 34745
rect 3972 34643 4006 34677
rect 3972 34575 4006 34609
rect 3972 34507 4006 34541
rect 3972 34439 4006 34473
rect 3972 34371 4006 34405
rect 3972 34303 4006 34337
rect 3972 34235 4006 34269
rect 3972 34167 4006 34201
rect 3972 34099 4006 34133
rect 3972 34031 4006 34065
rect 3972 33963 4006 33997
rect 3972 33895 4006 33929
rect 3972 33827 4006 33861
rect 3972 33759 4006 33793
rect 3972 33691 4006 33725
rect 3972 33623 4006 33657
rect 3972 33555 4006 33589
rect 3972 33487 4006 33521
rect 3972 33419 4006 33453
rect 3972 33351 4006 33385
rect 3972 33283 4006 33317
rect 3972 33215 4006 33249
rect 3972 33147 4006 33181
rect 3972 33079 4006 33113
rect 3972 33011 4006 33045
rect 3972 32943 4006 32977
rect 3972 32875 4006 32909
rect 3972 32807 4006 32841
rect 3972 32739 4006 32773
rect 3972 32671 4006 32705
rect 3972 32603 4006 32637
rect 3972 32535 4006 32569
rect 3972 32467 4006 32501
rect 3972 32399 4006 32433
rect 3972 32331 4006 32365
rect 3972 32263 4006 32297
rect 3972 32195 4006 32229
rect 3972 32127 4006 32161
rect 3972 32059 4006 32093
rect 3972 31991 4006 32025
rect 3972 31923 4006 31957
rect 3972 31855 4006 31889
rect 3972 31787 4006 31821
rect 3972 31719 4006 31753
rect 3972 31651 4006 31685
rect 3972 31583 4006 31617
rect 3972 31515 4006 31549
rect 3972 31447 4006 31481
rect 3972 31379 4006 31413
rect 3972 31311 4006 31345
rect 3972 31243 4006 31277
rect 3972 31175 4006 31209
rect 3972 31107 4006 31141
rect 3972 31039 4006 31073
rect 3972 30971 4006 31005
rect 3972 30903 4006 30937
rect 3972 30835 4006 30869
rect 3972 30767 4006 30801
rect 3972 30699 4006 30733
rect 3972 30631 4006 30665
rect 3972 30563 4006 30597
rect 3972 30495 4006 30529
rect 3972 30427 4006 30461
rect 3972 30359 4006 30393
rect 3972 30291 4006 30325
rect 3972 30223 4006 30257
rect 3972 30155 4006 30189
rect 3972 30087 4006 30121
rect 3972 30019 4006 30053
rect 3972 29951 4006 29985
rect 3972 29883 4006 29917
rect 3972 29815 4006 29849
rect 3972 29747 4006 29781
rect 3972 29679 4006 29713
rect 3972 29611 4006 29645
rect 3972 29543 4006 29577
rect 3972 29475 4006 29509
rect 3972 29407 4006 29441
rect 3972 29339 4006 29373
rect 3972 29271 4006 29305
rect 3972 29203 4006 29237
rect 3972 29135 4006 29169
rect 3972 29067 4006 29101
rect 3972 28999 4006 29033
rect 3972 28931 4006 28965
rect 3972 28863 4006 28897
rect 3972 28795 4006 28829
rect 3972 28727 4006 28761
rect 3972 28659 4006 28693
rect 3972 28591 4006 28625
rect 3972 28523 4006 28557
rect 3972 28455 4006 28489
rect 3972 28387 4006 28421
rect 3972 28319 4006 28353
rect 3972 28251 4006 28285
rect 3972 28183 4006 28217
rect 3972 28115 4006 28149
rect 3972 28047 4006 28081
rect 3972 27979 4006 28013
rect 3972 27911 4006 27945
rect 3972 27843 4006 27877
rect 3972 27775 4006 27809
rect 3972 27707 4006 27741
rect 3972 27639 4006 27673
rect 3972 27571 4006 27605
rect 3972 27503 4006 27537
rect 3972 27435 4006 27469
rect 3972 27367 4006 27401
rect 3972 27299 4006 27333
rect 3972 27231 4006 27265
rect 3972 27163 4006 27197
rect 3972 27095 4006 27129
rect 3972 27027 4006 27061
rect 3972 26959 4006 26993
rect 3972 26891 4006 26925
rect 3972 26823 4006 26857
rect 3972 26755 4006 26789
rect 3972 26687 4006 26721
rect 3972 26619 4006 26653
rect 3972 26551 4006 26585
rect 3972 26483 4006 26517
rect 3972 26415 4006 26449
rect 3972 26347 4006 26381
rect 3972 26279 4006 26313
rect 3972 26211 4006 26245
rect 3972 26143 4006 26177
rect 3972 26075 4006 26109
rect 3972 26007 4006 26041
rect 3972 25939 4006 25973
rect 3972 25871 4006 25905
rect 3972 25803 4006 25837
rect 3972 25735 4006 25769
rect 3972 25667 4006 25701
rect 3972 25599 4006 25633
rect 3972 25531 4006 25565
rect 3972 25463 4006 25497
rect 3972 25395 4006 25429
rect 3972 25327 4006 25361
rect 3972 25259 4006 25293
rect 3972 25191 4006 25225
rect 3972 25123 4006 25157
rect 3972 25055 4006 25089
rect 3972 24987 4006 25021
rect 3972 24919 4006 24953
rect 3972 24851 4006 24885
rect 3972 24783 4006 24817
rect 3972 24715 4006 24749
rect 3972 24647 4006 24681
rect 3972 24579 4006 24613
rect 3972 24511 4006 24545
rect 3972 24443 4006 24477
rect 3972 24375 4006 24409
rect 3972 24307 4006 24341
rect 3972 24239 4006 24273
rect 3972 24171 4006 24205
rect 3972 24103 4006 24137
rect 3972 24035 4006 24069
rect 3972 23967 4006 24001
rect 3972 23899 4006 23933
rect 3972 23831 4006 23865
rect 3972 23763 4006 23797
rect 3972 23695 4006 23729
rect 3972 23627 4006 23661
rect 3972 23559 4006 23593
rect 3972 23491 4006 23525
rect 3972 23423 4006 23457
rect 3972 23355 4006 23389
rect 3972 23287 4006 23321
rect 3972 23219 4006 23253
rect 3972 23151 4006 23185
rect 3972 23083 4006 23117
rect 3972 23015 4006 23049
rect 3972 22947 4006 22981
rect 3972 22879 4006 22913
rect 3972 22811 4006 22845
rect 3972 22743 4006 22777
rect 3972 22675 4006 22709
rect 3972 22607 4006 22641
rect 3972 22539 4006 22573
rect 3972 22471 4006 22505
rect 3972 22403 4006 22437
rect 3972 22335 4006 22369
rect 3972 22267 4006 22301
rect 3972 22199 4006 22233
rect 3972 22131 4006 22165
rect 3972 22063 4006 22097
rect 3972 21995 4006 22029
rect 3972 21927 4006 21961
rect 3972 21859 4006 21893
rect 3972 21791 4006 21825
rect 3972 21723 4006 21757
rect 3972 21655 4006 21689
rect 3972 21587 4006 21621
rect 3972 21519 4006 21553
rect 3972 21451 4006 21485
rect 3972 21383 4006 21417
rect 3972 21315 4006 21349
rect 3972 21247 4006 21281
rect 3972 21179 4006 21213
rect 3972 21111 4006 21145
rect 3972 21043 4006 21077
rect 3972 20975 4006 21009
rect 3972 20907 4006 20941
rect 3972 20839 4006 20873
rect 3972 20771 4006 20805
rect 3972 20703 4006 20737
rect 3972 20635 4006 20669
rect 3972 20567 4006 20601
rect 3972 20499 4006 20533
rect 3972 20431 4006 20465
rect 3972 20363 4006 20397
rect 3972 20295 4006 20329
rect 3972 20227 4006 20261
rect 3972 20159 4006 20193
rect 3972 20091 4006 20125
rect 3972 20023 4006 20057
rect 3972 19955 4006 19989
rect 3972 19887 4006 19921
rect 3972 19819 4006 19853
rect 3972 19751 4006 19785
rect 3972 19683 4006 19717
rect 3972 19615 4006 19649
rect 3972 19547 4006 19581
rect 3972 19479 4006 19513
rect 3972 19411 4006 19445
rect 3972 19343 4006 19377
rect 3972 19275 4006 19309
rect 3972 19207 4006 19241
rect 3972 19139 4006 19173
rect 3972 19071 4006 19105
rect 3972 19003 4006 19037
rect 3972 18935 4006 18969
rect 3972 18867 4006 18901
rect 3972 18799 4006 18833
rect 3972 18731 4006 18765
rect 3972 18663 4006 18697
rect 3972 18595 4006 18629
rect 3972 18527 4006 18561
rect 3972 18459 4006 18493
rect 3972 18391 4006 18425
rect 3972 18323 4006 18357
rect 3972 18255 4006 18289
rect 3972 18187 4006 18221
rect 3972 18119 4006 18153
rect 3972 18051 4006 18085
rect 3972 17983 4006 18017
rect 3972 17915 4006 17949
rect 3972 17847 4006 17881
rect 3972 17779 4006 17813
rect 3972 17711 4006 17745
rect 3972 17643 4006 17677
rect 3972 17575 4006 17609
rect 3972 17507 4006 17541
rect 3972 17439 4006 17473
rect 3972 17371 4006 17405
rect 3972 17303 4006 17337
rect 3972 17235 4006 17269
rect 3972 17167 4006 17201
rect 3972 17099 4006 17133
rect 3972 17031 4006 17065
rect 3972 16963 4006 16997
rect 3972 16895 4006 16929
rect 3972 16827 4006 16861
rect 3972 16759 4006 16793
rect 3972 16691 4006 16725
rect 3972 16623 4006 16657
rect 3972 16555 4006 16589
rect 3972 16487 4006 16521
rect 3972 16419 4006 16453
rect 3972 16351 4006 16385
rect 3972 16283 4006 16317
rect 3972 16215 4006 16249
rect 3972 16147 4006 16181
rect 3972 16079 4006 16113
rect 3972 16011 4006 16045
rect 3972 15943 4006 15977
rect 3972 15875 4006 15909
rect 3972 15807 4006 15841
rect 3972 15739 4006 15773
rect 3972 15671 4006 15705
rect 3972 15603 4006 15637
rect 3972 15535 4006 15569
rect 3972 15467 4006 15501
rect 3972 15399 4006 15433
rect 3972 15331 4006 15365
rect 3972 15263 4006 15297
rect 3972 15195 4006 15229
rect 3972 15127 4006 15161
rect 3972 15059 4006 15093
rect 3972 14991 4006 15025
rect 3972 14923 4006 14957
rect 3972 14855 4006 14889
rect 3972 14787 4006 14821
rect 3972 14719 4006 14753
rect 3972 14651 4006 14685
rect 3972 14583 4006 14617
rect 3972 14515 4006 14549
rect 3972 14447 4006 14481
rect 3972 14379 4006 14413
rect 3972 14311 4006 14345
rect 3972 14243 4006 14277
rect 3972 14175 4006 14209
rect 3972 14107 4006 14141
rect 3972 14039 4006 14073
rect 3972 13971 4006 14005
rect 3972 13903 4006 13937
rect 3972 13835 4006 13869
rect 3972 13767 4006 13801
rect 3972 13699 4006 13733
rect 3972 13631 4006 13665
rect 3972 13563 4006 13597
rect 3972 13495 4006 13529
rect 3972 13427 4006 13461
rect 3972 13359 4006 13393
rect 3972 13291 4006 13325
rect 3972 13223 4006 13257
rect 3972 13155 4006 13189
rect 3972 13087 4006 13121
rect 3972 13019 4006 13053
rect 3972 12951 4006 12985
rect 3972 12883 4006 12917
rect 3972 12815 4006 12849
rect 3972 12747 4006 12781
rect 3972 12679 4006 12713
rect 3972 12611 4006 12645
rect 3972 12543 4006 12577
rect 3972 12475 4006 12509
rect 3972 12407 4006 12441
rect 3972 12339 4006 12373
rect 3972 12271 4006 12305
rect 3972 12203 4006 12237
rect 3972 12135 4006 12169
rect 3972 12067 4006 12101
rect 3972 11999 4006 12033
rect 3972 11931 4006 11965
rect 3972 11863 4006 11897
rect 3972 11795 4006 11829
rect 3972 11727 4006 11761
rect 3972 11659 4006 11693
rect 3972 11591 4006 11625
rect 3972 11523 4006 11557
rect 3972 11455 4006 11489
rect 3972 11387 4006 11421
rect 3972 11319 4006 11353
rect 3972 11251 4006 11285
rect 3972 11183 4006 11217
rect 3972 11115 4006 11149
rect 3972 11047 4006 11081
rect 3972 10979 4006 11013
rect 3972 10911 4006 10945
rect 3972 10843 4006 10877
rect 3972 10775 4006 10809
rect 3972 10707 4006 10741
rect 3972 10639 4006 10673
rect 3972 10571 4006 10605
rect 3972 10503 4006 10537
rect 3972 10435 4006 10469
rect 3972 10367 4006 10401
rect 3972 10299 4006 10333
rect 3972 10231 4006 10265
rect 3972 10163 4006 10197
rect 3972 10095 4006 10129
rect 3972 10027 4006 10061
rect 3972 9959 4006 9993
rect 3972 9891 4006 9925
rect 3972 9823 4006 9857
rect 3972 9755 4006 9789
rect 3972 9687 4006 9721
rect 3972 9619 4006 9653
rect 3972 9551 4006 9585
rect 3972 9483 4006 9517
rect 3972 9415 4006 9449
rect 3972 9347 4006 9381
rect 3972 9279 4006 9313
rect 3972 9211 4006 9245
rect 3972 9143 4006 9177
rect 3972 9075 4006 9109
rect 3972 9007 4006 9041
rect 3972 8939 4006 8973
rect 3972 8871 4006 8905
rect 3972 8803 4006 8837
rect 3972 8735 4006 8769
rect 3972 8667 4006 8701
rect 3972 8599 4006 8633
rect 3972 8531 4006 8565
rect 3972 8463 4006 8497
rect 3972 8395 4006 8429
rect 3972 8327 4006 8361
rect 3972 8259 4006 8293
rect 3972 8191 4006 8225
rect 3972 8123 4006 8157
rect 3972 8055 4006 8089
rect 3972 7987 4006 8021
rect 3972 7919 4006 7953
rect 3972 7851 4006 7885
rect 3972 7783 4006 7817
rect 3972 7715 4006 7749
rect 3972 7647 4006 7681
rect 3972 7579 4006 7613
rect 3972 7511 4006 7545
rect 3972 7443 4006 7477
rect 3972 7375 4006 7409
rect 3972 7307 4006 7341
rect 3972 7239 4006 7273
rect 3972 7171 4006 7205
rect 3972 7103 4006 7137
rect 3972 7035 4006 7069
rect 3972 6967 4006 7001
rect 3972 6899 4006 6933
rect 3972 6831 4006 6865
rect 3972 6763 4006 6797
rect 3972 6695 4006 6729
rect 3972 6627 4006 6661
rect 3972 6559 4006 6593
rect 3972 6491 4006 6525
rect 3972 6423 4006 6457
rect 3972 6355 4006 6389
rect 3972 6287 4006 6321
rect 3972 6219 4006 6253
rect 3972 6151 4006 6185
rect 3972 6083 4006 6117
rect 3972 6015 4006 6049
rect 3972 5947 4006 5981
rect 3972 5879 4006 5913
rect 3972 5811 4006 5845
rect 3972 5743 4006 5777
rect 3972 5675 4006 5709
rect 3972 5607 4006 5641
rect 3972 5539 4006 5573
rect 3972 5471 4006 5505
rect 3972 5403 4006 5437
rect 3972 5335 4006 5369
rect 3972 5267 4006 5301
rect 3972 5199 4006 5233
rect 3972 5131 4006 5165
rect 3972 5063 4006 5097
rect 3972 4995 4006 5029
rect 3972 4927 4006 4961
rect 3972 4859 4006 4893
rect 3972 4791 4006 4825
rect 3972 4723 4006 4757
rect 3972 4655 4006 4689
rect 3972 4587 4006 4621
rect 3972 4519 4006 4553
rect 3972 4451 4006 4485
rect 3972 4383 4006 4417
rect 3972 4315 4006 4349
rect 3972 4247 4006 4281
rect 3972 4179 4006 4213
rect 3972 4111 4006 4145
rect 3972 4043 4006 4077
rect 3972 3975 4006 4009
rect 3972 3907 4006 3941
rect 3972 3839 4006 3873
rect 3972 3771 4006 3805
rect 3972 3703 4006 3737
rect 3972 3635 4006 3669
rect 3972 3567 4006 3601
rect 3972 3499 4006 3533
rect 1830 3383 1864 3417
rect -252 3295 -218 3329
rect 6114 38607 6148 38641
rect 6114 38539 6148 38573
rect 6114 38471 6148 38505
rect 6114 38403 6148 38437
rect 6114 38335 6148 38369
rect 6114 38267 6148 38301
rect 6114 38199 6148 38233
rect 6114 38131 6148 38165
rect 6114 38063 6148 38097
rect 6114 37995 6148 38029
rect 6114 37927 6148 37961
rect 6114 37859 6148 37893
rect 6114 37791 6148 37825
rect 6114 37723 6148 37757
rect 6114 37655 6148 37689
rect 6114 37587 6148 37621
rect 6114 37519 6148 37553
rect 6114 37451 6148 37485
rect 6114 37383 6148 37417
rect 6114 37315 6148 37349
rect 6114 37247 6148 37281
rect 6114 37179 6148 37213
rect 6114 37111 6148 37145
rect 6114 37043 6148 37077
rect 6114 36975 6148 37009
rect 6114 36907 6148 36941
rect 6114 36839 6148 36873
rect 6114 36771 6148 36805
rect 6114 36703 6148 36737
rect 6114 36635 6148 36669
rect 6114 36567 6148 36601
rect 6114 36499 6148 36533
rect 6114 36431 6148 36465
rect 6114 36363 6148 36397
rect 6114 36295 6148 36329
rect 6114 36227 6148 36261
rect 6114 36159 6148 36193
rect 6114 36091 6148 36125
rect 6114 36023 6148 36057
rect 6114 35955 6148 35989
rect 6114 35887 6148 35921
rect 6114 35819 6148 35853
rect 6114 35751 6148 35785
rect 6114 35683 6148 35717
rect 6114 35615 6148 35649
rect 6114 35547 6148 35581
rect 6114 35479 6148 35513
rect 6114 35411 6148 35445
rect 6114 35343 6148 35377
rect 6114 35275 6148 35309
rect 6114 35207 6148 35241
rect 6114 35139 6148 35173
rect 6114 35071 6148 35105
rect 6114 35003 6148 35037
rect 6114 34935 6148 34969
rect 6114 34867 6148 34901
rect 6114 34799 6148 34833
rect 6114 34731 6148 34765
rect 6114 34663 6148 34697
rect 6114 34595 6148 34629
rect 6114 34527 6148 34561
rect 6114 34459 6148 34493
rect 6114 34391 6148 34425
rect 6114 34323 6148 34357
rect 6114 34255 6148 34289
rect 6114 34187 6148 34221
rect 6114 34119 6148 34153
rect 6114 34051 6148 34085
rect 6114 33983 6148 34017
rect 6114 33915 6148 33949
rect 6114 33847 6148 33881
rect 6114 33779 6148 33813
rect 6114 33711 6148 33745
rect 6114 33643 6148 33677
rect 6114 33575 6148 33609
rect 6114 33507 6148 33541
rect 6114 33439 6148 33473
rect 6114 33371 6148 33405
rect 6114 33303 6148 33337
rect 6114 33235 6148 33269
rect 6114 33167 6148 33201
rect 6114 33099 6148 33133
rect 6114 33031 6148 33065
rect 6114 32963 6148 32997
rect 6114 32895 6148 32929
rect 6114 32827 6148 32861
rect 6114 32759 6148 32793
rect 6114 32691 6148 32725
rect 6114 32623 6148 32657
rect 6114 32555 6148 32589
rect 6114 32487 6148 32521
rect 6114 32419 6148 32453
rect 6114 32351 6148 32385
rect 6114 32283 6148 32317
rect 6114 32215 6148 32249
rect 6114 32147 6148 32181
rect 6114 32079 6148 32113
rect 6114 32011 6148 32045
rect 6114 31943 6148 31977
rect 6114 31875 6148 31909
rect 6114 31807 6148 31841
rect 6114 31739 6148 31773
rect 6114 31671 6148 31705
rect 6114 31603 6148 31637
rect 6114 31535 6148 31569
rect 6114 31467 6148 31501
rect 6114 31399 6148 31433
rect 6114 31331 6148 31365
rect 6114 31263 6148 31297
rect 6114 31195 6148 31229
rect 6114 31127 6148 31161
rect 6114 31059 6148 31093
rect 6114 30991 6148 31025
rect 6114 30923 6148 30957
rect 6114 30855 6148 30889
rect 6114 30787 6148 30821
rect 6114 30719 6148 30753
rect 6114 30651 6148 30685
rect 6114 30583 6148 30617
rect 6114 30515 6148 30549
rect 6114 30447 6148 30481
rect 6114 30379 6148 30413
rect 6114 30311 6148 30345
rect 6114 30243 6148 30277
rect 6114 30175 6148 30209
rect 6114 30107 6148 30141
rect 6114 30039 6148 30073
rect 6114 29971 6148 30005
rect 6114 29903 6148 29937
rect 6114 29835 6148 29869
rect 6114 29767 6148 29801
rect 6114 29699 6148 29733
rect 6114 29631 6148 29665
rect 6114 29563 6148 29597
rect 6114 29495 6148 29529
rect 6114 29427 6148 29461
rect 6114 29359 6148 29393
rect 6114 29291 6148 29325
rect 6114 29223 6148 29257
rect 6114 29155 6148 29189
rect 6114 29087 6148 29121
rect 6114 29019 6148 29053
rect 6114 28951 6148 28985
rect 6114 28883 6148 28917
rect 6114 28815 6148 28849
rect 6114 28747 6148 28781
rect 6114 28679 6148 28713
rect 6114 28611 6148 28645
rect 6114 28543 6148 28577
rect 6114 28475 6148 28509
rect 6114 28407 6148 28441
rect 6114 28339 6148 28373
rect 6114 28271 6148 28305
rect 6114 28203 6148 28237
rect 6114 28135 6148 28169
rect 6114 28067 6148 28101
rect 6114 27999 6148 28033
rect 6114 27931 6148 27965
rect 6114 27863 6148 27897
rect 6114 27795 6148 27829
rect 6114 27727 6148 27761
rect 6114 27659 6148 27693
rect 6114 27591 6148 27625
rect 6114 27523 6148 27557
rect 6114 27455 6148 27489
rect 6114 27387 6148 27421
rect 6114 27319 6148 27353
rect 6114 27251 6148 27285
rect 6114 27183 6148 27217
rect 6114 27115 6148 27149
rect 6114 27047 6148 27081
rect 6114 26979 6148 27013
rect 6114 26911 6148 26945
rect 6114 26843 6148 26877
rect 6114 26775 6148 26809
rect 6114 26707 6148 26741
rect 6114 26639 6148 26673
rect 6114 26571 6148 26605
rect 6114 26503 6148 26537
rect 6114 26435 6148 26469
rect 6114 26367 6148 26401
rect 6114 26299 6148 26333
rect 6114 26231 6148 26265
rect 6114 26163 6148 26197
rect 6114 26095 6148 26129
rect 6114 26027 6148 26061
rect 6114 25959 6148 25993
rect 6114 25891 6148 25925
rect 6114 25823 6148 25857
rect 6114 25755 6148 25789
rect 6114 25687 6148 25721
rect 6114 25619 6148 25653
rect 6114 25551 6148 25585
rect 6114 25483 6148 25517
rect 6114 25415 6148 25449
rect 6114 25347 6148 25381
rect 6114 25279 6148 25313
rect 6114 25211 6148 25245
rect 6114 25143 6148 25177
rect 6114 25075 6148 25109
rect 6114 25007 6148 25041
rect 6114 24939 6148 24973
rect 6114 24871 6148 24905
rect 6114 24803 6148 24837
rect 6114 24735 6148 24769
rect 6114 24667 6148 24701
rect 6114 24599 6148 24633
rect 6114 24531 6148 24565
rect 6114 24463 6148 24497
rect 6114 24395 6148 24429
rect 6114 24327 6148 24361
rect 6114 24259 6148 24293
rect 6114 24191 6148 24225
rect 6114 24123 6148 24157
rect 6114 24055 6148 24089
rect 6114 23987 6148 24021
rect 6114 23919 6148 23953
rect 6114 23851 6148 23885
rect 6114 23783 6148 23817
rect 6114 23715 6148 23749
rect 6114 23647 6148 23681
rect 6114 23579 6148 23613
rect 6114 23511 6148 23545
rect 6114 23443 6148 23477
rect 6114 23375 6148 23409
rect 6114 23307 6148 23341
rect 6114 23239 6148 23273
rect 6114 23171 6148 23205
rect 6114 23103 6148 23137
rect 6114 23035 6148 23069
rect 6114 22967 6148 23001
rect 6114 22899 6148 22933
rect 6114 22831 6148 22865
rect 6114 22763 6148 22797
rect 6114 22695 6148 22729
rect 6114 22627 6148 22661
rect 6114 22559 6148 22593
rect 6114 22491 6148 22525
rect 6114 22423 6148 22457
rect 6114 22355 6148 22389
rect 6114 22287 6148 22321
rect 6114 22219 6148 22253
rect 6114 22151 6148 22185
rect 6114 22083 6148 22117
rect 6114 22015 6148 22049
rect 6114 21947 6148 21981
rect 6114 21879 6148 21913
rect 6114 21811 6148 21845
rect 6114 21743 6148 21777
rect 6114 21675 6148 21709
rect 6114 21607 6148 21641
rect 6114 21539 6148 21573
rect 6114 21471 6148 21505
rect 6114 21403 6148 21437
rect 6114 21335 6148 21369
rect 6114 21267 6148 21301
rect 6114 21199 6148 21233
rect 6114 21131 6148 21165
rect 6114 21063 6148 21097
rect 6114 20995 6148 21029
rect 6114 20927 6148 20961
rect 6114 20859 6148 20893
rect 6114 20791 6148 20825
rect 6114 20723 6148 20757
rect 6114 20655 6148 20689
rect 6114 20587 6148 20621
rect 6114 20519 6148 20553
rect 6114 20451 6148 20485
rect 6114 20383 6148 20417
rect 6114 20315 6148 20349
rect 6114 20247 6148 20281
rect 6114 20179 6148 20213
rect 6114 20111 6148 20145
rect 6114 20043 6148 20077
rect 6114 19975 6148 20009
rect 6114 19907 6148 19941
rect 6114 19839 6148 19873
rect 6114 19771 6148 19805
rect 6114 19703 6148 19737
rect 6114 19635 6148 19669
rect 6114 19567 6148 19601
rect 6114 19499 6148 19533
rect 6114 19431 6148 19465
rect 6114 19363 6148 19397
rect 6114 19295 6148 19329
rect 6114 19227 6148 19261
rect 6114 19159 6148 19193
rect 6114 19091 6148 19125
rect 6114 19023 6148 19057
rect 6114 18955 6148 18989
rect 6114 18887 6148 18921
rect 6114 18819 6148 18853
rect 6114 18751 6148 18785
rect 6114 18683 6148 18717
rect 6114 18615 6148 18649
rect 6114 18547 6148 18581
rect 6114 18479 6148 18513
rect 6114 18411 6148 18445
rect 6114 18343 6148 18377
rect 6114 18275 6148 18309
rect 6114 18207 6148 18241
rect 6114 18139 6148 18173
rect 6114 18071 6148 18105
rect 6114 18003 6148 18037
rect 6114 17935 6148 17969
rect 6114 17867 6148 17901
rect 6114 17799 6148 17833
rect 6114 17731 6148 17765
rect 6114 17663 6148 17697
rect 6114 17595 6148 17629
rect 6114 17527 6148 17561
rect 6114 17459 6148 17493
rect 6114 17391 6148 17425
rect 6114 17323 6148 17357
rect 6114 17255 6148 17289
rect 6114 17187 6148 17221
rect 6114 17119 6148 17153
rect 6114 17051 6148 17085
rect 6114 16983 6148 17017
rect 6114 16915 6148 16949
rect 6114 16847 6148 16881
rect 6114 16779 6148 16813
rect 6114 16711 6148 16745
rect 6114 16643 6148 16677
rect 6114 16575 6148 16609
rect 6114 16507 6148 16541
rect 6114 16439 6148 16473
rect 6114 16371 6148 16405
rect 6114 16303 6148 16337
rect 6114 16235 6148 16269
rect 6114 16167 6148 16201
rect 6114 16099 6148 16133
rect 6114 16031 6148 16065
rect 6114 15963 6148 15997
rect 6114 15895 6148 15929
rect 6114 15827 6148 15861
rect 6114 15759 6148 15793
rect 6114 15691 6148 15725
rect 6114 15623 6148 15657
rect 6114 15555 6148 15589
rect 6114 15487 6148 15521
rect 6114 15419 6148 15453
rect 6114 15351 6148 15385
rect 6114 15283 6148 15317
rect 6114 15215 6148 15249
rect 6114 15147 6148 15181
rect 6114 15079 6148 15113
rect 6114 15011 6148 15045
rect 6114 14943 6148 14977
rect 6114 14875 6148 14909
rect 6114 14807 6148 14841
rect 6114 14739 6148 14773
rect 6114 14671 6148 14705
rect 6114 14603 6148 14637
rect 6114 14535 6148 14569
rect 6114 14467 6148 14501
rect 6114 14399 6148 14433
rect 6114 14331 6148 14365
rect 6114 14263 6148 14297
rect 6114 14195 6148 14229
rect 6114 14127 6148 14161
rect 6114 14059 6148 14093
rect 6114 13991 6148 14025
rect 6114 13923 6148 13957
rect 6114 13855 6148 13889
rect 6114 13787 6148 13821
rect 6114 13719 6148 13753
rect 6114 13651 6148 13685
rect 6114 13583 6148 13617
rect 6114 13515 6148 13549
rect 6114 13447 6148 13481
rect 6114 13379 6148 13413
rect 6114 13311 6148 13345
rect 6114 13243 6148 13277
rect 6114 13175 6148 13209
rect 6114 13107 6148 13141
rect 6114 13039 6148 13073
rect 6114 12971 6148 13005
rect 6114 12903 6148 12937
rect 6114 12835 6148 12869
rect 6114 12767 6148 12801
rect 6114 12699 6148 12733
rect 6114 12631 6148 12665
rect 6114 12563 6148 12597
rect 6114 12495 6148 12529
rect 6114 12427 6148 12461
rect 6114 12359 6148 12393
rect 6114 12291 6148 12325
rect 6114 12223 6148 12257
rect 6114 12155 6148 12189
rect 6114 12087 6148 12121
rect 6114 12019 6148 12053
rect 6114 11951 6148 11985
rect 6114 11883 6148 11917
rect 6114 11815 6148 11849
rect 6114 11747 6148 11781
rect 6114 11679 6148 11713
rect 6114 11611 6148 11645
rect 6114 11543 6148 11577
rect 6114 11475 6148 11509
rect 6114 11407 6148 11441
rect 6114 11339 6148 11373
rect 6114 11271 6148 11305
rect 6114 11203 6148 11237
rect 6114 11135 6148 11169
rect 6114 11067 6148 11101
rect 6114 10999 6148 11033
rect 6114 10931 6148 10965
rect 6114 10863 6148 10897
rect 6114 10795 6148 10829
rect 6114 10727 6148 10761
rect 6114 10659 6148 10693
rect 6114 10591 6148 10625
rect 6114 10523 6148 10557
rect 6114 10455 6148 10489
rect 6114 10387 6148 10421
rect 6114 10319 6148 10353
rect 6114 10251 6148 10285
rect 6114 10183 6148 10217
rect 6114 10115 6148 10149
rect 6114 10047 6148 10081
rect 6114 9979 6148 10013
rect 6114 9911 6148 9945
rect 6114 9843 6148 9877
rect 6114 9775 6148 9809
rect 6114 9707 6148 9741
rect 6114 9639 6148 9673
rect 6114 9571 6148 9605
rect 6114 9503 6148 9537
rect 6114 9435 6148 9469
rect 6114 9367 6148 9401
rect 6114 9299 6148 9333
rect 6114 9231 6148 9265
rect 6114 9163 6148 9197
rect 6114 9095 6148 9129
rect 6114 9027 6148 9061
rect 6114 8959 6148 8993
rect 6114 8891 6148 8925
rect 6114 8823 6148 8857
rect 6114 8755 6148 8789
rect 6114 8687 6148 8721
rect 6114 8619 6148 8653
rect 6114 8551 6148 8585
rect 6114 8483 6148 8517
rect 6114 8415 6148 8449
rect 6114 8347 6148 8381
rect 6114 8279 6148 8313
rect 6114 8211 6148 8245
rect 6114 8143 6148 8177
rect 6114 8075 6148 8109
rect 6114 8007 6148 8041
rect 6114 7939 6148 7973
rect 6114 7871 6148 7905
rect 6114 7803 6148 7837
rect 6114 7735 6148 7769
rect 6114 7667 6148 7701
rect 6114 7599 6148 7633
rect 6114 7531 6148 7565
rect 6114 7463 6148 7497
rect 6114 7395 6148 7429
rect 6114 7327 6148 7361
rect 6114 7259 6148 7293
rect 6114 7191 6148 7225
rect 6114 7123 6148 7157
rect 6114 7055 6148 7089
rect 6114 6987 6148 7021
rect 6114 6919 6148 6953
rect 6114 6851 6148 6885
rect 6114 6783 6148 6817
rect 6114 6715 6148 6749
rect 6114 6647 6148 6681
rect 6114 6579 6148 6613
rect 6114 6511 6148 6545
rect 6114 6443 6148 6477
rect 6114 6375 6148 6409
rect 6114 6307 6148 6341
rect 6114 6239 6148 6273
rect 6114 6171 6148 6205
rect 6114 6103 6148 6137
rect 6114 6035 6148 6069
rect 6114 5967 6148 6001
rect 6114 5899 6148 5933
rect 6114 5831 6148 5865
rect 6114 5763 6148 5797
rect 6114 5695 6148 5729
rect 6114 5627 6148 5661
rect 6114 5559 6148 5593
rect 6114 5491 6148 5525
rect 6114 5423 6148 5457
rect 6114 5355 6148 5389
rect 6114 5287 6148 5321
rect 6114 5219 6148 5253
rect 6114 5151 6148 5185
rect 6114 5083 6148 5117
rect 6114 5015 6148 5049
rect 6114 4947 6148 4981
rect 6114 4879 6148 4913
rect 6114 4811 6148 4845
rect 6114 4743 6148 4777
rect 6114 4675 6148 4709
rect 6114 4607 6148 4641
rect 6114 4539 6148 4573
rect 6114 4471 6148 4505
rect 6114 4403 6148 4437
rect 6114 4335 6148 4369
rect 6114 4267 6148 4301
rect 6114 4199 6148 4233
rect 6114 4131 6148 4165
rect 6114 4063 6148 4097
rect 6114 3995 6148 4029
rect 6114 3927 6148 3961
rect 6114 3859 6148 3893
rect 6114 3791 6148 3825
rect 6114 3723 6148 3757
rect 6114 3655 6148 3689
rect 6114 3587 6148 3621
rect 6114 3519 6148 3553
rect 3972 3431 4006 3465
rect 3972 3363 4006 3397
rect 1830 3315 1864 3349
rect 1830 3247 1864 3281
rect 6114 3451 6148 3485
rect 6114 3383 6148 3417
rect 3972 3295 4006 3329
rect 6114 3315 6148 3349
rect 6114 3247 6148 3281
rect -184 3179 -150 3213
rect -116 3179 -82 3213
rect -48 3179 -14 3213
rect 20 3179 54 3213
rect 88 3179 122 3213
rect 156 3179 190 3213
rect 224 3179 258 3213
rect 292 3179 326 3213
rect 360 3179 394 3213
rect 428 3179 462 3213
rect 496 3179 530 3213
rect 564 3179 598 3213
rect 632 3179 666 3213
rect 700 3179 734 3213
rect 768 3179 802 3213
rect 836 3179 870 3213
rect 904 3179 938 3213
rect 972 3179 1006 3213
rect 1040 3179 1074 3213
rect 1108 3179 1142 3213
rect 1176 3179 1210 3213
rect 1244 3179 1278 3213
rect 1312 3179 1346 3213
rect 1380 3179 1414 3213
rect 1448 3179 1482 3213
rect 1516 3179 1550 3213
rect 1584 3179 1618 3213
rect 1652 3179 1686 3213
rect 1720 3179 1754 3213
rect 1932 3179 1966 3213
rect 2000 3179 2034 3213
rect 2068 3179 2102 3213
rect 2136 3179 2170 3213
rect 2204 3179 2238 3213
rect 2272 3179 2306 3213
rect 2340 3179 2374 3213
rect 2408 3179 2442 3213
rect 2476 3179 2510 3213
rect 2544 3179 2578 3213
rect 2612 3179 2646 3213
rect 2680 3179 2714 3213
rect 2748 3179 2782 3213
rect 2816 3179 2850 3213
rect 2884 3179 2918 3213
rect 2952 3179 2986 3213
rect 3020 3179 3054 3213
rect 3088 3179 3122 3213
rect 3156 3179 3190 3213
rect 3224 3179 3258 3213
rect 3292 3179 3326 3213
rect 3360 3179 3394 3213
rect 3428 3179 3462 3213
rect 3496 3179 3530 3213
rect 3564 3179 3598 3213
rect 3632 3179 3666 3213
rect 3700 3179 3734 3213
rect 3768 3179 3802 3213
rect 3836 3179 3870 3213
rect 3904 3179 3938 3213
rect 4040 3179 4074 3213
rect 4108 3179 4142 3213
rect 4176 3179 4210 3213
rect 4244 3179 4278 3213
rect 4312 3179 4346 3213
rect 4380 3179 4414 3213
rect 4448 3179 4482 3213
rect 4516 3179 4550 3213
rect 4584 3179 4618 3213
rect 4652 3179 4686 3213
rect 4720 3179 4754 3213
rect 4788 3179 4822 3213
rect 4856 3179 4890 3213
rect 4924 3179 4958 3213
rect 4992 3179 5026 3213
rect 5060 3179 5094 3213
rect 5128 3179 5162 3213
rect 5196 3179 5230 3213
rect 5264 3179 5298 3213
rect 5332 3179 5366 3213
rect 5400 3179 5434 3213
rect 5468 3179 5502 3213
rect 5536 3179 5570 3213
rect 5604 3179 5638 3213
rect 5672 3179 5706 3213
rect 5740 3179 5774 3213
rect 5808 3179 5842 3213
rect 5876 3179 5910 3213
rect 5944 3179 5978 3213
rect 6012 3179 6046 3213
rect 9206 38723 9240 38757
rect 9274 38723 9308 38757
rect 9342 38723 9376 38757
rect 9410 38723 9444 38757
rect 9478 38723 9512 38757
rect 9546 38723 9580 38757
rect 9614 38723 9648 38757
rect 9682 38723 9716 38757
rect 9750 38723 9784 38757
rect 9818 38723 9852 38757
rect 9886 38723 9920 38757
rect 9954 38723 9988 38757
rect 10022 38723 10056 38757
rect 10090 38723 10124 38757
rect 10158 38723 10192 38757
rect 10294 38723 10328 38757
rect 10362 38723 10396 38757
rect 10430 38723 10464 38757
rect 10498 38723 10532 38757
rect 10566 38723 10600 38757
rect 10634 38723 10668 38757
rect 10702 38723 10736 38757
rect 10770 38723 10804 38757
rect 10838 38723 10872 38757
rect 10906 38723 10940 38757
rect 10974 38723 11008 38757
rect 11042 38723 11076 38757
rect 11110 38723 11144 38757
rect 11178 38723 11212 38757
rect 11246 38723 11280 38757
rect 11314 38723 11348 38757
rect 11512 38723 11546 38757
rect 11580 38723 11614 38757
rect 11648 38723 11682 38757
rect 11716 38723 11750 38757
rect 11784 38723 11818 38757
rect 11852 38723 11886 38757
rect 11920 38723 11954 38757
rect 11988 38723 12022 38757
rect 12056 38723 12090 38757
rect 12124 38723 12158 38757
rect 12192 38723 12226 38757
rect 12260 38723 12294 38757
rect 12328 38723 12362 38757
rect 12396 38723 12430 38757
rect 12464 38723 12498 38757
rect 12532 38723 12566 38757
rect 12600 38723 12634 38757
rect 12668 38723 12702 38757
rect 12736 38723 12770 38757
rect 12804 38723 12838 38757
rect 12872 38723 12906 38757
rect 12940 38723 12974 38757
rect 13008 38723 13042 38757
rect 13076 38723 13110 38757
rect 13144 38723 13178 38757
rect 13280 38723 13314 38757
rect 13348 38723 13382 38757
rect 13416 38723 13450 38757
rect 13484 38723 13518 38757
rect 13552 38723 13586 38757
rect 13620 38723 13654 38757
rect 13688 38723 13722 38757
rect 13756 38723 13790 38757
rect 13824 38723 13858 38757
rect 13892 38723 13926 38757
rect 13960 38723 13994 38757
rect 14028 38723 14062 38757
rect 14096 38723 14130 38757
rect 14164 38723 14198 38757
rect 14232 38723 14266 38757
rect 14300 38723 14334 38757
rect 14368 38723 14402 38757
rect 14436 38723 14470 38757
rect 14504 38723 14538 38757
rect 14572 38723 14606 38757
rect 14640 38723 14674 38757
rect 14708 38723 14742 38757
rect 14776 38723 14810 38757
rect 14844 38723 14878 38757
rect 9088 38655 9122 38689
rect 9088 38587 9122 38621
rect 9088 38519 9122 38553
rect 9088 38451 9122 38485
rect 9088 38383 9122 38417
rect 9088 38315 9122 38349
rect 9088 38247 9122 38281
rect 9088 38179 9122 38213
rect 9088 38111 9122 38145
rect 9088 38043 9122 38077
rect 9088 37975 9122 38009
rect 9088 37907 9122 37941
rect 9088 37839 9122 37873
rect 9088 37771 9122 37805
rect 9088 37703 9122 37737
rect 9088 37635 9122 37669
rect 9088 37567 9122 37601
rect 9088 37499 9122 37533
rect 9088 37431 9122 37465
rect 9088 37363 9122 37397
rect 9088 37295 9122 37329
rect 9088 37227 9122 37261
rect 9088 37159 9122 37193
rect 9088 37091 9122 37125
rect 9088 37023 9122 37057
rect 9088 36955 9122 36989
rect 9088 36887 9122 36921
rect 9088 36819 9122 36853
rect 9088 36751 9122 36785
rect 9088 36683 9122 36717
rect 9088 36615 9122 36649
rect 9088 36547 9122 36581
rect 9088 36479 9122 36513
rect 9088 36411 9122 36445
rect 9088 36343 9122 36377
rect 9088 36275 9122 36309
rect 9088 36207 9122 36241
rect 9088 36139 9122 36173
rect 9088 36071 9122 36105
rect 9088 36003 9122 36037
rect 9088 35935 9122 35969
rect 9088 35867 9122 35901
rect 9088 35799 9122 35833
rect 9088 35731 9122 35765
rect 9088 35663 9122 35697
rect 9088 35595 9122 35629
rect 9088 35527 9122 35561
rect 9088 35459 9122 35493
rect 9088 35391 9122 35425
rect 9088 35323 9122 35357
rect 9088 35255 9122 35289
rect 9088 35187 9122 35221
rect 9088 35119 9122 35153
rect 9088 35051 9122 35085
rect 9088 34983 9122 35017
rect 9088 34915 9122 34949
rect 9088 34847 9122 34881
rect 9088 34779 9122 34813
rect 9088 34711 9122 34745
rect 9088 34643 9122 34677
rect 9088 34575 9122 34609
rect 9088 34507 9122 34541
rect 9088 34439 9122 34473
rect 9088 34371 9122 34405
rect 9088 34303 9122 34337
rect 9088 34235 9122 34269
rect 9088 34167 9122 34201
rect 9088 34099 9122 34133
rect 9088 34031 9122 34065
rect 9088 33963 9122 33997
rect 9088 33895 9122 33929
rect 9088 33827 9122 33861
rect 9088 33759 9122 33793
rect 9088 33691 9122 33725
rect 9088 33623 9122 33657
rect 9088 33555 9122 33589
rect 9088 33487 9122 33521
rect 9088 33419 9122 33453
rect 9088 33351 9122 33385
rect 9088 33283 9122 33317
rect 9088 33215 9122 33249
rect 9088 33147 9122 33181
rect 9088 33079 9122 33113
rect 9088 33011 9122 33045
rect 9088 32943 9122 32977
rect 9088 32875 9122 32909
rect 9088 32807 9122 32841
rect 9088 32739 9122 32773
rect 9088 32671 9122 32705
rect 9088 32603 9122 32637
rect 9088 32535 9122 32569
rect 9088 32467 9122 32501
rect 9088 32399 9122 32433
rect 9088 32331 9122 32365
rect 9088 32263 9122 32297
rect 9088 32195 9122 32229
rect 9088 32127 9122 32161
rect 9088 32059 9122 32093
rect 9088 31991 9122 32025
rect 9088 31923 9122 31957
rect 9088 31855 9122 31889
rect 9088 31787 9122 31821
rect 9088 31719 9122 31753
rect 9088 31651 9122 31685
rect 9088 31583 9122 31617
rect 9088 31515 9122 31549
rect 9088 31447 9122 31481
rect 9088 31379 9122 31413
rect 9088 31311 9122 31345
rect 9088 31243 9122 31277
rect 9088 31175 9122 31209
rect 9088 31107 9122 31141
rect 9088 31039 9122 31073
rect 9088 30971 9122 31005
rect 9088 30903 9122 30937
rect 9088 30835 9122 30869
rect 9088 30767 9122 30801
rect 9088 30699 9122 30733
rect 9088 30631 9122 30665
rect 9088 30563 9122 30597
rect 9088 30495 9122 30529
rect 9088 30427 9122 30461
rect 9088 30359 9122 30393
rect 9088 30291 9122 30325
rect 9088 30223 9122 30257
rect 9088 30155 9122 30189
rect 9088 30087 9122 30121
rect 9088 30019 9122 30053
rect 9088 29951 9122 29985
rect 9088 29883 9122 29917
rect 9088 29815 9122 29849
rect 9088 29747 9122 29781
rect 9088 29679 9122 29713
rect 9088 29611 9122 29645
rect 9088 29543 9122 29577
rect 9088 29475 9122 29509
rect 9088 29407 9122 29441
rect 9088 29339 9122 29373
rect 9088 29271 9122 29305
rect 9088 29203 9122 29237
rect 9088 29135 9122 29169
rect 9088 29067 9122 29101
rect 9088 28999 9122 29033
rect 9088 28931 9122 28965
rect 9088 28863 9122 28897
rect 9088 28795 9122 28829
rect 9088 28727 9122 28761
rect 9088 28659 9122 28693
rect 9088 28591 9122 28625
rect 9088 28523 9122 28557
rect 9088 28455 9122 28489
rect 9088 28387 9122 28421
rect 9088 28319 9122 28353
rect 9088 28251 9122 28285
rect 9088 28183 9122 28217
rect 9088 28115 9122 28149
rect 9088 28047 9122 28081
rect 9088 27979 9122 28013
rect 9088 27911 9122 27945
rect 9088 27843 9122 27877
rect 9088 27775 9122 27809
rect 9088 27707 9122 27741
rect 9088 27639 9122 27673
rect 9088 27571 9122 27605
rect 9088 27503 9122 27537
rect 9088 27435 9122 27469
rect 9088 27367 9122 27401
rect 9088 27299 9122 27333
rect 9088 27231 9122 27265
rect 9088 27163 9122 27197
rect 9088 27095 9122 27129
rect 9088 27027 9122 27061
rect 9088 26959 9122 26993
rect 9088 26891 9122 26925
rect 9088 26823 9122 26857
rect 9088 26755 9122 26789
rect 9088 26687 9122 26721
rect 9088 26619 9122 26653
rect 9088 26551 9122 26585
rect 9088 26483 9122 26517
rect 9088 26415 9122 26449
rect 9088 26347 9122 26381
rect 9088 26279 9122 26313
rect 9088 26211 9122 26245
rect 9088 26143 9122 26177
rect 9088 26075 9122 26109
rect 9088 26007 9122 26041
rect 9088 25939 9122 25973
rect 9088 25871 9122 25905
rect 9088 25803 9122 25837
rect 9088 25735 9122 25769
rect 9088 25667 9122 25701
rect 9088 25599 9122 25633
rect 9088 25531 9122 25565
rect 9088 25463 9122 25497
rect 9088 25395 9122 25429
rect 9088 25327 9122 25361
rect 9088 25259 9122 25293
rect 9088 25191 9122 25225
rect 9088 25123 9122 25157
rect 9088 25055 9122 25089
rect 9088 24987 9122 25021
rect 9088 24919 9122 24953
rect 9088 24851 9122 24885
rect 9088 24783 9122 24817
rect 9088 24715 9122 24749
rect 9088 24647 9122 24681
rect 9088 24579 9122 24613
rect 9088 24511 9122 24545
rect 9088 24443 9122 24477
rect 9088 24375 9122 24409
rect 9088 24307 9122 24341
rect 9088 24239 9122 24273
rect 9088 24171 9122 24205
rect 9088 24103 9122 24137
rect 9088 24035 9122 24069
rect 9088 23967 9122 24001
rect 9088 23899 9122 23933
rect 9088 23831 9122 23865
rect 9088 23763 9122 23797
rect 9088 23695 9122 23729
rect 9088 23627 9122 23661
rect 9088 23559 9122 23593
rect 9088 23491 9122 23525
rect 9088 23423 9122 23457
rect 9088 23355 9122 23389
rect 9088 23287 9122 23321
rect 9088 23219 9122 23253
rect 9088 23151 9122 23185
rect 9088 23083 9122 23117
rect 9088 23015 9122 23049
rect 9088 22947 9122 22981
rect 9088 22879 9122 22913
rect 9088 22811 9122 22845
rect 9088 22743 9122 22777
rect 9088 22675 9122 22709
rect 9088 22607 9122 22641
rect 9088 22539 9122 22573
rect 9088 22471 9122 22505
rect 9088 22403 9122 22437
rect 9088 22335 9122 22369
rect 9088 22267 9122 22301
rect 9088 22199 9122 22233
rect 9088 22131 9122 22165
rect 9088 22063 9122 22097
rect 9088 21995 9122 22029
rect 9088 21927 9122 21961
rect 9088 21859 9122 21893
rect 9088 21791 9122 21825
rect 9088 21723 9122 21757
rect 9088 21655 9122 21689
rect 9088 21587 9122 21621
rect 9088 21519 9122 21553
rect 9088 21451 9122 21485
rect 9088 21383 9122 21417
rect 9088 21315 9122 21349
rect 9088 21247 9122 21281
rect 9088 21179 9122 21213
rect 9088 21111 9122 21145
rect 9088 21043 9122 21077
rect 9088 20975 9122 21009
rect 9088 20907 9122 20941
rect 9088 20839 9122 20873
rect 9088 20771 9122 20805
rect 9088 20703 9122 20737
rect 9088 20635 9122 20669
rect 9088 20567 9122 20601
rect 9088 20499 9122 20533
rect 9088 20431 9122 20465
rect 9088 20363 9122 20397
rect 9088 20295 9122 20329
rect 9088 20227 9122 20261
rect 9088 20159 9122 20193
rect 9088 20091 9122 20125
rect 9088 20023 9122 20057
rect 9088 19955 9122 19989
rect 9088 19887 9122 19921
rect 9088 19819 9122 19853
rect 9088 19751 9122 19785
rect 9088 19683 9122 19717
rect 9088 19615 9122 19649
rect 9088 19547 9122 19581
rect 9088 19479 9122 19513
rect 9088 19411 9122 19445
rect 9088 19343 9122 19377
rect 9088 19275 9122 19309
rect 9088 19207 9122 19241
rect 9088 19139 9122 19173
rect 9088 19071 9122 19105
rect 9088 19003 9122 19037
rect 9088 18935 9122 18969
rect 9088 18867 9122 18901
rect 9088 18799 9122 18833
rect 9088 18731 9122 18765
rect 9088 18663 9122 18697
rect 9088 18595 9122 18629
rect 9088 18527 9122 18561
rect 9088 18459 9122 18493
rect 9088 18391 9122 18425
rect 9088 18323 9122 18357
rect 9088 18255 9122 18289
rect 9088 18187 9122 18221
rect 9088 18119 9122 18153
rect 9088 18051 9122 18085
rect 9088 17983 9122 18017
rect 9088 17915 9122 17949
rect 9088 17847 9122 17881
rect 9088 17779 9122 17813
rect 9088 17711 9122 17745
rect 9088 17643 9122 17677
rect 9088 17575 9122 17609
rect 9088 17507 9122 17541
rect 9088 17439 9122 17473
rect 9088 17371 9122 17405
rect 9088 17303 9122 17337
rect 9088 17235 9122 17269
rect 9088 17167 9122 17201
rect 9088 17099 9122 17133
rect 9088 17031 9122 17065
rect 9088 16963 9122 16997
rect 9088 16895 9122 16929
rect 9088 16827 9122 16861
rect 9088 16759 9122 16793
rect 9088 16691 9122 16725
rect 9088 16623 9122 16657
rect 9088 16555 9122 16589
rect 9088 16487 9122 16521
rect 9088 16419 9122 16453
rect 9088 16351 9122 16385
rect 9088 16283 9122 16317
rect 9088 16215 9122 16249
rect 9088 16147 9122 16181
rect 9088 16079 9122 16113
rect 9088 16011 9122 16045
rect 9088 15943 9122 15977
rect 9088 15875 9122 15909
rect 9088 15807 9122 15841
rect 9088 15739 9122 15773
rect 9088 15671 9122 15705
rect 9088 15603 9122 15637
rect 9088 15535 9122 15569
rect 9088 15467 9122 15501
rect 9088 15399 9122 15433
rect 9088 15331 9122 15365
rect 9088 15263 9122 15297
rect 9088 15195 9122 15229
rect 9088 15127 9122 15161
rect 9088 15059 9122 15093
rect 9088 14991 9122 15025
rect 9088 14923 9122 14957
rect 9088 14855 9122 14889
rect 9088 14787 9122 14821
rect 9088 14719 9122 14753
rect 9088 14651 9122 14685
rect 9088 14583 9122 14617
rect 9088 14515 9122 14549
rect 9088 14447 9122 14481
rect 9088 14379 9122 14413
rect 9088 14311 9122 14345
rect 9088 14243 9122 14277
rect 9088 14175 9122 14209
rect 9088 14107 9122 14141
rect 9088 14039 9122 14073
rect 9088 13971 9122 14005
rect 9088 13903 9122 13937
rect 9088 13835 9122 13869
rect 9088 13767 9122 13801
rect 9088 13699 9122 13733
rect 9088 13631 9122 13665
rect 9088 13563 9122 13597
rect 9088 13495 9122 13529
rect 9088 13427 9122 13461
rect 9088 13359 9122 13393
rect 9088 13291 9122 13325
rect 9088 13223 9122 13257
rect 9088 13155 9122 13189
rect 9088 13087 9122 13121
rect 9088 13019 9122 13053
rect 9088 12951 9122 12985
rect 9088 12883 9122 12917
rect 9088 12815 9122 12849
rect 9088 12747 9122 12781
rect 9088 12679 9122 12713
rect 9088 12611 9122 12645
rect 9088 12543 9122 12577
rect 9088 12475 9122 12509
rect 9088 12407 9122 12441
rect 9088 12339 9122 12373
rect 9088 12271 9122 12305
rect 9088 12203 9122 12237
rect 9088 12135 9122 12169
rect 9088 12067 9122 12101
rect 9088 11999 9122 12033
rect 9088 11931 9122 11965
rect 9088 11863 9122 11897
rect 9088 11795 9122 11829
rect 9088 11727 9122 11761
rect 9088 11659 9122 11693
rect 9088 11591 9122 11625
rect 9088 11523 9122 11557
rect 9088 11455 9122 11489
rect 9088 11387 9122 11421
rect 9088 11319 9122 11353
rect 9088 11251 9122 11285
rect 9088 11183 9122 11217
rect 9088 11115 9122 11149
rect 9088 11047 9122 11081
rect 9088 10979 9122 11013
rect 9088 10911 9122 10945
rect 9088 10843 9122 10877
rect 9088 10775 9122 10809
rect 9088 10707 9122 10741
rect 9088 10639 9122 10673
rect 9088 10571 9122 10605
rect 9088 10503 9122 10537
rect 9088 10435 9122 10469
rect 9088 10367 9122 10401
rect 9088 10299 9122 10333
rect 9088 10231 9122 10265
rect 9088 10163 9122 10197
rect 9088 10095 9122 10129
rect 9088 10027 9122 10061
rect 9088 9959 9122 9993
rect 9088 9891 9122 9925
rect 9088 9823 9122 9857
rect 9088 9755 9122 9789
rect 9088 9687 9122 9721
rect 9088 9619 9122 9653
rect 9088 9551 9122 9585
rect 9088 9483 9122 9517
rect 9088 9415 9122 9449
rect 9088 9347 9122 9381
rect 9088 9279 9122 9313
rect 9088 9211 9122 9245
rect 9088 9143 9122 9177
rect 9088 9075 9122 9109
rect 9088 9007 9122 9041
rect 9088 8939 9122 8973
rect 9088 8871 9122 8905
rect 9088 8803 9122 8837
rect 9088 8735 9122 8769
rect 9088 8667 9122 8701
rect 9088 8599 9122 8633
rect 9088 8531 9122 8565
rect 9088 8463 9122 8497
rect 9088 8395 9122 8429
rect 9088 8327 9122 8361
rect 9088 8259 9122 8293
rect 9088 8191 9122 8225
rect 9088 8123 9122 8157
rect 9088 8055 9122 8089
rect 9088 7987 9122 8021
rect 9088 7919 9122 7953
rect 9088 7851 9122 7885
rect 9088 7783 9122 7817
rect 9088 7715 9122 7749
rect 9088 7647 9122 7681
rect 9088 7579 9122 7613
rect 9088 7511 9122 7545
rect 9088 7443 9122 7477
rect 9088 7375 9122 7409
rect 9088 7307 9122 7341
rect 9088 7239 9122 7273
rect 9088 7171 9122 7205
rect 9088 7103 9122 7137
rect 9088 7035 9122 7069
rect 9088 6967 9122 7001
rect 9088 6899 9122 6933
rect 9088 6831 9122 6865
rect 9088 6763 9122 6797
rect 9088 6695 9122 6729
rect 9088 6627 9122 6661
rect 9088 6559 9122 6593
rect 9088 6491 9122 6525
rect 9088 6423 9122 6457
rect 9088 6355 9122 6389
rect 9088 6287 9122 6321
rect 9088 6219 9122 6253
rect 9088 6151 9122 6185
rect 9088 6083 9122 6117
rect 9088 6015 9122 6049
rect 9088 5947 9122 5981
rect 9088 5879 9122 5913
rect 9088 5811 9122 5845
rect 9088 5743 9122 5777
rect 9088 5675 9122 5709
rect 9088 5607 9122 5641
rect 9088 5539 9122 5573
rect 9088 5471 9122 5505
rect 9088 5403 9122 5437
rect 9088 5335 9122 5369
rect 9088 5267 9122 5301
rect 9088 5199 9122 5233
rect 9088 5131 9122 5165
rect 9088 5063 9122 5097
rect 9088 4995 9122 5029
rect 9088 4927 9122 4961
rect 9088 4859 9122 4893
rect 9088 4791 9122 4825
rect 9088 4723 9122 4757
rect 9088 4655 9122 4689
rect 9088 4587 9122 4621
rect 9088 4519 9122 4553
rect 9088 4451 9122 4485
rect 9088 4383 9122 4417
rect 9088 4315 9122 4349
rect 9088 4247 9122 4281
rect 9088 4179 9122 4213
rect 9088 4111 9122 4145
rect 9088 4043 9122 4077
rect 9088 3975 9122 4009
rect 9088 3907 9122 3941
rect 9088 3839 9122 3873
rect 9088 3771 9122 3805
rect 9088 3703 9122 3737
rect 9088 3635 9122 3669
rect 9088 3567 9122 3601
rect 9088 3499 9122 3533
rect 10226 38607 10260 38641
rect 10226 38539 10260 38573
rect 10226 38471 10260 38505
rect 10226 38403 10260 38437
rect 10226 38335 10260 38369
rect 10226 38267 10260 38301
rect 10226 38199 10260 38233
rect 10226 38131 10260 38165
rect 10226 38063 10260 38097
rect 10226 37995 10260 38029
rect 10226 37927 10260 37961
rect 10226 37859 10260 37893
rect 10226 37791 10260 37825
rect 10226 37723 10260 37757
rect 10226 37655 10260 37689
rect 10226 37587 10260 37621
rect 10226 37519 10260 37553
rect 10226 37451 10260 37485
rect 10226 37383 10260 37417
rect 10226 37315 10260 37349
rect 10226 37247 10260 37281
rect 10226 37179 10260 37213
rect 10226 37111 10260 37145
rect 10226 37043 10260 37077
rect 10226 36975 10260 37009
rect 10226 36907 10260 36941
rect 10226 36839 10260 36873
rect 10226 36771 10260 36805
rect 10226 36703 10260 36737
rect 10226 36635 10260 36669
rect 10226 36567 10260 36601
rect 10226 36499 10260 36533
rect 10226 36431 10260 36465
rect 10226 36363 10260 36397
rect 10226 36295 10260 36329
rect 10226 36227 10260 36261
rect 10226 36159 10260 36193
rect 10226 36091 10260 36125
rect 10226 36023 10260 36057
rect 10226 35955 10260 35989
rect 10226 35887 10260 35921
rect 10226 35819 10260 35853
rect 10226 35751 10260 35785
rect 10226 35683 10260 35717
rect 10226 35615 10260 35649
rect 10226 35547 10260 35581
rect 10226 35479 10260 35513
rect 10226 35411 10260 35445
rect 10226 35343 10260 35377
rect 10226 35275 10260 35309
rect 10226 35207 10260 35241
rect 10226 35139 10260 35173
rect 10226 35071 10260 35105
rect 10226 35003 10260 35037
rect 10226 34935 10260 34969
rect 10226 34867 10260 34901
rect 10226 34799 10260 34833
rect 10226 34731 10260 34765
rect 10226 34663 10260 34697
rect 10226 34595 10260 34629
rect 10226 34527 10260 34561
rect 10226 34459 10260 34493
rect 10226 34391 10260 34425
rect 10226 34323 10260 34357
rect 10226 34255 10260 34289
rect 10226 34187 10260 34221
rect 10226 34119 10260 34153
rect 10226 34051 10260 34085
rect 10226 33983 10260 34017
rect 10226 33915 10260 33949
rect 10226 33847 10260 33881
rect 10226 33779 10260 33813
rect 10226 33711 10260 33745
rect 10226 33643 10260 33677
rect 10226 33575 10260 33609
rect 10226 33507 10260 33541
rect 10226 33439 10260 33473
rect 10226 33371 10260 33405
rect 10226 33303 10260 33337
rect 10226 33235 10260 33269
rect 10226 33167 10260 33201
rect 10226 33099 10260 33133
rect 10226 33031 10260 33065
rect 10226 32963 10260 32997
rect 10226 32895 10260 32929
rect 10226 32827 10260 32861
rect 10226 32759 10260 32793
rect 10226 32691 10260 32725
rect 10226 32623 10260 32657
rect 10226 32555 10260 32589
rect 10226 32487 10260 32521
rect 10226 32419 10260 32453
rect 10226 32351 10260 32385
rect 10226 32283 10260 32317
rect 10226 32215 10260 32249
rect 10226 32147 10260 32181
rect 10226 32079 10260 32113
rect 10226 32011 10260 32045
rect 10226 31943 10260 31977
rect 10226 31875 10260 31909
rect 10226 31807 10260 31841
rect 10226 31739 10260 31773
rect 10226 31671 10260 31705
rect 10226 31603 10260 31637
rect 10226 31535 10260 31569
rect 10226 31467 10260 31501
rect 10226 31399 10260 31433
rect 10226 31331 10260 31365
rect 10226 31263 10260 31297
rect 10226 31195 10260 31229
rect 10226 31127 10260 31161
rect 10226 31059 10260 31093
rect 10226 30991 10260 31025
rect 10226 30923 10260 30957
rect 10226 30855 10260 30889
rect 10226 30787 10260 30821
rect 10226 30719 10260 30753
rect 10226 30651 10260 30685
rect 10226 30583 10260 30617
rect 10226 30515 10260 30549
rect 10226 30447 10260 30481
rect 10226 30379 10260 30413
rect 10226 30311 10260 30345
rect 10226 30243 10260 30277
rect 10226 30175 10260 30209
rect 10226 30107 10260 30141
rect 10226 30039 10260 30073
rect 10226 29971 10260 30005
rect 10226 29903 10260 29937
rect 10226 29835 10260 29869
rect 10226 29767 10260 29801
rect 10226 29699 10260 29733
rect 10226 29631 10260 29665
rect 10226 29563 10260 29597
rect 10226 29495 10260 29529
rect 10226 29427 10260 29461
rect 10226 29359 10260 29393
rect 10226 29291 10260 29325
rect 10226 29223 10260 29257
rect 10226 29155 10260 29189
rect 10226 29087 10260 29121
rect 10226 29019 10260 29053
rect 10226 28951 10260 28985
rect 10226 28883 10260 28917
rect 10226 28815 10260 28849
rect 10226 28747 10260 28781
rect 10226 28679 10260 28713
rect 10226 28611 10260 28645
rect 10226 28543 10260 28577
rect 10226 28475 10260 28509
rect 10226 28407 10260 28441
rect 10226 28339 10260 28373
rect 10226 28271 10260 28305
rect 10226 28203 10260 28237
rect 10226 28135 10260 28169
rect 10226 28067 10260 28101
rect 10226 27999 10260 28033
rect 10226 27931 10260 27965
rect 10226 27863 10260 27897
rect 10226 27795 10260 27829
rect 10226 27727 10260 27761
rect 10226 27659 10260 27693
rect 10226 27591 10260 27625
rect 10226 27523 10260 27557
rect 10226 27455 10260 27489
rect 10226 27387 10260 27421
rect 10226 27319 10260 27353
rect 10226 27251 10260 27285
rect 10226 27183 10260 27217
rect 10226 27115 10260 27149
rect 10226 27047 10260 27081
rect 10226 26979 10260 27013
rect 10226 26911 10260 26945
rect 10226 26843 10260 26877
rect 10226 26775 10260 26809
rect 10226 26707 10260 26741
rect 10226 26639 10260 26673
rect 10226 26571 10260 26605
rect 10226 26503 10260 26537
rect 10226 26435 10260 26469
rect 10226 26367 10260 26401
rect 10226 26299 10260 26333
rect 10226 26231 10260 26265
rect 10226 26163 10260 26197
rect 10226 26095 10260 26129
rect 10226 26027 10260 26061
rect 10226 25959 10260 25993
rect 10226 25891 10260 25925
rect 10226 25823 10260 25857
rect 10226 25755 10260 25789
rect 10226 25687 10260 25721
rect 10226 25619 10260 25653
rect 10226 25551 10260 25585
rect 10226 25483 10260 25517
rect 10226 25415 10260 25449
rect 10226 25347 10260 25381
rect 10226 25279 10260 25313
rect 10226 25211 10260 25245
rect 10226 25143 10260 25177
rect 10226 25075 10260 25109
rect 10226 25007 10260 25041
rect 10226 24939 10260 24973
rect 10226 24871 10260 24905
rect 10226 24803 10260 24837
rect 10226 24735 10260 24769
rect 10226 24667 10260 24701
rect 10226 24599 10260 24633
rect 10226 24531 10260 24565
rect 10226 24463 10260 24497
rect 10226 24395 10260 24429
rect 10226 24327 10260 24361
rect 10226 24259 10260 24293
rect 10226 24191 10260 24225
rect 10226 24123 10260 24157
rect 10226 24055 10260 24089
rect 10226 23987 10260 24021
rect 10226 23919 10260 23953
rect 10226 23851 10260 23885
rect 10226 23783 10260 23817
rect 10226 23715 10260 23749
rect 10226 23647 10260 23681
rect 10226 23579 10260 23613
rect 10226 23511 10260 23545
rect 10226 23443 10260 23477
rect 10226 23375 10260 23409
rect 10226 23307 10260 23341
rect 10226 23239 10260 23273
rect 10226 23171 10260 23205
rect 10226 23103 10260 23137
rect 10226 23035 10260 23069
rect 10226 22967 10260 23001
rect 10226 22899 10260 22933
rect 10226 22831 10260 22865
rect 10226 22763 10260 22797
rect 10226 22695 10260 22729
rect 10226 22627 10260 22661
rect 10226 22559 10260 22593
rect 10226 22491 10260 22525
rect 10226 22423 10260 22457
rect 10226 22355 10260 22389
rect 10226 22287 10260 22321
rect 10226 22219 10260 22253
rect 10226 22151 10260 22185
rect 10226 22083 10260 22117
rect 10226 22015 10260 22049
rect 10226 21947 10260 21981
rect 10226 21879 10260 21913
rect 10226 21811 10260 21845
rect 10226 21743 10260 21777
rect 10226 21675 10260 21709
rect 10226 21607 10260 21641
rect 10226 21539 10260 21573
rect 10226 21471 10260 21505
rect 10226 21403 10260 21437
rect 10226 21335 10260 21369
rect 10226 21267 10260 21301
rect 10226 21199 10260 21233
rect 10226 21131 10260 21165
rect 10226 21063 10260 21097
rect 10226 20995 10260 21029
rect 10226 20927 10260 20961
rect 10226 20859 10260 20893
rect 10226 20791 10260 20825
rect 10226 20723 10260 20757
rect 10226 20655 10260 20689
rect 10226 20587 10260 20621
rect 10226 20519 10260 20553
rect 10226 20451 10260 20485
rect 10226 20383 10260 20417
rect 10226 20315 10260 20349
rect 10226 20247 10260 20281
rect 10226 20179 10260 20213
rect 10226 20111 10260 20145
rect 10226 20043 10260 20077
rect 10226 19975 10260 20009
rect 10226 19907 10260 19941
rect 10226 19839 10260 19873
rect 10226 19771 10260 19805
rect 10226 19703 10260 19737
rect 10226 19635 10260 19669
rect 10226 19567 10260 19601
rect 10226 19499 10260 19533
rect 10226 19431 10260 19465
rect 10226 19363 10260 19397
rect 10226 19295 10260 19329
rect 10226 19227 10260 19261
rect 10226 19159 10260 19193
rect 10226 19091 10260 19125
rect 10226 19023 10260 19057
rect 10226 18955 10260 18989
rect 10226 18887 10260 18921
rect 10226 18819 10260 18853
rect 10226 18751 10260 18785
rect 10226 18683 10260 18717
rect 10226 18615 10260 18649
rect 10226 18547 10260 18581
rect 10226 18479 10260 18513
rect 10226 18411 10260 18445
rect 10226 18343 10260 18377
rect 10226 18275 10260 18309
rect 10226 18207 10260 18241
rect 10226 18139 10260 18173
rect 10226 18071 10260 18105
rect 10226 18003 10260 18037
rect 10226 17935 10260 17969
rect 10226 17867 10260 17901
rect 10226 17799 10260 17833
rect 10226 17731 10260 17765
rect 10226 17663 10260 17697
rect 10226 17595 10260 17629
rect 10226 17527 10260 17561
rect 10226 17459 10260 17493
rect 10226 17391 10260 17425
rect 10226 17323 10260 17357
rect 10226 17255 10260 17289
rect 10226 17187 10260 17221
rect 10226 17119 10260 17153
rect 10226 17051 10260 17085
rect 10226 16983 10260 17017
rect 10226 16915 10260 16949
rect 10226 16847 10260 16881
rect 10226 16779 10260 16813
rect 10226 16711 10260 16745
rect 10226 16643 10260 16677
rect 10226 16575 10260 16609
rect 10226 16507 10260 16541
rect 10226 16439 10260 16473
rect 10226 16371 10260 16405
rect 10226 16303 10260 16337
rect 10226 16235 10260 16269
rect 10226 16167 10260 16201
rect 10226 16099 10260 16133
rect 10226 16031 10260 16065
rect 10226 15963 10260 15997
rect 10226 15895 10260 15929
rect 10226 15827 10260 15861
rect 10226 15759 10260 15793
rect 10226 15691 10260 15725
rect 10226 15623 10260 15657
rect 10226 15555 10260 15589
rect 10226 15487 10260 15521
rect 10226 15419 10260 15453
rect 10226 15351 10260 15385
rect 10226 15283 10260 15317
rect 10226 15215 10260 15249
rect 10226 15147 10260 15181
rect 10226 15079 10260 15113
rect 10226 15011 10260 15045
rect 10226 14943 10260 14977
rect 10226 14875 10260 14909
rect 10226 14807 10260 14841
rect 10226 14739 10260 14773
rect 10226 14671 10260 14705
rect 10226 14603 10260 14637
rect 10226 14535 10260 14569
rect 10226 14467 10260 14501
rect 10226 14399 10260 14433
rect 10226 14331 10260 14365
rect 10226 14263 10260 14297
rect 10226 14195 10260 14229
rect 10226 14127 10260 14161
rect 10226 14059 10260 14093
rect 10226 13991 10260 14025
rect 10226 13923 10260 13957
rect 10226 13855 10260 13889
rect 10226 13787 10260 13821
rect 10226 13719 10260 13753
rect 10226 13651 10260 13685
rect 10226 13583 10260 13617
rect 10226 13515 10260 13549
rect 10226 13447 10260 13481
rect 10226 13379 10260 13413
rect 10226 13311 10260 13345
rect 10226 13243 10260 13277
rect 10226 13175 10260 13209
rect 10226 13107 10260 13141
rect 10226 13039 10260 13073
rect 10226 12971 10260 13005
rect 10226 12903 10260 12937
rect 10226 12835 10260 12869
rect 10226 12767 10260 12801
rect 10226 12699 10260 12733
rect 10226 12631 10260 12665
rect 10226 12563 10260 12597
rect 10226 12495 10260 12529
rect 10226 12427 10260 12461
rect 10226 12359 10260 12393
rect 10226 12291 10260 12325
rect 10226 12223 10260 12257
rect 10226 12155 10260 12189
rect 10226 12087 10260 12121
rect 10226 12019 10260 12053
rect 10226 11951 10260 11985
rect 10226 11883 10260 11917
rect 10226 11815 10260 11849
rect 10226 11747 10260 11781
rect 10226 11679 10260 11713
rect 10226 11611 10260 11645
rect 10226 11543 10260 11577
rect 10226 11475 10260 11509
rect 10226 11407 10260 11441
rect 10226 11339 10260 11373
rect 10226 11271 10260 11305
rect 10226 11203 10260 11237
rect 10226 11135 10260 11169
rect 10226 11067 10260 11101
rect 10226 10999 10260 11033
rect 10226 10931 10260 10965
rect 10226 10863 10260 10897
rect 10226 10795 10260 10829
rect 10226 10727 10260 10761
rect 10226 10659 10260 10693
rect 10226 10591 10260 10625
rect 10226 10523 10260 10557
rect 10226 10455 10260 10489
rect 10226 10387 10260 10421
rect 10226 10319 10260 10353
rect 10226 10251 10260 10285
rect 10226 10183 10260 10217
rect 10226 10115 10260 10149
rect 10226 10047 10260 10081
rect 10226 9979 10260 10013
rect 10226 9911 10260 9945
rect 10226 9843 10260 9877
rect 10226 9775 10260 9809
rect 10226 9707 10260 9741
rect 10226 9639 10260 9673
rect 10226 9571 10260 9605
rect 10226 9503 10260 9537
rect 10226 9435 10260 9469
rect 10226 9367 10260 9401
rect 10226 9299 10260 9333
rect 10226 9231 10260 9265
rect 10226 9163 10260 9197
rect 10226 9095 10260 9129
rect 10226 9027 10260 9061
rect 10226 8959 10260 8993
rect 10226 8891 10260 8925
rect 10226 8823 10260 8857
rect 10226 8755 10260 8789
rect 10226 8687 10260 8721
rect 10226 8619 10260 8653
rect 10226 8551 10260 8585
rect 10226 8483 10260 8517
rect 10226 8415 10260 8449
rect 10226 8347 10260 8381
rect 10226 8279 10260 8313
rect 10226 8211 10260 8245
rect 10226 8143 10260 8177
rect 10226 8075 10260 8109
rect 10226 8007 10260 8041
rect 10226 7939 10260 7973
rect 10226 7871 10260 7905
rect 10226 7803 10260 7837
rect 10226 7735 10260 7769
rect 10226 7667 10260 7701
rect 10226 7599 10260 7633
rect 10226 7531 10260 7565
rect 10226 7463 10260 7497
rect 10226 7395 10260 7429
rect 10226 7327 10260 7361
rect 10226 7259 10260 7293
rect 10226 7191 10260 7225
rect 10226 7123 10260 7157
rect 10226 7055 10260 7089
rect 10226 6987 10260 7021
rect 10226 6919 10260 6953
rect 10226 6851 10260 6885
rect 10226 6783 10260 6817
rect 10226 6715 10260 6749
rect 10226 6647 10260 6681
rect 10226 6579 10260 6613
rect 10226 6511 10260 6545
rect 10226 6443 10260 6477
rect 10226 6375 10260 6409
rect 10226 6307 10260 6341
rect 10226 6239 10260 6273
rect 10226 6171 10260 6205
rect 10226 6103 10260 6137
rect 10226 6035 10260 6069
rect 10226 5967 10260 6001
rect 10226 5899 10260 5933
rect 10226 5831 10260 5865
rect 10226 5763 10260 5797
rect 10226 5695 10260 5729
rect 10226 5627 10260 5661
rect 10226 5559 10260 5593
rect 10226 5491 10260 5525
rect 10226 5423 10260 5457
rect 10226 5355 10260 5389
rect 10226 5287 10260 5321
rect 10226 5219 10260 5253
rect 10226 5151 10260 5185
rect 10226 5083 10260 5117
rect 10226 5015 10260 5049
rect 10226 4947 10260 4981
rect 10226 4879 10260 4913
rect 10226 4811 10260 4845
rect 10226 4743 10260 4777
rect 10226 4675 10260 4709
rect 10226 4607 10260 4641
rect 10226 4539 10260 4573
rect 10226 4471 10260 4505
rect 10226 4403 10260 4437
rect 10226 4335 10260 4369
rect 10226 4267 10260 4301
rect 10226 4199 10260 4233
rect 10226 4131 10260 4165
rect 10226 4063 10260 4097
rect 10226 3995 10260 4029
rect 10226 3927 10260 3961
rect 10226 3859 10260 3893
rect 10226 3791 10260 3825
rect 10226 3723 10260 3757
rect 10226 3655 10260 3689
rect 10226 3587 10260 3621
rect 10226 3519 10260 3553
rect 9088 3431 9122 3465
rect 9088 3363 9122 3397
rect 10226 3451 10260 3485
rect 11424 38655 11458 38689
rect 11424 38587 11458 38621
rect 11424 38519 11458 38553
rect 14940 38655 14974 38689
rect 13212 38596 13246 38630
rect 13212 38528 13246 38562
rect 11424 38451 11458 38485
rect 11424 38383 11458 38417
rect 11424 38315 11458 38349
rect 11424 38247 11458 38281
rect 11424 38179 11458 38213
rect 11424 38111 11458 38145
rect 11424 38043 11458 38077
rect 11424 37975 11458 38009
rect 11424 37907 11458 37941
rect 11424 37839 11458 37873
rect 11424 37771 11458 37805
rect 11424 37703 11458 37737
rect 11424 37635 11458 37669
rect 11424 37567 11458 37601
rect 11424 37499 11458 37533
rect 11424 37431 11458 37465
rect 11424 37363 11458 37397
rect 11424 37295 11458 37329
rect 11424 37227 11458 37261
rect 11424 37159 11458 37193
rect 11424 37091 11458 37125
rect 11424 37023 11458 37057
rect 11424 36955 11458 36989
rect 11424 36887 11458 36921
rect 11424 36819 11458 36853
rect 11424 36751 11458 36785
rect 11424 36683 11458 36717
rect 11424 36615 11458 36649
rect 11424 36547 11458 36581
rect 11424 36479 11458 36513
rect 11424 36411 11458 36445
rect 11424 36343 11458 36377
rect 11424 36275 11458 36309
rect 11424 36207 11458 36241
rect 11424 36139 11458 36173
rect 11424 36071 11458 36105
rect 11424 36003 11458 36037
rect 11424 35935 11458 35969
rect 11424 35867 11458 35901
rect 11424 35799 11458 35833
rect 11424 35731 11458 35765
rect 11424 35663 11458 35697
rect 11424 35595 11458 35629
rect 11424 35527 11458 35561
rect 11424 35459 11458 35493
rect 11424 35391 11458 35425
rect 11424 35323 11458 35357
rect 11424 35255 11458 35289
rect 11424 35187 11458 35221
rect 11424 35119 11458 35153
rect 11424 35051 11458 35085
rect 11424 34983 11458 35017
rect 11424 34915 11458 34949
rect 11424 34847 11458 34881
rect 11424 34779 11458 34813
rect 11424 34711 11458 34745
rect 11424 34643 11458 34677
rect 11424 34575 11458 34609
rect 11424 34507 11458 34541
rect 11424 34439 11458 34473
rect 11424 34371 11458 34405
rect 11424 34303 11458 34337
rect 11424 34235 11458 34269
rect 11424 34167 11458 34201
rect 11424 34099 11458 34133
rect 11424 34031 11458 34065
rect 11424 33963 11458 33997
rect 11424 33895 11458 33929
rect 11424 33827 11458 33861
rect 11424 33759 11458 33793
rect 11424 33691 11458 33725
rect 11424 33623 11458 33657
rect 11424 33555 11458 33589
rect 11424 33487 11458 33521
rect 11424 33419 11458 33453
rect 11424 33351 11458 33385
rect 11424 33283 11458 33317
rect 11424 33215 11458 33249
rect 11424 33147 11458 33181
rect 11424 33079 11458 33113
rect 11424 33011 11458 33045
rect 11424 32943 11458 32977
rect 11424 32875 11458 32909
rect 11424 32807 11458 32841
rect 11424 32739 11458 32773
rect 11424 32671 11458 32705
rect 11424 32603 11458 32637
rect 11424 32535 11458 32569
rect 11424 32467 11458 32501
rect 11424 32399 11458 32433
rect 11424 32331 11458 32365
rect 11424 32263 11458 32297
rect 11424 32195 11458 32229
rect 11424 32127 11458 32161
rect 11424 32059 11458 32093
rect 11424 31991 11458 32025
rect 11424 31923 11458 31957
rect 11424 31855 11458 31889
rect 11424 31787 11458 31821
rect 11424 31719 11458 31753
rect 11424 31651 11458 31685
rect 11424 31583 11458 31617
rect 11424 31515 11458 31549
rect 11424 31447 11458 31481
rect 11424 31379 11458 31413
rect 11424 31311 11458 31345
rect 11424 31243 11458 31277
rect 11424 31175 11458 31209
rect 11424 31107 11458 31141
rect 11424 31039 11458 31073
rect 11424 30971 11458 31005
rect 11424 30903 11458 30937
rect 11424 30835 11458 30869
rect 11424 30767 11458 30801
rect 11424 30699 11458 30733
rect 11424 30631 11458 30665
rect 11424 30563 11458 30597
rect 11424 30495 11458 30529
rect 11424 30427 11458 30461
rect 11424 30359 11458 30393
rect 11424 30291 11458 30325
rect 11424 30223 11458 30257
rect 11424 30155 11458 30189
rect 11424 30087 11458 30121
rect 11424 30019 11458 30053
rect 11424 29951 11458 29985
rect 11424 29883 11458 29917
rect 11424 29815 11458 29849
rect 11424 29747 11458 29781
rect 11424 29679 11458 29713
rect 11424 29611 11458 29645
rect 11424 29543 11458 29577
rect 11424 29475 11458 29509
rect 11424 29407 11458 29441
rect 11424 29339 11458 29373
rect 11424 29271 11458 29305
rect 11424 29203 11458 29237
rect 11424 29135 11458 29169
rect 11424 29067 11458 29101
rect 11424 28999 11458 29033
rect 11424 28931 11458 28965
rect 11424 28863 11458 28897
rect 11424 28795 11458 28829
rect 11424 28727 11458 28761
rect 11424 28659 11458 28693
rect 11424 28591 11458 28625
rect 11424 28523 11458 28557
rect 11424 28455 11458 28489
rect 11424 28387 11458 28421
rect 11424 28319 11458 28353
rect 11424 28251 11458 28285
rect 11424 28183 11458 28217
rect 11424 28115 11458 28149
rect 11424 28047 11458 28081
rect 11424 27979 11458 28013
rect 11424 27911 11458 27945
rect 11424 27843 11458 27877
rect 11424 27775 11458 27809
rect 11424 27707 11458 27741
rect 11424 27639 11458 27673
rect 11424 27571 11458 27605
rect 11424 27503 11458 27537
rect 11424 27435 11458 27469
rect 11424 27367 11458 27401
rect 11424 27299 11458 27333
rect 11424 27231 11458 27265
rect 11424 27163 11458 27197
rect 11424 27095 11458 27129
rect 11424 27027 11458 27061
rect 11424 26959 11458 26993
rect 11424 26891 11458 26925
rect 11424 26823 11458 26857
rect 11424 26755 11458 26789
rect 11424 26687 11458 26721
rect 11424 26619 11458 26653
rect 11424 26551 11458 26585
rect 11424 26483 11458 26517
rect 11424 26415 11458 26449
rect 11424 26347 11458 26381
rect 11424 26279 11458 26313
rect 11424 26211 11458 26245
rect 11424 26143 11458 26177
rect 11424 26075 11458 26109
rect 11424 26007 11458 26041
rect 11424 25939 11458 25973
rect 11424 25871 11458 25905
rect 11424 25803 11458 25837
rect 11424 25735 11458 25769
rect 11424 25667 11458 25701
rect 11424 25599 11458 25633
rect 11424 25531 11458 25565
rect 11424 25463 11458 25497
rect 11424 25395 11458 25429
rect 11424 25327 11458 25361
rect 11424 25259 11458 25293
rect 11424 25191 11458 25225
rect 11424 25123 11458 25157
rect 11424 25055 11458 25089
rect 11424 24987 11458 25021
rect 11424 24919 11458 24953
rect 11424 24851 11458 24885
rect 11424 24783 11458 24817
rect 11424 24715 11458 24749
rect 11424 24647 11458 24681
rect 11424 24579 11458 24613
rect 11424 24511 11458 24545
rect 11424 24443 11458 24477
rect 11424 24375 11458 24409
rect 11424 24307 11458 24341
rect 11424 24239 11458 24273
rect 11424 24171 11458 24205
rect 11424 24103 11458 24137
rect 11424 24035 11458 24069
rect 11424 23967 11458 24001
rect 11424 23899 11458 23933
rect 11424 23831 11458 23865
rect 11424 23763 11458 23797
rect 11424 23695 11458 23729
rect 11424 23627 11458 23661
rect 11424 23559 11458 23593
rect 11424 23491 11458 23525
rect 11424 23423 11458 23457
rect 11424 23355 11458 23389
rect 11424 23287 11458 23321
rect 11424 23219 11458 23253
rect 11424 23151 11458 23185
rect 11424 23083 11458 23117
rect 11424 23015 11458 23049
rect 11424 22947 11458 22981
rect 11424 22879 11458 22913
rect 11424 22811 11458 22845
rect 11424 22743 11458 22777
rect 11424 22675 11458 22709
rect 11424 22607 11458 22641
rect 11424 22539 11458 22573
rect 11424 22471 11458 22505
rect 11424 22403 11458 22437
rect 11424 22335 11458 22369
rect 11424 22267 11458 22301
rect 11424 22199 11458 22233
rect 11424 22131 11458 22165
rect 11424 22063 11458 22097
rect 11424 21995 11458 22029
rect 11424 21927 11458 21961
rect 11424 21859 11458 21893
rect 11424 21791 11458 21825
rect 11424 21723 11458 21757
rect 11424 21655 11458 21689
rect 11424 21587 11458 21621
rect 11424 21519 11458 21553
rect 11424 21451 11458 21485
rect 11424 21383 11458 21417
rect 11424 21315 11458 21349
rect 11424 21247 11458 21281
rect 11424 21179 11458 21213
rect 11424 21111 11458 21145
rect 11424 21043 11458 21077
rect 11424 20975 11458 21009
rect 11424 20907 11458 20941
rect 11424 20839 11458 20873
rect 11424 20771 11458 20805
rect 11424 20703 11458 20737
rect 11424 20635 11458 20669
rect 11424 20567 11458 20601
rect 11424 20499 11458 20533
rect 11424 20431 11458 20465
rect 11424 20363 11458 20397
rect 11424 20295 11458 20329
rect 11424 20227 11458 20261
rect 11424 20159 11458 20193
rect 11424 20091 11458 20125
rect 11424 20023 11458 20057
rect 11424 19955 11458 19989
rect 11424 19887 11458 19921
rect 11424 19819 11458 19853
rect 11424 19751 11458 19785
rect 11424 19683 11458 19717
rect 11424 19615 11458 19649
rect 11424 19547 11458 19581
rect 11424 19479 11458 19513
rect 11424 19411 11458 19445
rect 11424 19343 11458 19377
rect 11424 19275 11458 19309
rect 11424 19207 11458 19241
rect 11424 19139 11458 19173
rect 11424 19071 11458 19105
rect 11424 19003 11458 19037
rect 11424 18935 11458 18969
rect 11424 18867 11458 18901
rect 11424 18799 11458 18833
rect 11424 18731 11458 18765
rect 11424 18663 11458 18697
rect 11424 18595 11458 18629
rect 11424 18527 11458 18561
rect 11424 18459 11458 18493
rect 11424 18391 11458 18425
rect 11424 18323 11458 18357
rect 11424 18255 11458 18289
rect 11424 18187 11458 18221
rect 11424 18119 11458 18153
rect 11424 18051 11458 18085
rect 11424 17983 11458 18017
rect 11424 17915 11458 17949
rect 11424 17847 11458 17881
rect 11424 17779 11458 17813
rect 11424 17711 11458 17745
rect 11424 17643 11458 17677
rect 11424 17575 11458 17609
rect 11424 17507 11458 17541
rect 11424 17439 11458 17473
rect 11424 17371 11458 17405
rect 11424 17303 11458 17337
rect 11424 17235 11458 17269
rect 11424 17167 11458 17201
rect 11424 17099 11458 17133
rect 11424 17031 11458 17065
rect 11424 16963 11458 16997
rect 11424 16895 11458 16929
rect 11424 16827 11458 16861
rect 11424 16759 11458 16793
rect 11424 16691 11458 16725
rect 11424 16623 11458 16657
rect 11424 16555 11458 16589
rect 11424 16487 11458 16521
rect 11424 16419 11458 16453
rect 11424 16351 11458 16385
rect 11424 16283 11458 16317
rect 11424 16215 11458 16249
rect 11424 16147 11458 16181
rect 11424 16079 11458 16113
rect 11424 16011 11458 16045
rect 11424 15943 11458 15977
rect 11424 15875 11458 15909
rect 11424 15807 11458 15841
rect 11424 15739 11458 15773
rect 11424 15671 11458 15705
rect 11424 15603 11458 15637
rect 11424 15535 11458 15569
rect 11424 15467 11458 15501
rect 11424 15399 11458 15433
rect 11424 15331 11458 15365
rect 11424 15263 11458 15297
rect 11424 15195 11458 15229
rect 11424 15127 11458 15161
rect 11424 15059 11458 15093
rect 11424 14991 11458 15025
rect 11424 14923 11458 14957
rect 11424 14855 11458 14889
rect 11424 14787 11458 14821
rect 11424 14719 11458 14753
rect 11424 14651 11458 14685
rect 11424 14583 11458 14617
rect 11424 14515 11458 14549
rect 11424 14447 11458 14481
rect 11424 14379 11458 14413
rect 11424 14311 11458 14345
rect 11424 14243 11458 14277
rect 11424 14175 11458 14209
rect 11424 14107 11458 14141
rect 11424 14039 11458 14073
rect 11424 13971 11458 14005
rect 11424 13903 11458 13937
rect 11424 13835 11458 13869
rect 11424 13767 11458 13801
rect 11424 13699 11458 13733
rect 11424 13631 11458 13665
rect 11424 13563 11458 13597
rect 11424 13495 11458 13529
rect 11424 13427 11458 13461
rect 11424 13359 11458 13393
rect 11424 13291 11458 13325
rect 11424 13223 11458 13257
rect 11424 13155 11458 13189
rect 11424 13087 11458 13121
rect 11424 13019 11458 13053
rect 11424 12951 11458 12985
rect 11424 12883 11458 12917
rect 11424 12815 11458 12849
rect 11424 12747 11458 12781
rect 11424 12679 11458 12713
rect 11424 12611 11458 12645
rect 11424 12543 11458 12577
rect 11424 12475 11458 12509
rect 11424 12407 11458 12441
rect 11424 12339 11458 12373
rect 11424 12271 11458 12305
rect 11424 12203 11458 12237
rect 11424 12135 11458 12169
rect 11424 12067 11458 12101
rect 11424 11999 11458 12033
rect 11424 11931 11458 11965
rect 11424 11863 11458 11897
rect 11424 11795 11458 11829
rect 11424 11727 11458 11761
rect 11424 11659 11458 11693
rect 11424 11591 11458 11625
rect 11424 11523 11458 11557
rect 11424 11455 11458 11489
rect 11424 11387 11458 11421
rect 11424 11319 11458 11353
rect 11424 11251 11458 11285
rect 11424 11183 11458 11217
rect 11424 11115 11458 11149
rect 11424 11047 11458 11081
rect 11424 10979 11458 11013
rect 11424 10911 11458 10945
rect 11424 10843 11458 10877
rect 11424 10775 11458 10809
rect 11424 10707 11458 10741
rect 11424 10639 11458 10673
rect 11424 10571 11458 10605
rect 11424 10503 11458 10537
rect 11424 10435 11458 10469
rect 11424 10367 11458 10401
rect 11424 10299 11458 10333
rect 11424 10231 11458 10265
rect 11424 10163 11458 10197
rect 11424 10095 11458 10129
rect 11424 10027 11458 10061
rect 11424 9959 11458 9993
rect 11424 9891 11458 9925
rect 11424 9823 11458 9857
rect 11424 9755 11458 9789
rect 11424 9687 11458 9721
rect 11424 9619 11458 9653
rect 11424 9551 11458 9585
rect 11424 9483 11458 9517
rect 11424 9415 11458 9449
rect 11424 9347 11458 9381
rect 11424 9279 11458 9313
rect 11424 9211 11458 9245
rect 11424 9143 11458 9177
rect 11424 9075 11458 9109
rect 11424 9007 11458 9041
rect 11424 8939 11458 8973
rect 11424 8871 11458 8905
rect 11424 8803 11458 8837
rect 11424 8735 11458 8769
rect 11424 8667 11458 8701
rect 11424 8599 11458 8633
rect 11424 8531 11458 8565
rect 11424 8463 11458 8497
rect 11424 8395 11458 8429
rect 11424 8327 11458 8361
rect 11424 8259 11458 8293
rect 11424 8191 11458 8225
rect 11424 8123 11458 8157
rect 11424 8055 11458 8089
rect 11424 7987 11458 8021
rect 11424 7919 11458 7953
rect 11424 7851 11458 7885
rect 11424 7783 11458 7817
rect 11424 7715 11458 7749
rect 11424 7647 11458 7681
rect 11424 7579 11458 7613
rect 11424 7511 11458 7545
rect 11424 7443 11458 7477
rect 11424 7375 11458 7409
rect 11424 7307 11458 7341
rect 11424 7239 11458 7273
rect 11424 7171 11458 7205
rect 11424 7103 11458 7137
rect 11424 7035 11458 7069
rect 11424 6967 11458 7001
rect 11424 6899 11458 6933
rect 11424 6831 11458 6865
rect 11424 6763 11458 6797
rect 11424 6695 11458 6729
rect 11424 6627 11458 6661
rect 11424 6559 11458 6593
rect 11424 6491 11458 6525
rect 11424 6423 11458 6457
rect 11424 6355 11458 6389
rect 11424 6287 11458 6321
rect 11424 6219 11458 6253
rect 11424 6151 11458 6185
rect 11424 6083 11458 6117
rect 11424 6015 11458 6049
rect 11424 5947 11458 5981
rect 11424 5879 11458 5913
rect 11424 5811 11458 5845
rect 11424 5743 11458 5777
rect 11424 5675 11458 5709
rect 11424 5607 11458 5641
rect 11424 5539 11458 5573
rect 11424 5471 11458 5505
rect 11424 5403 11458 5437
rect 11424 5335 11458 5369
rect 11424 5267 11458 5301
rect 11424 5199 11458 5233
rect 11424 5131 11458 5165
rect 11424 5063 11458 5097
rect 11424 4995 11458 5029
rect 11424 4927 11458 4961
rect 11424 4859 11458 4893
rect 11424 4791 11458 4825
rect 11424 4723 11458 4757
rect 11424 4655 11458 4689
rect 11424 4587 11458 4621
rect 11424 4519 11458 4553
rect 11424 4451 11458 4485
rect 11424 4383 11458 4417
rect 11424 4315 11458 4349
rect 11424 4247 11458 4281
rect 11424 4179 11458 4213
rect 11424 4111 11458 4145
rect 11424 4043 11458 4077
rect 11424 3975 11458 4009
rect 11424 3907 11458 3941
rect 11424 3839 11458 3873
rect 11424 3771 11458 3805
rect 11424 3703 11458 3737
rect 11424 3635 11458 3669
rect 11424 3567 11458 3601
rect 11424 3499 11458 3533
rect 10226 3383 10260 3417
rect 9088 3295 9122 3329
rect 11424 3431 11458 3465
rect 11424 3363 11458 3397
rect 10226 3315 10260 3349
rect 10226 3247 10260 3281
rect 11424 3295 11458 3329
rect 9156 3179 9190 3213
rect 9224 3179 9258 3213
rect 9292 3179 9326 3213
rect 9360 3179 9394 3213
rect 9428 3179 9462 3213
rect 9496 3179 9530 3213
rect 9564 3179 9598 3213
rect 9632 3179 9666 3213
rect 9700 3179 9734 3213
rect 9768 3179 9802 3213
rect 9836 3179 9870 3213
rect 9904 3179 9938 3213
rect 9972 3179 10006 3213
rect 10040 3179 10074 3213
rect 10108 3179 10142 3213
rect 10336 3179 10370 3213
rect 10404 3179 10438 3213
rect 10472 3179 10506 3213
rect 10540 3179 10574 3213
rect 10608 3179 10642 3213
rect 10676 3179 10710 3213
rect 10744 3179 10778 3213
rect 10812 3179 10846 3213
rect 10880 3179 10914 3213
rect 10948 3179 10982 3213
rect 11016 3179 11050 3213
rect 11084 3179 11118 3213
rect 11152 3179 11186 3213
rect 11220 3179 11254 3213
rect 11288 3179 11322 3213
rect 11356 3179 11390 3213
rect 11424 3171 11458 3205
rect 11424 3103 11458 3137
rect 11424 3035 11458 3069
rect 11424 2967 11458 3001
rect 11424 2899 11458 2933
rect 11424 2831 11458 2865
rect 11424 2763 11458 2797
rect 11424 2695 11458 2729
rect 11424 2627 11458 2661
rect 11424 2559 11458 2593
rect 11424 2491 11458 2525
rect 11424 2423 11458 2457
rect 11424 2355 11458 2389
rect 11424 2287 11458 2321
rect 11424 2219 11458 2253
rect 11424 2151 11458 2185
rect 11424 2083 11458 2117
rect 11424 2015 11458 2049
rect 11424 1947 11458 1981
rect 11424 1879 11458 1913
rect 11424 1811 11458 1845
rect 11424 1743 11458 1777
rect 11424 1675 11458 1709
rect 11424 1607 11458 1641
rect 11424 1539 11458 1573
rect 11424 1471 11458 1505
rect 11424 1403 11458 1437
rect 11424 1335 11458 1369
rect 11424 1267 11458 1301
rect 11424 1199 11458 1233
rect 11424 1131 11458 1165
rect 11424 1063 11458 1097
rect 11424 995 11458 1029
rect 11424 927 11458 961
rect 11424 859 11458 893
rect 11424 791 11458 825
rect 11424 723 11458 757
rect 11424 655 11458 689
rect 11424 587 11458 621
rect 11424 519 11458 553
rect 11424 451 11458 485
rect 11424 383 11458 417
rect 14940 38587 14974 38621
rect 14940 38519 14974 38553
rect 13212 38460 13246 38494
rect 13212 38392 13246 38426
rect 13212 38324 13246 38358
rect 13212 38256 13246 38290
rect 13212 38188 13246 38222
rect 13212 38120 13246 38154
rect 13212 38052 13246 38086
rect 13212 37984 13246 38018
rect 13212 37916 13246 37950
rect 13212 37848 13246 37882
rect 13212 37780 13246 37814
rect 13212 37712 13246 37746
rect 13212 37644 13246 37678
rect 13212 37576 13246 37610
rect 13212 37508 13246 37542
rect 13212 37440 13246 37474
rect 13212 37372 13246 37406
rect 13212 37304 13246 37338
rect 13212 37236 13246 37270
rect 13212 37168 13246 37202
rect 13212 37100 13246 37134
rect 13212 37032 13246 37066
rect 13212 36964 13246 36998
rect 13212 36896 13246 36930
rect 13212 36828 13246 36862
rect 13212 36760 13246 36794
rect 13212 36692 13246 36726
rect 13212 36624 13246 36658
rect 13212 36556 13246 36590
rect 13212 36488 13246 36522
rect 13212 36420 13246 36454
rect 13212 36352 13246 36386
rect 13212 36284 13246 36318
rect 13212 36216 13246 36250
rect 13212 36148 13246 36182
rect 13212 36080 13246 36114
rect 13212 36012 13246 36046
rect 13212 35944 13246 35978
rect 13212 35876 13246 35910
rect 13212 35808 13246 35842
rect 13212 35740 13246 35774
rect 13212 35672 13246 35706
rect 13212 35604 13246 35638
rect 13212 35536 13246 35570
rect 13212 35468 13246 35502
rect 13212 35400 13246 35434
rect 13212 35332 13246 35366
rect 13212 35264 13246 35298
rect 13212 35196 13246 35230
rect 13212 35128 13246 35162
rect 13212 35060 13246 35094
rect 13212 34992 13246 35026
rect 13212 34924 13246 34958
rect 13212 34856 13246 34890
rect 13212 34788 13246 34822
rect 13212 34720 13246 34754
rect 13212 34652 13246 34686
rect 13212 34584 13246 34618
rect 13212 34516 13246 34550
rect 13212 34448 13246 34482
rect 13212 34380 13246 34414
rect 13212 34312 13246 34346
rect 13212 34244 13246 34278
rect 13212 34176 13246 34210
rect 13212 34108 13246 34142
rect 13212 34040 13246 34074
rect 13212 33972 13246 34006
rect 13212 33904 13246 33938
rect 13212 33836 13246 33870
rect 13212 33768 13246 33802
rect 13212 33700 13246 33734
rect 13212 33632 13246 33666
rect 13212 33564 13246 33598
rect 13212 33496 13246 33530
rect 13212 33428 13246 33462
rect 13212 33360 13246 33394
rect 13212 33292 13246 33326
rect 13212 33224 13246 33258
rect 13212 33156 13246 33190
rect 13212 33088 13246 33122
rect 13212 33020 13246 33054
rect 13212 32952 13246 32986
rect 13212 32884 13246 32918
rect 13212 32816 13246 32850
rect 13212 32748 13246 32782
rect 13212 32680 13246 32714
rect 13212 32612 13246 32646
rect 13212 32544 13246 32578
rect 13212 32476 13246 32510
rect 13212 32408 13246 32442
rect 13212 32340 13246 32374
rect 13212 32272 13246 32306
rect 13212 32204 13246 32238
rect 13212 32136 13246 32170
rect 13212 32068 13246 32102
rect 13212 32000 13246 32034
rect 13212 31932 13246 31966
rect 13212 31864 13246 31898
rect 13212 31796 13246 31830
rect 13212 31728 13246 31762
rect 13212 31660 13246 31694
rect 13212 31592 13246 31626
rect 13212 31524 13246 31558
rect 13212 31456 13246 31490
rect 13212 31388 13246 31422
rect 13212 31320 13246 31354
rect 13212 31252 13246 31286
rect 13212 31184 13246 31218
rect 13212 31116 13246 31150
rect 13212 31048 13246 31082
rect 13212 30980 13246 31014
rect 13212 30912 13246 30946
rect 13212 30844 13246 30878
rect 13212 30776 13246 30810
rect 13212 30708 13246 30742
rect 13212 30640 13246 30674
rect 13212 30572 13246 30606
rect 13212 30504 13246 30538
rect 13212 30436 13246 30470
rect 13212 30368 13246 30402
rect 13212 30300 13246 30334
rect 13212 30232 13246 30266
rect 13212 30164 13246 30198
rect 13212 30096 13246 30130
rect 13212 30028 13246 30062
rect 13212 29960 13246 29994
rect 13212 29892 13246 29926
rect 13212 29824 13246 29858
rect 13212 29756 13246 29790
rect 13212 29688 13246 29722
rect 13212 29620 13246 29654
rect 13212 29552 13246 29586
rect 13212 29484 13246 29518
rect 13212 29416 13246 29450
rect 13212 29348 13246 29382
rect 13212 29280 13246 29314
rect 13212 29212 13246 29246
rect 13212 29144 13246 29178
rect 13212 29076 13246 29110
rect 13212 29008 13246 29042
rect 13212 28940 13246 28974
rect 13212 28872 13246 28906
rect 13212 28804 13246 28838
rect 13212 28736 13246 28770
rect 13212 28668 13246 28702
rect 13212 28600 13246 28634
rect 13212 28532 13246 28566
rect 13212 28464 13246 28498
rect 13212 28396 13246 28430
rect 13212 28328 13246 28362
rect 13212 28260 13246 28294
rect 13212 28192 13246 28226
rect 13212 28124 13246 28158
rect 13212 28056 13246 28090
rect 13212 27988 13246 28022
rect 13212 27920 13246 27954
rect 13212 27852 13246 27886
rect 13212 27784 13246 27818
rect 13212 27716 13246 27750
rect 13212 27648 13246 27682
rect 13212 27580 13246 27614
rect 13212 27512 13246 27546
rect 13212 27444 13246 27478
rect 13212 27376 13246 27410
rect 13212 27308 13246 27342
rect 13212 27240 13246 27274
rect 13212 27172 13246 27206
rect 13212 27104 13246 27138
rect 13212 27036 13246 27070
rect 13212 26968 13246 27002
rect 13212 26900 13246 26934
rect 13212 26832 13246 26866
rect 13212 26764 13246 26798
rect 13212 26696 13246 26730
rect 13212 26628 13246 26662
rect 13212 26560 13246 26594
rect 13212 26492 13246 26526
rect 13212 26424 13246 26458
rect 13212 26356 13246 26390
rect 13212 26288 13246 26322
rect 13212 26220 13246 26254
rect 13212 26152 13246 26186
rect 13212 26084 13246 26118
rect 13212 26016 13246 26050
rect 13212 25948 13246 25982
rect 13212 25880 13246 25914
rect 13212 25812 13246 25846
rect 13212 25744 13246 25778
rect 13212 25676 13246 25710
rect 13212 25608 13246 25642
rect 13212 25540 13246 25574
rect 13212 25472 13246 25506
rect 13212 25404 13246 25438
rect 13212 25336 13246 25370
rect 13212 25268 13246 25302
rect 13212 25200 13246 25234
rect 13212 25132 13246 25166
rect 13212 25064 13246 25098
rect 13212 24996 13246 25030
rect 13212 24928 13246 24962
rect 13212 24860 13246 24894
rect 13212 24792 13246 24826
rect 13212 24724 13246 24758
rect 13212 24656 13246 24690
rect 13212 24588 13246 24622
rect 13212 24520 13246 24554
rect 13212 24452 13246 24486
rect 13212 24384 13246 24418
rect 13212 24316 13246 24350
rect 13212 24248 13246 24282
rect 13212 24180 13246 24214
rect 13212 24112 13246 24146
rect 13212 24044 13246 24078
rect 13212 23976 13246 24010
rect 13212 23908 13246 23942
rect 13212 23840 13246 23874
rect 13212 23772 13246 23806
rect 13212 23704 13246 23738
rect 13212 23636 13246 23670
rect 13212 23568 13246 23602
rect 13212 23500 13246 23534
rect 13212 23432 13246 23466
rect 13212 23364 13246 23398
rect 13212 23296 13246 23330
rect 13212 23228 13246 23262
rect 13212 23160 13246 23194
rect 13212 23092 13246 23126
rect 13212 23024 13246 23058
rect 13212 22956 13246 22990
rect 13212 22888 13246 22922
rect 13212 22820 13246 22854
rect 13212 22752 13246 22786
rect 13212 22684 13246 22718
rect 13212 22616 13246 22650
rect 13212 22548 13246 22582
rect 13212 22480 13246 22514
rect 13212 22412 13246 22446
rect 13212 22344 13246 22378
rect 13212 22276 13246 22310
rect 13212 22208 13246 22242
rect 13212 22140 13246 22174
rect 13212 22072 13246 22106
rect 13212 22004 13246 22038
rect 13212 21936 13246 21970
rect 13212 21868 13246 21902
rect 13212 21800 13246 21834
rect 13212 21732 13246 21766
rect 13212 21664 13246 21698
rect 13212 21596 13246 21630
rect 13212 21528 13246 21562
rect 13212 21460 13246 21494
rect 13212 21392 13246 21426
rect 13212 21324 13246 21358
rect 13212 21256 13246 21290
rect 13212 21188 13246 21222
rect 13212 21120 13246 21154
rect 13212 21052 13246 21086
rect 13212 20984 13246 21018
rect 13212 20916 13246 20950
rect 13212 20848 13246 20882
rect 13212 20780 13246 20814
rect 13212 20712 13246 20746
rect 13212 20644 13246 20678
rect 13212 20576 13246 20610
rect 13212 20508 13246 20542
rect 13212 20440 13246 20474
rect 13212 20372 13246 20406
rect 13212 20304 13246 20338
rect 13212 20236 13246 20270
rect 13212 20168 13246 20202
rect 13212 20100 13246 20134
rect 13212 20032 13246 20066
rect 13212 19964 13246 19998
rect 13212 19896 13246 19930
rect 13212 19828 13246 19862
rect 13212 19760 13246 19794
rect 13212 19692 13246 19726
rect 13212 19624 13246 19658
rect 13212 19556 13246 19590
rect 13212 19488 13246 19522
rect 13212 19420 13246 19454
rect 13212 19352 13246 19386
rect 13212 19284 13246 19318
rect 13212 19216 13246 19250
rect 13212 19148 13246 19182
rect 13212 19080 13246 19114
rect 13212 19012 13246 19046
rect 13212 18944 13246 18978
rect 13212 18876 13246 18910
rect 13212 18808 13246 18842
rect 13212 18740 13246 18774
rect 13212 18672 13246 18706
rect 13212 18604 13246 18638
rect 13212 18536 13246 18570
rect 13212 18468 13246 18502
rect 13212 18400 13246 18434
rect 13212 18332 13246 18366
rect 13212 18264 13246 18298
rect 13212 18196 13246 18230
rect 13212 18128 13246 18162
rect 13212 18060 13246 18094
rect 13212 17992 13246 18026
rect 13212 17924 13246 17958
rect 13212 17856 13246 17890
rect 13212 17788 13246 17822
rect 13212 17720 13246 17754
rect 13212 17652 13246 17686
rect 13212 17584 13246 17618
rect 13212 17516 13246 17550
rect 13212 17448 13246 17482
rect 13212 17380 13246 17414
rect 13212 17312 13246 17346
rect 13212 17244 13246 17278
rect 13212 17176 13246 17210
rect 13212 17108 13246 17142
rect 13212 17040 13246 17074
rect 13212 16972 13246 17006
rect 13212 16904 13246 16938
rect 13212 16836 13246 16870
rect 13212 16768 13246 16802
rect 13212 16700 13246 16734
rect 13212 16632 13246 16666
rect 13212 16564 13246 16598
rect 13212 16496 13246 16530
rect 13212 16428 13246 16462
rect 13212 16360 13246 16394
rect 13212 16292 13246 16326
rect 13212 16224 13246 16258
rect 13212 16156 13246 16190
rect 13212 16088 13246 16122
rect 13212 16020 13246 16054
rect 13212 15952 13246 15986
rect 13212 15884 13246 15918
rect 13212 15816 13246 15850
rect 13212 15748 13246 15782
rect 13212 15680 13246 15714
rect 13212 15612 13246 15646
rect 13212 15544 13246 15578
rect 13212 15476 13246 15510
rect 13212 15408 13246 15442
rect 13212 15340 13246 15374
rect 13212 15272 13246 15306
rect 13212 15204 13246 15238
rect 13212 15136 13246 15170
rect 13212 15068 13246 15102
rect 13212 15000 13246 15034
rect 13212 14932 13246 14966
rect 13212 14864 13246 14898
rect 13212 14796 13246 14830
rect 13212 14728 13246 14762
rect 13212 14660 13246 14694
rect 13212 14592 13246 14626
rect 13212 14524 13246 14558
rect 13212 14456 13246 14490
rect 13212 14388 13246 14422
rect 13212 14320 13246 14354
rect 13212 14252 13246 14286
rect 13212 14184 13246 14218
rect 13212 14116 13246 14150
rect 13212 14048 13246 14082
rect 13212 13980 13246 14014
rect 13212 13912 13246 13946
rect 13212 13844 13246 13878
rect 13212 13776 13246 13810
rect 13212 13708 13246 13742
rect 13212 13640 13246 13674
rect 13212 13572 13246 13606
rect 13212 13504 13246 13538
rect 13212 13436 13246 13470
rect 13212 13368 13246 13402
rect 13212 13300 13246 13334
rect 13212 13232 13246 13266
rect 13212 13164 13246 13198
rect 13212 13096 13246 13130
rect 13212 13028 13246 13062
rect 13212 12960 13246 12994
rect 13212 12892 13246 12926
rect 13212 12824 13246 12858
rect 13212 12756 13246 12790
rect 13212 12688 13246 12722
rect 13212 12620 13246 12654
rect 13212 12552 13246 12586
rect 13212 12484 13246 12518
rect 13212 12416 13246 12450
rect 13212 12348 13246 12382
rect 13212 12280 13246 12314
rect 13212 12212 13246 12246
rect 13212 12144 13246 12178
rect 13212 12076 13246 12110
rect 13212 12008 13246 12042
rect 13212 11940 13246 11974
rect 13212 11872 13246 11906
rect 13212 11804 13246 11838
rect 13212 11736 13246 11770
rect 13212 11668 13246 11702
rect 13212 11600 13246 11634
rect 13212 11532 13246 11566
rect 13212 11464 13246 11498
rect 13212 11396 13246 11430
rect 13212 11328 13246 11362
rect 13212 11260 13246 11294
rect 13212 11192 13246 11226
rect 13212 11124 13246 11158
rect 13212 11056 13246 11090
rect 13212 10988 13246 11022
rect 13212 10920 13246 10954
rect 13212 10852 13246 10886
rect 13212 10784 13246 10818
rect 13212 10716 13246 10750
rect 13212 10648 13246 10682
rect 13212 10580 13246 10614
rect 13212 10512 13246 10546
rect 13212 10444 13246 10478
rect 13212 10376 13246 10410
rect 13212 10308 13246 10342
rect 13212 10240 13246 10274
rect 13212 10172 13246 10206
rect 13212 10104 13246 10138
rect 13212 10036 13246 10070
rect 13212 9968 13246 10002
rect 13212 9900 13246 9934
rect 13212 9832 13246 9866
rect 13212 9764 13246 9798
rect 13212 9696 13246 9730
rect 13212 9628 13246 9662
rect 13212 9560 13246 9594
rect 13212 9492 13246 9526
rect 13212 9424 13246 9458
rect 13212 9356 13246 9390
rect 13212 9288 13246 9322
rect 13212 9220 13246 9254
rect 13212 9152 13246 9186
rect 13212 9084 13246 9118
rect 13212 9016 13246 9050
rect 13212 8948 13246 8982
rect 13212 8880 13246 8914
rect 13212 8812 13246 8846
rect 13212 8744 13246 8778
rect 13212 8676 13246 8710
rect 13212 8608 13246 8642
rect 13212 8540 13246 8574
rect 13212 8472 13246 8506
rect 13212 8404 13246 8438
rect 13212 8336 13246 8370
rect 13212 8268 13246 8302
rect 13212 8200 13246 8234
rect 13212 8132 13246 8166
rect 13212 8064 13246 8098
rect 13212 7996 13246 8030
rect 13212 7928 13246 7962
rect 13212 7860 13246 7894
rect 13212 7792 13246 7826
rect 13212 7724 13246 7758
rect 13212 7656 13246 7690
rect 13212 7588 13246 7622
rect 13212 7520 13246 7554
rect 13212 7452 13246 7486
rect 13212 7384 13246 7418
rect 13212 7316 13246 7350
rect 13212 7248 13246 7282
rect 13212 7180 13246 7214
rect 13212 7112 13246 7146
rect 13212 7044 13246 7078
rect 13212 6976 13246 7010
rect 13212 6908 13246 6942
rect 13212 6840 13246 6874
rect 13212 6772 13246 6806
rect 13212 6704 13246 6738
rect 13212 6636 13246 6670
rect 13212 6568 13246 6602
rect 13212 6500 13246 6534
rect 13212 6432 13246 6466
rect 13212 6364 13246 6398
rect 13212 6296 13246 6330
rect 13212 6228 13246 6262
rect 13212 6160 13246 6194
rect 13212 6092 13246 6126
rect 13212 6024 13246 6058
rect 13212 5956 13246 5990
rect 13212 5888 13246 5922
rect 13212 5820 13246 5854
rect 13212 5752 13246 5786
rect 13212 5684 13246 5718
rect 13212 5616 13246 5650
rect 13212 5548 13246 5582
rect 13212 5480 13246 5514
rect 13212 5412 13246 5446
rect 13212 5344 13246 5378
rect 13212 5276 13246 5310
rect 13212 5208 13246 5242
rect 13212 5140 13246 5174
rect 13212 5072 13246 5106
rect 13212 5004 13246 5038
rect 13212 4936 13246 4970
rect 13212 4868 13246 4902
rect 13212 4800 13246 4834
rect 13212 4732 13246 4766
rect 13212 4664 13246 4698
rect 13212 4596 13246 4630
rect 13212 4528 13246 4562
rect 13212 4460 13246 4494
rect 13212 4392 13246 4426
rect 13212 4324 13246 4358
rect 13212 4256 13246 4290
rect 13212 4188 13246 4222
rect 13212 4120 13246 4154
rect 13212 4052 13246 4086
rect 13212 3984 13246 4018
rect 13212 3916 13246 3950
rect 13212 3848 13246 3882
rect 13212 3780 13246 3814
rect 13212 3712 13246 3746
rect 13212 3644 13246 3678
rect 13212 3576 13246 3610
rect 13212 3508 13246 3542
rect 13212 3440 13246 3474
rect 13212 3372 13246 3406
rect 13212 3304 13246 3338
rect 13212 3236 13246 3270
rect 13212 3168 13246 3202
rect 13212 3100 13246 3134
rect 13212 3032 13246 3066
rect 13212 2964 13246 2998
rect 13212 2896 13246 2930
rect 13212 2828 13246 2862
rect 13212 2760 13246 2794
rect 13212 2692 13246 2726
rect 13212 2624 13246 2658
rect 13212 2556 13246 2590
rect 13212 2488 13246 2522
rect 13212 2420 13246 2454
rect 13212 2352 13246 2386
rect 13212 2284 13246 2318
rect 13212 2216 13246 2250
rect 13212 2148 13246 2182
rect 13212 2080 13246 2114
rect 13212 2012 13246 2046
rect 13212 1944 13246 1978
rect 13212 1876 13246 1910
rect 13212 1808 13246 1842
rect 13212 1740 13246 1774
rect 13212 1672 13246 1706
rect 13212 1604 13246 1638
rect 13212 1536 13246 1570
rect 13212 1468 13246 1502
rect 13212 1400 13246 1434
rect 13212 1332 13246 1366
rect 13212 1264 13246 1298
rect 13212 1196 13246 1230
rect 13212 1128 13246 1162
rect 13212 1060 13246 1094
rect 13212 992 13246 1026
rect 13212 924 13246 958
rect 13212 856 13246 890
rect 13212 788 13246 822
rect 13212 720 13246 754
rect 13212 652 13246 686
rect 13212 584 13246 618
rect 13212 516 13246 550
rect 13212 448 13246 482
rect 11424 315 11458 349
rect 11424 247 11458 281
rect 13212 380 13246 414
rect 14940 38451 14974 38485
rect 14940 38383 14974 38417
rect 14940 38315 14974 38349
rect 14940 38247 14974 38281
rect 14940 38179 14974 38213
rect 14940 38111 14974 38145
rect 14940 38043 14974 38077
rect 14940 37975 14974 38009
rect 14940 37907 14974 37941
rect 14940 37839 14974 37873
rect 14940 37771 14974 37805
rect 14940 37703 14974 37737
rect 14940 37635 14974 37669
rect 14940 37567 14974 37601
rect 14940 37499 14974 37533
rect 14940 37431 14974 37465
rect 14940 37363 14974 37397
rect 14940 37295 14974 37329
rect 14940 37227 14974 37261
rect 14940 37159 14974 37193
rect 14940 37091 14974 37125
rect 14940 37023 14974 37057
rect 14940 36955 14974 36989
rect 14940 36887 14974 36921
rect 14940 36819 14974 36853
rect 14940 36751 14974 36785
rect 14940 36683 14974 36717
rect 14940 36615 14974 36649
rect 14940 36547 14974 36581
rect 14940 36479 14974 36513
rect 14940 36411 14974 36445
rect 14940 36343 14974 36377
rect 14940 36275 14974 36309
rect 14940 36207 14974 36241
rect 14940 36139 14974 36173
rect 14940 36071 14974 36105
rect 14940 36003 14974 36037
rect 14940 35935 14974 35969
rect 14940 35867 14974 35901
rect 14940 35799 14974 35833
rect 14940 35731 14974 35765
rect 14940 35663 14974 35697
rect 14940 35595 14974 35629
rect 14940 35527 14974 35561
rect 14940 35459 14974 35493
rect 14940 35391 14974 35425
rect 14940 35323 14974 35357
rect 14940 35255 14974 35289
rect 14940 35187 14974 35221
rect 14940 35119 14974 35153
rect 14940 35051 14974 35085
rect 14940 34983 14974 35017
rect 14940 34915 14974 34949
rect 14940 34847 14974 34881
rect 14940 34779 14974 34813
rect 14940 34711 14974 34745
rect 14940 34643 14974 34677
rect 14940 34575 14974 34609
rect 14940 34507 14974 34541
rect 14940 34439 14974 34473
rect 14940 34371 14974 34405
rect 14940 34303 14974 34337
rect 14940 34235 14974 34269
rect 14940 34167 14974 34201
rect 14940 34099 14974 34133
rect 14940 34031 14974 34065
rect 14940 33963 14974 33997
rect 14940 33895 14974 33929
rect 14940 33827 14974 33861
rect 14940 33759 14974 33793
rect 14940 33691 14974 33725
rect 14940 33623 14974 33657
rect 14940 33555 14974 33589
rect 14940 33487 14974 33521
rect 14940 33419 14974 33453
rect 14940 33351 14974 33385
rect 14940 33283 14974 33317
rect 14940 33215 14974 33249
rect 14940 33147 14974 33181
rect 14940 33079 14974 33113
rect 14940 33011 14974 33045
rect 14940 32943 14974 32977
rect 14940 32875 14974 32909
rect 14940 32807 14974 32841
rect 14940 32739 14974 32773
rect 14940 32671 14974 32705
rect 14940 32603 14974 32637
rect 14940 32535 14974 32569
rect 14940 32467 14974 32501
rect 14940 32399 14974 32433
rect 14940 32331 14974 32365
rect 14940 32263 14974 32297
rect 14940 32195 14974 32229
rect 14940 32127 14974 32161
rect 14940 32059 14974 32093
rect 14940 31991 14974 32025
rect 14940 31923 14974 31957
rect 14940 31855 14974 31889
rect 14940 31787 14974 31821
rect 14940 31719 14974 31753
rect 14940 31651 14974 31685
rect 14940 31583 14974 31617
rect 14940 31515 14974 31549
rect 14940 31447 14974 31481
rect 14940 31379 14974 31413
rect 14940 31311 14974 31345
rect 14940 31243 14974 31277
rect 14940 31175 14974 31209
rect 14940 31107 14974 31141
rect 14940 31039 14974 31073
rect 14940 30971 14974 31005
rect 14940 30903 14974 30937
rect 14940 30835 14974 30869
rect 14940 30767 14974 30801
rect 14940 30699 14974 30733
rect 14940 30631 14974 30665
rect 14940 30563 14974 30597
rect 14940 30495 14974 30529
rect 14940 30427 14974 30461
rect 14940 30359 14974 30393
rect 14940 30291 14974 30325
rect 14940 30223 14974 30257
rect 14940 30155 14974 30189
rect 14940 30087 14974 30121
rect 14940 30019 14974 30053
rect 14940 29951 14974 29985
rect 14940 29883 14974 29917
rect 14940 29815 14974 29849
rect 14940 29747 14974 29781
rect 14940 29679 14974 29713
rect 14940 29611 14974 29645
rect 14940 29543 14974 29577
rect 14940 29475 14974 29509
rect 14940 29407 14974 29441
rect 14940 29339 14974 29373
rect 14940 29271 14974 29305
rect 14940 29203 14974 29237
rect 14940 29135 14974 29169
rect 14940 29067 14974 29101
rect 14940 28999 14974 29033
rect 14940 28931 14974 28965
rect 14940 28863 14974 28897
rect 14940 28795 14974 28829
rect 14940 28727 14974 28761
rect 14940 28659 14974 28693
rect 14940 28591 14974 28625
rect 14940 28523 14974 28557
rect 14940 28455 14974 28489
rect 14940 28387 14974 28421
rect 14940 28319 14974 28353
rect 14940 28251 14974 28285
rect 14940 28183 14974 28217
rect 14940 28115 14974 28149
rect 14940 28047 14974 28081
rect 14940 27979 14974 28013
rect 14940 27911 14974 27945
rect 14940 27843 14974 27877
rect 14940 27775 14974 27809
rect 14940 27707 14974 27741
rect 14940 27639 14974 27673
rect 14940 27571 14974 27605
rect 14940 27503 14974 27537
rect 14940 27435 14974 27469
rect 14940 27367 14974 27401
rect 14940 27299 14974 27333
rect 14940 27231 14974 27265
rect 14940 27163 14974 27197
rect 14940 27095 14974 27129
rect 14940 27027 14974 27061
rect 14940 26959 14974 26993
rect 14940 26891 14974 26925
rect 14940 26823 14974 26857
rect 14940 26755 14974 26789
rect 14940 26687 14974 26721
rect 14940 26619 14974 26653
rect 14940 26551 14974 26585
rect 14940 26483 14974 26517
rect 14940 26415 14974 26449
rect 14940 26347 14974 26381
rect 14940 26279 14974 26313
rect 14940 26211 14974 26245
rect 14940 26143 14974 26177
rect 14940 26075 14974 26109
rect 14940 26007 14974 26041
rect 14940 25939 14974 25973
rect 14940 25871 14974 25905
rect 14940 25803 14974 25837
rect 14940 25735 14974 25769
rect 14940 25667 14974 25701
rect 14940 25599 14974 25633
rect 14940 25531 14974 25565
rect 14940 25463 14974 25497
rect 14940 25395 14974 25429
rect 14940 25327 14974 25361
rect 14940 25259 14974 25293
rect 14940 25191 14974 25225
rect 14940 25123 14974 25157
rect 14940 25055 14974 25089
rect 14940 24987 14974 25021
rect 14940 24919 14974 24953
rect 14940 24851 14974 24885
rect 14940 24783 14974 24817
rect 14940 24715 14974 24749
rect 14940 24647 14974 24681
rect 14940 24579 14974 24613
rect 14940 24511 14974 24545
rect 14940 24443 14974 24477
rect 14940 24375 14974 24409
rect 14940 24307 14974 24341
rect 14940 24239 14974 24273
rect 14940 24171 14974 24205
rect 14940 24103 14974 24137
rect 14940 24035 14974 24069
rect 14940 23967 14974 24001
rect 14940 23899 14974 23933
rect 14940 23831 14974 23865
rect 14940 23763 14974 23797
rect 14940 23695 14974 23729
rect 14940 23627 14974 23661
rect 14940 23559 14974 23593
rect 14940 23491 14974 23525
rect 14940 23423 14974 23457
rect 14940 23355 14974 23389
rect 14940 23287 14974 23321
rect 14940 23219 14974 23253
rect 14940 23151 14974 23185
rect 14940 23083 14974 23117
rect 14940 23015 14974 23049
rect 14940 22947 14974 22981
rect 14940 22879 14974 22913
rect 14940 22811 14974 22845
rect 14940 22743 14974 22777
rect 14940 22675 14974 22709
rect 14940 22607 14974 22641
rect 14940 22539 14974 22573
rect 14940 22471 14974 22505
rect 14940 22403 14974 22437
rect 14940 22335 14974 22369
rect 14940 22267 14974 22301
rect 14940 22199 14974 22233
rect 14940 22131 14974 22165
rect 14940 22063 14974 22097
rect 14940 21995 14974 22029
rect 14940 21927 14974 21961
rect 14940 21859 14974 21893
rect 14940 21791 14974 21825
rect 14940 21723 14974 21757
rect 14940 21655 14974 21689
rect 14940 21587 14974 21621
rect 14940 21519 14974 21553
rect 14940 21451 14974 21485
rect 14940 21383 14974 21417
rect 14940 21315 14974 21349
rect 14940 21247 14974 21281
rect 14940 21179 14974 21213
rect 14940 21111 14974 21145
rect 14940 21043 14974 21077
rect 14940 20975 14974 21009
rect 14940 20907 14974 20941
rect 14940 20839 14974 20873
rect 14940 20771 14974 20805
rect 14940 20703 14974 20737
rect 14940 20635 14974 20669
rect 14940 20567 14974 20601
rect 14940 20499 14974 20533
rect 14940 20431 14974 20465
rect 14940 20363 14974 20397
rect 14940 20295 14974 20329
rect 14940 20227 14974 20261
rect 14940 20159 14974 20193
rect 14940 20091 14974 20125
rect 14940 20023 14974 20057
rect 14940 19955 14974 19989
rect 14940 19887 14974 19921
rect 14940 19819 14974 19853
rect 14940 19751 14974 19785
rect 14940 19683 14974 19717
rect 14940 19615 14974 19649
rect 14940 19547 14974 19581
rect 14940 19479 14974 19513
rect 14940 19411 14974 19445
rect 14940 19343 14974 19377
rect 14940 19275 14974 19309
rect 14940 19207 14974 19241
rect 14940 19139 14974 19173
rect 14940 19071 14974 19105
rect 14940 19003 14974 19037
rect 14940 18935 14974 18969
rect 14940 18867 14974 18901
rect 14940 18799 14974 18833
rect 14940 18731 14974 18765
rect 14940 18663 14974 18697
rect 14940 18595 14974 18629
rect 14940 18527 14974 18561
rect 14940 18459 14974 18493
rect 14940 18391 14974 18425
rect 14940 18323 14974 18357
rect 14940 18255 14974 18289
rect 14940 18187 14974 18221
rect 14940 18119 14974 18153
rect 14940 18051 14974 18085
rect 14940 17983 14974 18017
rect 14940 17915 14974 17949
rect 14940 17847 14974 17881
rect 14940 17779 14974 17813
rect 14940 17711 14974 17745
rect 14940 17643 14974 17677
rect 14940 17575 14974 17609
rect 14940 17507 14974 17541
rect 14940 17439 14974 17473
rect 14940 17371 14974 17405
rect 14940 17303 14974 17337
rect 14940 17235 14974 17269
rect 14940 17167 14974 17201
rect 14940 17099 14974 17133
rect 14940 17031 14974 17065
rect 14940 16963 14974 16997
rect 14940 16895 14974 16929
rect 14940 16827 14974 16861
rect 14940 16759 14974 16793
rect 14940 16691 14974 16725
rect 14940 16623 14974 16657
rect 14940 16555 14974 16589
rect 14940 16487 14974 16521
rect 14940 16419 14974 16453
rect 14940 16351 14974 16385
rect 14940 16283 14974 16317
rect 14940 16215 14974 16249
rect 14940 16147 14974 16181
rect 14940 16079 14974 16113
rect 14940 16011 14974 16045
rect 14940 15943 14974 15977
rect 14940 15875 14974 15909
rect 14940 15807 14974 15841
rect 14940 15739 14974 15773
rect 14940 15671 14974 15705
rect 14940 15603 14974 15637
rect 14940 15535 14974 15569
rect 14940 15467 14974 15501
rect 14940 15399 14974 15433
rect 14940 15331 14974 15365
rect 14940 15263 14974 15297
rect 14940 15195 14974 15229
rect 14940 15127 14974 15161
rect 14940 15059 14974 15093
rect 14940 14991 14974 15025
rect 14940 14923 14974 14957
rect 14940 14855 14974 14889
rect 14940 14787 14974 14821
rect 14940 14719 14974 14753
rect 14940 14651 14974 14685
rect 14940 14583 14974 14617
rect 14940 14515 14974 14549
rect 14940 14447 14974 14481
rect 14940 14379 14974 14413
rect 14940 14311 14974 14345
rect 14940 14243 14974 14277
rect 14940 14175 14974 14209
rect 14940 14107 14974 14141
rect 14940 14039 14974 14073
rect 14940 13971 14974 14005
rect 14940 13903 14974 13937
rect 14940 13835 14974 13869
rect 14940 13767 14974 13801
rect 14940 13699 14974 13733
rect 14940 13631 14974 13665
rect 14940 13563 14974 13597
rect 14940 13495 14974 13529
rect 14940 13427 14974 13461
rect 14940 13359 14974 13393
rect 14940 13291 14974 13325
rect 14940 13223 14974 13257
rect 14940 13155 14974 13189
rect 14940 13087 14974 13121
rect 14940 13019 14974 13053
rect 14940 12951 14974 12985
rect 14940 12883 14974 12917
rect 14940 12815 14974 12849
rect 14940 12747 14974 12781
rect 14940 12679 14974 12713
rect 14940 12611 14974 12645
rect 14940 12543 14974 12577
rect 14940 12475 14974 12509
rect 14940 12407 14974 12441
rect 14940 12339 14974 12373
rect 14940 12271 14974 12305
rect 14940 12203 14974 12237
rect 14940 12135 14974 12169
rect 14940 12067 14974 12101
rect 14940 11999 14974 12033
rect 14940 11931 14974 11965
rect 14940 11863 14974 11897
rect 14940 11795 14974 11829
rect 14940 11727 14974 11761
rect 14940 11659 14974 11693
rect 14940 11591 14974 11625
rect 14940 11523 14974 11557
rect 14940 11455 14974 11489
rect 14940 11387 14974 11421
rect 14940 11319 14974 11353
rect 14940 11251 14974 11285
rect 14940 11183 14974 11217
rect 14940 11115 14974 11149
rect 14940 11047 14974 11081
rect 14940 10979 14974 11013
rect 14940 10911 14974 10945
rect 14940 10843 14974 10877
rect 14940 10775 14974 10809
rect 14940 10707 14974 10741
rect 14940 10639 14974 10673
rect 14940 10571 14974 10605
rect 14940 10503 14974 10537
rect 14940 10435 14974 10469
rect 14940 10367 14974 10401
rect 14940 10299 14974 10333
rect 14940 10231 14974 10265
rect 14940 10163 14974 10197
rect 14940 10095 14974 10129
rect 14940 10027 14974 10061
rect 14940 9959 14974 9993
rect 14940 9891 14974 9925
rect 14940 9823 14974 9857
rect 14940 9755 14974 9789
rect 14940 9687 14974 9721
rect 14940 9619 14974 9653
rect 14940 9551 14974 9585
rect 14940 9483 14974 9517
rect 14940 9415 14974 9449
rect 14940 9347 14974 9381
rect 14940 9279 14974 9313
rect 14940 9211 14974 9245
rect 14940 9143 14974 9177
rect 14940 9075 14974 9109
rect 14940 9007 14974 9041
rect 14940 8939 14974 8973
rect 14940 8871 14974 8905
rect 14940 8803 14974 8837
rect 14940 8735 14974 8769
rect 14940 8667 14974 8701
rect 14940 8599 14974 8633
rect 14940 8531 14974 8565
rect 14940 8463 14974 8497
rect 14940 8395 14974 8429
rect 14940 8327 14974 8361
rect 14940 8259 14974 8293
rect 14940 8191 14974 8225
rect 14940 8123 14974 8157
rect 14940 8055 14974 8089
rect 14940 7987 14974 8021
rect 14940 7919 14974 7953
rect 14940 7851 14974 7885
rect 14940 7783 14974 7817
rect 14940 7715 14974 7749
rect 14940 7647 14974 7681
rect 14940 7579 14974 7613
rect 14940 7511 14974 7545
rect 14940 7443 14974 7477
rect 14940 7375 14974 7409
rect 14940 7307 14974 7341
rect 14940 7239 14974 7273
rect 14940 7171 14974 7205
rect 14940 7103 14974 7137
rect 14940 7035 14974 7069
rect 14940 6967 14974 7001
rect 14940 6899 14974 6933
rect 14940 6831 14974 6865
rect 14940 6763 14974 6797
rect 14940 6695 14974 6729
rect 14940 6627 14974 6661
rect 14940 6559 14974 6593
rect 14940 6491 14974 6525
rect 14940 6423 14974 6457
rect 14940 6355 14974 6389
rect 14940 6287 14974 6321
rect 14940 6219 14974 6253
rect 14940 6151 14974 6185
rect 14940 6083 14974 6117
rect 14940 6015 14974 6049
rect 14940 5947 14974 5981
rect 14940 5879 14974 5913
rect 14940 5811 14974 5845
rect 14940 5743 14974 5777
rect 14940 5675 14974 5709
rect 14940 5607 14974 5641
rect 14940 5539 14974 5573
rect 14940 5471 14974 5505
rect 14940 5403 14974 5437
rect 14940 5335 14974 5369
rect 14940 5267 14974 5301
rect 14940 5199 14974 5233
rect 14940 5131 14974 5165
rect 14940 5063 14974 5097
rect 14940 4995 14974 5029
rect 14940 4927 14974 4961
rect 14940 4859 14974 4893
rect 14940 4791 14974 4825
rect 14940 4723 14974 4757
rect 14940 4655 14974 4689
rect 14940 4587 14974 4621
rect 14940 4519 14974 4553
rect 14940 4451 14974 4485
rect 14940 4383 14974 4417
rect 14940 4315 14974 4349
rect 14940 4247 14974 4281
rect 14940 4179 14974 4213
rect 14940 4111 14974 4145
rect 14940 4043 14974 4077
rect 14940 3975 14974 4009
rect 14940 3907 14974 3941
rect 14940 3839 14974 3873
rect 14940 3771 14974 3805
rect 14940 3703 14974 3737
rect 14940 3635 14974 3669
rect 14940 3567 14974 3601
rect 14940 3499 14974 3533
rect 14940 3431 14974 3465
rect 14940 3363 14974 3397
rect 14940 3295 14974 3329
rect 14940 3171 14974 3205
rect 14940 3103 14974 3137
rect 14940 3035 14974 3069
rect 14940 2967 14974 3001
rect 14940 2899 14974 2933
rect 14940 2831 14974 2865
rect 14940 2763 14974 2797
rect 14940 2695 14974 2729
rect 14940 2627 14974 2661
rect 14940 2559 14974 2593
rect 14940 2491 14974 2525
rect 14940 2423 14974 2457
rect 14940 2355 14974 2389
rect 14940 2287 14974 2321
rect 14940 2219 14974 2253
rect 14940 2151 14974 2185
rect 14940 2083 14974 2117
rect 14940 2015 14974 2049
rect 14940 1947 14974 1981
rect 14940 1879 14974 1913
rect 14940 1811 14974 1845
rect 14940 1743 14974 1777
rect 14940 1675 14974 1709
rect 14940 1607 14974 1641
rect 14940 1539 14974 1573
rect 14940 1471 14974 1505
rect 14940 1403 14974 1437
rect 14940 1335 14974 1369
rect 14940 1267 14974 1301
rect 14940 1199 14974 1233
rect 14940 1131 14974 1165
rect 14940 1063 14974 1097
rect 14940 995 14974 1029
rect 14940 927 14974 961
rect 14940 859 14974 893
rect 14940 791 14974 825
rect 14940 723 14974 757
rect 14940 655 14974 689
rect 14940 587 14974 621
rect 14940 519 14974 553
rect 14940 451 14974 485
rect 13212 312 13246 346
rect 11424 179 11458 213
rect 11424 111 11458 145
rect 13212 244 13246 278
rect 14940 383 14974 417
rect 14940 315 14974 349
rect 13212 176 13246 210
rect 13212 108 13246 142
rect 14940 247 14974 281
rect 14940 179 14974 213
rect 14940 111 14974 145
rect 11492 40 11526 74
rect 11560 40 11594 74
rect 11628 40 11662 74
rect 11696 40 11730 74
rect 11764 40 11798 74
rect 11832 40 11866 74
rect 11900 40 11934 74
rect 11968 40 12002 74
rect 12036 40 12070 74
rect 12104 40 12138 74
rect 12172 40 12206 74
rect 12240 40 12274 74
rect 12308 40 12342 74
rect 12376 40 12410 74
rect 12444 40 12478 74
rect 12512 40 12546 74
rect 12580 40 12614 74
rect 12648 40 12682 74
rect 12716 40 12750 74
rect 12784 40 12818 74
rect 12852 40 12886 74
rect 12920 40 12954 74
rect 12988 40 13022 74
rect 13056 40 13090 74
rect 13124 40 13158 74
rect 13308 40 13342 74
rect 13376 40 13410 74
rect 13444 40 13478 74
rect 13512 40 13546 74
rect 13580 40 13614 74
rect 13648 40 13682 74
rect 13716 40 13750 74
rect 13784 40 13818 74
rect 13852 40 13886 74
rect 13920 40 13954 74
rect 13988 40 14022 74
rect 14056 40 14090 74
rect 14124 40 14158 74
rect 14192 40 14226 74
rect 14260 40 14294 74
rect 14328 40 14362 74
rect 14396 40 14430 74
rect 14464 40 14498 74
rect 14532 40 14566 74
rect 14600 40 14634 74
rect 14668 40 14702 74
rect 14736 40 14770 74
rect 14804 40 14838 74
rect 14872 40 14906 74
rect 11631 -189 11665 -155
rect 11699 -189 11733 -155
rect 11767 -189 11801 -155
rect 11835 -189 11869 -155
rect 11903 -189 11937 -155
rect 11971 -189 12005 -155
rect 12039 -189 12073 -155
rect 12107 -189 12141 -155
rect 12175 -189 12209 -155
rect 12243 -189 12277 -155
rect 12311 -189 12345 -155
rect 12379 -189 12413 -155
rect 12447 -189 12481 -155
rect 12515 -189 12549 -155
rect 12583 -189 12617 -155
rect 12651 -189 12685 -155
rect 12719 -189 12753 -155
rect 12787 -189 12821 -155
rect 12856 -189 12890 -155
rect 12925 -189 12959 -155
rect 12994 -189 13028 -155
rect 13063 -189 13097 -155
rect 13132 -189 13166 -155
rect 13201 -189 13235 -155
rect 13270 -189 13304 -155
rect 13339 -189 13373 -155
rect 13408 -189 13442 -155
rect 13477 -189 13511 -155
rect 13546 -189 13580 -155
rect 13615 -189 13649 -155
rect 13684 -189 13718 -155
rect 13753 -189 13787 -155
rect 13822 -189 13856 -155
rect 13891 -189 13925 -155
rect 13960 -189 13994 -155
rect 14029 -189 14063 -155
rect 14098 -189 14132 -155
rect 14167 -189 14201 -155
rect 14236 -189 14270 -155
rect 14305 -189 14339 -155
rect 14374 -189 14408 -155
rect 14443 -189 14477 -155
rect 14512 -189 14546 -155
rect 14581 -189 14615 -155
rect 14650 -189 14684 -155
rect 14719 -189 14753 -155
<< mvnsubdiffcont >>
rect 5940 2534 5974 2568
rect 5940 2466 5974 2500
rect 5940 2398 5974 2432
rect 5940 2330 5974 2364
rect 5940 2262 5974 2296
rect 5940 2194 5974 2228
rect 5940 2126 5974 2160
rect 5940 2058 5974 2092
rect 5940 1990 5974 2024
rect 5940 1922 5974 1956
rect 5940 1854 5974 1888
rect 5940 1786 5974 1820
rect 5940 1718 5974 1752
rect 5940 1650 5974 1684
rect 5940 1582 5974 1616
rect 5940 1514 5974 1548
rect 5940 1446 5974 1480
rect 5940 1378 5974 1412
rect 5940 1310 5974 1344
rect 5940 1242 5974 1276
rect 5940 1174 5974 1208
rect 5940 1106 5974 1140
rect 5940 1038 5974 1072
<< poly >>
rect 5168 2534 5234 2550
rect 5168 2500 5184 2534
rect 5218 2500 5234 2534
rect 5168 2465 5234 2500
rect 5168 2431 5184 2465
rect 5218 2431 5234 2465
rect 5168 2396 5234 2431
rect 5168 2362 5184 2396
rect 5218 2362 5234 2396
rect 5168 2327 5234 2362
rect 5168 2293 5184 2327
rect 5218 2293 5234 2327
rect 5168 2258 5234 2293
rect 5168 2224 5184 2258
rect 5218 2224 5234 2258
rect 5168 2189 5234 2224
rect 5168 2155 5184 2189
rect 5218 2155 5234 2189
rect 5168 2120 5234 2155
rect 5168 2086 5184 2120
rect 5218 2086 5234 2120
rect 5168 2051 5234 2086
rect 5168 2017 5184 2051
rect 5218 2017 5234 2051
rect 5168 1982 5234 2017
rect 5168 1948 5184 1982
rect 5218 1948 5234 1982
rect 5168 1913 5234 1948
rect 5168 1879 5184 1913
rect 5218 1879 5234 1913
rect 5168 1844 5234 1879
rect 5168 1810 5184 1844
rect 5218 1810 5234 1844
rect 5168 1776 5234 1810
rect 5168 1742 5184 1776
rect 5218 1742 5234 1776
rect 5168 1708 5234 1742
rect 5168 1674 5184 1708
rect 5218 1674 5234 1708
rect 5168 1640 5234 1674
rect 5168 1606 5184 1640
rect 5218 1606 5234 1640
rect 5168 1572 5234 1606
rect 5168 1538 5184 1572
rect 5218 1538 5234 1572
rect 5168 1504 5234 1538
rect 5168 1470 5184 1504
rect 5218 1470 5234 1504
rect 5168 1436 5234 1470
rect 5168 1402 5184 1436
rect 5218 1402 5234 1436
rect 5168 1368 5234 1402
rect 5168 1334 5184 1368
rect 5218 1334 5234 1368
rect 5168 1300 5234 1334
rect 5168 1266 5184 1300
rect 5218 1266 5234 1300
rect 5168 1232 5234 1266
rect 5168 1198 5184 1232
rect 5218 1198 5234 1232
rect 5168 1164 5234 1198
rect 5168 1130 5184 1164
rect 5218 1130 5234 1164
rect 5168 1096 5234 1130
rect 5168 1062 5184 1096
rect 5218 1062 5234 1096
rect 5168 1046 5234 1062
rect 11660 -917 14724 -901
rect 11660 -951 11676 -917
rect 11710 -951 11744 -917
rect 11778 -951 11812 -917
rect 11846 -951 11880 -917
rect 11914 -951 11948 -917
rect 11982 -951 12016 -917
rect 12050 -951 12084 -917
rect 12118 -951 12152 -917
rect 12186 -951 12220 -917
rect 12254 -951 12288 -917
rect 12322 -951 12356 -917
rect 12390 -951 12424 -917
rect 12458 -951 12492 -917
rect 12526 -951 12560 -917
rect 12594 -951 12628 -917
rect 12662 -951 12696 -917
rect 12730 -951 12764 -917
rect 12798 -951 12832 -917
rect 12866 -951 12900 -917
rect 12934 -951 12968 -917
rect 13002 -951 13036 -917
rect 13070 -951 13104 -917
rect 13138 -951 13172 -917
rect 13206 -951 13240 -917
rect 13274 -951 13308 -917
rect 13342 -951 13376 -917
rect 13410 -951 13444 -917
rect 13478 -951 13512 -917
rect 13546 -951 13580 -917
rect 13614 -951 13648 -917
rect 13682 -951 13716 -917
rect 13750 -951 13784 -917
rect 13818 -951 13852 -917
rect 13886 -951 13920 -917
rect 13954 -951 13988 -917
rect 14022 -951 14056 -917
rect 14090 -951 14124 -917
rect 14158 -951 14192 -917
rect 14226 -951 14260 -917
rect 14294 -951 14329 -917
rect 14363 -951 14398 -917
rect 14432 -951 14467 -917
rect 14501 -951 14536 -917
rect 14570 -951 14605 -917
rect 14639 -951 14674 -917
rect 14708 -951 14724 -917
rect 11660 -967 14724 -951
<< polycont >>
rect 5184 2500 5218 2534
rect 5184 2431 5218 2465
rect 5184 2362 5218 2396
rect 5184 2293 5218 2327
rect 5184 2224 5218 2258
rect 5184 2155 5218 2189
rect 5184 2086 5218 2120
rect 5184 2017 5218 2051
rect 5184 1948 5218 1982
rect 5184 1879 5218 1913
rect 5184 1810 5218 1844
rect 5184 1742 5218 1776
rect 5184 1674 5218 1708
rect 5184 1606 5218 1640
rect 5184 1538 5218 1572
rect 5184 1470 5218 1504
rect 5184 1402 5218 1436
rect 5184 1334 5218 1368
rect 5184 1266 5218 1300
rect 5184 1198 5218 1232
rect 5184 1130 5218 1164
rect 5184 1062 5218 1096
rect 11676 -951 11710 -917
rect 11744 -951 11778 -917
rect 11812 -951 11846 -917
rect 11880 -951 11914 -917
rect 11948 -951 11982 -917
rect 12016 -951 12050 -917
rect 12084 -951 12118 -917
rect 12152 -951 12186 -917
rect 12220 -951 12254 -917
rect 12288 -951 12322 -917
rect 12356 -951 12390 -917
rect 12424 -951 12458 -917
rect 12492 -951 12526 -917
rect 12560 -951 12594 -917
rect 12628 -951 12662 -917
rect 12696 -951 12730 -917
rect 12764 -951 12798 -917
rect 12832 -951 12866 -917
rect 12900 -951 12934 -917
rect 12968 -951 13002 -917
rect 13036 -951 13070 -917
rect 13104 -951 13138 -917
rect 13172 -951 13206 -917
rect 13240 -951 13274 -917
rect 13308 -951 13342 -917
rect 13376 -951 13410 -917
rect 13444 -951 13478 -917
rect 13512 -951 13546 -917
rect 13580 -951 13614 -917
rect 13648 -951 13682 -917
rect 13716 -951 13750 -917
rect 13784 -951 13818 -917
rect 13852 -951 13886 -917
rect 13920 -951 13954 -917
rect 13988 -951 14022 -917
rect 14056 -951 14090 -917
rect 14124 -951 14158 -917
rect 14192 -951 14226 -917
rect 14260 -951 14294 -917
rect 14329 -951 14363 -917
rect 14398 -951 14432 -917
rect 14467 -951 14501 -917
rect 14536 -951 14570 -917
rect 14605 -951 14639 -917
rect 14674 -951 14708 -917
<< locali >>
rect -258 38757 6154 38763
rect -258 38723 -176 38757
rect -108 38723 -99 38757
rect -40 38723 -6 38757
rect 45 38723 62 38757
rect 117 38723 130 38757
rect 189 38723 198 38757
rect 261 38723 266 38757
rect 333 38723 334 38757
rect 368 38723 371 38757
rect 436 38723 443 38757
rect 504 38723 515 38757
rect 572 38723 587 38757
rect 640 38723 659 38757
rect 708 38723 731 38757
rect 776 38723 803 38757
rect 844 38723 875 38757
rect 912 38723 946 38757
rect 981 38723 1014 38757
rect 1053 38723 1082 38757
rect 1125 38723 1150 38757
rect 1197 38723 1218 38757
rect 1269 38723 1286 38757
rect 1341 38723 1354 38757
rect 1413 38723 1422 38757
rect 1485 38723 1490 38757
rect 1557 38723 1558 38757
rect 1592 38723 1595 38757
rect 1660 38723 1667 38757
rect 1728 38723 1739 38757
rect 1796 38723 1811 38757
rect 1845 38723 1883 38757
rect 1932 38723 1955 38757
rect 2000 38723 2027 38757
rect 2068 38723 2100 38757
rect 2136 38723 2170 38757
rect 2207 38723 2238 38757
rect 2280 38723 2306 38757
rect 2353 38723 2374 38757
rect 2426 38723 2442 38757
rect 2499 38723 2510 38757
rect 2572 38723 2578 38757
rect 2645 38723 2646 38757
rect 2680 38723 2684 38757
rect 2748 38723 2757 38757
rect 2816 38723 2830 38757
rect 2884 38723 2903 38757
rect 2952 38723 2976 38757
rect 3020 38723 3049 38757
rect 3088 38723 3122 38757
rect 3156 38723 3190 38757
rect 3229 38723 3258 38757
rect 3302 38723 3326 38757
rect 3375 38723 3394 38757
rect 3448 38723 3462 38757
rect 3521 38723 3530 38757
rect 3594 38723 3598 38757
rect 3632 38723 3633 38757
rect 3700 38723 3706 38757
rect 3768 38723 3779 38757
rect 3836 38723 3852 38757
rect 3904 38723 3925 38757
rect 3959 38723 3998 38757
rect 4032 38723 4071 38757
rect 4108 38723 4142 38757
rect 4178 38723 4210 38757
rect 4251 38723 4278 38757
rect 4324 38723 4346 38757
rect 4397 38723 4414 38757
rect 4470 38723 4482 38757
rect 4543 38723 4550 38757
rect 4616 38723 4618 38757
rect 4652 38723 4655 38757
rect 4720 38723 4728 38757
rect 4788 38723 4801 38757
rect 4856 38723 4874 38757
rect 4924 38723 4947 38757
rect 4992 38723 5020 38757
rect 5060 38723 5093 38757
rect 5128 38723 5162 38757
rect 5200 38723 5230 38757
rect 5273 38723 5298 38757
rect 5346 38723 5366 38757
rect 5419 38723 5434 38757
rect 5492 38723 5502 38757
rect 5565 38723 5570 38757
rect 5672 38723 5677 38757
rect 5740 38723 5750 38757
rect 5808 38723 5823 38757
rect 5876 38723 5896 38757
rect 5944 38723 5969 38757
rect 6012 38723 6042 38757
rect 6080 38723 6154 38757
rect -258 38717 6154 38723
rect -258 38689 -212 38717
rect -258 38651 -252 38689
rect -218 38651 -212 38689
rect -258 38621 -212 38651
rect -258 38578 -252 38621
rect -218 38578 -212 38621
rect -258 38553 -212 38578
rect -258 38505 -252 38553
rect -218 38505 -212 38553
rect -258 38485 -212 38505
rect -258 38432 -252 38485
rect -218 38432 -212 38485
rect -258 38417 -212 38432
rect -258 38359 -252 38417
rect -218 38359 -212 38417
rect -258 38349 -212 38359
rect -258 38286 -252 38349
rect -218 38286 -212 38349
rect -258 38281 -212 38286
rect -258 38179 -252 38281
rect -218 38179 -212 38281
rect -258 38174 -212 38179
rect -258 38111 -252 38174
rect -218 38111 -212 38174
rect -258 38101 -212 38111
rect -258 38043 -252 38101
rect -218 38043 -212 38101
rect -258 38028 -212 38043
rect -258 37975 -252 38028
rect -218 37975 -212 38028
rect -258 37955 -212 37975
rect -258 37907 -252 37955
rect -218 37907 -212 37955
rect -258 37882 -212 37907
rect -258 37839 -252 37882
rect -218 37839 -212 37882
rect -258 37809 -212 37839
rect -258 37771 -252 37809
rect -218 37771 -212 37809
rect -258 37737 -212 37771
rect -258 37702 -252 37737
rect -218 37702 -212 37737
rect -258 37669 -212 37702
rect -258 37629 -252 37669
rect -218 37629 -212 37669
rect -258 37601 -212 37629
rect -258 37556 -252 37601
rect -218 37556 -212 37601
rect -258 37533 -212 37556
rect -258 37483 -252 37533
rect -218 37483 -212 37533
rect -258 37465 -212 37483
rect -258 37410 -252 37465
rect -218 37410 -212 37465
rect -258 37397 -212 37410
rect -258 37337 -252 37397
rect -218 37337 -212 37397
rect -258 37329 -212 37337
rect -258 37264 -252 37329
rect -218 37264 -212 37329
rect -258 37261 -212 37264
rect -258 37227 -252 37261
rect -218 37227 -212 37261
rect -258 37225 -212 37227
rect -258 37159 -252 37225
rect -218 37159 -212 37225
rect -258 37152 -212 37159
rect -258 37091 -252 37152
rect -218 37091 -212 37152
rect -258 37079 -212 37091
rect -258 37023 -252 37079
rect -218 37023 -212 37079
rect -258 37006 -212 37023
rect -258 36955 -252 37006
rect -218 36955 -212 37006
rect -258 36933 -212 36955
rect -258 36887 -252 36933
rect -218 36887 -212 36933
rect -258 36860 -212 36887
rect -258 36819 -252 36860
rect -218 36819 -212 36860
rect -258 36787 -212 36819
rect -258 36751 -252 36787
rect -218 36751 -212 36787
rect -258 36717 -212 36751
rect -258 36680 -252 36717
rect -218 36680 -212 36717
rect -258 36649 -212 36680
rect -258 36607 -252 36649
rect -218 36607 -212 36649
rect -258 36581 -212 36607
rect -258 36534 -252 36581
rect -218 36534 -212 36581
rect -258 36513 -212 36534
rect -258 36461 -252 36513
rect -218 36461 -212 36513
rect -258 36445 -212 36461
rect -258 36388 -252 36445
rect -218 36388 -212 36445
rect -258 36377 -212 36388
rect -258 36315 -252 36377
rect -218 36315 -212 36377
rect -258 36309 -212 36315
rect -258 36242 -252 36309
rect -218 36242 -212 36309
rect -258 36241 -212 36242
rect -258 36207 -252 36241
rect -218 36207 -212 36241
rect -258 36203 -212 36207
rect -258 36139 -252 36203
rect -218 36139 -212 36203
rect -258 36130 -212 36139
rect -258 36071 -252 36130
rect -218 36071 -212 36130
rect -258 36057 -212 36071
rect -258 36003 -252 36057
rect -218 36003 -212 36057
rect -258 35984 -212 36003
rect -258 35935 -252 35984
rect -218 35935 -212 35984
rect -258 35911 -212 35935
rect -258 35867 -252 35911
rect -218 35867 -212 35911
rect -258 35838 -212 35867
rect -258 35799 -252 35838
rect -218 35799 -212 35838
rect -258 35765 -212 35799
rect -258 35731 -252 35765
rect -218 35731 -212 35765
rect -258 35697 -212 35731
rect -258 35658 -252 35697
rect -218 35658 -212 35697
rect -258 35629 -212 35658
rect -258 35585 -252 35629
rect -218 35585 -212 35629
rect -258 35561 -212 35585
rect -258 35512 -252 35561
rect -218 35512 -212 35561
rect -258 35493 -212 35512
rect -258 35439 -252 35493
rect -218 35439 -212 35493
rect -258 35425 -212 35439
rect -258 35366 -252 35425
rect -218 35366 -212 35425
rect -258 35357 -212 35366
rect -258 35293 -252 35357
rect -218 35293 -212 35357
rect -258 35289 -212 35293
rect -258 35255 -252 35289
rect -218 35255 -212 35289
rect -258 35254 -212 35255
rect -258 35187 -252 35254
rect -218 35187 -212 35254
rect -258 35181 -212 35187
rect -258 35119 -252 35181
rect -218 35119 -212 35181
rect -258 35109 -212 35119
rect -258 35051 -252 35109
rect -218 35051 -212 35109
rect -258 35037 -212 35051
rect -258 34983 -252 35037
rect -218 34983 -212 35037
rect -258 34965 -212 34983
rect -258 34915 -252 34965
rect -218 34915 -212 34965
rect -258 34893 -212 34915
rect -258 34847 -252 34893
rect -218 34847 -212 34893
rect -258 34821 -212 34847
rect -258 34779 -252 34821
rect -218 34779 -212 34821
rect -258 34749 -212 34779
rect -258 34711 -252 34749
rect -218 34711 -212 34749
rect -258 34677 -212 34711
rect -258 34643 -252 34677
rect -218 34643 -212 34677
rect -258 34609 -212 34643
rect -258 34571 -252 34609
rect -218 34571 -212 34609
rect -258 34541 -212 34571
rect -258 34499 -252 34541
rect -218 34499 -212 34541
rect -258 34473 -212 34499
rect -258 34427 -252 34473
rect -218 34427 -212 34473
rect -258 34405 -212 34427
rect -258 34355 -252 34405
rect -218 34355 -212 34405
rect -258 34337 -212 34355
rect -258 34283 -252 34337
rect -218 34283 -212 34337
rect -258 34269 -212 34283
rect -258 34211 -252 34269
rect -218 34211 -212 34269
rect -258 34201 -212 34211
rect -258 34139 -252 34201
rect -218 34139 -212 34201
rect -258 34133 -212 34139
rect -258 34067 -252 34133
rect -218 34067 -212 34133
rect -258 34065 -212 34067
rect -258 34031 -252 34065
rect -218 34031 -212 34065
rect -258 34029 -212 34031
rect -258 33963 -252 34029
rect -218 33963 -212 34029
rect -258 33957 -212 33963
rect -258 33895 -252 33957
rect -218 33895 -212 33957
rect -258 33885 -212 33895
rect -258 33827 -252 33885
rect -218 33827 -212 33885
rect -258 33813 -212 33827
rect -258 33759 -252 33813
rect -218 33759 -212 33813
rect -258 33741 -212 33759
rect -258 33691 -252 33741
rect -218 33691 -212 33741
rect -258 33669 -212 33691
rect -258 33623 -252 33669
rect -218 33623 -212 33669
rect -258 33597 -212 33623
rect -258 33555 -252 33597
rect -218 33555 -212 33597
rect -258 33525 -212 33555
rect -258 33487 -252 33525
rect -218 33487 -212 33525
rect -258 33453 -212 33487
rect -258 33419 -252 33453
rect -218 33419 -212 33453
rect -258 33385 -212 33419
rect -258 33347 -252 33385
rect -218 33347 -212 33385
rect -258 33317 -212 33347
rect -258 33275 -252 33317
rect -218 33275 -212 33317
rect -258 33249 -212 33275
rect -258 33203 -252 33249
rect -218 33203 -212 33249
rect -258 33181 -212 33203
rect -258 33131 -252 33181
rect -218 33131 -212 33181
rect -258 33113 -212 33131
rect -258 33059 -252 33113
rect -218 33059 -212 33113
rect -258 33045 -212 33059
rect -258 32987 -252 33045
rect -218 32987 -212 33045
rect -258 32977 -212 32987
rect -258 32915 -252 32977
rect -218 32915 -212 32977
rect -258 32909 -212 32915
rect -258 32843 -252 32909
rect -218 32843 -212 32909
rect -258 32841 -212 32843
rect -258 32807 -252 32841
rect -218 32807 -212 32841
rect -258 32805 -212 32807
rect -258 32739 -252 32805
rect -218 32739 -212 32805
rect -258 32733 -212 32739
rect -258 32671 -252 32733
rect -218 32671 -212 32733
rect -258 32661 -212 32671
rect -258 32603 -252 32661
rect -218 32603 -212 32661
rect -258 32589 -212 32603
rect -258 32535 -252 32589
rect -218 32535 -212 32589
rect -258 32517 -212 32535
rect -258 32467 -252 32517
rect -218 32467 -212 32517
rect -258 32445 -212 32467
rect -258 32399 -252 32445
rect -218 32399 -212 32445
rect -258 32373 -212 32399
rect -258 32331 -252 32373
rect -218 32331 -212 32373
rect -258 32301 -212 32331
rect -258 32263 -252 32301
rect -218 32263 -212 32301
rect -258 32229 -212 32263
rect -258 32195 -252 32229
rect -218 32195 -212 32229
rect -258 32161 -212 32195
rect -258 32123 -252 32161
rect -218 32123 -212 32161
rect -258 32093 -212 32123
rect -258 32051 -252 32093
rect -218 32051 -212 32093
rect -258 32025 -212 32051
rect -258 31979 -252 32025
rect -218 31979 -212 32025
rect -258 31957 -212 31979
rect -258 31907 -252 31957
rect -218 31907 -212 31957
rect -258 31889 -212 31907
rect -258 31835 -252 31889
rect -218 31835 -212 31889
rect -258 31821 -212 31835
rect -258 31763 -252 31821
rect -218 31763 -212 31821
rect -258 31753 -212 31763
rect -258 31691 -252 31753
rect -218 31691 -212 31753
rect -258 31685 -212 31691
rect -258 31619 -252 31685
rect -218 31619 -212 31685
rect -258 31617 -212 31619
rect -258 31583 -252 31617
rect -218 31583 -212 31617
rect -258 31581 -212 31583
rect -258 31515 -252 31581
rect -218 31515 -212 31581
rect -258 31509 -212 31515
rect -258 31447 -252 31509
rect -218 31447 -212 31509
rect -258 31437 -212 31447
rect -258 31379 -252 31437
rect -218 31379 -212 31437
rect -258 31365 -212 31379
rect -258 31311 -252 31365
rect -218 31311 -212 31365
rect -258 31293 -212 31311
rect -258 31243 -252 31293
rect -218 31243 -212 31293
rect -258 31221 -212 31243
rect -258 31175 -252 31221
rect -218 31175 -212 31221
rect -258 31149 -212 31175
rect -258 31107 -252 31149
rect -218 31107 -212 31149
rect -258 31077 -212 31107
rect -258 31039 -252 31077
rect -218 31039 -212 31077
rect -258 31005 -212 31039
rect -258 30971 -252 31005
rect -218 30971 -212 31005
rect -258 30937 -212 30971
rect -258 30899 -252 30937
rect -218 30899 -212 30937
rect -258 30869 -212 30899
rect -258 30827 -252 30869
rect -218 30827 -212 30869
rect -258 30801 -212 30827
rect -258 30755 -252 30801
rect -218 30755 -212 30801
rect -258 30733 -212 30755
rect -258 30683 -252 30733
rect -218 30683 -212 30733
rect -258 30665 -212 30683
rect -258 30611 -252 30665
rect -218 30611 -212 30665
rect -258 30597 -212 30611
rect -258 30539 -252 30597
rect -218 30539 -212 30597
rect -258 30529 -212 30539
rect -258 30467 -252 30529
rect -218 30467 -212 30529
rect -258 30461 -212 30467
rect -258 30395 -252 30461
rect -218 30395 -212 30461
rect -258 30393 -212 30395
rect -258 30359 -252 30393
rect -218 30359 -212 30393
rect -258 30357 -212 30359
rect -258 30291 -252 30357
rect -218 30291 -212 30357
rect -258 30285 -212 30291
rect -258 30223 -252 30285
rect -218 30223 -212 30285
rect -258 30213 -212 30223
rect -258 30155 -252 30213
rect -218 30155 -212 30213
rect -258 30141 -212 30155
rect -258 30087 -252 30141
rect -218 30087 -212 30141
rect -258 30069 -212 30087
rect -258 30019 -252 30069
rect -218 30019 -212 30069
rect -258 29997 -212 30019
rect -258 29951 -252 29997
rect -218 29951 -212 29997
rect -258 29925 -212 29951
rect -258 29883 -252 29925
rect -218 29883 -212 29925
rect -258 29853 -212 29883
rect -258 29815 -252 29853
rect -218 29815 -212 29853
rect -258 29781 -212 29815
rect -258 29747 -252 29781
rect -218 29747 -212 29781
rect -258 29713 -212 29747
rect -258 29675 -252 29713
rect -218 29675 -212 29713
rect -258 29645 -212 29675
rect -258 29603 -252 29645
rect -218 29603 -212 29645
rect -258 29577 -212 29603
rect -258 29531 -252 29577
rect -218 29531 -212 29577
rect -258 29509 -212 29531
rect -258 29459 -252 29509
rect -218 29459 -212 29509
rect -258 29441 -212 29459
rect -258 29387 -252 29441
rect -218 29387 -212 29441
rect -258 29373 -212 29387
rect -258 29315 -252 29373
rect -218 29315 -212 29373
rect -258 29305 -212 29315
rect -258 29243 -252 29305
rect -218 29243 -212 29305
rect -258 29237 -212 29243
rect -258 29171 -252 29237
rect -218 29171 -212 29237
rect -258 29169 -212 29171
rect -258 29135 -252 29169
rect -218 29135 -212 29169
rect -258 29133 -212 29135
rect -258 29067 -252 29133
rect -218 29067 -212 29133
rect -258 29061 -212 29067
rect -258 28999 -252 29061
rect -218 28999 -212 29061
rect -258 28989 -212 28999
rect -258 28931 -252 28989
rect -218 28931 -212 28989
rect -258 28917 -212 28931
rect -258 28863 -252 28917
rect -218 28863 -212 28917
rect -258 28845 -212 28863
rect -258 28795 -252 28845
rect -218 28795 -212 28845
rect -258 28773 -212 28795
rect -258 28727 -252 28773
rect -218 28727 -212 28773
rect -258 28701 -212 28727
rect -258 28659 -252 28701
rect -218 28659 -212 28701
rect -258 28629 -212 28659
rect -258 28591 -252 28629
rect -218 28591 -212 28629
rect -258 28557 -212 28591
rect -258 28523 -252 28557
rect -218 28523 -212 28557
rect -258 28489 -212 28523
rect -258 28451 -252 28489
rect -218 28451 -212 28489
rect -258 28421 -212 28451
rect -258 28379 -252 28421
rect -218 28379 -212 28421
rect -258 28353 -212 28379
rect -258 28307 -252 28353
rect -218 28307 -212 28353
rect -258 28285 -212 28307
rect -258 28235 -252 28285
rect -218 28235 -212 28285
rect -258 28217 -212 28235
rect -258 28163 -252 28217
rect -218 28163 -212 28217
rect -258 28149 -212 28163
rect -258 28091 -252 28149
rect -218 28091 -212 28149
rect -258 28081 -212 28091
rect -258 28019 -252 28081
rect -218 28019 -212 28081
rect -258 28013 -212 28019
rect -258 27947 -252 28013
rect -218 27947 -212 28013
rect -258 27945 -212 27947
rect -258 27911 -252 27945
rect -218 27911 -212 27945
rect -258 27909 -212 27911
rect -258 27843 -252 27909
rect -218 27843 -212 27909
rect -258 27837 -212 27843
rect -258 27775 -252 27837
rect -218 27775 -212 27837
rect -258 27765 -212 27775
rect -258 27707 -252 27765
rect -218 27707 -212 27765
rect -258 27693 -212 27707
rect -258 27639 -252 27693
rect -218 27639 -212 27693
rect -258 27621 -212 27639
rect -258 27571 -252 27621
rect -218 27571 -212 27621
rect -258 27549 -212 27571
rect -258 27503 -252 27549
rect -218 27503 -212 27549
rect -258 27477 -212 27503
rect -258 27435 -252 27477
rect -218 27435 -212 27477
rect -258 27405 -212 27435
rect -258 27367 -252 27405
rect -218 27367 -212 27405
rect -258 27333 -212 27367
rect -258 27299 -252 27333
rect -218 27299 -212 27333
rect -258 27265 -212 27299
rect -258 27227 -252 27265
rect -218 27227 -212 27265
rect -258 27197 -212 27227
rect -258 27155 -252 27197
rect -218 27155 -212 27197
rect -258 27129 -212 27155
rect -258 27083 -252 27129
rect -218 27083 -212 27129
rect -258 27061 -212 27083
rect -258 27011 -252 27061
rect -218 27011 -212 27061
rect -258 26993 -212 27011
rect -258 26939 -252 26993
rect -218 26939 -212 26993
rect -258 26925 -212 26939
rect -258 26867 -252 26925
rect -218 26867 -212 26925
rect -258 26857 -212 26867
rect -258 26795 -252 26857
rect -218 26795 -212 26857
rect -258 26789 -212 26795
rect -258 26723 -252 26789
rect -218 26723 -212 26789
rect -258 26721 -212 26723
rect -258 26687 -252 26721
rect -218 26687 -212 26721
rect -258 26685 -212 26687
rect -258 26619 -252 26685
rect -218 26619 -212 26685
rect -258 26613 -212 26619
rect -258 26551 -252 26613
rect -218 26551 -212 26613
rect -258 26541 -212 26551
rect -258 26483 -252 26541
rect -218 26483 -212 26541
rect -258 26469 -212 26483
rect -258 26415 -252 26469
rect -218 26415 -212 26469
rect -258 26397 -212 26415
rect -258 26347 -252 26397
rect -218 26347 -212 26397
rect -258 26325 -212 26347
rect -258 26279 -252 26325
rect -218 26279 -212 26325
rect -258 26253 -212 26279
rect -258 26211 -252 26253
rect -218 26211 -212 26253
rect -258 26181 -212 26211
rect -258 26143 -252 26181
rect -218 26143 -212 26181
rect -258 26109 -212 26143
rect -258 26075 -252 26109
rect -218 26075 -212 26109
rect -258 26041 -212 26075
rect -258 26003 -252 26041
rect -218 26003 -212 26041
rect -258 25973 -212 26003
rect -258 25931 -252 25973
rect -218 25931 -212 25973
rect -258 25905 -212 25931
rect -258 25859 -252 25905
rect -218 25859 -212 25905
rect -258 25837 -212 25859
rect -258 25787 -252 25837
rect -218 25787 -212 25837
rect -258 25769 -212 25787
rect -258 25715 -252 25769
rect -218 25715 -212 25769
rect -258 25701 -212 25715
rect -258 25643 -252 25701
rect -218 25643 -212 25701
rect -258 25633 -212 25643
rect -258 25571 -252 25633
rect -218 25571 -212 25633
rect -258 25565 -212 25571
rect -258 25499 -252 25565
rect -218 25499 -212 25565
rect -258 25497 -212 25499
rect -258 25463 -252 25497
rect -218 25463 -212 25497
rect -258 25461 -212 25463
rect -258 25395 -252 25461
rect -218 25395 -212 25461
rect -258 25389 -212 25395
rect -258 25327 -252 25389
rect -218 25327 -212 25389
rect -258 25317 -212 25327
rect -258 25259 -252 25317
rect -218 25259 -212 25317
rect -258 25245 -212 25259
rect -258 25191 -252 25245
rect -218 25191 -212 25245
rect -258 25173 -212 25191
rect -258 25123 -252 25173
rect -218 25123 -212 25173
rect -258 25101 -212 25123
rect -258 25055 -252 25101
rect -218 25055 -212 25101
rect -258 25029 -212 25055
rect -258 24987 -252 25029
rect -218 24987 -212 25029
rect -258 24957 -212 24987
rect -258 24919 -252 24957
rect -218 24919 -212 24957
rect -258 24885 -212 24919
rect -258 24851 -252 24885
rect -218 24851 -212 24885
rect -258 24817 -212 24851
rect -258 24779 -252 24817
rect -218 24779 -212 24817
rect -258 24749 -212 24779
rect -258 24707 -252 24749
rect -218 24707 -212 24749
rect -258 24681 -212 24707
rect -258 24635 -252 24681
rect -218 24635 -212 24681
rect -258 24613 -212 24635
rect -258 24563 -252 24613
rect -218 24563 -212 24613
rect -258 24545 -212 24563
rect -258 24491 -252 24545
rect -218 24491 -212 24545
rect -258 24477 -212 24491
rect -258 24419 -252 24477
rect -218 24419 -212 24477
rect -258 24409 -212 24419
rect -258 24347 -252 24409
rect -218 24347 -212 24409
rect -258 24341 -212 24347
rect -258 24275 -252 24341
rect -218 24275 -212 24341
rect -258 24273 -212 24275
rect -258 24239 -252 24273
rect -218 24239 -212 24273
rect -258 24237 -212 24239
rect -258 24171 -252 24237
rect -218 24171 -212 24237
rect -258 24165 -212 24171
rect -258 24103 -252 24165
rect -218 24103 -212 24165
rect -258 24093 -212 24103
rect -258 24035 -252 24093
rect -218 24035 -212 24093
rect -258 24021 -212 24035
rect -258 23967 -252 24021
rect -218 23967 -212 24021
rect -258 23949 -212 23967
rect -258 23899 -252 23949
rect -218 23899 -212 23949
rect -258 23877 -212 23899
rect -258 23831 -252 23877
rect -218 23831 -212 23877
rect -258 23805 -212 23831
rect -258 23763 -252 23805
rect -218 23763 -212 23805
rect -258 23733 -212 23763
rect -258 23695 -252 23733
rect -218 23695 -212 23733
rect -258 23661 -212 23695
rect -258 23627 -252 23661
rect -218 23627 -212 23661
rect -258 23593 -212 23627
rect -258 23555 -252 23593
rect -218 23555 -212 23593
rect -258 23525 -212 23555
rect -258 23483 -252 23525
rect -218 23483 -212 23525
rect -258 23457 -212 23483
rect -258 23411 -252 23457
rect -218 23411 -212 23457
rect -258 23389 -212 23411
rect -258 23339 -252 23389
rect -218 23339 -212 23389
rect -258 23321 -212 23339
rect -258 23267 -252 23321
rect -218 23267 -212 23321
rect -258 23253 -212 23267
rect -258 23195 -252 23253
rect -218 23195 -212 23253
rect -258 23185 -212 23195
rect -258 23123 -252 23185
rect -218 23123 -212 23185
rect -258 23117 -212 23123
rect -258 23051 -252 23117
rect -218 23051 -212 23117
rect -258 23049 -212 23051
rect -258 23015 -252 23049
rect -218 23015 -212 23049
rect -258 23013 -212 23015
rect -258 22947 -252 23013
rect -218 22947 -212 23013
rect -258 22941 -212 22947
rect -258 22879 -252 22941
rect -218 22879 -212 22941
rect -258 22869 -212 22879
rect -258 22811 -252 22869
rect -218 22811 -212 22869
rect -258 22797 -212 22811
rect -258 22743 -252 22797
rect -218 22743 -212 22797
rect -258 22725 -212 22743
rect -258 22675 -252 22725
rect -218 22675 -212 22725
rect -258 22653 -212 22675
rect -258 22607 -252 22653
rect -218 22607 -212 22653
rect -258 22581 -212 22607
rect -258 22539 -252 22581
rect -218 22539 -212 22581
rect -258 22509 -212 22539
rect -258 22471 -252 22509
rect -218 22471 -212 22509
rect -258 22437 -212 22471
rect -258 22403 -252 22437
rect -218 22403 -212 22437
rect -258 22369 -212 22403
rect -258 22331 -252 22369
rect -218 22331 -212 22369
rect -258 22301 -212 22331
rect -258 22259 -252 22301
rect -218 22259 -212 22301
rect -258 22233 -212 22259
rect -258 22187 -252 22233
rect -218 22187 -212 22233
rect -258 22165 -212 22187
rect -258 22115 -252 22165
rect -218 22115 -212 22165
rect -258 22097 -212 22115
rect -258 22043 -252 22097
rect -218 22043 -212 22097
rect -258 22029 -212 22043
rect -258 21971 -252 22029
rect -218 21971 -212 22029
rect -258 21961 -212 21971
rect -258 21899 -252 21961
rect -218 21899 -212 21961
rect -258 21893 -212 21899
rect -258 21827 -252 21893
rect -218 21827 -212 21893
rect -258 21825 -212 21827
rect -258 21791 -252 21825
rect -218 21791 -212 21825
rect -258 21789 -212 21791
rect -258 21723 -252 21789
rect -218 21723 -212 21789
rect -258 21717 -212 21723
rect -258 21655 -252 21717
rect -218 21655 -212 21717
rect -258 21645 -212 21655
rect -258 21587 -252 21645
rect -218 21587 -212 21645
rect -258 21573 -212 21587
rect -258 21519 -252 21573
rect -218 21519 -212 21573
rect -258 21501 -212 21519
rect -258 21451 -252 21501
rect -218 21451 -212 21501
rect -258 21429 -212 21451
rect -258 21383 -252 21429
rect -218 21383 -212 21429
rect -258 21357 -212 21383
rect -258 21315 -252 21357
rect -218 21315 -212 21357
rect -258 21285 -212 21315
rect -258 21247 -252 21285
rect -218 21247 -212 21285
rect -258 21213 -212 21247
rect -258 21179 -252 21213
rect -218 21179 -212 21213
rect -258 21145 -212 21179
rect -258 21107 -252 21145
rect -218 21107 -212 21145
rect -258 21077 -212 21107
rect -258 21035 -252 21077
rect -218 21035 -212 21077
rect -258 21009 -212 21035
rect -258 20963 -252 21009
rect -218 20963 -212 21009
rect -258 20941 -212 20963
rect -258 20891 -252 20941
rect -218 20891 -212 20941
rect -258 20873 -212 20891
rect -258 20819 -252 20873
rect -218 20819 -212 20873
rect -258 20805 -212 20819
rect -258 20747 -252 20805
rect -218 20747 -212 20805
rect -258 20737 -212 20747
rect -258 20675 -252 20737
rect -218 20675 -212 20737
rect -258 20669 -212 20675
rect -258 20603 -252 20669
rect -218 20603 -212 20669
rect -258 20601 -212 20603
rect -258 20567 -252 20601
rect -218 20567 -212 20601
rect -258 20565 -212 20567
rect -258 20499 -252 20565
rect -218 20499 -212 20565
rect -258 20493 -212 20499
rect -258 20431 -252 20493
rect -218 20431 -212 20493
rect -258 20421 -212 20431
rect -258 20363 -252 20421
rect -218 20363 -212 20421
rect -258 20349 -212 20363
rect -258 20295 -252 20349
rect -218 20295 -212 20349
rect -258 20277 -212 20295
rect -258 20227 -252 20277
rect -218 20227 -212 20277
rect -258 20205 -212 20227
rect -258 20159 -252 20205
rect -218 20159 -212 20205
rect -258 20133 -212 20159
rect -258 20091 -252 20133
rect -218 20091 -212 20133
rect -258 20061 -212 20091
rect -258 20023 -252 20061
rect -218 20023 -212 20061
rect -258 19989 -212 20023
rect -258 19955 -252 19989
rect -218 19955 -212 19989
rect -258 19921 -212 19955
rect -258 19883 -252 19921
rect -218 19883 -212 19921
rect -258 19853 -212 19883
rect -258 19811 -252 19853
rect -218 19811 -212 19853
rect -258 19785 -212 19811
rect -258 19739 -252 19785
rect -218 19739 -212 19785
rect -258 19717 -212 19739
rect -258 19667 -252 19717
rect -218 19667 -212 19717
rect -258 19649 -212 19667
rect -258 19595 -252 19649
rect -218 19595 -212 19649
rect -258 19581 -212 19595
rect -258 19523 -252 19581
rect -218 19523 -212 19581
rect -258 19513 -212 19523
rect -258 19451 -252 19513
rect -218 19451 -212 19513
rect -258 19445 -212 19451
rect -258 19379 -252 19445
rect -218 19379 -212 19445
rect -258 19377 -212 19379
rect -258 19343 -252 19377
rect -218 19343 -212 19377
rect -258 19341 -212 19343
rect -258 19275 -252 19341
rect -218 19275 -212 19341
rect -258 19269 -212 19275
rect -258 19207 -252 19269
rect -218 19207 -212 19269
rect -258 19197 -212 19207
rect -258 19139 -252 19197
rect -218 19139 -212 19197
rect -258 19125 -212 19139
rect -258 19071 -252 19125
rect -218 19071 -212 19125
rect -258 19053 -212 19071
rect -258 19003 -252 19053
rect -218 19003 -212 19053
rect -258 18981 -212 19003
rect -258 18935 -252 18981
rect -218 18935 -212 18981
rect -258 18909 -212 18935
rect -258 18867 -252 18909
rect -218 18867 -212 18909
rect -258 18837 -212 18867
rect -258 18799 -252 18837
rect -218 18799 -212 18837
rect -258 18765 -212 18799
rect -258 18731 -252 18765
rect -218 18731 -212 18765
rect -258 18697 -212 18731
rect -258 18659 -252 18697
rect -218 18659 -212 18697
rect -258 18629 -212 18659
rect -258 18587 -252 18629
rect -218 18587 -212 18629
rect -258 18561 -212 18587
rect -258 18515 -252 18561
rect -218 18515 -212 18561
rect -258 18493 -212 18515
rect -258 18443 -252 18493
rect -218 18443 -212 18493
rect -258 18425 -212 18443
rect -258 18371 -252 18425
rect -218 18371 -212 18425
rect -258 18357 -212 18371
rect -258 18299 -252 18357
rect -218 18299 -212 18357
rect -258 18289 -212 18299
rect -258 18227 -252 18289
rect -218 18227 -212 18289
rect -258 18221 -212 18227
rect -258 18155 -252 18221
rect -218 18155 -212 18221
rect -258 18153 -212 18155
rect -258 18119 -252 18153
rect -218 18119 -212 18153
rect -258 18117 -212 18119
rect -258 18051 -252 18117
rect -218 18051 -212 18117
rect -258 18045 -212 18051
rect -258 17983 -252 18045
rect -218 17983 -212 18045
rect -258 17973 -212 17983
rect -258 17915 -252 17973
rect -218 17915 -212 17973
rect -258 17901 -212 17915
rect -258 17847 -252 17901
rect -218 17847 -212 17901
rect -258 17829 -212 17847
rect -258 17779 -252 17829
rect -218 17779 -212 17829
rect -258 17757 -212 17779
rect -258 17711 -252 17757
rect -218 17711 -212 17757
rect -258 17685 -212 17711
rect -258 17643 -252 17685
rect -218 17643 -212 17685
rect -258 17613 -212 17643
rect -258 17575 -252 17613
rect -218 17575 -212 17613
rect -258 17541 -212 17575
rect -258 17507 -252 17541
rect -218 17507 -212 17541
rect -258 17473 -212 17507
rect -258 17435 -252 17473
rect -218 17435 -212 17473
rect -258 17405 -212 17435
rect -258 17363 -252 17405
rect -218 17363 -212 17405
rect -258 17337 -212 17363
rect -258 17291 -252 17337
rect -218 17291 -212 17337
rect -258 17269 -212 17291
rect -258 17219 -252 17269
rect -218 17219 -212 17269
rect -258 17201 -212 17219
rect -258 17147 -252 17201
rect -218 17147 -212 17201
rect -258 17133 -212 17147
rect -258 17075 -252 17133
rect -218 17075 -212 17133
rect -258 17065 -212 17075
rect -258 17003 -252 17065
rect -218 17003 -212 17065
rect -258 16997 -212 17003
rect -258 16931 -252 16997
rect -218 16931 -212 16997
rect -258 16929 -212 16931
rect -258 16895 -252 16929
rect -218 16895 -212 16929
rect -258 16893 -212 16895
rect -258 16827 -252 16893
rect -218 16827 -212 16893
rect -258 16821 -212 16827
rect -258 16759 -252 16821
rect -218 16759 -212 16821
rect -258 16749 -212 16759
rect -258 16691 -252 16749
rect -218 16691 -212 16749
rect -258 16677 -212 16691
rect -258 16623 -252 16677
rect -218 16623 -212 16677
rect -258 16605 -212 16623
rect -258 16555 -252 16605
rect -218 16555 -212 16605
rect -258 16533 -212 16555
rect -258 16487 -252 16533
rect -218 16487 -212 16533
rect -258 16461 -212 16487
rect -258 16419 -252 16461
rect -218 16419 -212 16461
rect -258 16389 -212 16419
rect -258 16351 -252 16389
rect -218 16351 -212 16389
rect -258 16317 -212 16351
rect -258 16283 -252 16317
rect -218 16283 -212 16317
rect -258 16249 -212 16283
rect -258 16211 -252 16249
rect -218 16211 -212 16249
rect -258 16181 -212 16211
rect -258 16139 -252 16181
rect -218 16139 -212 16181
rect -258 16113 -212 16139
rect -258 16067 -252 16113
rect -218 16067 -212 16113
rect -258 16045 -212 16067
rect -258 15995 -252 16045
rect -218 15995 -212 16045
rect -258 15977 -212 15995
rect -258 15923 -252 15977
rect -218 15923 -212 15977
rect -258 15909 -212 15923
rect -258 15851 -252 15909
rect -218 15851 -212 15909
rect -258 15841 -212 15851
rect -258 15779 -252 15841
rect -218 15779 -212 15841
rect -258 15773 -212 15779
rect -258 15707 -252 15773
rect -218 15707 -212 15773
rect -258 15705 -212 15707
rect -258 15671 -252 15705
rect -218 15671 -212 15705
rect -258 15669 -212 15671
rect -258 15603 -252 15669
rect -218 15603 -212 15669
rect -258 15597 -212 15603
rect -258 15535 -252 15597
rect -218 15535 -212 15597
rect -258 15525 -212 15535
rect -258 15467 -252 15525
rect -218 15467 -212 15525
rect -258 15453 -212 15467
rect -258 15399 -252 15453
rect -218 15399 -212 15453
rect -258 15381 -212 15399
rect -258 15331 -252 15381
rect -218 15331 -212 15381
rect -258 15309 -212 15331
rect -258 15263 -252 15309
rect -218 15263 -212 15309
rect -258 15237 -212 15263
rect -258 15195 -252 15237
rect -218 15195 -212 15237
rect -258 15165 -212 15195
rect -258 15127 -252 15165
rect -218 15127 -212 15165
rect -258 15093 -212 15127
rect -258 15059 -252 15093
rect -218 15059 -212 15093
rect -258 15025 -212 15059
rect -258 14987 -252 15025
rect -218 14987 -212 15025
rect -258 14957 -212 14987
rect -258 14915 -252 14957
rect -218 14915 -212 14957
rect -258 14889 -212 14915
rect -258 14843 -252 14889
rect -218 14843 -212 14889
rect -258 14821 -212 14843
rect -258 14771 -252 14821
rect -218 14771 -212 14821
rect -258 14753 -212 14771
rect -258 14699 -252 14753
rect -218 14699 -212 14753
rect -258 14685 -212 14699
rect -258 14627 -252 14685
rect -218 14627 -212 14685
rect -258 14617 -212 14627
rect -258 14555 -252 14617
rect -218 14555 -212 14617
rect -258 14549 -212 14555
rect -258 14483 -252 14549
rect -218 14483 -212 14549
rect -258 14481 -212 14483
rect -258 14447 -252 14481
rect -218 14447 -212 14481
rect -258 14445 -212 14447
rect -258 14379 -252 14445
rect -218 14379 -212 14445
rect -258 14373 -212 14379
rect -258 14311 -252 14373
rect -218 14311 -212 14373
rect -258 14301 -212 14311
rect -258 14243 -252 14301
rect -218 14243 -212 14301
rect -258 14229 -212 14243
rect -258 14175 -252 14229
rect -218 14175 -212 14229
rect -258 14157 -212 14175
rect -258 14107 -252 14157
rect -218 14107 -212 14157
rect -258 14085 -212 14107
rect -258 14039 -252 14085
rect -218 14039 -212 14085
rect -258 14013 -212 14039
rect -258 13971 -252 14013
rect -218 13971 -212 14013
rect -258 13941 -212 13971
rect -258 13903 -252 13941
rect -218 13903 -212 13941
rect -258 13869 -212 13903
rect -258 13835 -252 13869
rect -218 13835 -212 13869
rect -258 13801 -212 13835
rect -258 13763 -252 13801
rect -218 13763 -212 13801
rect -258 13733 -212 13763
rect -258 13691 -252 13733
rect -218 13691 -212 13733
rect -258 13665 -212 13691
rect -258 13619 -252 13665
rect -218 13619 -212 13665
rect -258 13597 -212 13619
rect -258 13547 -252 13597
rect -218 13547 -212 13597
rect -258 13529 -212 13547
rect -258 13475 -252 13529
rect -218 13475 -212 13529
rect -258 13461 -212 13475
rect -258 13403 -252 13461
rect -218 13403 -212 13461
rect -258 13393 -212 13403
rect -258 13331 -252 13393
rect -218 13331 -212 13393
rect -258 13325 -212 13331
rect -258 13259 -252 13325
rect -218 13259 -212 13325
rect -258 13257 -212 13259
rect -258 13223 -252 13257
rect -218 13223 -212 13257
rect -258 13221 -212 13223
rect -258 13155 -252 13221
rect -218 13155 -212 13221
rect -258 13149 -212 13155
rect -258 13087 -252 13149
rect -218 13087 -212 13149
rect -258 13077 -212 13087
rect -258 13019 -252 13077
rect -218 13019 -212 13077
rect -258 13005 -212 13019
rect -258 12951 -252 13005
rect -218 12951 -212 13005
rect -258 12933 -212 12951
rect -258 12883 -252 12933
rect -218 12883 -212 12933
rect -258 12861 -212 12883
rect -258 12815 -252 12861
rect -218 12815 -212 12861
rect -258 12789 -212 12815
rect -258 12747 -252 12789
rect -218 12747 -212 12789
rect -258 12717 -212 12747
rect -258 12679 -252 12717
rect -218 12679 -212 12717
rect -258 12645 -212 12679
rect -258 12611 -252 12645
rect -218 12611 -212 12645
rect -258 12577 -212 12611
rect -258 12539 -252 12577
rect -218 12539 -212 12577
rect -258 12509 -212 12539
rect -258 12467 -252 12509
rect -218 12467 -212 12509
rect -258 12441 -212 12467
rect -258 12395 -252 12441
rect -218 12395 -212 12441
rect -258 12373 -212 12395
rect -258 12323 -252 12373
rect -218 12323 -212 12373
rect -258 12305 -212 12323
rect -258 12251 -252 12305
rect -218 12251 -212 12305
rect -258 12237 -212 12251
rect -258 12179 -252 12237
rect -218 12179 -212 12237
rect -258 12169 -212 12179
rect -258 12107 -252 12169
rect -218 12107 -212 12169
rect -258 12101 -212 12107
rect -258 12035 -252 12101
rect -218 12035 -212 12101
rect -258 12033 -212 12035
rect -258 11999 -252 12033
rect -218 11999 -212 12033
rect -258 11997 -212 11999
rect -258 11931 -252 11997
rect -218 11931 -212 11997
rect -258 11925 -212 11931
rect -258 11863 -252 11925
rect -218 11863 -212 11925
rect -258 11853 -212 11863
rect -258 11795 -252 11853
rect -218 11795 -212 11853
rect -258 11781 -212 11795
rect -258 11727 -252 11781
rect -218 11727 -212 11781
rect -258 11709 -212 11727
rect -258 11659 -252 11709
rect -218 11659 -212 11709
rect -258 11637 -212 11659
rect -258 11591 -252 11637
rect -218 11591 -212 11637
rect -258 11565 -212 11591
rect -258 11523 -252 11565
rect -218 11523 -212 11565
rect -258 11493 -212 11523
rect -258 11455 -252 11493
rect -218 11455 -212 11493
rect -258 11421 -212 11455
rect -258 11387 -252 11421
rect -218 11387 -212 11421
rect -258 11353 -212 11387
rect -258 11315 -252 11353
rect -218 11315 -212 11353
rect -258 11285 -212 11315
rect -258 11243 -252 11285
rect -218 11243 -212 11285
rect -258 11217 -212 11243
rect -258 11171 -252 11217
rect -218 11171 -212 11217
rect -258 11149 -212 11171
rect -258 11099 -252 11149
rect -218 11099 -212 11149
rect -258 11081 -212 11099
rect -258 11027 -252 11081
rect -218 11027 -212 11081
rect -258 11013 -212 11027
rect -258 10955 -252 11013
rect -218 10955 -212 11013
rect -258 10945 -212 10955
rect -258 10883 -252 10945
rect -218 10883 -212 10945
rect -258 10877 -212 10883
rect -258 10811 -252 10877
rect -218 10811 -212 10877
rect -258 10809 -212 10811
rect -258 10775 -252 10809
rect -218 10775 -212 10809
rect -258 10773 -212 10775
rect -258 10707 -252 10773
rect -218 10707 -212 10773
rect -258 10701 -212 10707
rect -258 10639 -252 10701
rect -218 10639 -212 10701
rect -258 10629 -212 10639
rect -258 10571 -252 10629
rect -218 10571 -212 10629
rect -258 10557 -212 10571
rect -258 10503 -252 10557
rect -218 10503 -212 10557
rect -258 10485 -212 10503
rect -258 10435 -252 10485
rect -218 10435 -212 10485
rect -258 10413 -212 10435
rect -258 10367 -252 10413
rect -218 10367 -212 10413
rect -258 10341 -212 10367
rect -258 10299 -252 10341
rect -218 10299 -212 10341
rect -258 10269 -212 10299
rect -258 10231 -252 10269
rect -218 10231 -212 10269
rect -258 10197 -212 10231
rect -258 10163 -252 10197
rect -218 10163 -212 10197
rect -258 10129 -212 10163
rect -258 10091 -252 10129
rect -218 10091 -212 10129
rect -258 10061 -212 10091
rect -258 10019 -252 10061
rect -218 10019 -212 10061
rect -258 9993 -212 10019
rect -258 9947 -252 9993
rect -218 9947 -212 9993
rect -258 9925 -212 9947
rect -258 9875 -252 9925
rect -218 9875 -212 9925
rect -258 9857 -212 9875
rect -258 9803 -252 9857
rect -218 9803 -212 9857
rect -258 9789 -212 9803
rect -258 9731 -252 9789
rect -218 9731 -212 9789
rect -258 9721 -212 9731
rect -258 9659 -252 9721
rect -218 9659 -212 9721
rect -258 9653 -212 9659
rect -258 9587 -252 9653
rect -218 9587 -212 9653
rect -258 9585 -212 9587
rect -258 9551 -252 9585
rect -218 9551 -212 9585
rect -258 9549 -212 9551
rect -258 9483 -252 9549
rect -218 9483 -212 9549
rect -258 9477 -212 9483
rect -258 9415 -252 9477
rect -218 9415 -212 9477
rect -258 9405 -212 9415
rect -258 9347 -252 9405
rect -218 9347 -212 9405
rect -258 9333 -212 9347
rect -258 9279 -252 9333
rect -218 9279 -212 9333
rect -258 9261 -212 9279
rect -258 9211 -252 9261
rect -218 9211 -212 9261
rect -258 9189 -212 9211
rect -258 9143 -252 9189
rect -218 9143 -212 9189
rect -258 9117 -212 9143
rect -258 9075 -252 9117
rect -218 9075 -212 9117
rect -258 9045 -212 9075
rect -258 9007 -252 9045
rect -218 9007 -212 9045
rect -258 8973 -212 9007
rect -258 8939 -252 8973
rect -218 8939 -212 8973
rect -258 8905 -212 8939
rect -258 8867 -252 8905
rect -218 8867 -212 8905
rect -258 8837 -212 8867
rect -258 8795 -252 8837
rect -218 8795 -212 8837
rect -258 8769 -212 8795
rect -258 8723 -252 8769
rect -218 8723 -212 8769
rect -258 8701 -212 8723
rect -258 8651 -252 8701
rect -218 8651 -212 8701
rect -258 8633 -212 8651
rect -258 8579 -252 8633
rect -218 8579 -212 8633
rect -258 8565 -212 8579
rect -258 8507 -252 8565
rect -218 8507 -212 8565
rect -258 8497 -212 8507
rect -258 8435 -252 8497
rect -218 8435 -212 8497
rect -258 8429 -212 8435
rect -258 8363 -252 8429
rect -218 8363 -212 8429
rect -258 8361 -212 8363
rect -258 8327 -252 8361
rect -218 8327 -212 8361
rect -258 8325 -212 8327
rect -258 8259 -252 8325
rect -218 8259 -212 8325
rect -258 8253 -212 8259
rect -258 8191 -252 8253
rect -218 8191 -212 8253
rect -258 8181 -212 8191
rect -258 8123 -252 8181
rect -218 8123 -212 8181
rect -258 8109 -212 8123
rect -258 8055 -252 8109
rect -218 8055 -212 8109
rect -258 8037 -212 8055
rect -258 7987 -252 8037
rect -218 7987 -212 8037
rect -258 7965 -212 7987
rect -258 7919 -252 7965
rect -218 7919 -212 7965
rect -258 7893 -212 7919
rect -258 7851 -252 7893
rect -218 7851 -212 7893
rect -258 7821 -212 7851
rect -258 7783 -252 7821
rect -218 7783 -212 7821
rect -258 7749 -212 7783
rect -258 7715 -252 7749
rect -218 7715 -212 7749
rect -258 7681 -212 7715
rect -258 7643 -252 7681
rect -218 7643 -212 7681
rect -258 7613 -212 7643
rect -258 7571 -252 7613
rect -218 7571 -212 7613
rect -258 7545 -212 7571
rect -258 7499 -252 7545
rect -218 7499 -212 7545
rect -258 7477 -212 7499
rect -258 7427 -252 7477
rect -218 7427 -212 7477
rect -258 7409 -212 7427
rect -258 7355 -252 7409
rect -218 7355 -212 7409
rect -258 7341 -212 7355
rect -258 7283 -252 7341
rect -218 7283 -212 7341
rect -258 7273 -212 7283
rect -258 7211 -252 7273
rect -218 7211 -212 7273
rect -258 7205 -212 7211
rect -258 7139 -252 7205
rect -218 7139 -212 7205
rect -258 7137 -212 7139
rect -258 7103 -252 7137
rect -218 7103 -212 7137
rect -258 7101 -212 7103
rect -258 7035 -252 7101
rect -218 7035 -212 7101
rect -258 7029 -212 7035
rect -258 6967 -252 7029
rect -218 6967 -212 7029
rect -258 6957 -212 6967
rect -258 6899 -252 6957
rect -218 6899 -212 6957
rect -258 6885 -212 6899
rect -258 6831 -252 6885
rect -218 6831 -212 6885
rect -258 6813 -212 6831
rect -258 6763 -252 6813
rect -218 6763 -212 6813
rect -258 6741 -212 6763
rect -258 6695 -252 6741
rect -218 6695 -212 6741
rect -258 6669 -212 6695
rect -258 6627 -252 6669
rect -218 6627 -212 6669
rect -258 6597 -212 6627
rect -258 6559 -252 6597
rect -218 6559 -212 6597
rect -258 6525 -212 6559
rect -258 6491 -252 6525
rect -218 6491 -212 6525
rect -258 6457 -212 6491
rect -258 6419 -252 6457
rect -218 6419 -212 6457
rect -258 6389 -212 6419
rect -258 6347 -252 6389
rect -218 6347 -212 6389
rect -258 6321 -212 6347
rect -258 6275 -252 6321
rect -218 6275 -212 6321
rect -258 6253 -212 6275
rect -258 6203 -252 6253
rect -218 6203 -212 6253
rect -258 6185 -212 6203
rect -258 6131 -252 6185
rect -218 6131 -212 6185
rect -258 6117 -212 6131
rect -258 6059 -252 6117
rect -218 6059 -212 6117
rect -258 6049 -212 6059
rect -258 5987 -252 6049
rect -218 5987 -212 6049
rect -258 5981 -212 5987
rect -258 5915 -252 5981
rect -218 5915 -212 5981
rect -258 5913 -212 5915
rect -258 5879 -252 5913
rect -218 5879 -212 5913
rect -258 5877 -212 5879
rect -258 5811 -252 5877
rect -218 5811 -212 5877
rect -258 5805 -212 5811
rect -258 5743 -252 5805
rect -218 5743 -212 5805
rect -258 5733 -212 5743
rect -258 5675 -252 5733
rect -218 5675 -212 5733
rect -258 5661 -212 5675
rect -258 5607 -252 5661
rect -218 5607 -212 5661
rect -258 5589 -212 5607
rect -258 5539 -252 5589
rect -218 5539 -212 5589
rect -258 5517 -212 5539
rect -258 5471 -252 5517
rect -218 5471 -212 5517
rect -258 5445 -212 5471
rect -258 5403 -252 5445
rect -218 5403 -212 5445
rect -258 5373 -212 5403
rect -258 5335 -252 5373
rect -218 5335 -212 5373
rect -258 5301 -212 5335
rect -258 5267 -252 5301
rect -218 5267 -212 5301
rect -258 5233 -212 5267
rect -258 5195 -252 5233
rect -218 5195 -212 5233
rect -258 5165 -212 5195
rect -258 5123 -252 5165
rect -218 5123 -212 5165
rect -258 5097 -212 5123
rect -258 5051 -252 5097
rect -218 5051 -212 5097
rect -258 5029 -212 5051
rect -258 4979 -252 5029
rect -218 4979 -212 5029
rect -258 4961 -212 4979
rect -258 4907 -252 4961
rect -218 4907 -212 4961
rect -258 4893 -212 4907
rect -258 4835 -252 4893
rect -218 4835 -212 4893
rect -258 4825 -212 4835
rect -258 4763 -252 4825
rect -218 4763 -212 4825
rect -258 4757 -212 4763
rect -258 4691 -252 4757
rect -218 4691 -212 4757
rect -258 4689 -212 4691
rect -258 4655 -252 4689
rect -218 4655 -212 4689
rect -258 4653 -212 4655
rect -258 4587 -252 4653
rect -218 4587 -212 4653
rect -258 4581 -212 4587
rect -258 4519 -252 4581
rect -218 4519 -212 4581
rect -258 4509 -212 4519
rect -258 4451 -252 4509
rect -218 4451 -212 4509
rect -258 4437 -212 4451
rect -258 4383 -252 4437
rect -218 4383 -212 4437
rect -258 4365 -212 4383
rect -258 4315 -252 4365
rect -218 4315 -212 4365
rect -258 4293 -212 4315
rect -258 4247 -252 4293
rect -218 4247 -212 4293
rect -258 4221 -212 4247
rect -258 4179 -252 4221
rect -218 4179 -212 4221
rect -258 4149 -212 4179
rect -258 4111 -252 4149
rect -218 4111 -212 4149
rect -258 4077 -212 4111
rect -258 4043 -252 4077
rect -218 4043 -212 4077
rect -258 4009 -212 4043
rect -258 3971 -252 4009
rect -218 3971 -212 4009
rect -258 3941 -212 3971
rect -258 3899 -252 3941
rect -218 3899 -212 3941
rect -258 3873 -212 3899
rect -258 3827 -252 3873
rect -218 3827 -212 3873
rect -258 3805 -212 3827
rect -258 3755 -252 3805
rect -218 3755 -212 3805
rect -258 3737 -212 3755
rect -258 3683 -252 3737
rect -218 3683 -212 3737
rect -258 3669 -212 3683
rect -258 3611 -252 3669
rect -218 3611 -212 3669
rect -258 3601 -212 3611
rect -258 3539 -252 3601
rect -218 3539 -212 3601
rect -258 3533 -212 3539
rect -258 3467 -252 3533
rect -218 3467 -212 3533
rect 1824 38685 1870 38717
rect 1824 38651 1830 38685
rect 1864 38651 1870 38685
rect 1824 38641 1870 38651
rect 1824 38578 1830 38641
rect 1864 38578 1870 38641
rect 1824 38573 1870 38578
rect 1824 38471 1830 38573
rect 1864 38471 1870 38573
rect 1824 38466 1870 38471
rect 1824 38403 1830 38466
rect 1864 38403 1870 38466
rect 1824 38393 1870 38403
rect 1824 38335 1830 38393
rect 1864 38335 1870 38393
rect 1824 38320 1870 38335
rect 1824 38267 1830 38320
rect 1864 38267 1870 38320
rect 1824 38247 1870 38267
rect 1824 38199 1830 38247
rect 1864 38199 1870 38247
rect 1824 38174 1870 38199
rect 1824 38131 1830 38174
rect 1864 38131 1870 38174
rect 1824 38101 1870 38131
rect 1824 38063 1830 38101
rect 1864 38063 1870 38101
rect 1824 38029 1870 38063
rect 1824 37994 1830 38029
rect 1864 37994 1870 38029
rect 1824 37961 1870 37994
rect 1824 37921 1830 37961
rect 1864 37921 1870 37961
rect 1824 37893 1870 37921
rect 1824 37848 1830 37893
rect 1864 37848 1870 37893
rect 1824 37825 1870 37848
rect 1824 37775 1830 37825
rect 1864 37775 1870 37825
rect 1824 37757 1870 37775
rect 1824 37702 1830 37757
rect 1864 37702 1870 37757
rect 1824 37689 1870 37702
rect 1824 37629 1830 37689
rect 1864 37629 1870 37689
rect 1824 37621 1870 37629
rect 1824 37556 1830 37621
rect 1864 37556 1870 37621
rect 1824 37553 1870 37556
rect 1824 37519 1830 37553
rect 1864 37519 1870 37553
rect 1824 37517 1870 37519
rect 1824 37451 1830 37517
rect 1864 37451 1870 37517
rect 1824 37444 1870 37451
rect 1824 37383 1830 37444
rect 1864 37383 1870 37444
rect 1824 37371 1870 37383
rect 1824 37315 1830 37371
rect 1864 37315 1870 37371
rect 1824 37298 1870 37315
rect 1824 37247 1830 37298
rect 1864 37247 1870 37298
rect 1824 37225 1870 37247
rect 1824 37179 1830 37225
rect 1864 37179 1870 37225
rect 1824 37152 1870 37179
rect 1824 37111 1830 37152
rect 1864 37111 1870 37152
rect 1824 37079 1870 37111
rect 1824 37043 1830 37079
rect 1864 37043 1870 37079
rect 1824 37009 1870 37043
rect 1824 36972 1830 37009
rect 1864 36972 1870 37009
rect 1824 36941 1870 36972
rect 1824 36899 1830 36941
rect 1864 36899 1870 36941
rect 1824 36873 1870 36899
rect 1824 36826 1830 36873
rect 1864 36826 1870 36873
rect 1824 36805 1870 36826
rect 1824 36753 1830 36805
rect 1864 36753 1870 36805
rect 1824 36737 1870 36753
rect 1824 36680 1830 36737
rect 1864 36680 1870 36737
rect 1824 36669 1870 36680
rect 1824 36607 1830 36669
rect 1864 36607 1870 36669
rect 1824 36601 1870 36607
rect 1824 36534 1830 36601
rect 1864 36534 1870 36601
rect 1824 36533 1870 36534
rect 1824 36499 1830 36533
rect 1864 36499 1870 36533
rect 1824 36495 1870 36499
rect 1824 36431 1830 36495
rect 1864 36431 1870 36495
rect 1824 36422 1870 36431
rect 1824 36363 1830 36422
rect 1864 36363 1870 36422
rect 1824 36349 1870 36363
rect 1824 36295 1830 36349
rect 1864 36295 1870 36349
rect 1824 36276 1870 36295
rect 1824 36227 1830 36276
rect 1864 36227 1870 36276
rect 1824 36203 1870 36227
rect 1824 36159 1830 36203
rect 1864 36159 1870 36203
rect 1824 36130 1870 36159
rect 1824 36091 1830 36130
rect 1864 36091 1870 36130
rect 1824 36057 1870 36091
rect 1824 36023 1830 36057
rect 1864 36023 1870 36057
rect 1824 35989 1870 36023
rect 1824 35950 1830 35989
rect 1864 35950 1870 35989
rect 1824 35921 1870 35950
rect 1824 35877 1830 35921
rect 1864 35877 1870 35921
rect 1824 35853 1870 35877
rect 1824 35804 1830 35853
rect 1864 35804 1870 35853
rect 1824 35785 1870 35804
rect 1824 35731 1830 35785
rect 1864 35731 1870 35785
rect 1824 35717 1870 35731
rect 1824 35658 1830 35717
rect 1864 35658 1870 35717
rect 1824 35649 1870 35658
rect 1824 35585 1830 35649
rect 1864 35585 1870 35649
rect 1824 35581 1870 35585
rect 1824 35547 1830 35581
rect 1864 35547 1870 35581
rect 1824 35546 1870 35547
rect 1824 35479 1830 35546
rect 1864 35479 1870 35546
rect 1824 35473 1870 35479
rect 1824 35411 1830 35473
rect 1864 35411 1870 35473
rect 1824 35400 1870 35411
rect 1824 35343 1830 35400
rect 1864 35343 1870 35400
rect 1824 35327 1870 35343
rect 1824 35275 1830 35327
rect 1864 35275 1870 35327
rect 1824 35254 1870 35275
rect 1824 35207 1830 35254
rect 1864 35207 1870 35254
rect 1824 35181 1870 35207
rect 1824 35139 1830 35181
rect 1864 35139 1870 35181
rect 1824 35109 1870 35139
rect 1824 35071 1830 35109
rect 1864 35071 1870 35109
rect 1824 35037 1870 35071
rect 1824 35003 1830 35037
rect 1864 35003 1870 35037
rect 1824 34969 1870 35003
rect 1824 34931 1830 34969
rect 1864 34931 1870 34969
rect 1824 34901 1870 34931
rect 1824 34859 1830 34901
rect 1864 34859 1870 34901
rect 1824 34833 1870 34859
rect 1824 34787 1830 34833
rect 1864 34787 1870 34833
rect 1824 34765 1870 34787
rect 1824 34715 1830 34765
rect 1864 34715 1870 34765
rect 1824 34697 1870 34715
rect 1824 34643 1830 34697
rect 1864 34643 1870 34697
rect 1824 34629 1870 34643
rect 1824 34571 1830 34629
rect 1864 34571 1870 34629
rect 1824 34561 1870 34571
rect 1824 34499 1830 34561
rect 1864 34499 1870 34561
rect 1824 34493 1870 34499
rect 1824 34427 1830 34493
rect 1864 34427 1870 34493
rect 1824 34425 1870 34427
rect 1824 34391 1830 34425
rect 1864 34391 1870 34425
rect 1824 34389 1870 34391
rect 1824 34323 1830 34389
rect 1864 34323 1870 34389
rect 1824 34317 1870 34323
rect 1824 34255 1830 34317
rect 1864 34255 1870 34317
rect 1824 34245 1870 34255
rect 1824 34187 1830 34245
rect 1864 34187 1870 34245
rect 1824 34173 1870 34187
rect 1824 34119 1830 34173
rect 1864 34119 1870 34173
rect 1824 34101 1870 34119
rect 1824 34051 1830 34101
rect 1864 34051 1870 34101
rect 1824 34029 1870 34051
rect 1824 33983 1830 34029
rect 1864 33983 1870 34029
rect 1824 33957 1870 33983
rect 1824 33915 1830 33957
rect 1864 33915 1870 33957
rect 1824 33885 1870 33915
rect 1824 33847 1830 33885
rect 1864 33847 1870 33885
rect 1824 33813 1870 33847
rect 1824 33779 1830 33813
rect 1864 33779 1870 33813
rect 1824 33745 1870 33779
rect 1824 33707 1830 33745
rect 1864 33707 1870 33745
rect 1824 33677 1870 33707
rect 1824 33635 1830 33677
rect 1864 33635 1870 33677
rect 1824 33609 1870 33635
rect 1824 33563 1830 33609
rect 1864 33563 1870 33609
rect 1824 33541 1870 33563
rect 1824 33491 1830 33541
rect 1864 33491 1870 33541
rect 1824 33473 1870 33491
rect 1824 33419 1830 33473
rect 1864 33419 1870 33473
rect 1824 33405 1870 33419
rect 1824 33347 1830 33405
rect 1864 33347 1870 33405
rect 1824 33337 1870 33347
rect 1824 33275 1830 33337
rect 1864 33275 1870 33337
rect 1824 33269 1870 33275
rect 1824 33203 1830 33269
rect 1864 33203 1870 33269
rect 1824 33201 1870 33203
rect 1824 33167 1830 33201
rect 1864 33167 1870 33201
rect 1824 33165 1870 33167
rect 1824 33099 1830 33165
rect 1864 33099 1870 33165
rect 1824 33093 1870 33099
rect 1824 33031 1830 33093
rect 1864 33031 1870 33093
rect 1824 33021 1870 33031
rect 1824 32963 1830 33021
rect 1864 32963 1870 33021
rect 1824 32949 1870 32963
rect 1824 32895 1830 32949
rect 1864 32895 1870 32949
rect 1824 32877 1870 32895
rect 1824 32827 1830 32877
rect 1864 32827 1870 32877
rect 1824 32805 1870 32827
rect 1824 32759 1830 32805
rect 1864 32759 1870 32805
rect 1824 32733 1870 32759
rect 1824 32691 1830 32733
rect 1864 32691 1870 32733
rect 1824 32661 1870 32691
rect 1824 32623 1830 32661
rect 1864 32623 1870 32661
rect 1824 32589 1870 32623
rect 1824 32555 1830 32589
rect 1864 32555 1870 32589
rect 1824 32521 1870 32555
rect 1824 32483 1830 32521
rect 1864 32483 1870 32521
rect 1824 32453 1870 32483
rect 1824 32411 1830 32453
rect 1864 32411 1870 32453
rect 1824 32385 1870 32411
rect 1824 32339 1830 32385
rect 1864 32339 1870 32385
rect 1824 32317 1870 32339
rect 1824 32267 1830 32317
rect 1864 32267 1870 32317
rect 1824 32249 1870 32267
rect 1824 32195 1830 32249
rect 1864 32195 1870 32249
rect 1824 32181 1870 32195
rect 1824 32123 1830 32181
rect 1864 32123 1870 32181
rect 1824 32113 1870 32123
rect 1824 32051 1830 32113
rect 1864 32051 1870 32113
rect 1824 32045 1870 32051
rect 1824 31979 1830 32045
rect 1864 31979 1870 32045
rect 1824 31977 1870 31979
rect 1824 31943 1830 31977
rect 1864 31943 1870 31977
rect 1824 31941 1870 31943
rect 1824 31875 1830 31941
rect 1864 31875 1870 31941
rect 1824 31869 1870 31875
rect 1824 31807 1830 31869
rect 1864 31807 1870 31869
rect 1824 31797 1870 31807
rect 1824 31739 1830 31797
rect 1864 31739 1870 31797
rect 1824 31725 1870 31739
rect 1824 31671 1830 31725
rect 1864 31671 1870 31725
rect 1824 31653 1870 31671
rect 1824 31603 1830 31653
rect 1864 31603 1870 31653
rect 1824 31581 1870 31603
rect 1824 31535 1830 31581
rect 1864 31535 1870 31581
rect 1824 31509 1870 31535
rect 1824 31467 1830 31509
rect 1864 31467 1870 31509
rect 1824 31437 1870 31467
rect 1824 31399 1830 31437
rect 1864 31399 1870 31437
rect 1824 31365 1870 31399
rect 1824 31331 1830 31365
rect 1864 31331 1870 31365
rect 1824 31297 1870 31331
rect 1824 31259 1830 31297
rect 1864 31259 1870 31297
rect 1824 31229 1870 31259
rect 1824 31187 1830 31229
rect 1864 31187 1870 31229
rect 1824 31161 1870 31187
rect 1824 31115 1830 31161
rect 1864 31115 1870 31161
rect 1824 31093 1870 31115
rect 1824 31043 1830 31093
rect 1864 31043 1870 31093
rect 1824 31025 1870 31043
rect 1824 30971 1830 31025
rect 1864 30971 1870 31025
rect 1824 30957 1870 30971
rect 1824 30899 1830 30957
rect 1864 30899 1870 30957
rect 1824 30889 1870 30899
rect 1824 30827 1830 30889
rect 1864 30827 1870 30889
rect 1824 30821 1870 30827
rect 1824 30755 1830 30821
rect 1864 30755 1870 30821
rect 1824 30753 1870 30755
rect 1824 30719 1830 30753
rect 1864 30719 1870 30753
rect 1824 30717 1870 30719
rect 1824 30651 1830 30717
rect 1864 30651 1870 30717
rect 1824 30645 1870 30651
rect 1824 30583 1830 30645
rect 1864 30583 1870 30645
rect 1824 30573 1870 30583
rect 1824 30515 1830 30573
rect 1864 30515 1870 30573
rect 1824 30501 1870 30515
rect 1824 30447 1830 30501
rect 1864 30447 1870 30501
rect 1824 30429 1870 30447
rect 1824 30379 1830 30429
rect 1864 30379 1870 30429
rect 1824 30357 1870 30379
rect 1824 30311 1830 30357
rect 1864 30311 1870 30357
rect 1824 30285 1870 30311
rect 1824 30243 1830 30285
rect 1864 30243 1870 30285
rect 1824 30213 1870 30243
rect 1824 30175 1830 30213
rect 1864 30175 1870 30213
rect 1824 30141 1870 30175
rect 1824 30107 1830 30141
rect 1864 30107 1870 30141
rect 1824 30073 1870 30107
rect 1824 30035 1830 30073
rect 1864 30035 1870 30073
rect 1824 30005 1870 30035
rect 1824 29963 1830 30005
rect 1864 29963 1870 30005
rect 1824 29937 1870 29963
rect 1824 29891 1830 29937
rect 1864 29891 1870 29937
rect 1824 29869 1870 29891
rect 1824 29819 1830 29869
rect 1864 29819 1870 29869
rect 1824 29801 1870 29819
rect 1824 29747 1830 29801
rect 1864 29747 1870 29801
rect 1824 29733 1870 29747
rect 1824 29675 1830 29733
rect 1864 29675 1870 29733
rect 1824 29665 1870 29675
rect 1824 29603 1830 29665
rect 1864 29603 1870 29665
rect 1824 29597 1870 29603
rect 1824 29531 1830 29597
rect 1864 29531 1870 29597
rect 1824 29529 1870 29531
rect 1824 29495 1830 29529
rect 1864 29495 1870 29529
rect 1824 29493 1870 29495
rect 1824 29427 1830 29493
rect 1864 29427 1870 29493
rect 1824 29421 1870 29427
rect 1824 29359 1830 29421
rect 1864 29359 1870 29421
rect 1824 29349 1870 29359
rect 1824 29291 1830 29349
rect 1864 29291 1870 29349
rect 1824 29277 1870 29291
rect 1824 29223 1830 29277
rect 1864 29223 1870 29277
rect 1824 29205 1870 29223
rect 1824 29155 1830 29205
rect 1864 29155 1870 29205
rect 1824 29133 1870 29155
rect 1824 29087 1830 29133
rect 1864 29087 1870 29133
rect 1824 29061 1870 29087
rect 1824 29019 1830 29061
rect 1864 29019 1870 29061
rect 1824 28989 1870 29019
rect 1824 28951 1830 28989
rect 1864 28951 1870 28989
rect 1824 28917 1870 28951
rect 1824 28883 1830 28917
rect 1864 28883 1870 28917
rect 1824 28849 1870 28883
rect 1824 28811 1830 28849
rect 1864 28811 1870 28849
rect 1824 28781 1870 28811
rect 1824 28739 1830 28781
rect 1864 28739 1870 28781
rect 1824 28713 1870 28739
rect 1824 28667 1830 28713
rect 1864 28667 1870 28713
rect 1824 28645 1870 28667
rect 1824 28595 1830 28645
rect 1864 28595 1870 28645
rect 1824 28577 1870 28595
rect 1824 28523 1830 28577
rect 1864 28523 1870 28577
rect 1824 28509 1870 28523
rect 1824 28451 1830 28509
rect 1864 28451 1870 28509
rect 1824 28441 1870 28451
rect 1824 28379 1830 28441
rect 1864 28379 1870 28441
rect 1824 28373 1870 28379
rect 1824 28307 1830 28373
rect 1864 28307 1870 28373
rect 1824 28305 1870 28307
rect 1824 28271 1830 28305
rect 1864 28271 1870 28305
rect 1824 28269 1870 28271
rect 1824 28203 1830 28269
rect 1864 28203 1870 28269
rect 1824 28197 1870 28203
rect 1824 28135 1830 28197
rect 1864 28135 1870 28197
rect 1824 28125 1870 28135
rect 1824 28067 1830 28125
rect 1864 28067 1870 28125
rect 1824 28053 1870 28067
rect 1824 27999 1830 28053
rect 1864 27999 1870 28053
rect 1824 27981 1870 27999
rect 1824 27931 1830 27981
rect 1864 27931 1870 27981
rect 1824 27909 1870 27931
rect 1824 27863 1830 27909
rect 1864 27863 1870 27909
rect 1824 27837 1870 27863
rect 1824 27795 1830 27837
rect 1864 27795 1870 27837
rect 1824 27765 1870 27795
rect 1824 27727 1830 27765
rect 1864 27727 1870 27765
rect 1824 27693 1870 27727
rect 1824 27659 1830 27693
rect 1864 27659 1870 27693
rect 1824 27625 1870 27659
rect 1824 27587 1830 27625
rect 1864 27587 1870 27625
rect 1824 27557 1870 27587
rect 1824 27515 1830 27557
rect 1864 27515 1870 27557
rect 1824 27489 1870 27515
rect 1824 27443 1830 27489
rect 1864 27443 1870 27489
rect 1824 27421 1870 27443
rect 1824 27371 1830 27421
rect 1864 27371 1870 27421
rect 1824 27353 1870 27371
rect 1824 27299 1830 27353
rect 1864 27299 1870 27353
rect 1824 27285 1870 27299
rect 1824 27227 1830 27285
rect 1864 27227 1870 27285
rect 1824 27217 1870 27227
rect 1824 27155 1830 27217
rect 1864 27155 1870 27217
rect 1824 27149 1870 27155
rect 1824 27083 1830 27149
rect 1864 27083 1870 27149
rect 1824 27081 1870 27083
rect 1824 27047 1830 27081
rect 1864 27047 1870 27081
rect 1824 27045 1870 27047
rect 1824 26979 1830 27045
rect 1864 26979 1870 27045
rect 1824 26973 1870 26979
rect 1824 26911 1830 26973
rect 1864 26911 1870 26973
rect 1824 26901 1870 26911
rect 1824 26843 1830 26901
rect 1864 26843 1870 26901
rect 1824 26829 1870 26843
rect 1824 26775 1830 26829
rect 1864 26775 1870 26829
rect 1824 26757 1870 26775
rect 1824 26707 1830 26757
rect 1864 26707 1870 26757
rect 1824 26685 1870 26707
rect 1824 26639 1830 26685
rect 1864 26639 1870 26685
rect 1824 26613 1870 26639
rect 1824 26571 1830 26613
rect 1864 26571 1870 26613
rect 1824 26541 1870 26571
rect 1824 26503 1830 26541
rect 1864 26503 1870 26541
rect 1824 26469 1870 26503
rect 1824 26435 1830 26469
rect 1864 26435 1870 26469
rect 1824 26401 1870 26435
rect 1824 26363 1830 26401
rect 1864 26363 1870 26401
rect 1824 26333 1870 26363
rect 1824 26291 1830 26333
rect 1864 26291 1870 26333
rect 1824 26265 1870 26291
rect 1824 26219 1830 26265
rect 1864 26219 1870 26265
rect 1824 26197 1870 26219
rect 1824 26147 1830 26197
rect 1864 26147 1870 26197
rect 1824 26129 1870 26147
rect 1824 26075 1830 26129
rect 1864 26075 1870 26129
rect 1824 26061 1870 26075
rect 1824 26003 1830 26061
rect 1864 26003 1870 26061
rect 1824 25993 1870 26003
rect 1824 25931 1830 25993
rect 1864 25931 1870 25993
rect 1824 25925 1870 25931
rect 1824 25859 1830 25925
rect 1864 25859 1870 25925
rect 1824 25857 1870 25859
rect 1824 25823 1830 25857
rect 1864 25823 1870 25857
rect 1824 25821 1870 25823
rect 1824 25755 1830 25821
rect 1864 25755 1870 25821
rect 1824 25749 1870 25755
rect 1824 25687 1830 25749
rect 1864 25687 1870 25749
rect 1824 25677 1870 25687
rect 1824 25619 1830 25677
rect 1864 25619 1870 25677
rect 1824 25605 1870 25619
rect 1824 25551 1830 25605
rect 1864 25551 1870 25605
rect 1824 25533 1870 25551
rect 1824 25483 1830 25533
rect 1864 25483 1870 25533
rect 1824 25461 1870 25483
rect 1824 25415 1830 25461
rect 1864 25415 1870 25461
rect 1824 25389 1870 25415
rect 1824 25347 1830 25389
rect 1864 25347 1870 25389
rect 1824 25317 1870 25347
rect 1824 25279 1830 25317
rect 1864 25279 1870 25317
rect 1824 25245 1870 25279
rect 1824 25211 1830 25245
rect 1864 25211 1870 25245
rect 1824 25177 1870 25211
rect 1824 25139 1830 25177
rect 1864 25139 1870 25177
rect 1824 25109 1870 25139
rect 1824 25067 1830 25109
rect 1864 25067 1870 25109
rect 1824 25041 1870 25067
rect 1824 24995 1830 25041
rect 1864 24995 1870 25041
rect 1824 24973 1870 24995
rect 1824 24923 1830 24973
rect 1864 24923 1870 24973
rect 1824 24905 1870 24923
rect 1824 24851 1830 24905
rect 1864 24851 1870 24905
rect 1824 24837 1870 24851
rect 1824 24779 1830 24837
rect 1864 24779 1870 24837
rect 1824 24769 1870 24779
rect 1824 24707 1830 24769
rect 1864 24707 1870 24769
rect 1824 24701 1870 24707
rect 1824 24635 1830 24701
rect 1864 24635 1870 24701
rect 1824 24633 1870 24635
rect 1824 24599 1830 24633
rect 1864 24599 1870 24633
rect 1824 24597 1870 24599
rect 1824 24531 1830 24597
rect 1864 24531 1870 24597
rect 1824 24525 1870 24531
rect 1824 24463 1830 24525
rect 1864 24463 1870 24525
rect 1824 24453 1870 24463
rect 1824 24395 1830 24453
rect 1864 24395 1870 24453
rect 1824 24381 1870 24395
rect 1824 24327 1830 24381
rect 1864 24327 1870 24381
rect 1824 24309 1870 24327
rect 1824 24259 1830 24309
rect 1864 24259 1870 24309
rect 1824 24237 1870 24259
rect 1824 24191 1830 24237
rect 1864 24191 1870 24237
rect 1824 24165 1870 24191
rect 1824 24123 1830 24165
rect 1864 24123 1870 24165
rect 1824 24093 1870 24123
rect 1824 24055 1830 24093
rect 1864 24055 1870 24093
rect 1824 24021 1870 24055
rect 1824 23987 1830 24021
rect 1864 23987 1870 24021
rect 1824 23953 1870 23987
rect 1824 23915 1830 23953
rect 1864 23915 1870 23953
rect 1824 23885 1870 23915
rect 1824 23843 1830 23885
rect 1864 23843 1870 23885
rect 1824 23817 1870 23843
rect 1824 23771 1830 23817
rect 1864 23771 1870 23817
rect 1824 23749 1870 23771
rect 1824 23699 1830 23749
rect 1864 23699 1870 23749
rect 1824 23681 1870 23699
rect 1824 23627 1830 23681
rect 1864 23627 1870 23681
rect 1824 23613 1870 23627
rect 1824 23555 1830 23613
rect 1864 23555 1870 23613
rect 1824 23545 1870 23555
rect 1824 23483 1830 23545
rect 1864 23483 1870 23545
rect 1824 23477 1870 23483
rect 1824 23411 1830 23477
rect 1864 23411 1870 23477
rect 1824 23409 1870 23411
rect 1824 23375 1830 23409
rect 1864 23375 1870 23409
rect 1824 23373 1870 23375
rect 1824 23307 1830 23373
rect 1864 23307 1870 23373
rect 1824 23301 1870 23307
rect 1824 23239 1830 23301
rect 1864 23239 1870 23301
rect 1824 23229 1870 23239
rect 1824 23171 1830 23229
rect 1864 23171 1870 23229
rect 1824 23157 1870 23171
rect 1824 23103 1830 23157
rect 1864 23103 1870 23157
rect 1824 23085 1870 23103
rect 1824 23035 1830 23085
rect 1864 23035 1870 23085
rect 1824 23013 1870 23035
rect 1824 22967 1830 23013
rect 1864 22967 1870 23013
rect 1824 22941 1870 22967
rect 1824 22899 1830 22941
rect 1864 22899 1870 22941
rect 1824 22869 1870 22899
rect 1824 22831 1830 22869
rect 1864 22831 1870 22869
rect 1824 22797 1870 22831
rect 1824 22763 1830 22797
rect 1864 22763 1870 22797
rect 1824 22729 1870 22763
rect 1824 22691 1830 22729
rect 1864 22691 1870 22729
rect 1824 22661 1870 22691
rect 1824 22619 1830 22661
rect 1864 22619 1870 22661
rect 1824 22593 1870 22619
rect 1824 22547 1830 22593
rect 1864 22547 1870 22593
rect 1824 22525 1870 22547
rect 1824 22475 1830 22525
rect 1864 22475 1870 22525
rect 1824 22457 1870 22475
rect 1824 22403 1830 22457
rect 1864 22403 1870 22457
rect 1824 22389 1870 22403
rect 1824 22331 1830 22389
rect 1864 22331 1870 22389
rect 1824 22321 1870 22331
rect 1824 22259 1830 22321
rect 1864 22259 1870 22321
rect 1824 22253 1870 22259
rect 1824 22187 1830 22253
rect 1864 22187 1870 22253
rect 1824 22185 1870 22187
rect 1824 22151 1830 22185
rect 1864 22151 1870 22185
rect 1824 22149 1870 22151
rect 1824 22083 1830 22149
rect 1864 22083 1870 22149
rect 1824 22077 1870 22083
rect 1824 22015 1830 22077
rect 1864 22015 1870 22077
rect 1824 22005 1870 22015
rect 1824 21947 1830 22005
rect 1864 21947 1870 22005
rect 1824 21933 1870 21947
rect 1824 21879 1830 21933
rect 1864 21879 1870 21933
rect 1824 21861 1870 21879
rect 1824 21811 1830 21861
rect 1864 21811 1870 21861
rect 1824 21789 1870 21811
rect 1824 21743 1830 21789
rect 1864 21743 1870 21789
rect 1824 21717 1870 21743
rect 1824 21675 1830 21717
rect 1864 21675 1870 21717
rect 1824 21645 1870 21675
rect 1824 21607 1830 21645
rect 1864 21607 1870 21645
rect 1824 21573 1870 21607
rect 1824 21539 1830 21573
rect 1864 21539 1870 21573
rect 1824 21505 1870 21539
rect 1824 21467 1830 21505
rect 1864 21467 1870 21505
rect 1824 21437 1870 21467
rect 1824 21395 1830 21437
rect 1864 21395 1870 21437
rect 1824 21369 1870 21395
rect 1824 21323 1830 21369
rect 1864 21323 1870 21369
rect 1824 21301 1870 21323
rect 1824 21251 1830 21301
rect 1864 21251 1870 21301
rect 1824 21233 1870 21251
rect 1824 21179 1830 21233
rect 1864 21179 1870 21233
rect 1824 21165 1870 21179
rect 1824 21107 1830 21165
rect 1864 21107 1870 21165
rect 1824 21097 1870 21107
rect 1824 21035 1830 21097
rect 1864 21035 1870 21097
rect 1824 21029 1870 21035
rect 1824 20963 1830 21029
rect 1864 20963 1870 21029
rect 1824 20961 1870 20963
rect 1824 20927 1830 20961
rect 1864 20927 1870 20961
rect 1824 20925 1870 20927
rect 1824 20859 1830 20925
rect 1864 20859 1870 20925
rect 1824 20853 1870 20859
rect 1824 20791 1830 20853
rect 1864 20791 1870 20853
rect 1824 20781 1870 20791
rect 1824 20723 1830 20781
rect 1864 20723 1870 20781
rect 1824 20709 1870 20723
rect 1824 20655 1830 20709
rect 1864 20655 1870 20709
rect 1824 20637 1870 20655
rect 1824 20587 1830 20637
rect 1864 20587 1870 20637
rect 1824 20565 1870 20587
rect 1824 20519 1830 20565
rect 1864 20519 1870 20565
rect 1824 20493 1870 20519
rect 1824 20451 1830 20493
rect 1864 20451 1870 20493
rect 1824 20421 1870 20451
rect 1824 20383 1830 20421
rect 1864 20383 1870 20421
rect 1824 20349 1870 20383
rect 1824 20315 1830 20349
rect 1864 20315 1870 20349
rect 1824 20281 1870 20315
rect 1824 20243 1830 20281
rect 1864 20243 1870 20281
rect 1824 20213 1870 20243
rect 1824 20171 1830 20213
rect 1864 20171 1870 20213
rect 1824 20145 1870 20171
rect 1824 20099 1830 20145
rect 1864 20099 1870 20145
rect 1824 20077 1870 20099
rect 1824 20027 1830 20077
rect 1864 20027 1870 20077
rect 1824 20009 1870 20027
rect 1824 19955 1830 20009
rect 1864 19955 1870 20009
rect 1824 19941 1870 19955
rect 1824 19883 1830 19941
rect 1864 19883 1870 19941
rect 1824 19873 1870 19883
rect 1824 19811 1830 19873
rect 1864 19811 1870 19873
rect 1824 19805 1870 19811
rect 1824 19739 1830 19805
rect 1864 19739 1870 19805
rect 1824 19737 1870 19739
rect 1824 19703 1830 19737
rect 1864 19703 1870 19737
rect 1824 19701 1870 19703
rect 1824 19635 1830 19701
rect 1864 19635 1870 19701
rect 1824 19629 1870 19635
rect 1824 19567 1830 19629
rect 1864 19567 1870 19629
rect 1824 19557 1870 19567
rect 1824 19499 1830 19557
rect 1864 19499 1870 19557
rect 1824 19485 1870 19499
rect 1824 19431 1830 19485
rect 1864 19431 1870 19485
rect 1824 19413 1870 19431
rect 1824 19363 1830 19413
rect 1864 19363 1870 19413
rect 1824 19341 1870 19363
rect 1824 19295 1830 19341
rect 1864 19295 1870 19341
rect 1824 19269 1870 19295
rect 1824 19227 1830 19269
rect 1864 19227 1870 19269
rect 1824 19197 1870 19227
rect 1824 19159 1830 19197
rect 1864 19159 1870 19197
rect 1824 19125 1870 19159
rect 1824 19091 1830 19125
rect 1864 19091 1870 19125
rect 1824 19057 1870 19091
rect 1824 19019 1830 19057
rect 1864 19019 1870 19057
rect 1824 18989 1870 19019
rect 1824 18947 1830 18989
rect 1864 18947 1870 18989
rect 1824 18921 1870 18947
rect 1824 18875 1830 18921
rect 1864 18875 1870 18921
rect 1824 18853 1870 18875
rect 1824 18803 1830 18853
rect 1864 18803 1870 18853
rect 1824 18785 1870 18803
rect 1824 18731 1830 18785
rect 1864 18731 1870 18785
rect 1824 18717 1870 18731
rect 1824 18659 1830 18717
rect 1864 18659 1870 18717
rect 1824 18649 1870 18659
rect 1824 18587 1830 18649
rect 1864 18587 1870 18649
rect 1824 18581 1870 18587
rect 1824 18515 1830 18581
rect 1864 18515 1870 18581
rect 1824 18513 1870 18515
rect 1824 18479 1830 18513
rect 1864 18479 1870 18513
rect 1824 18477 1870 18479
rect 1824 18411 1830 18477
rect 1864 18411 1870 18477
rect 1824 18405 1870 18411
rect 1824 18343 1830 18405
rect 1864 18343 1870 18405
rect 1824 18333 1870 18343
rect 1824 18275 1830 18333
rect 1864 18275 1870 18333
rect 1824 18261 1870 18275
rect 1824 18207 1830 18261
rect 1864 18207 1870 18261
rect 1824 18189 1870 18207
rect 1824 18139 1830 18189
rect 1864 18139 1870 18189
rect 1824 18117 1870 18139
rect 1824 18071 1830 18117
rect 1864 18071 1870 18117
rect 1824 18045 1870 18071
rect 1824 18003 1830 18045
rect 1864 18003 1870 18045
rect 1824 17973 1870 18003
rect 1824 17935 1830 17973
rect 1864 17935 1870 17973
rect 1824 17901 1870 17935
rect 1824 17867 1830 17901
rect 1864 17867 1870 17901
rect 1824 17833 1870 17867
rect 1824 17795 1830 17833
rect 1864 17795 1870 17833
rect 1824 17765 1870 17795
rect 1824 17723 1830 17765
rect 1864 17723 1870 17765
rect 1824 17697 1870 17723
rect 1824 17651 1830 17697
rect 1864 17651 1870 17697
rect 1824 17629 1870 17651
rect 1824 17579 1830 17629
rect 1864 17579 1870 17629
rect 1824 17561 1870 17579
rect 1824 17507 1830 17561
rect 1864 17507 1870 17561
rect 1824 17493 1870 17507
rect 1824 17435 1830 17493
rect 1864 17435 1870 17493
rect 1824 17425 1870 17435
rect 1824 17363 1830 17425
rect 1864 17363 1870 17425
rect 1824 17357 1870 17363
rect 1824 17291 1830 17357
rect 1864 17291 1870 17357
rect 1824 17289 1870 17291
rect 1824 17255 1830 17289
rect 1864 17255 1870 17289
rect 1824 17253 1870 17255
rect 1824 17187 1830 17253
rect 1864 17187 1870 17253
rect 1824 17181 1870 17187
rect 1824 17119 1830 17181
rect 1864 17119 1870 17181
rect 1824 17109 1870 17119
rect 1824 17051 1830 17109
rect 1864 17051 1870 17109
rect 1824 17037 1870 17051
rect 1824 16983 1830 17037
rect 1864 16983 1870 17037
rect 1824 16965 1870 16983
rect 1824 16915 1830 16965
rect 1864 16915 1870 16965
rect 1824 16893 1870 16915
rect 1824 16847 1830 16893
rect 1864 16847 1870 16893
rect 1824 16821 1870 16847
rect 1824 16779 1830 16821
rect 1864 16779 1870 16821
rect 1824 16749 1870 16779
rect 1824 16711 1830 16749
rect 1864 16711 1870 16749
rect 1824 16677 1870 16711
rect 1824 16643 1830 16677
rect 1864 16643 1870 16677
rect 1824 16609 1870 16643
rect 1824 16571 1830 16609
rect 1864 16571 1870 16609
rect 1824 16541 1870 16571
rect 1824 16499 1830 16541
rect 1864 16499 1870 16541
rect 1824 16473 1870 16499
rect 1824 16427 1830 16473
rect 1864 16427 1870 16473
rect 1824 16405 1870 16427
rect 1824 16355 1830 16405
rect 1864 16355 1870 16405
rect 1824 16337 1870 16355
rect 1824 16283 1830 16337
rect 1864 16283 1870 16337
rect 1824 16269 1870 16283
rect 1824 16211 1830 16269
rect 1864 16211 1870 16269
rect 1824 16201 1870 16211
rect 1824 16139 1830 16201
rect 1864 16139 1870 16201
rect 1824 16133 1870 16139
rect 1824 16067 1830 16133
rect 1864 16067 1870 16133
rect 1824 16065 1870 16067
rect 1824 16031 1830 16065
rect 1864 16031 1870 16065
rect 1824 16029 1870 16031
rect 1824 15963 1830 16029
rect 1864 15963 1870 16029
rect 1824 15957 1870 15963
rect 1824 15895 1830 15957
rect 1864 15895 1870 15957
rect 1824 15885 1870 15895
rect 1824 15827 1830 15885
rect 1864 15827 1870 15885
rect 1824 15813 1870 15827
rect 1824 15759 1830 15813
rect 1864 15759 1870 15813
rect 1824 15741 1870 15759
rect 1824 15691 1830 15741
rect 1864 15691 1870 15741
rect 1824 15669 1870 15691
rect 1824 15623 1830 15669
rect 1864 15623 1870 15669
rect 1824 15597 1870 15623
rect 1824 15555 1830 15597
rect 1864 15555 1870 15597
rect 1824 15525 1870 15555
rect 1824 15487 1830 15525
rect 1864 15487 1870 15525
rect 1824 15453 1870 15487
rect 1824 15419 1830 15453
rect 1864 15419 1870 15453
rect 1824 15385 1870 15419
rect 1824 15347 1830 15385
rect 1864 15347 1870 15385
rect 1824 15317 1870 15347
rect 1824 15275 1830 15317
rect 1864 15275 1870 15317
rect 1824 15249 1870 15275
rect 1824 15203 1830 15249
rect 1864 15203 1870 15249
rect 1824 15181 1870 15203
rect 1824 15131 1830 15181
rect 1864 15131 1870 15181
rect 1824 15113 1870 15131
rect 1824 15059 1830 15113
rect 1864 15059 1870 15113
rect 1824 15045 1870 15059
rect 1824 14987 1830 15045
rect 1864 14987 1870 15045
rect 1824 14977 1870 14987
rect 1824 14915 1830 14977
rect 1864 14915 1870 14977
rect 1824 14909 1870 14915
rect 1824 14843 1830 14909
rect 1864 14843 1870 14909
rect 1824 14841 1870 14843
rect 1824 14807 1830 14841
rect 1864 14807 1870 14841
rect 1824 14805 1870 14807
rect 1824 14739 1830 14805
rect 1864 14739 1870 14805
rect 1824 14733 1870 14739
rect 1824 14671 1830 14733
rect 1864 14671 1870 14733
rect 1824 14661 1870 14671
rect 1824 14603 1830 14661
rect 1864 14603 1870 14661
rect 1824 14589 1870 14603
rect 1824 14535 1830 14589
rect 1864 14535 1870 14589
rect 1824 14517 1870 14535
rect 1824 14467 1830 14517
rect 1864 14467 1870 14517
rect 1824 14445 1870 14467
rect 1824 14399 1830 14445
rect 1864 14399 1870 14445
rect 1824 14373 1870 14399
rect 1824 14331 1830 14373
rect 1864 14331 1870 14373
rect 1824 14301 1870 14331
rect 1824 14263 1830 14301
rect 1864 14263 1870 14301
rect 1824 14229 1870 14263
rect 1824 14195 1830 14229
rect 1864 14195 1870 14229
rect 1824 14161 1870 14195
rect 1824 14123 1830 14161
rect 1864 14123 1870 14161
rect 1824 14093 1870 14123
rect 1824 14051 1830 14093
rect 1864 14051 1870 14093
rect 1824 14025 1870 14051
rect 1824 13979 1830 14025
rect 1864 13979 1870 14025
rect 1824 13957 1870 13979
rect 1824 13907 1830 13957
rect 1864 13907 1870 13957
rect 1824 13889 1870 13907
rect 1824 13835 1830 13889
rect 1864 13835 1870 13889
rect 1824 13821 1870 13835
rect 1824 13763 1830 13821
rect 1864 13763 1870 13821
rect 1824 13753 1870 13763
rect 1824 13691 1830 13753
rect 1864 13691 1870 13753
rect 1824 13685 1870 13691
rect 1824 13619 1830 13685
rect 1864 13619 1870 13685
rect 1824 13617 1870 13619
rect 1824 13583 1830 13617
rect 1864 13583 1870 13617
rect 1824 13581 1870 13583
rect 1824 13515 1830 13581
rect 1864 13515 1870 13581
rect 1824 13509 1870 13515
rect 1824 13447 1830 13509
rect 1864 13447 1870 13509
rect 1824 13437 1870 13447
rect 1824 13379 1830 13437
rect 1864 13379 1870 13437
rect 1824 13365 1870 13379
rect 1824 13311 1830 13365
rect 1864 13311 1870 13365
rect 1824 13293 1870 13311
rect 1824 13243 1830 13293
rect 1864 13243 1870 13293
rect 1824 13221 1870 13243
rect 1824 13175 1830 13221
rect 1864 13175 1870 13221
rect 1824 13149 1870 13175
rect 1824 13107 1830 13149
rect 1864 13107 1870 13149
rect 1824 13077 1870 13107
rect 1824 13039 1830 13077
rect 1864 13039 1870 13077
rect 1824 13005 1870 13039
rect 1824 12971 1830 13005
rect 1864 12971 1870 13005
rect 1824 12937 1870 12971
rect 1824 12899 1830 12937
rect 1864 12899 1870 12937
rect 1824 12869 1870 12899
rect 1824 12827 1830 12869
rect 1864 12827 1870 12869
rect 1824 12801 1870 12827
rect 1824 12755 1830 12801
rect 1864 12755 1870 12801
rect 1824 12733 1870 12755
rect 1824 12683 1830 12733
rect 1864 12683 1870 12733
rect 1824 12665 1870 12683
rect 1824 12611 1830 12665
rect 1864 12611 1870 12665
rect 1824 12597 1870 12611
rect 1824 12539 1830 12597
rect 1864 12539 1870 12597
rect 1824 12529 1870 12539
rect 1824 12467 1830 12529
rect 1864 12467 1870 12529
rect 1824 12461 1870 12467
rect 1824 12395 1830 12461
rect 1864 12395 1870 12461
rect 1824 12393 1870 12395
rect 1824 12359 1830 12393
rect 1864 12359 1870 12393
rect 1824 12357 1870 12359
rect 1824 12291 1830 12357
rect 1864 12291 1870 12357
rect 1824 12285 1870 12291
rect 1824 12223 1830 12285
rect 1864 12223 1870 12285
rect 1824 12213 1870 12223
rect 1824 12155 1830 12213
rect 1864 12155 1870 12213
rect 1824 12141 1870 12155
rect 1824 12087 1830 12141
rect 1864 12087 1870 12141
rect 1824 12069 1870 12087
rect 1824 12019 1830 12069
rect 1864 12019 1870 12069
rect 1824 11997 1870 12019
rect 1824 11951 1830 11997
rect 1864 11951 1870 11997
rect 1824 11925 1870 11951
rect 1824 11883 1830 11925
rect 1864 11883 1870 11925
rect 1824 11853 1870 11883
rect 1824 11815 1830 11853
rect 1864 11815 1870 11853
rect 1824 11781 1870 11815
rect 1824 11747 1830 11781
rect 1864 11747 1870 11781
rect 1824 11713 1870 11747
rect 1824 11675 1830 11713
rect 1864 11675 1870 11713
rect 1824 11645 1870 11675
rect 1824 11603 1830 11645
rect 1864 11603 1870 11645
rect 1824 11577 1870 11603
rect 1824 11531 1830 11577
rect 1864 11531 1870 11577
rect 1824 11509 1870 11531
rect 1824 11459 1830 11509
rect 1864 11459 1870 11509
rect 1824 11441 1870 11459
rect 1824 11387 1830 11441
rect 1864 11387 1870 11441
rect 1824 11373 1870 11387
rect 1824 11315 1830 11373
rect 1864 11315 1870 11373
rect 1824 11305 1870 11315
rect 1824 11243 1830 11305
rect 1864 11243 1870 11305
rect 1824 11237 1870 11243
rect 1824 11171 1830 11237
rect 1864 11171 1870 11237
rect 1824 11169 1870 11171
rect 1824 11135 1830 11169
rect 1864 11135 1870 11169
rect 1824 11133 1870 11135
rect 1824 11067 1830 11133
rect 1864 11067 1870 11133
rect 1824 11061 1870 11067
rect 1824 10999 1830 11061
rect 1864 10999 1870 11061
rect 1824 10989 1870 10999
rect 1824 10931 1830 10989
rect 1864 10931 1870 10989
rect 1824 10917 1870 10931
rect 1824 10863 1830 10917
rect 1864 10863 1870 10917
rect 1824 10845 1870 10863
rect 1824 10795 1830 10845
rect 1864 10795 1870 10845
rect 1824 10773 1870 10795
rect 1824 10727 1830 10773
rect 1864 10727 1870 10773
rect 1824 10701 1870 10727
rect 1824 10659 1830 10701
rect 1864 10659 1870 10701
rect 1824 10629 1870 10659
rect 1824 10591 1830 10629
rect 1864 10591 1870 10629
rect 1824 10557 1870 10591
rect 1824 10523 1830 10557
rect 1864 10523 1870 10557
rect 1824 10489 1870 10523
rect 1824 10451 1830 10489
rect 1864 10451 1870 10489
rect 1824 10421 1870 10451
rect 1824 10379 1830 10421
rect 1864 10379 1870 10421
rect 1824 10353 1870 10379
rect 1824 10307 1830 10353
rect 1864 10307 1870 10353
rect 1824 10285 1870 10307
rect 1824 10235 1830 10285
rect 1864 10235 1870 10285
rect 1824 10217 1870 10235
rect 1824 10163 1830 10217
rect 1864 10163 1870 10217
rect 1824 10149 1870 10163
rect 1824 10091 1830 10149
rect 1864 10091 1870 10149
rect 1824 10081 1870 10091
rect 1824 10019 1830 10081
rect 1864 10019 1870 10081
rect 1824 10013 1870 10019
rect 1824 9947 1830 10013
rect 1864 9947 1870 10013
rect 1824 9945 1870 9947
rect 1824 9911 1830 9945
rect 1864 9911 1870 9945
rect 1824 9909 1870 9911
rect 1824 9843 1830 9909
rect 1864 9843 1870 9909
rect 1824 9837 1870 9843
rect 1824 9775 1830 9837
rect 1864 9775 1870 9837
rect 1824 9765 1870 9775
rect 1824 9707 1830 9765
rect 1864 9707 1870 9765
rect 1824 9693 1870 9707
rect 1824 9639 1830 9693
rect 1864 9639 1870 9693
rect 1824 9621 1870 9639
rect 1824 9571 1830 9621
rect 1864 9571 1870 9621
rect 1824 9549 1870 9571
rect 1824 9503 1830 9549
rect 1864 9503 1870 9549
rect 1824 9477 1870 9503
rect 1824 9435 1830 9477
rect 1864 9435 1870 9477
rect 1824 9405 1870 9435
rect 1824 9367 1830 9405
rect 1864 9367 1870 9405
rect 1824 9333 1870 9367
rect 1824 9299 1830 9333
rect 1864 9299 1870 9333
rect 1824 9265 1870 9299
rect 1824 9227 1830 9265
rect 1864 9227 1870 9265
rect 1824 9197 1870 9227
rect 1824 9155 1830 9197
rect 1864 9155 1870 9197
rect 1824 9129 1870 9155
rect 1824 9083 1830 9129
rect 1864 9083 1870 9129
rect 1824 9061 1870 9083
rect 1824 9011 1830 9061
rect 1864 9011 1870 9061
rect 1824 8993 1870 9011
rect 1824 8939 1830 8993
rect 1864 8939 1870 8993
rect 1824 8925 1870 8939
rect 1824 8867 1830 8925
rect 1864 8867 1870 8925
rect 1824 8857 1870 8867
rect 1824 8795 1830 8857
rect 1864 8795 1870 8857
rect 1824 8789 1870 8795
rect 1824 8723 1830 8789
rect 1864 8723 1870 8789
rect 1824 8721 1870 8723
rect 1824 8687 1830 8721
rect 1864 8687 1870 8721
rect 1824 8685 1870 8687
rect 1824 8619 1830 8685
rect 1864 8619 1870 8685
rect 1824 8613 1870 8619
rect 1824 8551 1830 8613
rect 1864 8551 1870 8613
rect 1824 8541 1870 8551
rect 1824 8483 1830 8541
rect 1864 8483 1870 8541
rect 1824 8469 1870 8483
rect 1824 8415 1830 8469
rect 1864 8415 1870 8469
rect 1824 8397 1870 8415
rect 1824 8347 1830 8397
rect 1864 8347 1870 8397
rect 1824 8325 1870 8347
rect 1824 8279 1830 8325
rect 1864 8279 1870 8325
rect 1824 8253 1870 8279
rect 1824 8211 1830 8253
rect 1864 8211 1870 8253
rect 1824 8181 1870 8211
rect 1824 8143 1830 8181
rect 1864 8143 1870 8181
rect 1824 8109 1870 8143
rect 1824 8075 1830 8109
rect 1864 8075 1870 8109
rect 1824 8041 1870 8075
rect 1824 8003 1830 8041
rect 1864 8003 1870 8041
rect 1824 7973 1870 8003
rect 1824 7931 1830 7973
rect 1864 7931 1870 7973
rect 1824 7905 1870 7931
rect 1824 7859 1830 7905
rect 1864 7859 1870 7905
rect 1824 7837 1870 7859
rect 1824 7787 1830 7837
rect 1864 7787 1870 7837
rect 1824 7769 1870 7787
rect 1824 7715 1830 7769
rect 1864 7715 1870 7769
rect 1824 7701 1870 7715
rect 1824 7643 1830 7701
rect 1864 7643 1870 7701
rect 1824 7633 1870 7643
rect 1824 7571 1830 7633
rect 1864 7571 1870 7633
rect 1824 7565 1870 7571
rect 1824 7499 1830 7565
rect 1864 7499 1870 7565
rect 1824 7497 1870 7499
rect 1824 7463 1830 7497
rect 1864 7463 1870 7497
rect 1824 7461 1870 7463
rect 1824 7395 1830 7461
rect 1864 7395 1870 7461
rect 1824 7389 1870 7395
rect 1824 7327 1830 7389
rect 1864 7327 1870 7389
rect 1824 7317 1870 7327
rect 1824 7259 1830 7317
rect 1864 7259 1870 7317
rect 1824 7245 1870 7259
rect 1824 7191 1830 7245
rect 1864 7191 1870 7245
rect 1824 7173 1870 7191
rect 1824 7123 1830 7173
rect 1864 7123 1870 7173
rect 1824 7101 1870 7123
rect 1824 7055 1830 7101
rect 1864 7055 1870 7101
rect 1824 7029 1870 7055
rect 1824 6987 1830 7029
rect 1864 6987 1870 7029
rect 1824 6957 1870 6987
rect 1824 6919 1830 6957
rect 1864 6919 1870 6957
rect 1824 6885 1870 6919
rect 1824 6851 1830 6885
rect 1864 6851 1870 6885
rect 1824 6817 1870 6851
rect 1824 6779 1830 6817
rect 1864 6779 1870 6817
rect 1824 6749 1870 6779
rect 1824 6707 1830 6749
rect 1864 6707 1870 6749
rect 1824 6681 1870 6707
rect 1824 6635 1830 6681
rect 1864 6635 1870 6681
rect 1824 6613 1870 6635
rect 1824 6563 1830 6613
rect 1864 6563 1870 6613
rect 1824 6545 1870 6563
rect 1824 6491 1830 6545
rect 1864 6491 1870 6545
rect 1824 6477 1870 6491
rect 1824 6419 1830 6477
rect 1864 6419 1870 6477
rect 1824 6409 1870 6419
rect 1824 6347 1830 6409
rect 1864 6347 1870 6409
rect 1824 6341 1870 6347
rect 1824 6275 1830 6341
rect 1864 6275 1870 6341
rect 1824 6273 1870 6275
rect 1824 6239 1830 6273
rect 1864 6239 1870 6273
rect 1824 6237 1870 6239
rect 1824 6171 1830 6237
rect 1864 6171 1870 6237
rect 1824 6165 1870 6171
rect 1824 6103 1830 6165
rect 1864 6103 1870 6165
rect 1824 6093 1870 6103
rect 1824 6035 1830 6093
rect 1864 6035 1870 6093
rect 1824 6021 1870 6035
rect 1824 5967 1830 6021
rect 1864 5967 1870 6021
rect 1824 5949 1870 5967
rect 1824 5899 1830 5949
rect 1864 5899 1870 5949
rect 1824 5877 1870 5899
rect 1824 5831 1830 5877
rect 1864 5831 1870 5877
rect 1824 5805 1870 5831
rect 1824 5763 1830 5805
rect 1864 5763 1870 5805
rect 1824 5733 1870 5763
rect 1824 5695 1830 5733
rect 1864 5695 1870 5733
rect 1824 5661 1870 5695
rect 1824 5627 1830 5661
rect 1864 5627 1870 5661
rect 1824 5593 1870 5627
rect 1824 5555 1830 5593
rect 1864 5555 1870 5593
rect 1824 5525 1870 5555
rect 1824 5483 1830 5525
rect 1864 5483 1870 5525
rect 1824 5457 1870 5483
rect 1824 5411 1830 5457
rect 1864 5411 1870 5457
rect 1824 5389 1870 5411
rect 1824 5339 1830 5389
rect 1864 5339 1870 5389
rect 1824 5321 1870 5339
rect 1824 5267 1830 5321
rect 1864 5267 1870 5321
rect 1824 5253 1870 5267
rect 1824 5195 1830 5253
rect 1864 5195 1870 5253
rect 1824 5185 1870 5195
rect 1824 5123 1830 5185
rect 1864 5123 1870 5185
rect 1824 5117 1870 5123
rect 1824 5051 1830 5117
rect 1864 5051 1870 5117
rect 1824 5049 1870 5051
rect 1824 5015 1830 5049
rect 1864 5015 1870 5049
rect 1824 5013 1870 5015
rect 1824 4947 1830 5013
rect 1864 4947 1870 5013
rect 1824 4941 1870 4947
rect 1824 4879 1830 4941
rect 1864 4879 1870 4941
rect 1824 4869 1870 4879
rect 1824 4811 1830 4869
rect 1864 4811 1870 4869
rect 1824 4797 1870 4811
rect 1824 4743 1830 4797
rect 1864 4743 1870 4797
rect 1824 4725 1870 4743
rect 1824 4675 1830 4725
rect 1864 4675 1870 4725
rect 1824 4653 1870 4675
rect 1824 4607 1830 4653
rect 1864 4607 1870 4653
rect 1824 4581 1870 4607
rect 1824 4539 1830 4581
rect 1864 4539 1870 4581
rect 1824 4509 1870 4539
rect 1824 4471 1830 4509
rect 1864 4471 1870 4509
rect 1824 4437 1870 4471
rect 1824 4403 1830 4437
rect 1864 4403 1870 4437
rect 1824 4369 1870 4403
rect 1824 4331 1830 4369
rect 1864 4331 1870 4369
rect 1824 4301 1870 4331
rect 1824 4259 1830 4301
rect 1864 4259 1870 4301
rect 1824 4233 1870 4259
rect 1824 4187 1830 4233
rect 1864 4187 1870 4233
rect 1824 4165 1870 4187
rect 1824 4115 1830 4165
rect 1864 4115 1870 4165
rect 1824 4097 1870 4115
rect 1824 4043 1830 4097
rect 1864 4043 1870 4097
rect 1824 4029 1870 4043
rect 1824 3971 1830 4029
rect 1864 3971 1870 4029
rect 1824 3961 1870 3971
rect 1824 3899 1830 3961
rect 1864 3899 1870 3961
rect 1824 3893 1870 3899
rect 1824 3827 1830 3893
rect 1864 3827 1870 3893
rect 1824 3825 1870 3827
rect 1824 3791 1830 3825
rect 1864 3791 1870 3825
rect 1824 3789 1870 3791
rect 1824 3723 1830 3789
rect 1864 3723 1870 3789
rect 1824 3717 1870 3723
rect 1824 3655 1830 3717
rect 1864 3655 1870 3717
rect 1824 3645 1870 3655
rect 1824 3587 1830 3645
rect 1864 3587 1870 3645
rect 1824 3573 1870 3587
rect 1824 3519 1830 3573
rect 1864 3519 1870 3573
rect 1824 3501 1870 3519
rect -258 3465 -212 3467
rect -258 3431 -252 3465
rect -218 3431 -212 3465
rect -258 3429 -212 3431
rect -258 3363 -252 3429
rect -218 3363 -212 3429
rect -258 3357 -212 3363
rect -142 3452 -126 3472
rect -92 3452 -76 3472
rect -142 3414 -76 3452
rect -142 3360 -126 3414
rect -92 3360 -76 3414
rect -24 3452 -8 3472
rect 26 3452 42 3472
rect -24 3414 42 3452
rect -24 3360 -8 3414
rect 26 3360 42 3414
rect 94 3452 110 3472
rect 144 3452 160 3472
rect 94 3414 160 3452
rect 94 3360 110 3414
rect 144 3360 160 3414
rect 212 3452 228 3472
rect 262 3452 278 3472
rect 212 3414 278 3452
rect 212 3360 228 3414
rect 262 3360 278 3414
rect 330 3452 346 3472
rect 380 3452 396 3472
rect 330 3414 396 3452
rect 330 3360 346 3414
rect 380 3360 396 3414
rect 448 3452 464 3472
rect 498 3452 514 3472
rect 448 3414 514 3452
rect 448 3360 464 3414
rect 498 3360 514 3414
rect 566 3452 582 3472
rect 616 3452 632 3472
rect 566 3414 632 3452
rect 566 3360 582 3414
rect 616 3360 632 3414
rect 684 3452 700 3472
rect 734 3452 750 3472
rect 684 3414 750 3452
rect 684 3360 700 3414
rect 734 3360 750 3414
rect 802 3452 818 3472
rect 852 3452 868 3472
rect 802 3414 868 3452
rect 802 3360 818 3414
rect 852 3360 868 3414
rect 920 3452 936 3472
rect 970 3452 986 3472
rect 920 3414 986 3452
rect 920 3360 936 3414
rect 970 3360 986 3414
rect 1038 3452 1054 3472
rect 1088 3452 1104 3472
rect 1038 3414 1104 3452
rect 1038 3360 1054 3414
rect 1088 3360 1104 3414
rect 1156 3452 1172 3472
rect 1206 3452 1222 3472
rect 1156 3414 1222 3452
rect 1156 3360 1172 3414
rect 1206 3360 1222 3414
rect 1274 3452 1290 3472
rect 1324 3452 1340 3472
rect 1274 3414 1340 3452
rect 1274 3360 1290 3414
rect 1324 3360 1340 3414
rect 1392 3452 1408 3472
rect 1442 3452 1458 3472
rect 1392 3414 1458 3452
rect 1392 3360 1408 3414
rect 1442 3360 1458 3414
rect 1510 3452 1526 3472
rect 1560 3452 1576 3472
rect 1510 3414 1576 3452
rect 1510 3360 1526 3414
rect 1560 3360 1576 3414
rect 1628 3452 1644 3472
rect 1678 3452 1694 3472
rect 1628 3414 1694 3452
rect 1628 3360 1644 3414
rect 1678 3360 1694 3414
rect 1824 3451 1830 3501
rect 1864 3451 1870 3501
rect 3966 38689 4012 38717
rect 3966 38651 3972 38689
rect 4006 38651 4012 38689
rect 3966 38621 4012 38651
rect 3966 38578 3972 38621
rect 4006 38578 4012 38621
rect 3966 38553 4012 38578
rect 3966 38505 3972 38553
rect 4006 38505 4012 38553
rect 3966 38485 4012 38505
rect 3966 38432 3972 38485
rect 4006 38432 4012 38485
rect 3966 38417 4012 38432
rect 3966 38359 3972 38417
rect 4006 38359 4012 38417
rect 3966 38349 4012 38359
rect 3966 38286 3972 38349
rect 4006 38286 4012 38349
rect 3966 38281 4012 38286
rect 3966 38179 3972 38281
rect 4006 38179 4012 38281
rect 3966 38174 4012 38179
rect 3966 38111 3972 38174
rect 4006 38111 4012 38174
rect 3966 38101 4012 38111
rect 3966 38043 3972 38101
rect 4006 38043 4012 38101
rect 3966 38028 4012 38043
rect 3966 37975 3972 38028
rect 4006 37975 4012 38028
rect 3966 37955 4012 37975
rect 3966 37907 3972 37955
rect 4006 37907 4012 37955
rect 3966 37882 4012 37907
rect 3966 37839 3972 37882
rect 4006 37839 4012 37882
rect 3966 37809 4012 37839
rect 3966 37771 3972 37809
rect 4006 37771 4012 37809
rect 3966 37737 4012 37771
rect 3966 37702 3972 37737
rect 4006 37702 4012 37737
rect 3966 37669 4012 37702
rect 3966 37629 3972 37669
rect 4006 37629 4012 37669
rect 3966 37601 4012 37629
rect 3966 37556 3972 37601
rect 4006 37556 4012 37601
rect 3966 37533 4012 37556
rect 3966 37483 3972 37533
rect 4006 37483 4012 37533
rect 3966 37465 4012 37483
rect 3966 37410 3972 37465
rect 4006 37410 4012 37465
rect 3966 37397 4012 37410
rect 3966 37337 3972 37397
rect 4006 37337 4012 37397
rect 3966 37329 4012 37337
rect 3966 37264 3972 37329
rect 4006 37264 4012 37329
rect 3966 37261 4012 37264
rect 3966 37227 3972 37261
rect 4006 37227 4012 37261
rect 3966 37225 4012 37227
rect 3966 37159 3972 37225
rect 4006 37159 4012 37225
rect 3966 37152 4012 37159
rect 3966 37091 3972 37152
rect 4006 37091 4012 37152
rect 3966 37079 4012 37091
rect 3966 37023 3972 37079
rect 4006 37023 4012 37079
rect 3966 37006 4012 37023
rect 3966 36955 3972 37006
rect 4006 36955 4012 37006
rect 3966 36933 4012 36955
rect 3966 36887 3972 36933
rect 4006 36887 4012 36933
rect 3966 36860 4012 36887
rect 3966 36819 3972 36860
rect 4006 36819 4012 36860
rect 3966 36787 4012 36819
rect 3966 36751 3972 36787
rect 4006 36751 4012 36787
rect 3966 36717 4012 36751
rect 3966 36680 3972 36717
rect 4006 36680 4012 36717
rect 3966 36649 4012 36680
rect 3966 36607 3972 36649
rect 4006 36607 4012 36649
rect 3966 36581 4012 36607
rect 3966 36534 3972 36581
rect 4006 36534 4012 36581
rect 3966 36513 4012 36534
rect 3966 36461 3972 36513
rect 4006 36461 4012 36513
rect 3966 36445 4012 36461
rect 3966 36388 3972 36445
rect 4006 36388 4012 36445
rect 3966 36377 4012 36388
rect 3966 36315 3972 36377
rect 4006 36315 4012 36377
rect 3966 36309 4012 36315
rect 3966 36242 3972 36309
rect 4006 36242 4012 36309
rect 3966 36241 4012 36242
rect 3966 36207 3972 36241
rect 4006 36207 4012 36241
rect 3966 36203 4012 36207
rect 3966 36139 3972 36203
rect 4006 36139 4012 36203
rect 3966 36130 4012 36139
rect 3966 36071 3972 36130
rect 4006 36071 4012 36130
rect 3966 36057 4012 36071
rect 3966 36003 3972 36057
rect 4006 36003 4012 36057
rect 3966 35984 4012 36003
rect 3966 35935 3972 35984
rect 4006 35935 4012 35984
rect 3966 35911 4012 35935
rect 3966 35867 3972 35911
rect 4006 35867 4012 35911
rect 3966 35838 4012 35867
rect 3966 35799 3972 35838
rect 4006 35799 4012 35838
rect 3966 35765 4012 35799
rect 3966 35731 3972 35765
rect 4006 35731 4012 35765
rect 3966 35697 4012 35731
rect 3966 35658 3972 35697
rect 4006 35658 4012 35697
rect 3966 35629 4012 35658
rect 3966 35585 3972 35629
rect 4006 35585 4012 35629
rect 3966 35561 4012 35585
rect 3966 35512 3972 35561
rect 4006 35512 4012 35561
rect 3966 35493 4012 35512
rect 3966 35439 3972 35493
rect 4006 35439 4012 35493
rect 3966 35425 4012 35439
rect 3966 35366 3972 35425
rect 4006 35366 4012 35425
rect 3966 35357 4012 35366
rect 3966 35293 3972 35357
rect 4006 35293 4012 35357
rect 3966 35289 4012 35293
rect 3966 35255 3972 35289
rect 4006 35255 4012 35289
rect 3966 35254 4012 35255
rect 3966 35187 3972 35254
rect 4006 35187 4012 35254
rect 3966 35181 4012 35187
rect 3966 35119 3972 35181
rect 4006 35119 4012 35181
rect 3966 35109 4012 35119
rect 3966 35051 3972 35109
rect 4006 35051 4012 35109
rect 3966 35037 4012 35051
rect 3966 34983 3972 35037
rect 4006 34983 4012 35037
rect 3966 34965 4012 34983
rect 3966 34915 3972 34965
rect 4006 34915 4012 34965
rect 3966 34893 4012 34915
rect 3966 34847 3972 34893
rect 4006 34847 4012 34893
rect 3966 34821 4012 34847
rect 3966 34779 3972 34821
rect 4006 34779 4012 34821
rect 3966 34749 4012 34779
rect 3966 34711 3972 34749
rect 4006 34711 4012 34749
rect 3966 34677 4012 34711
rect 3966 34643 3972 34677
rect 4006 34643 4012 34677
rect 3966 34609 4012 34643
rect 3966 34571 3972 34609
rect 4006 34571 4012 34609
rect 3966 34541 4012 34571
rect 3966 34499 3972 34541
rect 4006 34499 4012 34541
rect 3966 34473 4012 34499
rect 3966 34427 3972 34473
rect 4006 34427 4012 34473
rect 3966 34405 4012 34427
rect 3966 34355 3972 34405
rect 4006 34355 4012 34405
rect 3966 34337 4012 34355
rect 3966 34283 3972 34337
rect 4006 34283 4012 34337
rect 3966 34269 4012 34283
rect 3966 34211 3972 34269
rect 4006 34211 4012 34269
rect 3966 34201 4012 34211
rect 3966 34139 3972 34201
rect 4006 34139 4012 34201
rect 3966 34133 4012 34139
rect 3966 34067 3972 34133
rect 4006 34067 4012 34133
rect 3966 34065 4012 34067
rect 3966 34031 3972 34065
rect 4006 34031 4012 34065
rect 3966 34029 4012 34031
rect 3966 33963 3972 34029
rect 4006 33963 4012 34029
rect 3966 33957 4012 33963
rect 3966 33895 3972 33957
rect 4006 33895 4012 33957
rect 3966 33885 4012 33895
rect 3966 33827 3972 33885
rect 4006 33827 4012 33885
rect 3966 33813 4012 33827
rect 3966 33759 3972 33813
rect 4006 33759 4012 33813
rect 3966 33741 4012 33759
rect 3966 33691 3972 33741
rect 4006 33691 4012 33741
rect 3966 33669 4012 33691
rect 3966 33623 3972 33669
rect 4006 33623 4012 33669
rect 3966 33597 4012 33623
rect 3966 33555 3972 33597
rect 4006 33555 4012 33597
rect 3966 33525 4012 33555
rect 3966 33487 3972 33525
rect 4006 33487 4012 33525
rect 3966 33453 4012 33487
rect 3966 33419 3972 33453
rect 4006 33419 4012 33453
rect 3966 33385 4012 33419
rect 3966 33347 3972 33385
rect 4006 33347 4012 33385
rect 3966 33317 4012 33347
rect 3966 33275 3972 33317
rect 4006 33275 4012 33317
rect 3966 33249 4012 33275
rect 3966 33203 3972 33249
rect 4006 33203 4012 33249
rect 3966 33181 4012 33203
rect 3966 33131 3972 33181
rect 4006 33131 4012 33181
rect 3966 33113 4012 33131
rect 3966 33059 3972 33113
rect 4006 33059 4012 33113
rect 3966 33045 4012 33059
rect 3966 32987 3972 33045
rect 4006 32987 4012 33045
rect 3966 32977 4012 32987
rect 3966 32915 3972 32977
rect 4006 32915 4012 32977
rect 3966 32909 4012 32915
rect 3966 32843 3972 32909
rect 4006 32843 4012 32909
rect 3966 32841 4012 32843
rect 3966 32807 3972 32841
rect 4006 32807 4012 32841
rect 3966 32805 4012 32807
rect 3966 32739 3972 32805
rect 4006 32739 4012 32805
rect 3966 32733 4012 32739
rect 3966 32671 3972 32733
rect 4006 32671 4012 32733
rect 3966 32661 4012 32671
rect 3966 32603 3972 32661
rect 4006 32603 4012 32661
rect 3966 32589 4012 32603
rect 3966 32535 3972 32589
rect 4006 32535 4012 32589
rect 3966 32517 4012 32535
rect 3966 32467 3972 32517
rect 4006 32467 4012 32517
rect 3966 32445 4012 32467
rect 3966 32399 3972 32445
rect 4006 32399 4012 32445
rect 3966 32373 4012 32399
rect 3966 32331 3972 32373
rect 4006 32331 4012 32373
rect 3966 32301 4012 32331
rect 3966 32263 3972 32301
rect 4006 32263 4012 32301
rect 3966 32229 4012 32263
rect 3966 32195 3972 32229
rect 4006 32195 4012 32229
rect 3966 32161 4012 32195
rect 3966 32123 3972 32161
rect 4006 32123 4012 32161
rect 3966 32093 4012 32123
rect 3966 32051 3972 32093
rect 4006 32051 4012 32093
rect 3966 32025 4012 32051
rect 3966 31979 3972 32025
rect 4006 31979 4012 32025
rect 3966 31957 4012 31979
rect 3966 31907 3972 31957
rect 4006 31907 4012 31957
rect 3966 31889 4012 31907
rect 3966 31835 3972 31889
rect 4006 31835 4012 31889
rect 3966 31821 4012 31835
rect 3966 31763 3972 31821
rect 4006 31763 4012 31821
rect 3966 31753 4012 31763
rect 3966 31691 3972 31753
rect 4006 31691 4012 31753
rect 3966 31685 4012 31691
rect 3966 31619 3972 31685
rect 4006 31619 4012 31685
rect 3966 31617 4012 31619
rect 3966 31583 3972 31617
rect 4006 31583 4012 31617
rect 3966 31581 4012 31583
rect 3966 31515 3972 31581
rect 4006 31515 4012 31581
rect 3966 31509 4012 31515
rect 3966 31447 3972 31509
rect 4006 31447 4012 31509
rect 3966 31437 4012 31447
rect 3966 31379 3972 31437
rect 4006 31379 4012 31437
rect 3966 31365 4012 31379
rect 3966 31311 3972 31365
rect 4006 31311 4012 31365
rect 3966 31293 4012 31311
rect 3966 31243 3972 31293
rect 4006 31243 4012 31293
rect 3966 31221 4012 31243
rect 3966 31175 3972 31221
rect 4006 31175 4012 31221
rect 3966 31149 4012 31175
rect 3966 31107 3972 31149
rect 4006 31107 4012 31149
rect 3966 31077 4012 31107
rect 3966 31039 3972 31077
rect 4006 31039 4012 31077
rect 3966 31005 4012 31039
rect 3966 30971 3972 31005
rect 4006 30971 4012 31005
rect 3966 30937 4012 30971
rect 3966 30899 3972 30937
rect 4006 30899 4012 30937
rect 3966 30869 4012 30899
rect 3966 30827 3972 30869
rect 4006 30827 4012 30869
rect 3966 30801 4012 30827
rect 3966 30755 3972 30801
rect 4006 30755 4012 30801
rect 3966 30733 4012 30755
rect 3966 30683 3972 30733
rect 4006 30683 4012 30733
rect 3966 30665 4012 30683
rect 3966 30611 3972 30665
rect 4006 30611 4012 30665
rect 3966 30597 4012 30611
rect 3966 30539 3972 30597
rect 4006 30539 4012 30597
rect 3966 30529 4012 30539
rect 3966 30467 3972 30529
rect 4006 30467 4012 30529
rect 3966 30461 4012 30467
rect 3966 30395 3972 30461
rect 4006 30395 4012 30461
rect 3966 30393 4012 30395
rect 3966 30359 3972 30393
rect 4006 30359 4012 30393
rect 3966 30357 4012 30359
rect 3966 30291 3972 30357
rect 4006 30291 4012 30357
rect 3966 30285 4012 30291
rect 3966 30223 3972 30285
rect 4006 30223 4012 30285
rect 3966 30213 4012 30223
rect 3966 30155 3972 30213
rect 4006 30155 4012 30213
rect 3966 30141 4012 30155
rect 3966 30087 3972 30141
rect 4006 30087 4012 30141
rect 3966 30069 4012 30087
rect 3966 30019 3972 30069
rect 4006 30019 4012 30069
rect 3966 29997 4012 30019
rect 3966 29951 3972 29997
rect 4006 29951 4012 29997
rect 3966 29925 4012 29951
rect 3966 29883 3972 29925
rect 4006 29883 4012 29925
rect 3966 29853 4012 29883
rect 3966 29815 3972 29853
rect 4006 29815 4012 29853
rect 3966 29781 4012 29815
rect 3966 29747 3972 29781
rect 4006 29747 4012 29781
rect 3966 29713 4012 29747
rect 3966 29675 3972 29713
rect 4006 29675 4012 29713
rect 3966 29645 4012 29675
rect 3966 29603 3972 29645
rect 4006 29603 4012 29645
rect 3966 29577 4012 29603
rect 3966 29531 3972 29577
rect 4006 29531 4012 29577
rect 3966 29509 4012 29531
rect 3966 29459 3972 29509
rect 4006 29459 4012 29509
rect 3966 29441 4012 29459
rect 3966 29387 3972 29441
rect 4006 29387 4012 29441
rect 3966 29373 4012 29387
rect 3966 29315 3972 29373
rect 4006 29315 4012 29373
rect 3966 29305 4012 29315
rect 3966 29243 3972 29305
rect 4006 29243 4012 29305
rect 3966 29237 4012 29243
rect 3966 29171 3972 29237
rect 4006 29171 4012 29237
rect 3966 29169 4012 29171
rect 3966 29135 3972 29169
rect 4006 29135 4012 29169
rect 3966 29133 4012 29135
rect 3966 29067 3972 29133
rect 4006 29067 4012 29133
rect 3966 29061 4012 29067
rect 3966 28999 3972 29061
rect 4006 28999 4012 29061
rect 3966 28989 4012 28999
rect 3966 28931 3972 28989
rect 4006 28931 4012 28989
rect 3966 28917 4012 28931
rect 3966 28863 3972 28917
rect 4006 28863 4012 28917
rect 3966 28845 4012 28863
rect 3966 28795 3972 28845
rect 4006 28795 4012 28845
rect 3966 28773 4012 28795
rect 3966 28727 3972 28773
rect 4006 28727 4012 28773
rect 3966 28701 4012 28727
rect 3966 28659 3972 28701
rect 4006 28659 4012 28701
rect 3966 28629 4012 28659
rect 3966 28591 3972 28629
rect 4006 28591 4012 28629
rect 3966 28557 4012 28591
rect 3966 28523 3972 28557
rect 4006 28523 4012 28557
rect 3966 28489 4012 28523
rect 3966 28451 3972 28489
rect 4006 28451 4012 28489
rect 3966 28421 4012 28451
rect 3966 28379 3972 28421
rect 4006 28379 4012 28421
rect 3966 28353 4012 28379
rect 3966 28307 3972 28353
rect 4006 28307 4012 28353
rect 3966 28285 4012 28307
rect 3966 28235 3972 28285
rect 4006 28235 4012 28285
rect 3966 28217 4012 28235
rect 3966 28163 3972 28217
rect 4006 28163 4012 28217
rect 3966 28149 4012 28163
rect 3966 28091 3972 28149
rect 4006 28091 4012 28149
rect 3966 28081 4012 28091
rect 3966 28019 3972 28081
rect 4006 28019 4012 28081
rect 3966 28013 4012 28019
rect 3966 27947 3972 28013
rect 4006 27947 4012 28013
rect 3966 27945 4012 27947
rect 3966 27911 3972 27945
rect 4006 27911 4012 27945
rect 3966 27909 4012 27911
rect 3966 27843 3972 27909
rect 4006 27843 4012 27909
rect 3966 27837 4012 27843
rect 3966 27775 3972 27837
rect 4006 27775 4012 27837
rect 3966 27765 4012 27775
rect 3966 27707 3972 27765
rect 4006 27707 4012 27765
rect 3966 27693 4012 27707
rect 3966 27639 3972 27693
rect 4006 27639 4012 27693
rect 3966 27621 4012 27639
rect 3966 27571 3972 27621
rect 4006 27571 4012 27621
rect 3966 27549 4012 27571
rect 3966 27503 3972 27549
rect 4006 27503 4012 27549
rect 3966 27477 4012 27503
rect 3966 27435 3972 27477
rect 4006 27435 4012 27477
rect 3966 27405 4012 27435
rect 3966 27367 3972 27405
rect 4006 27367 4012 27405
rect 3966 27333 4012 27367
rect 3966 27299 3972 27333
rect 4006 27299 4012 27333
rect 3966 27265 4012 27299
rect 3966 27227 3972 27265
rect 4006 27227 4012 27265
rect 3966 27197 4012 27227
rect 3966 27155 3972 27197
rect 4006 27155 4012 27197
rect 3966 27129 4012 27155
rect 3966 27083 3972 27129
rect 4006 27083 4012 27129
rect 3966 27061 4012 27083
rect 3966 27011 3972 27061
rect 4006 27011 4012 27061
rect 3966 26993 4012 27011
rect 3966 26939 3972 26993
rect 4006 26939 4012 26993
rect 3966 26925 4012 26939
rect 3966 26867 3972 26925
rect 4006 26867 4012 26925
rect 3966 26857 4012 26867
rect 3966 26795 3972 26857
rect 4006 26795 4012 26857
rect 3966 26789 4012 26795
rect 3966 26723 3972 26789
rect 4006 26723 4012 26789
rect 3966 26721 4012 26723
rect 3966 26687 3972 26721
rect 4006 26687 4012 26721
rect 3966 26685 4012 26687
rect 3966 26619 3972 26685
rect 4006 26619 4012 26685
rect 3966 26613 4012 26619
rect 3966 26551 3972 26613
rect 4006 26551 4012 26613
rect 3966 26541 4012 26551
rect 3966 26483 3972 26541
rect 4006 26483 4012 26541
rect 3966 26469 4012 26483
rect 3966 26415 3972 26469
rect 4006 26415 4012 26469
rect 3966 26397 4012 26415
rect 3966 26347 3972 26397
rect 4006 26347 4012 26397
rect 3966 26325 4012 26347
rect 3966 26279 3972 26325
rect 4006 26279 4012 26325
rect 3966 26253 4012 26279
rect 3966 26211 3972 26253
rect 4006 26211 4012 26253
rect 3966 26181 4012 26211
rect 3966 26143 3972 26181
rect 4006 26143 4012 26181
rect 3966 26109 4012 26143
rect 3966 26075 3972 26109
rect 4006 26075 4012 26109
rect 3966 26041 4012 26075
rect 3966 26003 3972 26041
rect 4006 26003 4012 26041
rect 3966 25973 4012 26003
rect 3966 25931 3972 25973
rect 4006 25931 4012 25973
rect 3966 25905 4012 25931
rect 3966 25859 3972 25905
rect 4006 25859 4012 25905
rect 3966 25837 4012 25859
rect 3966 25787 3972 25837
rect 4006 25787 4012 25837
rect 3966 25769 4012 25787
rect 3966 25715 3972 25769
rect 4006 25715 4012 25769
rect 3966 25701 4012 25715
rect 3966 25643 3972 25701
rect 4006 25643 4012 25701
rect 3966 25633 4012 25643
rect 3966 25571 3972 25633
rect 4006 25571 4012 25633
rect 3966 25565 4012 25571
rect 3966 25499 3972 25565
rect 4006 25499 4012 25565
rect 3966 25497 4012 25499
rect 3966 25463 3972 25497
rect 4006 25463 4012 25497
rect 3966 25461 4012 25463
rect 3966 25395 3972 25461
rect 4006 25395 4012 25461
rect 3966 25389 4012 25395
rect 3966 25327 3972 25389
rect 4006 25327 4012 25389
rect 3966 25317 4012 25327
rect 3966 25259 3972 25317
rect 4006 25259 4012 25317
rect 3966 25245 4012 25259
rect 3966 25191 3972 25245
rect 4006 25191 4012 25245
rect 3966 25173 4012 25191
rect 3966 25123 3972 25173
rect 4006 25123 4012 25173
rect 3966 25101 4012 25123
rect 3966 25055 3972 25101
rect 4006 25055 4012 25101
rect 3966 25029 4012 25055
rect 3966 24987 3972 25029
rect 4006 24987 4012 25029
rect 3966 24957 4012 24987
rect 3966 24919 3972 24957
rect 4006 24919 4012 24957
rect 3966 24885 4012 24919
rect 3966 24851 3972 24885
rect 4006 24851 4012 24885
rect 3966 24817 4012 24851
rect 3966 24779 3972 24817
rect 4006 24779 4012 24817
rect 3966 24749 4012 24779
rect 3966 24707 3972 24749
rect 4006 24707 4012 24749
rect 3966 24681 4012 24707
rect 3966 24635 3972 24681
rect 4006 24635 4012 24681
rect 3966 24613 4012 24635
rect 3966 24563 3972 24613
rect 4006 24563 4012 24613
rect 3966 24545 4012 24563
rect 3966 24491 3972 24545
rect 4006 24491 4012 24545
rect 3966 24477 4012 24491
rect 3966 24419 3972 24477
rect 4006 24419 4012 24477
rect 3966 24409 4012 24419
rect 3966 24347 3972 24409
rect 4006 24347 4012 24409
rect 3966 24341 4012 24347
rect 3966 24275 3972 24341
rect 4006 24275 4012 24341
rect 3966 24273 4012 24275
rect 3966 24239 3972 24273
rect 4006 24239 4012 24273
rect 3966 24237 4012 24239
rect 3966 24171 3972 24237
rect 4006 24171 4012 24237
rect 3966 24165 4012 24171
rect 3966 24103 3972 24165
rect 4006 24103 4012 24165
rect 3966 24093 4012 24103
rect 3966 24035 3972 24093
rect 4006 24035 4012 24093
rect 3966 24021 4012 24035
rect 3966 23967 3972 24021
rect 4006 23967 4012 24021
rect 3966 23949 4012 23967
rect 3966 23899 3972 23949
rect 4006 23899 4012 23949
rect 3966 23877 4012 23899
rect 3966 23831 3972 23877
rect 4006 23831 4012 23877
rect 3966 23805 4012 23831
rect 3966 23763 3972 23805
rect 4006 23763 4012 23805
rect 3966 23733 4012 23763
rect 3966 23695 3972 23733
rect 4006 23695 4012 23733
rect 3966 23661 4012 23695
rect 3966 23627 3972 23661
rect 4006 23627 4012 23661
rect 3966 23593 4012 23627
rect 3966 23555 3972 23593
rect 4006 23555 4012 23593
rect 3966 23525 4012 23555
rect 3966 23483 3972 23525
rect 4006 23483 4012 23525
rect 3966 23457 4012 23483
rect 3966 23411 3972 23457
rect 4006 23411 4012 23457
rect 3966 23389 4012 23411
rect 3966 23339 3972 23389
rect 4006 23339 4012 23389
rect 3966 23321 4012 23339
rect 3966 23267 3972 23321
rect 4006 23267 4012 23321
rect 3966 23253 4012 23267
rect 3966 23195 3972 23253
rect 4006 23195 4012 23253
rect 3966 23185 4012 23195
rect 3966 23123 3972 23185
rect 4006 23123 4012 23185
rect 3966 23117 4012 23123
rect 3966 23051 3972 23117
rect 4006 23051 4012 23117
rect 3966 23049 4012 23051
rect 3966 23015 3972 23049
rect 4006 23015 4012 23049
rect 3966 23013 4012 23015
rect 3966 22947 3972 23013
rect 4006 22947 4012 23013
rect 3966 22941 4012 22947
rect 3966 22879 3972 22941
rect 4006 22879 4012 22941
rect 3966 22869 4012 22879
rect 3966 22811 3972 22869
rect 4006 22811 4012 22869
rect 3966 22797 4012 22811
rect 3966 22743 3972 22797
rect 4006 22743 4012 22797
rect 3966 22725 4012 22743
rect 3966 22675 3972 22725
rect 4006 22675 4012 22725
rect 3966 22653 4012 22675
rect 3966 22607 3972 22653
rect 4006 22607 4012 22653
rect 3966 22581 4012 22607
rect 3966 22539 3972 22581
rect 4006 22539 4012 22581
rect 3966 22509 4012 22539
rect 3966 22471 3972 22509
rect 4006 22471 4012 22509
rect 3966 22437 4012 22471
rect 3966 22403 3972 22437
rect 4006 22403 4012 22437
rect 3966 22369 4012 22403
rect 3966 22331 3972 22369
rect 4006 22331 4012 22369
rect 3966 22301 4012 22331
rect 3966 22259 3972 22301
rect 4006 22259 4012 22301
rect 3966 22233 4012 22259
rect 3966 22187 3972 22233
rect 4006 22187 4012 22233
rect 3966 22165 4012 22187
rect 3966 22115 3972 22165
rect 4006 22115 4012 22165
rect 3966 22097 4012 22115
rect 3966 22043 3972 22097
rect 4006 22043 4012 22097
rect 3966 22029 4012 22043
rect 3966 21971 3972 22029
rect 4006 21971 4012 22029
rect 3966 21961 4012 21971
rect 3966 21899 3972 21961
rect 4006 21899 4012 21961
rect 3966 21893 4012 21899
rect 3966 21827 3972 21893
rect 4006 21827 4012 21893
rect 3966 21825 4012 21827
rect 3966 21791 3972 21825
rect 4006 21791 4012 21825
rect 3966 21789 4012 21791
rect 3966 21723 3972 21789
rect 4006 21723 4012 21789
rect 3966 21717 4012 21723
rect 3966 21655 3972 21717
rect 4006 21655 4012 21717
rect 3966 21645 4012 21655
rect 3966 21587 3972 21645
rect 4006 21587 4012 21645
rect 3966 21573 4012 21587
rect 3966 21519 3972 21573
rect 4006 21519 4012 21573
rect 3966 21501 4012 21519
rect 3966 21451 3972 21501
rect 4006 21451 4012 21501
rect 3966 21429 4012 21451
rect 3966 21383 3972 21429
rect 4006 21383 4012 21429
rect 3966 21357 4012 21383
rect 3966 21315 3972 21357
rect 4006 21315 4012 21357
rect 3966 21285 4012 21315
rect 3966 21247 3972 21285
rect 4006 21247 4012 21285
rect 3966 21213 4012 21247
rect 3966 21179 3972 21213
rect 4006 21179 4012 21213
rect 3966 21145 4012 21179
rect 3966 21107 3972 21145
rect 4006 21107 4012 21145
rect 3966 21077 4012 21107
rect 3966 21035 3972 21077
rect 4006 21035 4012 21077
rect 3966 21009 4012 21035
rect 3966 20963 3972 21009
rect 4006 20963 4012 21009
rect 3966 20941 4012 20963
rect 3966 20891 3972 20941
rect 4006 20891 4012 20941
rect 3966 20873 4012 20891
rect 3966 20819 3972 20873
rect 4006 20819 4012 20873
rect 3966 20805 4012 20819
rect 3966 20747 3972 20805
rect 4006 20747 4012 20805
rect 3966 20737 4012 20747
rect 3966 20675 3972 20737
rect 4006 20675 4012 20737
rect 3966 20669 4012 20675
rect 3966 20603 3972 20669
rect 4006 20603 4012 20669
rect 3966 20601 4012 20603
rect 3966 20567 3972 20601
rect 4006 20567 4012 20601
rect 3966 20565 4012 20567
rect 3966 20499 3972 20565
rect 4006 20499 4012 20565
rect 3966 20493 4012 20499
rect 3966 20431 3972 20493
rect 4006 20431 4012 20493
rect 3966 20421 4012 20431
rect 3966 20363 3972 20421
rect 4006 20363 4012 20421
rect 3966 20349 4012 20363
rect 3966 20295 3972 20349
rect 4006 20295 4012 20349
rect 3966 20277 4012 20295
rect 3966 20227 3972 20277
rect 4006 20227 4012 20277
rect 3966 20205 4012 20227
rect 3966 20159 3972 20205
rect 4006 20159 4012 20205
rect 3966 20133 4012 20159
rect 3966 20091 3972 20133
rect 4006 20091 4012 20133
rect 3966 20061 4012 20091
rect 3966 20023 3972 20061
rect 4006 20023 4012 20061
rect 3966 19989 4012 20023
rect 3966 19955 3972 19989
rect 4006 19955 4012 19989
rect 3966 19921 4012 19955
rect 3966 19883 3972 19921
rect 4006 19883 4012 19921
rect 3966 19853 4012 19883
rect 3966 19811 3972 19853
rect 4006 19811 4012 19853
rect 3966 19785 4012 19811
rect 3966 19739 3972 19785
rect 4006 19739 4012 19785
rect 3966 19717 4012 19739
rect 3966 19667 3972 19717
rect 4006 19667 4012 19717
rect 3966 19649 4012 19667
rect 3966 19595 3972 19649
rect 4006 19595 4012 19649
rect 3966 19581 4012 19595
rect 3966 19523 3972 19581
rect 4006 19523 4012 19581
rect 3966 19513 4012 19523
rect 3966 19451 3972 19513
rect 4006 19451 4012 19513
rect 3966 19445 4012 19451
rect 3966 19379 3972 19445
rect 4006 19379 4012 19445
rect 3966 19377 4012 19379
rect 3966 19343 3972 19377
rect 4006 19343 4012 19377
rect 3966 19341 4012 19343
rect 3966 19275 3972 19341
rect 4006 19275 4012 19341
rect 3966 19269 4012 19275
rect 3966 19207 3972 19269
rect 4006 19207 4012 19269
rect 3966 19197 4012 19207
rect 3966 19139 3972 19197
rect 4006 19139 4012 19197
rect 3966 19125 4012 19139
rect 3966 19071 3972 19125
rect 4006 19071 4012 19125
rect 3966 19053 4012 19071
rect 3966 19003 3972 19053
rect 4006 19003 4012 19053
rect 3966 18981 4012 19003
rect 3966 18935 3972 18981
rect 4006 18935 4012 18981
rect 3966 18909 4012 18935
rect 3966 18867 3972 18909
rect 4006 18867 4012 18909
rect 3966 18837 4012 18867
rect 3966 18799 3972 18837
rect 4006 18799 4012 18837
rect 3966 18765 4012 18799
rect 3966 18731 3972 18765
rect 4006 18731 4012 18765
rect 3966 18697 4012 18731
rect 3966 18659 3972 18697
rect 4006 18659 4012 18697
rect 3966 18629 4012 18659
rect 3966 18587 3972 18629
rect 4006 18587 4012 18629
rect 3966 18561 4012 18587
rect 3966 18515 3972 18561
rect 4006 18515 4012 18561
rect 3966 18493 4012 18515
rect 3966 18443 3972 18493
rect 4006 18443 4012 18493
rect 3966 18425 4012 18443
rect 3966 18371 3972 18425
rect 4006 18371 4012 18425
rect 3966 18357 4012 18371
rect 3966 18299 3972 18357
rect 4006 18299 4012 18357
rect 3966 18289 4012 18299
rect 3966 18227 3972 18289
rect 4006 18227 4012 18289
rect 3966 18221 4012 18227
rect 3966 18155 3972 18221
rect 4006 18155 4012 18221
rect 3966 18153 4012 18155
rect 3966 18119 3972 18153
rect 4006 18119 4012 18153
rect 3966 18117 4012 18119
rect 3966 18051 3972 18117
rect 4006 18051 4012 18117
rect 3966 18045 4012 18051
rect 3966 17983 3972 18045
rect 4006 17983 4012 18045
rect 3966 17973 4012 17983
rect 3966 17915 3972 17973
rect 4006 17915 4012 17973
rect 3966 17901 4012 17915
rect 3966 17847 3972 17901
rect 4006 17847 4012 17901
rect 3966 17829 4012 17847
rect 3966 17779 3972 17829
rect 4006 17779 4012 17829
rect 3966 17757 4012 17779
rect 3966 17711 3972 17757
rect 4006 17711 4012 17757
rect 3966 17685 4012 17711
rect 3966 17643 3972 17685
rect 4006 17643 4012 17685
rect 3966 17613 4012 17643
rect 3966 17575 3972 17613
rect 4006 17575 4012 17613
rect 3966 17541 4012 17575
rect 3966 17507 3972 17541
rect 4006 17507 4012 17541
rect 3966 17473 4012 17507
rect 3966 17435 3972 17473
rect 4006 17435 4012 17473
rect 3966 17405 4012 17435
rect 3966 17363 3972 17405
rect 4006 17363 4012 17405
rect 3966 17337 4012 17363
rect 3966 17291 3972 17337
rect 4006 17291 4012 17337
rect 3966 17269 4012 17291
rect 3966 17219 3972 17269
rect 4006 17219 4012 17269
rect 3966 17201 4012 17219
rect 3966 17147 3972 17201
rect 4006 17147 4012 17201
rect 3966 17133 4012 17147
rect 3966 17075 3972 17133
rect 4006 17075 4012 17133
rect 3966 17065 4012 17075
rect 3966 17003 3972 17065
rect 4006 17003 4012 17065
rect 3966 16997 4012 17003
rect 3966 16931 3972 16997
rect 4006 16931 4012 16997
rect 3966 16929 4012 16931
rect 3966 16895 3972 16929
rect 4006 16895 4012 16929
rect 3966 16893 4012 16895
rect 3966 16827 3972 16893
rect 4006 16827 4012 16893
rect 3966 16821 4012 16827
rect 3966 16759 3972 16821
rect 4006 16759 4012 16821
rect 3966 16749 4012 16759
rect 3966 16691 3972 16749
rect 4006 16691 4012 16749
rect 3966 16677 4012 16691
rect 3966 16623 3972 16677
rect 4006 16623 4012 16677
rect 3966 16605 4012 16623
rect 3966 16555 3972 16605
rect 4006 16555 4012 16605
rect 3966 16533 4012 16555
rect 3966 16487 3972 16533
rect 4006 16487 4012 16533
rect 3966 16461 4012 16487
rect 3966 16419 3972 16461
rect 4006 16419 4012 16461
rect 3966 16389 4012 16419
rect 3966 16351 3972 16389
rect 4006 16351 4012 16389
rect 3966 16317 4012 16351
rect 3966 16283 3972 16317
rect 4006 16283 4012 16317
rect 3966 16249 4012 16283
rect 3966 16211 3972 16249
rect 4006 16211 4012 16249
rect 3966 16181 4012 16211
rect 3966 16139 3972 16181
rect 4006 16139 4012 16181
rect 3966 16113 4012 16139
rect 3966 16067 3972 16113
rect 4006 16067 4012 16113
rect 3966 16045 4012 16067
rect 3966 15995 3972 16045
rect 4006 15995 4012 16045
rect 3966 15977 4012 15995
rect 3966 15923 3972 15977
rect 4006 15923 4012 15977
rect 3966 15909 4012 15923
rect 3966 15851 3972 15909
rect 4006 15851 4012 15909
rect 3966 15841 4012 15851
rect 3966 15779 3972 15841
rect 4006 15779 4012 15841
rect 3966 15773 4012 15779
rect 3966 15707 3972 15773
rect 4006 15707 4012 15773
rect 3966 15705 4012 15707
rect 3966 15671 3972 15705
rect 4006 15671 4012 15705
rect 3966 15669 4012 15671
rect 3966 15603 3972 15669
rect 4006 15603 4012 15669
rect 3966 15597 4012 15603
rect 3966 15535 3972 15597
rect 4006 15535 4012 15597
rect 3966 15525 4012 15535
rect 3966 15467 3972 15525
rect 4006 15467 4012 15525
rect 3966 15453 4012 15467
rect 3966 15399 3972 15453
rect 4006 15399 4012 15453
rect 3966 15381 4012 15399
rect 3966 15331 3972 15381
rect 4006 15331 4012 15381
rect 3966 15309 4012 15331
rect 3966 15263 3972 15309
rect 4006 15263 4012 15309
rect 3966 15237 4012 15263
rect 3966 15195 3972 15237
rect 4006 15195 4012 15237
rect 3966 15165 4012 15195
rect 3966 15127 3972 15165
rect 4006 15127 4012 15165
rect 3966 15093 4012 15127
rect 3966 15059 3972 15093
rect 4006 15059 4012 15093
rect 3966 15025 4012 15059
rect 3966 14987 3972 15025
rect 4006 14987 4012 15025
rect 3966 14957 4012 14987
rect 3966 14915 3972 14957
rect 4006 14915 4012 14957
rect 3966 14889 4012 14915
rect 3966 14843 3972 14889
rect 4006 14843 4012 14889
rect 3966 14821 4012 14843
rect 3966 14771 3972 14821
rect 4006 14771 4012 14821
rect 3966 14753 4012 14771
rect 3966 14699 3972 14753
rect 4006 14699 4012 14753
rect 3966 14685 4012 14699
rect 3966 14627 3972 14685
rect 4006 14627 4012 14685
rect 3966 14617 4012 14627
rect 3966 14555 3972 14617
rect 4006 14555 4012 14617
rect 3966 14549 4012 14555
rect 3966 14483 3972 14549
rect 4006 14483 4012 14549
rect 3966 14481 4012 14483
rect 3966 14447 3972 14481
rect 4006 14447 4012 14481
rect 3966 14445 4012 14447
rect 3966 14379 3972 14445
rect 4006 14379 4012 14445
rect 3966 14373 4012 14379
rect 3966 14311 3972 14373
rect 4006 14311 4012 14373
rect 3966 14301 4012 14311
rect 3966 14243 3972 14301
rect 4006 14243 4012 14301
rect 3966 14229 4012 14243
rect 3966 14175 3972 14229
rect 4006 14175 4012 14229
rect 3966 14157 4012 14175
rect 3966 14107 3972 14157
rect 4006 14107 4012 14157
rect 3966 14085 4012 14107
rect 3966 14039 3972 14085
rect 4006 14039 4012 14085
rect 3966 14013 4012 14039
rect 3966 13971 3972 14013
rect 4006 13971 4012 14013
rect 3966 13941 4012 13971
rect 3966 13903 3972 13941
rect 4006 13903 4012 13941
rect 3966 13869 4012 13903
rect 3966 13835 3972 13869
rect 4006 13835 4012 13869
rect 3966 13801 4012 13835
rect 3966 13763 3972 13801
rect 4006 13763 4012 13801
rect 3966 13733 4012 13763
rect 3966 13691 3972 13733
rect 4006 13691 4012 13733
rect 3966 13665 4012 13691
rect 3966 13619 3972 13665
rect 4006 13619 4012 13665
rect 3966 13597 4012 13619
rect 3966 13547 3972 13597
rect 4006 13547 4012 13597
rect 3966 13529 4012 13547
rect 3966 13475 3972 13529
rect 4006 13475 4012 13529
rect 3966 13461 4012 13475
rect 3966 13403 3972 13461
rect 4006 13403 4012 13461
rect 3966 13393 4012 13403
rect 3966 13331 3972 13393
rect 4006 13331 4012 13393
rect 3966 13325 4012 13331
rect 3966 13259 3972 13325
rect 4006 13259 4012 13325
rect 3966 13257 4012 13259
rect 3966 13223 3972 13257
rect 4006 13223 4012 13257
rect 3966 13221 4012 13223
rect 3966 13155 3972 13221
rect 4006 13155 4012 13221
rect 3966 13149 4012 13155
rect 3966 13087 3972 13149
rect 4006 13087 4012 13149
rect 3966 13077 4012 13087
rect 3966 13019 3972 13077
rect 4006 13019 4012 13077
rect 3966 13005 4012 13019
rect 3966 12951 3972 13005
rect 4006 12951 4012 13005
rect 3966 12933 4012 12951
rect 3966 12883 3972 12933
rect 4006 12883 4012 12933
rect 3966 12861 4012 12883
rect 3966 12815 3972 12861
rect 4006 12815 4012 12861
rect 3966 12789 4012 12815
rect 3966 12747 3972 12789
rect 4006 12747 4012 12789
rect 3966 12717 4012 12747
rect 3966 12679 3972 12717
rect 4006 12679 4012 12717
rect 3966 12645 4012 12679
rect 3966 12611 3972 12645
rect 4006 12611 4012 12645
rect 3966 12577 4012 12611
rect 3966 12539 3972 12577
rect 4006 12539 4012 12577
rect 3966 12509 4012 12539
rect 3966 12467 3972 12509
rect 4006 12467 4012 12509
rect 3966 12441 4012 12467
rect 3966 12395 3972 12441
rect 4006 12395 4012 12441
rect 3966 12373 4012 12395
rect 3966 12323 3972 12373
rect 4006 12323 4012 12373
rect 3966 12305 4012 12323
rect 3966 12251 3972 12305
rect 4006 12251 4012 12305
rect 3966 12237 4012 12251
rect 3966 12179 3972 12237
rect 4006 12179 4012 12237
rect 3966 12169 4012 12179
rect 3966 12107 3972 12169
rect 4006 12107 4012 12169
rect 3966 12101 4012 12107
rect 3966 12035 3972 12101
rect 4006 12035 4012 12101
rect 3966 12033 4012 12035
rect 3966 11999 3972 12033
rect 4006 11999 4012 12033
rect 3966 11997 4012 11999
rect 3966 11931 3972 11997
rect 4006 11931 4012 11997
rect 3966 11925 4012 11931
rect 3966 11863 3972 11925
rect 4006 11863 4012 11925
rect 3966 11853 4012 11863
rect 3966 11795 3972 11853
rect 4006 11795 4012 11853
rect 3966 11781 4012 11795
rect 3966 11727 3972 11781
rect 4006 11727 4012 11781
rect 3966 11709 4012 11727
rect 3966 11659 3972 11709
rect 4006 11659 4012 11709
rect 3966 11637 4012 11659
rect 3966 11591 3972 11637
rect 4006 11591 4012 11637
rect 3966 11565 4012 11591
rect 3966 11523 3972 11565
rect 4006 11523 4012 11565
rect 3966 11493 4012 11523
rect 3966 11455 3972 11493
rect 4006 11455 4012 11493
rect 3966 11421 4012 11455
rect 3966 11387 3972 11421
rect 4006 11387 4012 11421
rect 3966 11353 4012 11387
rect 3966 11315 3972 11353
rect 4006 11315 4012 11353
rect 3966 11285 4012 11315
rect 3966 11243 3972 11285
rect 4006 11243 4012 11285
rect 3966 11217 4012 11243
rect 3966 11171 3972 11217
rect 4006 11171 4012 11217
rect 3966 11149 4012 11171
rect 3966 11099 3972 11149
rect 4006 11099 4012 11149
rect 3966 11081 4012 11099
rect 3966 11027 3972 11081
rect 4006 11027 4012 11081
rect 3966 11013 4012 11027
rect 3966 10955 3972 11013
rect 4006 10955 4012 11013
rect 3966 10945 4012 10955
rect 3966 10883 3972 10945
rect 4006 10883 4012 10945
rect 3966 10877 4012 10883
rect 3966 10811 3972 10877
rect 4006 10811 4012 10877
rect 3966 10809 4012 10811
rect 3966 10775 3972 10809
rect 4006 10775 4012 10809
rect 3966 10773 4012 10775
rect 3966 10707 3972 10773
rect 4006 10707 4012 10773
rect 3966 10701 4012 10707
rect 3966 10639 3972 10701
rect 4006 10639 4012 10701
rect 3966 10629 4012 10639
rect 3966 10571 3972 10629
rect 4006 10571 4012 10629
rect 3966 10557 4012 10571
rect 3966 10503 3972 10557
rect 4006 10503 4012 10557
rect 3966 10485 4012 10503
rect 3966 10435 3972 10485
rect 4006 10435 4012 10485
rect 3966 10413 4012 10435
rect 3966 10367 3972 10413
rect 4006 10367 4012 10413
rect 3966 10341 4012 10367
rect 3966 10299 3972 10341
rect 4006 10299 4012 10341
rect 3966 10269 4012 10299
rect 3966 10231 3972 10269
rect 4006 10231 4012 10269
rect 3966 10197 4012 10231
rect 3966 10163 3972 10197
rect 4006 10163 4012 10197
rect 3966 10129 4012 10163
rect 3966 10091 3972 10129
rect 4006 10091 4012 10129
rect 3966 10061 4012 10091
rect 3966 10019 3972 10061
rect 4006 10019 4012 10061
rect 3966 9993 4012 10019
rect 3966 9947 3972 9993
rect 4006 9947 4012 9993
rect 3966 9925 4012 9947
rect 3966 9875 3972 9925
rect 4006 9875 4012 9925
rect 3966 9857 4012 9875
rect 3966 9803 3972 9857
rect 4006 9803 4012 9857
rect 3966 9789 4012 9803
rect 3966 9731 3972 9789
rect 4006 9731 4012 9789
rect 3966 9721 4012 9731
rect 3966 9659 3972 9721
rect 4006 9659 4012 9721
rect 3966 9653 4012 9659
rect 3966 9587 3972 9653
rect 4006 9587 4012 9653
rect 3966 9585 4012 9587
rect 3966 9551 3972 9585
rect 4006 9551 4012 9585
rect 3966 9549 4012 9551
rect 3966 9483 3972 9549
rect 4006 9483 4012 9549
rect 3966 9477 4012 9483
rect 3966 9415 3972 9477
rect 4006 9415 4012 9477
rect 3966 9405 4012 9415
rect 3966 9347 3972 9405
rect 4006 9347 4012 9405
rect 3966 9333 4012 9347
rect 3966 9279 3972 9333
rect 4006 9279 4012 9333
rect 3966 9261 4012 9279
rect 3966 9211 3972 9261
rect 4006 9211 4012 9261
rect 3966 9189 4012 9211
rect 3966 9143 3972 9189
rect 4006 9143 4012 9189
rect 3966 9117 4012 9143
rect 3966 9075 3972 9117
rect 4006 9075 4012 9117
rect 3966 9045 4012 9075
rect 3966 9007 3972 9045
rect 4006 9007 4012 9045
rect 3966 8973 4012 9007
rect 3966 8939 3972 8973
rect 4006 8939 4012 8973
rect 3966 8905 4012 8939
rect 3966 8867 3972 8905
rect 4006 8867 4012 8905
rect 3966 8837 4012 8867
rect 3966 8795 3972 8837
rect 4006 8795 4012 8837
rect 3966 8769 4012 8795
rect 3966 8723 3972 8769
rect 4006 8723 4012 8769
rect 3966 8701 4012 8723
rect 3966 8651 3972 8701
rect 4006 8651 4012 8701
rect 3966 8633 4012 8651
rect 3966 8579 3972 8633
rect 4006 8579 4012 8633
rect 3966 8565 4012 8579
rect 3966 8507 3972 8565
rect 4006 8507 4012 8565
rect 3966 8497 4012 8507
rect 3966 8435 3972 8497
rect 4006 8435 4012 8497
rect 3966 8429 4012 8435
rect 3966 8363 3972 8429
rect 4006 8363 4012 8429
rect 3966 8361 4012 8363
rect 3966 8327 3972 8361
rect 4006 8327 4012 8361
rect 3966 8325 4012 8327
rect 3966 8259 3972 8325
rect 4006 8259 4012 8325
rect 3966 8253 4012 8259
rect 3966 8191 3972 8253
rect 4006 8191 4012 8253
rect 3966 8181 4012 8191
rect 3966 8123 3972 8181
rect 4006 8123 4012 8181
rect 3966 8109 4012 8123
rect 3966 8055 3972 8109
rect 4006 8055 4012 8109
rect 3966 8037 4012 8055
rect 3966 7987 3972 8037
rect 4006 7987 4012 8037
rect 3966 7965 4012 7987
rect 3966 7919 3972 7965
rect 4006 7919 4012 7965
rect 3966 7893 4012 7919
rect 3966 7851 3972 7893
rect 4006 7851 4012 7893
rect 3966 7821 4012 7851
rect 3966 7783 3972 7821
rect 4006 7783 4012 7821
rect 3966 7749 4012 7783
rect 3966 7715 3972 7749
rect 4006 7715 4012 7749
rect 3966 7681 4012 7715
rect 3966 7643 3972 7681
rect 4006 7643 4012 7681
rect 3966 7613 4012 7643
rect 3966 7571 3972 7613
rect 4006 7571 4012 7613
rect 3966 7545 4012 7571
rect 3966 7499 3972 7545
rect 4006 7499 4012 7545
rect 3966 7477 4012 7499
rect 3966 7427 3972 7477
rect 4006 7427 4012 7477
rect 3966 7409 4012 7427
rect 3966 7355 3972 7409
rect 4006 7355 4012 7409
rect 3966 7341 4012 7355
rect 3966 7283 3972 7341
rect 4006 7283 4012 7341
rect 3966 7273 4012 7283
rect 3966 7211 3972 7273
rect 4006 7211 4012 7273
rect 3966 7205 4012 7211
rect 3966 7139 3972 7205
rect 4006 7139 4012 7205
rect 3966 7137 4012 7139
rect 3966 7103 3972 7137
rect 4006 7103 4012 7137
rect 3966 7101 4012 7103
rect 3966 7035 3972 7101
rect 4006 7035 4012 7101
rect 3966 7029 4012 7035
rect 3966 6967 3972 7029
rect 4006 6967 4012 7029
rect 3966 6957 4012 6967
rect 3966 6899 3972 6957
rect 4006 6899 4012 6957
rect 3966 6885 4012 6899
rect 3966 6831 3972 6885
rect 4006 6831 4012 6885
rect 3966 6813 4012 6831
rect 3966 6763 3972 6813
rect 4006 6763 4012 6813
rect 3966 6741 4012 6763
rect 3966 6695 3972 6741
rect 4006 6695 4012 6741
rect 3966 6669 4012 6695
rect 3966 6627 3972 6669
rect 4006 6627 4012 6669
rect 3966 6597 4012 6627
rect 3966 6559 3972 6597
rect 4006 6559 4012 6597
rect 3966 6525 4012 6559
rect 3966 6491 3972 6525
rect 4006 6491 4012 6525
rect 3966 6457 4012 6491
rect 3966 6419 3972 6457
rect 4006 6419 4012 6457
rect 3966 6389 4012 6419
rect 3966 6347 3972 6389
rect 4006 6347 4012 6389
rect 3966 6321 4012 6347
rect 3966 6275 3972 6321
rect 4006 6275 4012 6321
rect 3966 6253 4012 6275
rect 3966 6203 3972 6253
rect 4006 6203 4012 6253
rect 3966 6185 4012 6203
rect 3966 6131 3972 6185
rect 4006 6131 4012 6185
rect 3966 6117 4012 6131
rect 3966 6059 3972 6117
rect 4006 6059 4012 6117
rect 3966 6049 4012 6059
rect 3966 5987 3972 6049
rect 4006 5987 4012 6049
rect 3966 5981 4012 5987
rect 3966 5915 3972 5981
rect 4006 5915 4012 5981
rect 3966 5913 4012 5915
rect 3966 5879 3972 5913
rect 4006 5879 4012 5913
rect 3966 5877 4012 5879
rect 3966 5811 3972 5877
rect 4006 5811 4012 5877
rect 3966 5805 4012 5811
rect 3966 5743 3972 5805
rect 4006 5743 4012 5805
rect 3966 5733 4012 5743
rect 3966 5675 3972 5733
rect 4006 5675 4012 5733
rect 3966 5661 4012 5675
rect 3966 5607 3972 5661
rect 4006 5607 4012 5661
rect 3966 5589 4012 5607
rect 3966 5539 3972 5589
rect 4006 5539 4012 5589
rect 3966 5517 4012 5539
rect 3966 5471 3972 5517
rect 4006 5471 4012 5517
rect 3966 5445 4012 5471
rect 3966 5403 3972 5445
rect 4006 5403 4012 5445
rect 3966 5373 4012 5403
rect 3966 5335 3972 5373
rect 4006 5335 4012 5373
rect 3966 5301 4012 5335
rect 3966 5267 3972 5301
rect 4006 5267 4012 5301
rect 3966 5233 4012 5267
rect 3966 5195 3972 5233
rect 4006 5195 4012 5233
rect 3966 5165 4012 5195
rect 3966 5123 3972 5165
rect 4006 5123 4012 5165
rect 3966 5097 4012 5123
rect 3966 5051 3972 5097
rect 4006 5051 4012 5097
rect 3966 5029 4012 5051
rect 3966 4979 3972 5029
rect 4006 4979 4012 5029
rect 3966 4961 4012 4979
rect 3966 4907 3972 4961
rect 4006 4907 4012 4961
rect 3966 4893 4012 4907
rect 3966 4835 3972 4893
rect 4006 4835 4012 4893
rect 3966 4825 4012 4835
rect 3966 4763 3972 4825
rect 4006 4763 4012 4825
rect 3966 4757 4012 4763
rect 3966 4691 3972 4757
rect 4006 4691 4012 4757
rect 3966 4689 4012 4691
rect 3966 4655 3972 4689
rect 4006 4655 4012 4689
rect 3966 4653 4012 4655
rect 3966 4587 3972 4653
rect 4006 4587 4012 4653
rect 3966 4581 4012 4587
rect 3966 4519 3972 4581
rect 4006 4519 4012 4581
rect 3966 4509 4012 4519
rect 3966 4451 3972 4509
rect 4006 4451 4012 4509
rect 3966 4437 4012 4451
rect 3966 4383 3972 4437
rect 4006 4383 4012 4437
rect 3966 4365 4012 4383
rect 3966 4315 3972 4365
rect 4006 4315 4012 4365
rect 3966 4293 4012 4315
rect 3966 4247 3972 4293
rect 4006 4247 4012 4293
rect 3966 4221 4012 4247
rect 3966 4179 3972 4221
rect 4006 4179 4012 4221
rect 3966 4149 4012 4179
rect 3966 4111 3972 4149
rect 4006 4111 4012 4149
rect 3966 4077 4012 4111
rect 3966 4043 3972 4077
rect 4006 4043 4012 4077
rect 3966 4009 4012 4043
rect 3966 3971 3972 4009
rect 4006 3971 4012 4009
rect 3966 3941 4012 3971
rect 3966 3899 3972 3941
rect 4006 3899 4012 3941
rect 3966 3873 4012 3899
rect 3966 3827 3972 3873
rect 4006 3827 4012 3873
rect 3966 3805 4012 3827
rect 3966 3755 3972 3805
rect 4006 3755 4012 3805
rect 3966 3737 4012 3755
rect 3966 3683 3972 3737
rect 4006 3683 4012 3737
rect 3966 3669 4012 3683
rect 3966 3611 3972 3669
rect 4006 3611 4012 3669
rect 3966 3601 4012 3611
rect 3966 3539 3972 3601
rect 4006 3539 4012 3601
rect 3966 3533 4012 3539
rect 1824 3429 1870 3451
rect 1824 3383 1830 3429
rect 1864 3383 1870 3429
rect -258 3295 -252 3357
rect -218 3295 -212 3357
rect -258 3285 -212 3295
rect -258 3251 -252 3285
rect -218 3251 -212 3285
rect -258 3219 -212 3251
rect 1824 3357 1870 3383
rect 2000 3452 2016 3472
rect 2050 3452 2066 3472
rect 2000 3414 2066 3452
rect 2000 3360 2016 3414
rect 2050 3360 2066 3414
rect 2118 3452 2134 3472
rect 2168 3452 2184 3472
rect 2118 3414 2184 3452
rect 2118 3360 2134 3414
rect 2168 3360 2184 3414
rect 2236 3452 2252 3472
rect 2286 3452 2302 3472
rect 2236 3414 2302 3452
rect 2236 3360 2252 3414
rect 2286 3360 2302 3414
rect 2354 3452 2370 3472
rect 2404 3452 2420 3472
rect 2354 3414 2420 3452
rect 2354 3360 2370 3414
rect 2404 3360 2420 3414
rect 2472 3452 2488 3472
rect 2522 3452 2538 3472
rect 2472 3414 2538 3452
rect 2472 3360 2488 3414
rect 2522 3360 2538 3414
rect 2590 3452 2606 3472
rect 2640 3452 2656 3472
rect 2590 3414 2656 3452
rect 2590 3360 2606 3414
rect 2640 3360 2656 3414
rect 2708 3452 2724 3472
rect 2758 3452 2774 3472
rect 2708 3414 2774 3452
rect 2708 3360 2724 3414
rect 2758 3360 2774 3414
rect 2826 3452 2842 3472
rect 2876 3452 2892 3472
rect 2826 3414 2892 3452
rect 2826 3360 2842 3414
rect 2876 3360 2892 3414
rect 2944 3452 2960 3472
rect 2994 3452 3010 3472
rect 2944 3414 3010 3452
rect 2944 3360 2960 3414
rect 2994 3360 3010 3414
rect 3062 3452 3078 3472
rect 3112 3452 3128 3472
rect 3062 3414 3128 3452
rect 3062 3360 3078 3414
rect 3112 3360 3128 3414
rect 3180 3452 3196 3472
rect 3230 3452 3246 3472
rect 3180 3414 3246 3452
rect 3180 3360 3196 3414
rect 3230 3360 3246 3414
rect 3298 3452 3314 3472
rect 3348 3452 3364 3472
rect 3298 3414 3364 3452
rect 3298 3360 3314 3414
rect 3348 3360 3364 3414
rect 3416 3452 3432 3472
rect 3466 3452 3482 3472
rect 3416 3414 3482 3452
rect 3416 3360 3432 3414
rect 3466 3360 3482 3414
rect 3534 3452 3550 3472
rect 3584 3452 3600 3472
rect 3534 3414 3600 3452
rect 3534 3360 3550 3414
rect 3584 3360 3600 3414
rect 3652 3452 3668 3472
rect 3702 3452 3718 3472
rect 3652 3414 3718 3452
rect 3652 3360 3668 3414
rect 3702 3360 3718 3414
rect 3770 3452 3786 3472
rect 3820 3452 3836 3472
rect 3770 3414 3836 3452
rect 3770 3360 3786 3414
rect 3820 3360 3836 3414
rect 3966 3467 3972 3533
rect 4006 3467 4012 3533
rect 6108 38685 6154 38717
rect 6108 38651 6114 38685
rect 6148 38651 6154 38685
rect 6108 38641 6154 38651
rect 6108 38579 6114 38641
rect 6148 38579 6154 38641
rect 6108 38573 6154 38579
rect 6108 38507 6114 38573
rect 6148 38507 6154 38573
rect 6108 38505 6154 38507
rect 6108 38471 6114 38505
rect 6148 38471 6154 38505
rect 6108 38469 6154 38471
rect 6108 38403 6114 38469
rect 6148 38403 6154 38469
rect 6108 38397 6154 38403
rect 6108 38335 6114 38397
rect 6148 38335 6154 38397
rect 6108 38325 6154 38335
rect 6108 38267 6114 38325
rect 6148 38267 6154 38325
rect 6108 38253 6154 38267
rect 6108 38199 6114 38253
rect 6148 38199 6154 38253
rect 6108 38181 6154 38199
rect 6108 38131 6114 38181
rect 6148 38131 6154 38181
rect 6108 38109 6154 38131
rect 6108 38063 6114 38109
rect 6148 38063 6154 38109
rect 6108 38037 6154 38063
rect 6108 37995 6114 38037
rect 6148 37995 6154 38037
rect 6108 37965 6154 37995
rect 6108 37927 6114 37965
rect 6148 37927 6154 37965
rect 6108 37893 6154 37927
rect 6108 37859 6114 37893
rect 6148 37859 6154 37893
rect 6108 37825 6154 37859
rect 6108 37787 6114 37825
rect 6148 37787 6154 37825
rect 6108 37757 6154 37787
rect 6108 37715 6114 37757
rect 6148 37715 6154 37757
rect 6108 37689 6154 37715
rect 6108 37643 6114 37689
rect 6148 37643 6154 37689
rect 6108 37621 6154 37643
rect 6108 37571 6114 37621
rect 6148 37571 6154 37621
rect 6108 37553 6154 37571
rect 6108 37499 6114 37553
rect 6148 37499 6154 37553
rect 6108 37485 6154 37499
rect 6108 37427 6114 37485
rect 6148 37427 6154 37485
rect 6108 37417 6154 37427
rect 6108 37355 6114 37417
rect 6148 37355 6154 37417
rect 6108 37349 6154 37355
rect 6108 37283 6114 37349
rect 6148 37283 6154 37349
rect 6108 37281 6154 37283
rect 6108 37247 6114 37281
rect 6148 37247 6154 37281
rect 6108 37245 6154 37247
rect 6108 37179 6114 37245
rect 6148 37179 6154 37245
rect 6108 37173 6154 37179
rect 6108 37111 6114 37173
rect 6148 37111 6154 37173
rect 6108 37101 6154 37111
rect 6108 37043 6114 37101
rect 6148 37043 6154 37101
rect 6108 37029 6154 37043
rect 6108 36975 6114 37029
rect 6148 36975 6154 37029
rect 6108 36957 6154 36975
rect 6108 36907 6114 36957
rect 6148 36907 6154 36957
rect 6108 36885 6154 36907
rect 6108 36839 6114 36885
rect 6148 36839 6154 36885
rect 6108 36813 6154 36839
rect 6108 36771 6114 36813
rect 6148 36771 6154 36813
rect 6108 36741 6154 36771
rect 6108 36703 6114 36741
rect 6148 36703 6154 36741
rect 6108 36669 6154 36703
rect 6108 36635 6114 36669
rect 6148 36635 6154 36669
rect 6108 36601 6154 36635
rect 6108 36563 6114 36601
rect 6148 36563 6154 36601
rect 6108 36533 6154 36563
rect 6108 36491 6114 36533
rect 6148 36491 6154 36533
rect 6108 36465 6154 36491
rect 6108 36419 6114 36465
rect 6148 36419 6154 36465
rect 6108 36397 6154 36419
rect 6108 36347 6114 36397
rect 6148 36347 6154 36397
rect 6108 36329 6154 36347
rect 6108 36275 6114 36329
rect 6148 36275 6154 36329
rect 6108 36261 6154 36275
rect 6108 36203 6114 36261
rect 6148 36203 6154 36261
rect 6108 36193 6154 36203
rect 6108 36131 6114 36193
rect 6148 36131 6154 36193
rect 6108 36125 6154 36131
rect 6108 36059 6114 36125
rect 6148 36059 6154 36125
rect 6108 36057 6154 36059
rect 6108 36023 6114 36057
rect 6148 36023 6154 36057
rect 6108 36021 6154 36023
rect 6108 35955 6114 36021
rect 6148 35955 6154 36021
rect 6108 35949 6154 35955
rect 6108 35887 6114 35949
rect 6148 35887 6154 35949
rect 6108 35877 6154 35887
rect 6108 35819 6114 35877
rect 6148 35819 6154 35877
rect 6108 35805 6154 35819
rect 6108 35751 6114 35805
rect 6148 35751 6154 35805
rect 6108 35733 6154 35751
rect 6108 35683 6114 35733
rect 6148 35683 6154 35733
rect 6108 35661 6154 35683
rect 6108 35615 6114 35661
rect 6148 35615 6154 35661
rect 6108 35589 6154 35615
rect 6108 35547 6114 35589
rect 6148 35547 6154 35589
rect 6108 35517 6154 35547
rect 6108 35479 6114 35517
rect 6148 35479 6154 35517
rect 6108 35445 6154 35479
rect 6108 35411 6114 35445
rect 6148 35411 6154 35445
rect 6108 35377 6154 35411
rect 6108 35339 6114 35377
rect 6148 35339 6154 35377
rect 6108 35309 6154 35339
rect 6108 35267 6114 35309
rect 6148 35267 6154 35309
rect 6108 35241 6154 35267
rect 6108 35195 6114 35241
rect 6148 35195 6154 35241
rect 6108 35173 6154 35195
rect 6108 35123 6114 35173
rect 6148 35123 6154 35173
rect 6108 35105 6154 35123
rect 6108 35051 6114 35105
rect 6148 35051 6154 35105
rect 6108 35037 6154 35051
rect 6108 34979 6114 35037
rect 6148 34979 6154 35037
rect 6108 34969 6154 34979
rect 6108 34907 6114 34969
rect 6148 34907 6154 34969
rect 6108 34901 6154 34907
rect 6108 34835 6114 34901
rect 6148 34835 6154 34901
rect 6108 34833 6154 34835
rect 6108 34799 6114 34833
rect 6148 34799 6154 34833
rect 6108 34797 6154 34799
rect 6108 34731 6114 34797
rect 6148 34731 6154 34797
rect 6108 34725 6154 34731
rect 6108 34663 6114 34725
rect 6148 34663 6154 34725
rect 6108 34653 6154 34663
rect 6108 34595 6114 34653
rect 6148 34595 6154 34653
rect 6108 34581 6154 34595
rect 6108 34527 6114 34581
rect 6148 34527 6154 34581
rect 6108 34509 6154 34527
rect 6108 34459 6114 34509
rect 6148 34459 6154 34509
rect 6108 34437 6154 34459
rect 6108 34391 6114 34437
rect 6148 34391 6154 34437
rect 6108 34365 6154 34391
rect 6108 34323 6114 34365
rect 6148 34323 6154 34365
rect 6108 34293 6154 34323
rect 6108 34255 6114 34293
rect 6148 34255 6154 34293
rect 6108 34221 6154 34255
rect 6108 34187 6114 34221
rect 6148 34187 6154 34221
rect 6108 34153 6154 34187
rect 6108 34115 6114 34153
rect 6148 34115 6154 34153
rect 6108 34085 6154 34115
rect 6108 34043 6114 34085
rect 6148 34043 6154 34085
rect 6108 34017 6154 34043
rect 6108 33971 6114 34017
rect 6148 33971 6154 34017
rect 6108 33949 6154 33971
rect 6108 33899 6114 33949
rect 6148 33899 6154 33949
rect 6108 33881 6154 33899
rect 6108 33827 6114 33881
rect 6148 33827 6154 33881
rect 6108 33813 6154 33827
rect 6108 33755 6114 33813
rect 6148 33755 6154 33813
rect 6108 33745 6154 33755
rect 6108 33683 6114 33745
rect 6148 33683 6154 33745
rect 6108 33677 6154 33683
rect 6108 33611 6114 33677
rect 6148 33611 6154 33677
rect 6108 33609 6154 33611
rect 6108 33575 6114 33609
rect 6148 33575 6154 33609
rect 6108 33573 6154 33575
rect 6108 33507 6114 33573
rect 6148 33507 6154 33573
rect 6108 33501 6154 33507
rect 6108 33439 6114 33501
rect 6148 33439 6154 33501
rect 6108 33429 6154 33439
rect 6108 33371 6114 33429
rect 6148 33371 6154 33429
rect 6108 33357 6154 33371
rect 6108 33303 6114 33357
rect 6148 33303 6154 33357
rect 6108 33285 6154 33303
rect 6108 33235 6114 33285
rect 6148 33235 6154 33285
rect 6108 33213 6154 33235
rect 6108 33167 6114 33213
rect 6148 33167 6154 33213
rect 6108 33141 6154 33167
rect 6108 33099 6114 33141
rect 6148 33099 6154 33141
rect 6108 33069 6154 33099
rect 6108 33031 6114 33069
rect 6148 33031 6154 33069
rect 6108 32997 6154 33031
rect 6108 32963 6114 32997
rect 6148 32963 6154 32997
rect 6108 32929 6154 32963
rect 6108 32891 6114 32929
rect 6148 32891 6154 32929
rect 6108 32861 6154 32891
rect 6108 32819 6114 32861
rect 6148 32819 6154 32861
rect 6108 32793 6154 32819
rect 6108 32747 6114 32793
rect 6148 32747 6154 32793
rect 6108 32725 6154 32747
rect 6108 32675 6114 32725
rect 6148 32675 6154 32725
rect 6108 32657 6154 32675
rect 6108 32603 6114 32657
rect 6148 32603 6154 32657
rect 6108 32589 6154 32603
rect 6108 32531 6114 32589
rect 6148 32531 6154 32589
rect 6108 32521 6154 32531
rect 6108 32459 6114 32521
rect 6148 32459 6154 32521
rect 6108 32453 6154 32459
rect 6108 32387 6114 32453
rect 6148 32387 6154 32453
rect 6108 32385 6154 32387
rect 6108 32351 6114 32385
rect 6148 32351 6154 32385
rect 6108 32349 6154 32351
rect 6108 32283 6114 32349
rect 6148 32283 6154 32349
rect 6108 32277 6154 32283
rect 6108 32215 6114 32277
rect 6148 32215 6154 32277
rect 6108 32205 6154 32215
rect 6108 32147 6114 32205
rect 6148 32147 6154 32205
rect 6108 32133 6154 32147
rect 6108 32079 6114 32133
rect 6148 32079 6154 32133
rect 6108 32061 6154 32079
rect 6108 32011 6114 32061
rect 6148 32011 6154 32061
rect 6108 31989 6154 32011
rect 6108 31943 6114 31989
rect 6148 31943 6154 31989
rect 6108 31917 6154 31943
rect 6108 31875 6114 31917
rect 6148 31875 6154 31917
rect 6108 31845 6154 31875
rect 6108 31807 6114 31845
rect 6148 31807 6154 31845
rect 6108 31773 6154 31807
rect 6108 31739 6114 31773
rect 6148 31739 6154 31773
rect 6108 31705 6154 31739
rect 6108 31667 6114 31705
rect 6148 31667 6154 31705
rect 6108 31637 6154 31667
rect 6108 31595 6114 31637
rect 6148 31595 6154 31637
rect 6108 31569 6154 31595
rect 6108 31523 6114 31569
rect 6148 31523 6154 31569
rect 6108 31501 6154 31523
rect 6108 31451 6114 31501
rect 6148 31451 6154 31501
rect 6108 31433 6154 31451
rect 6108 31379 6114 31433
rect 6148 31379 6154 31433
rect 6108 31365 6154 31379
rect 6108 31307 6114 31365
rect 6148 31307 6154 31365
rect 6108 31297 6154 31307
rect 6108 31235 6114 31297
rect 6148 31235 6154 31297
rect 6108 31229 6154 31235
rect 6108 31163 6114 31229
rect 6148 31163 6154 31229
rect 6108 31161 6154 31163
rect 6108 31127 6114 31161
rect 6148 31127 6154 31161
rect 6108 31125 6154 31127
rect 6108 31059 6114 31125
rect 6148 31059 6154 31125
rect 6108 31053 6154 31059
rect 6108 30991 6114 31053
rect 6148 30991 6154 31053
rect 6108 30981 6154 30991
rect 6108 30923 6114 30981
rect 6148 30923 6154 30981
rect 6108 30909 6154 30923
rect 6108 30855 6114 30909
rect 6148 30855 6154 30909
rect 6108 30837 6154 30855
rect 6108 30787 6114 30837
rect 6148 30787 6154 30837
rect 6108 30765 6154 30787
rect 6108 30719 6114 30765
rect 6148 30719 6154 30765
rect 6108 30693 6154 30719
rect 6108 30651 6114 30693
rect 6148 30651 6154 30693
rect 6108 30621 6154 30651
rect 6108 30583 6114 30621
rect 6148 30583 6154 30621
rect 6108 30549 6154 30583
rect 6108 30515 6114 30549
rect 6148 30515 6154 30549
rect 6108 30481 6154 30515
rect 6108 30443 6114 30481
rect 6148 30443 6154 30481
rect 6108 30413 6154 30443
rect 6108 30371 6114 30413
rect 6148 30371 6154 30413
rect 6108 30345 6154 30371
rect 6108 30299 6114 30345
rect 6148 30299 6154 30345
rect 6108 30277 6154 30299
rect 6108 30227 6114 30277
rect 6148 30227 6154 30277
rect 6108 30209 6154 30227
rect 6108 30155 6114 30209
rect 6148 30155 6154 30209
rect 6108 30141 6154 30155
rect 6108 30083 6114 30141
rect 6148 30083 6154 30141
rect 6108 30073 6154 30083
rect 6108 30011 6114 30073
rect 6148 30011 6154 30073
rect 6108 30005 6154 30011
rect 6108 29939 6114 30005
rect 6148 29939 6154 30005
rect 6108 29937 6154 29939
rect 6108 29903 6114 29937
rect 6148 29903 6154 29937
rect 6108 29901 6154 29903
rect 6108 29835 6114 29901
rect 6148 29835 6154 29901
rect 6108 29829 6154 29835
rect 6108 29767 6114 29829
rect 6148 29767 6154 29829
rect 6108 29757 6154 29767
rect 6108 29699 6114 29757
rect 6148 29699 6154 29757
rect 6108 29685 6154 29699
rect 6108 29631 6114 29685
rect 6148 29631 6154 29685
rect 6108 29613 6154 29631
rect 6108 29563 6114 29613
rect 6148 29563 6154 29613
rect 6108 29541 6154 29563
rect 6108 29495 6114 29541
rect 6148 29495 6154 29541
rect 6108 29469 6154 29495
rect 6108 29427 6114 29469
rect 6148 29427 6154 29469
rect 6108 29397 6154 29427
rect 6108 29359 6114 29397
rect 6148 29359 6154 29397
rect 6108 29325 6154 29359
rect 6108 29291 6114 29325
rect 6148 29291 6154 29325
rect 6108 29257 6154 29291
rect 6108 29219 6114 29257
rect 6148 29219 6154 29257
rect 6108 29189 6154 29219
rect 6108 29147 6114 29189
rect 6148 29147 6154 29189
rect 6108 29121 6154 29147
rect 6108 29075 6114 29121
rect 6148 29075 6154 29121
rect 6108 29053 6154 29075
rect 6108 29003 6114 29053
rect 6148 29003 6154 29053
rect 6108 28985 6154 29003
rect 6108 28931 6114 28985
rect 6148 28931 6154 28985
rect 6108 28917 6154 28931
rect 6108 28859 6114 28917
rect 6148 28859 6154 28917
rect 6108 28849 6154 28859
rect 6108 28787 6114 28849
rect 6148 28787 6154 28849
rect 6108 28781 6154 28787
rect 6108 28715 6114 28781
rect 6148 28715 6154 28781
rect 6108 28713 6154 28715
rect 6108 28679 6114 28713
rect 6148 28679 6154 28713
rect 6108 28677 6154 28679
rect 6108 28611 6114 28677
rect 6148 28611 6154 28677
rect 6108 28605 6154 28611
rect 6108 28543 6114 28605
rect 6148 28543 6154 28605
rect 6108 28533 6154 28543
rect 6108 28475 6114 28533
rect 6148 28475 6154 28533
rect 6108 28461 6154 28475
rect 6108 28407 6114 28461
rect 6148 28407 6154 28461
rect 6108 28389 6154 28407
rect 6108 28339 6114 28389
rect 6148 28339 6154 28389
rect 6108 28317 6154 28339
rect 6108 28271 6114 28317
rect 6148 28271 6154 28317
rect 6108 28245 6154 28271
rect 6108 28203 6114 28245
rect 6148 28203 6154 28245
rect 6108 28173 6154 28203
rect 6108 28135 6114 28173
rect 6148 28135 6154 28173
rect 6108 28101 6154 28135
rect 6108 28067 6114 28101
rect 6148 28067 6154 28101
rect 6108 28033 6154 28067
rect 6108 27995 6114 28033
rect 6148 27995 6154 28033
rect 6108 27965 6154 27995
rect 6108 27923 6114 27965
rect 6148 27923 6154 27965
rect 6108 27897 6154 27923
rect 6108 27851 6114 27897
rect 6148 27851 6154 27897
rect 6108 27829 6154 27851
rect 6108 27779 6114 27829
rect 6148 27779 6154 27829
rect 6108 27761 6154 27779
rect 6108 27707 6114 27761
rect 6148 27707 6154 27761
rect 6108 27693 6154 27707
rect 6108 27635 6114 27693
rect 6148 27635 6154 27693
rect 6108 27625 6154 27635
rect 6108 27563 6114 27625
rect 6148 27563 6154 27625
rect 6108 27557 6154 27563
rect 6108 27491 6114 27557
rect 6148 27491 6154 27557
rect 6108 27489 6154 27491
rect 6108 27455 6114 27489
rect 6148 27455 6154 27489
rect 6108 27453 6154 27455
rect 6108 27387 6114 27453
rect 6148 27387 6154 27453
rect 6108 27381 6154 27387
rect 6108 27319 6114 27381
rect 6148 27319 6154 27381
rect 6108 27309 6154 27319
rect 6108 27251 6114 27309
rect 6148 27251 6154 27309
rect 6108 27237 6154 27251
rect 6108 27183 6114 27237
rect 6148 27183 6154 27237
rect 6108 27165 6154 27183
rect 6108 27115 6114 27165
rect 6148 27115 6154 27165
rect 6108 27093 6154 27115
rect 6108 27047 6114 27093
rect 6148 27047 6154 27093
rect 6108 27021 6154 27047
rect 6108 26979 6114 27021
rect 6148 26979 6154 27021
rect 6108 26949 6154 26979
rect 6108 26911 6114 26949
rect 6148 26911 6154 26949
rect 6108 26877 6154 26911
rect 6108 26843 6114 26877
rect 6148 26843 6154 26877
rect 6108 26809 6154 26843
rect 6108 26771 6114 26809
rect 6148 26771 6154 26809
rect 6108 26741 6154 26771
rect 6108 26699 6114 26741
rect 6148 26699 6154 26741
rect 6108 26673 6154 26699
rect 6108 26627 6114 26673
rect 6148 26627 6154 26673
rect 6108 26605 6154 26627
rect 6108 26555 6114 26605
rect 6148 26555 6154 26605
rect 6108 26537 6154 26555
rect 6108 26483 6114 26537
rect 6148 26483 6154 26537
rect 6108 26469 6154 26483
rect 6108 26411 6114 26469
rect 6148 26411 6154 26469
rect 6108 26401 6154 26411
rect 6108 26339 6114 26401
rect 6148 26339 6154 26401
rect 6108 26333 6154 26339
rect 6108 26267 6114 26333
rect 6148 26267 6154 26333
rect 6108 26265 6154 26267
rect 6108 26231 6114 26265
rect 6148 26231 6154 26265
rect 6108 26229 6154 26231
rect 6108 26163 6114 26229
rect 6148 26163 6154 26229
rect 6108 26157 6154 26163
rect 6108 26095 6114 26157
rect 6148 26095 6154 26157
rect 6108 26085 6154 26095
rect 6108 26027 6114 26085
rect 6148 26027 6154 26085
rect 6108 26013 6154 26027
rect 6108 25959 6114 26013
rect 6148 25959 6154 26013
rect 6108 25941 6154 25959
rect 6108 25891 6114 25941
rect 6148 25891 6154 25941
rect 6108 25869 6154 25891
rect 6108 25823 6114 25869
rect 6148 25823 6154 25869
rect 6108 25797 6154 25823
rect 6108 25755 6114 25797
rect 6148 25755 6154 25797
rect 6108 25725 6154 25755
rect 6108 25687 6114 25725
rect 6148 25687 6154 25725
rect 6108 25653 6154 25687
rect 6108 25619 6114 25653
rect 6148 25619 6154 25653
rect 6108 25585 6154 25619
rect 6108 25547 6114 25585
rect 6148 25547 6154 25585
rect 6108 25517 6154 25547
rect 6108 25475 6114 25517
rect 6148 25475 6154 25517
rect 6108 25449 6154 25475
rect 6108 25403 6114 25449
rect 6148 25403 6154 25449
rect 6108 25381 6154 25403
rect 6108 25331 6114 25381
rect 6148 25331 6154 25381
rect 6108 25313 6154 25331
rect 6108 25259 6114 25313
rect 6148 25259 6154 25313
rect 6108 25245 6154 25259
rect 6108 25187 6114 25245
rect 6148 25187 6154 25245
rect 6108 25177 6154 25187
rect 6108 25115 6114 25177
rect 6148 25115 6154 25177
rect 6108 25109 6154 25115
rect 6108 25043 6114 25109
rect 6148 25043 6154 25109
rect 6108 25041 6154 25043
rect 6108 25007 6114 25041
rect 6148 25007 6154 25041
rect 6108 25005 6154 25007
rect 6108 24939 6114 25005
rect 6148 24939 6154 25005
rect 6108 24933 6154 24939
rect 6108 24871 6114 24933
rect 6148 24871 6154 24933
rect 6108 24861 6154 24871
rect 6108 24803 6114 24861
rect 6148 24803 6154 24861
rect 6108 24789 6154 24803
rect 6108 24735 6114 24789
rect 6148 24735 6154 24789
rect 6108 24717 6154 24735
rect 6108 24667 6114 24717
rect 6148 24667 6154 24717
rect 6108 24645 6154 24667
rect 6108 24599 6114 24645
rect 6148 24599 6154 24645
rect 6108 24573 6154 24599
rect 6108 24531 6114 24573
rect 6148 24531 6154 24573
rect 6108 24501 6154 24531
rect 6108 24463 6114 24501
rect 6148 24463 6154 24501
rect 6108 24429 6154 24463
rect 6108 24395 6114 24429
rect 6148 24395 6154 24429
rect 6108 24361 6154 24395
rect 6108 24323 6114 24361
rect 6148 24323 6154 24361
rect 6108 24293 6154 24323
rect 6108 24251 6114 24293
rect 6148 24251 6154 24293
rect 6108 24225 6154 24251
rect 6108 24179 6114 24225
rect 6148 24179 6154 24225
rect 6108 24157 6154 24179
rect 6108 24107 6114 24157
rect 6148 24107 6154 24157
rect 6108 24089 6154 24107
rect 6108 24035 6114 24089
rect 6148 24035 6154 24089
rect 6108 24021 6154 24035
rect 6108 23963 6114 24021
rect 6148 23963 6154 24021
rect 6108 23953 6154 23963
rect 6108 23891 6114 23953
rect 6148 23891 6154 23953
rect 6108 23885 6154 23891
rect 6108 23819 6114 23885
rect 6148 23819 6154 23885
rect 6108 23817 6154 23819
rect 6108 23783 6114 23817
rect 6148 23783 6154 23817
rect 6108 23781 6154 23783
rect 6108 23715 6114 23781
rect 6148 23715 6154 23781
rect 6108 23709 6154 23715
rect 6108 23647 6114 23709
rect 6148 23647 6154 23709
rect 6108 23637 6154 23647
rect 6108 23579 6114 23637
rect 6148 23579 6154 23637
rect 6108 23565 6154 23579
rect 6108 23511 6114 23565
rect 6148 23511 6154 23565
rect 6108 23493 6154 23511
rect 6108 23443 6114 23493
rect 6148 23443 6154 23493
rect 6108 23421 6154 23443
rect 6108 23375 6114 23421
rect 6148 23375 6154 23421
rect 6108 23349 6154 23375
rect 6108 23307 6114 23349
rect 6148 23307 6154 23349
rect 6108 23277 6154 23307
rect 6108 23239 6114 23277
rect 6148 23239 6154 23277
rect 6108 23205 6154 23239
rect 6108 23171 6114 23205
rect 6148 23171 6154 23205
rect 6108 23137 6154 23171
rect 6108 23099 6114 23137
rect 6148 23099 6154 23137
rect 6108 23069 6154 23099
rect 6108 23027 6114 23069
rect 6148 23027 6154 23069
rect 6108 23001 6154 23027
rect 6108 22955 6114 23001
rect 6148 22955 6154 23001
rect 6108 22933 6154 22955
rect 6108 22883 6114 22933
rect 6148 22883 6154 22933
rect 6108 22865 6154 22883
rect 6108 22811 6114 22865
rect 6148 22811 6154 22865
rect 6108 22797 6154 22811
rect 6108 22739 6114 22797
rect 6148 22739 6154 22797
rect 6108 22729 6154 22739
rect 6108 22667 6114 22729
rect 6148 22667 6154 22729
rect 6108 22661 6154 22667
rect 6108 22595 6114 22661
rect 6148 22595 6154 22661
rect 6108 22593 6154 22595
rect 6108 22559 6114 22593
rect 6148 22559 6154 22593
rect 6108 22557 6154 22559
rect 6108 22491 6114 22557
rect 6148 22491 6154 22557
rect 6108 22485 6154 22491
rect 6108 22423 6114 22485
rect 6148 22423 6154 22485
rect 6108 22413 6154 22423
rect 6108 22355 6114 22413
rect 6148 22355 6154 22413
rect 6108 22341 6154 22355
rect 6108 22287 6114 22341
rect 6148 22287 6154 22341
rect 6108 22269 6154 22287
rect 6108 22219 6114 22269
rect 6148 22219 6154 22269
rect 6108 22197 6154 22219
rect 6108 22151 6114 22197
rect 6148 22151 6154 22197
rect 6108 22125 6154 22151
rect 6108 22083 6114 22125
rect 6148 22083 6154 22125
rect 6108 22053 6154 22083
rect 6108 22015 6114 22053
rect 6148 22015 6154 22053
rect 6108 21981 6154 22015
rect 6108 21947 6114 21981
rect 6148 21947 6154 21981
rect 6108 21913 6154 21947
rect 6108 21875 6114 21913
rect 6148 21875 6154 21913
rect 6108 21845 6154 21875
rect 6108 21803 6114 21845
rect 6148 21803 6154 21845
rect 6108 21777 6154 21803
rect 6108 21731 6114 21777
rect 6148 21731 6154 21777
rect 6108 21709 6154 21731
rect 6108 21659 6114 21709
rect 6148 21659 6154 21709
rect 6108 21641 6154 21659
rect 6108 21587 6114 21641
rect 6148 21587 6154 21641
rect 6108 21573 6154 21587
rect 6108 21515 6114 21573
rect 6148 21515 6154 21573
rect 6108 21505 6154 21515
rect 6108 21443 6114 21505
rect 6148 21443 6154 21505
rect 6108 21437 6154 21443
rect 6108 21371 6114 21437
rect 6148 21371 6154 21437
rect 6108 21369 6154 21371
rect 6108 21335 6114 21369
rect 6148 21335 6154 21369
rect 6108 21333 6154 21335
rect 6108 21267 6114 21333
rect 6148 21267 6154 21333
rect 6108 21261 6154 21267
rect 6108 21199 6114 21261
rect 6148 21199 6154 21261
rect 6108 21189 6154 21199
rect 6108 21131 6114 21189
rect 6148 21131 6154 21189
rect 6108 21117 6154 21131
rect 6108 21063 6114 21117
rect 6148 21063 6154 21117
rect 6108 21045 6154 21063
rect 6108 20995 6114 21045
rect 6148 20995 6154 21045
rect 6108 20973 6154 20995
rect 6108 20927 6114 20973
rect 6148 20927 6154 20973
rect 6108 20901 6154 20927
rect 6108 20859 6114 20901
rect 6148 20859 6154 20901
rect 6108 20829 6154 20859
rect 6108 20791 6114 20829
rect 6148 20791 6154 20829
rect 6108 20757 6154 20791
rect 6108 20723 6114 20757
rect 6148 20723 6154 20757
rect 6108 20689 6154 20723
rect 6108 20651 6114 20689
rect 6148 20651 6154 20689
rect 6108 20621 6154 20651
rect 6108 20579 6114 20621
rect 6148 20579 6154 20621
rect 6108 20553 6154 20579
rect 6108 20507 6114 20553
rect 6148 20507 6154 20553
rect 6108 20485 6154 20507
rect 6108 20435 6114 20485
rect 6148 20435 6154 20485
rect 6108 20417 6154 20435
rect 6108 20363 6114 20417
rect 6148 20363 6154 20417
rect 6108 20349 6154 20363
rect 6108 20291 6114 20349
rect 6148 20291 6154 20349
rect 6108 20281 6154 20291
rect 6108 20219 6114 20281
rect 6148 20219 6154 20281
rect 6108 20213 6154 20219
rect 6108 20147 6114 20213
rect 6148 20147 6154 20213
rect 6108 20145 6154 20147
rect 6108 20111 6114 20145
rect 6148 20111 6154 20145
rect 6108 20109 6154 20111
rect 6108 20043 6114 20109
rect 6148 20043 6154 20109
rect 6108 20037 6154 20043
rect 6108 19975 6114 20037
rect 6148 19975 6154 20037
rect 6108 19965 6154 19975
rect 6108 19907 6114 19965
rect 6148 19907 6154 19965
rect 6108 19893 6154 19907
rect 6108 19839 6114 19893
rect 6148 19839 6154 19893
rect 6108 19821 6154 19839
rect 6108 19771 6114 19821
rect 6148 19771 6154 19821
rect 6108 19749 6154 19771
rect 6108 19703 6114 19749
rect 6148 19703 6154 19749
rect 6108 19677 6154 19703
rect 6108 19635 6114 19677
rect 6148 19635 6154 19677
rect 6108 19605 6154 19635
rect 6108 19567 6114 19605
rect 6148 19567 6154 19605
rect 6108 19533 6154 19567
rect 6108 19499 6114 19533
rect 6148 19499 6154 19533
rect 6108 19465 6154 19499
rect 6108 19427 6114 19465
rect 6148 19427 6154 19465
rect 6108 19397 6154 19427
rect 6108 19355 6114 19397
rect 6148 19355 6154 19397
rect 6108 19329 6154 19355
rect 6108 19283 6114 19329
rect 6148 19283 6154 19329
rect 6108 19261 6154 19283
rect 6108 19211 6114 19261
rect 6148 19211 6154 19261
rect 6108 19193 6154 19211
rect 6108 19139 6114 19193
rect 6148 19139 6154 19193
rect 6108 19125 6154 19139
rect 6108 19067 6114 19125
rect 6148 19067 6154 19125
rect 6108 19057 6154 19067
rect 6108 18995 6114 19057
rect 6148 18995 6154 19057
rect 6108 18989 6154 18995
rect 6108 18923 6114 18989
rect 6148 18923 6154 18989
rect 6108 18921 6154 18923
rect 6108 18887 6114 18921
rect 6148 18887 6154 18921
rect 6108 18885 6154 18887
rect 6108 18819 6114 18885
rect 6148 18819 6154 18885
rect 6108 18813 6154 18819
rect 6108 18751 6114 18813
rect 6148 18751 6154 18813
rect 6108 18741 6154 18751
rect 6108 18683 6114 18741
rect 6148 18683 6154 18741
rect 6108 18669 6154 18683
rect 6108 18615 6114 18669
rect 6148 18615 6154 18669
rect 6108 18597 6154 18615
rect 6108 18547 6114 18597
rect 6148 18547 6154 18597
rect 6108 18525 6154 18547
rect 6108 18479 6114 18525
rect 6148 18479 6154 18525
rect 6108 18453 6154 18479
rect 6108 18411 6114 18453
rect 6148 18411 6154 18453
rect 6108 18381 6154 18411
rect 6108 18343 6114 18381
rect 6148 18343 6154 18381
rect 6108 18309 6154 18343
rect 6108 18275 6114 18309
rect 6148 18275 6154 18309
rect 6108 18241 6154 18275
rect 6108 18203 6114 18241
rect 6148 18203 6154 18241
rect 6108 18173 6154 18203
rect 6108 18131 6114 18173
rect 6148 18131 6154 18173
rect 6108 18105 6154 18131
rect 6108 18059 6114 18105
rect 6148 18059 6154 18105
rect 6108 18037 6154 18059
rect 6108 17987 6114 18037
rect 6148 17987 6154 18037
rect 6108 17969 6154 17987
rect 6108 17915 6114 17969
rect 6148 17915 6154 17969
rect 6108 17901 6154 17915
rect 6108 17843 6114 17901
rect 6148 17843 6154 17901
rect 6108 17833 6154 17843
rect 6108 17771 6114 17833
rect 6148 17771 6154 17833
rect 6108 17765 6154 17771
rect 6108 17699 6114 17765
rect 6148 17699 6154 17765
rect 6108 17697 6154 17699
rect 6108 17663 6114 17697
rect 6148 17663 6154 17697
rect 6108 17661 6154 17663
rect 6108 17595 6114 17661
rect 6148 17595 6154 17661
rect 6108 17589 6154 17595
rect 6108 17527 6114 17589
rect 6148 17527 6154 17589
rect 6108 17517 6154 17527
rect 6108 17459 6114 17517
rect 6148 17459 6154 17517
rect 6108 17445 6154 17459
rect 6108 17391 6114 17445
rect 6148 17391 6154 17445
rect 6108 17373 6154 17391
rect 6108 17323 6114 17373
rect 6148 17323 6154 17373
rect 6108 17301 6154 17323
rect 6108 17255 6114 17301
rect 6148 17255 6154 17301
rect 6108 17229 6154 17255
rect 6108 17187 6114 17229
rect 6148 17187 6154 17229
rect 6108 17157 6154 17187
rect 6108 17119 6114 17157
rect 6148 17119 6154 17157
rect 6108 17085 6154 17119
rect 6108 17051 6114 17085
rect 6148 17051 6154 17085
rect 6108 17017 6154 17051
rect 6108 16979 6114 17017
rect 6148 16979 6154 17017
rect 6108 16949 6154 16979
rect 6108 16907 6114 16949
rect 6148 16907 6154 16949
rect 6108 16881 6154 16907
rect 6108 16835 6114 16881
rect 6148 16835 6154 16881
rect 6108 16813 6154 16835
rect 6108 16763 6114 16813
rect 6148 16763 6154 16813
rect 6108 16745 6154 16763
rect 6108 16691 6114 16745
rect 6148 16691 6154 16745
rect 6108 16677 6154 16691
rect 6108 16619 6114 16677
rect 6148 16619 6154 16677
rect 6108 16609 6154 16619
rect 6108 16547 6114 16609
rect 6148 16547 6154 16609
rect 6108 16541 6154 16547
rect 6108 16475 6114 16541
rect 6148 16475 6154 16541
rect 6108 16473 6154 16475
rect 6108 16439 6114 16473
rect 6148 16439 6154 16473
rect 6108 16437 6154 16439
rect 6108 16371 6114 16437
rect 6148 16371 6154 16437
rect 6108 16365 6154 16371
rect 6108 16303 6114 16365
rect 6148 16303 6154 16365
rect 6108 16293 6154 16303
rect 6108 16235 6114 16293
rect 6148 16235 6154 16293
rect 6108 16221 6154 16235
rect 6108 16167 6114 16221
rect 6148 16167 6154 16221
rect 6108 16149 6154 16167
rect 6108 16099 6114 16149
rect 6148 16099 6154 16149
rect 6108 16077 6154 16099
rect 6108 16031 6114 16077
rect 6148 16031 6154 16077
rect 6108 16005 6154 16031
rect 6108 15963 6114 16005
rect 6148 15963 6154 16005
rect 6108 15933 6154 15963
rect 6108 15895 6114 15933
rect 6148 15895 6154 15933
rect 6108 15861 6154 15895
rect 6108 15827 6114 15861
rect 6148 15827 6154 15861
rect 6108 15793 6154 15827
rect 6108 15755 6114 15793
rect 6148 15755 6154 15793
rect 6108 15725 6154 15755
rect 6108 15683 6114 15725
rect 6148 15683 6154 15725
rect 6108 15657 6154 15683
rect 6108 15611 6114 15657
rect 6148 15611 6154 15657
rect 6108 15589 6154 15611
rect 6108 15539 6114 15589
rect 6148 15539 6154 15589
rect 6108 15521 6154 15539
rect 6108 15467 6114 15521
rect 6148 15467 6154 15521
rect 6108 15453 6154 15467
rect 6108 15395 6114 15453
rect 6148 15395 6154 15453
rect 6108 15385 6154 15395
rect 6108 15323 6114 15385
rect 6148 15323 6154 15385
rect 6108 15317 6154 15323
rect 6108 15251 6114 15317
rect 6148 15251 6154 15317
rect 6108 15249 6154 15251
rect 6108 15215 6114 15249
rect 6148 15215 6154 15249
rect 6108 15213 6154 15215
rect 6108 15147 6114 15213
rect 6148 15147 6154 15213
rect 6108 15141 6154 15147
rect 6108 15079 6114 15141
rect 6148 15079 6154 15141
rect 6108 15069 6154 15079
rect 6108 15011 6114 15069
rect 6148 15011 6154 15069
rect 6108 14997 6154 15011
rect 6108 14943 6114 14997
rect 6148 14943 6154 14997
rect 6108 14925 6154 14943
rect 6108 14875 6114 14925
rect 6148 14875 6154 14925
rect 6108 14853 6154 14875
rect 6108 14807 6114 14853
rect 6148 14807 6154 14853
rect 6108 14781 6154 14807
rect 6108 14739 6114 14781
rect 6148 14739 6154 14781
rect 6108 14709 6154 14739
rect 6108 14671 6114 14709
rect 6148 14671 6154 14709
rect 6108 14637 6154 14671
rect 6108 14603 6114 14637
rect 6148 14603 6154 14637
rect 6108 14569 6154 14603
rect 6108 14531 6114 14569
rect 6148 14531 6154 14569
rect 6108 14501 6154 14531
rect 6108 14459 6114 14501
rect 6148 14459 6154 14501
rect 6108 14433 6154 14459
rect 6108 14387 6114 14433
rect 6148 14387 6154 14433
rect 6108 14365 6154 14387
rect 6108 14315 6114 14365
rect 6148 14315 6154 14365
rect 6108 14297 6154 14315
rect 6108 14243 6114 14297
rect 6148 14243 6154 14297
rect 6108 14229 6154 14243
rect 6108 14171 6114 14229
rect 6148 14171 6154 14229
rect 6108 14161 6154 14171
rect 6108 14099 6114 14161
rect 6148 14099 6154 14161
rect 6108 14093 6154 14099
rect 6108 14027 6114 14093
rect 6148 14027 6154 14093
rect 6108 14025 6154 14027
rect 6108 13991 6114 14025
rect 6148 13991 6154 14025
rect 6108 13989 6154 13991
rect 6108 13923 6114 13989
rect 6148 13923 6154 13989
rect 6108 13917 6154 13923
rect 6108 13855 6114 13917
rect 6148 13855 6154 13917
rect 6108 13845 6154 13855
rect 6108 13787 6114 13845
rect 6148 13787 6154 13845
rect 6108 13773 6154 13787
rect 6108 13719 6114 13773
rect 6148 13719 6154 13773
rect 6108 13701 6154 13719
rect 6108 13651 6114 13701
rect 6148 13651 6154 13701
rect 6108 13629 6154 13651
rect 6108 13583 6114 13629
rect 6148 13583 6154 13629
rect 6108 13557 6154 13583
rect 6108 13515 6114 13557
rect 6148 13515 6154 13557
rect 6108 13485 6154 13515
rect 6108 13447 6114 13485
rect 6148 13447 6154 13485
rect 6108 13413 6154 13447
rect 6108 13379 6114 13413
rect 6148 13379 6154 13413
rect 6108 13345 6154 13379
rect 6108 13307 6114 13345
rect 6148 13307 6154 13345
rect 6108 13277 6154 13307
rect 6108 13235 6114 13277
rect 6148 13235 6154 13277
rect 6108 13209 6154 13235
rect 6108 13163 6114 13209
rect 6148 13163 6154 13209
rect 6108 13141 6154 13163
rect 6108 13091 6114 13141
rect 6148 13091 6154 13141
rect 6108 13073 6154 13091
rect 6108 13019 6114 13073
rect 6148 13019 6154 13073
rect 6108 13005 6154 13019
rect 6108 12947 6114 13005
rect 6148 12947 6154 13005
rect 6108 12937 6154 12947
rect 6108 12875 6114 12937
rect 6148 12875 6154 12937
rect 6108 12869 6154 12875
rect 6108 12803 6114 12869
rect 6148 12803 6154 12869
rect 6108 12801 6154 12803
rect 6108 12767 6114 12801
rect 6148 12767 6154 12801
rect 6108 12765 6154 12767
rect 6108 12699 6114 12765
rect 6148 12699 6154 12765
rect 6108 12693 6154 12699
rect 6108 12631 6114 12693
rect 6148 12631 6154 12693
rect 6108 12621 6154 12631
rect 6108 12563 6114 12621
rect 6148 12563 6154 12621
rect 6108 12549 6154 12563
rect 6108 12495 6114 12549
rect 6148 12495 6154 12549
rect 6108 12477 6154 12495
rect 6108 12427 6114 12477
rect 6148 12427 6154 12477
rect 6108 12405 6154 12427
rect 6108 12359 6114 12405
rect 6148 12359 6154 12405
rect 6108 12333 6154 12359
rect 6108 12291 6114 12333
rect 6148 12291 6154 12333
rect 6108 12261 6154 12291
rect 6108 12223 6114 12261
rect 6148 12223 6154 12261
rect 6108 12189 6154 12223
rect 6108 12155 6114 12189
rect 6148 12155 6154 12189
rect 6108 12121 6154 12155
rect 6108 12083 6114 12121
rect 6148 12083 6154 12121
rect 6108 12053 6154 12083
rect 6108 12011 6114 12053
rect 6148 12011 6154 12053
rect 6108 11985 6154 12011
rect 6108 11939 6114 11985
rect 6148 11939 6154 11985
rect 6108 11917 6154 11939
rect 6108 11867 6114 11917
rect 6148 11867 6154 11917
rect 6108 11849 6154 11867
rect 6108 11795 6114 11849
rect 6148 11795 6154 11849
rect 6108 11781 6154 11795
rect 6108 11723 6114 11781
rect 6148 11723 6154 11781
rect 6108 11713 6154 11723
rect 6108 11651 6114 11713
rect 6148 11651 6154 11713
rect 6108 11645 6154 11651
rect 6108 11579 6114 11645
rect 6148 11579 6154 11645
rect 6108 11577 6154 11579
rect 6108 11543 6114 11577
rect 6148 11543 6154 11577
rect 6108 11541 6154 11543
rect 6108 11475 6114 11541
rect 6148 11475 6154 11541
rect 6108 11469 6154 11475
rect 6108 11407 6114 11469
rect 6148 11407 6154 11469
rect 6108 11397 6154 11407
rect 6108 11339 6114 11397
rect 6148 11339 6154 11397
rect 6108 11325 6154 11339
rect 6108 11271 6114 11325
rect 6148 11271 6154 11325
rect 6108 11253 6154 11271
rect 6108 11203 6114 11253
rect 6148 11203 6154 11253
rect 6108 11181 6154 11203
rect 6108 11135 6114 11181
rect 6148 11135 6154 11181
rect 6108 11109 6154 11135
rect 6108 11067 6114 11109
rect 6148 11067 6154 11109
rect 6108 11037 6154 11067
rect 6108 10999 6114 11037
rect 6148 10999 6154 11037
rect 6108 10965 6154 10999
rect 6108 10931 6114 10965
rect 6148 10931 6154 10965
rect 6108 10897 6154 10931
rect 6108 10859 6114 10897
rect 6148 10859 6154 10897
rect 6108 10829 6154 10859
rect 6108 10787 6114 10829
rect 6148 10787 6154 10829
rect 6108 10761 6154 10787
rect 6108 10715 6114 10761
rect 6148 10715 6154 10761
rect 6108 10693 6154 10715
rect 6108 10643 6114 10693
rect 6148 10643 6154 10693
rect 6108 10625 6154 10643
rect 6108 10571 6114 10625
rect 6148 10571 6154 10625
rect 6108 10557 6154 10571
rect 6108 10499 6114 10557
rect 6148 10499 6154 10557
rect 6108 10489 6154 10499
rect 6108 10427 6114 10489
rect 6148 10427 6154 10489
rect 6108 10421 6154 10427
rect 6108 10355 6114 10421
rect 6148 10355 6154 10421
rect 6108 10353 6154 10355
rect 6108 10319 6114 10353
rect 6148 10319 6154 10353
rect 6108 10317 6154 10319
rect 6108 10251 6114 10317
rect 6148 10251 6154 10317
rect 6108 10245 6154 10251
rect 6108 10183 6114 10245
rect 6148 10183 6154 10245
rect 6108 10173 6154 10183
rect 6108 10115 6114 10173
rect 6148 10115 6154 10173
rect 6108 10101 6154 10115
rect 6108 10047 6114 10101
rect 6148 10047 6154 10101
rect 6108 10029 6154 10047
rect 6108 9979 6114 10029
rect 6148 9979 6154 10029
rect 6108 9957 6154 9979
rect 6108 9911 6114 9957
rect 6148 9911 6154 9957
rect 6108 9885 6154 9911
rect 6108 9843 6114 9885
rect 6148 9843 6154 9885
rect 6108 9813 6154 9843
rect 6108 9775 6114 9813
rect 6148 9775 6154 9813
rect 6108 9741 6154 9775
rect 6108 9707 6114 9741
rect 6148 9707 6154 9741
rect 6108 9673 6154 9707
rect 6108 9635 6114 9673
rect 6148 9635 6154 9673
rect 6108 9605 6154 9635
rect 6108 9563 6114 9605
rect 6148 9563 6154 9605
rect 6108 9537 6154 9563
rect 6108 9491 6114 9537
rect 6148 9491 6154 9537
rect 6108 9469 6154 9491
rect 6108 9419 6114 9469
rect 6148 9419 6154 9469
rect 6108 9401 6154 9419
rect 6108 9347 6114 9401
rect 6148 9347 6154 9401
rect 6108 9333 6154 9347
rect 6108 9275 6114 9333
rect 6148 9275 6154 9333
rect 6108 9265 6154 9275
rect 6108 9203 6114 9265
rect 6148 9203 6154 9265
rect 6108 9197 6154 9203
rect 6108 9131 6114 9197
rect 6148 9131 6154 9197
rect 6108 9129 6154 9131
rect 6108 9095 6114 9129
rect 6148 9095 6154 9129
rect 6108 9093 6154 9095
rect 6108 9027 6114 9093
rect 6148 9027 6154 9093
rect 6108 9021 6154 9027
rect 6108 8959 6114 9021
rect 6148 8959 6154 9021
rect 6108 8949 6154 8959
rect 6108 8891 6114 8949
rect 6148 8891 6154 8949
rect 6108 8877 6154 8891
rect 6108 8823 6114 8877
rect 6148 8823 6154 8877
rect 6108 8805 6154 8823
rect 6108 8755 6114 8805
rect 6148 8755 6154 8805
rect 6108 8733 6154 8755
rect 6108 8687 6114 8733
rect 6148 8687 6154 8733
rect 6108 8661 6154 8687
rect 6108 8619 6114 8661
rect 6148 8619 6154 8661
rect 6108 8589 6154 8619
rect 6108 8551 6114 8589
rect 6148 8551 6154 8589
rect 6108 8517 6154 8551
rect 6108 8483 6114 8517
rect 6148 8483 6154 8517
rect 6108 8449 6154 8483
rect 6108 8411 6114 8449
rect 6148 8411 6154 8449
rect 6108 8381 6154 8411
rect 6108 8339 6114 8381
rect 6148 8339 6154 8381
rect 6108 8313 6154 8339
rect 6108 8267 6114 8313
rect 6148 8267 6154 8313
rect 6108 8245 6154 8267
rect 6108 8195 6114 8245
rect 6148 8195 6154 8245
rect 6108 8177 6154 8195
rect 6108 8123 6114 8177
rect 6148 8123 6154 8177
rect 6108 8109 6154 8123
rect 6108 8051 6114 8109
rect 6148 8051 6154 8109
rect 6108 8041 6154 8051
rect 6108 7979 6114 8041
rect 6148 7979 6154 8041
rect 6108 7973 6154 7979
rect 6108 7907 6114 7973
rect 6148 7907 6154 7973
rect 6108 7905 6154 7907
rect 6108 7871 6114 7905
rect 6148 7871 6154 7905
rect 6108 7869 6154 7871
rect 6108 7803 6114 7869
rect 6148 7803 6154 7869
rect 6108 7797 6154 7803
rect 6108 7735 6114 7797
rect 6148 7735 6154 7797
rect 6108 7725 6154 7735
rect 6108 7667 6114 7725
rect 6148 7667 6154 7725
rect 6108 7653 6154 7667
rect 6108 7599 6114 7653
rect 6148 7599 6154 7653
rect 6108 7581 6154 7599
rect 6108 7531 6114 7581
rect 6148 7531 6154 7581
rect 6108 7509 6154 7531
rect 6108 7463 6114 7509
rect 6148 7463 6154 7509
rect 6108 7437 6154 7463
rect 6108 7395 6114 7437
rect 6148 7395 6154 7437
rect 6108 7365 6154 7395
rect 6108 7327 6114 7365
rect 6148 7327 6154 7365
rect 6108 7293 6154 7327
rect 6108 7259 6114 7293
rect 6148 7259 6154 7293
rect 6108 7225 6154 7259
rect 6108 7187 6114 7225
rect 6148 7187 6154 7225
rect 6108 7157 6154 7187
rect 6108 7115 6114 7157
rect 6148 7115 6154 7157
rect 6108 7089 6154 7115
rect 6108 7043 6114 7089
rect 6148 7043 6154 7089
rect 6108 7021 6154 7043
rect 6108 6971 6114 7021
rect 6148 6971 6154 7021
rect 6108 6953 6154 6971
rect 6108 6899 6114 6953
rect 6148 6899 6154 6953
rect 6108 6885 6154 6899
rect 6108 6827 6114 6885
rect 6148 6827 6154 6885
rect 6108 6817 6154 6827
rect 6108 6755 6114 6817
rect 6148 6755 6154 6817
rect 6108 6749 6154 6755
rect 6108 6682 6114 6749
rect 6148 6682 6154 6749
rect 6108 6681 6154 6682
rect 6108 6647 6114 6681
rect 6148 6647 6154 6681
rect 6108 6643 6154 6647
rect 6108 6579 6114 6643
rect 6148 6579 6154 6643
rect 6108 6570 6154 6579
rect 6108 6511 6114 6570
rect 6148 6511 6154 6570
rect 6108 6497 6154 6511
rect 6108 6443 6114 6497
rect 6148 6443 6154 6497
rect 6108 6424 6154 6443
rect 6108 6375 6114 6424
rect 6148 6375 6154 6424
rect 6108 6351 6154 6375
rect 6108 6307 6114 6351
rect 6148 6307 6154 6351
rect 6108 6278 6154 6307
rect 6108 6239 6114 6278
rect 6148 6239 6154 6278
rect 6108 6205 6154 6239
rect 6108 6171 6114 6205
rect 6148 6171 6154 6205
rect 6108 6137 6154 6171
rect 6108 6098 6114 6137
rect 6148 6098 6154 6137
rect 6108 6069 6154 6098
rect 6108 6025 6114 6069
rect 6148 6025 6154 6069
rect 6108 6001 6154 6025
rect 6108 5952 6114 6001
rect 6148 5952 6154 6001
rect 6108 5933 6154 5952
rect 6108 5879 6114 5933
rect 6148 5879 6154 5933
rect 6108 5865 6154 5879
rect 6108 5806 6114 5865
rect 6148 5806 6154 5865
rect 6108 5797 6154 5806
rect 6108 5733 6114 5797
rect 6148 5733 6154 5797
rect 6108 5729 6154 5733
rect 6108 5695 6114 5729
rect 6148 5695 6154 5729
rect 6108 5694 6154 5695
rect 6108 5627 6114 5694
rect 6148 5627 6154 5694
rect 6108 5621 6154 5627
rect 6108 5559 6114 5621
rect 6148 5559 6154 5621
rect 6108 5548 6154 5559
rect 6108 5491 6114 5548
rect 6148 5491 6154 5548
rect 6108 5475 6154 5491
rect 6108 5423 6114 5475
rect 6148 5423 6154 5475
rect 6108 5402 6154 5423
rect 6108 5355 6114 5402
rect 6148 5355 6154 5402
rect 6108 5329 6154 5355
rect 6108 5287 6114 5329
rect 6148 5287 6154 5329
rect 6108 5256 6154 5287
rect 6108 5219 6114 5256
rect 6148 5219 6154 5256
rect 6108 5185 6154 5219
rect 6108 5149 6114 5185
rect 6148 5149 6154 5185
rect 6108 5117 6154 5149
rect 6108 5076 6114 5117
rect 6148 5076 6154 5117
rect 6108 5049 6154 5076
rect 6108 5003 6114 5049
rect 6148 5003 6154 5049
rect 6108 4981 6154 5003
rect 6108 4930 6114 4981
rect 6148 4930 6154 4981
rect 6108 4913 6154 4930
rect 6108 4857 6114 4913
rect 6148 4857 6154 4913
rect 6108 4845 6154 4857
rect 6108 4784 6114 4845
rect 6148 4784 6154 4845
rect 6108 4777 6154 4784
rect 6108 4711 6114 4777
rect 6148 4711 6154 4777
rect 6108 4709 6154 4711
rect 6108 4675 6114 4709
rect 6148 4675 6154 4709
rect 6108 4672 6154 4675
rect 6108 4607 6114 4672
rect 6148 4607 6154 4672
rect 6108 4599 6154 4607
rect 6108 4539 6114 4599
rect 6148 4539 6154 4599
rect 6108 4526 6154 4539
rect 6108 4471 6114 4526
rect 6148 4471 6154 4526
rect 6108 4453 6154 4471
rect 6108 4403 6114 4453
rect 6148 4403 6154 4453
rect 6108 4380 6154 4403
rect 6108 4335 6114 4380
rect 6148 4335 6154 4380
rect 6108 4307 6154 4335
rect 6108 4267 6114 4307
rect 6148 4267 6154 4307
rect 6108 4234 6154 4267
rect 6108 4199 6114 4234
rect 6148 4199 6154 4234
rect 6108 4165 6154 4199
rect 6108 4127 6114 4165
rect 6148 4127 6154 4165
rect 6108 4097 6154 4127
rect 6108 4054 6114 4097
rect 6148 4054 6154 4097
rect 6108 4029 6154 4054
rect 6108 3981 6114 4029
rect 6148 3981 6154 4029
rect 6108 3961 6154 3981
rect 6108 3908 6114 3961
rect 6148 3908 6154 3961
rect 6108 3893 6154 3908
rect 6108 3835 6114 3893
rect 6148 3835 6154 3893
rect 6108 3825 6154 3835
rect 6108 3762 6114 3825
rect 6148 3762 6154 3825
rect 6108 3757 6154 3762
rect 6108 3655 6114 3757
rect 6148 3655 6154 3757
rect 6108 3650 6154 3655
rect 6108 3587 6114 3650
rect 6148 3587 6154 3650
rect 6108 3577 6154 3587
rect 6108 3519 6114 3577
rect 6148 3519 6154 3577
rect 6108 3504 6154 3519
rect 3966 3465 4012 3467
rect 3966 3431 3972 3465
rect 4006 3431 4012 3465
rect 3966 3429 4012 3431
rect 3966 3363 3972 3429
rect 4006 3363 4012 3429
rect 1824 3315 1830 3357
rect 1864 3315 1870 3357
rect 1824 3285 1870 3315
rect 1824 3247 1830 3285
rect 1864 3247 1870 3285
rect 1824 3219 1870 3247
rect 3966 3357 4012 3363
rect 4142 3453 4158 3473
rect 4192 3453 4208 3473
rect 4142 3415 4208 3453
rect 4142 3361 4158 3415
rect 4192 3361 4208 3415
rect 4260 3453 4276 3473
rect 4310 3453 4326 3473
rect 4260 3415 4326 3453
rect 4260 3361 4276 3415
rect 4310 3361 4326 3415
rect 4378 3453 4394 3473
rect 4428 3453 4444 3473
rect 4378 3415 4444 3453
rect 4378 3361 4394 3415
rect 4428 3361 4444 3415
rect 4496 3453 4512 3473
rect 4546 3453 4562 3473
rect 4496 3415 4562 3453
rect 4496 3361 4512 3415
rect 4546 3361 4562 3415
rect 4614 3453 4630 3473
rect 4664 3453 4680 3473
rect 4614 3415 4680 3453
rect 4614 3361 4630 3415
rect 4664 3361 4680 3415
rect 4732 3453 4748 3473
rect 4782 3453 4798 3473
rect 4732 3415 4798 3453
rect 4732 3361 4748 3415
rect 4782 3361 4798 3415
rect 4850 3453 4866 3473
rect 4900 3453 4916 3473
rect 4850 3415 4916 3453
rect 4850 3361 4866 3415
rect 4900 3361 4916 3415
rect 4968 3453 4984 3473
rect 5018 3453 5034 3473
rect 4968 3415 5034 3453
rect 4968 3361 4984 3415
rect 5018 3361 5034 3415
rect 5086 3453 5102 3472
rect 5136 3453 5152 3472
rect 5086 3415 5152 3453
rect 5086 3361 5102 3415
rect 5136 3361 5152 3415
rect 5086 3360 5152 3361
rect 5204 3452 5220 3472
rect 5254 3452 5270 3472
rect 5204 3414 5270 3452
rect 5204 3361 5220 3414
rect 5254 3361 5270 3414
rect 5204 3360 5270 3361
rect 5322 3452 5338 3472
rect 5372 3452 5388 3472
rect 5322 3414 5388 3452
rect 5322 3361 5338 3414
rect 5372 3361 5388 3414
rect 5322 3360 5388 3361
rect 5440 3452 5456 3472
rect 5490 3452 5506 3472
rect 5440 3414 5506 3452
rect 5440 3361 5456 3414
rect 5490 3361 5506 3414
rect 5440 3360 5506 3361
rect 5558 3452 5574 3472
rect 5608 3452 5624 3472
rect 5558 3414 5624 3452
rect 5558 3361 5574 3414
rect 5608 3361 5624 3414
rect 5558 3360 5624 3361
rect 5676 3452 5692 3472
rect 5726 3452 5742 3472
rect 5676 3414 5742 3452
rect 5676 3361 5692 3414
rect 5726 3361 5742 3414
rect 5676 3360 5742 3361
rect 5794 3452 5810 3472
rect 5844 3452 5860 3472
rect 5794 3414 5860 3452
rect 5794 3361 5810 3414
rect 5844 3361 5860 3414
rect 5794 3360 5860 3361
rect 5912 3452 5928 3472
rect 5962 3452 5978 3472
rect 5912 3414 5978 3452
rect 5912 3361 5928 3414
rect 5962 3361 5978 3414
rect 5912 3360 5978 3361
rect 6108 3451 6114 3504
rect 6148 3451 6154 3504
rect 6108 3431 6154 3451
rect 6108 3383 6114 3431
rect 6148 3383 6154 3431
rect 3966 3295 3972 3357
rect 4006 3295 4012 3357
rect 3966 3285 4012 3295
rect 3966 3251 3972 3285
rect 4006 3251 4012 3285
rect 3966 3219 4012 3251
rect 6108 3358 6154 3383
rect 6108 3315 6114 3358
rect 6148 3315 6154 3358
rect 6108 3285 6154 3315
rect 6108 3247 6114 3285
rect 6148 3247 6154 3285
rect 6108 3219 6154 3247
rect -258 3213 6154 3219
rect -258 3179 -184 3213
rect -146 3179 -116 3213
rect -73 3179 -48 3213
rect 0 3179 20 3213
rect 73 3179 88 3213
rect 146 3179 156 3213
rect 219 3179 224 3213
rect 326 3179 331 3213
rect 394 3179 404 3213
rect 462 3179 477 3213
rect 530 3179 550 3213
rect 598 3179 623 3213
rect 666 3179 696 3213
rect 734 3179 768 3213
rect 803 3179 836 3213
rect 876 3179 904 3213
rect 949 3179 972 3213
rect 1022 3179 1040 3213
rect 1095 3179 1108 3213
rect 1168 3179 1176 3213
rect 1241 3179 1244 3213
rect 1278 3179 1280 3213
rect 1346 3179 1353 3213
rect 1414 3179 1426 3213
rect 1482 3179 1499 3213
rect 1550 3179 1572 3213
rect 1618 3179 1645 3213
rect 1686 3179 1718 3213
rect 1754 3179 1791 3213
rect 1825 3179 1864 3213
rect 1898 3179 1932 3213
rect 1971 3179 2000 3213
rect 2044 3179 2068 3213
rect 2116 3179 2136 3213
rect 2188 3179 2204 3213
rect 2260 3179 2272 3213
rect 2332 3179 2340 3213
rect 2404 3179 2408 3213
rect 2510 3179 2514 3213
rect 2578 3179 2586 3213
rect 2646 3179 2658 3213
rect 2714 3179 2730 3213
rect 2782 3179 2802 3213
rect 2850 3179 2874 3213
rect 2918 3179 2946 3213
rect 2986 3179 3018 3213
rect 3054 3179 3088 3213
rect 3124 3179 3156 3213
rect 3196 3179 3224 3213
rect 3268 3179 3292 3213
rect 3340 3179 3360 3213
rect 3412 3179 3428 3213
rect 3484 3179 3496 3213
rect 3556 3179 3564 3213
rect 3628 3179 3632 3213
rect 3734 3179 3738 3213
rect 3802 3179 3810 3213
rect 3870 3179 3882 3213
rect 3938 3179 3954 3213
rect 3988 3179 4026 3213
rect 4074 3179 4098 3213
rect 4142 3179 4170 3213
rect 4210 3179 4242 3213
rect 4278 3179 4312 3213
rect 4348 3179 4380 3213
rect 4420 3179 4448 3213
rect 4492 3179 4516 3213
rect 4564 3179 4584 3213
rect 4636 3179 4652 3213
rect 4708 3179 4720 3213
rect 4780 3179 4788 3213
rect 4852 3179 4856 3213
rect 4958 3179 4962 3213
rect 5026 3179 5034 3213
rect 5094 3179 5106 3213
rect 5162 3179 5178 3213
rect 5230 3179 5250 3213
rect 5298 3179 5322 3213
rect 5366 3179 5394 3213
rect 5434 3179 5466 3213
rect 5502 3179 5536 3213
rect 5572 3179 5604 3213
rect 5644 3179 5672 3213
rect 5716 3179 5740 3213
rect 5788 3179 5808 3213
rect 5860 3179 5876 3213
rect 5932 3179 5944 3213
rect 6004 3179 6012 3213
rect 6076 3179 6154 3213
rect -258 3173 6154 3179
rect 9082 38757 14980 38762
rect 9082 38756 9206 38757
rect 9240 38756 9274 38757
rect 9082 38722 9162 38756
rect 9196 38723 9206 38756
rect 9271 38723 9274 38756
rect 9308 38756 9342 38757
rect 9308 38723 9312 38756
rect 9376 38723 9410 38757
rect 9444 38756 9478 38757
rect 9512 38756 9546 38757
rect 9580 38756 9614 38757
rect 9648 38756 9682 38757
rect 9716 38756 9750 38757
rect 9784 38756 9818 38757
rect 9456 38723 9478 38756
rect 9528 38723 9546 38756
rect 9600 38723 9614 38756
rect 9672 38723 9682 38756
rect 9744 38723 9750 38756
rect 9816 38723 9818 38756
rect 9852 38756 9886 38757
rect 9920 38756 9954 38757
rect 9988 38756 10022 38757
rect 10056 38756 10090 38757
rect 10124 38756 10158 38757
rect 10192 38756 10294 38757
rect 10328 38756 10362 38757
rect 9852 38723 9854 38756
rect 9920 38723 9926 38756
rect 9988 38723 9998 38756
rect 10056 38723 10070 38756
rect 10124 38723 10142 38756
rect 10192 38723 10214 38756
rect 9196 38722 9237 38723
rect 9271 38722 9312 38723
rect 9346 38722 9422 38723
rect 9456 38722 9494 38723
rect 9528 38722 9566 38723
rect 9600 38722 9638 38723
rect 9672 38722 9710 38723
rect 9744 38722 9782 38723
rect 9816 38722 9854 38723
rect 9888 38722 9926 38723
rect 9960 38722 9998 38723
rect 10032 38722 10070 38723
rect 10104 38722 10142 38723
rect 10176 38722 10214 38723
rect 10248 38722 10286 38756
rect 10328 38723 10358 38756
rect 10396 38723 10430 38757
rect 10464 38723 10498 38757
rect 10532 38756 10566 38757
rect 10600 38756 10634 38757
rect 10668 38756 10702 38757
rect 10736 38756 10770 38757
rect 10804 38756 10838 38757
rect 10872 38756 10906 38757
rect 10940 38756 10974 38757
rect 11008 38756 11042 38757
rect 10536 38723 10566 38756
rect 10608 38723 10634 38756
rect 10680 38723 10702 38756
rect 10752 38723 10770 38756
rect 10824 38723 10838 38756
rect 10896 38723 10906 38756
rect 10968 38723 10974 38756
rect 11040 38723 11042 38756
rect 11076 38756 11110 38757
rect 11144 38756 11178 38757
rect 11212 38756 11246 38757
rect 11280 38756 11314 38757
rect 11348 38756 11512 38757
rect 11076 38723 11078 38756
rect 11144 38723 11150 38756
rect 11212 38723 11222 38756
rect 11280 38723 11294 38756
rect 11348 38723 11366 38756
rect 10320 38722 10358 38723
rect 10392 38722 10430 38723
rect 10464 38722 10502 38723
rect 10536 38722 10574 38723
rect 10608 38722 10646 38723
rect 10680 38722 10718 38723
rect 10752 38722 10790 38723
rect 10824 38722 10862 38723
rect 10896 38722 10934 38723
rect 10968 38722 11006 38723
rect 11040 38722 11078 38723
rect 11112 38722 11150 38723
rect 11184 38722 11222 38723
rect 11256 38722 11294 38723
rect 11328 38722 11366 38723
rect 11400 38722 11438 38756
rect 11472 38722 11510 38756
rect 11546 38723 11580 38757
rect 11614 38756 11648 38757
rect 11682 38756 11716 38757
rect 11750 38756 11784 38757
rect 11818 38756 11852 38757
rect 11886 38756 11920 38757
rect 11954 38756 11988 38757
rect 12022 38756 12056 38757
rect 11617 38723 11648 38756
rect 11690 38723 11716 38756
rect 11763 38723 11784 38756
rect 11836 38723 11852 38756
rect 11909 38723 11920 38756
rect 11982 38723 11988 38756
rect 12055 38723 12056 38756
rect 12090 38756 12124 38757
rect 12158 38756 12192 38757
rect 12226 38756 12260 38757
rect 12294 38756 12328 38757
rect 12362 38756 12396 38757
rect 12430 38756 12464 38757
rect 12090 38723 12094 38756
rect 12158 38723 12167 38756
rect 12226 38723 12240 38756
rect 12294 38723 12313 38756
rect 12362 38723 12386 38756
rect 12430 38723 12459 38756
rect 12498 38723 12532 38757
rect 12566 38723 12600 38757
rect 12634 38756 12668 38757
rect 12702 38756 12736 38757
rect 12770 38756 12804 38757
rect 12838 38756 12872 38757
rect 12906 38756 12940 38757
rect 12974 38756 13008 38757
rect 12639 38723 12668 38756
rect 12712 38723 12736 38756
rect 12785 38723 12804 38756
rect 12858 38723 12872 38756
rect 12931 38723 12940 38756
rect 13004 38723 13008 38756
rect 13042 38756 13076 38757
rect 13110 38756 13144 38757
rect 13178 38756 13280 38757
rect 13314 38756 13348 38757
rect 13382 38756 13416 38757
rect 13450 38756 13484 38757
rect 13042 38723 13043 38756
rect 13110 38723 13116 38756
rect 13178 38723 13189 38756
rect 11544 38722 11583 38723
rect 11617 38722 11656 38723
rect 11690 38722 11729 38723
rect 11763 38722 11802 38723
rect 11836 38722 11875 38723
rect 11909 38722 11948 38723
rect 11982 38722 12021 38723
rect 12055 38722 12094 38723
rect 12128 38722 12167 38723
rect 12201 38722 12240 38723
rect 12274 38722 12313 38723
rect 12347 38722 12386 38723
rect 12420 38722 12459 38723
rect 12493 38722 12532 38723
rect 12566 38722 12605 38723
rect 12639 38722 12678 38723
rect 12712 38722 12751 38723
rect 12785 38722 12824 38723
rect 12858 38722 12897 38723
rect 12931 38722 12970 38723
rect 13004 38722 13043 38723
rect 13077 38722 13116 38723
rect 13150 38722 13189 38723
rect 13223 38722 13262 38756
rect 13314 38723 13335 38756
rect 13382 38723 13408 38756
rect 13450 38723 13481 38756
rect 13518 38723 13552 38757
rect 13586 38756 13620 38757
rect 13654 38756 13688 38757
rect 13722 38756 13756 38757
rect 13790 38756 13824 38757
rect 13858 38756 13892 38757
rect 13926 38756 13960 38757
rect 13994 38756 14028 38757
rect 13588 38723 13620 38756
rect 13661 38723 13688 38756
rect 13734 38723 13756 38756
rect 13807 38723 13824 38756
rect 13880 38723 13892 38756
rect 13953 38723 13960 38756
rect 14026 38723 14028 38756
rect 14062 38756 14096 38757
rect 14130 38756 14164 38757
rect 14198 38756 14232 38757
rect 14266 38756 14300 38757
rect 14334 38756 14368 38757
rect 14402 38756 14436 38757
rect 14470 38756 14504 38757
rect 14062 38723 14065 38756
rect 14130 38723 14138 38756
rect 14198 38723 14211 38756
rect 14266 38723 14284 38756
rect 14334 38723 14357 38756
rect 14402 38723 14430 38756
rect 14470 38723 14503 38756
rect 14538 38723 14572 38757
rect 14606 38756 14640 38757
rect 14674 38756 14708 38757
rect 14742 38756 14776 38757
rect 14810 38756 14844 38757
rect 14878 38756 14980 38757
rect 14610 38723 14640 38756
rect 14683 38723 14708 38756
rect 14756 38723 14776 38756
rect 14829 38723 14844 38756
rect 13296 38722 13335 38723
rect 13369 38722 13408 38723
rect 13442 38722 13481 38723
rect 13515 38722 13554 38723
rect 13588 38722 13627 38723
rect 13661 38722 13700 38723
rect 13734 38722 13773 38723
rect 13807 38722 13846 38723
rect 13880 38722 13919 38723
rect 13953 38722 13992 38723
rect 14026 38722 14065 38723
rect 14099 38722 14138 38723
rect 14172 38722 14211 38723
rect 14245 38722 14284 38723
rect 14318 38722 14357 38723
rect 14391 38722 14430 38723
rect 14464 38722 14503 38723
rect 14537 38722 14576 38723
rect 14610 38722 14649 38723
rect 14683 38722 14722 38723
rect 14756 38722 14795 38723
rect 14829 38722 14868 38723
rect 14902 38722 14980 38756
rect 9082 38716 14980 38722
rect 9082 38689 9128 38716
rect 9082 38650 9088 38689
rect 9122 38650 9128 38689
rect 9082 38621 9128 38650
rect 9082 38577 9088 38621
rect 9122 38577 9128 38621
rect 9082 38553 9128 38577
rect 9082 38504 9088 38553
rect 9122 38504 9128 38553
rect 9082 38485 9128 38504
rect 9082 38431 9088 38485
rect 9122 38431 9128 38485
rect 9082 38417 9128 38431
rect 9082 38358 9088 38417
rect 9122 38358 9128 38417
rect 9082 38349 9128 38358
rect 9082 38285 9088 38349
rect 9122 38285 9128 38349
rect 9082 38281 9128 38285
rect 9082 38247 9088 38281
rect 9122 38247 9128 38281
rect 9082 38246 9128 38247
rect 9082 38179 9088 38246
rect 9122 38179 9128 38246
rect 9082 38173 9128 38179
rect 9082 38111 9088 38173
rect 9122 38111 9128 38173
rect 9082 38100 9128 38111
rect 9082 38043 9088 38100
rect 9122 38043 9128 38100
rect 9082 38027 9128 38043
rect 9082 37975 9088 38027
rect 9122 37975 9128 38027
rect 9082 37954 9128 37975
rect 9082 37907 9088 37954
rect 9122 37907 9128 37954
rect 9082 37881 9128 37907
rect 9082 37839 9088 37881
rect 9122 37839 9128 37881
rect 9082 37808 9128 37839
rect 9082 37771 9088 37808
rect 9122 37771 9128 37808
rect 9082 37737 9128 37771
rect 9082 37701 9088 37737
rect 9122 37701 9128 37737
rect 9082 37669 9128 37701
rect 9082 37628 9088 37669
rect 9122 37628 9128 37669
rect 9082 37601 9128 37628
rect 9082 37555 9088 37601
rect 9122 37555 9128 37601
rect 9082 37533 9128 37555
rect 9082 37482 9088 37533
rect 9122 37482 9128 37533
rect 9082 37465 9128 37482
rect 9082 37409 9088 37465
rect 9122 37409 9128 37465
rect 9082 37397 9128 37409
rect 9082 37336 9088 37397
rect 9122 37336 9128 37397
rect 9082 37329 9128 37336
rect 9082 37263 9088 37329
rect 9122 37263 9128 37329
rect 9082 37261 9128 37263
rect 9082 37227 9088 37261
rect 9122 37227 9128 37261
rect 9082 37224 9128 37227
rect 9082 37159 9088 37224
rect 9122 37159 9128 37224
rect 9082 37151 9128 37159
rect 9082 37091 9088 37151
rect 9122 37091 9128 37151
rect 9082 37078 9128 37091
rect 9082 37023 9088 37078
rect 9122 37023 9128 37078
rect 9082 37005 9128 37023
rect 9082 36955 9088 37005
rect 9122 36955 9128 37005
rect 9082 36932 9128 36955
rect 9082 36887 9088 36932
rect 9122 36887 9128 36932
rect 9082 36859 9128 36887
rect 9082 36819 9088 36859
rect 9122 36819 9128 36859
rect 9082 36786 9128 36819
rect 9082 36751 9088 36786
rect 9122 36751 9128 36786
rect 9082 36717 9128 36751
rect 9082 36679 9088 36717
rect 9122 36679 9128 36717
rect 9082 36649 9128 36679
rect 9082 36606 9088 36649
rect 9122 36606 9128 36649
rect 9082 36581 9128 36606
rect 9082 36533 9088 36581
rect 9122 36533 9128 36581
rect 9082 36513 9128 36533
rect 9082 36460 9088 36513
rect 9122 36460 9128 36513
rect 9082 36445 9128 36460
rect 9082 36387 9088 36445
rect 9122 36387 9128 36445
rect 9082 36377 9128 36387
rect 9082 36314 9088 36377
rect 9122 36314 9128 36377
rect 9082 36309 9128 36314
rect 9082 36207 9088 36309
rect 9122 36207 9128 36309
rect 9082 36202 9128 36207
rect 9082 36139 9088 36202
rect 9122 36139 9128 36202
rect 9082 36129 9128 36139
rect 9082 36071 9088 36129
rect 9122 36071 9128 36129
rect 9082 36056 9128 36071
rect 9082 36003 9088 36056
rect 9122 36003 9128 36056
rect 9082 35983 9128 36003
rect 9082 35935 9088 35983
rect 9122 35935 9128 35983
rect 9082 35910 9128 35935
rect 9082 35867 9088 35910
rect 9122 35867 9128 35910
rect 9082 35837 9128 35867
rect 9082 35799 9088 35837
rect 9122 35799 9128 35837
rect 9082 35765 9128 35799
rect 9082 35730 9088 35765
rect 9122 35730 9128 35765
rect 9082 35697 9128 35730
rect 9082 35657 9088 35697
rect 9122 35657 9128 35697
rect 9082 35629 9128 35657
rect 9082 35584 9088 35629
rect 9122 35584 9128 35629
rect 9082 35561 9128 35584
rect 9082 35511 9088 35561
rect 9122 35511 9128 35561
rect 9082 35493 9128 35511
rect 9082 35438 9088 35493
rect 9122 35438 9128 35493
rect 9082 35425 9128 35438
rect 9082 35365 9088 35425
rect 9122 35365 9128 35425
rect 9082 35357 9128 35365
rect 9082 35292 9088 35357
rect 9122 35292 9128 35357
rect 9082 35289 9128 35292
rect 9082 35255 9088 35289
rect 9122 35255 9128 35289
rect 9082 35253 9128 35255
rect 9082 35187 9088 35253
rect 9122 35187 9128 35253
rect 9082 35180 9128 35187
rect 9082 35119 9088 35180
rect 9122 35119 9128 35180
rect 9082 35108 9128 35119
rect 9082 35051 9088 35108
rect 9122 35051 9128 35108
rect 9082 35036 9128 35051
rect 9082 34983 9088 35036
rect 9122 34983 9128 35036
rect 9082 34964 9128 34983
rect 9082 34915 9088 34964
rect 9122 34915 9128 34964
rect 9082 34892 9128 34915
rect 9082 34847 9088 34892
rect 9122 34847 9128 34892
rect 9082 34820 9128 34847
rect 9082 34779 9088 34820
rect 9122 34779 9128 34820
rect 9082 34748 9128 34779
rect 9082 34711 9088 34748
rect 9122 34711 9128 34748
rect 9082 34677 9128 34711
rect 9082 34642 9088 34677
rect 9122 34642 9128 34677
rect 9082 34609 9128 34642
rect 9082 34570 9088 34609
rect 9122 34570 9128 34609
rect 9082 34541 9128 34570
rect 9082 34498 9088 34541
rect 9122 34498 9128 34541
rect 9082 34473 9128 34498
rect 9082 34426 9088 34473
rect 9122 34426 9128 34473
rect 9082 34405 9128 34426
rect 9082 34354 9088 34405
rect 9122 34354 9128 34405
rect 9082 34337 9128 34354
rect 9082 34282 9088 34337
rect 9122 34282 9128 34337
rect 9082 34269 9128 34282
rect 9082 34210 9088 34269
rect 9122 34210 9128 34269
rect 9082 34201 9128 34210
rect 9082 34138 9088 34201
rect 9122 34138 9128 34201
rect 9082 34133 9128 34138
rect 9082 34066 9088 34133
rect 9122 34066 9128 34133
rect 9082 34065 9128 34066
rect 9082 34031 9088 34065
rect 9122 34031 9128 34065
rect 9082 34028 9128 34031
rect 9082 33963 9088 34028
rect 9122 33963 9128 34028
rect 9082 33956 9128 33963
rect 9082 33895 9088 33956
rect 9122 33895 9128 33956
rect 9082 33884 9128 33895
rect 9082 33827 9088 33884
rect 9122 33827 9128 33884
rect 9082 33812 9128 33827
rect 9082 33759 9088 33812
rect 9122 33759 9128 33812
rect 9082 33740 9128 33759
rect 9082 33691 9088 33740
rect 9122 33691 9128 33740
rect 9082 33668 9128 33691
rect 9082 33623 9088 33668
rect 9122 33623 9128 33668
rect 9082 33596 9128 33623
rect 9082 33555 9088 33596
rect 9122 33555 9128 33596
rect 9082 33524 9128 33555
rect 9082 33487 9088 33524
rect 9122 33487 9128 33524
rect 9082 33453 9128 33487
rect 9082 33418 9088 33453
rect 9122 33418 9128 33453
rect 9082 33385 9128 33418
rect 9082 33346 9088 33385
rect 9122 33346 9128 33385
rect 9082 33317 9128 33346
rect 9082 33274 9088 33317
rect 9122 33274 9128 33317
rect 9082 33249 9128 33274
rect 9082 33202 9088 33249
rect 9122 33202 9128 33249
rect 9082 33181 9128 33202
rect 9082 33130 9088 33181
rect 9122 33130 9128 33181
rect 9082 33113 9128 33130
rect 9082 33058 9088 33113
rect 9122 33058 9128 33113
rect 9082 33045 9128 33058
rect 9082 32986 9088 33045
rect 9122 32986 9128 33045
rect 9082 32977 9128 32986
rect 9082 32914 9088 32977
rect 9122 32914 9128 32977
rect 9082 32909 9128 32914
rect 9082 32842 9088 32909
rect 9122 32842 9128 32909
rect 9082 32841 9128 32842
rect 9082 32807 9088 32841
rect 9122 32807 9128 32841
rect 9082 32804 9128 32807
rect 9082 32739 9088 32804
rect 9122 32739 9128 32804
rect 9082 32732 9128 32739
rect 9082 32671 9088 32732
rect 9122 32671 9128 32732
rect 9082 32660 9128 32671
rect 9082 32603 9088 32660
rect 9122 32603 9128 32660
rect 9082 32588 9128 32603
rect 9082 32535 9088 32588
rect 9122 32535 9128 32588
rect 9082 32516 9128 32535
rect 9082 32467 9088 32516
rect 9122 32467 9128 32516
rect 9082 32444 9128 32467
rect 9082 32399 9088 32444
rect 9122 32399 9128 32444
rect 9082 32372 9128 32399
rect 9082 32331 9088 32372
rect 9122 32331 9128 32372
rect 9082 32300 9128 32331
rect 9082 32263 9088 32300
rect 9122 32263 9128 32300
rect 9082 32229 9128 32263
rect 9082 32194 9088 32229
rect 9122 32194 9128 32229
rect 9082 32161 9128 32194
rect 9082 32122 9088 32161
rect 9122 32122 9128 32161
rect 9082 32093 9128 32122
rect 9082 32050 9088 32093
rect 9122 32050 9128 32093
rect 9082 32025 9128 32050
rect 9082 31978 9088 32025
rect 9122 31978 9128 32025
rect 9082 31957 9128 31978
rect 9082 31906 9088 31957
rect 9122 31906 9128 31957
rect 9082 31889 9128 31906
rect 9082 31834 9088 31889
rect 9122 31834 9128 31889
rect 9082 31821 9128 31834
rect 9082 31762 9088 31821
rect 9122 31762 9128 31821
rect 9082 31753 9128 31762
rect 9082 31690 9088 31753
rect 9122 31690 9128 31753
rect 9082 31685 9128 31690
rect 9082 31618 9088 31685
rect 9122 31618 9128 31685
rect 9082 31617 9128 31618
rect 9082 31583 9088 31617
rect 9122 31583 9128 31617
rect 9082 31580 9128 31583
rect 9082 31515 9088 31580
rect 9122 31515 9128 31580
rect 9082 31508 9128 31515
rect 9082 31447 9088 31508
rect 9122 31447 9128 31508
rect 9082 31436 9128 31447
rect 9082 31379 9088 31436
rect 9122 31379 9128 31436
rect 9082 31364 9128 31379
rect 9082 31311 9088 31364
rect 9122 31311 9128 31364
rect 9082 31292 9128 31311
rect 9082 31243 9088 31292
rect 9122 31243 9128 31292
rect 9082 31220 9128 31243
rect 9082 31175 9088 31220
rect 9122 31175 9128 31220
rect 9082 31148 9128 31175
rect 9082 31107 9088 31148
rect 9122 31107 9128 31148
rect 9082 31076 9128 31107
rect 9082 31039 9088 31076
rect 9122 31039 9128 31076
rect 9082 31005 9128 31039
rect 9082 30970 9088 31005
rect 9122 30970 9128 31005
rect 9082 30937 9128 30970
rect 9082 30898 9088 30937
rect 9122 30898 9128 30937
rect 9082 30869 9128 30898
rect 9082 30826 9088 30869
rect 9122 30826 9128 30869
rect 9082 30801 9128 30826
rect 9082 30754 9088 30801
rect 9122 30754 9128 30801
rect 9082 30733 9128 30754
rect 9082 30682 9088 30733
rect 9122 30682 9128 30733
rect 9082 30665 9128 30682
rect 9082 30610 9088 30665
rect 9122 30610 9128 30665
rect 9082 30597 9128 30610
rect 9082 30538 9088 30597
rect 9122 30538 9128 30597
rect 9082 30529 9128 30538
rect 9082 30466 9088 30529
rect 9122 30466 9128 30529
rect 9082 30461 9128 30466
rect 9082 30394 9088 30461
rect 9122 30394 9128 30461
rect 9082 30393 9128 30394
rect 9082 30359 9088 30393
rect 9122 30359 9128 30393
rect 9082 30356 9128 30359
rect 9082 30291 9088 30356
rect 9122 30291 9128 30356
rect 9082 30284 9128 30291
rect 9082 30223 9088 30284
rect 9122 30223 9128 30284
rect 9082 30212 9128 30223
rect 9082 30155 9088 30212
rect 9122 30155 9128 30212
rect 9082 30140 9128 30155
rect 9082 30087 9088 30140
rect 9122 30087 9128 30140
rect 9082 30068 9128 30087
rect 9082 30019 9088 30068
rect 9122 30019 9128 30068
rect 9082 29996 9128 30019
rect 9082 29951 9088 29996
rect 9122 29951 9128 29996
rect 9082 29924 9128 29951
rect 9082 29883 9088 29924
rect 9122 29883 9128 29924
rect 9082 29852 9128 29883
rect 9082 29815 9088 29852
rect 9122 29815 9128 29852
rect 9082 29781 9128 29815
rect 9082 29746 9088 29781
rect 9122 29746 9128 29781
rect 9082 29713 9128 29746
rect 9082 29674 9088 29713
rect 9122 29674 9128 29713
rect 9082 29645 9128 29674
rect 9082 29602 9088 29645
rect 9122 29602 9128 29645
rect 9082 29577 9128 29602
rect 9082 29530 9088 29577
rect 9122 29530 9128 29577
rect 9082 29509 9128 29530
rect 9082 29458 9088 29509
rect 9122 29458 9128 29509
rect 9082 29441 9128 29458
rect 9082 29386 9088 29441
rect 9122 29386 9128 29441
rect 9082 29373 9128 29386
rect 9082 29314 9088 29373
rect 9122 29314 9128 29373
rect 9082 29305 9128 29314
rect 9082 29242 9088 29305
rect 9122 29242 9128 29305
rect 9082 29237 9128 29242
rect 9082 29170 9088 29237
rect 9122 29170 9128 29237
rect 9082 29169 9128 29170
rect 9082 29135 9088 29169
rect 9122 29135 9128 29169
rect 9082 29132 9128 29135
rect 9082 29067 9088 29132
rect 9122 29067 9128 29132
rect 9082 29060 9128 29067
rect 9082 28999 9088 29060
rect 9122 28999 9128 29060
rect 9082 28988 9128 28999
rect 9082 28931 9088 28988
rect 9122 28931 9128 28988
rect 9082 28916 9128 28931
rect 9082 28863 9088 28916
rect 9122 28863 9128 28916
rect 9082 28844 9128 28863
rect 9082 28795 9088 28844
rect 9122 28795 9128 28844
rect 9082 28772 9128 28795
rect 9082 28727 9088 28772
rect 9122 28727 9128 28772
rect 9082 28700 9128 28727
rect 9082 28659 9088 28700
rect 9122 28659 9128 28700
rect 9082 28628 9128 28659
rect 9082 28591 9088 28628
rect 9122 28591 9128 28628
rect 9082 28557 9128 28591
rect 9082 28522 9088 28557
rect 9122 28522 9128 28557
rect 9082 28489 9128 28522
rect 9082 28450 9088 28489
rect 9122 28450 9128 28489
rect 9082 28421 9128 28450
rect 9082 28378 9088 28421
rect 9122 28378 9128 28421
rect 9082 28353 9128 28378
rect 9082 28306 9088 28353
rect 9122 28306 9128 28353
rect 9082 28285 9128 28306
rect 9082 28234 9088 28285
rect 9122 28234 9128 28285
rect 9082 28217 9128 28234
rect 9082 28162 9088 28217
rect 9122 28162 9128 28217
rect 9082 28149 9128 28162
rect 9082 28090 9088 28149
rect 9122 28090 9128 28149
rect 9082 28081 9128 28090
rect 9082 28018 9088 28081
rect 9122 28018 9128 28081
rect 9082 28013 9128 28018
rect 9082 27946 9088 28013
rect 9122 27946 9128 28013
rect 9082 27945 9128 27946
rect 9082 27911 9088 27945
rect 9122 27911 9128 27945
rect 9082 27908 9128 27911
rect 9082 27843 9088 27908
rect 9122 27843 9128 27908
rect 9082 27836 9128 27843
rect 9082 27775 9088 27836
rect 9122 27775 9128 27836
rect 9082 27764 9128 27775
rect 9082 27707 9088 27764
rect 9122 27707 9128 27764
rect 9082 27692 9128 27707
rect 9082 27639 9088 27692
rect 9122 27639 9128 27692
rect 9082 27620 9128 27639
rect 9082 27571 9088 27620
rect 9122 27571 9128 27620
rect 9082 27548 9128 27571
rect 9082 27503 9088 27548
rect 9122 27503 9128 27548
rect 9082 27476 9128 27503
rect 9082 27435 9088 27476
rect 9122 27435 9128 27476
rect 9082 27404 9128 27435
rect 9082 27367 9088 27404
rect 9122 27367 9128 27404
rect 9082 27333 9128 27367
rect 9082 27298 9088 27333
rect 9122 27298 9128 27333
rect 9082 27265 9128 27298
rect 9082 27226 9088 27265
rect 9122 27226 9128 27265
rect 9082 27197 9128 27226
rect 9082 27154 9088 27197
rect 9122 27154 9128 27197
rect 9082 27129 9128 27154
rect 9082 27082 9088 27129
rect 9122 27082 9128 27129
rect 9082 27061 9128 27082
rect 9082 27010 9088 27061
rect 9122 27010 9128 27061
rect 9082 26993 9128 27010
rect 9082 26938 9088 26993
rect 9122 26938 9128 26993
rect 9082 26925 9128 26938
rect 9082 26866 9088 26925
rect 9122 26866 9128 26925
rect 9082 26857 9128 26866
rect 9082 26794 9088 26857
rect 9122 26794 9128 26857
rect 9082 26789 9128 26794
rect 9082 26722 9088 26789
rect 9122 26722 9128 26789
rect 9082 26721 9128 26722
rect 9082 26687 9088 26721
rect 9122 26687 9128 26721
rect 9082 26684 9128 26687
rect 9082 26619 9088 26684
rect 9122 26619 9128 26684
rect 9082 26612 9128 26619
rect 9082 26551 9088 26612
rect 9122 26551 9128 26612
rect 9082 26540 9128 26551
rect 9082 26483 9088 26540
rect 9122 26483 9128 26540
rect 9082 26468 9128 26483
rect 9082 26415 9088 26468
rect 9122 26415 9128 26468
rect 9082 26396 9128 26415
rect 9082 26347 9088 26396
rect 9122 26347 9128 26396
rect 9082 26324 9128 26347
rect 9082 26279 9088 26324
rect 9122 26279 9128 26324
rect 9082 26252 9128 26279
rect 9082 26211 9088 26252
rect 9122 26211 9128 26252
rect 9082 26180 9128 26211
rect 9082 26143 9088 26180
rect 9122 26143 9128 26180
rect 9082 26109 9128 26143
rect 9082 26074 9088 26109
rect 9122 26074 9128 26109
rect 9082 26041 9128 26074
rect 9082 26002 9088 26041
rect 9122 26002 9128 26041
rect 9082 25973 9128 26002
rect 9082 25930 9088 25973
rect 9122 25930 9128 25973
rect 9082 25905 9128 25930
rect 9082 25858 9088 25905
rect 9122 25858 9128 25905
rect 9082 25837 9128 25858
rect 9082 25786 9088 25837
rect 9122 25786 9128 25837
rect 9082 25769 9128 25786
rect 9082 25714 9088 25769
rect 9122 25714 9128 25769
rect 9082 25701 9128 25714
rect 9082 25642 9088 25701
rect 9122 25642 9128 25701
rect 9082 25633 9128 25642
rect 9082 25570 9088 25633
rect 9122 25570 9128 25633
rect 9082 25565 9128 25570
rect 9082 25498 9088 25565
rect 9122 25498 9128 25565
rect 9082 25497 9128 25498
rect 9082 25463 9088 25497
rect 9122 25463 9128 25497
rect 9082 25460 9128 25463
rect 9082 25395 9088 25460
rect 9122 25395 9128 25460
rect 9082 25388 9128 25395
rect 9082 25327 9088 25388
rect 9122 25327 9128 25388
rect 9082 25316 9128 25327
rect 9082 25259 9088 25316
rect 9122 25259 9128 25316
rect 9082 25244 9128 25259
rect 9082 25191 9088 25244
rect 9122 25191 9128 25244
rect 9082 25172 9128 25191
rect 9082 25123 9088 25172
rect 9122 25123 9128 25172
rect 9082 25100 9128 25123
rect 9082 25055 9088 25100
rect 9122 25055 9128 25100
rect 9082 25028 9128 25055
rect 9082 24987 9088 25028
rect 9122 24987 9128 25028
rect 9082 24956 9128 24987
rect 9082 24919 9088 24956
rect 9122 24919 9128 24956
rect 9082 24885 9128 24919
rect 9082 24850 9088 24885
rect 9122 24850 9128 24885
rect 9082 24817 9128 24850
rect 9082 24778 9088 24817
rect 9122 24778 9128 24817
rect 9082 24749 9128 24778
rect 9082 24706 9088 24749
rect 9122 24706 9128 24749
rect 9082 24681 9128 24706
rect 9082 24634 9088 24681
rect 9122 24634 9128 24681
rect 9082 24613 9128 24634
rect 9082 24562 9088 24613
rect 9122 24562 9128 24613
rect 9082 24545 9128 24562
rect 9082 24490 9088 24545
rect 9122 24490 9128 24545
rect 9082 24477 9128 24490
rect 9082 24418 9088 24477
rect 9122 24418 9128 24477
rect 9082 24409 9128 24418
rect 9082 24346 9088 24409
rect 9122 24346 9128 24409
rect 9082 24341 9128 24346
rect 9082 24274 9088 24341
rect 9122 24274 9128 24341
rect 9082 24273 9128 24274
rect 9082 24239 9088 24273
rect 9122 24239 9128 24273
rect 9082 24236 9128 24239
rect 9082 24171 9088 24236
rect 9122 24171 9128 24236
rect 9082 24164 9128 24171
rect 9082 24103 9088 24164
rect 9122 24103 9128 24164
rect 9082 24092 9128 24103
rect 9082 24035 9088 24092
rect 9122 24035 9128 24092
rect 9082 24020 9128 24035
rect 9082 23967 9088 24020
rect 9122 23967 9128 24020
rect 9082 23948 9128 23967
rect 9082 23899 9088 23948
rect 9122 23899 9128 23948
rect 9082 23876 9128 23899
rect 9082 23831 9088 23876
rect 9122 23831 9128 23876
rect 9082 23804 9128 23831
rect 9082 23763 9088 23804
rect 9122 23763 9128 23804
rect 9082 23732 9128 23763
rect 9082 23695 9088 23732
rect 9122 23695 9128 23732
rect 9082 23661 9128 23695
rect 9082 23626 9088 23661
rect 9122 23626 9128 23661
rect 9082 23593 9128 23626
rect 9082 23554 9088 23593
rect 9122 23554 9128 23593
rect 9082 23525 9128 23554
rect 9082 23482 9088 23525
rect 9122 23482 9128 23525
rect 9082 23457 9128 23482
rect 9082 23410 9088 23457
rect 9122 23410 9128 23457
rect 9082 23389 9128 23410
rect 9082 23338 9088 23389
rect 9122 23338 9128 23389
rect 9082 23321 9128 23338
rect 9082 23266 9088 23321
rect 9122 23266 9128 23321
rect 9082 23253 9128 23266
rect 9082 23194 9088 23253
rect 9122 23194 9128 23253
rect 9082 23185 9128 23194
rect 9082 23122 9088 23185
rect 9122 23122 9128 23185
rect 9082 23117 9128 23122
rect 9082 23050 9088 23117
rect 9122 23050 9128 23117
rect 9082 23049 9128 23050
rect 9082 23015 9088 23049
rect 9122 23015 9128 23049
rect 9082 23012 9128 23015
rect 9082 22947 9088 23012
rect 9122 22947 9128 23012
rect 9082 22940 9128 22947
rect 9082 22879 9088 22940
rect 9122 22879 9128 22940
rect 9082 22868 9128 22879
rect 9082 22811 9088 22868
rect 9122 22811 9128 22868
rect 9082 22796 9128 22811
rect 9082 22743 9088 22796
rect 9122 22743 9128 22796
rect 9082 22724 9128 22743
rect 9082 22675 9088 22724
rect 9122 22675 9128 22724
rect 9082 22652 9128 22675
rect 9082 22607 9088 22652
rect 9122 22607 9128 22652
rect 9082 22580 9128 22607
rect 9082 22539 9088 22580
rect 9122 22539 9128 22580
rect 9082 22508 9128 22539
rect 9082 22471 9088 22508
rect 9122 22471 9128 22508
rect 9082 22437 9128 22471
rect 9082 22402 9088 22437
rect 9122 22402 9128 22437
rect 9082 22369 9128 22402
rect 9082 22330 9088 22369
rect 9122 22330 9128 22369
rect 9082 22301 9128 22330
rect 9082 22258 9088 22301
rect 9122 22258 9128 22301
rect 9082 22233 9128 22258
rect 9082 22186 9088 22233
rect 9122 22186 9128 22233
rect 9082 22165 9128 22186
rect 9082 22114 9088 22165
rect 9122 22114 9128 22165
rect 9082 22097 9128 22114
rect 9082 22042 9088 22097
rect 9122 22042 9128 22097
rect 9082 22029 9128 22042
rect 9082 21970 9088 22029
rect 9122 21970 9128 22029
rect 9082 21961 9128 21970
rect 9082 21898 9088 21961
rect 9122 21898 9128 21961
rect 9082 21893 9128 21898
rect 9082 21826 9088 21893
rect 9122 21826 9128 21893
rect 9082 21825 9128 21826
rect 9082 21791 9088 21825
rect 9122 21791 9128 21825
rect 9082 21788 9128 21791
rect 9082 21723 9088 21788
rect 9122 21723 9128 21788
rect 9082 21716 9128 21723
rect 9082 21655 9088 21716
rect 9122 21655 9128 21716
rect 9082 21644 9128 21655
rect 9082 21587 9088 21644
rect 9122 21587 9128 21644
rect 9082 21572 9128 21587
rect 9082 21519 9088 21572
rect 9122 21519 9128 21572
rect 9082 21500 9128 21519
rect 9082 21451 9088 21500
rect 9122 21451 9128 21500
rect 9082 21428 9128 21451
rect 9082 21383 9088 21428
rect 9122 21383 9128 21428
rect 9082 21356 9128 21383
rect 9082 21315 9088 21356
rect 9122 21315 9128 21356
rect 9082 21284 9128 21315
rect 9082 21247 9088 21284
rect 9122 21247 9128 21284
rect 9082 21213 9128 21247
rect 9082 21178 9088 21213
rect 9122 21178 9128 21213
rect 9082 21145 9128 21178
rect 9082 21106 9088 21145
rect 9122 21106 9128 21145
rect 9082 21077 9128 21106
rect 9082 21034 9088 21077
rect 9122 21034 9128 21077
rect 9082 21009 9128 21034
rect 9082 20962 9088 21009
rect 9122 20962 9128 21009
rect 9082 20941 9128 20962
rect 9082 20890 9088 20941
rect 9122 20890 9128 20941
rect 9082 20873 9128 20890
rect 9082 20818 9088 20873
rect 9122 20818 9128 20873
rect 9082 20805 9128 20818
rect 9082 20746 9088 20805
rect 9122 20746 9128 20805
rect 9082 20737 9128 20746
rect 9082 20674 9088 20737
rect 9122 20674 9128 20737
rect 9082 20669 9128 20674
rect 9082 20602 9088 20669
rect 9122 20602 9128 20669
rect 9082 20601 9128 20602
rect 9082 20567 9088 20601
rect 9122 20567 9128 20601
rect 9082 20564 9128 20567
rect 9082 20499 9088 20564
rect 9122 20499 9128 20564
rect 9082 20492 9128 20499
rect 9082 20431 9088 20492
rect 9122 20431 9128 20492
rect 9082 20420 9128 20431
rect 9082 20363 9088 20420
rect 9122 20363 9128 20420
rect 9082 20348 9128 20363
rect 9082 20295 9088 20348
rect 9122 20295 9128 20348
rect 9082 20276 9128 20295
rect 9082 20227 9088 20276
rect 9122 20227 9128 20276
rect 9082 20204 9128 20227
rect 9082 20159 9088 20204
rect 9122 20159 9128 20204
rect 9082 20132 9128 20159
rect 9082 20091 9088 20132
rect 9122 20091 9128 20132
rect 9082 20060 9128 20091
rect 9082 20023 9088 20060
rect 9122 20023 9128 20060
rect 9082 19989 9128 20023
rect 9082 19954 9088 19989
rect 9122 19954 9128 19989
rect 9082 19921 9128 19954
rect 9082 19882 9088 19921
rect 9122 19882 9128 19921
rect 9082 19853 9128 19882
rect 9082 19810 9088 19853
rect 9122 19810 9128 19853
rect 9082 19785 9128 19810
rect 9082 19738 9088 19785
rect 9122 19738 9128 19785
rect 9082 19717 9128 19738
rect 9082 19666 9088 19717
rect 9122 19666 9128 19717
rect 9082 19649 9128 19666
rect 9082 19594 9088 19649
rect 9122 19594 9128 19649
rect 9082 19581 9128 19594
rect 9082 19522 9088 19581
rect 9122 19522 9128 19581
rect 9082 19513 9128 19522
rect 9082 19450 9088 19513
rect 9122 19450 9128 19513
rect 9082 19445 9128 19450
rect 9082 19378 9088 19445
rect 9122 19378 9128 19445
rect 9082 19377 9128 19378
rect 9082 19343 9088 19377
rect 9122 19343 9128 19377
rect 9082 19340 9128 19343
rect 9082 19275 9088 19340
rect 9122 19275 9128 19340
rect 9082 19268 9128 19275
rect 9082 19207 9088 19268
rect 9122 19207 9128 19268
rect 9082 19196 9128 19207
rect 9082 19139 9088 19196
rect 9122 19139 9128 19196
rect 9082 19124 9128 19139
rect 9082 19071 9088 19124
rect 9122 19071 9128 19124
rect 9082 19052 9128 19071
rect 9082 19003 9088 19052
rect 9122 19003 9128 19052
rect 9082 18980 9128 19003
rect 9082 18935 9088 18980
rect 9122 18935 9128 18980
rect 9082 18908 9128 18935
rect 9082 18867 9088 18908
rect 9122 18867 9128 18908
rect 9082 18836 9128 18867
rect 9082 18799 9088 18836
rect 9122 18799 9128 18836
rect 9082 18765 9128 18799
rect 9082 18730 9088 18765
rect 9122 18730 9128 18765
rect 9082 18697 9128 18730
rect 9082 18658 9088 18697
rect 9122 18658 9128 18697
rect 9082 18629 9128 18658
rect 9082 18586 9088 18629
rect 9122 18586 9128 18629
rect 9082 18561 9128 18586
rect 9082 18514 9088 18561
rect 9122 18514 9128 18561
rect 9082 18493 9128 18514
rect 9082 18442 9088 18493
rect 9122 18442 9128 18493
rect 9082 18425 9128 18442
rect 9082 18370 9088 18425
rect 9122 18370 9128 18425
rect 9082 18357 9128 18370
rect 9082 18298 9088 18357
rect 9122 18298 9128 18357
rect 9082 18289 9128 18298
rect 9082 18226 9088 18289
rect 9122 18226 9128 18289
rect 9082 18221 9128 18226
rect 9082 18154 9088 18221
rect 9122 18154 9128 18221
rect 9082 18153 9128 18154
rect 9082 18119 9088 18153
rect 9122 18119 9128 18153
rect 9082 18116 9128 18119
rect 9082 18051 9088 18116
rect 9122 18051 9128 18116
rect 9082 18044 9128 18051
rect 9082 17983 9088 18044
rect 9122 17983 9128 18044
rect 9082 17972 9128 17983
rect 9082 17915 9088 17972
rect 9122 17915 9128 17972
rect 9082 17900 9128 17915
rect 9082 17847 9088 17900
rect 9122 17847 9128 17900
rect 9082 17828 9128 17847
rect 9082 17779 9088 17828
rect 9122 17779 9128 17828
rect 9082 17756 9128 17779
rect 9082 17711 9088 17756
rect 9122 17711 9128 17756
rect 9082 17684 9128 17711
rect 9082 17643 9088 17684
rect 9122 17643 9128 17684
rect 9082 17612 9128 17643
rect 9082 17575 9088 17612
rect 9122 17575 9128 17612
rect 9082 17541 9128 17575
rect 9082 17506 9088 17541
rect 9122 17506 9128 17541
rect 9082 17473 9128 17506
rect 9082 17434 9088 17473
rect 9122 17434 9128 17473
rect 9082 17405 9128 17434
rect 9082 17362 9088 17405
rect 9122 17362 9128 17405
rect 9082 17337 9128 17362
rect 9082 17290 9088 17337
rect 9122 17290 9128 17337
rect 9082 17269 9128 17290
rect 9082 17218 9088 17269
rect 9122 17218 9128 17269
rect 9082 17201 9128 17218
rect 9082 17146 9088 17201
rect 9122 17146 9128 17201
rect 9082 17133 9128 17146
rect 9082 17074 9088 17133
rect 9122 17074 9128 17133
rect 9082 17065 9128 17074
rect 9082 17002 9088 17065
rect 9122 17002 9128 17065
rect 9082 16997 9128 17002
rect 9082 16930 9088 16997
rect 9122 16930 9128 16997
rect 9082 16929 9128 16930
rect 9082 16895 9088 16929
rect 9122 16895 9128 16929
rect 9082 16892 9128 16895
rect 9082 16827 9088 16892
rect 9122 16827 9128 16892
rect 9082 16820 9128 16827
rect 9082 16759 9088 16820
rect 9122 16759 9128 16820
rect 9082 16748 9128 16759
rect 9082 16691 9088 16748
rect 9122 16691 9128 16748
rect 9082 16676 9128 16691
rect 9082 16623 9088 16676
rect 9122 16623 9128 16676
rect 9082 16604 9128 16623
rect 9082 16555 9088 16604
rect 9122 16555 9128 16604
rect 9082 16532 9128 16555
rect 9082 16487 9088 16532
rect 9122 16487 9128 16532
rect 9082 16460 9128 16487
rect 9082 16419 9088 16460
rect 9122 16419 9128 16460
rect 9082 16388 9128 16419
rect 9082 16351 9088 16388
rect 9122 16351 9128 16388
rect 9082 16317 9128 16351
rect 9082 16282 9088 16317
rect 9122 16282 9128 16317
rect 9082 16249 9128 16282
rect 9082 16210 9088 16249
rect 9122 16210 9128 16249
rect 9082 16181 9128 16210
rect 9082 16138 9088 16181
rect 9122 16138 9128 16181
rect 9082 16113 9128 16138
rect 9082 16066 9088 16113
rect 9122 16066 9128 16113
rect 9082 16045 9128 16066
rect 9082 15994 9088 16045
rect 9122 15994 9128 16045
rect 9082 15977 9128 15994
rect 9082 15922 9088 15977
rect 9122 15922 9128 15977
rect 9082 15909 9128 15922
rect 9082 15850 9088 15909
rect 9122 15850 9128 15909
rect 9082 15841 9128 15850
rect 9082 15778 9088 15841
rect 9122 15778 9128 15841
rect 9082 15773 9128 15778
rect 9082 15706 9088 15773
rect 9122 15706 9128 15773
rect 9082 15705 9128 15706
rect 9082 15671 9088 15705
rect 9122 15671 9128 15705
rect 9082 15668 9128 15671
rect 9082 15603 9088 15668
rect 9122 15603 9128 15668
rect 9082 15596 9128 15603
rect 9082 15535 9088 15596
rect 9122 15535 9128 15596
rect 9082 15524 9128 15535
rect 9082 15467 9088 15524
rect 9122 15467 9128 15524
rect 9082 15452 9128 15467
rect 9082 15399 9088 15452
rect 9122 15399 9128 15452
rect 9082 15380 9128 15399
rect 9082 15331 9088 15380
rect 9122 15331 9128 15380
rect 9082 15308 9128 15331
rect 9082 15263 9088 15308
rect 9122 15263 9128 15308
rect 9082 15236 9128 15263
rect 9082 15195 9088 15236
rect 9122 15195 9128 15236
rect 9082 15164 9128 15195
rect 9082 15127 9088 15164
rect 9122 15127 9128 15164
rect 9082 15093 9128 15127
rect 9082 15058 9088 15093
rect 9122 15058 9128 15093
rect 9082 15025 9128 15058
rect 9082 14986 9088 15025
rect 9122 14986 9128 15025
rect 9082 14957 9128 14986
rect 9082 14914 9088 14957
rect 9122 14914 9128 14957
rect 9082 14889 9128 14914
rect 9082 14842 9088 14889
rect 9122 14842 9128 14889
rect 9082 14821 9128 14842
rect 9082 14770 9088 14821
rect 9122 14770 9128 14821
rect 9082 14753 9128 14770
rect 9082 14698 9088 14753
rect 9122 14698 9128 14753
rect 9082 14685 9128 14698
rect 9082 14626 9088 14685
rect 9122 14626 9128 14685
rect 9082 14617 9128 14626
rect 9082 14554 9088 14617
rect 9122 14554 9128 14617
rect 9082 14549 9128 14554
rect 9082 14482 9088 14549
rect 9122 14482 9128 14549
rect 9082 14481 9128 14482
rect 9082 14447 9088 14481
rect 9122 14447 9128 14481
rect 9082 14444 9128 14447
rect 9082 14379 9088 14444
rect 9122 14379 9128 14444
rect 9082 14372 9128 14379
rect 9082 14311 9088 14372
rect 9122 14311 9128 14372
rect 9082 14300 9128 14311
rect 9082 14243 9088 14300
rect 9122 14243 9128 14300
rect 9082 14228 9128 14243
rect 9082 14175 9088 14228
rect 9122 14175 9128 14228
rect 9082 14156 9128 14175
rect 9082 14107 9088 14156
rect 9122 14107 9128 14156
rect 9082 14084 9128 14107
rect 9082 14039 9088 14084
rect 9122 14039 9128 14084
rect 9082 14012 9128 14039
rect 9082 13971 9088 14012
rect 9122 13971 9128 14012
rect 9082 13940 9128 13971
rect 9082 13903 9088 13940
rect 9122 13903 9128 13940
rect 9082 13869 9128 13903
rect 9082 13834 9088 13869
rect 9122 13834 9128 13869
rect 9082 13801 9128 13834
rect 9082 13762 9088 13801
rect 9122 13762 9128 13801
rect 9082 13733 9128 13762
rect 9082 13690 9088 13733
rect 9122 13690 9128 13733
rect 9082 13665 9128 13690
rect 9082 13618 9088 13665
rect 9122 13618 9128 13665
rect 9082 13597 9128 13618
rect 9082 13546 9088 13597
rect 9122 13546 9128 13597
rect 9082 13529 9128 13546
rect 9082 13474 9088 13529
rect 9122 13474 9128 13529
rect 9082 13461 9128 13474
rect 9082 13402 9088 13461
rect 9122 13402 9128 13461
rect 9082 13393 9128 13402
rect 9082 13330 9088 13393
rect 9122 13330 9128 13393
rect 9082 13325 9128 13330
rect 9082 13258 9088 13325
rect 9122 13258 9128 13325
rect 9082 13257 9128 13258
rect 9082 13223 9088 13257
rect 9122 13223 9128 13257
rect 9082 13220 9128 13223
rect 9082 13155 9088 13220
rect 9122 13155 9128 13220
rect 9082 13148 9128 13155
rect 9082 13087 9088 13148
rect 9122 13087 9128 13148
rect 9082 13076 9128 13087
rect 9082 13019 9088 13076
rect 9122 13019 9128 13076
rect 9082 13004 9128 13019
rect 9082 12951 9088 13004
rect 9122 12951 9128 13004
rect 9082 12932 9128 12951
rect 9082 12883 9088 12932
rect 9122 12883 9128 12932
rect 9082 12860 9128 12883
rect 9082 12815 9088 12860
rect 9122 12815 9128 12860
rect 9082 12788 9128 12815
rect 9082 12747 9088 12788
rect 9122 12747 9128 12788
rect 9082 12716 9128 12747
rect 9082 12679 9088 12716
rect 9122 12679 9128 12716
rect 9082 12645 9128 12679
rect 9082 12610 9088 12645
rect 9122 12610 9128 12645
rect 9082 12577 9128 12610
rect 9082 12538 9088 12577
rect 9122 12538 9128 12577
rect 9082 12509 9128 12538
rect 9082 12466 9088 12509
rect 9122 12466 9128 12509
rect 9082 12441 9128 12466
rect 9082 12394 9088 12441
rect 9122 12394 9128 12441
rect 9082 12373 9128 12394
rect 9082 12322 9088 12373
rect 9122 12322 9128 12373
rect 9082 12305 9128 12322
rect 9082 12250 9088 12305
rect 9122 12250 9128 12305
rect 9082 12237 9128 12250
rect 9082 12178 9088 12237
rect 9122 12178 9128 12237
rect 9082 12169 9128 12178
rect 9082 12106 9088 12169
rect 9122 12106 9128 12169
rect 9082 12101 9128 12106
rect 9082 12034 9088 12101
rect 9122 12034 9128 12101
rect 9082 12033 9128 12034
rect 9082 11999 9088 12033
rect 9122 11999 9128 12033
rect 9082 11996 9128 11999
rect 9082 11931 9088 11996
rect 9122 11931 9128 11996
rect 9082 11924 9128 11931
rect 9082 11863 9088 11924
rect 9122 11863 9128 11924
rect 9082 11852 9128 11863
rect 9082 11795 9088 11852
rect 9122 11795 9128 11852
rect 9082 11780 9128 11795
rect 9082 11727 9088 11780
rect 9122 11727 9128 11780
rect 9082 11708 9128 11727
rect 9082 11659 9088 11708
rect 9122 11659 9128 11708
rect 9082 11636 9128 11659
rect 9082 11591 9088 11636
rect 9122 11591 9128 11636
rect 9082 11564 9128 11591
rect 9082 11523 9088 11564
rect 9122 11523 9128 11564
rect 9082 11492 9128 11523
rect 9082 11455 9088 11492
rect 9122 11455 9128 11492
rect 9082 11421 9128 11455
rect 9082 11386 9088 11421
rect 9122 11386 9128 11421
rect 9082 11353 9128 11386
rect 9082 11314 9088 11353
rect 9122 11314 9128 11353
rect 9082 11285 9128 11314
rect 9082 11242 9088 11285
rect 9122 11242 9128 11285
rect 9082 11217 9128 11242
rect 9082 11170 9088 11217
rect 9122 11170 9128 11217
rect 9082 11149 9128 11170
rect 9082 11098 9088 11149
rect 9122 11098 9128 11149
rect 9082 11081 9128 11098
rect 9082 11026 9088 11081
rect 9122 11026 9128 11081
rect 9082 11013 9128 11026
rect 9082 10954 9088 11013
rect 9122 10954 9128 11013
rect 9082 10945 9128 10954
rect 9082 10882 9088 10945
rect 9122 10882 9128 10945
rect 9082 10877 9128 10882
rect 9082 10810 9088 10877
rect 9122 10810 9128 10877
rect 9082 10809 9128 10810
rect 9082 10775 9088 10809
rect 9122 10775 9128 10809
rect 9082 10772 9128 10775
rect 9082 10707 9088 10772
rect 9122 10707 9128 10772
rect 9082 10700 9128 10707
rect 9082 10639 9088 10700
rect 9122 10639 9128 10700
rect 9082 10628 9128 10639
rect 9082 10571 9088 10628
rect 9122 10571 9128 10628
rect 9082 10556 9128 10571
rect 9082 10503 9088 10556
rect 9122 10503 9128 10556
rect 9082 10484 9128 10503
rect 9082 10435 9088 10484
rect 9122 10435 9128 10484
rect 9082 10412 9128 10435
rect 9082 10367 9088 10412
rect 9122 10367 9128 10412
rect 9082 10340 9128 10367
rect 9082 10299 9088 10340
rect 9122 10299 9128 10340
rect 9082 10268 9128 10299
rect 9082 10231 9088 10268
rect 9122 10231 9128 10268
rect 9082 10197 9128 10231
rect 9082 10162 9088 10197
rect 9122 10162 9128 10197
rect 9082 10129 9128 10162
rect 9082 10090 9088 10129
rect 9122 10090 9128 10129
rect 9082 10061 9128 10090
rect 9082 10018 9088 10061
rect 9122 10018 9128 10061
rect 9082 9993 9128 10018
rect 9082 9946 9088 9993
rect 9122 9946 9128 9993
rect 9082 9925 9128 9946
rect 9082 9874 9088 9925
rect 9122 9874 9128 9925
rect 9082 9857 9128 9874
rect 9082 9802 9088 9857
rect 9122 9802 9128 9857
rect 9082 9789 9128 9802
rect 9082 9730 9088 9789
rect 9122 9730 9128 9789
rect 9082 9721 9128 9730
rect 9082 9658 9088 9721
rect 9122 9658 9128 9721
rect 9082 9653 9128 9658
rect 9082 9586 9088 9653
rect 9122 9586 9128 9653
rect 9082 9585 9128 9586
rect 9082 9551 9088 9585
rect 9122 9551 9128 9585
rect 9082 9548 9128 9551
rect 9082 9483 9088 9548
rect 9122 9483 9128 9548
rect 9082 9476 9128 9483
rect 9082 9415 9088 9476
rect 9122 9415 9128 9476
rect 9082 9404 9128 9415
rect 9082 9347 9088 9404
rect 9122 9347 9128 9404
rect 9082 9332 9128 9347
rect 9082 9279 9088 9332
rect 9122 9279 9128 9332
rect 9082 9260 9128 9279
rect 9082 9211 9088 9260
rect 9122 9211 9128 9260
rect 9082 9188 9128 9211
rect 9082 9143 9088 9188
rect 9122 9143 9128 9188
rect 9082 9116 9128 9143
rect 9082 9075 9088 9116
rect 9122 9075 9128 9116
rect 9082 9044 9128 9075
rect 9082 9007 9088 9044
rect 9122 9007 9128 9044
rect 9082 8973 9128 9007
rect 9082 8938 9088 8973
rect 9122 8938 9128 8973
rect 9082 8905 9128 8938
rect 9082 8866 9088 8905
rect 9122 8866 9128 8905
rect 9082 8837 9128 8866
rect 9082 8794 9088 8837
rect 9122 8794 9128 8837
rect 9082 8769 9128 8794
rect 9082 8722 9088 8769
rect 9122 8722 9128 8769
rect 9082 8701 9128 8722
rect 9082 8650 9088 8701
rect 9122 8650 9128 8701
rect 9082 8633 9128 8650
rect 9082 8578 9088 8633
rect 9122 8578 9128 8633
rect 9082 8565 9128 8578
rect 9082 8506 9088 8565
rect 9122 8506 9128 8565
rect 9082 8497 9128 8506
rect 9082 8434 9088 8497
rect 9122 8434 9128 8497
rect 9082 8429 9128 8434
rect 9082 8362 9088 8429
rect 9122 8362 9128 8429
rect 9082 8361 9128 8362
rect 9082 8327 9088 8361
rect 9122 8327 9128 8361
rect 9082 8324 9128 8327
rect 9082 8259 9088 8324
rect 9122 8259 9128 8324
rect 9082 8252 9128 8259
rect 9082 8191 9088 8252
rect 9122 8191 9128 8252
rect 9082 8180 9128 8191
rect 9082 8123 9088 8180
rect 9122 8123 9128 8180
rect 9082 8108 9128 8123
rect 9082 8055 9088 8108
rect 9122 8055 9128 8108
rect 9082 8036 9128 8055
rect 9082 7987 9088 8036
rect 9122 7987 9128 8036
rect 9082 7964 9128 7987
rect 9082 7919 9088 7964
rect 9122 7919 9128 7964
rect 9082 7892 9128 7919
rect 9082 7851 9088 7892
rect 9122 7851 9128 7892
rect 9082 7820 9128 7851
rect 9082 7783 9088 7820
rect 9122 7783 9128 7820
rect 9082 7749 9128 7783
rect 9082 7714 9088 7749
rect 9122 7714 9128 7749
rect 9082 7681 9128 7714
rect 9082 7642 9088 7681
rect 9122 7642 9128 7681
rect 9082 7613 9128 7642
rect 9082 7570 9088 7613
rect 9122 7570 9128 7613
rect 9082 7545 9128 7570
rect 9082 7498 9088 7545
rect 9122 7498 9128 7545
rect 9082 7477 9128 7498
rect 9082 7426 9088 7477
rect 9122 7426 9128 7477
rect 9082 7409 9128 7426
rect 9082 7354 9088 7409
rect 9122 7354 9128 7409
rect 9082 7341 9128 7354
rect 9082 7282 9088 7341
rect 9122 7282 9128 7341
rect 9082 7273 9128 7282
rect 9082 7210 9088 7273
rect 9122 7210 9128 7273
rect 9082 7205 9128 7210
rect 9082 7138 9088 7205
rect 9122 7138 9128 7205
rect 9082 7137 9128 7138
rect 9082 7103 9088 7137
rect 9122 7103 9128 7137
rect 9082 7100 9128 7103
rect 9082 7035 9088 7100
rect 9122 7035 9128 7100
rect 9082 7028 9128 7035
rect 9082 6967 9088 7028
rect 9122 6967 9128 7028
rect 9082 6956 9128 6967
rect 9082 6899 9088 6956
rect 9122 6899 9128 6956
rect 9082 6884 9128 6899
rect 9082 6831 9088 6884
rect 9122 6831 9128 6884
rect 9082 6812 9128 6831
rect 9082 6763 9088 6812
rect 9122 6763 9128 6812
rect 9082 6740 9128 6763
rect 9082 6695 9088 6740
rect 9122 6695 9128 6740
rect 9082 6668 9128 6695
rect 9082 6627 9088 6668
rect 9122 6627 9128 6668
rect 9082 6596 9128 6627
rect 9082 6559 9088 6596
rect 9122 6559 9128 6596
rect 9082 6525 9128 6559
rect 9082 6490 9088 6525
rect 9122 6490 9128 6525
rect 9082 6457 9128 6490
rect 9082 6418 9088 6457
rect 9122 6418 9128 6457
rect 9082 6389 9128 6418
rect 9082 6346 9088 6389
rect 9122 6346 9128 6389
rect 9082 6321 9128 6346
rect 9082 6274 9088 6321
rect 9122 6274 9128 6321
rect 9082 6253 9128 6274
rect 9082 6202 9088 6253
rect 9122 6202 9128 6253
rect 9082 6185 9128 6202
rect 9082 6130 9088 6185
rect 9122 6130 9128 6185
rect 9082 6117 9128 6130
rect 9082 6058 9088 6117
rect 9122 6058 9128 6117
rect 9082 6049 9128 6058
rect 9082 5986 9088 6049
rect 9122 5986 9128 6049
rect 9082 5981 9128 5986
rect 9082 5914 9088 5981
rect 9122 5914 9128 5981
rect 9082 5913 9128 5914
rect 9082 5879 9088 5913
rect 9122 5879 9128 5913
rect 9082 5876 9128 5879
rect 9082 5811 9088 5876
rect 9122 5811 9128 5876
rect 9082 5804 9128 5811
rect 9082 5743 9088 5804
rect 9122 5743 9128 5804
rect 9082 5732 9128 5743
rect 9082 5675 9088 5732
rect 9122 5675 9128 5732
rect 9082 5660 9128 5675
rect 9082 5607 9088 5660
rect 9122 5607 9128 5660
rect 9082 5588 9128 5607
rect 9082 5539 9088 5588
rect 9122 5539 9128 5588
rect 9082 5516 9128 5539
rect 9082 5471 9088 5516
rect 9122 5471 9128 5516
rect 9082 5444 9128 5471
rect 9082 5403 9088 5444
rect 9122 5403 9128 5444
rect 9082 5372 9128 5403
rect 9082 5335 9088 5372
rect 9122 5335 9128 5372
rect 9082 5301 9128 5335
rect 9082 5266 9088 5301
rect 9122 5266 9128 5301
rect 9082 5233 9128 5266
rect 9082 5194 9088 5233
rect 9122 5194 9128 5233
rect 9082 5165 9128 5194
rect 9082 5122 9088 5165
rect 9122 5122 9128 5165
rect 9082 5097 9128 5122
rect 9082 5050 9088 5097
rect 9122 5050 9128 5097
rect 9082 5029 9128 5050
rect 9082 4978 9088 5029
rect 9122 4978 9128 5029
rect 9082 4961 9128 4978
rect 9082 4906 9088 4961
rect 9122 4906 9128 4961
rect 9082 4893 9128 4906
rect 9082 4834 9088 4893
rect 9122 4834 9128 4893
rect 9082 4825 9128 4834
rect 9082 4762 9088 4825
rect 9122 4762 9128 4825
rect 9082 4757 9128 4762
rect 9082 4690 9088 4757
rect 9122 4690 9128 4757
rect 9082 4689 9128 4690
rect 9082 4655 9088 4689
rect 9122 4655 9128 4689
rect 9082 4652 9128 4655
rect 9082 4587 9088 4652
rect 9122 4587 9128 4652
rect 9082 4580 9128 4587
rect 9082 4519 9088 4580
rect 9122 4519 9128 4580
rect 9082 4508 9128 4519
rect 9082 4451 9088 4508
rect 9122 4451 9128 4508
rect 9082 4436 9128 4451
rect 9082 4383 9088 4436
rect 9122 4383 9128 4436
rect 9082 4364 9128 4383
rect 9082 4315 9088 4364
rect 9122 4315 9128 4364
rect 9082 4292 9128 4315
rect 9082 4247 9088 4292
rect 9122 4247 9128 4292
rect 9082 4220 9128 4247
rect 9082 4179 9088 4220
rect 9122 4179 9128 4220
rect 9082 4148 9128 4179
rect 9082 4111 9088 4148
rect 9122 4111 9128 4148
rect 9082 4077 9128 4111
rect 9082 4042 9088 4077
rect 9122 4042 9128 4077
rect 9082 4009 9128 4042
rect 9082 3970 9088 4009
rect 9122 3970 9128 4009
rect 9082 3941 9128 3970
rect 9082 3898 9088 3941
rect 9122 3898 9128 3941
rect 9082 3873 9128 3898
rect 9082 3826 9088 3873
rect 9122 3826 9128 3873
rect 9082 3805 9128 3826
rect 9082 3754 9088 3805
rect 9122 3754 9128 3805
rect 9082 3737 9128 3754
rect 9082 3682 9088 3737
rect 9122 3682 9128 3737
rect 9082 3669 9128 3682
rect 9082 3610 9088 3669
rect 9122 3610 9128 3669
rect 9082 3601 9128 3610
rect 9082 3538 9088 3601
rect 9122 3538 9128 3601
rect 9082 3533 9128 3538
rect 9082 3466 9088 3533
rect 9122 3466 9128 3533
rect 10220 38684 10266 38716
rect 10220 38650 10226 38684
rect 10260 38650 10266 38684
rect 10220 38641 10266 38650
rect 10220 38577 10226 38641
rect 10260 38577 10266 38641
rect 10220 38573 10266 38577
rect 10220 38539 10226 38573
rect 10260 38539 10266 38573
rect 10220 38538 10266 38539
rect 10220 38471 10226 38538
rect 10260 38471 10266 38538
rect 10220 38465 10266 38471
rect 10220 38403 10226 38465
rect 10260 38403 10266 38465
rect 10220 38392 10266 38403
rect 10220 38335 10226 38392
rect 10260 38335 10266 38392
rect 10220 38319 10266 38335
rect 10220 38267 10226 38319
rect 10260 38267 10266 38319
rect 10220 38246 10266 38267
rect 10220 38199 10226 38246
rect 10260 38199 10266 38246
rect 10220 38173 10266 38199
rect 10220 38131 10226 38173
rect 10260 38131 10266 38173
rect 10220 38100 10266 38131
rect 10220 38063 10226 38100
rect 10260 38063 10266 38100
rect 10220 38029 10266 38063
rect 10220 37993 10226 38029
rect 10260 37993 10266 38029
rect 10220 37961 10266 37993
rect 10220 37920 10226 37961
rect 10260 37920 10266 37961
rect 10220 37893 10266 37920
rect 10220 37847 10226 37893
rect 10260 37847 10266 37893
rect 10220 37825 10266 37847
rect 10220 37774 10226 37825
rect 10260 37774 10266 37825
rect 10220 37757 10266 37774
rect 10220 37701 10226 37757
rect 10260 37701 10266 37757
rect 10220 37689 10266 37701
rect 10220 37628 10226 37689
rect 10260 37628 10266 37689
rect 10220 37621 10266 37628
rect 10220 37555 10226 37621
rect 10260 37555 10266 37621
rect 10220 37553 10266 37555
rect 10220 37519 10226 37553
rect 10260 37519 10266 37553
rect 10220 37516 10266 37519
rect 10220 37451 10226 37516
rect 10260 37451 10266 37516
rect 10220 37443 10266 37451
rect 10220 37383 10226 37443
rect 10260 37383 10266 37443
rect 10220 37370 10266 37383
rect 10220 37315 10226 37370
rect 10260 37315 10266 37370
rect 10220 37297 10266 37315
rect 10220 37247 10226 37297
rect 10260 37247 10266 37297
rect 10220 37224 10266 37247
rect 10220 37179 10226 37224
rect 10260 37179 10266 37224
rect 10220 37151 10266 37179
rect 10220 37111 10226 37151
rect 10260 37111 10266 37151
rect 10220 37078 10266 37111
rect 10220 37043 10226 37078
rect 10260 37043 10266 37078
rect 10220 37009 10266 37043
rect 10220 36971 10226 37009
rect 10260 36971 10266 37009
rect 10220 36941 10266 36971
rect 10220 36898 10226 36941
rect 10260 36898 10266 36941
rect 10220 36873 10266 36898
rect 10220 36825 10226 36873
rect 10260 36825 10266 36873
rect 10220 36805 10266 36825
rect 10220 36752 10226 36805
rect 10260 36752 10266 36805
rect 10220 36737 10266 36752
rect 10220 36679 10226 36737
rect 10260 36679 10266 36737
rect 10220 36669 10266 36679
rect 10220 36606 10226 36669
rect 10260 36606 10266 36669
rect 10220 36601 10266 36606
rect 10220 36499 10226 36601
rect 10260 36499 10266 36601
rect 10220 36494 10266 36499
rect 10220 36431 10226 36494
rect 10260 36431 10266 36494
rect 10220 36421 10266 36431
rect 10220 36363 10226 36421
rect 10260 36363 10266 36421
rect 10220 36348 10266 36363
rect 10220 36295 10226 36348
rect 10260 36295 10266 36348
rect 10220 36275 10266 36295
rect 10220 36227 10226 36275
rect 10260 36227 10266 36275
rect 10220 36202 10266 36227
rect 10220 36159 10226 36202
rect 10260 36159 10266 36202
rect 10220 36129 10266 36159
rect 10220 36091 10226 36129
rect 10260 36091 10266 36129
rect 10220 36057 10266 36091
rect 10220 36022 10226 36057
rect 10260 36022 10266 36057
rect 10220 35989 10266 36022
rect 10220 35949 10226 35989
rect 10260 35949 10266 35989
rect 10220 35921 10266 35949
rect 10220 35876 10226 35921
rect 10260 35876 10266 35921
rect 10220 35853 10266 35876
rect 10220 35803 10226 35853
rect 10260 35803 10266 35853
rect 10220 35785 10266 35803
rect 10220 35730 10226 35785
rect 10260 35730 10266 35785
rect 10220 35717 10266 35730
rect 10220 35657 10226 35717
rect 10260 35657 10266 35717
rect 10220 35649 10266 35657
rect 10220 35584 10226 35649
rect 10260 35584 10266 35649
rect 10220 35581 10266 35584
rect 10220 35547 10226 35581
rect 10260 35547 10266 35581
rect 10220 35545 10266 35547
rect 10220 35479 10226 35545
rect 10260 35479 10266 35545
rect 10220 35472 10266 35479
rect 10220 35411 10226 35472
rect 10260 35411 10266 35472
rect 10220 35399 10266 35411
rect 10220 35343 10226 35399
rect 10260 35343 10266 35399
rect 10220 35326 10266 35343
rect 10220 35275 10226 35326
rect 10260 35275 10266 35326
rect 10220 35253 10266 35275
rect 10220 35207 10226 35253
rect 10260 35207 10266 35253
rect 10220 35180 10266 35207
rect 10220 35139 10226 35180
rect 10260 35139 10266 35180
rect 10220 35108 10266 35139
rect 10220 35071 10226 35108
rect 10260 35071 10266 35108
rect 10220 35037 10266 35071
rect 10220 35002 10226 35037
rect 10260 35002 10266 35037
rect 10220 34969 10266 35002
rect 10220 34930 10226 34969
rect 10260 34930 10266 34969
rect 10220 34901 10266 34930
rect 10220 34858 10226 34901
rect 10260 34858 10266 34901
rect 10220 34833 10266 34858
rect 10220 34786 10226 34833
rect 10260 34786 10266 34833
rect 10220 34765 10266 34786
rect 10220 34714 10226 34765
rect 10260 34714 10266 34765
rect 10220 34697 10266 34714
rect 10220 34642 10226 34697
rect 10260 34642 10266 34697
rect 10220 34629 10266 34642
rect 10220 34570 10226 34629
rect 10260 34570 10266 34629
rect 10220 34561 10266 34570
rect 10220 34498 10226 34561
rect 10260 34498 10266 34561
rect 10220 34493 10266 34498
rect 10220 34426 10226 34493
rect 10260 34426 10266 34493
rect 10220 34425 10266 34426
rect 10220 34391 10226 34425
rect 10260 34391 10266 34425
rect 10220 34388 10266 34391
rect 10220 34323 10226 34388
rect 10260 34323 10266 34388
rect 10220 34316 10266 34323
rect 10220 34255 10226 34316
rect 10260 34255 10266 34316
rect 10220 34244 10266 34255
rect 10220 34187 10226 34244
rect 10260 34187 10266 34244
rect 10220 34172 10266 34187
rect 10220 34119 10226 34172
rect 10260 34119 10266 34172
rect 10220 34100 10266 34119
rect 10220 34051 10226 34100
rect 10260 34051 10266 34100
rect 10220 34028 10266 34051
rect 10220 33983 10226 34028
rect 10260 33983 10266 34028
rect 10220 33956 10266 33983
rect 10220 33915 10226 33956
rect 10260 33915 10266 33956
rect 10220 33884 10266 33915
rect 10220 33847 10226 33884
rect 10260 33847 10266 33884
rect 10220 33813 10266 33847
rect 10220 33778 10226 33813
rect 10260 33778 10266 33813
rect 10220 33745 10266 33778
rect 10220 33706 10226 33745
rect 10260 33706 10266 33745
rect 10220 33677 10266 33706
rect 10220 33634 10226 33677
rect 10260 33634 10266 33677
rect 10220 33609 10266 33634
rect 10220 33562 10226 33609
rect 10260 33562 10266 33609
rect 10220 33541 10266 33562
rect 10220 33490 10226 33541
rect 10260 33490 10266 33541
rect 10220 33473 10266 33490
rect 10220 33418 10226 33473
rect 10260 33418 10266 33473
rect 10220 33405 10266 33418
rect 10220 33346 10226 33405
rect 10260 33346 10266 33405
rect 10220 33337 10266 33346
rect 10220 33274 10226 33337
rect 10260 33274 10266 33337
rect 10220 33269 10266 33274
rect 10220 33202 10226 33269
rect 10260 33202 10266 33269
rect 10220 33201 10266 33202
rect 10220 33167 10226 33201
rect 10260 33167 10266 33201
rect 10220 33164 10266 33167
rect 10220 33099 10226 33164
rect 10260 33099 10266 33164
rect 10220 33092 10266 33099
rect 10220 33031 10226 33092
rect 10260 33031 10266 33092
rect 10220 33020 10266 33031
rect 10220 32963 10226 33020
rect 10260 32963 10266 33020
rect 10220 32948 10266 32963
rect 10220 32895 10226 32948
rect 10260 32895 10266 32948
rect 10220 32876 10266 32895
rect 10220 32827 10226 32876
rect 10260 32827 10266 32876
rect 10220 32804 10266 32827
rect 10220 32759 10226 32804
rect 10260 32759 10266 32804
rect 10220 32732 10266 32759
rect 10220 32691 10226 32732
rect 10260 32691 10266 32732
rect 10220 32660 10266 32691
rect 10220 32623 10226 32660
rect 10260 32623 10266 32660
rect 10220 32589 10266 32623
rect 10220 32554 10226 32589
rect 10260 32554 10266 32589
rect 10220 32521 10266 32554
rect 10220 32482 10226 32521
rect 10260 32482 10266 32521
rect 10220 32453 10266 32482
rect 10220 32410 10226 32453
rect 10260 32410 10266 32453
rect 10220 32385 10266 32410
rect 10220 32338 10226 32385
rect 10260 32338 10266 32385
rect 10220 32317 10266 32338
rect 10220 32266 10226 32317
rect 10260 32266 10266 32317
rect 10220 32249 10266 32266
rect 10220 32194 10226 32249
rect 10260 32194 10266 32249
rect 10220 32181 10266 32194
rect 10220 32122 10226 32181
rect 10260 32122 10266 32181
rect 10220 32113 10266 32122
rect 10220 32050 10226 32113
rect 10260 32050 10266 32113
rect 10220 32045 10266 32050
rect 10220 31978 10226 32045
rect 10260 31978 10266 32045
rect 10220 31977 10266 31978
rect 10220 31943 10226 31977
rect 10260 31943 10266 31977
rect 10220 31940 10266 31943
rect 10220 31875 10226 31940
rect 10260 31875 10266 31940
rect 10220 31868 10266 31875
rect 10220 31807 10226 31868
rect 10260 31807 10266 31868
rect 10220 31796 10266 31807
rect 10220 31739 10226 31796
rect 10260 31739 10266 31796
rect 10220 31724 10266 31739
rect 10220 31671 10226 31724
rect 10260 31671 10266 31724
rect 10220 31652 10266 31671
rect 10220 31603 10226 31652
rect 10260 31603 10266 31652
rect 10220 31580 10266 31603
rect 10220 31535 10226 31580
rect 10260 31535 10266 31580
rect 10220 31508 10266 31535
rect 10220 31467 10226 31508
rect 10260 31467 10266 31508
rect 10220 31436 10266 31467
rect 10220 31399 10226 31436
rect 10260 31399 10266 31436
rect 10220 31365 10266 31399
rect 10220 31330 10226 31365
rect 10260 31330 10266 31365
rect 10220 31297 10266 31330
rect 10220 31258 10226 31297
rect 10260 31258 10266 31297
rect 10220 31229 10266 31258
rect 10220 31186 10226 31229
rect 10260 31186 10266 31229
rect 10220 31161 10266 31186
rect 10220 31114 10226 31161
rect 10260 31114 10266 31161
rect 10220 31093 10266 31114
rect 10220 31042 10226 31093
rect 10260 31042 10266 31093
rect 10220 31025 10266 31042
rect 10220 30970 10226 31025
rect 10260 30970 10266 31025
rect 10220 30957 10266 30970
rect 10220 30898 10226 30957
rect 10260 30898 10266 30957
rect 10220 30889 10266 30898
rect 10220 30826 10226 30889
rect 10260 30826 10266 30889
rect 10220 30821 10266 30826
rect 10220 30754 10226 30821
rect 10260 30754 10266 30821
rect 10220 30753 10266 30754
rect 10220 30719 10226 30753
rect 10260 30719 10266 30753
rect 10220 30716 10266 30719
rect 10220 30651 10226 30716
rect 10260 30651 10266 30716
rect 10220 30644 10266 30651
rect 10220 30583 10226 30644
rect 10260 30583 10266 30644
rect 10220 30572 10266 30583
rect 10220 30515 10226 30572
rect 10260 30515 10266 30572
rect 10220 30500 10266 30515
rect 10220 30447 10226 30500
rect 10260 30447 10266 30500
rect 10220 30428 10266 30447
rect 10220 30379 10226 30428
rect 10260 30379 10266 30428
rect 10220 30356 10266 30379
rect 10220 30311 10226 30356
rect 10260 30311 10266 30356
rect 10220 30284 10266 30311
rect 10220 30243 10226 30284
rect 10260 30243 10266 30284
rect 10220 30212 10266 30243
rect 10220 30175 10226 30212
rect 10260 30175 10266 30212
rect 10220 30141 10266 30175
rect 10220 30106 10226 30141
rect 10260 30106 10266 30141
rect 10220 30073 10266 30106
rect 10220 30034 10226 30073
rect 10260 30034 10266 30073
rect 10220 30005 10266 30034
rect 10220 29962 10226 30005
rect 10260 29962 10266 30005
rect 10220 29937 10266 29962
rect 10220 29890 10226 29937
rect 10260 29890 10266 29937
rect 10220 29869 10266 29890
rect 10220 29818 10226 29869
rect 10260 29818 10266 29869
rect 10220 29801 10266 29818
rect 10220 29746 10226 29801
rect 10260 29746 10266 29801
rect 10220 29733 10266 29746
rect 10220 29674 10226 29733
rect 10260 29674 10266 29733
rect 10220 29665 10266 29674
rect 10220 29602 10226 29665
rect 10260 29602 10266 29665
rect 10220 29597 10266 29602
rect 10220 29530 10226 29597
rect 10260 29530 10266 29597
rect 10220 29529 10266 29530
rect 10220 29495 10226 29529
rect 10260 29495 10266 29529
rect 10220 29492 10266 29495
rect 10220 29427 10226 29492
rect 10260 29427 10266 29492
rect 10220 29420 10266 29427
rect 10220 29359 10226 29420
rect 10260 29359 10266 29420
rect 10220 29348 10266 29359
rect 10220 29291 10226 29348
rect 10260 29291 10266 29348
rect 10220 29276 10266 29291
rect 10220 29223 10226 29276
rect 10260 29223 10266 29276
rect 10220 29204 10266 29223
rect 10220 29155 10226 29204
rect 10260 29155 10266 29204
rect 10220 29132 10266 29155
rect 10220 29087 10226 29132
rect 10260 29087 10266 29132
rect 10220 29060 10266 29087
rect 10220 29019 10226 29060
rect 10260 29019 10266 29060
rect 10220 28988 10266 29019
rect 10220 28951 10226 28988
rect 10260 28951 10266 28988
rect 10220 28917 10266 28951
rect 10220 28882 10226 28917
rect 10260 28882 10266 28917
rect 10220 28849 10266 28882
rect 10220 28810 10226 28849
rect 10260 28810 10266 28849
rect 10220 28781 10266 28810
rect 10220 28738 10226 28781
rect 10260 28738 10266 28781
rect 10220 28713 10266 28738
rect 10220 28666 10226 28713
rect 10260 28666 10266 28713
rect 10220 28645 10266 28666
rect 10220 28594 10226 28645
rect 10260 28594 10266 28645
rect 10220 28577 10266 28594
rect 10220 28522 10226 28577
rect 10260 28522 10266 28577
rect 10220 28509 10266 28522
rect 10220 28450 10226 28509
rect 10260 28450 10266 28509
rect 10220 28441 10266 28450
rect 10220 28378 10226 28441
rect 10260 28378 10266 28441
rect 10220 28373 10266 28378
rect 10220 28306 10226 28373
rect 10260 28306 10266 28373
rect 10220 28305 10266 28306
rect 10220 28271 10226 28305
rect 10260 28271 10266 28305
rect 10220 28268 10266 28271
rect 10220 28203 10226 28268
rect 10260 28203 10266 28268
rect 10220 28196 10266 28203
rect 10220 28135 10226 28196
rect 10260 28135 10266 28196
rect 10220 28124 10266 28135
rect 10220 28067 10226 28124
rect 10260 28067 10266 28124
rect 10220 28052 10266 28067
rect 10220 27999 10226 28052
rect 10260 27999 10266 28052
rect 10220 27980 10266 27999
rect 10220 27931 10226 27980
rect 10260 27931 10266 27980
rect 10220 27908 10266 27931
rect 10220 27863 10226 27908
rect 10260 27863 10266 27908
rect 10220 27836 10266 27863
rect 10220 27795 10226 27836
rect 10260 27795 10266 27836
rect 10220 27764 10266 27795
rect 10220 27727 10226 27764
rect 10260 27727 10266 27764
rect 10220 27693 10266 27727
rect 10220 27658 10226 27693
rect 10260 27658 10266 27693
rect 10220 27625 10266 27658
rect 10220 27586 10226 27625
rect 10260 27586 10266 27625
rect 10220 27557 10266 27586
rect 10220 27514 10226 27557
rect 10260 27514 10266 27557
rect 10220 27489 10266 27514
rect 10220 27442 10226 27489
rect 10260 27442 10266 27489
rect 10220 27421 10266 27442
rect 10220 27370 10226 27421
rect 10260 27370 10266 27421
rect 10220 27353 10266 27370
rect 10220 27298 10226 27353
rect 10260 27298 10266 27353
rect 10220 27285 10266 27298
rect 10220 27226 10226 27285
rect 10260 27226 10266 27285
rect 10220 27217 10266 27226
rect 10220 27154 10226 27217
rect 10260 27154 10266 27217
rect 10220 27149 10266 27154
rect 10220 27082 10226 27149
rect 10260 27082 10266 27149
rect 10220 27081 10266 27082
rect 10220 27047 10226 27081
rect 10260 27047 10266 27081
rect 10220 27044 10266 27047
rect 10220 26979 10226 27044
rect 10260 26979 10266 27044
rect 10220 26972 10266 26979
rect 10220 26911 10226 26972
rect 10260 26911 10266 26972
rect 10220 26900 10266 26911
rect 10220 26843 10226 26900
rect 10260 26843 10266 26900
rect 10220 26828 10266 26843
rect 10220 26775 10226 26828
rect 10260 26775 10266 26828
rect 10220 26756 10266 26775
rect 10220 26707 10226 26756
rect 10260 26707 10266 26756
rect 10220 26684 10266 26707
rect 10220 26639 10226 26684
rect 10260 26639 10266 26684
rect 10220 26612 10266 26639
rect 10220 26571 10226 26612
rect 10260 26571 10266 26612
rect 10220 26540 10266 26571
rect 10220 26503 10226 26540
rect 10260 26503 10266 26540
rect 10220 26469 10266 26503
rect 10220 26434 10226 26469
rect 10260 26434 10266 26469
rect 10220 26401 10266 26434
rect 10220 26362 10226 26401
rect 10260 26362 10266 26401
rect 10220 26333 10266 26362
rect 10220 26290 10226 26333
rect 10260 26290 10266 26333
rect 10220 26265 10266 26290
rect 10220 26218 10226 26265
rect 10260 26218 10266 26265
rect 10220 26197 10266 26218
rect 10220 26146 10226 26197
rect 10260 26146 10266 26197
rect 10220 26129 10266 26146
rect 10220 26074 10226 26129
rect 10260 26074 10266 26129
rect 10220 26061 10266 26074
rect 10220 26002 10226 26061
rect 10260 26002 10266 26061
rect 10220 25993 10266 26002
rect 10220 25930 10226 25993
rect 10260 25930 10266 25993
rect 10220 25925 10266 25930
rect 10220 25858 10226 25925
rect 10260 25858 10266 25925
rect 10220 25857 10266 25858
rect 10220 25823 10226 25857
rect 10260 25823 10266 25857
rect 10220 25820 10266 25823
rect 10220 25755 10226 25820
rect 10260 25755 10266 25820
rect 10220 25748 10266 25755
rect 10220 25687 10226 25748
rect 10260 25687 10266 25748
rect 10220 25676 10266 25687
rect 10220 25619 10226 25676
rect 10260 25619 10266 25676
rect 10220 25604 10266 25619
rect 10220 25551 10226 25604
rect 10260 25551 10266 25604
rect 10220 25532 10266 25551
rect 10220 25483 10226 25532
rect 10260 25483 10266 25532
rect 10220 25460 10266 25483
rect 10220 25415 10226 25460
rect 10260 25415 10266 25460
rect 10220 25388 10266 25415
rect 10220 25347 10226 25388
rect 10260 25347 10266 25388
rect 10220 25316 10266 25347
rect 10220 25279 10226 25316
rect 10260 25279 10266 25316
rect 10220 25245 10266 25279
rect 10220 25210 10226 25245
rect 10260 25210 10266 25245
rect 10220 25177 10266 25210
rect 10220 25138 10226 25177
rect 10260 25138 10266 25177
rect 10220 25109 10266 25138
rect 10220 25066 10226 25109
rect 10260 25066 10266 25109
rect 10220 25041 10266 25066
rect 10220 24994 10226 25041
rect 10260 24994 10266 25041
rect 10220 24973 10266 24994
rect 10220 24922 10226 24973
rect 10260 24922 10266 24973
rect 10220 24905 10266 24922
rect 10220 24850 10226 24905
rect 10260 24850 10266 24905
rect 10220 24837 10266 24850
rect 10220 24778 10226 24837
rect 10260 24778 10266 24837
rect 10220 24769 10266 24778
rect 10220 24706 10226 24769
rect 10260 24706 10266 24769
rect 10220 24701 10266 24706
rect 10220 24634 10226 24701
rect 10260 24634 10266 24701
rect 10220 24633 10266 24634
rect 10220 24599 10226 24633
rect 10260 24599 10266 24633
rect 10220 24596 10266 24599
rect 10220 24531 10226 24596
rect 10260 24531 10266 24596
rect 10220 24524 10266 24531
rect 10220 24463 10226 24524
rect 10260 24463 10266 24524
rect 10220 24452 10266 24463
rect 10220 24395 10226 24452
rect 10260 24395 10266 24452
rect 10220 24380 10266 24395
rect 10220 24327 10226 24380
rect 10260 24327 10266 24380
rect 10220 24308 10266 24327
rect 10220 24259 10226 24308
rect 10260 24259 10266 24308
rect 10220 24236 10266 24259
rect 10220 24191 10226 24236
rect 10260 24191 10266 24236
rect 10220 24164 10266 24191
rect 10220 24123 10226 24164
rect 10260 24123 10266 24164
rect 10220 24092 10266 24123
rect 10220 24055 10226 24092
rect 10260 24055 10266 24092
rect 10220 24021 10266 24055
rect 10220 23986 10226 24021
rect 10260 23986 10266 24021
rect 10220 23953 10266 23986
rect 10220 23914 10226 23953
rect 10260 23914 10266 23953
rect 10220 23885 10266 23914
rect 10220 23842 10226 23885
rect 10260 23842 10266 23885
rect 10220 23817 10266 23842
rect 10220 23770 10226 23817
rect 10260 23770 10266 23817
rect 10220 23749 10266 23770
rect 10220 23698 10226 23749
rect 10260 23698 10266 23749
rect 10220 23681 10266 23698
rect 10220 23626 10226 23681
rect 10260 23626 10266 23681
rect 10220 23613 10266 23626
rect 10220 23554 10226 23613
rect 10260 23554 10266 23613
rect 10220 23545 10266 23554
rect 10220 23482 10226 23545
rect 10260 23482 10266 23545
rect 10220 23477 10266 23482
rect 10220 23410 10226 23477
rect 10260 23410 10266 23477
rect 10220 23409 10266 23410
rect 10220 23375 10226 23409
rect 10260 23375 10266 23409
rect 10220 23372 10266 23375
rect 10220 23307 10226 23372
rect 10260 23307 10266 23372
rect 10220 23300 10266 23307
rect 10220 23239 10226 23300
rect 10260 23239 10266 23300
rect 10220 23228 10266 23239
rect 10220 23171 10226 23228
rect 10260 23171 10266 23228
rect 10220 23156 10266 23171
rect 10220 23103 10226 23156
rect 10260 23103 10266 23156
rect 10220 23084 10266 23103
rect 10220 23035 10226 23084
rect 10260 23035 10266 23084
rect 10220 23012 10266 23035
rect 10220 22967 10226 23012
rect 10260 22967 10266 23012
rect 10220 22940 10266 22967
rect 10220 22899 10226 22940
rect 10260 22899 10266 22940
rect 10220 22868 10266 22899
rect 10220 22831 10226 22868
rect 10260 22831 10266 22868
rect 10220 22797 10266 22831
rect 10220 22762 10226 22797
rect 10260 22762 10266 22797
rect 10220 22729 10266 22762
rect 10220 22690 10226 22729
rect 10260 22690 10266 22729
rect 10220 22661 10266 22690
rect 10220 22618 10226 22661
rect 10260 22618 10266 22661
rect 10220 22593 10266 22618
rect 10220 22546 10226 22593
rect 10260 22546 10266 22593
rect 10220 22525 10266 22546
rect 10220 22474 10226 22525
rect 10260 22474 10266 22525
rect 10220 22457 10266 22474
rect 10220 22402 10226 22457
rect 10260 22402 10266 22457
rect 10220 22389 10266 22402
rect 10220 22330 10226 22389
rect 10260 22330 10266 22389
rect 10220 22321 10266 22330
rect 10220 22258 10226 22321
rect 10260 22258 10266 22321
rect 10220 22253 10266 22258
rect 10220 22186 10226 22253
rect 10260 22186 10266 22253
rect 10220 22185 10266 22186
rect 10220 22151 10226 22185
rect 10260 22151 10266 22185
rect 10220 22148 10266 22151
rect 10220 22083 10226 22148
rect 10260 22083 10266 22148
rect 10220 22076 10266 22083
rect 10220 22015 10226 22076
rect 10260 22015 10266 22076
rect 10220 22004 10266 22015
rect 10220 21947 10226 22004
rect 10260 21947 10266 22004
rect 10220 21932 10266 21947
rect 10220 21879 10226 21932
rect 10260 21879 10266 21932
rect 10220 21860 10266 21879
rect 10220 21811 10226 21860
rect 10260 21811 10266 21860
rect 10220 21788 10266 21811
rect 10220 21743 10226 21788
rect 10260 21743 10266 21788
rect 10220 21716 10266 21743
rect 10220 21675 10226 21716
rect 10260 21675 10266 21716
rect 10220 21644 10266 21675
rect 10220 21607 10226 21644
rect 10260 21607 10266 21644
rect 10220 21573 10266 21607
rect 10220 21538 10226 21573
rect 10260 21538 10266 21573
rect 10220 21505 10266 21538
rect 10220 21466 10226 21505
rect 10260 21466 10266 21505
rect 10220 21437 10266 21466
rect 10220 21394 10226 21437
rect 10260 21394 10266 21437
rect 10220 21369 10266 21394
rect 10220 21322 10226 21369
rect 10260 21322 10266 21369
rect 10220 21301 10266 21322
rect 10220 21250 10226 21301
rect 10260 21250 10266 21301
rect 10220 21233 10266 21250
rect 10220 21178 10226 21233
rect 10260 21178 10266 21233
rect 10220 21165 10266 21178
rect 10220 21106 10226 21165
rect 10260 21106 10266 21165
rect 10220 21097 10266 21106
rect 10220 21034 10226 21097
rect 10260 21034 10266 21097
rect 10220 21029 10266 21034
rect 10220 20962 10226 21029
rect 10260 20962 10266 21029
rect 10220 20961 10266 20962
rect 10220 20927 10226 20961
rect 10260 20927 10266 20961
rect 10220 20924 10266 20927
rect 10220 20859 10226 20924
rect 10260 20859 10266 20924
rect 10220 20852 10266 20859
rect 10220 20791 10226 20852
rect 10260 20791 10266 20852
rect 10220 20780 10266 20791
rect 10220 20723 10226 20780
rect 10260 20723 10266 20780
rect 10220 20708 10266 20723
rect 10220 20655 10226 20708
rect 10260 20655 10266 20708
rect 10220 20636 10266 20655
rect 10220 20587 10226 20636
rect 10260 20587 10266 20636
rect 10220 20564 10266 20587
rect 10220 20519 10226 20564
rect 10260 20519 10266 20564
rect 10220 20492 10266 20519
rect 10220 20451 10226 20492
rect 10260 20451 10266 20492
rect 10220 20420 10266 20451
rect 10220 20383 10226 20420
rect 10260 20383 10266 20420
rect 10220 20349 10266 20383
rect 10220 20314 10226 20349
rect 10260 20314 10266 20349
rect 10220 20281 10266 20314
rect 10220 20242 10226 20281
rect 10260 20242 10266 20281
rect 10220 20213 10266 20242
rect 10220 20170 10226 20213
rect 10260 20170 10266 20213
rect 10220 20145 10266 20170
rect 10220 20098 10226 20145
rect 10260 20098 10266 20145
rect 10220 20077 10266 20098
rect 10220 20026 10226 20077
rect 10260 20026 10266 20077
rect 10220 20009 10266 20026
rect 10220 19954 10226 20009
rect 10260 19954 10266 20009
rect 10220 19941 10266 19954
rect 10220 19882 10226 19941
rect 10260 19882 10266 19941
rect 10220 19873 10266 19882
rect 10220 19810 10226 19873
rect 10260 19810 10266 19873
rect 10220 19805 10266 19810
rect 10220 19738 10226 19805
rect 10260 19738 10266 19805
rect 10220 19737 10266 19738
rect 10220 19703 10226 19737
rect 10260 19703 10266 19737
rect 10220 19700 10266 19703
rect 10220 19635 10226 19700
rect 10260 19635 10266 19700
rect 10220 19628 10266 19635
rect 10220 19567 10226 19628
rect 10260 19567 10266 19628
rect 10220 19556 10266 19567
rect 10220 19499 10226 19556
rect 10260 19499 10266 19556
rect 10220 19484 10266 19499
rect 10220 19431 10226 19484
rect 10260 19431 10266 19484
rect 10220 19412 10266 19431
rect 10220 19363 10226 19412
rect 10260 19363 10266 19412
rect 10220 19340 10266 19363
rect 10220 19295 10226 19340
rect 10260 19295 10266 19340
rect 10220 19268 10266 19295
rect 10220 19227 10226 19268
rect 10260 19227 10266 19268
rect 10220 19196 10266 19227
rect 10220 19159 10226 19196
rect 10260 19159 10266 19196
rect 10220 19125 10266 19159
rect 10220 19090 10226 19125
rect 10260 19090 10266 19125
rect 10220 19057 10266 19090
rect 10220 19018 10226 19057
rect 10260 19018 10266 19057
rect 10220 18989 10266 19018
rect 10220 18946 10226 18989
rect 10260 18946 10266 18989
rect 10220 18921 10266 18946
rect 10220 18874 10226 18921
rect 10260 18874 10266 18921
rect 10220 18853 10266 18874
rect 10220 18802 10226 18853
rect 10260 18802 10266 18853
rect 10220 18785 10266 18802
rect 10220 18730 10226 18785
rect 10260 18730 10266 18785
rect 10220 18717 10266 18730
rect 10220 18658 10226 18717
rect 10260 18658 10266 18717
rect 10220 18649 10266 18658
rect 10220 18586 10226 18649
rect 10260 18586 10266 18649
rect 10220 18581 10266 18586
rect 10220 18514 10226 18581
rect 10260 18514 10266 18581
rect 10220 18513 10266 18514
rect 10220 18479 10226 18513
rect 10260 18479 10266 18513
rect 10220 18476 10266 18479
rect 10220 18411 10226 18476
rect 10260 18411 10266 18476
rect 10220 18404 10266 18411
rect 10220 18343 10226 18404
rect 10260 18343 10266 18404
rect 10220 18332 10266 18343
rect 10220 18275 10226 18332
rect 10260 18275 10266 18332
rect 10220 18260 10266 18275
rect 10220 18207 10226 18260
rect 10260 18207 10266 18260
rect 10220 18188 10266 18207
rect 10220 18139 10226 18188
rect 10260 18139 10266 18188
rect 10220 18116 10266 18139
rect 10220 18071 10226 18116
rect 10260 18071 10266 18116
rect 10220 18044 10266 18071
rect 10220 18003 10226 18044
rect 10260 18003 10266 18044
rect 10220 17972 10266 18003
rect 10220 17935 10226 17972
rect 10260 17935 10266 17972
rect 10220 17901 10266 17935
rect 10220 17866 10226 17901
rect 10260 17866 10266 17901
rect 10220 17833 10266 17866
rect 10220 17794 10226 17833
rect 10260 17794 10266 17833
rect 10220 17765 10266 17794
rect 10220 17722 10226 17765
rect 10260 17722 10266 17765
rect 10220 17697 10266 17722
rect 10220 17650 10226 17697
rect 10260 17650 10266 17697
rect 10220 17629 10266 17650
rect 10220 17578 10226 17629
rect 10260 17578 10266 17629
rect 10220 17561 10266 17578
rect 10220 17506 10226 17561
rect 10260 17506 10266 17561
rect 10220 17493 10266 17506
rect 10220 17434 10226 17493
rect 10260 17434 10266 17493
rect 10220 17425 10266 17434
rect 10220 17362 10226 17425
rect 10260 17362 10266 17425
rect 10220 17357 10266 17362
rect 10220 17290 10226 17357
rect 10260 17290 10266 17357
rect 10220 17289 10266 17290
rect 10220 17255 10226 17289
rect 10260 17255 10266 17289
rect 10220 17252 10266 17255
rect 10220 17187 10226 17252
rect 10260 17187 10266 17252
rect 10220 17180 10266 17187
rect 10220 17119 10226 17180
rect 10260 17119 10266 17180
rect 10220 17108 10266 17119
rect 10220 17051 10226 17108
rect 10260 17051 10266 17108
rect 10220 17036 10266 17051
rect 10220 16983 10226 17036
rect 10260 16983 10266 17036
rect 10220 16964 10266 16983
rect 10220 16915 10226 16964
rect 10260 16915 10266 16964
rect 10220 16892 10266 16915
rect 10220 16847 10226 16892
rect 10260 16847 10266 16892
rect 10220 16820 10266 16847
rect 10220 16779 10226 16820
rect 10260 16779 10266 16820
rect 10220 16748 10266 16779
rect 10220 16711 10226 16748
rect 10260 16711 10266 16748
rect 10220 16677 10266 16711
rect 10220 16642 10226 16677
rect 10260 16642 10266 16677
rect 10220 16609 10266 16642
rect 10220 16570 10226 16609
rect 10260 16570 10266 16609
rect 10220 16541 10266 16570
rect 10220 16498 10226 16541
rect 10260 16498 10266 16541
rect 10220 16473 10266 16498
rect 10220 16426 10226 16473
rect 10260 16426 10266 16473
rect 10220 16405 10266 16426
rect 10220 16354 10226 16405
rect 10260 16354 10266 16405
rect 10220 16337 10266 16354
rect 10220 16282 10226 16337
rect 10260 16282 10266 16337
rect 10220 16269 10266 16282
rect 10220 16210 10226 16269
rect 10260 16210 10266 16269
rect 10220 16201 10266 16210
rect 10220 16138 10226 16201
rect 10260 16138 10266 16201
rect 10220 16133 10266 16138
rect 10220 16066 10226 16133
rect 10260 16066 10266 16133
rect 10220 16065 10266 16066
rect 10220 16031 10226 16065
rect 10260 16031 10266 16065
rect 10220 16028 10266 16031
rect 10220 15963 10226 16028
rect 10260 15963 10266 16028
rect 10220 15956 10266 15963
rect 10220 15895 10226 15956
rect 10260 15895 10266 15956
rect 10220 15884 10266 15895
rect 10220 15827 10226 15884
rect 10260 15827 10266 15884
rect 10220 15812 10266 15827
rect 10220 15759 10226 15812
rect 10260 15759 10266 15812
rect 10220 15740 10266 15759
rect 10220 15691 10226 15740
rect 10260 15691 10266 15740
rect 10220 15668 10266 15691
rect 10220 15623 10226 15668
rect 10260 15623 10266 15668
rect 10220 15596 10266 15623
rect 10220 15555 10226 15596
rect 10260 15555 10266 15596
rect 10220 15524 10266 15555
rect 10220 15487 10226 15524
rect 10260 15487 10266 15524
rect 10220 15453 10266 15487
rect 10220 15418 10226 15453
rect 10260 15418 10266 15453
rect 10220 15385 10266 15418
rect 10220 15346 10226 15385
rect 10260 15346 10266 15385
rect 10220 15317 10266 15346
rect 10220 15274 10226 15317
rect 10260 15274 10266 15317
rect 10220 15249 10266 15274
rect 10220 15202 10226 15249
rect 10260 15202 10266 15249
rect 10220 15181 10266 15202
rect 10220 15130 10226 15181
rect 10260 15130 10266 15181
rect 10220 15113 10266 15130
rect 10220 15058 10226 15113
rect 10260 15058 10266 15113
rect 10220 15045 10266 15058
rect 10220 14986 10226 15045
rect 10260 14986 10266 15045
rect 10220 14977 10266 14986
rect 10220 14914 10226 14977
rect 10260 14914 10266 14977
rect 10220 14909 10266 14914
rect 10220 14842 10226 14909
rect 10260 14842 10266 14909
rect 10220 14841 10266 14842
rect 10220 14807 10226 14841
rect 10260 14807 10266 14841
rect 10220 14804 10266 14807
rect 10220 14739 10226 14804
rect 10260 14739 10266 14804
rect 10220 14732 10266 14739
rect 10220 14671 10226 14732
rect 10260 14671 10266 14732
rect 10220 14660 10266 14671
rect 10220 14603 10226 14660
rect 10260 14603 10266 14660
rect 10220 14588 10266 14603
rect 10220 14535 10226 14588
rect 10260 14535 10266 14588
rect 10220 14516 10266 14535
rect 10220 14467 10226 14516
rect 10260 14467 10266 14516
rect 10220 14444 10266 14467
rect 10220 14399 10226 14444
rect 10260 14399 10266 14444
rect 10220 14372 10266 14399
rect 10220 14331 10226 14372
rect 10260 14331 10266 14372
rect 10220 14300 10266 14331
rect 10220 14263 10226 14300
rect 10260 14263 10266 14300
rect 10220 14229 10266 14263
rect 10220 14194 10226 14229
rect 10260 14194 10266 14229
rect 10220 14161 10266 14194
rect 10220 14122 10226 14161
rect 10260 14122 10266 14161
rect 10220 14093 10266 14122
rect 10220 14050 10226 14093
rect 10260 14050 10266 14093
rect 10220 14025 10266 14050
rect 10220 13978 10226 14025
rect 10260 13978 10266 14025
rect 10220 13957 10266 13978
rect 10220 13906 10226 13957
rect 10260 13906 10266 13957
rect 10220 13889 10266 13906
rect 10220 13834 10226 13889
rect 10260 13834 10266 13889
rect 10220 13821 10266 13834
rect 10220 13762 10226 13821
rect 10260 13762 10266 13821
rect 10220 13753 10266 13762
rect 10220 13690 10226 13753
rect 10260 13690 10266 13753
rect 10220 13685 10266 13690
rect 10220 13618 10226 13685
rect 10260 13618 10266 13685
rect 10220 13617 10266 13618
rect 10220 13583 10226 13617
rect 10260 13583 10266 13617
rect 10220 13580 10266 13583
rect 10220 13515 10226 13580
rect 10260 13515 10266 13580
rect 10220 13508 10266 13515
rect 10220 13447 10226 13508
rect 10260 13447 10266 13508
rect 10220 13436 10266 13447
rect 10220 13379 10226 13436
rect 10260 13379 10266 13436
rect 10220 13364 10266 13379
rect 10220 13311 10226 13364
rect 10260 13311 10266 13364
rect 10220 13292 10266 13311
rect 10220 13243 10226 13292
rect 10260 13243 10266 13292
rect 10220 13220 10266 13243
rect 10220 13175 10226 13220
rect 10260 13175 10266 13220
rect 10220 13148 10266 13175
rect 10220 13107 10226 13148
rect 10260 13107 10266 13148
rect 10220 13076 10266 13107
rect 10220 13039 10226 13076
rect 10260 13039 10266 13076
rect 10220 13005 10266 13039
rect 10220 12970 10226 13005
rect 10260 12970 10266 13005
rect 10220 12937 10266 12970
rect 10220 12898 10226 12937
rect 10260 12898 10266 12937
rect 10220 12869 10266 12898
rect 10220 12826 10226 12869
rect 10260 12826 10266 12869
rect 10220 12801 10266 12826
rect 10220 12754 10226 12801
rect 10260 12754 10266 12801
rect 10220 12733 10266 12754
rect 10220 12682 10226 12733
rect 10260 12682 10266 12733
rect 10220 12665 10266 12682
rect 10220 12610 10226 12665
rect 10260 12610 10266 12665
rect 10220 12597 10266 12610
rect 10220 12538 10226 12597
rect 10260 12538 10266 12597
rect 10220 12529 10266 12538
rect 10220 12466 10226 12529
rect 10260 12466 10266 12529
rect 10220 12461 10266 12466
rect 10220 12394 10226 12461
rect 10260 12394 10266 12461
rect 10220 12393 10266 12394
rect 10220 12359 10226 12393
rect 10260 12359 10266 12393
rect 10220 12356 10266 12359
rect 10220 12291 10226 12356
rect 10260 12291 10266 12356
rect 10220 12284 10266 12291
rect 10220 12223 10226 12284
rect 10260 12223 10266 12284
rect 10220 12212 10266 12223
rect 10220 12155 10226 12212
rect 10260 12155 10266 12212
rect 10220 12140 10266 12155
rect 10220 12087 10226 12140
rect 10260 12087 10266 12140
rect 10220 12068 10266 12087
rect 10220 12019 10226 12068
rect 10260 12019 10266 12068
rect 10220 11996 10266 12019
rect 10220 11951 10226 11996
rect 10260 11951 10266 11996
rect 10220 11924 10266 11951
rect 10220 11883 10226 11924
rect 10260 11883 10266 11924
rect 10220 11852 10266 11883
rect 10220 11815 10226 11852
rect 10260 11815 10266 11852
rect 10220 11781 10266 11815
rect 10220 11746 10226 11781
rect 10260 11746 10266 11781
rect 10220 11713 10266 11746
rect 10220 11674 10226 11713
rect 10260 11674 10266 11713
rect 10220 11645 10266 11674
rect 10220 11602 10226 11645
rect 10260 11602 10266 11645
rect 10220 11577 10266 11602
rect 10220 11530 10226 11577
rect 10260 11530 10266 11577
rect 10220 11509 10266 11530
rect 10220 11458 10226 11509
rect 10260 11458 10266 11509
rect 10220 11441 10266 11458
rect 10220 11386 10226 11441
rect 10260 11386 10266 11441
rect 10220 11373 10266 11386
rect 10220 11314 10226 11373
rect 10260 11314 10266 11373
rect 10220 11305 10266 11314
rect 10220 11242 10226 11305
rect 10260 11242 10266 11305
rect 10220 11237 10266 11242
rect 10220 11170 10226 11237
rect 10260 11170 10266 11237
rect 10220 11169 10266 11170
rect 10220 11135 10226 11169
rect 10260 11135 10266 11169
rect 10220 11132 10266 11135
rect 10220 11067 10226 11132
rect 10260 11067 10266 11132
rect 10220 11060 10266 11067
rect 10220 10999 10226 11060
rect 10260 10999 10266 11060
rect 10220 10988 10266 10999
rect 10220 10931 10226 10988
rect 10260 10931 10266 10988
rect 10220 10916 10266 10931
rect 10220 10863 10226 10916
rect 10260 10863 10266 10916
rect 10220 10844 10266 10863
rect 10220 10795 10226 10844
rect 10260 10795 10266 10844
rect 10220 10772 10266 10795
rect 10220 10727 10226 10772
rect 10260 10727 10266 10772
rect 10220 10700 10266 10727
rect 10220 10659 10226 10700
rect 10260 10659 10266 10700
rect 10220 10628 10266 10659
rect 10220 10591 10226 10628
rect 10260 10591 10266 10628
rect 10220 10557 10266 10591
rect 10220 10522 10226 10557
rect 10260 10522 10266 10557
rect 10220 10489 10266 10522
rect 10220 10450 10226 10489
rect 10260 10450 10266 10489
rect 10220 10421 10266 10450
rect 10220 10378 10226 10421
rect 10260 10378 10266 10421
rect 10220 10353 10266 10378
rect 10220 10306 10226 10353
rect 10260 10306 10266 10353
rect 10220 10285 10266 10306
rect 10220 10234 10226 10285
rect 10260 10234 10266 10285
rect 10220 10217 10266 10234
rect 10220 10162 10226 10217
rect 10260 10162 10266 10217
rect 10220 10149 10266 10162
rect 10220 10090 10226 10149
rect 10260 10090 10266 10149
rect 10220 10081 10266 10090
rect 10220 10018 10226 10081
rect 10260 10018 10266 10081
rect 10220 10013 10266 10018
rect 10220 9946 10226 10013
rect 10260 9946 10266 10013
rect 10220 9945 10266 9946
rect 10220 9911 10226 9945
rect 10260 9911 10266 9945
rect 10220 9908 10266 9911
rect 10220 9843 10226 9908
rect 10260 9843 10266 9908
rect 10220 9836 10266 9843
rect 10220 9775 10226 9836
rect 10260 9775 10266 9836
rect 10220 9764 10266 9775
rect 10220 9707 10226 9764
rect 10260 9707 10266 9764
rect 10220 9692 10266 9707
rect 10220 9639 10226 9692
rect 10260 9639 10266 9692
rect 10220 9620 10266 9639
rect 10220 9571 10226 9620
rect 10260 9571 10266 9620
rect 10220 9548 10266 9571
rect 10220 9503 10226 9548
rect 10260 9503 10266 9548
rect 10220 9476 10266 9503
rect 10220 9435 10226 9476
rect 10260 9435 10266 9476
rect 10220 9404 10266 9435
rect 10220 9367 10226 9404
rect 10260 9367 10266 9404
rect 10220 9333 10266 9367
rect 10220 9298 10226 9333
rect 10260 9298 10266 9333
rect 10220 9265 10266 9298
rect 10220 9226 10226 9265
rect 10260 9226 10266 9265
rect 10220 9197 10266 9226
rect 10220 9154 10226 9197
rect 10260 9154 10266 9197
rect 10220 9129 10266 9154
rect 10220 9082 10226 9129
rect 10260 9082 10266 9129
rect 10220 9061 10266 9082
rect 10220 9010 10226 9061
rect 10260 9010 10266 9061
rect 10220 8993 10266 9010
rect 10220 8938 10226 8993
rect 10260 8938 10266 8993
rect 10220 8925 10266 8938
rect 10220 8866 10226 8925
rect 10260 8866 10266 8925
rect 10220 8857 10266 8866
rect 10220 8794 10226 8857
rect 10260 8794 10266 8857
rect 10220 8789 10266 8794
rect 10220 8722 10226 8789
rect 10260 8722 10266 8789
rect 10220 8721 10266 8722
rect 10220 8687 10226 8721
rect 10260 8687 10266 8721
rect 10220 8684 10266 8687
rect 10220 8619 10226 8684
rect 10260 8619 10266 8684
rect 10220 8612 10266 8619
rect 10220 8551 10226 8612
rect 10260 8551 10266 8612
rect 10220 8540 10266 8551
rect 10220 8483 10226 8540
rect 10260 8483 10266 8540
rect 10220 8468 10266 8483
rect 10220 8415 10226 8468
rect 10260 8415 10266 8468
rect 10220 8396 10266 8415
rect 10220 8347 10226 8396
rect 10260 8347 10266 8396
rect 10220 8324 10266 8347
rect 10220 8279 10226 8324
rect 10260 8279 10266 8324
rect 10220 8252 10266 8279
rect 10220 8211 10226 8252
rect 10260 8211 10266 8252
rect 10220 8180 10266 8211
rect 10220 8143 10226 8180
rect 10260 8143 10266 8180
rect 10220 8109 10266 8143
rect 10220 8074 10226 8109
rect 10260 8074 10266 8109
rect 10220 8041 10266 8074
rect 10220 8002 10226 8041
rect 10260 8002 10266 8041
rect 10220 7973 10266 8002
rect 10220 7930 10226 7973
rect 10260 7930 10266 7973
rect 10220 7905 10266 7930
rect 10220 7858 10226 7905
rect 10260 7858 10266 7905
rect 10220 7837 10266 7858
rect 10220 7786 10226 7837
rect 10260 7786 10266 7837
rect 10220 7769 10266 7786
rect 10220 7714 10226 7769
rect 10260 7714 10266 7769
rect 10220 7701 10266 7714
rect 10220 7642 10226 7701
rect 10260 7642 10266 7701
rect 10220 7633 10266 7642
rect 10220 7570 10226 7633
rect 10260 7570 10266 7633
rect 10220 7565 10266 7570
rect 10220 7498 10226 7565
rect 10260 7498 10266 7565
rect 10220 7497 10266 7498
rect 10220 7463 10226 7497
rect 10260 7463 10266 7497
rect 10220 7460 10266 7463
rect 10220 7395 10226 7460
rect 10260 7395 10266 7460
rect 10220 7388 10266 7395
rect 10220 7327 10226 7388
rect 10260 7327 10266 7388
rect 10220 7316 10266 7327
rect 10220 7259 10226 7316
rect 10260 7259 10266 7316
rect 10220 7244 10266 7259
rect 10220 7191 10226 7244
rect 10260 7191 10266 7244
rect 10220 7172 10266 7191
rect 10220 7123 10226 7172
rect 10260 7123 10266 7172
rect 10220 7100 10266 7123
rect 10220 7055 10226 7100
rect 10260 7055 10266 7100
rect 10220 7028 10266 7055
rect 10220 6987 10226 7028
rect 10260 6987 10266 7028
rect 10220 6956 10266 6987
rect 10220 6919 10226 6956
rect 10260 6919 10266 6956
rect 10220 6885 10266 6919
rect 10220 6850 10226 6885
rect 10260 6850 10266 6885
rect 10220 6817 10266 6850
rect 10220 6778 10226 6817
rect 10260 6778 10266 6817
rect 10220 6749 10266 6778
rect 10220 6706 10226 6749
rect 10260 6706 10266 6749
rect 10220 6681 10266 6706
rect 10220 6634 10226 6681
rect 10260 6634 10266 6681
rect 10220 6613 10266 6634
rect 10220 6562 10226 6613
rect 10260 6562 10266 6613
rect 10220 6545 10266 6562
rect 10220 6490 10226 6545
rect 10260 6490 10266 6545
rect 10220 6477 10266 6490
rect 10220 6418 10226 6477
rect 10260 6418 10266 6477
rect 10220 6409 10266 6418
rect 10220 6346 10226 6409
rect 10260 6346 10266 6409
rect 10220 6341 10266 6346
rect 10220 6274 10226 6341
rect 10260 6274 10266 6341
rect 10220 6273 10266 6274
rect 10220 6239 10226 6273
rect 10260 6239 10266 6273
rect 10220 6236 10266 6239
rect 10220 6171 10226 6236
rect 10260 6171 10266 6236
rect 10220 6164 10266 6171
rect 10220 6103 10226 6164
rect 10260 6103 10266 6164
rect 10220 6092 10266 6103
rect 10220 6035 10226 6092
rect 10260 6035 10266 6092
rect 10220 6020 10266 6035
rect 10220 5967 10226 6020
rect 10260 5967 10266 6020
rect 10220 5948 10266 5967
rect 10220 5899 10226 5948
rect 10260 5899 10266 5948
rect 10220 5876 10266 5899
rect 10220 5831 10226 5876
rect 10260 5831 10266 5876
rect 10220 5804 10266 5831
rect 10220 5763 10226 5804
rect 10260 5763 10266 5804
rect 10220 5732 10266 5763
rect 10220 5695 10226 5732
rect 10260 5695 10266 5732
rect 10220 5661 10266 5695
rect 10220 5626 10226 5661
rect 10260 5626 10266 5661
rect 10220 5593 10266 5626
rect 10220 5554 10226 5593
rect 10260 5554 10266 5593
rect 10220 5525 10266 5554
rect 10220 5482 10226 5525
rect 10260 5482 10266 5525
rect 10220 5457 10266 5482
rect 10220 5410 10226 5457
rect 10260 5410 10266 5457
rect 10220 5389 10266 5410
rect 10220 5338 10226 5389
rect 10260 5338 10266 5389
rect 10220 5321 10266 5338
rect 10220 5266 10226 5321
rect 10260 5266 10266 5321
rect 10220 5253 10266 5266
rect 10220 5194 10226 5253
rect 10260 5194 10266 5253
rect 10220 5185 10266 5194
rect 10220 5122 10226 5185
rect 10260 5122 10266 5185
rect 10220 5117 10266 5122
rect 10220 5050 10226 5117
rect 10260 5050 10266 5117
rect 10220 5049 10266 5050
rect 10220 5015 10226 5049
rect 10260 5015 10266 5049
rect 10220 5012 10266 5015
rect 10220 4947 10226 5012
rect 10260 4947 10266 5012
rect 10220 4940 10266 4947
rect 10220 4879 10226 4940
rect 10260 4879 10266 4940
rect 10220 4868 10266 4879
rect 10220 4811 10226 4868
rect 10260 4811 10266 4868
rect 10220 4796 10266 4811
rect 10220 4743 10226 4796
rect 10260 4743 10266 4796
rect 10220 4724 10266 4743
rect 10220 4675 10226 4724
rect 10260 4675 10266 4724
rect 10220 4652 10266 4675
rect 10220 4607 10226 4652
rect 10260 4607 10266 4652
rect 10220 4580 10266 4607
rect 10220 4539 10226 4580
rect 10260 4539 10266 4580
rect 10220 4508 10266 4539
rect 10220 4471 10226 4508
rect 10260 4471 10266 4508
rect 10220 4437 10266 4471
rect 10220 4402 10226 4437
rect 10260 4402 10266 4437
rect 10220 4369 10266 4402
rect 10220 4330 10226 4369
rect 10260 4330 10266 4369
rect 10220 4301 10266 4330
rect 10220 4258 10226 4301
rect 10260 4258 10266 4301
rect 10220 4233 10266 4258
rect 10220 4186 10226 4233
rect 10260 4186 10266 4233
rect 10220 4165 10266 4186
rect 10220 4114 10226 4165
rect 10260 4114 10266 4165
rect 10220 4097 10266 4114
rect 10220 4042 10226 4097
rect 10260 4042 10266 4097
rect 10220 4029 10266 4042
rect 10220 3970 10226 4029
rect 10260 3970 10266 4029
rect 10220 3961 10266 3970
rect 10220 3898 10226 3961
rect 10260 3898 10266 3961
rect 10220 3893 10266 3898
rect 10220 3826 10226 3893
rect 10260 3826 10266 3893
rect 10220 3825 10266 3826
rect 10220 3791 10226 3825
rect 10260 3791 10266 3825
rect 10220 3788 10266 3791
rect 10220 3723 10226 3788
rect 10260 3723 10266 3788
rect 10220 3716 10266 3723
rect 10220 3655 10226 3716
rect 10260 3655 10266 3716
rect 10220 3644 10266 3655
rect 10220 3587 10226 3644
rect 10260 3587 10266 3644
rect 10220 3572 10266 3587
rect 10220 3519 10226 3572
rect 10260 3519 10266 3572
rect 10220 3500 10266 3519
rect 9082 3465 9128 3466
rect 9082 3431 9088 3465
rect 9122 3431 9128 3465
rect 9082 3428 9128 3431
rect 9082 3363 9088 3428
rect 9122 3363 9128 3428
rect 9082 3356 9128 3363
rect 9198 3453 9214 3473
rect 9248 3453 9264 3473
rect 9198 3415 9264 3453
rect 9198 3361 9214 3415
rect 9248 3361 9264 3415
rect 9316 3453 9332 3473
rect 9366 3453 9382 3473
rect 9316 3415 9382 3453
rect 9316 3361 9332 3415
rect 9366 3361 9382 3415
rect 9434 3453 9450 3473
rect 9484 3453 9500 3473
rect 9434 3415 9500 3453
rect 9434 3361 9450 3415
rect 9484 3361 9500 3415
rect 9552 3453 9568 3473
rect 9602 3453 9618 3473
rect 9552 3415 9618 3453
rect 9552 3361 9568 3415
rect 9602 3361 9618 3415
rect 9670 3453 9686 3473
rect 9720 3453 9736 3473
rect 9670 3415 9736 3453
rect 9670 3361 9686 3415
rect 9720 3361 9736 3415
rect 9788 3453 9804 3473
rect 9838 3453 9854 3473
rect 9788 3415 9854 3453
rect 9788 3361 9804 3415
rect 9838 3361 9854 3415
rect 9906 3453 9922 3473
rect 9956 3453 9972 3473
rect 9906 3415 9972 3453
rect 9906 3361 9922 3415
rect 9956 3361 9972 3415
rect 10024 3453 10040 3473
rect 10074 3453 10090 3473
rect 10024 3415 10090 3453
rect 10024 3361 10040 3415
rect 10074 3361 10090 3415
rect 10220 3451 10226 3500
rect 10260 3451 10266 3500
rect 11418 38689 11464 38716
rect 11418 38650 11424 38689
rect 11458 38650 11464 38689
rect 11418 38621 11464 38650
rect 11418 38577 11424 38621
rect 11458 38577 11464 38621
rect 13206 38684 13252 38716
rect 13206 38650 13212 38684
rect 13246 38650 13252 38684
rect 13206 38630 13252 38650
rect 12942 38581 12964 38615
rect 12998 38581 13026 38615
rect 13060 38612 13076 38615
rect 11418 38553 11464 38577
rect 11418 38504 11424 38553
rect 11458 38504 11464 38553
rect 11418 38485 11464 38504
rect 13010 38578 13038 38581
rect 13072 38578 13076 38612
rect 13010 38517 13076 38578
rect 13010 38494 13038 38517
rect 11418 38431 11424 38485
rect 11458 38431 11464 38485
rect 13072 38494 13076 38517
rect 13206 38577 13212 38630
rect 13246 38577 13252 38630
rect 14934 38689 14980 38716
rect 14934 38650 14940 38689
rect 14974 38650 14980 38689
rect 14934 38621 14980 38650
rect 13206 38562 13252 38577
rect 13206 38504 13212 38562
rect 13246 38504 13252 38562
rect 13206 38494 13252 38504
rect 13382 38612 13398 38615
rect 13382 38578 13392 38612
rect 13432 38581 13466 38615
rect 13500 38581 13516 38615
rect 13426 38578 13448 38581
rect 13382 38517 13448 38578
rect 13382 38494 13392 38517
rect 11418 38417 11464 38431
rect 11418 38358 11424 38417
rect 11458 38358 11464 38417
rect 11418 38349 11464 38358
rect 11418 38285 11424 38349
rect 11458 38285 11464 38349
rect 11418 38281 11464 38285
rect 11418 38247 11424 38281
rect 11458 38247 11464 38281
rect 11418 38246 11464 38247
rect 11418 38179 11424 38246
rect 11458 38179 11464 38246
rect 11418 38173 11464 38179
rect 11418 38111 11424 38173
rect 11458 38111 11464 38173
rect 11418 38100 11464 38111
rect 11418 38043 11424 38100
rect 11458 38043 11464 38100
rect 11418 38027 11464 38043
rect 11418 37975 11424 38027
rect 11458 37975 11464 38027
rect 11418 37954 11464 37975
rect 11418 37907 11424 37954
rect 11458 37907 11464 37954
rect 11418 37881 11464 37907
rect 11418 37839 11424 37881
rect 11458 37839 11464 37881
rect 11418 37808 11464 37839
rect 11418 37771 11424 37808
rect 11458 37771 11464 37808
rect 11418 37737 11464 37771
rect 11418 37701 11424 37737
rect 11458 37701 11464 37737
rect 11418 37669 11464 37701
rect 11418 37628 11424 37669
rect 11458 37628 11464 37669
rect 11418 37601 11464 37628
rect 11418 37555 11424 37601
rect 11458 37555 11464 37601
rect 11418 37533 11464 37555
rect 11418 37482 11424 37533
rect 11458 37482 11464 37533
rect 11418 37465 11464 37482
rect 11418 37409 11424 37465
rect 11458 37409 11464 37465
rect 11418 37397 11464 37409
rect 11418 37336 11424 37397
rect 11458 37336 11464 37397
rect 11418 37329 11464 37336
rect 11418 37263 11424 37329
rect 11458 37263 11464 37329
rect 11418 37261 11464 37263
rect 11418 37227 11424 37261
rect 11458 37227 11464 37261
rect 11418 37224 11464 37227
rect 11418 37159 11424 37224
rect 11458 37159 11464 37224
rect 11418 37151 11464 37159
rect 11418 37091 11424 37151
rect 11458 37091 11464 37151
rect 11418 37078 11464 37091
rect 11418 37023 11424 37078
rect 11458 37023 11464 37078
rect 11418 37005 11464 37023
rect 11418 36955 11424 37005
rect 11458 36955 11464 37005
rect 11418 36932 11464 36955
rect 11418 36887 11424 36932
rect 11458 36887 11464 36932
rect 11418 36859 11464 36887
rect 11418 36819 11424 36859
rect 11458 36819 11464 36859
rect 11418 36786 11464 36819
rect 11418 36751 11424 36786
rect 11458 36751 11464 36786
rect 11418 36717 11464 36751
rect 11418 36679 11424 36717
rect 11458 36679 11464 36717
rect 11418 36649 11464 36679
rect 11418 36606 11424 36649
rect 11458 36606 11464 36649
rect 11418 36581 11464 36606
rect 11418 36533 11424 36581
rect 11458 36533 11464 36581
rect 11418 36513 11464 36533
rect 11418 36460 11424 36513
rect 11458 36460 11464 36513
rect 11418 36445 11464 36460
rect 11418 36387 11424 36445
rect 11458 36387 11464 36445
rect 11418 36377 11464 36387
rect 11418 36314 11424 36377
rect 11458 36314 11464 36377
rect 11418 36309 11464 36314
rect 11418 36207 11424 36309
rect 11458 36207 11464 36309
rect 11418 36202 11464 36207
rect 11418 36139 11424 36202
rect 11458 36139 11464 36202
rect 11418 36129 11464 36139
rect 11418 36071 11424 36129
rect 11458 36071 11464 36129
rect 11418 36056 11464 36071
rect 11418 36003 11424 36056
rect 11458 36003 11464 36056
rect 11418 35983 11464 36003
rect 11418 35935 11424 35983
rect 11458 35935 11464 35983
rect 11418 35910 11464 35935
rect 11418 35867 11424 35910
rect 11458 35867 11464 35910
rect 11418 35837 11464 35867
rect 11418 35799 11424 35837
rect 11458 35799 11464 35837
rect 11418 35765 11464 35799
rect 11418 35730 11424 35765
rect 11458 35730 11464 35765
rect 11418 35697 11464 35730
rect 11418 35657 11424 35697
rect 11458 35657 11464 35697
rect 11418 35629 11464 35657
rect 11418 35584 11424 35629
rect 11458 35584 11464 35629
rect 11418 35561 11464 35584
rect 11418 35511 11424 35561
rect 11458 35511 11464 35561
rect 11418 35493 11464 35511
rect 11418 35438 11424 35493
rect 11458 35438 11464 35493
rect 11418 35425 11464 35438
rect 11418 35365 11424 35425
rect 11458 35365 11464 35425
rect 11418 35357 11464 35365
rect 11418 35292 11424 35357
rect 11458 35292 11464 35357
rect 11418 35289 11464 35292
rect 11418 35255 11424 35289
rect 11458 35255 11464 35289
rect 11418 35253 11464 35255
rect 11418 35187 11424 35253
rect 11458 35187 11464 35253
rect 11418 35180 11464 35187
rect 11418 35119 11424 35180
rect 11458 35119 11464 35180
rect 11418 35108 11464 35119
rect 11418 35051 11424 35108
rect 11458 35051 11464 35108
rect 11418 35036 11464 35051
rect 11418 34983 11424 35036
rect 11458 34983 11464 35036
rect 11418 34964 11464 34983
rect 11418 34915 11424 34964
rect 11458 34915 11464 34964
rect 11418 34892 11464 34915
rect 11418 34847 11424 34892
rect 11458 34847 11464 34892
rect 11418 34820 11464 34847
rect 11418 34779 11424 34820
rect 11458 34779 11464 34820
rect 11418 34748 11464 34779
rect 11418 34711 11424 34748
rect 11458 34711 11464 34748
rect 11418 34677 11464 34711
rect 11418 34642 11424 34677
rect 11458 34642 11464 34677
rect 11418 34609 11464 34642
rect 11418 34570 11424 34609
rect 11458 34570 11464 34609
rect 11418 34541 11464 34570
rect 11418 34498 11424 34541
rect 11458 34498 11464 34541
rect 11418 34473 11464 34498
rect 11418 34426 11424 34473
rect 11458 34426 11464 34473
rect 11418 34405 11464 34426
rect 11418 34354 11424 34405
rect 11458 34354 11464 34405
rect 11418 34337 11464 34354
rect 11418 34282 11424 34337
rect 11458 34282 11464 34337
rect 11418 34269 11464 34282
rect 11418 34210 11424 34269
rect 11458 34210 11464 34269
rect 11418 34201 11464 34210
rect 11418 34138 11424 34201
rect 11458 34138 11464 34201
rect 11418 34133 11464 34138
rect 11418 34066 11424 34133
rect 11458 34066 11464 34133
rect 11418 34065 11464 34066
rect 11418 34031 11424 34065
rect 11458 34031 11464 34065
rect 11418 34028 11464 34031
rect 11418 33963 11424 34028
rect 11458 33963 11464 34028
rect 11418 33956 11464 33963
rect 11418 33895 11424 33956
rect 11458 33895 11464 33956
rect 11418 33884 11464 33895
rect 11418 33827 11424 33884
rect 11458 33827 11464 33884
rect 11418 33812 11464 33827
rect 11418 33759 11424 33812
rect 11458 33759 11464 33812
rect 11418 33740 11464 33759
rect 11418 33691 11424 33740
rect 11458 33691 11464 33740
rect 11418 33668 11464 33691
rect 11418 33623 11424 33668
rect 11458 33623 11464 33668
rect 11418 33596 11464 33623
rect 11418 33555 11424 33596
rect 11458 33555 11464 33596
rect 11418 33524 11464 33555
rect 11418 33487 11424 33524
rect 11458 33487 11464 33524
rect 11418 33453 11464 33487
rect 11418 33418 11424 33453
rect 11458 33418 11464 33453
rect 11418 33385 11464 33418
rect 11418 33346 11424 33385
rect 11458 33346 11464 33385
rect 11418 33317 11464 33346
rect 11418 33274 11424 33317
rect 11458 33274 11464 33317
rect 11418 33249 11464 33274
rect 11418 33202 11424 33249
rect 11458 33202 11464 33249
rect 11418 33181 11464 33202
rect 11418 33130 11424 33181
rect 11458 33130 11464 33181
rect 11418 33113 11464 33130
rect 11418 33058 11424 33113
rect 11458 33058 11464 33113
rect 11418 33045 11464 33058
rect 11418 32986 11424 33045
rect 11458 32986 11464 33045
rect 11418 32977 11464 32986
rect 11418 32914 11424 32977
rect 11458 32914 11464 32977
rect 11418 32909 11464 32914
rect 11418 32842 11424 32909
rect 11458 32842 11464 32909
rect 11418 32841 11464 32842
rect 11418 32807 11424 32841
rect 11458 32807 11464 32841
rect 11418 32804 11464 32807
rect 11418 32739 11424 32804
rect 11458 32739 11464 32804
rect 11418 32732 11464 32739
rect 11418 32671 11424 32732
rect 11458 32671 11464 32732
rect 11418 32660 11464 32671
rect 11418 32603 11424 32660
rect 11458 32603 11464 32660
rect 11418 32588 11464 32603
rect 11418 32535 11424 32588
rect 11458 32535 11464 32588
rect 11418 32516 11464 32535
rect 11418 32467 11424 32516
rect 11458 32467 11464 32516
rect 11418 32444 11464 32467
rect 11418 32399 11424 32444
rect 11458 32399 11464 32444
rect 11418 32372 11464 32399
rect 11418 32331 11424 32372
rect 11458 32331 11464 32372
rect 11418 32300 11464 32331
rect 11418 32263 11424 32300
rect 11458 32263 11464 32300
rect 11418 32229 11464 32263
rect 11418 32194 11424 32229
rect 11458 32194 11464 32229
rect 11418 32161 11464 32194
rect 11418 32122 11424 32161
rect 11458 32122 11464 32161
rect 11418 32093 11464 32122
rect 11418 32050 11424 32093
rect 11458 32050 11464 32093
rect 11418 32025 11464 32050
rect 11418 31978 11424 32025
rect 11458 31978 11464 32025
rect 11418 31957 11464 31978
rect 11418 31906 11424 31957
rect 11458 31906 11464 31957
rect 11418 31889 11464 31906
rect 11418 31834 11424 31889
rect 11458 31834 11464 31889
rect 11418 31821 11464 31834
rect 11418 31762 11424 31821
rect 11458 31762 11464 31821
rect 11418 31753 11464 31762
rect 11418 31690 11424 31753
rect 11458 31690 11464 31753
rect 11418 31685 11464 31690
rect 11418 31618 11424 31685
rect 11458 31618 11464 31685
rect 11418 31617 11464 31618
rect 11418 31583 11424 31617
rect 11458 31583 11464 31617
rect 11418 31580 11464 31583
rect 11418 31515 11424 31580
rect 11458 31515 11464 31580
rect 11418 31508 11464 31515
rect 11418 31447 11424 31508
rect 11458 31447 11464 31508
rect 11418 31436 11464 31447
rect 11418 31379 11424 31436
rect 11458 31379 11464 31436
rect 11418 31364 11464 31379
rect 11418 31311 11424 31364
rect 11458 31311 11464 31364
rect 11418 31292 11464 31311
rect 11418 31243 11424 31292
rect 11458 31243 11464 31292
rect 11418 31220 11464 31243
rect 11418 31175 11424 31220
rect 11458 31175 11464 31220
rect 11418 31148 11464 31175
rect 11418 31107 11424 31148
rect 11458 31107 11464 31148
rect 11418 31076 11464 31107
rect 11418 31039 11424 31076
rect 11458 31039 11464 31076
rect 11418 31005 11464 31039
rect 11418 30970 11424 31005
rect 11458 30970 11464 31005
rect 11418 30937 11464 30970
rect 11418 30898 11424 30937
rect 11458 30898 11464 30937
rect 11418 30869 11464 30898
rect 11418 30826 11424 30869
rect 11458 30826 11464 30869
rect 11418 30801 11464 30826
rect 11418 30754 11424 30801
rect 11458 30754 11464 30801
rect 11418 30733 11464 30754
rect 11418 30682 11424 30733
rect 11458 30682 11464 30733
rect 11418 30665 11464 30682
rect 11418 30610 11424 30665
rect 11458 30610 11464 30665
rect 11418 30597 11464 30610
rect 11418 30538 11424 30597
rect 11458 30538 11464 30597
rect 11418 30529 11464 30538
rect 11418 30466 11424 30529
rect 11458 30466 11464 30529
rect 11418 30461 11464 30466
rect 11418 30394 11424 30461
rect 11458 30394 11464 30461
rect 11418 30393 11464 30394
rect 11418 30359 11424 30393
rect 11458 30359 11464 30393
rect 11418 30356 11464 30359
rect 11418 30291 11424 30356
rect 11458 30291 11464 30356
rect 11418 30284 11464 30291
rect 11418 30223 11424 30284
rect 11458 30223 11464 30284
rect 11418 30212 11464 30223
rect 11418 30155 11424 30212
rect 11458 30155 11464 30212
rect 11418 30140 11464 30155
rect 11418 30087 11424 30140
rect 11458 30087 11464 30140
rect 11418 30068 11464 30087
rect 11418 30019 11424 30068
rect 11458 30019 11464 30068
rect 11418 29996 11464 30019
rect 11418 29951 11424 29996
rect 11458 29951 11464 29996
rect 11418 29924 11464 29951
rect 11418 29883 11424 29924
rect 11458 29883 11464 29924
rect 11418 29852 11464 29883
rect 11418 29815 11424 29852
rect 11458 29815 11464 29852
rect 11418 29781 11464 29815
rect 11418 29746 11424 29781
rect 11458 29746 11464 29781
rect 11418 29713 11464 29746
rect 11418 29674 11424 29713
rect 11458 29674 11464 29713
rect 11418 29645 11464 29674
rect 11418 29602 11424 29645
rect 11458 29602 11464 29645
rect 11418 29577 11464 29602
rect 11418 29530 11424 29577
rect 11458 29530 11464 29577
rect 11418 29509 11464 29530
rect 11418 29458 11424 29509
rect 11458 29458 11464 29509
rect 11418 29441 11464 29458
rect 11418 29386 11424 29441
rect 11458 29386 11464 29441
rect 11418 29373 11464 29386
rect 11418 29314 11424 29373
rect 11458 29314 11464 29373
rect 11418 29305 11464 29314
rect 11418 29242 11424 29305
rect 11458 29242 11464 29305
rect 11418 29237 11464 29242
rect 11418 29170 11424 29237
rect 11458 29170 11464 29237
rect 11418 29169 11464 29170
rect 11418 29135 11424 29169
rect 11458 29135 11464 29169
rect 11418 29132 11464 29135
rect 11418 29067 11424 29132
rect 11458 29067 11464 29132
rect 11418 29060 11464 29067
rect 11418 28999 11424 29060
rect 11458 28999 11464 29060
rect 11418 28988 11464 28999
rect 11418 28931 11424 28988
rect 11458 28931 11464 28988
rect 11418 28916 11464 28931
rect 11418 28863 11424 28916
rect 11458 28863 11464 28916
rect 11418 28844 11464 28863
rect 11418 28795 11424 28844
rect 11458 28795 11464 28844
rect 11418 28772 11464 28795
rect 11418 28727 11424 28772
rect 11458 28727 11464 28772
rect 11418 28700 11464 28727
rect 11418 28659 11424 28700
rect 11458 28659 11464 28700
rect 11418 28628 11464 28659
rect 11418 28591 11424 28628
rect 11458 28591 11464 28628
rect 11418 28557 11464 28591
rect 11418 28522 11424 28557
rect 11458 28522 11464 28557
rect 11418 28489 11464 28522
rect 11418 28450 11424 28489
rect 11458 28450 11464 28489
rect 11418 28421 11464 28450
rect 11418 28378 11424 28421
rect 11458 28378 11464 28421
rect 11418 28353 11464 28378
rect 11418 28306 11424 28353
rect 11458 28306 11464 28353
rect 11418 28285 11464 28306
rect 11418 28234 11424 28285
rect 11458 28234 11464 28285
rect 11418 28217 11464 28234
rect 11418 28162 11424 28217
rect 11458 28162 11464 28217
rect 11418 28149 11464 28162
rect 11418 28090 11424 28149
rect 11458 28090 11464 28149
rect 11418 28081 11464 28090
rect 11418 28018 11424 28081
rect 11458 28018 11464 28081
rect 11418 28013 11464 28018
rect 11418 27946 11424 28013
rect 11458 27946 11464 28013
rect 11418 27945 11464 27946
rect 11418 27911 11424 27945
rect 11458 27911 11464 27945
rect 11418 27908 11464 27911
rect 11418 27843 11424 27908
rect 11458 27843 11464 27908
rect 11418 27836 11464 27843
rect 11418 27775 11424 27836
rect 11458 27775 11464 27836
rect 11418 27764 11464 27775
rect 11418 27707 11424 27764
rect 11458 27707 11464 27764
rect 11418 27692 11464 27707
rect 11418 27639 11424 27692
rect 11458 27639 11464 27692
rect 11418 27620 11464 27639
rect 11418 27571 11424 27620
rect 11458 27571 11464 27620
rect 11418 27548 11464 27571
rect 11418 27503 11424 27548
rect 11458 27503 11464 27548
rect 11418 27476 11464 27503
rect 11418 27435 11424 27476
rect 11458 27435 11464 27476
rect 11418 27404 11464 27435
rect 11418 27367 11424 27404
rect 11458 27367 11464 27404
rect 11418 27333 11464 27367
rect 11418 27298 11424 27333
rect 11458 27298 11464 27333
rect 11418 27265 11464 27298
rect 11418 27226 11424 27265
rect 11458 27226 11464 27265
rect 11418 27197 11464 27226
rect 11418 27154 11424 27197
rect 11458 27154 11464 27197
rect 11418 27129 11464 27154
rect 11418 27082 11424 27129
rect 11458 27082 11464 27129
rect 11418 27061 11464 27082
rect 11418 27010 11424 27061
rect 11458 27010 11464 27061
rect 11418 26993 11464 27010
rect 11418 26938 11424 26993
rect 11458 26938 11464 26993
rect 11418 26925 11464 26938
rect 11418 26866 11424 26925
rect 11458 26866 11464 26925
rect 11418 26857 11464 26866
rect 11418 26794 11424 26857
rect 11458 26794 11464 26857
rect 11418 26789 11464 26794
rect 11418 26722 11424 26789
rect 11458 26722 11464 26789
rect 11418 26721 11464 26722
rect 11418 26687 11424 26721
rect 11458 26687 11464 26721
rect 11418 26684 11464 26687
rect 11418 26619 11424 26684
rect 11458 26619 11464 26684
rect 11418 26612 11464 26619
rect 11418 26551 11424 26612
rect 11458 26551 11464 26612
rect 11418 26540 11464 26551
rect 11418 26483 11424 26540
rect 11458 26483 11464 26540
rect 11418 26468 11464 26483
rect 11418 26415 11424 26468
rect 11458 26415 11464 26468
rect 11418 26396 11464 26415
rect 11418 26347 11424 26396
rect 11458 26347 11464 26396
rect 11418 26324 11464 26347
rect 11418 26279 11424 26324
rect 11458 26279 11464 26324
rect 11418 26252 11464 26279
rect 11418 26211 11424 26252
rect 11458 26211 11464 26252
rect 11418 26180 11464 26211
rect 11418 26143 11424 26180
rect 11458 26143 11464 26180
rect 11418 26109 11464 26143
rect 11418 26074 11424 26109
rect 11458 26074 11464 26109
rect 11418 26041 11464 26074
rect 11418 26002 11424 26041
rect 11458 26002 11464 26041
rect 11418 25973 11464 26002
rect 11418 25930 11424 25973
rect 11458 25930 11464 25973
rect 11418 25905 11464 25930
rect 11418 25858 11424 25905
rect 11458 25858 11464 25905
rect 11418 25837 11464 25858
rect 11418 25786 11424 25837
rect 11458 25786 11464 25837
rect 11418 25769 11464 25786
rect 11418 25714 11424 25769
rect 11458 25714 11464 25769
rect 11418 25701 11464 25714
rect 11418 25642 11424 25701
rect 11458 25642 11464 25701
rect 11418 25633 11464 25642
rect 11418 25570 11424 25633
rect 11458 25570 11464 25633
rect 11418 25565 11464 25570
rect 11418 25498 11424 25565
rect 11458 25498 11464 25565
rect 11418 25497 11464 25498
rect 11418 25463 11424 25497
rect 11458 25463 11464 25497
rect 11418 25460 11464 25463
rect 11418 25395 11424 25460
rect 11458 25395 11464 25460
rect 11418 25388 11464 25395
rect 11418 25327 11424 25388
rect 11458 25327 11464 25388
rect 11418 25316 11464 25327
rect 11418 25259 11424 25316
rect 11458 25259 11464 25316
rect 11418 25244 11464 25259
rect 11418 25191 11424 25244
rect 11458 25191 11464 25244
rect 11418 25172 11464 25191
rect 11418 25123 11424 25172
rect 11458 25123 11464 25172
rect 11418 25100 11464 25123
rect 11418 25055 11424 25100
rect 11458 25055 11464 25100
rect 11418 25028 11464 25055
rect 11418 24987 11424 25028
rect 11458 24987 11464 25028
rect 11418 24956 11464 24987
rect 11418 24919 11424 24956
rect 11458 24919 11464 24956
rect 11418 24885 11464 24919
rect 11418 24850 11424 24885
rect 11458 24850 11464 24885
rect 11418 24817 11464 24850
rect 11418 24778 11424 24817
rect 11458 24778 11464 24817
rect 11418 24749 11464 24778
rect 11418 24706 11424 24749
rect 11458 24706 11464 24749
rect 11418 24681 11464 24706
rect 11418 24634 11424 24681
rect 11458 24634 11464 24681
rect 11418 24613 11464 24634
rect 11418 24562 11424 24613
rect 11458 24562 11464 24613
rect 11418 24545 11464 24562
rect 11418 24490 11424 24545
rect 11458 24490 11464 24545
rect 11418 24477 11464 24490
rect 11418 24418 11424 24477
rect 11458 24418 11464 24477
rect 11418 24409 11464 24418
rect 11418 24346 11424 24409
rect 11458 24346 11464 24409
rect 11418 24341 11464 24346
rect 11418 24274 11424 24341
rect 11458 24274 11464 24341
rect 11418 24273 11464 24274
rect 11418 24239 11424 24273
rect 11458 24239 11464 24273
rect 11418 24236 11464 24239
rect 11418 24171 11424 24236
rect 11458 24171 11464 24236
rect 11418 24164 11464 24171
rect 11418 24103 11424 24164
rect 11458 24103 11464 24164
rect 11418 24092 11464 24103
rect 11418 24035 11424 24092
rect 11458 24035 11464 24092
rect 11418 24020 11464 24035
rect 11418 23967 11424 24020
rect 11458 23967 11464 24020
rect 11418 23948 11464 23967
rect 11418 23899 11424 23948
rect 11458 23899 11464 23948
rect 11418 23876 11464 23899
rect 11418 23831 11424 23876
rect 11458 23831 11464 23876
rect 11418 23804 11464 23831
rect 11418 23763 11424 23804
rect 11458 23763 11464 23804
rect 11418 23732 11464 23763
rect 11418 23695 11424 23732
rect 11458 23695 11464 23732
rect 11418 23661 11464 23695
rect 11418 23626 11424 23661
rect 11458 23626 11464 23661
rect 11418 23593 11464 23626
rect 11418 23554 11424 23593
rect 11458 23554 11464 23593
rect 11418 23525 11464 23554
rect 11418 23482 11424 23525
rect 11458 23482 11464 23525
rect 11418 23457 11464 23482
rect 11418 23410 11424 23457
rect 11458 23410 11464 23457
rect 11418 23389 11464 23410
rect 11418 23338 11424 23389
rect 11458 23338 11464 23389
rect 11418 23321 11464 23338
rect 11418 23266 11424 23321
rect 11458 23266 11464 23321
rect 11418 23253 11464 23266
rect 11418 23194 11424 23253
rect 11458 23194 11464 23253
rect 11418 23185 11464 23194
rect 11418 23122 11424 23185
rect 11458 23122 11464 23185
rect 11418 23117 11464 23122
rect 11418 23050 11424 23117
rect 11458 23050 11464 23117
rect 11418 23049 11464 23050
rect 11418 23015 11424 23049
rect 11458 23015 11464 23049
rect 11418 23012 11464 23015
rect 11418 22947 11424 23012
rect 11458 22947 11464 23012
rect 11418 22940 11464 22947
rect 11418 22879 11424 22940
rect 11458 22879 11464 22940
rect 11418 22868 11464 22879
rect 11418 22811 11424 22868
rect 11458 22811 11464 22868
rect 11418 22796 11464 22811
rect 11418 22743 11424 22796
rect 11458 22743 11464 22796
rect 11418 22724 11464 22743
rect 11418 22675 11424 22724
rect 11458 22675 11464 22724
rect 11418 22652 11464 22675
rect 11418 22607 11424 22652
rect 11458 22607 11464 22652
rect 11418 22580 11464 22607
rect 11418 22539 11424 22580
rect 11458 22539 11464 22580
rect 11418 22508 11464 22539
rect 11418 22471 11424 22508
rect 11458 22471 11464 22508
rect 11418 22437 11464 22471
rect 11418 22402 11424 22437
rect 11458 22402 11464 22437
rect 11418 22369 11464 22402
rect 11418 22330 11424 22369
rect 11458 22330 11464 22369
rect 11418 22301 11464 22330
rect 11418 22258 11424 22301
rect 11458 22258 11464 22301
rect 11418 22233 11464 22258
rect 11418 22186 11424 22233
rect 11458 22186 11464 22233
rect 11418 22165 11464 22186
rect 11418 22114 11424 22165
rect 11458 22114 11464 22165
rect 11418 22097 11464 22114
rect 11418 22042 11424 22097
rect 11458 22042 11464 22097
rect 11418 22029 11464 22042
rect 11418 21970 11424 22029
rect 11458 21970 11464 22029
rect 11418 21961 11464 21970
rect 11418 21898 11424 21961
rect 11458 21898 11464 21961
rect 11418 21893 11464 21898
rect 11418 21826 11424 21893
rect 11458 21826 11464 21893
rect 11418 21825 11464 21826
rect 11418 21791 11424 21825
rect 11458 21791 11464 21825
rect 11418 21788 11464 21791
rect 11418 21723 11424 21788
rect 11458 21723 11464 21788
rect 11418 21716 11464 21723
rect 11418 21655 11424 21716
rect 11458 21655 11464 21716
rect 11418 21644 11464 21655
rect 11418 21587 11424 21644
rect 11458 21587 11464 21644
rect 11418 21572 11464 21587
rect 11418 21519 11424 21572
rect 11458 21519 11464 21572
rect 11418 21500 11464 21519
rect 11418 21451 11424 21500
rect 11458 21451 11464 21500
rect 11418 21428 11464 21451
rect 11418 21383 11424 21428
rect 11458 21383 11464 21428
rect 11418 21356 11464 21383
rect 11418 21315 11424 21356
rect 11458 21315 11464 21356
rect 11418 21284 11464 21315
rect 11418 21247 11424 21284
rect 11458 21247 11464 21284
rect 11418 21213 11464 21247
rect 11418 21178 11424 21213
rect 11458 21178 11464 21213
rect 11418 21145 11464 21178
rect 11418 21106 11424 21145
rect 11458 21106 11464 21145
rect 11418 21077 11464 21106
rect 11418 21034 11424 21077
rect 11458 21034 11464 21077
rect 11418 21009 11464 21034
rect 11418 20962 11424 21009
rect 11458 20962 11464 21009
rect 11418 20941 11464 20962
rect 11418 20890 11424 20941
rect 11458 20890 11464 20941
rect 11418 20873 11464 20890
rect 11418 20818 11424 20873
rect 11458 20818 11464 20873
rect 11418 20805 11464 20818
rect 11418 20746 11424 20805
rect 11458 20746 11464 20805
rect 11418 20737 11464 20746
rect 11418 20674 11424 20737
rect 11458 20674 11464 20737
rect 11418 20669 11464 20674
rect 11418 20602 11424 20669
rect 11458 20602 11464 20669
rect 11418 20601 11464 20602
rect 11418 20567 11424 20601
rect 11458 20567 11464 20601
rect 11418 20564 11464 20567
rect 11418 20499 11424 20564
rect 11458 20499 11464 20564
rect 11418 20492 11464 20499
rect 11418 20431 11424 20492
rect 11458 20431 11464 20492
rect 11418 20420 11464 20431
rect 11418 20363 11424 20420
rect 11458 20363 11464 20420
rect 11418 20348 11464 20363
rect 11418 20295 11424 20348
rect 11458 20295 11464 20348
rect 11418 20276 11464 20295
rect 11418 20227 11424 20276
rect 11458 20227 11464 20276
rect 11418 20204 11464 20227
rect 11418 20159 11424 20204
rect 11458 20159 11464 20204
rect 11418 20132 11464 20159
rect 11418 20091 11424 20132
rect 11458 20091 11464 20132
rect 11418 20060 11464 20091
rect 11418 20023 11424 20060
rect 11458 20023 11464 20060
rect 11418 19989 11464 20023
rect 11418 19954 11424 19989
rect 11458 19954 11464 19989
rect 11418 19921 11464 19954
rect 11418 19882 11424 19921
rect 11458 19882 11464 19921
rect 11418 19853 11464 19882
rect 11418 19810 11424 19853
rect 11458 19810 11464 19853
rect 11418 19785 11464 19810
rect 11418 19738 11424 19785
rect 11458 19738 11464 19785
rect 11418 19717 11464 19738
rect 11418 19666 11424 19717
rect 11458 19666 11464 19717
rect 11418 19649 11464 19666
rect 11418 19594 11424 19649
rect 11458 19594 11464 19649
rect 11418 19581 11464 19594
rect 11418 19522 11424 19581
rect 11458 19522 11464 19581
rect 11418 19513 11464 19522
rect 11418 19450 11424 19513
rect 11458 19450 11464 19513
rect 11418 19445 11464 19450
rect 11418 19378 11424 19445
rect 11458 19378 11464 19445
rect 11418 19377 11464 19378
rect 11418 19343 11424 19377
rect 11458 19343 11464 19377
rect 11418 19340 11464 19343
rect 11418 19275 11424 19340
rect 11458 19275 11464 19340
rect 11418 19268 11464 19275
rect 11418 19207 11424 19268
rect 11458 19207 11464 19268
rect 11418 19196 11464 19207
rect 11418 19139 11424 19196
rect 11458 19139 11464 19196
rect 11418 19124 11464 19139
rect 11418 19071 11424 19124
rect 11458 19071 11464 19124
rect 11418 19052 11464 19071
rect 11418 19003 11424 19052
rect 11458 19003 11464 19052
rect 11418 18980 11464 19003
rect 11418 18935 11424 18980
rect 11458 18935 11464 18980
rect 11418 18908 11464 18935
rect 11418 18867 11424 18908
rect 11458 18867 11464 18908
rect 11418 18836 11464 18867
rect 11418 18799 11424 18836
rect 11458 18799 11464 18836
rect 11418 18765 11464 18799
rect 11418 18730 11424 18765
rect 11458 18730 11464 18765
rect 11418 18697 11464 18730
rect 11418 18658 11424 18697
rect 11458 18658 11464 18697
rect 11418 18629 11464 18658
rect 11418 18586 11424 18629
rect 11458 18586 11464 18629
rect 11418 18561 11464 18586
rect 11418 18514 11424 18561
rect 11458 18514 11464 18561
rect 11418 18493 11464 18514
rect 11418 18442 11424 18493
rect 11458 18442 11464 18493
rect 11418 18425 11464 18442
rect 11418 18370 11424 18425
rect 11458 18370 11464 18425
rect 11418 18357 11464 18370
rect 11418 18298 11424 18357
rect 11458 18298 11464 18357
rect 11418 18289 11464 18298
rect 11418 18226 11424 18289
rect 11458 18226 11464 18289
rect 11418 18221 11464 18226
rect 11418 18154 11424 18221
rect 11458 18154 11464 18221
rect 11418 18153 11464 18154
rect 11418 18119 11424 18153
rect 11458 18119 11464 18153
rect 11418 18116 11464 18119
rect 11418 18051 11424 18116
rect 11458 18051 11464 18116
rect 11418 18044 11464 18051
rect 11418 17983 11424 18044
rect 11458 17983 11464 18044
rect 11418 17972 11464 17983
rect 11418 17915 11424 17972
rect 11458 17915 11464 17972
rect 11418 17900 11464 17915
rect 11418 17847 11424 17900
rect 11458 17847 11464 17900
rect 11418 17828 11464 17847
rect 11418 17779 11424 17828
rect 11458 17779 11464 17828
rect 11418 17756 11464 17779
rect 11418 17711 11424 17756
rect 11458 17711 11464 17756
rect 11418 17684 11464 17711
rect 11418 17643 11424 17684
rect 11458 17643 11464 17684
rect 11418 17612 11464 17643
rect 11418 17575 11424 17612
rect 11458 17575 11464 17612
rect 11418 17541 11464 17575
rect 11418 17506 11424 17541
rect 11458 17506 11464 17541
rect 11418 17473 11464 17506
rect 11418 17434 11424 17473
rect 11458 17434 11464 17473
rect 11418 17405 11464 17434
rect 11418 17362 11424 17405
rect 11458 17362 11464 17405
rect 11418 17337 11464 17362
rect 11418 17290 11424 17337
rect 11458 17290 11464 17337
rect 11418 17269 11464 17290
rect 11418 17218 11424 17269
rect 11458 17218 11464 17269
rect 11418 17201 11464 17218
rect 11418 17146 11424 17201
rect 11458 17146 11464 17201
rect 11418 17133 11464 17146
rect 11418 17074 11424 17133
rect 11458 17074 11464 17133
rect 11418 17065 11464 17074
rect 11418 17002 11424 17065
rect 11458 17002 11464 17065
rect 11418 16997 11464 17002
rect 11418 16930 11424 16997
rect 11458 16930 11464 16997
rect 11418 16929 11464 16930
rect 11418 16895 11424 16929
rect 11458 16895 11464 16929
rect 11418 16892 11464 16895
rect 11418 16827 11424 16892
rect 11458 16827 11464 16892
rect 11418 16820 11464 16827
rect 11418 16759 11424 16820
rect 11458 16759 11464 16820
rect 11418 16748 11464 16759
rect 11418 16691 11424 16748
rect 11458 16691 11464 16748
rect 11418 16676 11464 16691
rect 11418 16623 11424 16676
rect 11458 16623 11464 16676
rect 11418 16604 11464 16623
rect 11418 16555 11424 16604
rect 11458 16555 11464 16604
rect 11418 16532 11464 16555
rect 11418 16487 11424 16532
rect 11458 16487 11464 16532
rect 11418 16460 11464 16487
rect 11418 16419 11424 16460
rect 11458 16419 11464 16460
rect 11418 16388 11464 16419
rect 11418 16351 11424 16388
rect 11458 16351 11464 16388
rect 11418 16317 11464 16351
rect 11418 16282 11424 16317
rect 11458 16282 11464 16317
rect 11418 16249 11464 16282
rect 11418 16210 11424 16249
rect 11458 16210 11464 16249
rect 11418 16181 11464 16210
rect 11418 16138 11424 16181
rect 11458 16138 11464 16181
rect 11418 16113 11464 16138
rect 11418 16066 11424 16113
rect 11458 16066 11464 16113
rect 11418 16045 11464 16066
rect 11418 15994 11424 16045
rect 11458 15994 11464 16045
rect 11418 15977 11464 15994
rect 11418 15922 11424 15977
rect 11458 15922 11464 15977
rect 11418 15909 11464 15922
rect 11418 15850 11424 15909
rect 11458 15850 11464 15909
rect 11418 15841 11464 15850
rect 11418 15778 11424 15841
rect 11458 15778 11464 15841
rect 11418 15773 11464 15778
rect 11418 15706 11424 15773
rect 11458 15706 11464 15773
rect 11418 15705 11464 15706
rect 11418 15671 11424 15705
rect 11458 15671 11464 15705
rect 11418 15668 11464 15671
rect 11418 15603 11424 15668
rect 11458 15603 11464 15668
rect 11418 15596 11464 15603
rect 11418 15535 11424 15596
rect 11458 15535 11464 15596
rect 11418 15524 11464 15535
rect 11418 15467 11424 15524
rect 11458 15467 11464 15524
rect 11418 15452 11464 15467
rect 11418 15399 11424 15452
rect 11458 15399 11464 15452
rect 11418 15380 11464 15399
rect 11418 15331 11424 15380
rect 11458 15331 11464 15380
rect 11418 15308 11464 15331
rect 11418 15263 11424 15308
rect 11458 15263 11464 15308
rect 11418 15236 11464 15263
rect 11418 15195 11424 15236
rect 11458 15195 11464 15236
rect 11418 15164 11464 15195
rect 11418 15127 11424 15164
rect 11458 15127 11464 15164
rect 11418 15093 11464 15127
rect 11418 15058 11424 15093
rect 11458 15058 11464 15093
rect 11418 15025 11464 15058
rect 11418 14986 11424 15025
rect 11458 14986 11464 15025
rect 11418 14957 11464 14986
rect 11418 14914 11424 14957
rect 11458 14914 11464 14957
rect 11418 14889 11464 14914
rect 11418 14842 11424 14889
rect 11458 14842 11464 14889
rect 11418 14821 11464 14842
rect 11418 14770 11424 14821
rect 11458 14770 11464 14821
rect 11418 14753 11464 14770
rect 11418 14698 11424 14753
rect 11458 14698 11464 14753
rect 11418 14685 11464 14698
rect 11418 14626 11424 14685
rect 11458 14626 11464 14685
rect 11418 14617 11464 14626
rect 11418 14554 11424 14617
rect 11458 14554 11464 14617
rect 11418 14549 11464 14554
rect 11418 14482 11424 14549
rect 11458 14482 11464 14549
rect 11418 14481 11464 14482
rect 11418 14447 11424 14481
rect 11458 14447 11464 14481
rect 11418 14444 11464 14447
rect 11418 14379 11424 14444
rect 11458 14379 11464 14444
rect 11418 14372 11464 14379
rect 11418 14311 11424 14372
rect 11458 14311 11464 14372
rect 11418 14300 11464 14311
rect 11418 14243 11424 14300
rect 11458 14243 11464 14300
rect 11418 14228 11464 14243
rect 11418 14175 11424 14228
rect 11458 14175 11464 14228
rect 11418 14156 11464 14175
rect 11418 14107 11424 14156
rect 11458 14107 11464 14156
rect 11418 14084 11464 14107
rect 11418 14039 11424 14084
rect 11458 14039 11464 14084
rect 11418 14012 11464 14039
rect 11418 13971 11424 14012
rect 11458 13971 11464 14012
rect 11418 13940 11464 13971
rect 11418 13903 11424 13940
rect 11458 13903 11464 13940
rect 11418 13869 11464 13903
rect 11418 13834 11424 13869
rect 11458 13834 11464 13869
rect 11418 13801 11464 13834
rect 11418 13762 11424 13801
rect 11458 13762 11464 13801
rect 11418 13733 11464 13762
rect 11418 13690 11424 13733
rect 11458 13690 11464 13733
rect 11418 13665 11464 13690
rect 11418 13618 11424 13665
rect 11458 13618 11464 13665
rect 11418 13597 11464 13618
rect 11418 13546 11424 13597
rect 11458 13546 11464 13597
rect 11418 13529 11464 13546
rect 11418 13474 11424 13529
rect 11458 13474 11464 13529
rect 11418 13461 11464 13474
rect 11418 13402 11424 13461
rect 11458 13402 11464 13461
rect 11418 13393 11464 13402
rect 11418 13330 11424 13393
rect 11458 13330 11464 13393
rect 11418 13325 11464 13330
rect 11418 13258 11424 13325
rect 11458 13258 11464 13325
rect 11418 13257 11464 13258
rect 11418 13223 11424 13257
rect 11458 13223 11464 13257
rect 11418 13220 11464 13223
rect 11418 13155 11424 13220
rect 11458 13155 11464 13220
rect 11418 13148 11464 13155
rect 11418 13087 11424 13148
rect 11458 13087 11464 13148
rect 11418 13076 11464 13087
rect 11418 13019 11424 13076
rect 11458 13019 11464 13076
rect 11418 13004 11464 13019
rect 11418 12951 11424 13004
rect 11458 12951 11464 13004
rect 11418 12932 11464 12951
rect 11418 12883 11424 12932
rect 11458 12883 11464 12932
rect 11418 12860 11464 12883
rect 11418 12815 11424 12860
rect 11458 12815 11464 12860
rect 11418 12788 11464 12815
rect 11418 12747 11424 12788
rect 11458 12747 11464 12788
rect 11418 12716 11464 12747
rect 11418 12679 11424 12716
rect 11458 12679 11464 12716
rect 11418 12645 11464 12679
rect 11418 12610 11424 12645
rect 11458 12610 11464 12645
rect 11418 12577 11464 12610
rect 11418 12538 11424 12577
rect 11458 12538 11464 12577
rect 11418 12509 11464 12538
rect 11418 12466 11424 12509
rect 11458 12466 11464 12509
rect 11418 12441 11464 12466
rect 11418 12394 11424 12441
rect 11458 12394 11464 12441
rect 11418 12373 11464 12394
rect 11418 12322 11424 12373
rect 11458 12322 11464 12373
rect 11418 12305 11464 12322
rect 11418 12250 11424 12305
rect 11458 12250 11464 12305
rect 11418 12237 11464 12250
rect 11418 12178 11424 12237
rect 11458 12178 11464 12237
rect 11418 12169 11464 12178
rect 11418 12106 11424 12169
rect 11458 12106 11464 12169
rect 11418 12101 11464 12106
rect 11418 12034 11424 12101
rect 11458 12034 11464 12101
rect 11418 12033 11464 12034
rect 11418 11999 11424 12033
rect 11458 11999 11464 12033
rect 11418 11996 11464 11999
rect 11418 11931 11424 11996
rect 11458 11931 11464 11996
rect 11418 11924 11464 11931
rect 11418 11863 11424 11924
rect 11458 11863 11464 11924
rect 11418 11852 11464 11863
rect 11418 11795 11424 11852
rect 11458 11795 11464 11852
rect 11418 11780 11464 11795
rect 11418 11727 11424 11780
rect 11458 11727 11464 11780
rect 11418 11708 11464 11727
rect 11418 11659 11424 11708
rect 11458 11659 11464 11708
rect 11418 11636 11464 11659
rect 11418 11591 11424 11636
rect 11458 11591 11464 11636
rect 11418 11564 11464 11591
rect 11418 11523 11424 11564
rect 11458 11523 11464 11564
rect 11418 11492 11464 11523
rect 11418 11455 11424 11492
rect 11458 11455 11464 11492
rect 11418 11421 11464 11455
rect 11418 11386 11424 11421
rect 11458 11386 11464 11421
rect 11418 11353 11464 11386
rect 11418 11314 11424 11353
rect 11458 11314 11464 11353
rect 11418 11285 11464 11314
rect 11418 11242 11424 11285
rect 11458 11242 11464 11285
rect 11418 11217 11464 11242
rect 11418 11170 11424 11217
rect 11458 11170 11464 11217
rect 11418 11149 11464 11170
rect 11418 11098 11424 11149
rect 11458 11098 11464 11149
rect 11418 11081 11464 11098
rect 11418 11026 11424 11081
rect 11458 11026 11464 11081
rect 11418 11013 11464 11026
rect 11418 10954 11424 11013
rect 11458 10954 11464 11013
rect 11418 10945 11464 10954
rect 11418 10882 11424 10945
rect 11458 10882 11464 10945
rect 11418 10877 11464 10882
rect 11418 10810 11424 10877
rect 11458 10810 11464 10877
rect 11418 10809 11464 10810
rect 11418 10775 11424 10809
rect 11458 10775 11464 10809
rect 11418 10772 11464 10775
rect 11418 10707 11424 10772
rect 11458 10707 11464 10772
rect 11418 10700 11464 10707
rect 11418 10639 11424 10700
rect 11458 10639 11464 10700
rect 11418 10628 11464 10639
rect 11418 10571 11424 10628
rect 11458 10571 11464 10628
rect 11418 10556 11464 10571
rect 11418 10503 11424 10556
rect 11458 10503 11464 10556
rect 11418 10484 11464 10503
rect 11418 10435 11424 10484
rect 11458 10435 11464 10484
rect 11418 10412 11464 10435
rect 11418 10367 11424 10412
rect 11458 10367 11464 10412
rect 11418 10340 11464 10367
rect 11418 10299 11424 10340
rect 11458 10299 11464 10340
rect 11418 10268 11464 10299
rect 11418 10231 11424 10268
rect 11458 10231 11464 10268
rect 11418 10197 11464 10231
rect 11418 10162 11424 10197
rect 11458 10162 11464 10197
rect 11418 10129 11464 10162
rect 11418 10090 11424 10129
rect 11458 10090 11464 10129
rect 11418 10061 11464 10090
rect 11418 10018 11424 10061
rect 11458 10018 11464 10061
rect 11418 9993 11464 10018
rect 11418 9946 11424 9993
rect 11458 9946 11464 9993
rect 11418 9925 11464 9946
rect 11418 9874 11424 9925
rect 11458 9874 11464 9925
rect 11418 9857 11464 9874
rect 11418 9802 11424 9857
rect 11458 9802 11464 9857
rect 11418 9789 11464 9802
rect 11418 9730 11424 9789
rect 11458 9730 11464 9789
rect 11418 9721 11464 9730
rect 11418 9658 11424 9721
rect 11458 9658 11464 9721
rect 11418 9653 11464 9658
rect 11418 9586 11424 9653
rect 11458 9586 11464 9653
rect 11418 9585 11464 9586
rect 11418 9551 11424 9585
rect 11458 9551 11464 9585
rect 11418 9548 11464 9551
rect 11418 9483 11424 9548
rect 11458 9483 11464 9548
rect 11418 9476 11464 9483
rect 11418 9415 11424 9476
rect 11458 9415 11464 9476
rect 11418 9404 11464 9415
rect 11418 9347 11424 9404
rect 11458 9347 11464 9404
rect 11418 9332 11464 9347
rect 11418 9279 11424 9332
rect 11458 9279 11464 9332
rect 11418 9260 11464 9279
rect 11418 9211 11424 9260
rect 11458 9211 11464 9260
rect 11418 9188 11464 9211
rect 11418 9143 11424 9188
rect 11458 9143 11464 9188
rect 11418 9116 11464 9143
rect 11418 9075 11424 9116
rect 11458 9075 11464 9116
rect 11418 9044 11464 9075
rect 11418 9007 11424 9044
rect 11458 9007 11464 9044
rect 11418 8973 11464 9007
rect 11418 8938 11424 8973
rect 11458 8938 11464 8973
rect 11418 8905 11464 8938
rect 11418 8866 11424 8905
rect 11458 8866 11464 8905
rect 11418 8837 11464 8866
rect 11418 8794 11424 8837
rect 11458 8794 11464 8837
rect 11418 8769 11464 8794
rect 11418 8722 11424 8769
rect 11458 8722 11464 8769
rect 11418 8701 11464 8722
rect 11418 8650 11424 8701
rect 11458 8650 11464 8701
rect 11418 8633 11464 8650
rect 11418 8578 11424 8633
rect 11458 8578 11464 8633
rect 11418 8565 11464 8578
rect 11418 8506 11424 8565
rect 11458 8506 11464 8565
rect 11418 8497 11464 8506
rect 11418 8434 11424 8497
rect 11458 8434 11464 8497
rect 11418 8429 11464 8434
rect 11418 8362 11424 8429
rect 11458 8362 11464 8429
rect 11418 8361 11464 8362
rect 11418 8327 11424 8361
rect 11458 8327 11464 8361
rect 11418 8324 11464 8327
rect 11418 8259 11424 8324
rect 11458 8259 11464 8324
rect 11418 8252 11464 8259
rect 11418 8191 11424 8252
rect 11458 8191 11464 8252
rect 11418 8180 11464 8191
rect 11418 8123 11424 8180
rect 11458 8123 11464 8180
rect 11418 8108 11464 8123
rect 11418 8055 11424 8108
rect 11458 8055 11464 8108
rect 11418 8036 11464 8055
rect 11418 7987 11424 8036
rect 11458 7987 11464 8036
rect 11418 7964 11464 7987
rect 11418 7919 11424 7964
rect 11458 7919 11464 7964
rect 11418 7892 11464 7919
rect 11418 7851 11424 7892
rect 11458 7851 11464 7892
rect 11418 7820 11464 7851
rect 11418 7783 11424 7820
rect 11458 7783 11464 7820
rect 11418 7749 11464 7783
rect 11418 7714 11424 7749
rect 11458 7714 11464 7749
rect 11418 7681 11464 7714
rect 11418 7642 11424 7681
rect 11458 7642 11464 7681
rect 11418 7613 11464 7642
rect 11418 7570 11424 7613
rect 11458 7570 11464 7613
rect 11418 7545 11464 7570
rect 11418 7498 11424 7545
rect 11458 7498 11464 7545
rect 11418 7477 11464 7498
rect 11418 7426 11424 7477
rect 11458 7426 11464 7477
rect 11418 7409 11464 7426
rect 11418 7354 11424 7409
rect 11458 7354 11464 7409
rect 11418 7341 11464 7354
rect 11418 7282 11424 7341
rect 11458 7282 11464 7341
rect 11418 7273 11464 7282
rect 11418 7210 11424 7273
rect 11458 7210 11464 7273
rect 11418 7205 11464 7210
rect 11418 7138 11424 7205
rect 11458 7138 11464 7205
rect 11418 7137 11464 7138
rect 11418 7103 11424 7137
rect 11458 7103 11464 7137
rect 11418 7100 11464 7103
rect 11418 7035 11424 7100
rect 11458 7035 11464 7100
rect 11418 7028 11464 7035
rect 11418 6967 11424 7028
rect 11458 6967 11464 7028
rect 11418 6956 11464 6967
rect 11418 6899 11424 6956
rect 11458 6899 11464 6956
rect 11418 6884 11464 6899
rect 11418 6831 11424 6884
rect 11458 6831 11464 6884
rect 11418 6812 11464 6831
rect 11418 6763 11424 6812
rect 11458 6763 11464 6812
rect 11418 6740 11464 6763
rect 11418 6695 11424 6740
rect 11458 6695 11464 6740
rect 11418 6668 11464 6695
rect 11418 6627 11424 6668
rect 11458 6627 11464 6668
rect 11418 6596 11464 6627
rect 11418 6559 11424 6596
rect 11458 6559 11464 6596
rect 11418 6525 11464 6559
rect 11418 6490 11424 6525
rect 11458 6490 11464 6525
rect 11418 6457 11464 6490
rect 11418 6418 11424 6457
rect 11458 6418 11464 6457
rect 11418 6389 11464 6418
rect 11418 6346 11424 6389
rect 11458 6346 11464 6389
rect 11418 6321 11464 6346
rect 11418 6274 11424 6321
rect 11458 6274 11464 6321
rect 11418 6253 11464 6274
rect 11418 6202 11424 6253
rect 11458 6202 11464 6253
rect 11418 6185 11464 6202
rect 11418 6130 11424 6185
rect 11458 6130 11464 6185
rect 11418 6117 11464 6130
rect 11418 6058 11424 6117
rect 11458 6058 11464 6117
rect 11418 6049 11464 6058
rect 11418 5986 11424 6049
rect 11458 5986 11464 6049
rect 11418 5981 11464 5986
rect 11418 5914 11424 5981
rect 11458 5914 11464 5981
rect 11418 5913 11464 5914
rect 11418 5879 11424 5913
rect 11458 5879 11464 5913
rect 11418 5876 11464 5879
rect 11418 5811 11424 5876
rect 11458 5811 11464 5876
rect 11418 5804 11464 5811
rect 11418 5743 11424 5804
rect 11458 5743 11464 5804
rect 11418 5732 11464 5743
rect 11418 5675 11424 5732
rect 11458 5675 11464 5732
rect 11418 5660 11464 5675
rect 11418 5607 11424 5660
rect 11458 5607 11464 5660
rect 11418 5588 11464 5607
rect 11418 5539 11424 5588
rect 11458 5539 11464 5588
rect 11418 5516 11464 5539
rect 11418 5471 11424 5516
rect 11458 5471 11464 5516
rect 11418 5444 11464 5471
rect 11418 5403 11424 5444
rect 11458 5403 11464 5444
rect 11418 5372 11464 5403
rect 11418 5335 11424 5372
rect 11458 5335 11464 5372
rect 11418 5301 11464 5335
rect 11418 5266 11424 5301
rect 11458 5266 11464 5301
rect 11418 5233 11464 5266
rect 11418 5194 11424 5233
rect 11458 5194 11464 5233
rect 11418 5165 11464 5194
rect 11418 5122 11424 5165
rect 11458 5122 11464 5165
rect 11418 5097 11464 5122
rect 11418 5050 11424 5097
rect 11458 5050 11464 5097
rect 11418 5029 11464 5050
rect 11418 4978 11424 5029
rect 11458 4978 11464 5029
rect 11418 4961 11464 4978
rect 11418 4906 11424 4961
rect 11458 4906 11464 4961
rect 11418 4893 11464 4906
rect 11418 4834 11424 4893
rect 11458 4834 11464 4893
rect 11418 4825 11464 4834
rect 11418 4762 11424 4825
rect 11458 4762 11464 4825
rect 11418 4757 11464 4762
rect 11418 4690 11424 4757
rect 11458 4690 11464 4757
rect 11418 4689 11464 4690
rect 11418 4655 11424 4689
rect 11458 4655 11464 4689
rect 11418 4652 11464 4655
rect 11418 4587 11424 4652
rect 11458 4587 11464 4652
rect 11418 4580 11464 4587
rect 11418 4519 11424 4580
rect 11458 4519 11464 4580
rect 11418 4508 11464 4519
rect 11418 4451 11424 4508
rect 11458 4451 11464 4508
rect 11418 4436 11464 4451
rect 11418 4383 11424 4436
rect 11458 4383 11464 4436
rect 11418 4364 11464 4383
rect 11418 4315 11424 4364
rect 11458 4315 11464 4364
rect 11418 4292 11464 4315
rect 11418 4247 11424 4292
rect 11458 4247 11464 4292
rect 11418 4220 11464 4247
rect 11418 4179 11424 4220
rect 11458 4179 11464 4220
rect 11418 4148 11464 4179
rect 11418 4111 11424 4148
rect 11458 4111 11464 4148
rect 11418 4077 11464 4111
rect 11418 4042 11424 4077
rect 11458 4042 11464 4077
rect 11418 4009 11464 4042
rect 11418 3970 11424 4009
rect 11458 3970 11464 4009
rect 11418 3941 11464 3970
rect 11418 3898 11424 3941
rect 11458 3898 11464 3941
rect 11418 3873 11464 3898
rect 11418 3826 11424 3873
rect 11458 3826 11464 3873
rect 11418 3805 11464 3826
rect 11418 3754 11424 3805
rect 11458 3754 11464 3805
rect 11418 3737 11464 3754
rect 11418 3682 11424 3737
rect 11458 3682 11464 3737
rect 11418 3669 11464 3682
rect 11418 3610 11424 3669
rect 11458 3610 11464 3669
rect 11418 3601 11464 3610
rect 11418 3538 11424 3601
rect 11458 3538 11464 3601
rect 11418 3533 11464 3538
rect 10220 3428 10266 3451
rect 10220 3383 10226 3428
rect 10260 3383 10266 3428
rect 9082 3295 9088 3356
rect 9122 3295 9128 3356
rect 9082 3284 9128 3295
rect 9082 3250 9088 3284
rect 9122 3250 9128 3284
rect 9082 3218 9128 3250
rect 10220 3356 10266 3383
rect 10396 3453 10412 3473
rect 10446 3453 10462 3473
rect 10396 3415 10462 3453
rect 10396 3361 10412 3415
rect 10446 3361 10462 3415
rect 10514 3453 10530 3473
rect 10564 3453 10580 3473
rect 10514 3415 10580 3453
rect 10514 3361 10530 3415
rect 10564 3361 10580 3415
rect 10632 3453 10648 3473
rect 10682 3453 10698 3473
rect 10632 3415 10698 3453
rect 10632 3361 10648 3415
rect 10682 3361 10698 3415
rect 10750 3453 10766 3473
rect 10800 3453 10816 3473
rect 10750 3415 10816 3453
rect 10750 3361 10766 3415
rect 10800 3361 10816 3415
rect 10868 3453 10884 3473
rect 10918 3453 10934 3473
rect 10868 3415 10934 3453
rect 10868 3361 10884 3415
rect 10918 3361 10934 3415
rect 10986 3453 11002 3473
rect 11036 3453 11052 3473
rect 10986 3415 11052 3453
rect 10986 3361 11002 3415
rect 11036 3361 11052 3415
rect 11104 3453 11120 3473
rect 11154 3453 11170 3473
rect 11104 3415 11170 3453
rect 11104 3361 11120 3415
rect 11154 3361 11170 3415
rect 11222 3453 11238 3473
rect 11272 3453 11288 3473
rect 11222 3415 11288 3453
rect 11222 3361 11238 3415
rect 11272 3361 11288 3415
rect 11418 3466 11424 3533
rect 11458 3466 11464 3533
rect 11418 3465 11464 3466
rect 11418 3431 11424 3465
rect 11458 3431 11464 3465
rect 11418 3428 11464 3431
rect 11418 3363 11424 3428
rect 11458 3363 11464 3428
rect 10220 3315 10226 3356
rect 10260 3315 10266 3356
rect 10220 3284 10266 3315
rect 10220 3247 10226 3284
rect 10260 3247 10266 3284
rect 10220 3218 10266 3247
rect 11418 3356 11464 3363
rect 11418 3295 11424 3356
rect 11458 3295 11464 3356
rect 11418 3284 11464 3295
rect 11418 3250 11424 3284
rect 11458 3250 11464 3284
rect 11418 3218 11464 3250
rect 9082 3213 11464 3218
rect 9082 3179 9156 3213
rect 9190 3212 9224 3213
rect 9258 3212 9292 3213
rect 9326 3212 9360 3213
rect 9394 3212 9428 3213
rect 9462 3212 9496 3213
rect 9530 3212 9564 3213
rect 9194 3179 9224 3212
rect 9268 3179 9292 3212
rect 9341 3179 9360 3212
rect 9414 3179 9428 3212
rect 9487 3179 9496 3212
rect 9560 3179 9564 3212
rect 9598 3212 9632 3213
rect 9666 3212 9700 3213
rect 9734 3212 9768 3213
rect 9802 3212 9836 3213
rect 9870 3212 9904 3213
rect 9938 3212 9972 3213
rect 10006 3212 10040 3213
rect 9598 3179 9599 3212
rect 9666 3179 9672 3212
rect 9734 3179 9745 3212
rect 9802 3179 9818 3212
rect 9870 3179 9891 3212
rect 9938 3179 9964 3212
rect 10006 3179 10037 3212
rect 10074 3179 10108 3213
rect 10142 3212 10336 3213
rect 10370 3212 10404 3213
rect 9082 3178 9160 3179
rect 9194 3178 9234 3179
rect 9268 3178 9307 3179
rect 9341 3178 9380 3179
rect 9414 3178 9453 3179
rect 9487 3178 9526 3179
rect 9560 3178 9599 3179
rect 9633 3178 9672 3179
rect 9706 3178 9745 3179
rect 9779 3178 9818 3179
rect 9852 3178 9891 3179
rect 9925 3178 9964 3179
rect 9998 3178 10037 3179
rect 10071 3178 10110 3179
rect 10144 3178 10183 3212
rect 10217 3178 10256 3212
rect 10290 3178 10329 3212
rect 10370 3179 10402 3212
rect 10438 3179 10472 3213
rect 10506 3212 10540 3213
rect 10574 3212 10608 3213
rect 10642 3212 10676 3213
rect 10710 3212 10744 3213
rect 10778 3212 10812 3213
rect 10846 3212 10880 3213
rect 10914 3212 10948 3213
rect 10509 3179 10540 3212
rect 10582 3179 10608 3212
rect 10655 3179 10676 3212
rect 10728 3179 10744 3212
rect 10801 3179 10812 3212
rect 10874 3179 10880 3212
rect 10947 3179 10948 3212
rect 10982 3212 11016 3213
rect 11050 3212 11084 3213
rect 11118 3212 11152 3213
rect 11186 3212 11220 3213
rect 11254 3212 11288 3213
rect 11322 3212 11356 3213
rect 10982 3179 10986 3212
rect 11050 3179 11059 3212
rect 11118 3179 11132 3212
rect 11186 3179 11205 3212
rect 11254 3179 11278 3212
rect 11322 3179 11351 3212
rect 11390 3205 11464 3213
rect 11390 3179 11424 3205
rect 10363 3178 10402 3179
rect 10436 3178 10475 3179
rect 10509 3178 10548 3179
rect 10582 3178 10621 3179
rect 10655 3178 10694 3179
rect 10728 3178 10767 3179
rect 10801 3178 10840 3179
rect 10874 3178 10913 3179
rect 10947 3178 10986 3179
rect 11020 3178 11059 3179
rect 11093 3178 11132 3179
rect 11166 3178 11205 3179
rect 11239 3178 11278 3179
rect 11312 3178 11351 3179
rect 11385 3178 11424 3179
rect 9082 3172 11424 3178
rect 11418 3171 11424 3172
rect 11458 3171 11464 3205
rect 11418 3140 11464 3171
rect 11418 3103 11424 3140
rect 11458 3103 11464 3140
rect 11418 3069 11464 3103
rect 11418 3033 11424 3069
rect 11458 3033 11464 3069
rect 11418 3001 11464 3033
rect 11418 2960 11424 3001
rect 11458 2960 11464 3001
rect 11418 2933 11464 2960
rect 11418 2887 11424 2933
rect 11458 2887 11464 2933
rect 11418 2865 11464 2887
rect 11418 2814 11424 2865
rect 11458 2814 11464 2865
rect 11418 2797 11464 2814
rect 11418 2741 11424 2797
rect 11458 2741 11464 2797
rect 11418 2729 11464 2741
rect 11418 2668 11424 2729
rect 11458 2668 11464 2729
rect 11418 2661 11464 2668
rect 5452 2561 5500 2595
rect 5534 2561 5583 2595
rect 5617 2561 5666 2595
rect 5700 2561 5749 2595
rect 5783 2561 5832 2595
rect 5940 2589 5974 2602
rect 5184 2549 5218 2550
rect 5184 2476 5218 2500
rect 5940 2515 5974 2534
rect 5940 2441 5974 2466
rect 5184 2403 5218 2431
rect 5312 2405 5357 2439
rect 5391 2405 5436 2439
rect 5470 2405 5515 2439
rect 5549 2405 5595 2439
rect 5629 2405 5675 2439
rect 5709 2405 5755 2439
rect 5184 2330 5218 2362
rect 5184 2258 5218 2293
rect 5940 2367 5974 2398
rect 5940 2296 5974 2330
rect 5452 2249 5500 2283
rect 5534 2249 5583 2283
rect 5617 2249 5666 2283
rect 5700 2249 5749 2283
rect 5783 2249 5832 2283
rect 5184 2189 5218 2223
rect 5184 2120 5218 2150
rect 5940 2228 5974 2259
rect 5940 2160 5974 2185
rect 5312 2093 5357 2127
rect 5391 2093 5436 2127
rect 5470 2093 5515 2127
rect 5549 2093 5595 2127
rect 5629 2093 5675 2127
rect 5709 2093 5755 2127
rect 5184 2051 5218 2077
rect 5184 1982 5218 2004
rect 5940 2092 5974 2111
rect 5940 2024 5974 2037
rect 5452 1937 5500 1971
rect 5534 1937 5583 1971
rect 5617 1937 5666 1971
rect 5700 1937 5749 1971
rect 5783 1937 5832 1971
rect 5940 1956 5974 1963
rect 5184 1913 5218 1931
rect 5184 1844 5218 1858
rect 5940 1888 5974 1889
rect 5940 1849 5974 1854
rect 5184 1776 5218 1785
rect 5312 1781 5357 1815
rect 5391 1781 5436 1815
rect 5470 1781 5515 1815
rect 5549 1781 5595 1815
rect 5629 1781 5675 1815
rect 5709 1781 5755 1815
rect 5184 1708 5218 1712
rect 5184 1673 5218 1674
rect 5940 1775 5974 1786
rect 5940 1701 5974 1718
rect 5452 1625 5500 1659
rect 5534 1625 5583 1659
rect 5617 1625 5666 1659
rect 5700 1625 5749 1659
rect 5783 1625 5832 1659
rect 5940 1627 5974 1650
rect 5184 1600 5218 1606
rect 5184 1527 5218 1538
rect 5940 1553 5974 1582
rect 5184 1454 5218 1470
rect 5312 1469 5357 1503
rect 5391 1469 5436 1503
rect 5470 1469 5515 1503
rect 5549 1469 5595 1503
rect 5629 1469 5675 1503
rect 5709 1469 5755 1503
rect 5940 1480 5974 1514
rect 5184 1381 5218 1402
rect 5940 1412 5974 1445
rect 5184 1308 5218 1334
rect 5452 1313 5500 1347
rect 5534 1313 5583 1347
rect 5617 1313 5666 1347
rect 5700 1313 5749 1347
rect 5783 1313 5832 1347
rect 5940 1344 5974 1372
rect 5184 1236 5218 1266
rect 5184 1164 5218 1198
rect 5940 1276 5974 1299
rect 5940 1208 5974 1226
rect 5312 1157 5357 1191
rect 5391 1157 5436 1191
rect 5470 1157 5515 1191
rect 5549 1157 5595 1191
rect 5629 1157 5675 1191
rect 5709 1157 5755 1191
rect 5184 1096 5218 1130
rect 5184 1046 5218 1058
rect 5940 1140 5974 1153
rect 5940 1072 5974 1080
rect 5452 1001 5500 1035
rect 5534 1001 5583 1035
rect 5617 1001 5666 1035
rect 5700 1001 5749 1035
rect 5783 1001 5832 1035
rect 5940 994 5974 1007
rect 11418 2595 11424 2661
rect 11458 2595 11464 2661
rect 11418 2593 11464 2595
rect 11418 2559 11424 2593
rect 11458 2559 11464 2593
rect 11418 2556 11464 2559
rect 11418 2491 11424 2556
rect 11458 2491 11464 2556
rect 11418 2483 11464 2491
rect 11418 2423 11424 2483
rect 11458 2423 11464 2483
rect 11418 2410 11464 2423
rect 11418 2355 11424 2410
rect 11458 2355 11464 2410
rect 11418 2337 11464 2355
rect 11418 2287 11424 2337
rect 11458 2287 11464 2337
rect 11418 2264 11464 2287
rect 11418 2219 11424 2264
rect 11458 2219 11464 2264
rect 11418 2191 11464 2219
rect 11418 2151 11424 2191
rect 11458 2151 11464 2191
rect 11418 2118 11464 2151
rect 11418 2083 11424 2118
rect 11458 2083 11464 2118
rect 11418 2049 11464 2083
rect 11418 2011 11424 2049
rect 11458 2011 11464 2049
rect 11418 1981 11464 2011
rect 11418 1938 11424 1981
rect 11458 1938 11464 1981
rect 11418 1913 11464 1938
rect 11418 1865 11424 1913
rect 11458 1865 11464 1913
rect 11418 1845 11464 1865
rect 11418 1792 11424 1845
rect 11458 1792 11464 1845
rect 11418 1777 11464 1792
rect 11418 1719 11424 1777
rect 11458 1719 11464 1777
rect 11418 1709 11464 1719
rect 11418 1646 11424 1709
rect 11458 1646 11464 1709
rect 11418 1641 11464 1646
rect 11418 1539 11424 1641
rect 11458 1539 11464 1641
rect 11418 1534 11464 1539
rect 11418 1471 11424 1534
rect 11458 1471 11464 1534
rect 11418 1461 11464 1471
rect 11418 1403 11424 1461
rect 11458 1403 11464 1461
rect 11418 1388 11464 1403
rect 11418 1335 11424 1388
rect 11458 1335 11464 1388
rect 11418 1315 11464 1335
rect 11418 1267 11424 1315
rect 11458 1267 11464 1315
rect 11418 1242 11464 1267
rect 11418 1199 11424 1242
rect 11458 1199 11464 1242
rect 11418 1169 11464 1199
rect 11418 1131 11424 1169
rect 11458 1131 11464 1169
rect 11418 1097 11464 1131
rect 11418 1062 11424 1097
rect 11458 1062 11464 1097
rect 11418 1029 11464 1062
rect 11418 989 11424 1029
rect 11458 989 11464 1029
rect 11418 961 11464 989
rect 11418 916 11424 961
rect 11458 916 11464 961
rect 11418 893 11464 916
rect 11418 843 11424 893
rect 11458 843 11464 893
rect 11418 825 11464 843
rect 11418 770 11424 825
rect 11458 770 11464 825
rect 11418 757 11464 770
rect 11418 697 11424 757
rect 11458 697 11464 757
rect 11418 689 11464 697
rect 11418 624 11424 689
rect 11458 624 11464 689
rect 11418 621 11464 624
rect 11418 587 11424 621
rect 11458 587 11464 621
rect 11418 585 11464 587
rect 11418 519 11424 585
rect 11458 519 11464 585
rect 11418 512 11464 519
rect 11418 451 11424 512
rect 11458 451 11464 512
rect 11418 439 11464 451
rect 11418 383 11424 439
rect 11458 383 11464 439
rect 13206 38431 13212 38494
rect 13246 38431 13252 38494
rect 13426 38494 13448 38517
rect 14934 38578 14940 38621
rect 14974 38578 14980 38621
rect 14934 38553 14980 38578
rect 14934 38506 14940 38553
rect 14974 38506 14980 38553
rect 14934 38485 14980 38506
rect 13206 38426 13252 38431
rect 13206 38324 13212 38426
rect 13246 38324 13252 38426
rect 13206 38319 13252 38324
rect 13206 38256 13212 38319
rect 13246 38256 13252 38319
rect 13206 38246 13252 38256
rect 13206 38188 13212 38246
rect 13246 38188 13252 38246
rect 13206 38173 13252 38188
rect 13206 38120 13212 38173
rect 13246 38120 13252 38173
rect 13206 38100 13252 38120
rect 13206 38052 13212 38100
rect 13246 38052 13252 38100
rect 13206 38027 13252 38052
rect 13206 37984 13212 38027
rect 13246 37984 13252 38027
rect 13206 37954 13252 37984
rect 13206 37916 13212 37954
rect 13246 37916 13252 37954
rect 13206 37882 13252 37916
rect 13206 37847 13212 37882
rect 13246 37847 13252 37882
rect 13206 37814 13252 37847
rect 13206 37774 13212 37814
rect 13246 37774 13252 37814
rect 13206 37746 13252 37774
rect 13206 37701 13212 37746
rect 13246 37701 13252 37746
rect 13206 37678 13252 37701
rect 13206 37628 13212 37678
rect 13246 37628 13252 37678
rect 13206 37610 13252 37628
rect 13206 37555 13212 37610
rect 13246 37555 13252 37610
rect 13206 37542 13252 37555
rect 13206 37482 13212 37542
rect 13246 37482 13252 37542
rect 13206 37474 13252 37482
rect 13206 37409 13212 37474
rect 13246 37409 13252 37474
rect 13206 37406 13252 37409
rect 13206 37372 13212 37406
rect 13246 37372 13252 37406
rect 13206 37370 13252 37372
rect 13206 37304 13212 37370
rect 13246 37304 13252 37370
rect 13206 37298 13252 37304
rect 13206 37236 13212 37298
rect 13246 37236 13252 37298
rect 13206 37226 13252 37236
rect 13206 37168 13212 37226
rect 13246 37168 13252 37226
rect 13206 37154 13252 37168
rect 13206 37100 13212 37154
rect 13246 37100 13252 37154
rect 13206 37082 13252 37100
rect 13206 37032 13212 37082
rect 13246 37032 13252 37082
rect 13206 37010 13252 37032
rect 13206 36964 13212 37010
rect 13246 36964 13252 37010
rect 13206 36938 13252 36964
rect 13206 36896 13212 36938
rect 13246 36896 13252 36938
rect 13206 36866 13252 36896
rect 13206 36828 13212 36866
rect 13246 36828 13252 36866
rect 13206 36794 13252 36828
rect 13206 36760 13212 36794
rect 13246 36760 13252 36794
rect 13206 36726 13252 36760
rect 13206 36688 13212 36726
rect 13246 36688 13252 36726
rect 13206 36658 13252 36688
rect 13206 36616 13212 36658
rect 13246 36616 13252 36658
rect 13206 36590 13252 36616
rect 13206 36544 13212 36590
rect 13246 36544 13252 36590
rect 13206 36522 13252 36544
rect 13206 36472 13212 36522
rect 13246 36472 13252 36522
rect 13206 36454 13252 36472
rect 13206 36400 13212 36454
rect 13246 36400 13252 36454
rect 13206 36386 13252 36400
rect 13206 36328 13212 36386
rect 13246 36328 13252 36386
rect 13206 36318 13252 36328
rect 13206 36256 13212 36318
rect 13246 36256 13252 36318
rect 13206 36250 13252 36256
rect 13206 36184 13212 36250
rect 13246 36184 13252 36250
rect 13206 36182 13252 36184
rect 13206 36148 13212 36182
rect 13246 36148 13252 36182
rect 13206 36146 13252 36148
rect 13206 36080 13212 36146
rect 13246 36080 13252 36146
rect 13206 36074 13252 36080
rect 13206 36012 13212 36074
rect 13246 36012 13252 36074
rect 13206 36002 13252 36012
rect 13206 35944 13212 36002
rect 13246 35944 13252 36002
rect 13206 35930 13252 35944
rect 13206 35876 13212 35930
rect 13246 35876 13252 35930
rect 13206 35858 13252 35876
rect 13206 35808 13212 35858
rect 13246 35808 13252 35858
rect 13206 35786 13252 35808
rect 13206 35740 13212 35786
rect 13246 35740 13252 35786
rect 13206 35714 13252 35740
rect 13206 35672 13212 35714
rect 13246 35672 13252 35714
rect 13206 35642 13252 35672
rect 13206 35604 13212 35642
rect 13246 35604 13252 35642
rect 13206 35570 13252 35604
rect 13206 35536 13212 35570
rect 13246 35536 13252 35570
rect 13206 35502 13252 35536
rect 13206 35464 13212 35502
rect 13246 35464 13252 35502
rect 13206 35434 13252 35464
rect 13206 35392 13212 35434
rect 13246 35392 13252 35434
rect 13206 35366 13252 35392
rect 13206 35320 13212 35366
rect 13246 35320 13252 35366
rect 13206 35298 13252 35320
rect 13206 35248 13212 35298
rect 13246 35248 13252 35298
rect 13206 35230 13252 35248
rect 13206 35176 13212 35230
rect 13246 35176 13252 35230
rect 13206 35162 13252 35176
rect 13206 35104 13212 35162
rect 13246 35104 13252 35162
rect 13206 35094 13252 35104
rect 13206 35032 13212 35094
rect 13246 35032 13252 35094
rect 13206 35026 13252 35032
rect 13206 34960 13212 35026
rect 13246 34960 13252 35026
rect 13206 34958 13252 34960
rect 13206 34924 13212 34958
rect 13246 34924 13252 34958
rect 13206 34922 13252 34924
rect 13206 34856 13212 34922
rect 13246 34856 13252 34922
rect 13206 34850 13252 34856
rect 13206 34788 13212 34850
rect 13246 34788 13252 34850
rect 13206 34778 13252 34788
rect 13206 34720 13212 34778
rect 13246 34720 13252 34778
rect 13206 34706 13252 34720
rect 13206 34652 13212 34706
rect 13246 34652 13252 34706
rect 13206 34634 13252 34652
rect 13206 34584 13212 34634
rect 13246 34584 13252 34634
rect 13206 34562 13252 34584
rect 13206 34516 13212 34562
rect 13246 34516 13252 34562
rect 13206 34490 13252 34516
rect 13206 34448 13212 34490
rect 13246 34448 13252 34490
rect 13206 34418 13252 34448
rect 13206 34380 13212 34418
rect 13246 34380 13252 34418
rect 13206 34346 13252 34380
rect 13206 34312 13212 34346
rect 13246 34312 13252 34346
rect 13206 34278 13252 34312
rect 13206 34240 13212 34278
rect 13246 34240 13252 34278
rect 13206 34210 13252 34240
rect 13206 34168 13212 34210
rect 13246 34168 13252 34210
rect 13206 34142 13252 34168
rect 13206 34096 13212 34142
rect 13246 34096 13252 34142
rect 13206 34074 13252 34096
rect 13206 34024 13212 34074
rect 13246 34024 13252 34074
rect 13206 34006 13252 34024
rect 13206 33952 13212 34006
rect 13246 33952 13252 34006
rect 13206 33938 13252 33952
rect 13206 33880 13212 33938
rect 13246 33880 13252 33938
rect 13206 33870 13252 33880
rect 13206 33808 13212 33870
rect 13246 33808 13252 33870
rect 13206 33802 13252 33808
rect 13206 33736 13212 33802
rect 13246 33736 13252 33802
rect 13206 33734 13252 33736
rect 13206 33700 13212 33734
rect 13246 33700 13252 33734
rect 13206 33698 13252 33700
rect 13206 33632 13212 33698
rect 13246 33632 13252 33698
rect 13206 33626 13252 33632
rect 13206 33564 13212 33626
rect 13246 33564 13252 33626
rect 13206 33554 13252 33564
rect 13206 33496 13212 33554
rect 13246 33496 13252 33554
rect 13206 33482 13252 33496
rect 13206 33428 13212 33482
rect 13246 33428 13252 33482
rect 13206 33410 13252 33428
rect 13206 33360 13212 33410
rect 13246 33360 13252 33410
rect 13206 33338 13252 33360
rect 13206 33292 13212 33338
rect 13246 33292 13252 33338
rect 13206 33266 13252 33292
rect 13206 33224 13212 33266
rect 13246 33224 13252 33266
rect 13206 33194 13252 33224
rect 13206 33156 13212 33194
rect 13246 33156 13252 33194
rect 13206 33122 13252 33156
rect 13206 33088 13212 33122
rect 13246 33088 13252 33122
rect 13206 33054 13252 33088
rect 13206 33016 13212 33054
rect 13246 33016 13252 33054
rect 13206 32986 13252 33016
rect 13206 32944 13212 32986
rect 13246 32944 13252 32986
rect 13206 32918 13252 32944
rect 13206 32872 13212 32918
rect 13246 32872 13252 32918
rect 13206 32850 13252 32872
rect 13206 32800 13212 32850
rect 13246 32800 13252 32850
rect 13206 32782 13252 32800
rect 13206 32728 13212 32782
rect 13246 32728 13252 32782
rect 13206 32714 13252 32728
rect 13206 32656 13212 32714
rect 13246 32656 13252 32714
rect 13206 32646 13252 32656
rect 13206 32584 13212 32646
rect 13246 32584 13252 32646
rect 13206 32578 13252 32584
rect 13206 32512 13212 32578
rect 13246 32512 13252 32578
rect 13206 32510 13252 32512
rect 13206 32476 13212 32510
rect 13246 32476 13252 32510
rect 13206 32474 13252 32476
rect 13206 32408 13212 32474
rect 13246 32408 13252 32474
rect 13206 32402 13252 32408
rect 13206 32340 13212 32402
rect 13246 32340 13252 32402
rect 13206 32330 13252 32340
rect 13206 32272 13212 32330
rect 13246 32272 13252 32330
rect 13206 32258 13252 32272
rect 13206 32204 13212 32258
rect 13246 32204 13252 32258
rect 13206 32186 13252 32204
rect 13206 32136 13212 32186
rect 13246 32136 13252 32186
rect 13206 32114 13252 32136
rect 13206 32068 13212 32114
rect 13246 32068 13252 32114
rect 13206 32042 13252 32068
rect 13206 32000 13212 32042
rect 13246 32000 13252 32042
rect 13206 31970 13252 32000
rect 13206 31932 13212 31970
rect 13246 31932 13252 31970
rect 13206 31898 13252 31932
rect 13206 31864 13212 31898
rect 13246 31864 13252 31898
rect 13206 31830 13252 31864
rect 13206 31792 13212 31830
rect 13246 31792 13252 31830
rect 13206 31762 13252 31792
rect 13206 31720 13212 31762
rect 13246 31720 13252 31762
rect 13206 31694 13252 31720
rect 13206 31648 13212 31694
rect 13246 31648 13252 31694
rect 13206 31626 13252 31648
rect 13206 31576 13212 31626
rect 13246 31576 13252 31626
rect 13206 31558 13252 31576
rect 13206 31504 13212 31558
rect 13246 31504 13252 31558
rect 13206 31490 13252 31504
rect 13206 31432 13212 31490
rect 13246 31432 13252 31490
rect 13206 31422 13252 31432
rect 13206 31360 13212 31422
rect 13246 31360 13252 31422
rect 13206 31354 13252 31360
rect 13206 31288 13212 31354
rect 13246 31288 13252 31354
rect 13206 31286 13252 31288
rect 13206 31252 13212 31286
rect 13246 31252 13252 31286
rect 13206 31250 13252 31252
rect 13206 31184 13212 31250
rect 13246 31184 13252 31250
rect 13206 31178 13252 31184
rect 13206 31116 13212 31178
rect 13246 31116 13252 31178
rect 13206 31106 13252 31116
rect 13206 31048 13212 31106
rect 13246 31048 13252 31106
rect 13206 31034 13252 31048
rect 13206 30980 13212 31034
rect 13246 30980 13252 31034
rect 13206 30962 13252 30980
rect 13206 30912 13212 30962
rect 13246 30912 13252 30962
rect 13206 30890 13252 30912
rect 13206 30844 13212 30890
rect 13246 30844 13252 30890
rect 13206 30818 13252 30844
rect 13206 30776 13212 30818
rect 13246 30776 13252 30818
rect 13206 30746 13252 30776
rect 13206 30708 13212 30746
rect 13246 30708 13252 30746
rect 13206 30674 13252 30708
rect 13206 30640 13212 30674
rect 13246 30640 13252 30674
rect 13206 30606 13252 30640
rect 13206 30568 13212 30606
rect 13246 30568 13252 30606
rect 13206 30538 13252 30568
rect 13206 30496 13212 30538
rect 13246 30496 13252 30538
rect 13206 30470 13252 30496
rect 13206 30424 13212 30470
rect 13246 30424 13252 30470
rect 13206 30402 13252 30424
rect 13206 30352 13212 30402
rect 13246 30352 13252 30402
rect 13206 30334 13252 30352
rect 13206 30280 13212 30334
rect 13246 30280 13252 30334
rect 13206 30266 13252 30280
rect 13206 30208 13212 30266
rect 13246 30208 13252 30266
rect 13206 30198 13252 30208
rect 13206 30136 13212 30198
rect 13246 30136 13252 30198
rect 13206 30130 13252 30136
rect 13206 30064 13212 30130
rect 13246 30064 13252 30130
rect 13206 30062 13252 30064
rect 13206 30028 13212 30062
rect 13246 30028 13252 30062
rect 13206 30026 13252 30028
rect 13206 29960 13212 30026
rect 13246 29960 13252 30026
rect 13206 29954 13252 29960
rect 13206 29892 13212 29954
rect 13246 29892 13252 29954
rect 13206 29882 13252 29892
rect 13206 29824 13212 29882
rect 13246 29824 13252 29882
rect 13206 29810 13252 29824
rect 13206 29756 13212 29810
rect 13246 29756 13252 29810
rect 13206 29738 13252 29756
rect 13206 29688 13212 29738
rect 13246 29688 13252 29738
rect 13206 29666 13252 29688
rect 13206 29620 13212 29666
rect 13246 29620 13252 29666
rect 13206 29594 13252 29620
rect 13206 29552 13212 29594
rect 13246 29552 13252 29594
rect 13206 29522 13252 29552
rect 13206 29484 13212 29522
rect 13246 29484 13252 29522
rect 13206 29450 13252 29484
rect 13206 29416 13212 29450
rect 13246 29416 13252 29450
rect 13206 29382 13252 29416
rect 13206 29344 13212 29382
rect 13246 29344 13252 29382
rect 13206 29314 13252 29344
rect 13206 29272 13212 29314
rect 13246 29272 13252 29314
rect 13206 29246 13252 29272
rect 13206 29200 13212 29246
rect 13246 29200 13252 29246
rect 13206 29178 13252 29200
rect 13206 29128 13212 29178
rect 13246 29128 13252 29178
rect 13206 29110 13252 29128
rect 13206 29056 13212 29110
rect 13246 29056 13252 29110
rect 13206 29042 13252 29056
rect 13206 28984 13212 29042
rect 13246 28984 13252 29042
rect 13206 28974 13252 28984
rect 13206 28912 13212 28974
rect 13246 28912 13252 28974
rect 13206 28906 13252 28912
rect 13206 28840 13212 28906
rect 13246 28840 13252 28906
rect 13206 28838 13252 28840
rect 13206 28804 13212 28838
rect 13246 28804 13252 28838
rect 13206 28802 13252 28804
rect 13206 28736 13212 28802
rect 13246 28736 13252 28802
rect 13206 28730 13252 28736
rect 13206 28668 13212 28730
rect 13246 28668 13252 28730
rect 13206 28658 13252 28668
rect 13206 28600 13212 28658
rect 13246 28600 13252 28658
rect 13206 28586 13252 28600
rect 13206 28532 13212 28586
rect 13246 28532 13252 28586
rect 13206 28514 13252 28532
rect 13206 28464 13212 28514
rect 13246 28464 13252 28514
rect 13206 28442 13252 28464
rect 13206 28396 13212 28442
rect 13246 28396 13252 28442
rect 13206 28370 13252 28396
rect 13206 28328 13212 28370
rect 13246 28328 13252 28370
rect 13206 28298 13252 28328
rect 13206 28260 13212 28298
rect 13246 28260 13252 28298
rect 13206 28226 13252 28260
rect 13206 28192 13212 28226
rect 13246 28192 13252 28226
rect 13206 28158 13252 28192
rect 13206 28120 13212 28158
rect 13246 28120 13252 28158
rect 13206 28090 13252 28120
rect 13206 28048 13212 28090
rect 13246 28048 13252 28090
rect 13206 28022 13252 28048
rect 13206 27976 13212 28022
rect 13246 27976 13252 28022
rect 13206 27954 13252 27976
rect 13206 27904 13212 27954
rect 13246 27904 13252 27954
rect 13206 27886 13252 27904
rect 13206 27832 13212 27886
rect 13246 27832 13252 27886
rect 13206 27818 13252 27832
rect 13206 27760 13212 27818
rect 13246 27760 13252 27818
rect 13206 27750 13252 27760
rect 13206 27688 13212 27750
rect 13246 27688 13252 27750
rect 13206 27682 13252 27688
rect 13206 27616 13212 27682
rect 13246 27616 13252 27682
rect 13206 27614 13252 27616
rect 13206 27580 13212 27614
rect 13246 27580 13252 27614
rect 13206 27578 13252 27580
rect 13206 27512 13212 27578
rect 13246 27512 13252 27578
rect 13206 27506 13252 27512
rect 13206 27444 13212 27506
rect 13246 27444 13252 27506
rect 13206 27434 13252 27444
rect 13206 27376 13212 27434
rect 13246 27376 13252 27434
rect 13206 27362 13252 27376
rect 13206 27308 13212 27362
rect 13246 27308 13252 27362
rect 13206 27290 13252 27308
rect 13206 27240 13212 27290
rect 13246 27240 13252 27290
rect 13206 27218 13252 27240
rect 13206 27172 13212 27218
rect 13246 27172 13252 27218
rect 13206 27146 13252 27172
rect 13206 27104 13212 27146
rect 13246 27104 13252 27146
rect 13206 27074 13252 27104
rect 13206 27036 13212 27074
rect 13246 27036 13252 27074
rect 13206 27002 13252 27036
rect 13206 26968 13212 27002
rect 13246 26968 13252 27002
rect 13206 26934 13252 26968
rect 13206 26896 13212 26934
rect 13246 26896 13252 26934
rect 13206 26866 13252 26896
rect 13206 26824 13212 26866
rect 13246 26824 13252 26866
rect 13206 26798 13252 26824
rect 13206 26752 13212 26798
rect 13246 26752 13252 26798
rect 13206 26730 13252 26752
rect 13206 26680 13212 26730
rect 13246 26680 13252 26730
rect 13206 26662 13252 26680
rect 13206 26608 13212 26662
rect 13246 26608 13252 26662
rect 13206 26594 13252 26608
rect 13206 26536 13212 26594
rect 13246 26536 13252 26594
rect 13206 26526 13252 26536
rect 13206 26464 13212 26526
rect 13246 26464 13252 26526
rect 13206 26458 13252 26464
rect 13206 26392 13212 26458
rect 13246 26392 13252 26458
rect 13206 26390 13252 26392
rect 13206 26356 13212 26390
rect 13246 26356 13252 26390
rect 13206 26354 13252 26356
rect 13206 26288 13212 26354
rect 13246 26288 13252 26354
rect 13206 26282 13252 26288
rect 13206 26220 13212 26282
rect 13246 26220 13252 26282
rect 13206 26210 13252 26220
rect 13206 26152 13212 26210
rect 13246 26152 13252 26210
rect 13206 26138 13252 26152
rect 13206 26084 13212 26138
rect 13246 26084 13252 26138
rect 13206 26066 13252 26084
rect 13206 26016 13212 26066
rect 13246 26016 13252 26066
rect 13206 25994 13252 26016
rect 13206 25948 13212 25994
rect 13246 25948 13252 25994
rect 13206 25922 13252 25948
rect 13206 25880 13212 25922
rect 13246 25880 13252 25922
rect 13206 25850 13252 25880
rect 13206 25812 13212 25850
rect 13246 25812 13252 25850
rect 13206 25778 13252 25812
rect 13206 25744 13212 25778
rect 13246 25744 13252 25778
rect 13206 25710 13252 25744
rect 13206 25672 13212 25710
rect 13246 25672 13252 25710
rect 13206 25642 13252 25672
rect 13206 25600 13212 25642
rect 13246 25600 13252 25642
rect 13206 25574 13252 25600
rect 13206 25528 13212 25574
rect 13246 25528 13252 25574
rect 13206 25506 13252 25528
rect 13206 25456 13212 25506
rect 13246 25456 13252 25506
rect 13206 25438 13252 25456
rect 13206 25384 13212 25438
rect 13246 25384 13252 25438
rect 13206 25370 13252 25384
rect 13206 25312 13212 25370
rect 13246 25312 13252 25370
rect 13206 25302 13252 25312
rect 13206 25240 13212 25302
rect 13246 25240 13252 25302
rect 13206 25234 13252 25240
rect 13206 25168 13212 25234
rect 13246 25168 13252 25234
rect 13206 25166 13252 25168
rect 13206 25132 13212 25166
rect 13246 25132 13252 25166
rect 13206 25130 13252 25132
rect 13206 25064 13212 25130
rect 13246 25064 13252 25130
rect 13206 25058 13252 25064
rect 13206 24996 13212 25058
rect 13246 24996 13252 25058
rect 13206 24986 13252 24996
rect 13206 24928 13212 24986
rect 13246 24928 13252 24986
rect 13206 24914 13252 24928
rect 13206 24860 13212 24914
rect 13246 24860 13252 24914
rect 13206 24842 13252 24860
rect 13206 24792 13212 24842
rect 13246 24792 13252 24842
rect 13206 24770 13252 24792
rect 13206 24724 13212 24770
rect 13246 24724 13252 24770
rect 13206 24698 13252 24724
rect 13206 24656 13212 24698
rect 13246 24656 13252 24698
rect 13206 24626 13252 24656
rect 13206 24588 13212 24626
rect 13246 24588 13252 24626
rect 13206 24554 13252 24588
rect 13206 24520 13212 24554
rect 13246 24520 13252 24554
rect 13206 24486 13252 24520
rect 13206 24448 13212 24486
rect 13246 24448 13252 24486
rect 13206 24418 13252 24448
rect 13206 24376 13212 24418
rect 13246 24376 13252 24418
rect 13206 24350 13252 24376
rect 13206 24304 13212 24350
rect 13246 24304 13252 24350
rect 13206 24282 13252 24304
rect 13206 24232 13212 24282
rect 13246 24232 13252 24282
rect 13206 24214 13252 24232
rect 13206 24160 13212 24214
rect 13246 24160 13252 24214
rect 13206 24146 13252 24160
rect 13206 24088 13212 24146
rect 13246 24088 13252 24146
rect 13206 24078 13252 24088
rect 13206 24016 13212 24078
rect 13246 24016 13252 24078
rect 13206 24010 13252 24016
rect 13206 23944 13212 24010
rect 13246 23944 13252 24010
rect 13206 23942 13252 23944
rect 13206 23908 13212 23942
rect 13246 23908 13252 23942
rect 13206 23906 13252 23908
rect 13206 23840 13212 23906
rect 13246 23840 13252 23906
rect 13206 23834 13252 23840
rect 13206 23772 13212 23834
rect 13246 23772 13252 23834
rect 13206 23762 13252 23772
rect 13206 23704 13212 23762
rect 13246 23704 13252 23762
rect 13206 23690 13252 23704
rect 13206 23636 13212 23690
rect 13246 23636 13252 23690
rect 13206 23618 13252 23636
rect 13206 23568 13212 23618
rect 13246 23568 13252 23618
rect 13206 23546 13252 23568
rect 13206 23500 13212 23546
rect 13246 23500 13252 23546
rect 13206 23474 13252 23500
rect 13206 23432 13212 23474
rect 13246 23432 13252 23474
rect 13206 23402 13252 23432
rect 13206 23364 13212 23402
rect 13246 23364 13252 23402
rect 13206 23330 13252 23364
rect 13206 23296 13212 23330
rect 13246 23296 13252 23330
rect 13206 23262 13252 23296
rect 13206 23224 13212 23262
rect 13246 23224 13252 23262
rect 13206 23194 13252 23224
rect 13206 23152 13212 23194
rect 13246 23152 13252 23194
rect 13206 23126 13252 23152
rect 13206 23080 13212 23126
rect 13246 23080 13252 23126
rect 13206 23058 13252 23080
rect 13206 23008 13212 23058
rect 13246 23008 13252 23058
rect 13206 22990 13252 23008
rect 13206 22936 13212 22990
rect 13246 22936 13252 22990
rect 13206 22922 13252 22936
rect 13206 22864 13212 22922
rect 13246 22864 13252 22922
rect 13206 22854 13252 22864
rect 13206 22792 13212 22854
rect 13246 22792 13252 22854
rect 13206 22786 13252 22792
rect 13206 22720 13212 22786
rect 13246 22720 13252 22786
rect 13206 22718 13252 22720
rect 13206 22684 13212 22718
rect 13246 22684 13252 22718
rect 13206 22682 13252 22684
rect 13206 22616 13212 22682
rect 13246 22616 13252 22682
rect 13206 22610 13252 22616
rect 13206 22548 13212 22610
rect 13246 22548 13252 22610
rect 13206 22538 13252 22548
rect 13206 22480 13212 22538
rect 13246 22480 13252 22538
rect 13206 22466 13252 22480
rect 13206 22412 13212 22466
rect 13246 22412 13252 22466
rect 13206 22394 13252 22412
rect 13206 22344 13212 22394
rect 13246 22344 13252 22394
rect 13206 22322 13252 22344
rect 13206 22276 13212 22322
rect 13246 22276 13252 22322
rect 13206 22250 13252 22276
rect 13206 22208 13212 22250
rect 13246 22208 13252 22250
rect 13206 22178 13252 22208
rect 13206 22140 13212 22178
rect 13246 22140 13252 22178
rect 13206 22106 13252 22140
rect 13206 22072 13212 22106
rect 13246 22072 13252 22106
rect 13206 22038 13252 22072
rect 13206 22000 13212 22038
rect 13246 22000 13252 22038
rect 13206 21970 13252 22000
rect 13206 21928 13212 21970
rect 13246 21928 13252 21970
rect 13206 21902 13252 21928
rect 13206 21856 13212 21902
rect 13246 21856 13252 21902
rect 13206 21834 13252 21856
rect 13206 21784 13212 21834
rect 13246 21784 13252 21834
rect 13206 21766 13252 21784
rect 13206 21712 13212 21766
rect 13246 21712 13252 21766
rect 13206 21698 13252 21712
rect 13206 21640 13212 21698
rect 13246 21640 13252 21698
rect 13206 21630 13252 21640
rect 13206 21568 13212 21630
rect 13246 21568 13252 21630
rect 13206 21562 13252 21568
rect 13206 21496 13212 21562
rect 13246 21496 13252 21562
rect 13206 21494 13252 21496
rect 13206 21460 13212 21494
rect 13246 21460 13252 21494
rect 13206 21458 13252 21460
rect 13206 21392 13212 21458
rect 13246 21392 13252 21458
rect 13206 21386 13252 21392
rect 13206 21324 13212 21386
rect 13246 21324 13252 21386
rect 13206 21314 13252 21324
rect 13206 21256 13212 21314
rect 13246 21256 13252 21314
rect 13206 21242 13252 21256
rect 13206 21188 13212 21242
rect 13246 21188 13252 21242
rect 13206 21170 13252 21188
rect 13206 21120 13212 21170
rect 13246 21120 13252 21170
rect 13206 21098 13252 21120
rect 13206 21052 13212 21098
rect 13246 21052 13252 21098
rect 13206 21026 13252 21052
rect 13206 20984 13212 21026
rect 13246 20984 13252 21026
rect 13206 20954 13252 20984
rect 13206 20916 13212 20954
rect 13246 20916 13252 20954
rect 13206 20882 13252 20916
rect 13206 20848 13212 20882
rect 13246 20848 13252 20882
rect 13206 20814 13252 20848
rect 13206 20776 13212 20814
rect 13246 20776 13252 20814
rect 13206 20746 13252 20776
rect 13206 20704 13212 20746
rect 13246 20704 13252 20746
rect 13206 20678 13252 20704
rect 13206 20632 13212 20678
rect 13246 20632 13252 20678
rect 13206 20610 13252 20632
rect 13206 20560 13212 20610
rect 13246 20560 13252 20610
rect 13206 20542 13252 20560
rect 13206 20488 13212 20542
rect 13246 20488 13252 20542
rect 13206 20474 13252 20488
rect 13206 20416 13212 20474
rect 13246 20416 13252 20474
rect 13206 20406 13252 20416
rect 13206 20344 13212 20406
rect 13246 20344 13252 20406
rect 13206 20338 13252 20344
rect 13206 20272 13212 20338
rect 13246 20272 13252 20338
rect 13206 20270 13252 20272
rect 13206 20236 13212 20270
rect 13246 20236 13252 20270
rect 13206 20234 13252 20236
rect 13206 20168 13212 20234
rect 13246 20168 13252 20234
rect 13206 20162 13252 20168
rect 13206 20100 13212 20162
rect 13246 20100 13252 20162
rect 13206 20090 13252 20100
rect 13206 20032 13212 20090
rect 13246 20032 13252 20090
rect 13206 20018 13252 20032
rect 13206 19964 13212 20018
rect 13246 19964 13252 20018
rect 13206 19946 13252 19964
rect 13206 19896 13212 19946
rect 13246 19896 13252 19946
rect 13206 19874 13252 19896
rect 13206 19828 13212 19874
rect 13246 19828 13252 19874
rect 13206 19802 13252 19828
rect 13206 19760 13212 19802
rect 13246 19760 13252 19802
rect 13206 19730 13252 19760
rect 13206 19692 13212 19730
rect 13246 19692 13252 19730
rect 13206 19658 13252 19692
rect 13206 19624 13212 19658
rect 13246 19624 13252 19658
rect 13206 19590 13252 19624
rect 13206 19552 13212 19590
rect 13246 19552 13252 19590
rect 13206 19522 13252 19552
rect 13206 19480 13212 19522
rect 13246 19480 13252 19522
rect 13206 19454 13252 19480
rect 13206 19408 13212 19454
rect 13246 19408 13252 19454
rect 13206 19386 13252 19408
rect 13206 19336 13212 19386
rect 13246 19336 13252 19386
rect 13206 19318 13252 19336
rect 13206 19264 13212 19318
rect 13246 19264 13252 19318
rect 13206 19250 13252 19264
rect 13206 19192 13212 19250
rect 13246 19192 13252 19250
rect 13206 19182 13252 19192
rect 13206 19120 13212 19182
rect 13246 19120 13252 19182
rect 13206 19114 13252 19120
rect 13206 19048 13212 19114
rect 13246 19048 13252 19114
rect 13206 19046 13252 19048
rect 13206 19012 13212 19046
rect 13246 19012 13252 19046
rect 13206 19010 13252 19012
rect 13206 18944 13212 19010
rect 13246 18944 13252 19010
rect 13206 18938 13252 18944
rect 13206 18876 13212 18938
rect 13246 18876 13252 18938
rect 13206 18866 13252 18876
rect 13206 18808 13212 18866
rect 13246 18808 13252 18866
rect 13206 18794 13252 18808
rect 13206 18740 13212 18794
rect 13246 18740 13252 18794
rect 13206 18722 13252 18740
rect 13206 18672 13212 18722
rect 13246 18672 13252 18722
rect 13206 18650 13252 18672
rect 13206 18604 13212 18650
rect 13246 18604 13252 18650
rect 13206 18578 13252 18604
rect 13206 18536 13212 18578
rect 13246 18536 13252 18578
rect 13206 18506 13252 18536
rect 13206 18468 13212 18506
rect 13246 18468 13252 18506
rect 13206 18434 13252 18468
rect 13206 18400 13212 18434
rect 13246 18400 13252 18434
rect 13206 18366 13252 18400
rect 13206 18328 13212 18366
rect 13246 18328 13252 18366
rect 13206 18298 13252 18328
rect 13206 18256 13212 18298
rect 13246 18256 13252 18298
rect 13206 18230 13252 18256
rect 13206 18184 13212 18230
rect 13246 18184 13252 18230
rect 13206 18162 13252 18184
rect 13206 18112 13212 18162
rect 13246 18112 13252 18162
rect 13206 18094 13252 18112
rect 13206 18040 13212 18094
rect 13246 18040 13252 18094
rect 13206 18026 13252 18040
rect 13206 17968 13212 18026
rect 13246 17968 13252 18026
rect 13206 17958 13252 17968
rect 13206 17896 13212 17958
rect 13246 17896 13252 17958
rect 13206 17890 13252 17896
rect 13206 17824 13212 17890
rect 13246 17824 13252 17890
rect 13206 17822 13252 17824
rect 13206 17788 13212 17822
rect 13246 17788 13252 17822
rect 13206 17786 13252 17788
rect 13206 17720 13212 17786
rect 13246 17720 13252 17786
rect 13206 17714 13252 17720
rect 13206 17652 13212 17714
rect 13246 17652 13252 17714
rect 13206 17642 13252 17652
rect 13206 17584 13212 17642
rect 13246 17584 13252 17642
rect 13206 17570 13252 17584
rect 13206 17516 13212 17570
rect 13246 17516 13252 17570
rect 13206 17498 13252 17516
rect 13206 17448 13212 17498
rect 13246 17448 13252 17498
rect 13206 17426 13252 17448
rect 13206 17380 13212 17426
rect 13246 17380 13252 17426
rect 13206 17354 13252 17380
rect 13206 17312 13212 17354
rect 13246 17312 13252 17354
rect 13206 17282 13252 17312
rect 13206 17244 13212 17282
rect 13246 17244 13252 17282
rect 13206 17210 13252 17244
rect 13206 17176 13212 17210
rect 13246 17176 13252 17210
rect 13206 17142 13252 17176
rect 13206 17104 13212 17142
rect 13246 17104 13252 17142
rect 13206 17074 13252 17104
rect 13206 17032 13212 17074
rect 13246 17032 13252 17074
rect 13206 17006 13252 17032
rect 13206 16960 13212 17006
rect 13246 16960 13252 17006
rect 13206 16938 13252 16960
rect 13206 16888 13212 16938
rect 13246 16888 13252 16938
rect 13206 16870 13252 16888
rect 13206 16816 13212 16870
rect 13246 16816 13252 16870
rect 13206 16802 13252 16816
rect 13206 16744 13212 16802
rect 13246 16744 13252 16802
rect 13206 16734 13252 16744
rect 13206 16672 13212 16734
rect 13246 16672 13252 16734
rect 13206 16666 13252 16672
rect 13206 16600 13212 16666
rect 13246 16600 13252 16666
rect 13206 16598 13252 16600
rect 13206 16564 13212 16598
rect 13246 16564 13252 16598
rect 13206 16562 13252 16564
rect 13206 16496 13212 16562
rect 13246 16496 13252 16562
rect 13206 16490 13252 16496
rect 13206 16428 13212 16490
rect 13246 16428 13252 16490
rect 13206 16418 13252 16428
rect 13206 16360 13212 16418
rect 13246 16360 13252 16418
rect 13206 16346 13252 16360
rect 13206 16292 13212 16346
rect 13246 16292 13252 16346
rect 13206 16274 13252 16292
rect 13206 16224 13212 16274
rect 13246 16224 13252 16274
rect 13206 16202 13252 16224
rect 13206 16156 13212 16202
rect 13246 16156 13252 16202
rect 13206 16130 13252 16156
rect 13206 16088 13212 16130
rect 13246 16088 13252 16130
rect 13206 16058 13252 16088
rect 13206 16020 13212 16058
rect 13246 16020 13252 16058
rect 13206 15986 13252 16020
rect 13206 15952 13212 15986
rect 13246 15952 13252 15986
rect 13206 15918 13252 15952
rect 13206 15880 13212 15918
rect 13246 15880 13252 15918
rect 13206 15850 13252 15880
rect 13206 15808 13212 15850
rect 13246 15808 13252 15850
rect 13206 15782 13252 15808
rect 13206 15736 13212 15782
rect 13246 15736 13252 15782
rect 13206 15714 13252 15736
rect 13206 15664 13212 15714
rect 13246 15664 13252 15714
rect 13206 15646 13252 15664
rect 13206 15592 13212 15646
rect 13246 15592 13252 15646
rect 13206 15578 13252 15592
rect 13206 15520 13212 15578
rect 13246 15520 13252 15578
rect 13206 15510 13252 15520
rect 13206 15448 13212 15510
rect 13246 15448 13252 15510
rect 13206 15442 13252 15448
rect 13206 15376 13212 15442
rect 13246 15376 13252 15442
rect 13206 15374 13252 15376
rect 13206 15340 13212 15374
rect 13246 15340 13252 15374
rect 13206 15338 13252 15340
rect 13206 15272 13212 15338
rect 13246 15272 13252 15338
rect 13206 15266 13252 15272
rect 13206 15204 13212 15266
rect 13246 15204 13252 15266
rect 13206 15194 13252 15204
rect 13206 15136 13212 15194
rect 13246 15136 13252 15194
rect 13206 15122 13252 15136
rect 13206 15068 13212 15122
rect 13246 15068 13252 15122
rect 13206 15050 13252 15068
rect 13206 15000 13212 15050
rect 13246 15000 13252 15050
rect 13206 14978 13252 15000
rect 13206 14932 13212 14978
rect 13246 14932 13252 14978
rect 13206 14906 13252 14932
rect 13206 14864 13212 14906
rect 13246 14864 13252 14906
rect 13206 14834 13252 14864
rect 13206 14796 13212 14834
rect 13246 14796 13252 14834
rect 13206 14762 13252 14796
rect 13206 14728 13212 14762
rect 13246 14728 13252 14762
rect 13206 14694 13252 14728
rect 13206 14656 13212 14694
rect 13246 14656 13252 14694
rect 13206 14626 13252 14656
rect 13206 14584 13212 14626
rect 13246 14584 13252 14626
rect 13206 14558 13252 14584
rect 13206 14512 13212 14558
rect 13246 14512 13252 14558
rect 13206 14490 13252 14512
rect 13206 14440 13212 14490
rect 13246 14440 13252 14490
rect 13206 14422 13252 14440
rect 13206 14368 13212 14422
rect 13246 14368 13252 14422
rect 13206 14354 13252 14368
rect 13206 14296 13212 14354
rect 13246 14296 13252 14354
rect 13206 14286 13252 14296
rect 13206 14224 13212 14286
rect 13246 14224 13252 14286
rect 13206 14218 13252 14224
rect 13206 14152 13212 14218
rect 13246 14152 13252 14218
rect 13206 14150 13252 14152
rect 13206 14116 13212 14150
rect 13246 14116 13252 14150
rect 13206 14114 13252 14116
rect 13206 14048 13212 14114
rect 13246 14048 13252 14114
rect 13206 14042 13252 14048
rect 13206 13980 13212 14042
rect 13246 13980 13252 14042
rect 13206 13970 13252 13980
rect 13206 13912 13212 13970
rect 13246 13912 13252 13970
rect 13206 13898 13252 13912
rect 13206 13844 13212 13898
rect 13246 13844 13252 13898
rect 13206 13826 13252 13844
rect 13206 13776 13212 13826
rect 13246 13776 13252 13826
rect 13206 13754 13252 13776
rect 13206 13708 13212 13754
rect 13246 13708 13252 13754
rect 13206 13682 13252 13708
rect 13206 13640 13212 13682
rect 13246 13640 13252 13682
rect 13206 13610 13252 13640
rect 13206 13572 13212 13610
rect 13246 13572 13252 13610
rect 13206 13538 13252 13572
rect 13206 13504 13212 13538
rect 13246 13504 13252 13538
rect 13206 13470 13252 13504
rect 13206 13432 13212 13470
rect 13246 13432 13252 13470
rect 13206 13402 13252 13432
rect 13206 13360 13212 13402
rect 13246 13360 13252 13402
rect 13206 13334 13252 13360
rect 13206 13288 13212 13334
rect 13246 13288 13252 13334
rect 13206 13266 13252 13288
rect 13206 13216 13212 13266
rect 13246 13216 13252 13266
rect 13206 13198 13252 13216
rect 13206 13144 13212 13198
rect 13246 13144 13252 13198
rect 13206 13130 13252 13144
rect 13206 13072 13212 13130
rect 13246 13072 13252 13130
rect 13206 13062 13252 13072
rect 13206 13000 13212 13062
rect 13246 13000 13252 13062
rect 13206 12994 13252 13000
rect 13206 12928 13212 12994
rect 13246 12928 13252 12994
rect 13206 12926 13252 12928
rect 13206 12892 13212 12926
rect 13246 12892 13252 12926
rect 13206 12890 13252 12892
rect 13206 12824 13212 12890
rect 13246 12824 13252 12890
rect 13206 12818 13252 12824
rect 13206 12756 13212 12818
rect 13246 12756 13252 12818
rect 13206 12746 13252 12756
rect 13206 12688 13212 12746
rect 13246 12688 13252 12746
rect 13206 12674 13252 12688
rect 13206 12620 13212 12674
rect 13246 12620 13252 12674
rect 13206 12602 13252 12620
rect 13206 12552 13212 12602
rect 13246 12552 13252 12602
rect 13206 12530 13252 12552
rect 13206 12484 13212 12530
rect 13246 12484 13252 12530
rect 13206 12458 13252 12484
rect 13206 12416 13212 12458
rect 13246 12416 13252 12458
rect 13206 12386 13252 12416
rect 13206 12348 13212 12386
rect 13246 12348 13252 12386
rect 13206 12314 13252 12348
rect 13206 12280 13212 12314
rect 13246 12280 13252 12314
rect 13206 12246 13252 12280
rect 13206 12208 13212 12246
rect 13246 12208 13252 12246
rect 13206 12178 13252 12208
rect 13206 12136 13212 12178
rect 13246 12136 13252 12178
rect 13206 12110 13252 12136
rect 13206 12064 13212 12110
rect 13246 12064 13252 12110
rect 13206 12042 13252 12064
rect 13206 11992 13212 12042
rect 13246 11992 13252 12042
rect 13206 11974 13252 11992
rect 13206 11920 13212 11974
rect 13246 11920 13252 11974
rect 13206 11906 13252 11920
rect 13206 11848 13212 11906
rect 13246 11848 13252 11906
rect 13206 11838 13252 11848
rect 13206 11776 13212 11838
rect 13246 11776 13252 11838
rect 13206 11770 13252 11776
rect 13206 11704 13212 11770
rect 13246 11704 13252 11770
rect 13206 11702 13252 11704
rect 13206 11668 13212 11702
rect 13246 11668 13252 11702
rect 13206 11666 13252 11668
rect 13206 11600 13212 11666
rect 13246 11600 13252 11666
rect 13206 11594 13252 11600
rect 13206 11532 13212 11594
rect 13246 11532 13252 11594
rect 13206 11522 13252 11532
rect 13206 11464 13212 11522
rect 13246 11464 13252 11522
rect 13206 11450 13252 11464
rect 13206 11396 13212 11450
rect 13246 11396 13252 11450
rect 13206 11378 13252 11396
rect 13206 11328 13212 11378
rect 13246 11328 13252 11378
rect 13206 11306 13252 11328
rect 13206 11260 13212 11306
rect 13246 11260 13252 11306
rect 13206 11234 13252 11260
rect 13206 11192 13212 11234
rect 13246 11192 13252 11234
rect 13206 11162 13252 11192
rect 13206 11124 13212 11162
rect 13246 11124 13252 11162
rect 13206 11090 13252 11124
rect 13206 11056 13212 11090
rect 13246 11056 13252 11090
rect 13206 11022 13252 11056
rect 13206 10984 13212 11022
rect 13246 10984 13252 11022
rect 13206 10954 13252 10984
rect 13206 10912 13212 10954
rect 13246 10912 13252 10954
rect 13206 10886 13252 10912
rect 13206 10840 13212 10886
rect 13246 10840 13252 10886
rect 13206 10818 13252 10840
rect 13206 10768 13212 10818
rect 13246 10768 13252 10818
rect 13206 10750 13252 10768
rect 13206 10696 13212 10750
rect 13246 10696 13252 10750
rect 13206 10682 13252 10696
rect 13206 10624 13212 10682
rect 13246 10624 13252 10682
rect 13206 10614 13252 10624
rect 13206 10552 13212 10614
rect 13246 10552 13252 10614
rect 13206 10546 13252 10552
rect 13206 10480 13212 10546
rect 13246 10480 13252 10546
rect 13206 10478 13252 10480
rect 13206 10444 13212 10478
rect 13246 10444 13252 10478
rect 13206 10442 13252 10444
rect 13206 10376 13212 10442
rect 13246 10376 13252 10442
rect 13206 10370 13252 10376
rect 13206 10308 13212 10370
rect 13246 10308 13252 10370
rect 13206 10298 13252 10308
rect 13206 10240 13212 10298
rect 13246 10240 13252 10298
rect 13206 10226 13252 10240
rect 13206 10172 13212 10226
rect 13246 10172 13252 10226
rect 13206 10154 13252 10172
rect 13206 10104 13212 10154
rect 13246 10104 13252 10154
rect 13206 10082 13252 10104
rect 13206 10036 13212 10082
rect 13246 10036 13252 10082
rect 13206 10010 13252 10036
rect 13206 9968 13212 10010
rect 13246 9968 13252 10010
rect 13206 9938 13252 9968
rect 13206 9900 13212 9938
rect 13246 9900 13252 9938
rect 13206 9866 13252 9900
rect 13206 9832 13212 9866
rect 13246 9832 13252 9866
rect 13206 9798 13252 9832
rect 13206 9760 13212 9798
rect 13246 9760 13252 9798
rect 13206 9730 13252 9760
rect 13206 9688 13212 9730
rect 13246 9688 13252 9730
rect 13206 9662 13252 9688
rect 13206 9616 13212 9662
rect 13246 9616 13252 9662
rect 13206 9594 13252 9616
rect 13206 9544 13212 9594
rect 13246 9544 13252 9594
rect 13206 9526 13252 9544
rect 13206 9472 13212 9526
rect 13246 9472 13252 9526
rect 13206 9458 13252 9472
rect 13206 9400 13212 9458
rect 13246 9400 13252 9458
rect 13206 9390 13252 9400
rect 13206 9328 13212 9390
rect 13246 9328 13252 9390
rect 13206 9322 13252 9328
rect 13206 9256 13212 9322
rect 13246 9256 13252 9322
rect 13206 9254 13252 9256
rect 13206 9220 13212 9254
rect 13246 9220 13252 9254
rect 13206 9218 13252 9220
rect 13206 9152 13212 9218
rect 13246 9152 13252 9218
rect 13206 9146 13252 9152
rect 13206 9084 13212 9146
rect 13246 9084 13252 9146
rect 13206 9074 13252 9084
rect 13206 9016 13212 9074
rect 13246 9016 13252 9074
rect 13206 9002 13252 9016
rect 13206 8948 13212 9002
rect 13246 8948 13252 9002
rect 13206 8930 13252 8948
rect 13206 8880 13212 8930
rect 13246 8880 13252 8930
rect 13206 8858 13252 8880
rect 13206 8812 13212 8858
rect 13246 8812 13252 8858
rect 13206 8786 13252 8812
rect 13206 8744 13212 8786
rect 13246 8744 13252 8786
rect 13206 8714 13252 8744
rect 13206 8676 13212 8714
rect 13246 8676 13252 8714
rect 13206 8642 13252 8676
rect 13206 8608 13212 8642
rect 13246 8608 13252 8642
rect 13206 8574 13252 8608
rect 13206 8536 13212 8574
rect 13246 8536 13252 8574
rect 13206 8506 13252 8536
rect 13206 8464 13212 8506
rect 13246 8464 13252 8506
rect 13206 8438 13252 8464
rect 13206 8392 13212 8438
rect 13246 8392 13252 8438
rect 13206 8370 13252 8392
rect 13206 8320 13212 8370
rect 13246 8320 13252 8370
rect 13206 8302 13252 8320
rect 13206 8248 13212 8302
rect 13246 8248 13252 8302
rect 13206 8234 13252 8248
rect 13206 8176 13212 8234
rect 13246 8176 13252 8234
rect 13206 8166 13252 8176
rect 13206 8104 13212 8166
rect 13246 8104 13252 8166
rect 13206 8098 13252 8104
rect 13206 8032 13212 8098
rect 13246 8032 13252 8098
rect 13206 8030 13252 8032
rect 13206 7996 13212 8030
rect 13246 7996 13252 8030
rect 13206 7994 13252 7996
rect 13206 7928 13212 7994
rect 13246 7928 13252 7994
rect 13206 7922 13252 7928
rect 13206 7860 13212 7922
rect 13246 7860 13252 7922
rect 13206 7850 13252 7860
rect 13206 7792 13212 7850
rect 13246 7792 13252 7850
rect 13206 7778 13252 7792
rect 13206 7724 13212 7778
rect 13246 7724 13252 7778
rect 13206 7706 13252 7724
rect 13206 7656 13212 7706
rect 13246 7656 13252 7706
rect 13206 7634 13252 7656
rect 13206 7588 13212 7634
rect 13246 7588 13252 7634
rect 13206 7562 13252 7588
rect 13206 7520 13212 7562
rect 13246 7520 13252 7562
rect 13206 7490 13252 7520
rect 13206 7452 13212 7490
rect 13246 7452 13252 7490
rect 13206 7418 13252 7452
rect 13206 7384 13212 7418
rect 13246 7384 13252 7418
rect 13206 7350 13252 7384
rect 13206 7312 13212 7350
rect 13246 7312 13252 7350
rect 13206 7282 13252 7312
rect 13206 7240 13212 7282
rect 13246 7240 13252 7282
rect 13206 7214 13252 7240
rect 13206 7168 13212 7214
rect 13246 7168 13252 7214
rect 13206 7146 13252 7168
rect 13206 7096 13212 7146
rect 13246 7096 13252 7146
rect 13206 7078 13252 7096
rect 13206 7024 13212 7078
rect 13246 7024 13252 7078
rect 13206 7010 13252 7024
rect 13206 6952 13212 7010
rect 13246 6952 13252 7010
rect 13206 6942 13252 6952
rect 13206 6880 13212 6942
rect 13246 6880 13252 6942
rect 13206 6874 13252 6880
rect 13206 6808 13212 6874
rect 13246 6808 13252 6874
rect 13206 6806 13252 6808
rect 13206 6772 13212 6806
rect 13246 6772 13252 6806
rect 13206 6770 13252 6772
rect 13206 6704 13212 6770
rect 13246 6704 13252 6770
rect 13206 6698 13252 6704
rect 13206 6636 13212 6698
rect 13246 6636 13252 6698
rect 13206 6626 13252 6636
rect 13206 6568 13212 6626
rect 13246 6568 13252 6626
rect 13206 6554 13252 6568
rect 13206 6500 13212 6554
rect 13246 6500 13252 6554
rect 13206 6482 13252 6500
rect 13206 6432 13212 6482
rect 13246 6432 13252 6482
rect 13206 6410 13252 6432
rect 13206 6364 13212 6410
rect 13246 6364 13252 6410
rect 13206 6338 13252 6364
rect 13206 6296 13212 6338
rect 13246 6296 13252 6338
rect 13206 6266 13252 6296
rect 13206 6228 13212 6266
rect 13246 6228 13252 6266
rect 13206 6194 13252 6228
rect 13206 6160 13212 6194
rect 13246 6160 13252 6194
rect 13206 6126 13252 6160
rect 13206 6088 13212 6126
rect 13246 6088 13252 6126
rect 13206 6058 13252 6088
rect 13206 6016 13212 6058
rect 13246 6016 13252 6058
rect 13206 5990 13252 6016
rect 13206 5944 13212 5990
rect 13246 5944 13252 5990
rect 13206 5922 13252 5944
rect 13206 5872 13212 5922
rect 13246 5872 13252 5922
rect 13206 5854 13252 5872
rect 13206 5800 13212 5854
rect 13246 5800 13252 5854
rect 13206 5786 13252 5800
rect 13206 5728 13212 5786
rect 13246 5728 13252 5786
rect 13206 5718 13252 5728
rect 13206 5656 13212 5718
rect 13246 5656 13252 5718
rect 13206 5650 13252 5656
rect 13206 5584 13212 5650
rect 13246 5584 13252 5650
rect 13206 5582 13252 5584
rect 13206 5548 13212 5582
rect 13246 5548 13252 5582
rect 13206 5546 13252 5548
rect 13206 5480 13212 5546
rect 13246 5480 13252 5546
rect 13206 5474 13252 5480
rect 13206 5412 13212 5474
rect 13246 5412 13252 5474
rect 13206 5402 13252 5412
rect 13206 5344 13212 5402
rect 13246 5344 13252 5402
rect 13206 5330 13252 5344
rect 13206 5276 13212 5330
rect 13246 5276 13252 5330
rect 13206 5258 13252 5276
rect 13206 5208 13212 5258
rect 13246 5208 13252 5258
rect 13206 5186 13252 5208
rect 13206 5140 13212 5186
rect 13246 5140 13252 5186
rect 13206 5114 13252 5140
rect 13206 5072 13212 5114
rect 13246 5072 13252 5114
rect 13206 5042 13252 5072
rect 13206 5004 13212 5042
rect 13246 5004 13252 5042
rect 13206 4970 13252 5004
rect 13206 4936 13212 4970
rect 13246 4936 13252 4970
rect 13206 4902 13252 4936
rect 13206 4864 13212 4902
rect 13246 4864 13252 4902
rect 13206 4834 13252 4864
rect 13206 4792 13212 4834
rect 13246 4792 13252 4834
rect 13206 4766 13252 4792
rect 13206 4720 13212 4766
rect 13246 4720 13252 4766
rect 13206 4698 13252 4720
rect 13206 4648 13212 4698
rect 13246 4648 13252 4698
rect 13206 4630 13252 4648
rect 13206 4576 13212 4630
rect 13246 4576 13252 4630
rect 13206 4562 13252 4576
rect 13206 4504 13212 4562
rect 13246 4504 13252 4562
rect 13206 4494 13252 4504
rect 13206 4432 13212 4494
rect 13246 4432 13252 4494
rect 13206 4426 13252 4432
rect 13206 4360 13212 4426
rect 13246 4360 13252 4426
rect 13206 4358 13252 4360
rect 13206 4324 13212 4358
rect 13246 4324 13252 4358
rect 13206 4322 13252 4324
rect 13206 4256 13212 4322
rect 13246 4256 13252 4322
rect 13206 4250 13252 4256
rect 13206 4188 13212 4250
rect 13246 4188 13252 4250
rect 13206 4178 13252 4188
rect 13206 4120 13212 4178
rect 13246 4120 13252 4178
rect 13206 4106 13252 4120
rect 13206 4052 13212 4106
rect 13246 4052 13252 4106
rect 13206 4034 13252 4052
rect 13206 3984 13212 4034
rect 13246 3984 13252 4034
rect 13206 3962 13252 3984
rect 13206 3916 13212 3962
rect 13246 3916 13252 3962
rect 13206 3890 13252 3916
rect 13206 3848 13212 3890
rect 13246 3848 13252 3890
rect 13206 3818 13252 3848
rect 13206 3780 13212 3818
rect 13246 3780 13252 3818
rect 13206 3746 13252 3780
rect 13206 3712 13212 3746
rect 13246 3712 13252 3746
rect 13206 3678 13252 3712
rect 13206 3640 13212 3678
rect 13246 3640 13252 3678
rect 13206 3610 13252 3640
rect 13206 3568 13212 3610
rect 13246 3568 13252 3610
rect 13206 3542 13252 3568
rect 13206 3496 13212 3542
rect 13246 3496 13252 3542
rect 13206 3474 13252 3496
rect 13206 3424 13212 3474
rect 13246 3424 13252 3474
rect 13206 3406 13252 3424
rect 13206 3352 13212 3406
rect 13246 3352 13252 3406
rect 13206 3338 13252 3352
rect 13206 3280 13212 3338
rect 13246 3280 13252 3338
rect 13206 3270 13252 3280
rect 13206 3208 13212 3270
rect 13246 3208 13252 3270
rect 13206 3202 13252 3208
rect 13206 3136 13212 3202
rect 13246 3136 13252 3202
rect 13206 3134 13252 3136
rect 13206 3100 13212 3134
rect 13246 3100 13252 3134
rect 13206 3098 13252 3100
rect 13206 3032 13212 3098
rect 13246 3032 13252 3098
rect 13206 3026 13252 3032
rect 13206 2964 13212 3026
rect 13246 2964 13252 3026
rect 13206 2954 13252 2964
rect 13206 2896 13212 2954
rect 13246 2896 13252 2954
rect 13206 2882 13252 2896
rect 13206 2828 13212 2882
rect 13246 2828 13252 2882
rect 13206 2810 13252 2828
rect 13206 2760 13212 2810
rect 13246 2760 13252 2810
rect 13206 2738 13252 2760
rect 13206 2692 13212 2738
rect 13246 2692 13252 2738
rect 13206 2666 13252 2692
rect 13206 2624 13212 2666
rect 13246 2624 13252 2666
rect 13206 2594 13252 2624
rect 13206 2556 13212 2594
rect 13246 2556 13252 2594
rect 13206 2522 13252 2556
rect 13206 2488 13212 2522
rect 13246 2488 13252 2522
rect 13206 2454 13252 2488
rect 13206 2416 13212 2454
rect 13246 2416 13252 2454
rect 13206 2386 13252 2416
rect 13206 2344 13212 2386
rect 13246 2344 13252 2386
rect 13206 2318 13252 2344
rect 13206 2272 13212 2318
rect 13246 2272 13252 2318
rect 13206 2250 13252 2272
rect 13206 2200 13212 2250
rect 13246 2200 13252 2250
rect 13206 2182 13252 2200
rect 13206 2128 13212 2182
rect 13246 2128 13252 2182
rect 13206 2114 13252 2128
rect 13206 2056 13212 2114
rect 13246 2056 13252 2114
rect 13206 2046 13252 2056
rect 13206 1984 13212 2046
rect 13246 1984 13252 2046
rect 13206 1978 13252 1984
rect 13206 1912 13212 1978
rect 13246 1912 13252 1978
rect 13206 1910 13252 1912
rect 13206 1876 13212 1910
rect 13246 1876 13252 1910
rect 13206 1874 13252 1876
rect 13206 1808 13212 1874
rect 13246 1808 13252 1874
rect 13206 1802 13252 1808
rect 13206 1740 13212 1802
rect 13246 1740 13252 1802
rect 13206 1730 13252 1740
rect 13206 1672 13212 1730
rect 13246 1672 13252 1730
rect 13206 1658 13252 1672
rect 13206 1604 13212 1658
rect 13246 1604 13252 1658
rect 13206 1586 13252 1604
rect 13206 1536 13212 1586
rect 13246 1536 13252 1586
rect 13206 1514 13252 1536
rect 13206 1468 13212 1514
rect 13246 1468 13252 1514
rect 13206 1442 13252 1468
rect 13206 1400 13212 1442
rect 13246 1400 13252 1442
rect 13206 1370 13252 1400
rect 13206 1332 13212 1370
rect 13246 1332 13252 1370
rect 13206 1298 13252 1332
rect 13206 1264 13212 1298
rect 13246 1264 13252 1298
rect 13206 1230 13252 1264
rect 13206 1192 13212 1230
rect 13246 1192 13252 1230
rect 13206 1162 13252 1192
rect 13206 1120 13212 1162
rect 13246 1120 13252 1162
rect 13206 1094 13252 1120
rect 13206 1048 13212 1094
rect 13246 1048 13252 1094
rect 13206 1026 13252 1048
rect 13206 976 13212 1026
rect 13246 976 13252 1026
rect 13206 958 13252 976
rect 13206 904 13212 958
rect 13246 904 13252 958
rect 13206 890 13252 904
rect 13206 832 13212 890
rect 13246 832 13252 890
rect 13206 822 13252 832
rect 13206 760 13212 822
rect 13246 760 13252 822
rect 13206 754 13252 760
rect 13206 688 13212 754
rect 13246 688 13252 754
rect 13206 686 13252 688
rect 13206 652 13212 686
rect 13246 652 13252 686
rect 13206 650 13252 652
rect 13206 584 13212 650
rect 13246 584 13252 650
rect 13206 578 13252 584
rect 13206 516 13212 578
rect 13246 516 13252 578
rect 13206 506 13252 516
rect 13206 448 13212 506
rect 13246 448 13252 506
rect 13206 434 13252 448
rect 11418 366 11464 383
rect 11418 315 11424 366
rect 11458 315 11464 366
rect 11418 293 11464 315
rect 11418 247 11424 293
rect 11458 247 11464 293
rect 11594 383 11610 403
rect 11644 383 11660 403
rect 11594 345 11660 383
rect 11594 291 11610 345
rect 11644 325 11660 345
rect 13206 380 13212 434
rect 13246 380 13252 434
rect 14934 38434 14940 38485
rect 14974 38434 14980 38485
rect 14934 38417 14980 38434
rect 14934 38362 14940 38417
rect 14974 38362 14980 38417
rect 14934 38349 14980 38362
rect 14934 38290 14940 38349
rect 14974 38290 14980 38349
rect 14934 38281 14980 38290
rect 14934 38218 14940 38281
rect 14974 38218 14980 38281
rect 14934 38213 14980 38218
rect 14934 38146 14940 38213
rect 14974 38146 14980 38213
rect 14934 38145 14980 38146
rect 14934 38111 14940 38145
rect 14974 38111 14980 38145
rect 14934 38108 14980 38111
rect 14934 38043 14940 38108
rect 14974 38043 14980 38108
rect 14934 38036 14980 38043
rect 14934 37975 14940 38036
rect 14974 37975 14980 38036
rect 14934 37964 14980 37975
rect 14934 37907 14940 37964
rect 14974 37907 14980 37964
rect 14934 37892 14980 37907
rect 14934 37839 14940 37892
rect 14974 37839 14980 37892
rect 14934 37820 14980 37839
rect 14934 37771 14940 37820
rect 14974 37771 14980 37820
rect 14934 37748 14980 37771
rect 14934 37703 14940 37748
rect 14974 37703 14980 37748
rect 14934 37676 14980 37703
rect 14934 37635 14940 37676
rect 14974 37635 14980 37676
rect 14934 37604 14980 37635
rect 14934 37567 14940 37604
rect 14974 37567 14980 37604
rect 14934 37533 14980 37567
rect 14934 37498 14940 37533
rect 14974 37498 14980 37533
rect 14934 37465 14980 37498
rect 14934 37426 14940 37465
rect 14974 37426 14980 37465
rect 14934 37397 14980 37426
rect 14934 37354 14940 37397
rect 14974 37354 14980 37397
rect 14934 37329 14980 37354
rect 14934 37282 14940 37329
rect 14974 37282 14980 37329
rect 14934 37261 14980 37282
rect 14934 37210 14940 37261
rect 14974 37210 14980 37261
rect 14934 37193 14980 37210
rect 14934 37138 14940 37193
rect 14974 37138 14980 37193
rect 14934 37125 14980 37138
rect 14934 37066 14940 37125
rect 14974 37066 14980 37125
rect 14934 37057 14980 37066
rect 14934 36994 14940 37057
rect 14974 36994 14980 37057
rect 14934 36989 14980 36994
rect 14934 36922 14940 36989
rect 14974 36922 14980 36989
rect 14934 36921 14980 36922
rect 14934 36887 14940 36921
rect 14974 36887 14980 36921
rect 14934 36884 14980 36887
rect 14934 36819 14940 36884
rect 14974 36819 14980 36884
rect 14934 36812 14980 36819
rect 14934 36751 14940 36812
rect 14974 36751 14980 36812
rect 14934 36740 14980 36751
rect 14934 36683 14940 36740
rect 14974 36683 14980 36740
rect 14934 36668 14980 36683
rect 14934 36615 14940 36668
rect 14974 36615 14980 36668
rect 14934 36596 14980 36615
rect 14934 36547 14940 36596
rect 14974 36547 14980 36596
rect 14934 36524 14980 36547
rect 14934 36479 14940 36524
rect 14974 36479 14980 36524
rect 14934 36452 14980 36479
rect 14934 36411 14940 36452
rect 14974 36411 14980 36452
rect 14934 36380 14980 36411
rect 14934 36343 14940 36380
rect 14974 36343 14980 36380
rect 14934 36309 14980 36343
rect 14934 36274 14940 36309
rect 14974 36274 14980 36309
rect 14934 36241 14980 36274
rect 14934 36202 14940 36241
rect 14974 36202 14980 36241
rect 14934 36173 14980 36202
rect 14934 36130 14940 36173
rect 14974 36130 14980 36173
rect 14934 36105 14980 36130
rect 14934 36058 14940 36105
rect 14974 36058 14980 36105
rect 14934 36037 14980 36058
rect 14934 35986 14940 36037
rect 14974 35986 14980 36037
rect 14934 35969 14980 35986
rect 14934 35914 14940 35969
rect 14974 35914 14980 35969
rect 14934 35901 14980 35914
rect 14934 35842 14940 35901
rect 14974 35842 14980 35901
rect 14934 35833 14980 35842
rect 14934 35770 14940 35833
rect 14974 35770 14980 35833
rect 14934 35765 14980 35770
rect 14934 35698 14940 35765
rect 14974 35698 14980 35765
rect 14934 35697 14980 35698
rect 14934 35663 14940 35697
rect 14974 35663 14980 35697
rect 14934 35660 14980 35663
rect 14934 35595 14940 35660
rect 14974 35595 14980 35660
rect 14934 35588 14980 35595
rect 14934 35527 14940 35588
rect 14974 35527 14980 35588
rect 14934 35516 14980 35527
rect 14934 35459 14940 35516
rect 14974 35459 14980 35516
rect 14934 35444 14980 35459
rect 14934 35391 14940 35444
rect 14974 35391 14980 35444
rect 14934 35372 14980 35391
rect 14934 35323 14940 35372
rect 14974 35323 14980 35372
rect 14934 35300 14980 35323
rect 14934 35255 14940 35300
rect 14974 35255 14980 35300
rect 14934 35228 14980 35255
rect 14934 35187 14940 35228
rect 14974 35187 14980 35228
rect 14934 35156 14980 35187
rect 14934 35119 14940 35156
rect 14974 35119 14980 35156
rect 14934 35085 14980 35119
rect 14934 35050 14940 35085
rect 14974 35050 14980 35085
rect 14934 35017 14980 35050
rect 14934 34978 14940 35017
rect 14974 34978 14980 35017
rect 14934 34949 14980 34978
rect 14934 34906 14940 34949
rect 14974 34906 14980 34949
rect 14934 34881 14980 34906
rect 14934 34834 14940 34881
rect 14974 34834 14980 34881
rect 14934 34813 14980 34834
rect 14934 34762 14940 34813
rect 14974 34762 14980 34813
rect 14934 34745 14980 34762
rect 14934 34690 14940 34745
rect 14974 34690 14980 34745
rect 14934 34677 14980 34690
rect 14934 34618 14940 34677
rect 14974 34618 14980 34677
rect 14934 34609 14980 34618
rect 14934 34546 14940 34609
rect 14974 34546 14980 34609
rect 14934 34541 14980 34546
rect 14934 34474 14940 34541
rect 14974 34474 14980 34541
rect 14934 34473 14980 34474
rect 14934 34439 14940 34473
rect 14974 34439 14980 34473
rect 14934 34436 14980 34439
rect 14934 34371 14940 34436
rect 14974 34371 14980 34436
rect 14934 34364 14980 34371
rect 14934 34303 14940 34364
rect 14974 34303 14980 34364
rect 14934 34292 14980 34303
rect 14934 34235 14940 34292
rect 14974 34235 14980 34292
rect 14934 34220 14980 34235
rect 14934 34167 14940 34220
rect 14974 34167 14980 34220
rect 14934 34148 14980 34167
rect 14934 34099 14940 34148
rect 14974 34099 14980 34148
rect 14934 34076 14980 34099
rect 14934 34031 14940 34076
rect 14974 34031 14980 34076
rect 14934 34004 14980 34031
rect 14934 33963 14940 34004
rect 14974 33963 14980 34004
rect 14934 33932 14980 33963
rect 14934 33895 14940 33932
rect 14974 33895 14980 33932
rect 14934 33861 14980 33895
rect 14934 33826 14940 33861
rect 14974 33826 14980 33861
rect 14934 33793 14980 33826
rect 14934 33754 14940 33793
rect 14974 33754 14980 33793
rect 14934 33725 14980 33754
rect 14934 33682 14940 33725
rect 14974 33682 14980 33725
rect 14934 33657 14980 33682
rect 14934 33610 14940 33657
rect 14974 33610 14980 33657
rect 14934 33589 14980 33610
rect 14934 33538 14940 33589
rect 14974 33538 14980 33589
rect 14934 33521 14980 33538
rect 14934 33466 14940 33521
rect 14974 33466 14980 33521
rect 14934 33453 14980 33466
rect 14934 33394 14940 33453
rect 14974 33394 14980 33453
rect 14934 33385 14980 33394
rect 14934 33322 14940 33385
rect 14974 33322 14980 33385
rect 14934 33317 14980 33322
rect 14934 33250 14940 33317
rect 14974 33250 14980 33317
rect 14934 33249 14980 33250
rect 14934 33215 14940 33249
rect 14974 33215 14980 33249
rect 14934 33212 14980 33215
rect 14934 33147 14940 33212
rect 14974 33147 14980 33212
rect 14934 33140 14980 33147
rect 14934 33079 14940 33140
rect 14974 33079 14980 33140
rect 14934 33068 14980 33079
rect 14934 33011 14940 33068
rect 14974 33011 14980 33068
rect 14934 32996 14980 33011
rect 14934 32943 14940 32996
rect 14974 32943 14980 32996
rect 14934 32924 14980 32943
rect 14934 32875 14940 32924
rect 14974 32875 14980 32924
rect 14934 32852 14980 32875
rect 14934 32807 14940 32852
rect 14974 32807 14980 32852
rect 14934 32780 14980 32807
rect 14934 32739 14940 32780
rect 14974 32739 14980 32780
rect 14934 32708 14980 32739
rect 14934 32671 14940 32708
rect 14974 32671 14980 32708
rect 14934 32637 14980 32671
rect 14934 32602 14940 32637
rect 14974 32602 14980 32637
rect 14934 32569 14980 32602
rect 14934 32530 14940 32569
rect 14974 32530 14980 32569
rect 14934 32501 14980 32530
rect 14934 32458 14940 32501
rect 14974 32458 14980 32501
rect 14934 32433 14980 32458
rect 14934 32386 14940 32433
rect 14974 32386 14980 32433
rect 14934 32365 14980 32386
rect 14934 32314 14940 32365
rect 14974 32314 14980 32365
rect 14934 32297 14980 32314
rect 14934 32242 14940 32297
rect 14974 32242 14980 32297
rect 14934 32229 14980 32242
rect 14934 32170 14940 32229
rect 14974 32170 14980 32229
rect 14934 32161 14980 32170
rect 14934 32098 14940 32161
rect 14974 32098 14980 32161
rect 14934 32093 14980 32098
rect 14934 32026 14940 32093
rect 14974 32026 14980 32093
rect 14934 32025 14980 32026
rect 14934 31991 14940 32025
rect 14974 31991 14980 32025
rect 14934 31988 14980 31991
rect 14934 31923 14940 31988
rect 14974 31923 14980 31988
rect 14934 31916 14980 31923
rect 14934 31855 14940 31916
rect 14974 31855 14980 31916
rect 14934 31844 14980 31855
rect 14934 31787 14940 31844
rect 14974 31787 14980 31844
rect 14934 31772 14980 31787
rect 14934 31719 14940 31772
rect 14974 31719 14980 31772
rect 14934 31700 14980 31719
rect 14934 31651 14940 31700
rect 14974 31651 14980 31700
rect 14934 31628 14980 31651
rect 14934 31583 14940 31628
rect 14974 31583 14980 31628
rect 14934 31556 14980 31583
rect 14934 31515 14940 31556
rect 14974 31515 14980 31556
rect 14934 31484 14980 31515
rect 14934 31447 14940 31484
rect 14974 31447 14980 31484
rect 14934 31413 14980 31447
rect 14934 31378 14940 31413
rect 14974 31378 14980 31413
rect 14934 31345 14980 31378
rect 14934 31306 14940 31345
rect 14974 31306 14980 31345
rect 14934 31277 14980 31306
rect 14934 31234 14940 31277
rect 14974 31234 14980 31277
rect 14934 31209 14980 31234
rect 14934 31162 14940 31209
rect 14974 31162 14980 31209
rect 14934 31141 14980 31162
rect 14934 31090 14940 31141
rect 14974 31090 14980 31141
rect 14934 31073 14980 31090
rect 14934 31018 14940 31073
rect 14974 31018 14980 31073
rect 14934 31005 14980 31018
rect 14934 30946 14940 31005
rect 14974 30946 14980 31005
rect 14934 30937 14980 30946
rect 14934 30874 14940 30937
rect 14974 30874 14980 30937
rect 14934 30869 14980 30874
rect 14934 30802 14940 30869
rect 14974 30802 14980 30869
rect 14934 30801 14980 30802
rect 14934 30767 14940 30801
rect 14974 30767 14980 30801
rect 14934 30764 14980 30767
rect 14934 30699 14940 30764
rect 14974 30699 14980 30764
rect 14934 30692 14980 30699
rect 14934 30631 14940 30692
rect 14974 30631 14980 30692
rect 14934 30620 14980 30631
rect 14934 30563 14940 30620
rect 14974 30563 14980 30620
rect 14934 30548 14980 30563
rect 14934 30495 14940 30548
rect 14974 30495 14980 30548
rect 14934 30476 14980 30495
rect 14934 30427 14940 30476
rect 14974 30427 14980 30476
rect 14934 30404 14980 30427
rect 14934 30359 14940 30404
rect 14974 30359 14980 30404
rect 14934 30332 14980 30359
rect 14934 30291 14940 30332
rect 14974 30291 14980 30332
rect 14934 30260 14980 30291
rect 14934 30223 14940 30260
rect 14974 30223 14980 30260
rect 14934 30189 14980 30223
rect 14934 30154 14940 30189
rect 14974 30154 14980 30189
rect 14934 30121 14980 30154
rect 14934 30082 14940 30121
rect 14974 30082 14980 30121
rect 14934 30053 14980 30082
rect 14934 30010 14940 30053
rect 14974 30010 14980 30053
rect 14934 29985 14980 30010
rect 14934 29938 14940 29985
rect 14974 29938 14980 29985
rect 14934 29917 14980 29938
rect 14934 29866 14940 29917
rect 14974 29866 14980 29917
rect 14934 29849 14980 29866
rect 14934 29794 14940 29849
rect 14974 29794 14980 29849
rect 14934 29781 14980 29794
rect 14934 29722 14940 29781
rect 14974 29722 14980 29781
rect 14934 29713 14980 29722
rect 14934 29650 14940 29713
rect 14974 29650 14980 29713
rect 14934 29645 14980 29650
rect 14934 29578 14940 29645
rect 14974 29578 14980 29645
rect 14934 29577 14980 29578
rect 14934 29543 14940 29577
rect 14974 29543 14980 29577
rect 14934 29540 14980 29543
rect 14934 29475 14940 29540
rect 14974 29475 14980 29540
rect 14934 29468 14980 29475
rect 14934 29407 14940 29468
rect 14974 29407 14980 29468
rect 14934 29396 14980 29407
rect 14934 29339 14940 29396
rect 14974 29339 14980 29396
rect 14934 29324 14980 29339
rect 14934 29271 14940 29324
rect 14974 29271 14980 29324
rect 14934 29252 14980 29271
rect 14934 29203 14940 29252
rect 14974 29203 14980 29252
rect 14934 29180 14980 29203
rect 14934 29135 14940 29180
rect 14974 29135 14980 29180
rect 14934 29108 14980 29135
rect 14934 29067 14940 29108
rect 14974 29067 14980 29108
rect 14934 29036 14980 29067
rect 14934 28999 14940 29036
rect 14974 28999 14980 29036
rect 14934 28965 14980 28999
rect 14934 28930 14940 28965
rect 14974 28930 14980 28965
rect 14934 28897 14980 28930
rect 14934 28858 14940 28897
rect 14974 28858 14980 28897
rect 14934 28829 14980 28858
rect 14934 28786 14940 28829
rect 14974 28786 14980 28829
rect 14934 28761 14980 28786
rect 14934 28714 14940 28761
rect 14974 28714 14980 28761
rect 14934 28693 14980 28714
rect 14934 28642 14940 28693
rect 14974 28642 14980 28693
rect 14934 28625 14980 28642
rect 14934 28570 14940 28625
rect 14974 28570 14980 28625
rect 14934 28557 14980 28570
rect 14934 28498 14940 28557
rect 14974 28498 14980 28557
rect 14934 28489 14980 28498
rect 14934 28426 14940 28489
rect 14974 28426 14980 28489
rect 14934 28421 14980 28426
rect 14934 28354 14940 28421
rect 14974 28354 14980 28421
rect 14934 28353 14980 28354
rect 14934 28319 14940 28353
rect 14974 28319 14980 28353
rect 14934 28316 14980 28319
rect 14934 28251 14940 28316
rect 14974 28251 14980 28316
rect 14934 28244 14980 28251
rect 14934 28183 14940 28244
rect 14974 28183 14980 28244
rect 14934 28172 14980 28183
rect 14934 28115 14940 28172
rect 14974 28115 14980 28172
rect 14934 28100 14980 28115
rect 14934 28047 14940 28100
rect 14974 28047 14980 28100
rect 14934 28028 14980 28047
rect 14934 27979 14940 28028
rect 14974 27979 14980 28028
rect 14934 27956 14980 27979
rect 14934 27911 14940 27956
rect 14974 27911 14980 27956
rect 14934 27884 14980 27911
rect 14934 27843 14940 27884
rect 14974 27843 14980 27884
rect 14934 27812 14980 27843
rect 14934 27775 14940 27812
rect 14974 27775 14980 27812
rect 14934 27741 14980 27775
rect 14934 27706 14940 27741
rect 14974 27706 14980 27741
rect 14934 27673 14980 27706
rect 14934 27634 14940 27673
rect 14974 27634 14980 27673
rect 14934 27605 14980 27634
rect 14934 27562 14940 27605
rect 14974 27562 14980 27605
rect 14934 27537 14980 27562
rect 14934 27490 14940 27537
rect 14974 27490 14980 27537
rect 14934 27469 14980 27490
rect 14934 27418 14940 27469
rect 14974 27418 14980 27469
rect 14934 27401 14980 27418
rect 14934 27346 14940 27401
rect 14974 27346 14980 27401
rect 14934 27333 14980 27346
rect 14934 27274 14940 27333
rect 14974 27274 14980 27333
rect 14934 27265 14980 27274
rect 14934 27202 14940 27265
rect 14974 27202 14980 27265
rect 14934 27197 14980 27202
rect 14934 27130 14940 27197
rect 14974 27130 14980 27197
rect 14934 27129 14980 27130
rect 14934 27095 14940 27129
rect 14974 27095 14980 27129
rect 14934 27092 14980 27095
rect 14934 27027 14940 27092
rect 14974 27027 14980 27092
rect 14934 27020 14980 27027
rect 14934 26959 14940 27020
rect 14974 26959 14980 27020
rect 14934 26948 14980 26959
rect 14934 26891 14940 26948
rect 14974 26891 14980 26948
rect 14934 26876 14980 26891
rect 14934 26823 14940 26876
rect 14974 26823 14980 26876
rect 14934 26804 14980 26823
rect 14934 26755 14940 26804
rect 14974 26755 14980 26804
rect 14934 26732 14980 26755
rect 14934 26687 14940 26732
rect 14974 26687 14980 26732
rect 14934 26660 14980 26687
rect 14934 26619 14940 26660
rect 14974 26619 14980 26660
rect 14934 26588 14980 26619
rect 14934 26551 14940 26588
rect 14974 26551 14980 26588
rect 14934 26517 14980 26551
rect 14934 26482 14940 26517
rect 14974 26482 14980 26517
rect 14934 26449 14980 26482
rect 14934 26410 14940 26449
rect 14974 26410 14980 26449
rect 14934 26381 14980 26410
rect 14934 26338 14940 26381
rect 14974 26338 14980 26381
rect 14934 26313 14980 26338
rect 14934 26266 14940 26313
rect 14974 26266 14980 26313
rect 14934 26245 14980 26266
rect 14934 26194 14940 26245
rect 14974 26194 14980 26245
rect 14934 26177 14980 26194
rect 14934 26122 14940 26177
rect 14974 26122 14980 26177
rect 14934 26109 14980 26122
rect 14934 26050 14940 26109
rect 14974 26050 14980 26109
rect 14934 26041 14980 26050
rect 14934 25978 14940 26041
rect 14974 25978 14980 26041
rect 14934 25973 14980 25978
rect 14934 25906 14940 25973
rect 14974 25906 14980 25973
rect 14934 25905 14980 25906
rect 14934 25871 14940 25905
rect 14974 25871 14980 25905
rect 14934 25868 14980 25871
rect 14934 25803 14940 25868
rect 14974 25803 14980 25868
rect 14934 25796 14980 25803
rect 14934 25735 14940 25796
rect 14974 25735 14980 25796
rect 14934 25724 14980 25735
rect 14934 25667 14940 25724
rect 14974 25667 14980 25724
rect 14934 25652 14980 25667
rect 14934 25599 14940 25652
rect 14974 25599 14980 25652
rect 14934 25580 14980 25599
rect 14934 25531 14940 25580
rect 14974 25531 14980 25580
rect 14934 25508 14980 25531
rect 14934 25463 14940 25508
rect 14974 25463 14980 25508
rect 14934 25436 14980 25463
rect 14934 25395 14940 25436
rect 14974 25395 14980 25436
rect 14934 25364 14980 25395
rect 14934 25327 14940 25364
rect 14974 25327 14980 25364
rect 14934 25293 14980 25327
rect 14934 25258 14940 25293
rect 14974 25258 14980 25293
rect 14934 25225 14980 25258
rect 14934 25186 14940 25225
rect 14974 25186 14980 25225
rect 14934 25157 14980 25186
rect 14934 25114 14940 25157
rect 14974 25114 14980 25157
rect 14934 25089 14980 25114
rect 14934 25042 14940 25089
rect 14974 25042 14980 25089
rect 14934 25021 14980 25042
rect 14934 24970 14940 25021
rect 14974 24970 14980 25021
rect 14934 24953 14980 24970
rect 14934 24898 14940 24953
rect 14974 24898 14980 24953
rect 14934 24885 14980 24898
rect 14934 24826 14940 24885
rect 14974 24826 14980 24885
rect 14934 24817 14980 24826
rect 14934 24754 14940 24817
rect 14974 24754 14980 24817
rect 14934 24749 14980 24754
rect 14934 24682 14940 24749
rect 14974 24682 14980 24749
rect 14934 24681 14980 24682
rect 14934 24647 14940 24681
rect 14974 24647 14980 24681
rect 14934 24644 14980 24647
rect 14934 24579 14940 24644
rect 14974 24579 14980 24644
rect 14934 24572 14980 24579
rect 14934 24511 14940 24572
rect 14974 24511 14980 24572
rect 14934 24500 14980 24511
rect 14934 24443 14940 24500
rect 14974 24443 14980 24500
rect 14934 24428 14980 24443
rect 14934 24375 14940 24428
rect 14974 24375 14980 24428
rect 14934 24356 14980 24375
rect 14934 24307 14940 24356
rect 14974 24307 14980 24356
rect 14934 24284 14980 24307
rect 14934 24239 14940 24284
rect 14974 24239 14980 24284
rect 14934 24212 14980 24239
rect 14934 24171 14940 24212
rect 14974 24171 14980 24212
rect 14934 24140 14980 24171
rect 14934 24103 14940 24140
rect 14974 24103 14980 24140
rect 14934 24069 14980 24103
rect 14934 24034 14940 24069
rect 14974 24034 14980 24069
rect 14934 24001 14980 24034
rect 14934 23962 14940 24001
rect 14974 23962 14980 24001
rect 14934 23933 14980 23962
rect 14934 23890 14940 23933
rect 14974 23890 14980 23933
rect 14934 23865 14980 23890
rect 14934 23818 14940 23865
rect 14974 23818 14980 23865
rect 14934 23797 14980 23818
rect 14934 23746 14940 23797
rect 14974 23746 14980 23797
rect 14934 23729 14980 23746
rect 14934 23674 14940 23729
rect 14974 23674 14980 23729
rect 14934 23661 14980 23674
rect 14934 23602 14940 23661
rect 14974 23602 14980 23661
rect 14934 23593 14980 23602
rect 14934 23530 14940 23593
rect 14974 23530 14980 23593
rect 14934 23525 14980 23530
rect 14934 23458 14940 23525
rect 14974 23458 14980 23525
rect 14934 23457 14980 23458
rect 14934 23423 14940 23457
rect 14974 23423 14980 23457
rect 14934 23420 14980 23423
rect 14934 23355 14940 23420
rect 14974 23355 14980 23420
rect 14934 23348 14980 23355
rect 14934 23287 14940 23348
rect 14974 23287 14980 23348
rect 14934 23276 14980 23287
rect 14934 23219 14940 23276
rect 14974 23219 14980 23276
rect 14934 23204 14980 23219
rect 14934 23151 14940 23204
rect 14974 23151 14980 23204
rect 14934 23132 14980 23151
rect 14934 23083 14940 23132
rect 14974 23083 14980 23132
rect 14934 23060 14980 23083
rect 14934 23015 14940 23060
rect 14974 23015 14980 23060
rect 14934 22988 14980 23015
rect 14934 22947 14940 22988
rect 14974 22947 14980 22988
rect 14934 22916 14980 22947
rect 14934 22879 14940 22916
rect 14974 22879 14980 22916
rect 14934 22845 14980 22879
rect 14934 22810 14940 22845
rect 14974 22810 14980 22845
rect 14934 22777 14980 22810
rect 14934 22738 14940 22777
rect 14974 22738 14980 22777
rect 14934 22709 14980 22738
rect 14934 22666 14940 22709
rect 14974 22666 14980 22709
rect 14934 22641 14980 22666
rect 14934 22594 14940 22641
rect 14974 22594 14980 22641
rect 14934 22573 14980 22594
rect 14934 22522 14940 22573
rect 14974 22522 14980 22573
rect 14934 22505 14980 22522
rect 14934 22450 14940 22505
rect 14974 22450 14980 22505
rect 14934 22437 14980 22450
rect 14934 22378 14940 22437
rect 14974 22378 14980 22437
rect 14934 22369 14980 22378
rect 14934 22306 14940 22369
rect 14974 22306 14980 22369
rect 14934 22301 14980 22306
rect 14934 22234 14940 22301
rect 14974 22234 14980 22301
rect 14934 22233 14980 22234
rect 14934 22199 14940 22233
rect 14974 22199 14980 22233
rect 14934 22196 14980 22199
rect 14934 22131 14940 22196
rect 14974 22131 14980 22196
rect 14934 22124 14980 22131
rect 14934 22063 14940 22124
rect 14974 22063 14980 22124
rect 14934 22052 14980 22063
rect 14934 21995 14940 22052
rect 14974 21995 14980 22052
rect 14934 21980 14980 21995
rect 14934 21927 14940 21980
rect 14974 21927 14980 21980
rect 14934 21908 14980 21927
rect 14934 21859 14940 21908
rect 14974 21859 14980 21908
rect 14934 21836 14980 21859
rect 14934 21791 14940 21836
rect 14974 21791 14980 21836
rect 14934 21764 14980 21791
rect 14934 21723 14940 21764
rect 14974 21723 14980 21764
rect 14934 21692 14980 21723
rect 14934 21655 14940 21692
rect 14974 21655 14980 21692
rect 14934 21621 14980 21655
rect 14934 21586 14940 21621
rect 14974 21586 14980 21621
rect 14934 21553 14980 21586
rect 14934 21514 14940 21553
rect 14974 21514 14980 21553
rect 14934 21485 14980 21514
rect 14934 21442 14940 21485
rect 14974 21442 14980 21485
rect 14934 21417 14980 21442
rect 14934 21370 14940 21417
rect 14974 21370 14980 21417
rect 14934 21349 14980 21370
rect 14934 21298 14940 21349
rect 14974 21298 14980 21349
rect 14934 21281 14980 21298
rect 14934 21226 14940 21281
rect 14974 21226 14980 21281
rect 14934 21213 14980 21226
rect 14934 21154 14940 21213
rect 14974 21154 14980 21213
rect 14934 21145 14980 21154
rect 14934 21082 14940 21145
rect 14974 21082 14980 21145
rect 14934 21077 14980 21082
rect 14934 21010 14940 21077
rect 14974 21010 14980 21077
rect 14934 21009 14980 21010
rect 14934 20975 14940 21009
rect 14974 20975 14980 21009
rect 14934 20972 14980 20975
rect 14934 20907 14940 20972
rect 14974 20907 14980 20972
rect 14934 20900 14980 20907
rect 14934 20839 14940 20900
rect 14974 20839 14980 20900
rect 14934 20828 14980 20839
rect 14934 20771 14940 20828
rect 14974 20771 14980 20828
rect 14934 20756 14980 20771
rect 14934 20703 14940 20756
rect 14974 20703 14980 20756
rect 14934 20684 14980 20703
rect 14934 20635 14940 20684
rect 14974 20635 14980 20684
rect 14934 20612 14980 20635
rect 14934 20567 14940 20612
rect 14974 20567 14980 20612
rect 14934 20540 14980 20567
rect 14934 20499 14940 20540
rect 14974 20499 14980 20540
rect 14934 20468 14980 20499
rect 14934 20431 14940 20468
rect 14974 20431 14980 20468
rect 14934 20397 14980 20431
rect 14934 20362 14940 20397
rect 14974 20362 14980 20397
rect 14934 20329 14980 20362
rect 14934 20290 14940 20329
rect 14974 20290 14980 20329
rect 14934 20261 14980 20290
rect 14934 20218 14940 20261
rect 14974 20218 14980 20261
rect 14934 20193 14980 20218
rect 14934 20146 14940 20193
rect 14974 20146 14980 20193
rect 14934 20125 14980 20146
rect 14934 20074 14940 20125
rect 14974 20074 14980 20125
rect 14934 20057 14980 20074
rect 14934 20002 14940 20057
rect 14974 20002 14980 20057
rect 14934 19989 14980 20002
rect 14934 19930 14940 19989
rect 14974 19930 14980 19989
rect 14934 19921 14980 19930
rect 14934 19858 14940 19921
rect 14974 19858 14980 19921
rect 14934 19853 14980 19858
rect 14934 19786 14940 19853
rect 14974 19786 14980 19853
rect 14934 19785 14980 19786
rect 14934 19751 14940 19785
rect 14974 19751 14980 19785
rect 14934 19748 14980 19751
rect 14934 19683 14940 19748
rect 14974 19683 14980 19748
rect 14934 19676 14980 19683
rect 14934 19615 14940 19676
rect 14974 19615 14980 19676
rect 14934 19604 14980 19615
rect 14934 19547 14940 19604
rect 14974 19547 14980 19604
rect 14934 19532 14980 19547
rect 14934 19479 14940 19532
rect 14974 19479 14980 19532
rect 14934 19460 14980 19479
rect 14934 19411 14940 19460
rect 14974 19411 14980 19460
rect 14934 19388 14980 19411
rect 14934 19343 14940 19388
rect 14974 19343 14980 19388
rect 14934 19316 14980 19343
rect 14934 19275 14940 19316
rect 14974 19275 14980 19316
rect 14934 19244 14980 19275
rect 14934 19207 14940 19244
rect 14974 19207 14980 19244
rect 14934 19173 14980 19207
rect 14934 19138 14940 19173
rect 14974 19138 14980 19173
rect 14934 19105 14980 19138
rect 14934 19066 14940 19105
rect 14974 19066 14980 19105
rect 14934 19037 14980 19066
rect 14934 18994 14940 19037
rect 14974 18994 14980 19037
rect 14934 18969 14980 18994
rect 14934 18922 14940 18969
rect 14974 18922 14980 18969
rect 14934 18901 14980 18922
rect 14934 18850 14940 18901
rect 14974 18850 14980 18901
rect 14934 18833 14980 18850
rect 14934 18778 14940 18833
rect 14974 18778 14980 18833
rect 14934 18765 14980 18778
rect 14934 18706 14940 18765
rect 14974 18706 14980 18765
rect 14934 18697 14980 18706
rect 14934 18634 14940 18697
rect 14974 18634 14980 18697
rect 14934 18629 14980 18634
rect 14934 18562 14940 18629
rect 14974 18562 14980 18629
rect 14934 18561 14980 18562
rect 14934 18527 14940 18561
rect 14974 18527 14980 18561
rect 14934 18524 14980 18527
rect 14934 18459 14940 18524
rect 14974 18459 14980 18524
rect 14934 18452 14980 18459
rect 14934 18391 14940 18452
rect 14974 18391 14980 18452
rect 14934 18380 14980 18391
rect 14934 18323 14940 18380
rect 14974 18323 14980 18380
rect 14934 18308 14980 18323
rect 14934 18255 14940 18308
rect 14974 18255 14980 18308
rect 14934 18236 14980 18255
rect 14934 18187 14940 18236
rect 14974 18187 14980 18236
rect 14934 18164 14980 18187
rect 14934 18119 14940 18164
rect 14974 18119 14980 18164
rect 14934 18092 14980 18119
rect 14934 18051 14940 18092
rect 14974 18051 14980 18092
rect 14934 18020 14980 18051
rect 14934 17983 14940 18020
rect 14974 17983 14980 18020
rect 14934 17949 14980 17983
rect 14934 17914 14940 17949
rect 14974 17914 14980 17949
rect 14934 17881 14980 17914
rect 14934 17842 14940 17881
rect 14974 17842 14980 17881
rect 14934 17813 14980 17842
rect 14934 17770 14940 17813
rect 14974 17770 14980 17813
rect 14934 17745 14980 17770
rect 14934 17698 14940 17745
rect 14974 17698 14980 17745
rect 14934 17677 14980 17698
rect 14934 17626 14940 17677
rect 14974 17626 14980 17677
rect 14934 17609 14980 17626
rect 14934 17554 14940 17609
rect 14974 17554 14980 17609
rect 14934 17541 14980 17554
rect 14934 17482 14940 17541
rect 14974 17482 14980 17541
rect 14934 17473 14980 17482
rect 14934 17410 14940 17473
rect 14974 17410 14980 17473
rect 14934 17405 14980 17410
rect 14934 17338 14940 17405
rect 14974 17338 14980 17405
rect 14934 17337 14980 17338
rect 14934 17303 14940 17337
rect 14974 17303 14980 17337
rect 14934 17300 14980 17303
rect 14934 17235 14940 17300
rect 14974 17235 14980 17300
rect 14934 17228 14980 17235
rect 14934 17167 14940 17228
rect 14974 17167 14980 17228
rect 14934 17156 14980 17167
rect 14934 17099 14940 17156
rect 14974 17099 14980 17156
rect 14934 17084 14980 17099
rect 14934 17031 14940 17084
rect 14974 17031 14980 17084
rect 14934 17012 14980 17031
rect 14934 16963 14940 17012
rect 14974 16963 14980 17012
rect 14934 16940 14980 16963
rect 14934 16895 14940 16940
rect 14974 16895 14980 16940
rect 14934 16868 14980 16895
rect 14934 16827 14940 16868
rect 14974 16827 14980 16868
rect 14934 16796 14980 16827
rect 14934 16759 14940 16796
rect 14974 16759 14980 16796
rect 14934 16725 14980 16759
rect 14934 16690 14940 16725
rect 14974 16690 14980 16725
rect 14934 16657 14980 16690
rect 14934 16618 14940 16657
rect 14974 16618 14980 16657
rect 14934 16589 14980 16618
rect 14934 16546 14940 16589
rect 14974 16546 14980 16589
rect 14934 16521 14980 16546
rect 14934 16474 14940 16521
rect 14974 16474 14980 16521
rect 14934 16453 14980 16474
rect 14934 16402 14940 16453
rect 14974 16402 14980 16453
rect 14934 16385 14980 16402
rect 14934 16330 14940 16385
rect 14974 16330 14980 16385
rect 14934 16317 14980 16330
rect 14934 16258 14940 16317
rect 14974 16258 14980 16317
rect 14934 16249 14980 16258
rect 14934 16186 14940 16249
rect 14974 16186 14980 16249
rect 14934 16181 14980 16186
rect 14934 16114 14940 16181
rect 14974 16114 14980 16181
rect 14934 16113 14980 16114
rect 14934 16079 14940 16113
rect 14974 16079 14980 16113
rect 14934 16076 14980 16079
rect 14934 16011 14940 16076
rect 14974 16011 14980 16076
rect 14934 16004 14980 16011
rect 14934 15943 14940 16004
rect 14974 15943 14980 16004
rect 14934 15932 14980 15943
rect 14934 15875 14940 15932
rect 14974 15875 14980 15932
rect 14934 15860 14980 15875
rect 14934 15807 14940 15860
rect 14974 15807 14980 15860
rect 14934 15788 14980 15807
rect 14934 15739 14940 15788
rect 14974 15739 14980 15788
rect 14934 15716 14980 15739
rect 14934 15671 14940 15716
rect 14974 15671 14980 15716
rect 14934 15644 14980 15671
rect 14934 15603 14940 15644
rect 14974 15603 14980 15644
rect 14934 15572 14980 15603
rect 14934 15535 14940 15572
rect 14974 15535 14980 15572
rect 14934 15501 14980 15535
rect 14934 15466 14940 15501
rect 14974 15466 14980 15501
rect 14934 15433 14980 15466
rect 14934 15394 14940 15433
rect 14974 15394 14980 15433
rect 14934 15365 14980 15394
rect 14934 15322 14940 15365
rect 14974 15322 14980 15365
rect 14934 15297 14980 15322
rect 14934 15250 14940 15297
rect 14974 15250 14980 15297
rect 14934 15229 14980 15250
rect 14934 15178 14940 15229
rect 14974 15178 14980 15229
rect 14934 15161 14980 15178
rect 14934 15106 14940 15161
rect 14974 15106 14980 15161
rect 14934 15093 14980 15106
rect 14934 15034 14940 15093
rect 14974 15034 14980 15093
rect 14934 15025 14980 15034
rect 14934 14962 14940 15025
rect 14974 14962 14980 15025
rect 14934 14957 14980 14962
rect 14934 14890 14940 14957
rect 14974 14890 14980 14957
rect 14934 14889 14980 14890
rect 14934 14855 14940 14889
rect 14974 14855 14980 14889
rect 14934 14852 14980 14855
rect 14934 14787 14940 14852
rect 14974 14787 14980 14852
rect 14934 14780 14980 14787
rect 14934 14719 14940 14780
rect 14974 14719 14980 14780
rect 14934 14708 14980 14719
rect 14934 14651 14940 14708
rect 14974 14651 14980 14708
rect 14934 14636 14980 14651
rect 14934 14583 14940 14636
rect 14974 14583 14980 14636
rect 14934 14564 14980 14583
rect 14934 14515 14940 14564
rect 14974 14515 14980 14564
rect 14934 14492 14980 14515
rect 14934 14447 14940 14492
rect 14974 14447 14980 14492
rect 14934 14420 14980 14447
rect 14934 14379 14940 14420
rect 14974 14379 14980 14420
rect 14934 14348 14980 14379
rect 14934 14311 14940 14348
rect 14974 14311 14980 14348
rect 14934 14277 14980 14311
rect 14934 14242 14940 14277
rect 14974 14242 14980 14277
rect 14934 14209 14980 14242
rect 14934 14170 14940 14209
rect 14974 14170 14980 14209
rect 14934 14141 14980 14170
rect 14934 14098 14940 14141
rect 14974 14098 14980 14141
rect 14934 14073 14980 14098
rect 14934 14026 14940 14073
rect 14974 14026 14980 14073
rect 14934 14005 14980 14026
rect 14934 13954 14940 14005
rect 14974 13954 14980 14005
rect 14934 13937 14980 13954
rect 14934 13882 14940 13937
rect 14974 13882 14980 13937
rect 14934 13869 14980 13882
rect 14934 13810 14940 13869
rect 14974 13810 14980 13869
rect 14934 13801 14980 13810
rect 14934 13738 14940 13801
rect 14974 13738 14980 13801
rect 14934 13733 14980 13738
rect 14934 13666 14940 13733
rect 14974 13666 14980 13733
rect 14934 13665 14980 13666
rect 14934 13631 14940 13665
rect 14974 13631 14980 13665
rect 14934 13628 14980 13631
rect 14934 13563 14940 13628
rect 14974 13563 14980 13628
rect 14934 13556 14980 13563
rect 14934 13495 14940 13556
rect 14974 13495 14980 13556
rect 14934 13484 14980 13495
rect 14934 13427 14940 13484
rect 14974 13427 14980 13484
rect 14934 13412 14980 13427
rect 14934 13359 14940 13412
rect 14974 13359 14980 13412
rect 14934 13340 14980 13359
rect 14934 13291 14940 13340
rect 14974 13291 14980 13340
rect 14934 13268 14980 13291
rect 14934 13223 14940 13268
rect 14974 13223 14980 13268
rect 14934 13196 14980 13223
rect 14934 13155 14940 13196
rect 14974 13155 14980 13196
rect 14934 13124 14980 13155
rect 14934 13087 14940 13124
rect 14974 13087 14980 13124
rect 14934 13053 14980 13087
rect 14934 13018 14940 13053
rect 14974 13018 14980 13053
rect 14934 12985 14980 13018
rect 14934 12946 14940 12985
rect 14974 12946 14980 12985
rect 14934 12917 14980 12946
rect 14934 12874 14940 12917
rect 14974 12874 14980 12917
rect 14934 12849 14980 12874
rect 14934 12802 14940 12849
rect 14974 12802 14980 12849
rect 14934 12781 14980 12802
rect 14934 12730 14940 12781
rect 14974 12730 14980 12781
rect 14934 12713 14980 12730
rect 14934 12658 14940 12713
rect 14974 12658 14980 12713
rect 14934 12645 14980 12658
rect 14934 12586 14940 12645
rect 14974 12586 14980 12645
rect 14934 12577 14980 12586
rect 14934 12514 14940 12577
rect 14974 12514 14980 12577
rect 14934 12509 14980 12514
rect 14934 12442 14940 12509
rect 14974 12442 14980 12509
rect 14934 12441 14980 12442
rect 14934 12407 14940 12441
rect 14974 12407 14980 12441
rect 14934 12404 14980 12407
rect 14934 12339 14940 12404
rect 14974 12339 14980 12404
rect 14934 12332 14980 12339
rect 14934 12271 14940 12332
rect 14974 12271 14980 12332
rect 14934 12260 14980 12271
rect 14934 12203 14940 12260
rect 14974 12203 14980 12260
rect 14934 12188 14980 12203
rect 14934 12135 14940 12188
rect 14974 12135 14980 12188
rect 14934 12116 14980 12135
rect 14934 12067 14940 12116
rect 14974 12067 14980 12116
rect 14934 12044 14980 12067
rect 14934 11999 14940 12044
rect 14974 11999 14980 12044
rect 14934 11972 14980 11999
rect 14934 11931 14940 11972
rect 14974 11931 14980 11972
rect 14934 11900 14980 11931
rect 14934 11863 14940 11900
rect 14974 11863 14980 11900
rect 14934 11829 14980 11863
rect 14934 11794 14940 11829
rect 14974 11794 14980 11829
rect 14934 11761 14980 11794
rect 14934 11722 14940 11761
rect 14974 11722 14980 11761
rect 14934 11693 14980 11722
rect 14934 11650 14940 11693
rect 14974 11650 14980 11693
rect 14934 11625 14980 11650
rect 14934 11578 14940 11625
rect 14974 11578 14980 11625
rect 14934 11557 14980 11578
rect 14934 11506 14940 11557
rect 14974 11506 14980 11557
rect 14934 11489 14980 11506
rect 14934 11434 14940 11489
rect 14974 11434 14980 11489
rect 14934 11421 14980 11434
rect 14934 11362 14940 11421
rect 14974 11362 14980 11421
rect 14934 11353 14980 11362
rect 14934 11290 14940 11353
rect 14974 11290 14980 11353
rect 14934 11285 14980 11290
rect 14934 11218 14940 11285
rect 14974 11218 14980 11285
rect 14934 11217 14980 11218
rect 14934 11183 14940 11217
rect 14974 11183 14980 11217
rect 14934 11180 14980 11183
rect 14934 11115 14940 11180
rect 14974 11115 14980 11180
rect 14934 11108 14980 11115
rect 14934 11047 14940 11108
rect 14974 11047 14980 11108
rect 14934 11036 14980 11047
rect 14934 10979 14940 11036
rect 14974 10979 14980 11036
rect 14934 10964 14980 10979
rect 14934 10911 14940 10964
rect 14974 10911 14980 10964
rect 14934 10892 14980 10911
rect 14934 10843 14940 10892
rect 14974 10843 14980 10892
rect 14934 10820 14980 10843
rect 14934 10775 14940 10820
rect 14974 10775 14980 10820
rect 14934 10748 14980 10775
rect 14934 10707 14940 10748
rect 14974 10707 14980 10748
rect 14934 10676 14980 10707
rect 14934 10639 14940 10676
rect 14974 10639 14980 10676
rect 14934 10605 14980 10639
rect 14934 10570 14940 10605
rect 14974 10570 14980 10605
rect 14934 10537 14980 10570
rect 14934 10498 14940 10537
rect 14974 10498 14980 10537
rect 14934 10469 14980 10498
rect 14934 10426 14940 10469
rect 14974 10426 14980 10469
rect 14934 10401 14980 10426
rect 14934 10354 14940 10401
rect 14974 10354 14980 10401
rect 14934 10333 14980 10354
rect 14934 10282 14940 10333
rect 14974 10282 14980 10333
rect 14934 10265 14980 10282
rect 14934 10210 14940 10265
rect 14974 10210 14980 10265
rect 14934 10197 14980 10210
rect 14934 10138 14940 10197
rect 14974 10138 14980 10197
rect 14934 10129 14980 10138
rect 14934 10066 14940 10129
rect 14974 10066 14980 10129
rect 14934 10061 14980 10066
rect 14934 9994 14940 10061
rect 14974 9994 14980 10061
rect 14934 9993 14980 9994
rect 14934 9959 14940 9993
rect 14974 9959 14980 9993
rect 14934 9956 14980 9959
rect 14934 9891 14940 9956
rect 14974 9891 14980 9956
rect 14934 9884 14980 9891
rect 14934 9823 14940 9884
rect 14974 9823 14980 9884
rect 14934 9812 14980 9823
rect 14934 9755 14940 9812
rect 14974 9755 14980 9812
rect 14934 9740 14980 9755
rect 14934 9687 14940 9740
rect 14974 9687 14980 9740
rect 14934 9668 14980 9687
rect 14934 9619 14940 9668
rect 14974 9619 14980 9668
rect 14934 9596 14980 9619
rect 14934 9551 14940 9596
rect 14974 9551 14980 9596
rect 14934 9524 14980 9551
rect 14934 9483 14940 9524
rect 14974 9483 14980 9524
rect 14934 9452 14980 9483
rect 14934 9415 14940 9452
rect 14974 9415 14980 9452
rect 14934 9381 14980 9415
rect 14934 9346 14940 9381
rect 14974 9346 14980 9381
rect 14934 9313 14980 9346
rect 14934 9274 14940 9313
rect 14974 9274 14980 9313
rect 14934 9245 14980 9274
rect 14934 9202 14940 9245
rect 14974 9202 14980 9245
rect 14934 9177 14980 9202
rect 14934 9130 14940 9177
rect 14974 9130 14980 9177
rect 14934 9109 14980 9130
rect 14934 9058 14940 9109
rect 14974 9058 14980 9109
rect 14934 9041 14980 9058
rect 14934 8986 14940 9041
rect 14974 8986 14980 9041
rect 14934 8973 14980 8986
rect 14934 8914 14940 8973
rect 14974 8914 14980 8973
rect 14934 8905 14980 8914
rect 14934 8842 14940 8905
rect 14974 8842 14980 8905
rect 14934 8837 14980 8842
rect 14934 8770 14940 8837
rect 14974 8770 14980 8837
rect 14934 8769 14980 8770
rect 14934 8735 14940 8769
rect 14974 8735 14980 8769
rect 14934 8732 14980 8735
rect 14934 8667 14940 8732
rect 14974 8667 14980 8732
rect 14934 8660 14980 8667
rect 14934 8599 14940 8660
rect 14974 8599 14980 8660
rect 14934 8588 14980 8599
rect 14934 8531 14940 8588
rect 14974 8531 14980 8588
rect 14934 8516 14980 8531
rect 14934 8463 14940 8516
rect 14974 8463 14980 8516
rect 14934 8444 14980 8463
rect 14934 8395 14940 8444
rect 14974 8395 14980 8444
rect 14934 8372 14980 8395
rect 14934 8327 14940 8372
rect 14974 8327 14980 8372
rect 14934 8300 14980 8327
rect 14934 8259 14940 8300
rect 14974 8259 14980 8300
rect 14934 8228 14980 8259
rect 14934 8191 14940 8228
rect 14974 8191 14980 8228
rect 14934 8157 14980 8191
rect 14934 8122 14940 8157
rect 14974 8122 14980 8157
rect 14934 8089 14980 8122
rect 14934 8050 14940 8089
rect 14974 8050 14980 8089
rect 14934 8021 14980 8050
rect 14934 7978 14940 8021
rect 14974 7978 14980 8021
rect 14934 7953 14980 7978
rect 14934 7906 14940 7953
rect 14974 7906 14980 7953
rect 14934 7885 14980 7906
rect 14934 7834 14940 7885
rect 14974 7834 14980 7885
rect 14934 7817 14980 7834
rect 14934 7762 14940 7817
rect 14974 7762 14980 7817
rect 14934 7749 14980 7762
rect 14934 7690 14940 7749
rect 14974 7690 14980 7749
rect 14934 7681 14980 7690
rect 14934 7618 14940 7681
rect 14974 7618 14980 7681
rect 14934 7613 14980 7618
rect 14934 7546 14940 7613
rect 14974 7546 14980 7613
rect 14934 7545 14980 7546
rect 14934 7511 14940 7545
rect 14974 7511 14980 7545
rect 14934 7508 14980 7511
rect 14934 7443 14940 7508
rect 14974 7443 14980 7508
rect 14934 7436 14980 7443
rect 14934 7375 14940 7436
rect 14974 7375 14980 7436
rect 14934 7364 14980 7375
rect 14934 7307 14940 7364
rect 14974 7307 14980 7364
rect 14934 7292 14980 7307
rect 14934 7239 14940 7292
rect 14974 7239 14980 7292
rect 14934 7220 14980 7239
rect 14934 7171 14940 7220
rect 14974 7171 14980 7220
rect 14934 7148 14980 7171
rect 14934 7103 14940 7148
rect 14974 7103 14980 7148
rect 14934 7076 14980 7103
rect 14934 7035 14940 7076
rect 14974 7035 14980 7076
rect 14934 7004 14980 7035
rect 14934 6967 14940 7004
rect 14974 6967 14980 7004
rect 14934 6933 14980 6967
rect 14934 6898 14940 6933
rect 14974 6898 14980 6933
rect 14934 6865 14980 6898
rect 14934 6826 14940 6865
rect 14974 6826 14980 6865
rect 14934 6797 14980 6826
rect 14934 6754 14940 6797
rect 14974 6754 14980 6797
rect 14934 6729 14980 6754
rect 14934 6682 14940 6729
rect 14974 6682 14980 6729
rect 14934 6661 14980 6682
rect 14934 6610 14940 6661
rect 14974 6610 14980 6661
rect 14934 6593 14980 6610
rect 14934 6538 14940 6593
rect 14974 6538 14980 6593
rect 14934 6525 14980 6538
rect 14934 6466 14940 6525
rect 14974 6466 14980 6525
rect 14934 6457 14980 6466
rect 14934 6394 14940 6457
rect 14974 6394 14980 6457
rect 14934 6389 14980 6394
rect 14934 6322 14940 6389
rect 14974 6322 14980 6389
rect 14934 6321 14980 6322
rect 14934 6287 14940 6321
rect 14974 6287 14980 6321
rect 14934 6284 14980 6287
rect 14934 6219 14940 6284
rect 14974 6219 14980 6284
rect 14934 6212 14980 6219
rect 14934 6151 14940 6212
rect 14974 6151 14980 6212
rect 14934 6140 14980 6151
rect 14934 6083 14940 6140
rect 14974 6083 14980 6140
rect 14934 6068 14980 6083
rect 14934 6015 14940 6068
rect 14974 6015 14980 6068
rect 14934 5996 14980 6015
rect 14934 5947 14940 5996
rect 14974 5947 14980 5996
rect 14934 5924 14980 5947
rect 14934 5879 14940 5924
rect 14974 5879 14980 5924
rect 14934 5852 14980 5879
rect 14934 5811 14940 5852
rect 14974 5811 14980 5852
rect 14934 5780 14980 5811
rect 14934 5743 14940 5780
rect 14974 5743 14980 5780
rect 14934 5709 14980 5743
rect 14934 5674 14940 5709
rect 14974 5674 14980 5709
rect 14934 5641 14980 5674
rect 14934 5602 14940 5641
rect 14974 5602 14980 5641
rect 14934 5573 14980 5602
rect 14934 5530 14940 5573
rect 14974 5530 14980 5573
rect 14934 5505 14980 5530
rect 14934 5458 14940 5505
rect 14974 5458 14980 5505
rect 14934 5437 14980 5458
rect 14934 5386 14940 5437
rect 14974 5386 14980 5437
rect 14934 5369 14980 5386
rect 14934 5314 14940 5369
rect 14974 5314 14980 5369
rect 14934 5301 14980 5314
rect 14934 5242 14940 5301
rect 14974 5242 14980 5301
rect 14934 5233 14980 5242
rect 14934 5170 14940 5233
rect 14974 5170 14980 5233
rect 14934 5165 14980 5170
rect 14934 5098 14940 5165
rect 14974 5098 14980 5165
rect 14934 5097 14980 5098
rect 14934 5063 14940 5097
rect 14974 5063 14980 5097
rect 14934 5060 14980 5063
rect 14934 4995 14940 5060
rect 14974 4995 14980 5060
rect 14934 4988 14980 4995
rect 14934 4927 14940 4988
rect 14974 4927 14980 4988
rect 14934 4916 14980 4927
rect 14934 4859 14940 4916
rect 14974 4859 14980 4916
rect 14934 4844 14980 4859
rect 14934 4791 14940 4844
rect 14974 4791 14980 4844
rect 14934 4772 14980 4791
rect 14934 4723 14940 4772
rect 14974 4723 14980 4772
rect 14934 4700 14980 4723
rect 14934 4655 14940 4700
rect 14974 4655 14980 4700
rect 14934 4628 14980 4655
rect 14934 4587 14940 4628
rect 14974 4587 14980 4628
rect 14934 4556 14980 4587
rect 14934 4519 14940 4556
rect 14974 4519 14980 4556
rect 14934 4485 14980 4519
rect 14934 4450 14940 4485
rect 14974 4450 14980 4485
rect 14934 4417 14980 4450
rect 14934 4378 14940 4417
rect 14974 4378 14980 4417
rect 14934 4349 14980 4378
rect 14934 4306 14940 4349
rect 14974 4306 14980 4349
rect 14934 4281 14980 4306
rect 14934 4234 14940 4281
rect 14974 4234 14980 4281
rect 14934 4213 14980 4234
rect 14934 4162 14940 4213
rect 14974 4162 14980 4213
rect 14934 4145 14980 4162
rect 14934 4090 14940 4145
rect 14974 4090 14980 4145
rect 14934 4077 14980 4090
rect 14934 4018 14940 4077
rect 14974 4018 14980 4077
rect 14934 4009 14980 4018
rect 14934 3946 14940 4009
rect 14974 3946 14980 4009
rect 14934 3941 14980 3946
rect 14934 3874 14940 3941
rect 14974 3874 14980 3941
rect 14934 3873 14980 3874
rect 14934 3839 14940 3873
rect 14974 3839 14980 3873
rect 14934 3836 14980 3839
rect 14934 3771 14940 3836
rect 14974 3771 14980 3836
rect 14934 3764 14980 3771
rect 14934 3703 14940 3764
rect 14974 3703 14980 3764
rect 14934 3692 14980 3703
rect 14934 3635 14940 3692
rect 14974 3635 14980 3692
rect 14934 3620 14980 3635
rect 14934 3567 14940 3620
rect 14974 3567 14980 3620
rect 14934 3548 14980 3567
rect 14934 3499 14940 3548
rect 14974 3499 14980 3548
rect 14934 3476 14980 3499
rect 14934 3431 14940 3476
rect 14974 3431 14980 3476
rect 14934 3404 14980 3431
rect 14934 3363 14940 3404
rect 14974 3363 14980 3404
rect 14934 3332 14980 3363
rect 14934 3295 14940 3332
rect 14974 3295 14980 3332
rect 14934 3260 14980 3295
rect 14934 3226 14940 3260
rect 14974 3226 14980 3260
rect 14934 3205 14980 3226
rect 14934 3154 14940 3205
rect 14974 3154 14980 3205
rect 14934 3137 14980 3154
rect 14934 3082 14940 3137
rect 14974 3082 14980 3137
rect 14934 3069 14980 3082
rect 14934 3010 14940 3069
rect 14974 3010 14980 3069
rect 14934 3001 14980 3010
rect 14934 2938 14940 3001
rect 14974 2938 14980 3001
rect 14934 2933 14980 2938
rect 14934 2866 14940 2933
rect 14974 2866 14980 2933
rect 14934 2865 14980 2866
rect 14934 2831 14940 2865
rect 14974 2831 14980 2865
rect 14934 2828 14980 2831
rect 14934 2763 14940 2828
rect 14974 2763 14980 2828
rect 14934 2756 14980 2763
rect 14934 2695 14940 2756
rect 14974 2695 14980 2756
rect 14934 2684 14980 2695
rect 14934 2627 14940 2684
rect 14974 2627 14980 2684
rect 14934 2612 14980 2627
rect 14934 2559 14940 2612
rect 14974 2559 14980 2612
rect 14934 2540 14980 2559
rect 14934 2491 14940 2540
rect 14974 2491 14980 2540
rect 14934 2468 14980 2491
rect 14934 2423 14940 2468
rect 14974 2423 14980 2468
rect 14934 2396 14980 2423
rect 14934 2355 14940 2396
rect 14974 2355 14980 2396
rect 14934 2324 14980 2355
rect 14934 2287 14940 2324
rect 14974 2287 14980 2324
rect 14934 2253 14980 2287
rect 14934 2218 14940 2253
rect 14974 2218 14980 2253
rect 14934 2185 14980 2218
rect 14934 2146 14940 2185
rect 14974 2146 14980 2185
rect 14934 2117 14980 2146
rect 14934 2074 14940 2117
rect 14974 2074 14980 2117
rect 14934 2049 14980 2074
rect 14934 2002 14940 2049
rect 14974 2002 14980 2049
rect 14934 1981 14980 2002
rect 14934 1930 14940 1981
rect 14974 1930 14980 1981
rect 14934 1913 14980 1930
rect 14934 1858 14940 1913
rect 14974 1858 14980 1913
rect 14934 1845 14980 1858
rect 14934 1786 14940 1845
rect 14974 1786 14980 1845
rect 14934 1777 14980 1786
rect 14934 1714 14940 1777
rect 14974 1714 14980 1777
rect 14934 1709 14980 1714
rect 14934 1642 14940 1709
rect 14974 1642 14980 1709
rect 14934 1641 14980 1642
rect 14934 1607 14940 1641
rect 14974 1607 14980 1641
rect 14934 1604 14980 1607
rect 14934 1539 14940 1604
rect 14974 1539 14980 1604
rect 14934 1532 14980 1539
rect 14934 1471 14940 1532
rect 14974 1471 14980 1532
rect 14934 1460 14980 1471
rect 14934 1403 14940 1460
rect 14974 1403 14980 1460
rect 14934 1387 14980 1403
rect 14934 1335 14940 1387
rect 14974 1335 14980 1387
rect 14934 1314 14980 1335
rect 14934 1267 14940 1314
rect 14974 1267 14980 1314
rect 14934 1241 14980 1267
rect 14934 1199 14940 1241
rect 14974 1199 14980 1241
rect 14934 1168 14980 1199
rect 14934 1131 14940 1168
rect 14974 1131 14980 1168
rect 14934 1097 14980 1131
rect 14934 1061 14940 1097
rect 14974 1061 14980 1097
rect 14934 1029 14980 1061
rect 14934 988 14940 1029
rect 14974 988 14980 1029
rect 14934 961 14980 988
rect 14934 915 14940 961
rect 14974 915 14980 961
rect 14934 893 14980 915
rect 14934 842 14940 893
rect 14974 842 14980 893
rect 14934 825 14980 842
rect 14934 769 14940 825
rect 14974 769 14980 825
rect 14934 757 14980 769
rect 14934 696 14940 757
rect 14974 696 14980 757
rect 14934 689 14980 696
rect 14934 623 14940 689
rect 14974 623 14980 689
rect 14934 621 14980 623
rect 14934 587 14940 621
rect 14974 587 14980 621
rect 14934 584 14980 587
rect 14934 519 14940 584
rect 14974 519 14980 584
rect 14934 511 14980 519
rect 14934 451 14940 511
rect 14974 451 14980 511
rect 14934 438 14980 451
rect 13206 362 13252 380
rect 11644 291 11724 325
rect 11758 291 11774 325
rect 13206 312 13212 362
rect 13246 312 13252 362
rect 14798 383 14817 403
rect 14851 383 14864 403
rect 14798 345 14864 383
rect 14798 325 14817 345
rect 14680 324 14696 325
rect 14730 324 14814 325
rect 11418 220 11464 247
rect 11418 179 11424 220
rect 11458 179 11464 220
rect 11418 147 11464 179
rect 11418 111 11424 147
rect 11458 111 11464 147
rect 11418 80 11464 111
rect 13206 290 13252 312
rect 14682 291 14696 324
rect 14754 291 14814 324
rect 14851 311 14864 345
rect 14848 291 14864 311
rect 14934 383 14940 438
rect 14974 383 14980 438
rect 14934 365 14980 383
rect 14934 315 14940 365
rect 14974 315 14980 365
rect 14934 292 14980 315
rect 14682 290 14720 291
rect 13206 244 13212 290
rect 13246 244 13252 290
rect 13206 218 13252 244
rect 13206 176 13212 218
rect 13246 176 13252 218
rect 13206 146 13252 176
rect 13206 108 13212 146
rect 13246 108 13252 146
rect 13206 80 13252 108
rect 14934 247 14940 292
rect 14974 247 14980 292
rect 14934 219 14980 247
rect 14934 179 14940 219
rect 14974 179 14980 219
rect 14934 146 14980 179
rect 14934 111 14940 146
rect 14974 111 14980 146
rect 14934 80 14980 111
rect 11418 74 14980 80
rect 11418 40 11492 74
rect 11530 40 11560 74
rect 11604 40 11628 74
rect 11678 40 11696 74
rect 11752 40 11764 74
rect 11826 40 11832 74
rect 11934 40 11940 74
rect 12002 40 12014 74
rect 12070 40 12088 74
rect 12138 40 12162 74
rect 12206 40 12236 74
rect 12274 40 12308 74
rect 12344 40 12376 74
rect 12418 40 12444 74
rect 12492 40 12512 74
rect 12565 40 12580 74
rect 12638 40 12648 74
rect 12711 40 12716 74
rect 12818 40 12823 74
rect 12886 40 12896 74
rect 12954 40 12969 74
rect 13022 40 13042 74
rect 13090 40 13115 74
rect 13158 40 13188 74
rect 13222 40 13261 74
rect 13295 40 13308 74
rect 13368 40 13376 74
rect 13441 40 13444 74
rect 13478 40 13480 74
rect 13546 40 13553 74
rect 13614 40 13626 74
rect 13682 40 13699 74
rect 13750 40 13772 74
rect 13818 40 13845 74
rect 13886 40 13918 74
rect 13954 40 13988 74
rect 14025 40 14056 74
rect 14098 40 14124 74
rect 14171 40 14192 74
rect 14244 40 14260 74
rect 14317 40 14328 74
rect 14390 40 14396 74
rect 14463 40 14464 74
rect 14498 40 14502 74
rect 14566 40 14575 74
rect 14634 40 14648 74
rect 14702 40 14721 74
rect 14770 40 14794 74
rect 14838 40 14867 74
rect 14906 40 14980 74
rect 11418 34 14980 40
rect 11665 -189 11679 -155
rect 11733 -189 11751 -155
rect 11801 -189 11823 -155
rect 11869 -189 11896 -155
rect 11937 -189 11969 -155
rect 12005 -189 12039 -155
rect 12076 -189 12107 -155
rect 12149 -189 12175 -155
rect 12222 -189 12243 -155
rect 12295 -189 12311 -155
rect 12368 -189 12379 -155
rect 12441 -189 12447 -155
rect 12514 -189 12515 -155
rect 12549 -189 12553 -155
rect 12617 -189 12626 -155
rect 12685 -189 12699 -155
rect 12753 -189 12772 -155
rect 12821 -189 12845 -155
rect 12890 -189 12918 -155
rect 12959 -189 12991 -155
rect 13028 -189 13063 -155
rect 13098 -189 13132 -155
rect 13171 -189 13201 -155
rect 13244 -189 13270 -155
rect 13317 -189 13339 -155
rect 13390 -189 13408 -155
rect 13463 -189 13477 -155
rect 13536 -189 13546 -155
rect 13609 -189 13615 -155
rect 13682 -189 13684 -155
rect 13718 -189 13721 -155
rect 13787 -189 13794 -155
rect 13856 -189 13867 -155
rect 13925 -189 13940 -155
rect 13994 -189 14013 -155
rect 14063 -189 14086 -155
rect 14132 -189 14159 -155
rect 14201 -189 14232 -155
rect 14270 -189 14305 -155
rect 14339 -189 14374 -155
rect 14412 -189 14443 -155
rect 14485 -189 14512 -155
rect 14558 -189 14581 -155
rect 14631 -189 14650 -155
rect 14704 -189 14719 -155
rect 11771 -348 11805 -300
rect 11615 -473 11649 -432
rect 11615 -548 11649 -507
rect 11615 -623 11649 -582
rect 11615 -698 11649 -657
rect 11771 -430 11805 -382
rect 12083 -348 12117 -300
rect 11771 -512 11805 -464
rect 11771 -594 11805 -546
rect 11771 -677 11805 -628
rect 11927 -473 11961 -432
rect 11927 -548 11961 -507
rect 11927 -623 11961 -582
rect 11927 -698 11961 -657
rect 11615 -773 11649 -732
rect 12083 -430 12117 -382
rect 12395 -348 12429 -300
rect 12083 -512 12117 -464
rect 12083 -594 12117 -546
rect 12083 -677 12117 -628
rect 12239 -473 12273 -432
rect 12239 -548 12273 -507
rect 12239 -623 12273 -582
rect 12239 -698 12273 -657
rect 11927 -773 11961 -732
rect 12395 -430 12429 -382
rect 12707 -348 12741 -300
rect 12395 -512 12429 -464
rect 12395 -594 12429 -546
rect 12395 -677 12429 -628
rect 12551 -473 12585 -432
rect 12551 -548 12585 -507
rect 12551 -623 12585 -582
rect 12551 -698 12585 -657
rect 12239 -773 12273 -732
rect 12707 -430 12741 -382
rect 13018 -348 13052 -300
rect 12707 -512 12741 -464
rect 12707 -594 12741 -546
rect 12707 -677 12741 -628
rect 12863 -473 12897 -432
rect 12863 -548 12897 -507
rect 12863 -623 12897 -582
rect 12863 -698 12897 -657
rect 12551 -773 12585 -732
rect 13018 -430 13052 -382
rect 13331 -348 13365 -300
rect 13018 -512 13052 -464
rect 13018 -594 13052 -546
rect 13018 -677 13052 -628
rect 13175 -473 13209 -432
rect 13175 -548 13209 -507
rect 13175 -623 13209 -582
rect 13175 -698 13209 -657
rect 12863 -773 12897 -732
rect 13331 -430 13365 -382
rect 13643 -348 13677 -300
rect 13331 -512 13365 -464
rect 13331 -594 13365 -546
rect 13331 -677 13365 -628
rect 13487 -473 13521 -432
rect 13487 -548 13521 -507
rect 13487 -623 13521 -582
rect 13487 -698 13521 -657
rect 13175 -773 13209 -732
rect 13643 -430 13677 -382
rect 13955 -348 13989 -300
rect 13643 -512 13677 -464
rect 13643 -594 13677 -546
rect 13643 -677 13677 -628
rect 13799 -473 13833 -432
rect 13799 -548 13833 -507
rect 13799 -623 13833 -582
rect 13799 -698 13833 -657
rect 13487 -773 13521 -732
rect 13955 -430 13989 -382
rect 14267 -348 14301 -300
rect 13955 -512 13989 -464
rect 13955 -594 13989 -546
rect 13955 -677 13989 -628
rect 14111 -473 14145 -432
rect 14111 -548 14145 -507
rect 14111 -623 14145 -582
rect 14111 -698 14145 -657
rect 13799 -773 13833 -732
rect 14267 -430 14301 -382
rect 14579 -348 14613 -300
rect 14267 -512 14301 -464
rect 14267 -594 14301 -546
rect 14267 -677 14301 -628
rect 14423 -473 14457 -432
rect 14423 -548 14457 -507
rect 14423 -623 14457 -582
rect 14423 -698 14457 -657
rect 14111 -773 14145 -732
rect 14579 -430 14613 -382
rect 14579 -512 14613 -464
rect 14579 -594 14613 -546
rect 14579 -677 14613 -628
rect 14735 -444 14769 -396
rect 14735 -526 14769 -478
rect 14735 -608 14769 -560
rect 14735 -690 14769 -642
rect 14423 -773 14457 -732
rect 14735 -773 14769 -724
rect 11660 -951 11676 -917
rect 11724 -951 11744 -917
rect 11796 -951 11812 -917
rect 11868 -951 11880 -917
rect 11940 -951 11948 -917
rect 12012 -951 12016 -917
rect 12118 -951 12123 -917
rect 12186 -951 12196 -917
rect 12254 -951 12269 -917
rect 12322 -951 12342 -917
rect 12390 -951 12415 -917
rect 12458 -951 12488 -917
rect 12526 -951 12560 -917
rect 12595 -951 12628 -917
rect 12668 -951 12696 -917
rect 12741 -951 12764 -917
rect 12814 -951 12832 -917
rect 12887 -951 12900 -917
rect 12960 -951 12968 -917
rect 13033 -951 13036 -917
rect 13070 -951 13072 -917
rect 13138 -951 13145 -917
rect 13206 -951 13218 -917
rect 13274 -951 13291 -917
rect 13342 -951 13364 -917
rect 13410 -951 13437 -917
rect 13478 -951 13510 -917
rect 13546 -951 13580 -917
rect 13617 -951 13648 -917
rect 13690 -951 13716 -917
rect 13763 -951 13784 -917
rect 13836 -951 13852 -917
rect 13909 -951 13920 -917
rect 13982 -951 13988 -917
rect 14055 -951 14056 -917
rect 14090 -951 14094 -917
rect 14158 -951 14167 -917
rect 14226 -951 14240 -917
rect 14294 -951 14313 -917
rect 14363 -951 14386 -917
rect 14432 -951 14459 -917
rect 14501 -951 14532 -917
rect 14570 -951 14605 -917
rect 14639 -951 14674 -917
rect 14712 -951 14724 -917
<< viali >>
rect -176 38723 -142 38757
rect -99 38723 -74 38757
rect -74 38723 -65 38757
rect 11 38723 28 38757
rect 28 38723 45 38757
rect 83 38723 96 38757
rect 96 38723 117 38757
rect 155 38723 164 38757
rect 164 38723 189 38757
rect 227 38723 232 38757
rect 232 38723 261 38757
rect 299 38723 300 38757
rect 300 38723 333 38757
rect 371 38723 402 38757
rect 402 38723 405 38757
rect 443 38723 470 38757
rect 470 38723 477 38757
rect 515 38723 538 38757
rect 538 38723 549 38757
rect 587 38723 606 38757
rect 606 38723 621 38757
rect 659 38723 674 38757
rect 674 38723 693 38757
rect 731 38723 742 38757
rect 742 38723 765 38757
rect 803 38723 810 38757
rect 810 38723 837 38757
rect 875 38723 878 38757
rect 878 38723 909 38757
rect 947 38723 980 38757
rect 980 38723 981 38757
rect 1019 38723 1048 38757
rect 1048 38723 1053 38757
rect 1091 38723 1116 38757
rect 1116 38723 1125 38757
rect 1163 38723 1184 38757
rect 1184 38723 1197 38757
rect 1235 38723 1252 38757
rect 1252 38723 1269 38757
rect 1307 38723 1320 38757
rect 1320 38723 1341 38757
rect 1379 38723 1388 38757
rect 1388 38723 1413 38757
rect 1451 38723 1456 38757
rect 1456 38723 1485 38757
rect 1523 38723 1524 38757
rect 1524 38723 1557 38757
rect 1595 38723 1626 38757
rect 1626 38723 1629 38757
rect 1667 38723 1694 38757
rect 1694 38723 1701 38757
rect 1739 38723 1762 38757
rect 1762 38723 1773 38757
rect 1811 38723 1845 38757
rect 1883 38723 1898 38757
rect 1898 38723 1917 38757
rect 1955 38723 1966 38757
rect 1966 38723 1989 38757
rect 2027 38723 2034 38757
rect 2034 38723 2061 38757
rect 2100 38723 2102 38757
rect 2102 38723 2134 38757
rect 2173 38723 2204 38757
rect 2204 38723 2207 38757
rect 2246 38723 2272 38757
rect 2272 38723 2280 38757
rect 2319 38723 2340 38757
rect 2340 38723 2353 38757
rect 2392 38723 2408 38757
rect 2408 38723 2426 38757
rect 2465 38723 2476 38757
rect 2476 38723 2499 38757
rect 2538 38723 2544 38757
rect 2544 38723 2572 38757
rect 2611 38723 2612 38757
rect 2612 38723 2645 38757
rect 2684 38723 2714 38757
rect 2714 38723 2718 38757
rect 2757 38723 2782 38757
rect 2782 38723 2791 38757
rect 2830 38723 2850 38757
rect 2850 38723 2864 38757
rect 2903 38723 2918 38757
rect 2918 38723 2937 38757
rect 2976 38723 2986 38757
rect 2986 38723 3010 38757
rect 3049 38723 3054 38757
rect 3054 38723 3083 38757
rect 3122 38723 3156 38757
rect 3195 38723 3224 38757
rect 3224 38723 3229 38757
rect 3268 38723 3292 38757
rect 3292 38723 3302 38757
rect 3341 38723 3360 38757
rect 3360 38723 3375 38757
rect 3414 38723 3428 38757
rect 3428 38723 3448 38757
rect 3487 38723 3496 38757
rect 3496 38723 3521 38757
rect 3560 38723 3564 38757
rect 3564 38723 3594 38757
rect 3633 38723 3666 38757
rect 3666 38723 3667 38757
rect 3706 38723 3734 38757
rect 3734 38723 3740 38757
rect 3779 38723 3802 38757
rect 3802 38723 3813 38757
rect 3852 38723 3870 38757
rect 3870 38723 3886 38757
rect 3925 38723 3959 38757
rect 3998 38723 4032 38757
rect 4071 38723 4074 38757
rect 4074 38723 4105 38757
rect 4144 38723 4176 38757
rect 4176 38723 4178 38757
rect 4217 38723 4244 38757
rect 4244 38723 4251 38757
rect 4290 38723 4312 38757
rect 4312 38723 4324 38757
rect 4363 38723 4380 38757
rect 4380 38723 4397 38757
rect 4436 38723 4448 38757
rect 4448 38723 4470 38757
rect 4509 38723 4516 38757
rect 4516 38723 4543 38757
rect 4582 38723 4584 38757
rect 4584 38723 4616 38757
rect 4655 38723 4686 38757
rect 4686 38723 4689 38757
rect 4728 38723 4754 38757
rect 4754 38723 4762 38757
rect 4801 38723 4822 38757
rect 4822 38723 4835 38757
rect 4874 38723 4890 38757
rect 4890 38723 4908 38757
rect 4947 38723 4958 38757
rect 4958 38723 4981 38757
rect 5020 38723 5026 38757
rect 5026 38723 5054 38757
rect 5093 38723 5094 38757
rect 5094 38723 5127 38757
rect 5166 38723 5196 38757
rect 5196 38723 5200 38757
rect 5239 38723 5264 38757
rect 5264 38723 5273 38757
rect 5312 38723 5332 38757
rect 5332 38723 5346 38757
rect 5385 38723 5400 38757
rect 5400 38723 5419 38757
rect 5458 38723 5468 38757
rect 5468 38723 5492 38757
rect 5531 38723 5536 38757
rect 5536 38723 5565 38757
rect 5604 38723 5638 38757
rect 5677 38723 5706 38757
rect 5706 38723 5711 38757
rect 5750 38723 5774 38757
rect 5774 38723 5784 38757
rect 5823 38723 5842 38757
rect 5842 38723 5857 38757
rect 5896 38723 5910 38757
rect 5910 38723 5930 38757
rect 5969 38723 5978 38757
rect 5978 38723 6003 38757
rect 6042 38723 6046 38757
rect 6046 38723 6076 38757
rect -252 38655 -218 38685
rect -252 38651 -218 38655
rect -252 38587 -218 38612
rect -252 38578 -218 38587
rect -252 38519 -218 38539
rect -252 38505 -218 38519
rect -252 38451 -218 38466
rect -252 38432 -218 38451
rect -252 38383 -218 38393
rect -252 38359 -218 38383
rect -252 38315 -218 38320
rect -252 38286 -218 38315
rect -252 38213 -218 38247
rect -252 38145 -218 38174
rect -252 38140 -218 38145
rect -252 38077 -218 38101
rect -252 38067 -218 38077
rect -252 38009 -218 38028
rect -252 37994 -218 38009
rect -252 37941 -218 37955
rect -252 37921 -218 37941
rect -252 37873 -218 37882
rect -252 37848 -218 37873
rect -252 37805 -218 37809
rect -252 37775 -218 37805
rect -252 37703 -218 37736
rect -252 37702 -218 37703
rect -252 37635 -218 37663
rect -252 37629 -218 37635
rect -252 37567 -218 37590
rect -252 37556 -218 37567
rect -252 37499 -218 37517
rect -252 37483 -218 37499
rect -252 37431 -218 37444
rect -252 37410 -218 37431
rect -252 37363 -218 37371
rect -252 37337 -218 37363
rect -252 37295 -218 37298
rect -252 37264 -218 37295
rect -252 37193 -218 37225
rect -252 37191 -218 37193
rect -252 37125 -218 37152
rect -252 37118 -218 37125
rect -252 37057 -218 37079
rect -252 37045 -218 37057
rect -252 36989 -218 37006
rect -252 36972 -218 36989
rect -252 36921 -218 36933
rect -252 36899 -218 36921
rect -252 36853 -218 36860
rect -252 36826 -218 36853
rect -252 36785 -218 36787
rect -252 36753 -218 36785
rect -252 36683 -218 36714
rect -252 36680 -218 36683
rect -252 36615 -218 36641
rect -252 36607 -218 36615
rect -252 36547 -218 36568
rect -252 36534 -218 36547
rect -252 36479 -218 36495
rect -252 36461 -218 36479
rect -252 36411 -218 36422
rect -252 36388 -218 36411
rect -252 36343 -218 36349
rect -252 36315 -218 36343
rect -252 36275 -218 36276
rect -252 36242 -218 36275
rect -252 36173 -218 36203
rect -252 36169 -218 36173
rect -252 36105 -218 36130
rect -252 36096 -218 36105
rect -252 36037 -218 36057
rect -252 36023 -218 36037
rect -252 35969 -218 35984
rect -252 35950 -218 35969
rect -252 35901 -218 35911
rect -252 35877 -218 35901
rect -252 35833 -218 35838
rect -252 35804 -218 35833
rect -252 35731 -218 35765
rect -252 35663 -218 35692
rect -252 35658 -218 35663
rect -252 35595 -218 35619
rect -252 35585 -218 35595
rect -252 35527 -218 35546
rect -252 35512 -218 35527
rect -252 35459 -218 35473
rect -252 35439 -218 35459
rect -252 35391 -218 35400
rect -252 35366 -218 35391
rect -252 35323 -218 35327
rect -252 35293 -218 35323
rect -252 35221 -218 35254
rect -252 35220 -218 35221
rect -252 35153 -218 35181
rect -252 35147 -218 35153
rect -252 35085 -218 35109
rect -252 35075 -218 35085
rect -252 35017 -218 35037
rect -252 35003 -218 35017
rect -252 34949 -218 34965
rect -252 34931 -218 34949
rect -252 34881 -218 34893
rect -252 34859 -218 34881
rect -252 34813 -218 34821
rect -252 34787 -218 34813
rect -252 34745 -218 34749
rect -252 34715 -218 34745
rect -252 34643 -218 34677
rect -252 34575 -218 34605
rect -252 34571 -218 34575
rect -252 34507 -218 34533
rect -252 34499 -218 34507
rect -252 34439 -218 34461
rect -252 34427 -218 34439
rect -252 34371 -218 34389
rect -252 34355 -218 34371
rect -252 34303 -218 34317
rect -252 34283 -218 34303
rect -252 34235 -218 34245
rect -252 34211 -218 34235
rect -252 34167 -218 34173
rect -252 34139 -218 34167
rect -252 34099 -218 34101
rect -252 34067 -218 34099
rect -252 33997 -218 34029
rect -252 33995 -218 33997
rect -252 33929 -218 33957
rect -252 33923 -218 33929
rect -252 33861 -218 33885
rect -252 33851 -218 33861
rect -252 33793 -218 33813
rect -252 33779 -218 33793
rect -252 33725 -218 33741
rect -252 33707 -218 33725
rect -252 33657 -218 33669
rect -252 33635 -218 33657
rect -252 33589 -218 33597
rect -252 33563 -218 33589
rect -252 33521 -218 33525
rect -252 33491 -218 33521
rect -252 33419 -218 33453
rect -252 33351 -218 33381
rect -252 33347 -218 33351
rect -252 33283 -218 33309
rect -252 33275 -218 33283
rect -252 33215 -218 33237
rect -252 33203 -218 33215
rect -252 33147 -218 33165
rect -252 33131 -218 33147
rect -252 33079 -218 33093
rect -252 33059 -218 33079
rect -252 33011 -218 33021
rect -252 32987 -218 33011
rect -252 32943 -218 32949
rect -252 32915 -218 32943
rect -252 32875 -218 32877
rect -252 32843 -218 32875
rect -252 32773 -218 32805
rect -252 32771 -218 32773
rect -252 32705 -218 32733
rect -252 32699 -218 32705
rect -252 32637 -218 32661
rect -252 32627 -218 32637
rect -252 32569 -218 32589
rect -252 32555 -218 32569
rect -252 32501 -218 32517
rect -252 32483 -218 32501
rect -252 32433 -218 32445
rect -252 32411 -218 32433
rect -252 32365 -218 32373
rect -252 32339 -218 32365
rect -252 32297 -218 32301
rect -252 32267 -218 32297
rect -252 32195 -218 32229
rect -252 32127 -218 32157
rect -252 32123 -218 32127
rect -252 32059 -218 32085
rect -252 32051 -218 32059
rect -252 31991 -218 32013
rect -252 31979 -218 31991
rect -252 31923 -218 31941
rect -252 31907 -218 31923
rect -252 31855 -218 31869
rect -252 31835 -218 31855
rect -252 31787 -218 31797
rect -252 31763 -218 31787
rect -252 31719 -218 31725
rect -252 31691 -218 31719
rect -252 31651 -218 31653
rect -252 31619 -218 31651
rect -252 31549 -218 31581
rect -252 31547 -218 31549
rect -252 31481 -218 31509
rect -252 31475 -218 31481
rect -252 31413 -218 31437
rect -252 31403 -218 31413
rect -252 31345 -218 31365
rect -252 31331 -218 31345
rect -252 31277 -218 31293
rect -252 31259 -218 31277
rect -252 31209 -218 31221
rect -252 31187 -218 31209
rect -252 31141 -218 31149
rect -252 31115 -218 31141
rect -252 31073 -218 31077
rect -252 31043 -218 31073
rect -252 30971 -218 31005
rect -252 30903 -218 30933
rect -252 30899 -218 30903
rect -252 30835 -218 30861
rect -252 30827 -218 30835
rect -252 30767 -218 30789
rect -252 30755 -218 30767
rect -252 30699 -218 30717
rect -252 30683 -218 30699
rect -252 30631 -218 30645
rect -252 30611 -218 30631
rect -252 30563 -218 30573
rect -252 30539 -218 30563
rect -252 30495 -218 30501
rect -252 30467 -218 30495
rect -252 30427 -218 30429
rect -252 30395 -218 30427
rect -252 30325 -218 30357
rect -252 30323 -218 30325
rect -252 30257 -218 30285
rect -252 30251 -218 30257
rect -252 30189 -218 30213
rect -252 30179 -218 30189
rect -252 30121 -218 30141
rect -252 30107 -218 30121
rect -252 30053 -218 30069
rect -252 30035 -218 30053
rect -252 29985 -218 29997
rect -252 29963 -218 29985
rect -252 29917 -218 29925
rect -252 29891 -218 29917
rect -252 29849 -218 29853
rect -252 29819 -218 29849
rect -252 29747 -218 29781
rect -252 29679 -218 29709
rect -252 29675 -218 29679
rect -252 29611 -218 29637
rect -252 29603 -218 29611
rect -252 29543 -218 29565
rect -252 29531 -218 29543
rect -252 29475 -218 29493
rect -252 29459 -218 29475
rect -252 29407 -218 29421
rect -252 29387 -218 29407
rect -252 29339 -218 29349
rect -252 29315 -218 29339
rect -252 29271 -218 29277
rect -252 29243 -218 29271
rect -252 29203 -218 29205
rect -252 29171 -218 29203
rect -252 29101 -218 29133
rect -252 29099 -218 29101
rect -252 29033 -218 29061
rect -252 29027 -218 29033
rect -252 28965 -218 28989
rect -252 28955 -218 28965
rect -252 28897 -218 28917
rect -252 28883 -218 28897
rect -252 28829 -218 28845
rect -252 28811 -218 28829
rect -252 28761 -218 28773
rect -252 28739 -218 28761
rect -252 28693 -218 28701
rect -252 28667 -218 28693
rect -252 28625 -218 28629
rect -252 28595 -218 28625
rect -252 28523 -218 28557
rect -252 28455 -218 28485
rect -252 28451 -218 28455
rect -252 28387 -218 28413
rect -252 28379 -218 28387
rect -252 28319 -218 28341
rect -252 28307 -218 28319
rect -252 28251 -218 28269
rect -252 28235 -218 28251
rect -252 28183 -218 28197
rect -252 28163 -218 28183
rect -252 28115 -218 28125
rect -252 28091 -218 28115
rect -252 28047 -218 28053
rect -252 28019 -218 28047
rect -252 27979 -218 27981
rect -252 27947 -218 27979
rect -252 27877 -218 27909
rect -252 27875 -218 27877
rect -252 27809 -218 27837
rect -252 27803 -218 27809
rect -252 27741 -218 27765
rect -252 27731 -218 27741
rect -252 27673 -218 27693
rect -252 27659 -218 27673
rect -252 27605 -218 27621
rect -252 27587 -218 27605
rect -252 27537 -218 27549
rect -252 27515 -218 27537
rect -252 27469 -218 27477
rect -252 27443 -218 27469
rect -252 27401 -218 27405
rect -252 27371 -218 27401
rect -252 27299 -218 27333
rect -252 27231 -218 27261
rect -252 27227 -218 27231
rect -252 27163 -218 27189
rect -252 27155 -218 27163
rect -252 27095 -218 27117
rect -252 27083 -218 27095
rect -252 27027 -218 27045
rect -252 27011 -218 27027
rect -252 26959 -218 26973
rect -252 26939 -218 26959
rect -252 26891 -218 26901
rect -252 26867 -218 26891
rect -252 26823 -218 26829
rect -252 26795 -218 26823
rect -252 26755 -218 26757
rect -252 26723 -218 26755
rect -252 26653 -218 26685
rect -252 26651 -218 26653
rect -252 26585 -218 26613
rect -252 26579 -218 26585
rect -252 26517 -218 26541
rect -252 26507 -218 26517
rect -252 26449 -218 26469
rect -252 26435 -218 26449
rect -252 26381 -218 26397
rect -252 26363 -218 26381
rect -252 26313 -218 26325
rect -252 26291 -218 26313
rect -252 26245 -218 26253
rect -252 26219 -218 26245
rect -252 26177 -218 26181
rect -252 26147 -218 26177
rect -252 26075 -218 26109
rect -252 26007 -218 26037
rect -252 26003 -218 26007
rect -252 25939 -218 25965
rect -252 25931 -218 25939
rect -252 25871 -218 25893
rect -252 25859 -218 25871
rect -252 25803 -218 25821
rect -252 25787 -218 25803
rect -252 25735 -218 25749
rect -252 25715 -218 25735
rect -252 25667 -218 25677
rect -252 25643 -218 25667
rect -252 25599 -218 25605
rect -252 25571 -218 25599
rect -252 25531 -218 25533
rect -252 25499 -218 25531
rect -252 25429 -218 25461
rect -252 25427 -218 25429
rect -252 25361 -218 25389
rect -252 25355 -218 25361
rect -252 25293 -218 25317
rect -252 25283 -218 25293
rect -252 25225 -218 25245
rect -252 25211 -218 25225
rect -252 25157 -218 25173
rect -252 25139 -218 25157
rect -252 25089 -218 25101
rect -252 25067 -218 25089
rect -252 25021 -218 25029
rect -252 24995 -218 25021
rect -252 24953 -218 24957
rect -252 24923 -218 24953
rect -252 24851 -218 24885
rect -252 24783 -218 24813
rect -252 24779 -218 24783
rect -252 24715 -218 24741
rect -252 24707 -218 24715
rect -252 24647 -218 24669
rect -252 24635 -218 24647
rect -252 24579 -218 24597
rect -252 24563 -218 24579
rect -252 24511 -218 24525
rect -252 24491 -218 24511
rect -252 24443 -218 24453
rect -252 24419 -218 24443
rect -252 24375 -218 24381
rect -252 24347 -218 24375
rect -252 24307 -218 24309
rect -252 24275 -218 24307
rect -252 24205 -218 24237
rect -252 24203 -218 24205
rect -252 24137 -218 24165
rect -252 24131 -218 24137
rect -252 24069 -218 24093
rect -252 24059 -218 24069
rect -252 24001 -218 24021
rect -252 23987 -218 24001
rect -252 23933 -218 23949
rect -252 23915 -218 23933
rect -252 23865 -218 23877
rect -252 23843 -218 23865
rect -252 23797 -218 23805
rect -252 23771 -218 23797
rect -252 23729 -218 23733
rect -252 23699 -218 23729
rect -252 23627 -218 23661
rect -252 23559 -218 23589
rect -252 23555 -218 23559
rect -252 23491 -218 23517
rect -252 23483 -218 23491
rect -252 23423 -218 23445
rect -252 23411 -218 23423
rect -252 23355 -218 23373
rect -252 23339 -218 23355
rect -252 23287 -218 23301
rect -252 23267 -218 23287
rect -252 23219 -218 23229
rect -252 23195 -218 23219
rect -252 23151 -218 23157
rect -252 23123 -218 23151
rect -252 23083 -218 23085
rect -252 23051 -218 23083
rect -252 22981 -218 23013
rect -252 22979 -218 22981
rect -252 22913 -218 22941
rect -252 22907 -218 22913
rect -252 22845 -218 22869
rect -252 22835 -218 22845
rect -252 22777 -218 22797
rect -252 22763 -218 22777
rect -252 22709 -218 22725
rect -252 22691 -218 22709
rect -252 22641 -218 22653
rect -252 22619 -218 22641
rect -252 22573 -218 22581
rect -252 22547 -218 22573
rect -252 22505 -218 22509
rect -252 22475 -218 22505
rect -252 22403 -218 22437
rect -252 22335 -218 22365
rect -252 22331 -218 22335
rect -252 22267 -218 22293
rect -252 22259 -218 22267
rect -252 22199 -218 22221
rect -252 22187 -218 22199
rect -252 22131 -218 22149
rect -252 22115 -218 22131
rect -252 22063 -218 22077
rect -252 22043 -218 22063
rect -252 21995 -218 22005
rect -252 21971 -218 21995
rect -252 21927 -218 21933
rect -252 21899 -218 21927
rect -252 21859 -218 21861
rect -252 21827 -218 21859
rect -252 21757 -218 21789
rect -252 21755 -218 21757
rect -252 21689 -218 21717
rect -252 21683 -218 21689
rect -252 21621 -218 21645
rect -252 21611 -218 21621
rect -252 21553 -218 21573
rect -252 21539 -218 21553
rect -252 21485 -218 21501
rect -252 21467 -218 21485
rect -252 21417 -218 21429
rect -252 21395 -218 21417
rect -252 21349 -218 21357
rect -252 21323 -218 21349
rect -252 21281 -218 21285
rect -252 21251 -218 21281
rect -252 21179 -218 21213
rect -252 21111 -218 21141
rect -252 21107 -218 21111
rect -252 21043 -218 21069
rect -252 21035 -218 21043
rect -252 20975 -218 20997
rect -252 20963 -218 20975
rect -252 20907 -218 20925
rect -252 20891 -218 20907
rect -252 20839 -218 20853
rect -252 20819 -218 20839
rect -252 20771 -218 20781
rect -252 20747 -218 20771
rect -252 20703 -218 20709
rect -252 20675 -218 20703
rect -252 20635 -218 20637
rect -252 20603 -218 20635
rect -252 20533 -218 20565
rect -252 20531 -218 20533
rect -252 20465 -218 20493
rect -252 20459 -218 20465
rect -252 20397 -218 20421
rect -252 20387 -218 20397
rect -252 20329 -218 20349
rect -252 20315 -218 20329
rect -252 20261 -218 20277
rect -252 20243 -218 20261
rect -252 20193 -218 20205
rect -252 20171 -218 20193
rect -252 20125 -218 20133
rect -252 20099 -218 20125
rect -252 20057 -218 20061
rect -252 20027 -218 20057
rect -252 19955 -218 19989
rect -252 19887 -218 19917
rect -252 19883 -218 19887
rect -252 19819 -218 19845
rect -252 19811 -218 19819
rect -252 19751 -218 19773
rect -252 19739 -218 19751
rect -252 19683 -218 19701
rect -252 19667 -218 19683
rect -252 19615 -218 19629
rect -252 19595 -218 19615
rect -252 19547 -218 19557
rect -252 19523 -218 19547
rect -252 19479 -218 19485
rect -252 19451 -218 19479
rect -252 19411 -218 19413
rect -252 19379 -218 19411
rect -252 19309 -218 19341
rect -252 19307 -218 19309
rect -252 19241 -218 19269
rect -252 19235 -218 19241
rect -252 19173 -218 19197
rect -252 19163 -218 19173
rect -252 19105 -218 19125
rect -252 19091 -218 19105
rect -252 19037 -218 19053
rect -252 19019 -218 19037
rect -252 18969 -218 18981
rect -252 18947 -218 18969
rect -252 18901 -218 18909
rect -252 18875 -218 18901
rect -252 18833 -218 18837
rect -252 18803 -218 18833
rect -252 18731 -218 18765
rect -252 18663 -218 18693
rect -252 18659 -218 18663
rect -252 18595 -218 18621
rect -252 18587 -218 18595
rect -252 18527 -218 18549
rect -252 18515 -218 18527
rect -252 18459 -218 18477
rect -252 18443 -218 18459
rect -252 18391 -218 18405
rect -252 18371 -218 18391
rect -252 18323 -218 18333
rect -252 18299 -218 18323
rect -252 18255 -218 18261
rect -252 18227 -218 18255
rect -252 18187 -218 18189
rect -252 18155 -218 18187
rect -252 18085 -218 18117
rect -252 18083 -218 18085
rect -252 18017 -218 18045
rect -252 18011 -218 18017
rect -252 17949 -218 17973
rect -252 17939 -218 17949
rect -252 17881 -218 17901
rect -252 17867 -218 17881
rect -252 17813 -218 17829
rect -252 17795 -218 17813
rect -252 17745 -218 17757
rect -252 17723 -218 17745
rect -252 17677 -218 17685
rect -252 17651 -218 17677
rect -252 17609 -218 17613
rect -252 17579 -218 17609
rect -252 17507 -218 17541
rect -252 17439 -218 17469
rect -252 17435 -218 17439
rect -252 17371 -218 17397
rect -252 17363 -218 17371
rect -252 17303 -218 17325
rect -252 17291 -218 17303
rect -252 17235 -218 17253
rect -252 17219 -218 17235
rect -252 17167 -218 17181
rect -252 17147 -218 17167
rect -252 17099 -218 17109
rect -252 17075 -218 17099
rect -252 17031 -218 17037
rect -252 17003 -218 17031
rect -252 16963 -218 16965
rect -252 16931 -218 16963
rect -252 16861 -218 16893
rect -252 16859 -218 16861
rect -252 16793 -218 16821
rect -252 16787 -218 16793
rect -252 16725 -218 16749
rect -252 16715 -218 16725
rect -252 16657 -218 16677
rect -252 16643 -218 16657
rect -252 16589 -218 16605
rect -252 16571 -218 16589
rect -252 16521 -218 16533
rect -252 16499 -218 16521
rect -252 16453 -218 16461
rect -252 16427 -218 16453
rect -252 16385 -218 16389
rect -252 16355 -218 16385
rect -252 16283 -218 16317
rect -252 16215 -218 16245
rect -252 16211 -218 16215
rect -252 16147 -218 16173
rect -252 16139 -218 16147
rect -252 16079 -218 16101
rect -252 16067 -218 16079
rect -252 16011 -218 16029
rect -252 15995 -218 16011
rect -252 15943 -218 15957
rect -252 15923 -218 15943
rect -252 15875 -218 15885
rect -252 15851 -218 15875
rect -252 15807 -218 15813
rect -252 15779 -218 15807
rect -252 15739 -218 15741
rect -252 15707 -218 15739
rect -252 15637 -218 15669
rect -252 15635 -218 15637
rect -252 15569 -218 15597
rect -252 15563 -218 15569
rect -252 15501 -218 15525
rect -252 15491 -218 15501
rect -252 15433 -218 15453
rect -252 15419 -218 15433
rect -252 15365 -218 15381
rect -252 15347 -218 15365
rect -252 15297 -218 15309
rect -252 15275 -218 15297
rect -252 15229 -218 15237
rect -252 15203 -218 15229
rect -252 15161 -218 15165
rect -252 15131 -218 15161
rect -252 15059 -218 15093
rect -252 14991 -218 15021
rect -252 14987 -218 14991
rect -252 14923 -218 14949
rect -252 14915 -218 14923
rect -252 14855 -218 14877
rect -252 14843 -218 14855
rect -252 14787 -218 14805
rect -252 14771 -218 14787
rect -252 14719 -218 14733
rect -252 14699 -218 14719
rect -252 14651 -218 14661
rect -252 14627 -218 14651
rect -252 14583 -218 14589
rect -252 14555 -218 14583
rect -252 14515 -218 14517
rect -252 14483 -218 14515
rect -252 14413 -218 14445
rect -252 14411 -218 14413
rect -252 14345 -218 14373
rect -252 14339 -218 14345
rect -252 14277 -218 14301
rect -252 14267 -218 14277
rect -252 14209 -218 14229
rect -252 14195 -218 14209
rect -252 14141 -218 14157
rect -252 14123 -218 14141
rect -252 14073 -218 14085
rect -252 14051 -218 14073
rect -252 14005 -218 14013
rect -252 13979 -218 14005
rect -252 13937 -218 13941
rect -252 13907 -218 13937
rect -252 13835 -218 13869
rect -252 13767 -218 13797
rect -252 13763 -218 13767
rect -252 13699 -218 13725
rect -252 13691 -218 13699
rect -252 13631 -218 13653
rect -252 13619 -218 13631
rect -252 13563 -218 13581
rect -252 13547 -218 13563
rect -252 13495 -218 13509
rect -252 13475 -218 13495
rect -252 13427 -218 13437
rect -252 13403 -218 13427
rect -252 13359 -218 13365
rect -252 13331 -218 13359
rect -252 13291 -218 13293
rect -252 13259 -218 13291
rect -252 13189 -218 13221
rect -252 13187 -218 13189
rect -252 13121 -218 13149
rect -252 13115 -218 13121
rect -252 13053 -218 13077
rect -252 13043 -218 13053
rect -252 12985 -218 13005
rect -252 12971 -218 12985
rect -252 12917 -218 12933
rect -252 12899 -218 12917
rect -252 12849 -218 12861
rect -252 12827 -218 12849
rect -252 12781 -218 12789
rect -252 12755 -218 12781
rect -252 12713 -218 12717
rect -252 12683 -218 12713
rect -252 12611 -218 12645
rect -252 12543 -218 12573
rect -252 12539 -218 12543
rect -252 12475 -218 12501
rect -252 12467 -218 12475
rect -252 12407 -218 12429
rect -252 12395 -218 12407
rect -252 12339 -218 12357
rect -252 12323 -218 12339
rect -252 12271 -218 12285
rect -252 12251 -218 12271
rect -252 12203 -218 12213
rect -252 12179 -218 12203
rect -252 12135 -218 12141
rect -252 12107 -218 12135
rect -252 12067 -218 12069
rect -252 12035 -218 12067
rect -252 11965 -218 11997
rect -252 11963 -218 11965
rect -252 11897 -218 11925
rect -252 11891 -218 11897
rect -252 11829 -218 11853
rect -252 11819 -218 11829
rect -252 11761 -218 11781
rect -252 11747 -218 11761
rect -252 11693 -218 11709
rect -252 11675 -218 11693
rect -252 11625 -218 11637
rect -252 11603 -218 11625
rect -252 11557 -218 11565
rect -252 11531 -218 11557
rect -252 11489 -218 11493
rect -252 11459 -218 11489
rect -252 11387 -218 11421
rect -252 11319 -218 11349
rect -252 11315 -218 11319
rect -252 11251 -218 11277
rect -252 11243 -218 11251
rect -252 11183 -218 11205
rect -252 11171 -218 11183
rect -252 11115 -218 11133
rect -252 11099 -218 11115
rect -252 11047 -218 11061
rect -252 11027 -218 11047
rect -252 10979 -218 10989
rect -252 10955 -218 10979
rect -252 10911 -218 10917
rect -252 10883 -218 10911
rect -252 10843 -218 10845
rect -252 10811 -218 10843
rect -252 10741 -218 10773
rect -252 10739 -218 10741
rect -252 10673 -218 10701
rect -252 10667 -218 10673
rect -252 10605 -218 10629
rect -252 10595 -218 10605
rect -252 10537 -218 10557
rect -252 10523 -218 10537
rect -252 10469 -218 10485
rect -252 10451 -218 10469
rect -252 10401 -218 10413
rect -252 10379 -218 10401
rect -252 10333 -218 10341
rect -252 10307 -218 10333
rect -252 10265 -218 10269
rect -252 10235 -218 10265
rect -252 10163 -218 10197
rect -252 10095 -218 10125
rect -252 10091 -218 10095
rect -252 10027 -218 10053
rect -252 10019 -218 10027
rect -252 9959 -218 9981
rect -252 9947 -218 9959
rect -252 9891 -218 9909
rect -252 9875 -218 9891
rect -252 9823 -218 9837
rect -252 9803 -218 9823
rect -252 9755 -218 9765
rect -252 9731 -218 9755
rect -252 9687 -218 9693
rect -252 9659 -218 9687
rect -252 9619 -218 9621
rect -252 9587 -218 9619
rect -252 9517 -218 9549
rect -252 9515 -218 9517
rect -252 9449 -218 9477
rect -252 9443 -218 9449
rect -252 9381 -218 9405
rect -252 9371 -218 9381
rect -252 9313 -218 9333
rect -252 9299 -218 9313
rect -252 9245 -218 9261
rect -252 9227 -218 9245
rect -252 9177 -218 9189
rect -252 9155 -218 9177
rect -252 9109 -218 9117
rect -252 9083 -218 9109
rect -252 9041 -218 9045
rect -252 9011 -218 9041
rect -252 8939 -218 8973
rect -252 8871 -218 8901
rect -252 8867 -218 8871
rect -252 8803 -218 8829
rect -252 8795 -218 8803
rect -252 8735 -218 8757
rect -252 8723 -218 8735
rect -252 8667 -218 8685
rect -252 8651 -218 8667
rect -252 8599 -218 8613
rect -252 8579 -218 8599
rect -252 8531 -218 8541
rect -252 8507 -218 8531
rect -252 8463 -218 8469
rect -252 8435 -218 8463
rect -252 8395 -218 8397
rect -252 8363 -218 8395
rect -252 8293 -218 8325
rect -252 8291 -218 8293
rect -252 8225 -218 8253
rect -252 8219 -218 8225
rect -252 8157 -218 8181
rect -252 8147 -218 8157
rect -252 8089 -218 8109
rect -252 8075 -218 8089
rect -252 8021 -218 8037
rect -252 8003 -218 8021
rect -252 7953 -218 7965
rect -252 7931 -218 7953
rect -252 7885 -218 7893
rect -252 7859 -218 7885
rect -252 7817 -218 7821
rect -252 7787 -218 7817
rect -252 7715 -218 7749
rect -252 7647 -218 7677
rect -252 7643 -218 7647
rect -252 7579 -218 7605
rect -252 7571 -218 7579
rect -252 7511 -218 7533
rect -252 7499 -218 7511
rect -252 7443 -218 7461
rect -252 7427 -218 7443
rect -252 7375 -218 7389
rect -252 7355 -218 7375
rect -252 7307 -218 7317
rect -252 7283 -218 7307
rect -252 7239 -218 7245
rect -252 7211 -218 7239
rect -252 7171 -218 7173
rect -252 7139 -218 7171
rect -252 7069 -218 7101
rect -252 7067 -218 7069
rect -252 7001 -218 7029
rect -252 6995 -218 7001
rect -252 6933 -218 6957
rect -252 6923 -218 6933
rect -252 6865 -218 6885
rect -252 6851 -218 6865
rect -252 6797 -218 6813
rect -252 6779 -218 6797
rect -252 6729 -218 6741
rect -252 6707 -218 6729
rect -252 6661 -218 6669
rect -252 6635 -218 6661
rect -252 6593 -218 6597
rect -252 6563 -218 6593
rect -252 6491 -218 6525
rect -252 6423 -218 6453
rect -252 6419 -218 6423
rect -252 6355 -218 6381
rect -252 6347 -218 6355
rect -252 6287 -218 6309
rect -252 6275 -218 6287
rect -252 6219 -218 6237
rect -252 6203 -218 6219
rect -252 6151 -218 6165
rect -252 6131 -218 6151
rect -252 6083 -218 6093
rect -252 6059 -218 6083
rect -252 6015 -218 6021
rect -252 5987 -218 6015
rect -252 5947 -218 5949
rect -252 5915 -218 5947
rect -252 5845 -218 5877
rect -252 5843 -218 5845
rect -252 5777 -218 5805
rect -252 5771 -218 5777
rect -252 5709 -218 5733
rect -252 5699 -218 5709
rect -252 5641 -218 5661
rect -252 5627 -218 5641
rect -252 5573 -218 5589
rect -252 5555 -218 5573
rect -252 5505 -218 5517
rect -252 5483 -218 5505
rect -252 5437 -218 5445
rect -252 5411 -218 5437
rect -252 5369 -218 5373
rect -252 5339 -218 5369
rect -252 5267 -218 5301
rect -252 5199 -218 5229
rect -252 5195 -218 5199
rect -252 5131 -218 5157
rect -252 5123 -218 5131
rect -252 5063 -218 5085
rect -252 5051 -218 5063
rect -252 4995 -218 5013
rect -252 4979 -218 4995
rect -252 4927 -218 4941
rect -252 4907 -218 4927
rect -252 4859 -218 4869
rect -252 4835 -218 4859
rect -252 4791 -218 4797
rect -252 4763 -218 4791
rect -252 4723 -218 4725
rect -252 4691 -218 4723
rect -252 4621 -218 4653
rect -252 4619 -218 4621
rect -252 4553 -218 4581
rect -252 4547 -218 4553
rect -252 4485 -218 4509
rect -252 4475 -218 4485
rect -252 4417 -218 4437
rect -252 4403 -218 4417
rect -252 4349 -218 4365
rect -252 4331 -218 4349
rect -252 4281 -218 4293
rect -252 4259 -218 4281
rect -252 4213 -218 4221
rect -252 4187 -218 4213
rect -252 4145 -218 4149
rect -252 4115 -218 4145
rect -252 4043 -218 4077
rect -252 3975 -218 4005
rect -252 3971 -218 3975
rect -252 3907 -218 3933
rect -252 3899 -218 3907
rect -252 3839 -218 3861
rect -252 3827 -218 3839
rect -252 3771 -218 3789
rect -252 3755 -218 3771
rect -252 3703 -218 3717
rect -252 3683 -218 3703
rect -252 3635 -218 3645
rect -252 3611 -218 3635
rect -252 3567 -218 3573
rect -252 3539 -218 3567
rect -252 3499 -218 3501
rect -252 3467 -218 3499
rect 1830 38651 1864 38685
rect 1830 38607 1864 38612
rect 1830 38578 1864 38607
rect 1830 38505 1864 38539
rect 1830 38437 1864 38466
rect 1830 38432 1864 38437
rect 1830 38369 1864 38393
rect 1830 38359 1864 38369
rect 1830 38301 1864 38320
rect 1830 38286 1864 38301
rect 1830 38233 1864 38247
rect 1830 38213 1864 38233
rect 1830 38165 1864 38174
rect 1830 38140 1864 38165
rect 1830 38097 1864 38101
rect 1830 38067 1864 38097
rect 1830 37995 1864 38028
rect 1830 37994 1864 37995
rect 1830 37927 1864 37955
rect 1830 37921 1864 37927
rect 1830 37859 1864 37882
rect 1830 37848 1864 37859
rect 1830 37791 1864 37809
rect 1830 37775 1864 37791
rect 1830 37723 1864 37736
rect 1830 37702 1864 37723
rect 1830 37655 1864 37663
rect 1830 37629 1864 37655
rect 1830 37587 1864 37590
rect 1830 37556 1864 37587
rect 1830 37485 1864 37517
rect 1830 37483 1864 37485
rect 1830 37417 1864 37444
rect 1830 37410 1864 37417
rect 1830 37349 1864 37371
rect 1830 37337 1864 37349
rect 1830 37281 1864 37298
rect 1830 37264 1864 37281
rect 1830 37213 1864 37225
rect 1830 37191 1864 37213
rect 1830 37145 1864 37152
rect 1830 37118 1864 37145
rect 1830 37077 1864 37079
rect 1830 37045 1864 37077
rect 1830 36975 1864 37006
rect 1830 36972 1864 36975
rect 1830 36907 1864 36933
rect 1830 36899 1864 36907
rect 1830 36839 1864 36860
rect 1830 36826 1864 36839
rect 1830 36771 1864 36787
rect 1830 36753 1864 36771
rect 1830 36703 1864 36714
rect 1830 36680 1864 36703
rect 1830 36635 1864 36641
rect 1830 36607 1864 36635
rect 1830 36567 1864 36568
rect 1830 36534 1864 36567
rect 1830 36465 1864 36495
rect 1830 36461 1864 36465
rect 1830 36397 1864 36422
rect 1830 36388 1864 36397
rect 1830 36329 1864 36349
rect 1830 36315 1864 36329
rect 1830 36261 1864 36276
rect 1830 36242 1864 36261
rect 1830 36193 1864 36203
rect 1830 36169 1864 36193
rect 1830 36125 1864 36130
rect 1830 36096 1864 36125
rect 1830 36023 1864 36057
rect 1830 35955 1864 35984
rect 1830 35950 1864 35955
rect 1830 35887 1864 35911
rect 1830 35877 1864 35887
rect 1830 35819 1864 35838
rect 1830 35804 1864 35819
rect 1830 35751 1864 35765
rect 1830 35731 1864 35751
rect 1830 35683 1864 35692
rect 1830 35658 1864 35683
rect 1830 35615 1864 35619
rect 1830 35585 1864 35615
rect 1830 35513 1864 35546
rect 1830 35512 1864 35513
rect 1830 35445 1864 35473
rect 1830 35439 1864 35445
rect 1830 35377 1864 35400
rect 1830 35366 1864 35377
rect 1830 35309 1864 35327
rect 1830 35293 1864 35309
rect 1830 35241 1864 35254
rect 1830 35220 1864 35241
rect 1830 35173 1864 35181
rect 1830 35147 1864 35173
rect 1830 35105 1864 35109
rect 1830 35075 1864 35105
rect 1830 35003 1864 35037
rect 1830 34935 1864 34965
rect 1830 34931 1864 34935
rect 1830 34867 1864 34893
rect 1830 34859 1864 34867
rect 1830 34799 1864 34821
rect 1830 34787 1864 34799
rect 1830 34731 1864 34749
rect 1830 34715 1864 34731
rect 1830 34663 1864 34677
rect 1830 34643 1864 34663
rect 1830 34595 1864 34605
rect 1830 34571 1864 34595
rect 1830 34527 1864 34533
rect 1830 34499 1864 34527
rect 1830 34459 1864 34461
rect 1830 34427 1864 34459
rect 1830 34357 1864 34389
rect 1830 34355 1864 34357
rect 1830 34289 1864 34317
rect 1830 34283 1864 34289
rect 1830 34221 1864 34245
rect 1830 34211 1864 34221
rect 1830 34153 1864 34173
rect 1830 34139 1864 34153
rect 1830 34085 1864 34101
rect 1830 34067 1864 34085
rect 1830 34017 1864 34029
rect 1830 33995 1864 34017
rect 1830 33949 1864 33957
rect 1830 33923 1864 33949
rect 1830 33881 1864 33885
rect 1830 33851 1864 33881
rect 1830 33779 1864 33813
rect 1830 33711 1864 33741
rect 1830 33707 1864 33711
rect 1830 33643 1864 33669
rect 1830 33635 1864 33643
rect 1830 33575 1864 33597
rect 1830 33563 1864 33575
rect 1830 33507 1864 33525
rect 1830 33491 1864 33507
rect 1830 33439 1864 33453
rect 1830 33419 1864 33439
rect 1830 33371 1864 33381
rect 1830 33347 1864 33371
rect 1830 33303 1864 33309
rect 1830 33275 1864 33303
rect 1830 33235 1864 33237
rect 1830 33203 1864 33235
rect 1830 33133 1864 33165
rect 1830 33131 1864 33133
rect 1830 33065 1864 33093
rect 1830 33059 1864 33065
rect 1830 32997 1864 33021
rect 1830 32987 1864 32997
rect 1830 32929 1864 32949
rect 1830 32915 1864 32929
rect 1830 32861 1864 32877
rect 1830 32843 1864 32861
rect 1830 32793 1864 32805
rect 1830 32771 1864 32793
rect 1830 32725 1864 32733
rect 1830 32699 1864 32725
rect 1830 32657 1864 32661
rect 1830 32627 1864 32657
rect 1830 32555 1864 32589
rect 1830 32487 1864 32517
rect 1830 32483 1864 32487
rect 1830 32419 1864 32445
rect 1830 32411 1864 32419
rect 1830 32351 1864 32373
rect 1830 32339 1864 32351
rect 1830 32283 1864 32301
rect 1830 32267 1864 32283
rect 1830 32215 1864 32229
rect 1830 32195 1864 32215
rect 1830 32147 1864 32157
rect 1830 32123 1864 32147
rect 1830 32079 1864 32085
rect 1830 32051 1864 32079
rect 1830 32011 1864 32013
rect 1830 31979 1864 32011
rect 1830 31909 1864 31941
rect 1830 31907 1864 31909
rect 1830 31841 1864 31869
rect 1830 31835 1864 31841
rect 1830 31773 1864 31797
rect 1830 31763 1864 31773
rect 1830 31705 1864 31725
rect 1830 31691 1864 31705
rect 1830 31637 1864 31653
rect 1830 31619 1864 31637
rect 1830 31569 1864 31581
rect 1830 31547 1864 31569
rect 1830 31501 1864 31509
rect 1830 31475 1864 31501
rect 1830 31433 1864 31437
rect 1830 31403 1864 31433
rect 1830 31331 1864 31365
rect 1830 31263 1864 31293
rect 1830 31259 1864 31263
rect 1830 31195 1864 31221
rect 1830 31187 1864 31195
rect 1830 31127 1864 31149
rect 1830 31115 1864 31127
rect 1830 31059 1864 31077
rect 1830 31043 1864 31059
rect 1830 30991 1864 31005
rect 1830 30971 1864 30991
rect 1830 30923 1864 30933
rect 1830 30899 1864 30923
rect 1830 30855 1864 30861
rect 1830 30827 1864 30855
rect 1830 30787 1864 30789
rect 1830 30755 1864 30787
rect 1830 30685 1864 30717
rect 1830 30683 1864 30685
rect 1830 30617 1864 30645
rect 1830 30611 1864 30617
rect 1830 30549 1864 30573
rect 1830 30539 1864 30549
rect 1830 30481 1864 30501
rect 1830 30467 1864 30481
rect 1830 30413 1864 30429
rect 1830 30395 1864 30413
rect 1830 30345 1864 30357
rect 1830 30323 1864 30345
rect 1830 30277 1864 30285
rect 1830 30251 1864 30277
rect 1830 30209 1864 30213
rect 1830 30179 1864 30209
rect 1830 30107 1864 30141
rect 1830 30039 1864 30069
rect 1830 30035 1864 30039
rect 1830 29971 1864 29997
rect 1830 29963 1864 29971
rect 1830 29903 1864 29925
rect 1830 29891 1864 29903
rect 1830 29835 1864 29853
rect 1830 29819 1864 29835
rect 1830 29767 1864 29781
rect 1830 29747 1864 29767
rect 1830 29699 1864 29709
rect 1830 29675 1864 29699
rect 1830 29631 1864 29637
rect 1830 29603 1864 29631
rect 1830 29563 1864 29565
rect 1830 29531 1864 29563
rect 1830 29461 1864 29493
rect 1830 29459 1864 29461
rect 1830 29393 1864 29421
rect 1830 29387 1864 29393
rect 1830 29325 1864 29349
rect 1830 29315 1864 29325
rect 1830 29257 1864 29277
rect 1830 29243 1864 29257
rect 1830 29189 1864 29205
rect 1830 29171 1864 29189
rect 1830 29121 1864 29133
rect 1830 29099 1864 29121
rect 1830 29053 1864 29061
rect 1830 29027 1864 29053
rect 1830 28985 1864 28989
rect 1830 28955 1864 28985
rect 1830 28883 1864 28917
rect 1830 28815 1864 28845
rect 1830 28811 1864 28815
rect 1830 28747 1864 28773
rect 1830 28739 1864 28747
rect 1830 28679 1864 28701
rect 1830 28667 1864 28679
rect 1830 28611 1864 28629
rect 1830 28595 1864 28611
rect 1830 28543 1864 28557
rect 1830 28523 1864 28543
rect 1830 28475 1864 28485
rect 1830 28451 1864 28475
rect 1830 28407 1864 28413
rect 1830 28379 1864 28407
rect 1830 28339 1864 28341
rect 1830 28307 1864 28339
rect 1830 28237 1864 28269
rect 1830 28235 1864 28237
rect 1830 28169 1864 28197
rect 1830 28163 1864 28169
rect 1830 28101 1864 28125
rect 1830 28091 1864 28101
rect 1830 28033 1864 28053
rect 1830 28019 1864 28033
rect 1830 27965 1864 27981
rect 1830 27947 1864 27965
rect 1830 27897 1864 27909
rect 1830 27875 1864 27897
rect 1830 27829 1864 27837
rect 1830 27803 1864 27829
rect 1830 27761 1864 27765
rect 1830 27731 1864 27761
rect 1830 27659 1864 27693
rect 1830 27591 1864 27621
rect 1830 27587 1864 27591
rect 1830 27523 1864 27549
rect 1830 27515 1864 27523
rect 1830 27455 1864 27477
rect 1830 27443 1864 27455
rect 1830 27387 1864 27405
rect 1830 27371 1864 27387
rect 1830 27319 1864 27333
rect 1830 27299 1864 27319
rect 1830 27251 1864 27261
rect 1830 27227 1864 27251
rect 1830 27183 1864 27189
rect 1830 27155 1864 27183
rect 1830 27115 1864 27117
rect 1830 27083 1864 27115
rect 1830 27013 1864 27045
rect 1830 27011 1864 27013
rect 1830 26945 1864 26973
rect 1830 26939 1864 26945
rect 1830 26877 1864 26901
rect 1830 26867 1864 26877
rect 1830 26809 1864 26829
rect 1830 26795 1864 26809
rect 1830 26741 1864 26757
rect 1830 26723 1864 26741
rect 1830 26673 1864 26685
rect 1830 26651 1864 26673
rect 1830 26605 1864 26613
rect 1830 26579 1864 26605
rect 1830 26537 1864 26541
rect 1830 26507 1864 26537
rect 1830 26435 1864 26469
rect 1830 26367 1864 26397
rect 1830 26363 1864 26367
rect 1830 26299 1864 26325
rect 1830 26291 1864 26299
rect 1830 26231 1864 26253
rect 1830 26219 1864 26231
rect 1830 26163 1864 26181
rect 1830 26147 1864 26163
rect 1830 26095 1864 26109
rect 1830 26075 1864 26095
rect 1830 26027 1864 26037
rect 1830 26003 1864 26027
rect 1830 25959 1864 25965
rect 1830 25931 1864 25959
rect 1830 25891 1864 25893
rect 1830 25859 1864 25891
rect 1830 25789 1864 25821
rect 1830 25787 1864 25789
rect 1830 25721 1864 25749
rect 1830 25715 1864 25721
rect 1830 25653 1864 25677
rect 1830 25643 1864 25653
rect 1830 25585 1864 25605
rect 1830 25571 1864 25585
rect 1830 25517 1864 25533
rect 1830 25499 1864 25517
rect 1830 25449 1864 25461
rect 1830 25427 1864 25449
rect 1830 25381 1864 25389
rect 1830 25355 1864 25381
rect 1830 25313 1864 25317
rect 1830 25283 1864 25313
rect 1830 25211 1864 25245
rect 1830 25143 1864 25173
rect 1830 25139 1864 25143
rect 1830 25075 1864 25101
rect 1830 25067 1864 25075
rect 1830 25007 1864 25029
rect 1830 24995 1864 25007
rect 1830 24939 1864 24957
rect 1830 24923 1864 24939
rect 1830 24871 1864 24885
rect 1830 24851 1864 24871
rect 1830 24803 1864 24813
rect 1830 24779 1864 24803
rect 1830 24735 1864 24741
rect 1830 24707 1864 24735
rect 1830 24667 1864 24669
rect 1830 24635 1864 24667
rect 1830 24565 1864 24597
rect 1830 24563 1864 24565
rect 1830 24497 1864 24525
rect 1830 24491 1864 24497
rect 1830 24429 1864 24453
rect 1830 24419 1864 24429
rect 1830 24361 1864 24381
rect 1830 24347 1864 24361
rect 1830 24293 1864 24309
rect 1830 24275 1864 24293
rect 1830 24225 1864 24237
rect 1830 24203 1864 24225
rect 1830 24157 1864 24165
rect 1830 24131 1864 24157
rect 1830 24089 1864 24093
rect 1830 24059 1864 24089
rect 1830 23987 1864 24021
rect 1830 23919 1864 23949
rect 1830 23915 1864 23919
rect 1830 23851 1864 23877
rect 1830 23843 1864 23851
rect 1830 23783 1864 23805
rect 1830 23771 1864 23783
rect 1830 23715 1864 23733
rect 1830 23699 1864 23715
rect 1830 23647 1864 23661
rect 1830 23627 1864 23647
rect 1830 23579 1864 23589
rect 1830 23555 1864 23579
rect 1830 23511 1864 23517
rect 1830 23483 1864 23511
rect 1830 23443 1864 23445
rect 1830 23411 1864 23443
rect 1830 23341 1864 23373
rect 1830 23339 1864 23341
rect 1830 23273 1864 23301
rect 1830 23267 1864 23273
rect 1830 23205 1864 23229
rect 1830 23195 1864 23205
rect 1830 23137 1864 23157
rect 1830 23123 1864 23137
rect 1830 23069 1864 23085
rect 1830 23051 1864 23069
rect 1830 23001 1864 23013
rect 1830 22979 1864 23001
rect 1830 22933 1864 22941
rect 1830 22907 1864 22933
rect 1830 22865 1864 22869
rect 1830 22835 1864 22865
rect 1830 22763 1864 22797
rect 1830 22695 1864 22725
rect 1830 22691 1864 22695
rect 1830 22627 1864 22653
rect 1830 22619 1864 22627
rect 1830 22559 1864 22581
rect 1830 22547 1864 22559
rect 1830 22491 1864 22509
rect 1830 22475 1864 22491
rect 1830 22423 1864 22437
rect 1830 22403 1864 22423
rect 1830 22355 1864 22365
rect 1830 22331 1864 22355
rect 1830 22287 1864 22293
rect 1830 22259 1864 22287
rect 1830 22219 1864 22221
rect 1830 22187 1864 22219
rect 1830 22117 1864 22149
rect 1830 22115 1864 22117
rect 1830 22049 1864 22077
rect 1830 22043 1864 22049
rect 1830 21981 1864 22005
rect 1830 21971 1864 21981
rect 1830 21913 1864 21933
rect 1830 21899 1864 21913
rect 1830 21845 1864 21861
rect 1830 21827 1864 21845
rect 1830 21777 1864 21789
rect 1830 21755 1864 21777
rect 1830 21709 1864 21717
rect 1830 21683 1864 21709
rect 1830 21641 1864 21645
rect 1830 21611 1864 21641
rect 1830 21539 1864 21573
rect 1830 21471 1864 21501
rect 1830 21467 1864 21471
rect 1830 21403 1864 21429
rect 1830 21395 1864 21403
rect 1830 21335 1864 21357
rect 1830 21323 1864 21335
rect 1830 21267 1864 21285
rect 1830 21251 1864 21267
rect 1830 21199 1864 21213
rect 1830 21179 1864 21199
rect 1830 21131 1864 21141
rect 1830 21107 1864 21131
rect 1830 21063 1864 21069
rect 1830 21035 1864 21063
rect 1830 20995 1864 20997
rect 1830 20963 1864 20995
rect 1830 20893 1864 20925
rect 1830 20891 1864 20893
rect 1830 20825 1864 20853
rect 1830 20819 1864 20825
rect 1830 20757 1864 20781
rect 1830 20747 1864 20757
rect 1830 20689 1864 20709
rect 1830 20675 1864 20689
rect 1830 20621 1864 20637
rect 1830 20603 1864 20621
rect 1830 20553 1864 20565
rect 1830 20531 1864 20553
rect 1830 20485 1864 20493
rect 1830 20459 1864 20485
rect 1830 20417 1864 20421
rect 1830 20387 1864 20417
rect 1830 20315 1864 20349
rect 1830 20247 1864 20277
rect 1830 20243 1864 20247
rect 1830 20179 1864 20205
rect 1830 20171 1864 20179
rect 1830 20111 1864 20133
rect 1830 20099 1864 20111
rect 1830 20043 1864 20061
rect 1830 20027 1864 20043
rect 1830 19975 1864 19989
rect 1830 19955 1864 19975
rect 1830 19907 1864 19917
rect 1830 19883 1864 19907
rect 1830 19839 1864 19845
rect 1830 19811 1864 19839
rect 1830 19771 1864 19773
rect 1830 19739 1864 19771
rect 1830 19669 1864 19701
rect 1830 19667 1864 19669
rect 1830 19601 1864 19629
rect 1830 19595 1864 19601
rect 1830 19533 1864 19557
rect 1830 19523 1864 19533
rect 1830 19465 1864 19485
rect 1830 19451 1864 19465
rect 1830 19397 1864 19413
rect 1830 19379 1864 19397
rect 1830 19329 1864 19341
rect 1830 19307 1864 19329
rect 1830 19261 1864 19269
rect 1830 19235 1864 19261
rect 1830 19193 1864 19197
rect 1830 19163 1864 19193
rect 1830 19091 1864 19125
rect 1830 19023 1864 19053
rect 1830 19019 1864 19023
rect 1830 18955 1864 18981
rect 1830 18947 1864 18955
rect 1830 18887 1864 18909
rect 1830 18875 1864 18887
rect 1830 18819 1864 18837
rect 1830 18803 1864 18819
rect 1830 18751 1864 18765
rect 1830 18731 1864 18751
rect 1830 18683 1864 18693
rect 1830 18659 1864 18683
rect 1830 18615 1864 18621
rect 1830 18587 1864 18615
rect 1830 18547 1864 18549
rect 1830 18515 1864 18547
rect 1830 18445 1864 18477
rect 1830 18443 1864 18445
rect 1830 18377 1864 18405
rect 1830 18371 1864 18377
rect 1830 18309 1864 18333
rect 1830 18299 1864 18309
rect 1830 18241 1864 18261
rect 1830 18227 1864 18241
rect 1830 18173 1864 18189
rect 1830 18155 1864 18173
rect 1830 18105 1864 18117
rect 1830 18083 1864 18105
rect 1830 18037 1864 18045
rect 1830 18011 1864 18037
rect 1830 17969 1864 17973
rect 1830 17939 1864 17969
rect 1830 17867 1864 17901
rect 1830 17799 1864 17829
rect 1830 17795 1864 17799
rect 1830 17731 1864 17757
rect 1830 17723 1864 17731
rect 1830 17663 1864 17685
rect 1830 17651 1864 17663
rect 1830 17595 1864 17613
rect 1830 17579 1864 17595
rect 1830 17527 1864 17541
rect 1830 17507 1864 17527
rect 1830 17459 1864 17469
rect 1830 17435 1864 17459
rect 1830 17391 1864 17397
rect 1830 17363 1864 17391
rect 1830 17323 1864 17325
rect 1830 17291 1864 17323
rect 1830 17221 1864 17253
rect 1830 17219 1864 17221
rect 1830 17153 1864 17181
rect 1830 17147 1864 17153
rect 1830 17085 1864 17109
rect 1830 17075 1864 17085
rect 1830 17017 1864 17037
rect 1830 17003 1864 17017
rect 1830 16949 1864 16965
rect 1830 16931 1864 16949
rect 1830 16881 1864 16893
rect 1830 16859 1864 16881
rect 1830 16813 1864 16821
rect 1830 16787 1864 16813
rect 1830 16745 1864 16749
rect 1830 16715 1864 16745
rect 1830 16643 1864 16677
rect 1830 16575 1864 16605
rect 1830 16571 1864 16575
rect 1830 16507 1864 16533
rect 1830 16499 1864 16507
rect 1830 16439 1864 16461
rect 1830 16427 1864 16439
rect 1830 16371 1864 16389
rect 1830 16355 1864 16371
rect 1830 16303 1864 16317
rect 1830 16283 1864 16303
rect 1830 16235 1864 16245
rect 1830 16211 1864 16235
rect 1830 16167 1864 16173
rect 1830 16139 1864 16167
rect 1830 16099 1864 16101
rect 1830 16067 1864 16099
rect 1830 15997 1864 16029
rect 1830 15995 1864 15997
rect 1830 15929 1864 15957
rect 1830 15923 1864 15929
rect 1830 15861 1864 15885
rect 1830 15851 1864 15861
rect 1830 15793 1864 15813
rect 1830 15779 1864 15793
rect 1830 15725 1864 15741
rect 1830 15707 1864 15725
rect 1830 15657 1864 15669
rect 1830 15635 1864 15657
rect 1830 15589 1864 15597
rect 1830 15563 1864 15589
rect 1830 15521 1864 15525
rect 1830 15491 1864 15521
rect 1830 15419 1864 15453
rect 1830 15351 1864 15381
rect 1830 15347 1864 15351
rect 1830 15283 1864 15309
rect 1830 15275 1864 15283
rect 1830 15215 1864 15237
rect 1830 15203 1864 15215
rect 1830 15147 1864 15165
rect 1830 15131 1864 15147
rect 1830 15079 1864 15093
rect 1830 15059 1864 15079
rect 1830 15011 1864 15021
rect 1830 14987 1864 15011
rect 1830 14943 1864 14949
rect 1830 14915 1864 14943
rect 1830 14875 1864 14877
rect 1830 14843 1864 14875
rect 1830 14773 1864 14805
rect 1830 14771 1864 14773
rect 1830 14705 1864 14733
rect 1830 14699 1864 14705
rect 1830 14637 1864 14661
rect 1830 14627 1864 14637
rect 1830 14569 1864 14589
rect 1830 14555 1864 14569
rect 1830 14501 1864 14517
rect 1830 14483 1864 14501
rect 1830 14433 1864 14445
rect 1830 14411 1864 14433
rect 1830 14365 1864 14373
rect 1830 14339 1864 14365
rect 1830 14297 1864 14301
rect 1830 14267 1864 14297
rect 1830 14195 1864 14229
rect 1830 14127 1864 14157
rect 1830 14123 1864 14127
rect 1830 14059 1864 14085
rect 1830 14051 1864 14059
rect 1830 13991 1864 14013
rect 1830 13979 1864 13991
rect 1830 13923 1864 13941
rect 1830 13907 1864 13923
rect 1830 13855 1864 13869
rect 1830 13835 1864 13855
rect 1830 13787 1864 13797
rect 1830 13763 1864 13787
rect 1830 13719 1864 13725
rect 1830 13691 1864 13719
rect 1830 13651 1864 13653
rect 1830 13619 1864 13651
rect 1830 13549 1864 13581
rect 1830 13547 1864 13549
rect 1830 13481 1864 13509
rect 1830 13475 1864 13481
rect 1830 13413 1864 13437
rect 1830 13403 1864 13413
rect 1830 13345 1864 13365
rect 1830 13331 1864 13345
rect 1830 13277 1864 13293
rect 1830 13259 1864 13277
rect 1830 13209 1864 13221
rect 1830 13187 1864 13209
rect 1830 13141 1864 13149
rect 1830 13115 1864 13141
rect 1830 13073 1864 13077
rect 1830 13043 1864 13073
rect 1830 12971 1864 13005
rect 1830 12903 1864 12933
rect 1830 12899 1864 12903
rect 1830 12835 1864 12861
rect 1830 12827 1864 12835
rect 1830 12767 1864 12789
rect 1830 12755 1864 12767
rect 1830 12699 1864 12717
rect 1830 12683 1864 12699
rect 1830 12631 1864 12645
rect 1830 12611 1864 12631
rect 1830 12563 1864 12573
rect 1830 12539 1864 12563
rect 1830 12495 1864 12501
rect 1830 12467 1864 12495
rect 1830 12427 1864 12429
rect 1830 12395 1864 12427
rect 1830 12325 1864 12357
rect 1830 12323 1864 12325
rect 1830 12257 1864 12285
rect 1830 12251 1864 12257
rect 1830 12189 1864 12213
rect 1830 12179 1864 12189
rect 1830 12121 1864 12141
rect 1830 12107 1864 12121
rect 1830 12053 1864 12069
rect 1830 12035 1864 12053
rect 1830 11985 1864 11997
rect 1830 11963 1864 11985
rect 1830 11917 1864 11925
rect 1830 11891 1864 11917
rect 1830 11849 1864 11853
rect 1830 11819 1864 11849
rect 1830 11747 1864 11781
rect 1830 11679 1864 11709
rect 1830 11675 1864 11679
rect 1830 11611 1864 11637
rect 1830 11603 1864 11611
rect 1830 11543 1864 11565
rect 1830 11531 1864 11543
rect 1830 11475 1864 11493
rect 1830 11459 1864 11475
rect 1830 11407 1864 11421
rect 1830 11387 1864 11407
rect 1830 11339 1864 11349
rect 1830 11315 1864 11339
rect 1830 11271 1864 11277
rect 1830 11243 1864 11271
rect 1830 11203 1864 11205
rect 1830 11171 1864 11203
rect 1830 11101 1864 11133
rect 1830 11099 1864 11101
rect 1830 11033 1864 11061
rect 1830 11027 1864 11033
rect 1830 10965 1864 10989
rect 1830 10955 1864 10965
rect 1830 10897 1864 10917
rect 1830 10883 1864 10897
rect 1830 10829 1864 10845
rect 1830 10811 1864 10829
rect 1830 10761 1864 10773
rect 1830 10739 1864 10761
rect 1830 10693 1864 10701
rect 1830 10667 1864 10693
rect 1830 10625 1864 10629
rect 1830 10595 1864 10625
rect 1830 10523 1864 10557
rect 1830 10455 1864 10485
rect 1830 10451 1864 10455
rect 1830 10387 1864 10413
rect 1830 10379 1864 10387
rect 1830 10319 1864 10341
rect 1830 10307 1864 10319
rect 1830 10251 1864 10269
rect 1830 10235 1864 10251
rect 1830 10183 1864 10197
rect 1830 10163 1864 10183
rect 1830 10115 1864 10125
rect 1830 10091 1864 10115
rect 1830 10047 1864 10053
rect 1830 10019 1864 10047
rect 1830 9979 1864 9981
rect 1830 9947 1864 9979
rect 1830 9877 1864 9909
rect 1830 9875 1864 9877
rect 1830 9809 1864 9837
rect 1830 9803 1864 9809
rect 1830 9741 1864 9765
rect 1830 9731 1864 9741
rect 1830 9673 1864 9693
rect 1830 9659 1864 9673
rect 1830 9605 1864 9621
rect 1830 9587 1864 9605
rect 1830 9537 1864 9549
rect 1830 9515 1864 9537
rect 1830 9469 1864 9477
rect 1830 9443 1864 9469
rect 1830 9401 1864 9405
rect 1830 9371 1864 9401
rect 1830 9299 1864 9333
rect 1830 9231 1864 9261
rect 1830 9227 1864 9231
rect 1830 9163 1864 9189
rect 1830 9155 1864 9163
rect 1830 9095 1864 9117
rect 1830 9083 1864 9095
rect 1830 9027 1864 9045
rect 1830 9011 1864 9027
rect 1830 8959 1864 8973
rect 1830 8939 1864 8959
rect 1830 8891 1864 8901
rect 1830 8867 1864 8891
rect 1830 8823 1864 8829
rect 1830 8795 1864 8823
rect 1830 8755 1864 8757
rect 1830 8723 1864 8755
rect 1830 8653 1864 8685
rect 1830 8651 1864 8653
rect 1830 8585 1864 8613
rect 1830 8579 1864 8585
rect 1830 8517 1864 8541
rect 1830 8507 1864 8517
rect 1830 8449 1864 8469
rect 1830 8435 1864 8449
rect 1830 8381 1864 8397
rect 1830 8363 1864 8381
rect 1830 8313 1864 8325
rect 1830 8291 1864 8313
rect 1830 8245 1864 8253
rect 1830 8219 1864 8245
rect 1830 8177 1864 8181
rect 1830 8147 1864 8177
rect 1830 8075 1864 8109
rect 1830 8007 1864 8037
rect 1830 8003 1864 8007
rect 1830 7939 1864 7965
rect 1830 7931 1864 7939
rect 1830 7871 1864 7893
rect 1830 7859 1864 7871
rect 1830 7803 1864 7821
rect 1830 7787 1864 7803
rect 1830 7735 1864 7749
rect 1830 7715 1864 7735
rect 1830 7667 1864 7677
rect 1830 7643 1864 7667
rect 1830 7599 1864 7605
rect 1830 7571 1864 7599
rect 1830 7531 1864 7533
rect 1830 7499 1864 7531
rect 1830 7429 1864 7461
rect 1830 7427 1864 7429
rect 1830 7361 1864 7389
rect 1830 7355 1864 7361
rect 1830 7293 1864 7317
rect 1830 7283 1864 7293
rect 1830 7225 1864 7245
rect 1830 7211 1864 7225
rect 1830 7157 1864 7173
rect 1830 7139 1864 7157
rect 1830 7089 1864 7101
rect 1830 7067 1864 7089
rect 1830 7021 1864 7029
rect 1830 6995 1864 7021
rect 1830 6953 1864 6957
rect 1830 6923 1864 6953
rect 1830 6851 1864 6885
rect 1830 6783 1864 6813
rect 1830 6779 1864 6783
rect 1830 6715 1864 6741
rect 1830 6707 1864 6715
rect 1830 6647 1864 6669
rect 1830 6635 1864 6647
rect 1830 6579 1864 6597
rect 1830 6563 1864 6579
rect 1830 6511 1864 6525
rect 1830 6491 1864 6511
rect 1830 6443 1864 6453
rect 1830 6419 1864 6443
rect 1830 6375 1864 6381
rect 1830 6347 1864 6375
rect 1830 6307 1864 6309
rect 1830 6275 1864 6307
rect 1830 6205 1864 6237
rect 1830 6203 1864 6205
rect 1830 6137 1864 6165
rect 1830 6131 1864 6137
rect 1830 6069 1864 6093
rect 1830 6059 1864 6069
rect 1830 6001 1864 6021
rect 1830 5987 1864 6001
rect 1830 5933 1864 5949
rect 1830 5915 1864 5933
rect 1830 5865 1864 5877
rect 1830 5843 1864 5865
rect 1830 5797 1864 5805
rect 1830 5771 1864 5797
rect 1830 5729 1864 5733
rect 1830 5699 1864 5729
rect 1830 5627 1864 5661
rect 1830 5559 1864 5589
rect 1830 5555 1864 5559
rect 1830 5491 1864 5517
rect 1830 5483 1864 5491
rect 1830 5423 1864 5445
rect 1830 5411 1864 5423
rect 1830 5355 1864 5373
rect 1830 5339 1864 5355
rect 1830 5287 1864 5301
rect 1830 5267 1864 5287
rect 1830 5219 1864 5229
rect 1830 5195 1864 5219
rect 1830 5151 1864 5157
rect 1830 5123 1864 5151
rect 1830 5083 1864 5085
rect 1830 5051 1864 5083
rect 1830 4981 1864 5013
rect 1830 4979 1864 4981
rect 1830 4913 1864 4941
rect 1830 4907 1864 4913
rect 1830 4845 1864 4869
rect 1830 4835 1864 4845
rect 1830 4777 1864 4797
rect 1830 4763 1864 4777
rect 1830 4709 1864 4725
rect 1830 4691 1864 4709
rect 1830 4641 1864 4653
rect 1830 4619 1864 4641
rect 1830 4573 1864 4581
rect 1830 4547 1864 4573
rect 1830 4505 1864 4509
rect 1830 4475 1864 4505
rect 1830 4403 1864 4437
rect 1830 4335 1864 4365
rect 1830 4331 1864 4335
rect 1830 4267 1864 4293
rect 1830 4259 1864 4267
rect 1830 4199 1864 4221
rect 1830 4187 1864 4199
rect 1830 4131 1864 4149
rect 1830 4115 1864 4131
rect 1830 4063 1864 4077
rect 1830 4043 1864 4063
rect 1830 3995 1864 4005
rect 1830 3971 1864 3995
rect 1830 3927 1864 3933
rect 1830 3899 1864 3927
rect 1830 3859 1864 3861
rect 1830 3827 1864 3859
rect 1830 3757 1864 3789
rect 1830 3755 1864 3757
rect 1830 3689 1864 3717
rect 1830 3683 1864 3689
rect 1830 3621 1864 3645
rect 1830 3611 1864 3621
rect 1830 3553 1864 3573
rect 1830 3539 1864 3553
rect -252 3397 -218 3429
rect -252 3395 -218 3397
rect -126 3452 -92 3486
rect -126 3394 -92 3414
rect -126 3380 -92 3394
rect -8 3452 26 3486
rect -8 3394 26 3414
rect -8 3380 26 3394
rect 110 3452 144 3486
rect 110 3394 144 3414
rect 110 3380 144 3394
rect 228 3452 262 3486
rect 228 3394 262 3414
rect 228 3380 262 3394
rect 346 3452 380 3486
rect 346 3394 380 3414
rect 346 3380 380 3394
rect 464 3452 498 3486
rect 464 3394 498 3414
rect 464 3380 498 3394
rect 582 3452 616 3486
rect 582 3394 616 3414
rect 582 3380 616 3394
rect 700 3452 734 3486
rect 700 3394 734 3414
rect 700 3380 734 3394
rect 818 3452 852 3486
rect 818 3394 852 3414
rect 818 3380 852 3394
rect 936 3452 970 3486
rect 936 3394 970 3414
rect 936 3380 970 3394
rect 1054 3452 1088 3486
rect 1054 3394 1088 3414
rect 1054 3380 1088 3394
rect 1172 3452 1206 3486
rect 1172 3394 1206 3414
rect 1172 3380 1206 3394
rect 1290 3452 1324 3486
rect 1290 3394 1324 3414
rect 1290 3380 1324 3394
rect 1408 3452 1442 3486
rect 1408 3394 1442 3414
rect 1408 3380 1442 3394
rect 1526 3452 1560 3486
rect 1526 3394 1560 3414
rect 1526 3380 1560 3394
rect 1644 3452 1678 3486
rect 1644 3394 1678 3414
rect 1644 3380 1678 3394
rect 1830 3485 1864 3501
rect 1830 3467 1864 3485
rect 3972 38655 4006 38685
rect 3972 38651 4006 38655
rect 3972 38587 4006 38612
rect 3972 38578 4006 38587
rect 3972 38519 4006 38539
rect 3972 38505 4006 38519
rect 3972 38451 4006 38466
rect 3972 38432 4006 38451
rect 3972 38383 4006 38393
rect 3972 38359 4006 38383
rect 3972 38315 4006 38320
rect 3972 38286 4006 38315
rect 3972 38213 4006 38247
rect 3972 38145 4006 38174
rect 3972 38140 4006 38145
rect 3972 38077 4006 38101
rect 3972 38067 4006 38077
rect 3972 38009 4006 38028
rect 3972 37994 4006 38009
rect 3972 37941 4006 37955
rect 3972 37921 4006 37941
rect 3972 37873 4006 37882
rect 3972 37848 4006 37873
rect 3972 37805 4006 37809
rect 3972 37775 4006 37805
rect 3972 37703 4006 37736
rect 3972 37702 4006 37703
rect 3972 37635 4006 37663
rect 3972 37629 4006 37635
rect 3972 37567 4006 37590
rect 3972 37556 4006 37567
rect 3972 37499 4006 37517
rect 3972 37483 4006 37499
rect 3972 37431 4006 37444
rect 3972 37410 4006 37431
rect 3972 37363 4006 37371
rect 3972 37337 4006 37363
rect 3972 37295 4006 37298
rect 3972 37264 4006 37295
rect 3972 37193 4006 37225
rect 3972 37191 4006 37193
rect 3972 37125 4006 37152
rect 3972 37118 4006 37125
rect 3972 37057 4006 37079
rect 3972 37045 4006 37057
rect 3972 36989 4006 37006
rect 3972 36972 4006 36989
rect 3972 36921 4006 36933
rect 3972 36899 4006 36921
rect 3972 36853 4006 36860
rect 3972 36826 4006 36853
rect 3972 36785 4006 36787
rect 3972 36753 4006 36785
rect 3972 36683 4006 36714
rect 3972 36680 4006 36683
rect 3972 36615 4006 36641
rect 3972 36607 4006 36615
rect 3972 36547 4006 36568
rect 3972 36534 4006 36547
rect 3972 36479 4006 36495
rect 3972 36461 4006 36479
rect 3972 36411 4006 36422
rect 3972 36388 4006 36411
rect 3972 36343 4006 36349
rect 3972 36315 4006 36343
rect 3972 36275 4006 36276
rect 3972 36242 4006 36275
rect 3972 36173 4006 36203
rect 3972 36169 4006 36173
rect 3972 36105 4006 36130
rect 3972 36096 4006 36105
rect 3972 36037 4006 36057
rect 3972 36023 4006 36037
rect 3972 35969 4006 35984
rect 3972 35950 4006 35969
rect 3972 35901 4006 35911
rect 3972 35877 4006 35901
rect 3972 35833 4006 35838
rect 3972 35804 4006 35833
rect 3972 35731 4006 35765
rect 3972 35663 4006 35692
rect 3972 35658 4006 35663
rect 3972 35595 4006 35619
rect 3972 35585 4006 35595
rect 3972 35527 4006 35546
rect 3972 35512 4006 35527
rect 3972 35459 4006 35473
rect 3972 35439 4006 35459
rect 3972 35391 4006 35400
rect 3972 35366 4006 35391
rect 3972 35323 4006 35327
rect 3972 35293 4006 35323
rect 3972 35221 4006 35254
rect 3972 35220 4006 35221
rect 3972 35153 4006 35181
rect 3972 35147 4006 35153
rect 3972 35085 4006 35109
rect 3972 35075 4006 35085
rect 3972 35017 4006 35037
rect 3972 35003 4006 35017
rect 3972 34949 4006 34965
rect 3972 34931 4006 34949
rect 3972 34881 4006 34893
rect 3972 34859 4006 34881
rect 3972 34813 4006 34821
rect 3972 34787 4006 34813
rect 3972 34745 4006 34749
rect 3972 34715 4006 34745
rect 3972 34643 4006 34677
rect 3972 34575 4006 34605
rect 3972 34571 4006 34575
rect 3972 34507 4006 34533
rect 3972 34499 4006 34507
rect 3972 34439 4006 34461
rect 3972 34427 4006 34439
rect 3972 34371 4006 34389
rect 3972 34355 4006 34371
rect 3972 34303 4006 34317
rect 3972 34283 4006 34303
rect 3972 34235 4006 34245
rect 3972 34211 4006 34235
rect 3972 34167 4006 34173
rect 3972 34139 4006 34167
rect 3972 34099 4006 34101
rect 3972 34067 4006 34099
rect 3972 33997 4006 34029
rect 3972 33995 4006 33997
rect 3972 33929 4006 33957
rect 3972 33923 4006 33929
rect 3972 33861 4006 33885
rect 3972 33851 4006 33861
rect 3972 33793 4006 33813
rect 3972 33779 4006 33793
rect 3972 33725 4006 33741
rect 3972 33707 4006 33725
rect 3972 33657 4006 33669
rect 3972 33635 4006 33657
rect 3972 33589 4006 33597
rect 3972 33563 4006 33589
rect 3972 33521 4006 33525
rect 3972 33491 4006 33521
rect 3972 33419 4006 33453
rect 3972 33351 4006 33381
rect 3972 33347 4006 33351
rect 3972 33283 4006 33309
rect 3972 33275 4006 33283
rect 3972 33215 4006 33237
rect 3972 33203 4006 33215
rect 3972 33147 4006 33165
rect 3972 33131 4006 33147
rect 3972 33079 4006 33093
rect 3972 33059 4006 33079
rect 3972 33011 4006 33021
rect 3972 32987 4006 33011
rect 3972 32943 4006 32949
rect 3972 32915 4006 32943
rect 3972 32875 4006 32877
rect 3972 32843 4006 32875
rect 3972 32773 4006 32805
rect 3972 32771 4006 32773
rect 3972 32705 4006 32733
rect 3972 32699 4006 32705
rect 3972 32637 4006 32661
rect 3972 32627 4006 32637
rect 3972 32569 4006 32589
rect 3972 32555 4006 32569
rect 3972 32501 4006 32517
rect 3972 32483 4006 32501
rect 3972 32433 4006 32445
rect 3972 32411 4006 32433
rect 3972 32365 4006 32373
rect 3972 32339 4006 32365
rect 3972 32297 4006 32301
rect 3972 32267 4006 32297
rect 3972 32195 4006 32229
rect 3972 32127 4006 32157
rect 3972 32123 4006 32127
rect 3972 32059 4006 32085
rect 3972 32051 4006 32059
rect 3972 31991 4006 32013
rect 3972 31979 4006 31991
rect 3972 31923 4006 31941
rect 3972 31907 4006 31923
rect 3972 31855 4006 31869
rect 3972 31835 4006 31855
rect 3972 31787 4006 31797
rect 3972 31763 4006 31787
rect 3972 31719 4006 31725
rect 3972 31691 4006 31719
rect 3972 31651 4006 31653
rect 3972 31619 4006 31651
rect 3972 31549 4006 31581
rect 3972 31547 4006 31549
rect 3972 31481 4006 31509
rect 3972 31475 4006 31481
rect 3972 31413 4006 31437
rect 3972 31403 4006 31413
rect 3972 31345 4006 31365
rect 3972 31331 4006 31345
rect 3972 31277 4006 31293
rect 3972 31259 4006 31277
rect 3972 31209 4006 31221
rect 3972 31187 4006 31209
rect 3972 31141 4006 31149
rect 3972 31115 4006 31141
rect 3972 31073 4006 31077
rect 3972 31043 4006 31073
rect 3972 30971 4006 31005
rect 3972 30903 4006 30933
rect 3972 30899 4006 30903
rect 3972 30835 4006 30861
rect 3972 30827 4006 30835
rect 3972 30767 4006 30789
rect 3972 30755 4006 30767
rect 3972 30699 4006 30717
rect 3972 30683 4006 30699
rect 3972 30631 4006 30645
rect 3972 30611 4006 30631
rect 3972 30563 4006 30573
rect 3972 30539 4006 30563
rect 3972 30495 4006 30501
rect 3972 30467 4006 30495
rect 3972 30427 4006 30429
rect 3972 30395 4006 30427
rect 3972 30325 4006 30357
rect 3972 30323 4006 30325
rect 3972 30257 4006 30285
rect 3972 30251 4006 30257
rect 3972 30189 4006 30213
rect 3972 30179 4006 30189
rect 3972 30121 4006 30141
rect 3972 30107 4006 30121
rect 3972 30053 4006 30069
rect 3972 30035 4006 30053
rect 3972 29985 4006 29997
rect 3972 29963 4006 29985
rect 3972 29917 4006 29925
rect 3972 29891 4006 29917
rect 3972 29849 4006 29853
rect 3972 29819 4006 29849
rect 3972 29747 4006 29781
rect 3972 29679 4006 29709
rect 3972 29675 4006 29679
rect 3972 29611 4006 29637
rect 3972 29603 4006 29611
rect 3972 29543 4006 29565
rect 3972 29531 4006 29543
rect 3972 29475 4006 29493
rect 3972 29459 4006 29475
rect 3972 29407 4006 29421
rect 3972 29387 4006 29407
rect 3972 29339 4006 29349
rect 3972 29315 4006 29339
rect 3972 29271 4006 29277
rect 3972 29243 4006 29271
rect 3972 29203 4006 29205
rect 3972 29171 4006 29203
rect 3972 29101 4006 29133
rect 3972 29099 4006 29101
rect 3972 29033 4006 29061
rect 3972 29027 4006 29033
rect 3972 28965 4006 28989
rect 3972 28955 4006 28965
rect 3972 28897 4006 28917
rect 3972 28883 4006 28897
rect 3972 28829 4006 28845
rect 3972 28811 4006 28829
rect 3972 28761 4006 28773
rect 3972 28739 4006 28761
rect 3972 28693 4006 28701
rect 3972 28667 4006 28693
rect 3972 28625 4006 28629
rect 3972 28595 4006 28625
rect 3972 28523 4006 28557
rect 3972 28455 4006 28485
rect 3972 28451 4006 28455
rect 3972 28387 4006 28413
rect 3972 28379 4006 28387
rect 3972 28319 4006 28341
rect 3972 28307 4006 28319
rect 3972 28251 4006 28269
rect 3972 28235 4006 28251
rect 3972 28183 4006 28197
rect 3972 28163 4006 28183
rect 3972 28115 4006 28125
rect 3972 28091 4006 28115
rect 3972 28047 4006 28053
rect 3972 28019 4006 28047
rect 3972 27979 4006 27981
rect 3972 27947 4006 27979
rect 3972 27877 4006 27909
rect 3972 27875 4006 27877
rect 3972 27809 4006 27837
rect 3972 27803 4006 27809
rect 3972 27741 4006 27765
rect 3972 27731 4006 27741
rect 3972 27673 4006 27693
rect 3972 27659 4006 27673
rect 3972 27605 4006 27621
rect 3972 27587 4006 27605
rect 3972 27537 4006 27549
rect 3972 27515 4006 27537
rect 3972 27469 4006 27477
rect 3972 27443 4006 27469
rect 3972 27401 4006 27405
rect 3972 27371 4006 27401
rect 3972 27299 4006 27333
rect 3972 27231 4006 27261
rect 3972 27227 4006 27231
rect 3972 27163 4006 27189
rect 3972 27155 4006 27163
rect 3972 27095 4006 27117
rect 3972 27083 4006 27095
rect 3972 27027 4006 27045
rect 3972 27011 4006 27027
rect 3972 26959 4006 26973
rect 3972 26939 4006 26959
rect 3972 26891 4006 26901
rect 3972 26867 4006 26891
rect 3972 26823 4006 26829
rect 3972 26795 4006 26823
rect 3972 26755 4006 26757
rect 3972 26723 4006 26755
rect 3972 26653 4006 26685
rect 3972 26651 4006 26653
rect 3972 26585 4006 26613
rect 3972 26579 4006 26585
rect 3972 26517 4006 26541
rect 3972 26507 4006 26517
rect 3972 26449 4006 26469
rect 3972 26435 4006 26449
rect 3972 26381 4006 26397
rect 3972 26363 4006 26381
rect 3972 26313 4006 26325
rect 3972 26291 4006 26313
rect 3972 26245 4006 26253
rect 3972 26219 4006 26245
rect 3972 26177 4006 26181
rect 3972 26147 4006 26177
rect 3972 26075 4006 26109
rect 3972 26007 4006 26037
rect 3972 26003 4006 26007
rect 3972 25939 4006 25965
rect 3972 25931 4006 25939
rect 3972 25871 4006 25893
rect 3972 25859 4006 25871
rect 3972 25803 4006 25821
rect 3972 25787 4006 25803
rect 3972 25735 4006 25749
rect 3972 25715 4006 25735
rect 3972 25667 4006 25677
rect 3972 25643 4006 25667
rect 3972 25599 4006 25605
rect 3972 25571 4006 25599
rect 3972 25531 4006 25533
rect 3972 25499 4006 25531
rect 3972 25429 4006 25461
rect 3972 25427 4006 25429
rect 3972 25361 4006 25389
rect 3972 25355 4006 25361
rect 3972 25293 4006 25317
rect 3972 25283 4006 25293
rect 3972 25225 4006 25245
rect 3972 25211 4006 25225
rect 3972 25157 4006 25173
rect 3972 25139 4006 25157
rect 3972 25089 4006 25101
rect 3972 25067 4006 25089
rect 3972 25021 4006 25029
rect 3972 24995 4006 25021
rect 3972 24953 4006 24957
rect 3972 24923 4006 24953
rect 3972 24851 4006 24885
rect 3972 24783 4006 24813
rect 3972 24779 4006 24783
rect 3972 24715 4006 24741
rect 3972 24707 4006 24715
rect 3972 24647 4006 24669
rect 3972 24635 4006 24647
rect 3972 24579 4006 24597
rect 3972 24563 4006 24579
rect 3972 24511 4006 24525
rect 3972 24491 4006 24511
rect 3972 24443 4006 24453
rect 3972 24419 4006 24443
rect 3972 24375 4006 24381
rect 3972 24347 4006 24375
rect 3972 24307 4006 24309
rect 3972 24275 4006 24307
rect 3972 24205 4006 24237
rect 3972 24203 4006 24205
rect 3972 24137 4006 24165
rect 3972 24131 4006 24137
rect 3972 24069 4006 24093
rect 3972 24059 4006 24069
rect 3972 24001 4006 24021
rect 3972 23987 4006 24001
rect 3972 23933 4006 23949
rect 3972 23915 4006 23933
rect 3972 23865 4006 23877
rect 3972 23843 4006 23865
rect 3972 23797 4006 23805
rect 3972 23771 4006 23797
rect 3972 23729 4006 23733
rect 3972 23699 4006 23729
rect 3972 23627 4006 23661
rect 3972 23559 4006 23589
rect 3972 23555 4006 23559
rect 3972 23491 4006 23517
rect 3972 23483 4006 23491
rect 3972 23423 4006 23445
rect 3972 23411 4006 23423
rect 3972 23355 4006 23373
rect 3972 23339 4006 23355
rect 3972 23287 4006 23301
rect 3972 23267 4006 23287
rect 3972 23219 4006 23229
rect 3972 23195 4006 23219
rect 3972 23151 4006 23157
rect 3972 23123 4006 23151
rect 3972 23083 4006 23085
rect 3972 23051 4006 23083
rect 3972 22981 4006 23013
rect 3972 22979 4006 22981
rect 3972 22913 4006 22941
rect 3972 22907 4006 22913
rect 3972 22845 4006 22869
rect 3972 22835 4006 22845
rect 3972 22777 4006 22797
rect 3972 22763 4006 22777
rect 3972 22709 4006 22725
rect 3972 22691 4006 22709
rect 3972 22641 4006 22653
rect 3972 22619 4006 22641
rect 3972 22573 4006 22581
rect 3972 22547 4006 22573
rect 3972 22505 4006 22509
rect 3972 22475 4006 22505
rect 3972 22403 4006 22437
rect 3972 22335 4006 22365
rect 3972 22331 4006 22335
rect 3972 22267 4006 22293
rect 3972 22259 4006 22267
rect 3972 22199 4006 22221
rect 3972 22187 4006 22199
rect 3972 22131 4006 22149
rect 3972 22115 4006 22131
rect 3972 22063 4006 22077
rect 3972 22043 4006 22063
rect 3972 21995 4006 22005
rect 3972 21971 4006 21995
rect 3972 21927 4006 21933
rect 3972 21899 4006 21927
rect 3972 21859 4006 21861
rect 3972 21827 4006 21859
rect 3972 21757 4006 21789
rect 3972 21755 4006 21757
rect 3972 21689 4006 21717
rect 3972 21683 4006 21689
rect 3972 21621 4006 21645
rect 3972 21611 4006 21621
rect 3972 21553 4006 21573
rect 3972 21539 4006 21553
rect 3972 21485 4006 21501
rect 3972 21467 4006 21485
rect 3972 21417 4006 21429
rect 3972 21395 4006 21417
rect 3972 21349 4006 21357
rect 3972 21323 4006 21349
rect 3972 21281 4006 21285
rect 3972 21251 4006 21281
rect 3972 21179 4006 21213
rect 3972 21111 4006 21141
rect 3972 21107 4006 21111
rect 3972 21043 4006 21069
rect 3972 21035 4006 21043
rect 3972 20975 4006 20997
rect 3972 20963 4006 20975
rect 3972 20907 4006 20925
rect 3972 20891 4006 20907
rect 3972 20839 4006 20853
rect 3972 20819 4006 20839
rect 3972 20771 4006 20781
rect 3972 20747 4006 20771
rect 3972 20703 4006 20709
rect 3972 20675 4006 20703
rect 3972 20635 4006 20637
rect 3972 20603 4006 20635
rect 3972 20533 4006 20565
rect 3972 20531 4006 20533
rect 3972 20465 4006 20493
rect 3972 20459 4006 20465
rect 3972 20397 4006 20421
rect 3972 20387 4006 20397
rect 3972 20329 4006 20349
rect 3972 20315 4006 20329
rect 3972 20261 4006 20277
rect 3972 20243 4006 20261
rect 3972 20193 4006 20205
rect 3972 20171 4006 20193
rect 3972 20125 4006 20133
rect 3972 20099 4006 20125
rect 3972 20057 4006 20061
rect 3972 20027 4006 20057
rect 3972 19955 4006 19989
rect 3972 19887 4006 19917
rect 3972 19883 4006 19887
rect 3972 19819 4006 19845
rect 3972 19811 4006 19819
rect 3972 19751 4006 19773
rect 3972 19739 4006 19751
rect 3972 19683 4006 19701
rect 3972 19667 4006 19683
rect 3972 19615 4006 19629
rect 3972 19595 4006 19615
rect 3972 19547 4006 19557
rect 3972 19523 4006 19547
rect 3972 19479 4006 19485
rect 3972 19451 4006 19479
rect 3972 19411 4006 19413
rect 3972 19379 4006 19411
rect 3972 19309 4006 19341
rect 3972 19307 4006 19309
rect 3972 19241 4006 19269
rect 3972 19235 4006 19241
rect 3972 19173 4006 19197
rect 3972 19163 4006 19173
rect 3972 19105 4006 19125
rect 3972 19091 4006 19105
rect 3972 19037 4006 19053
rect 3972 19019 4006 19037
rect 3972 18969 4006 18981
rect 3972 18947 4006 18969
rect 3972 18901 4006 18909
rect 3972 18875 4006 18901
rect 3972 18833 4006 18837
rect 3972 18803 4006 18833
rect 3972 18731 4006 18765
rect 3972 18663 4006 18693
rect 3972 18659 4006 18663
rect 3972 18595 4006 18621
rect 3972 18587 4006 18595
rect 3972 18527 4006 18549
rect 3972 18515 4006 18527
rect 3972 18459 4006 18477
rect 3972 18443 4006 18459
rect 3972 18391 4006 18405
rect 3972 18371 4006 18391
rect 3972 18323 4006 18333
rect 3972 18299 4006 18323
rect 3972 18255 4006 18261
rect 3972 18227 4006 18255
rect 3972 18187 4006 18189
rect 3972 18155 4006 18187
rect 3972 18085 4006 18117
rect 3972 18083 4006 18085
rect 3972 18017 4006 18045
rect 3972 18011 4006 18017
rect 3972 17949 4006 17973
rect 3972 17939 4006 17949
rect 3972 17881 4006 17901
rect 3972 17867 4006 17881
rect 3972 17813 4006 17829
rect 3972 17795 4006 17813
rect 3972 17745 4006 17757
rect 3972 17723 4006 17745
rect 3972 17677 4006 17685
rect 3972 17651 4006 17677
rect 3972 17609 4006 17613
rect 3972 17579 4006 17609
rect 3972 17507 4006 17541
rect 3972 17439 4006 17469
rect 3972 17435 4006 17439
rect 3972 17371 4006 17397
rect 3972 17363 4006 17371
rect 3972 17303 4006 17325
rect 3972 17291 4006 17303
rect 3972 17235 4006 17253
rect 3972 17219 4006 17235
rect 3972 17167 4006 17181
rect 3972 17147 4006 17167
rect 3972 17099 4006 17109
rect 3972 17075 4006 17099
rect 3972 17031 4006 17037
rect 3972 17003 4006 17031
rect 3972 16963 4006 16965
rect 3972 16931 4006 16963
rect 3972 16861 4006 16893
rect 3972 16859 4006 16861
rect 3972 16793 4006 16821
rect 3972 16787 4006 16793
rect 3972 16725 4006 16749
rect 3972 16715 4006 16725
rect 3972 16657 4006 16677
rect 3972 16643 4006 16657
rect 3972 16589 4006 16605
rect 3972 16571 4006 16589
rect 3972 16521 4006 16533
rect 3972 16499 4006 16521
rect 3972 16453 4006 16461
rect 3972 16427 4006 16453
rect 3972 16385 4006 16389
rect 3972 16355 4006 16385
rect 3972 16283 4006 16317
rect 3972 16215 4006 16245
rect 3972 16211 4006 16215
rect 3972 16147 4006 16173
rect 3972 16139 4006 16147
rect 3972 16079 4006 16101
rect 3972 16067 4006 16079
rect 3972 16011 4006 16029
rect 3972 15995 4006 16011
rect 3972 15943 4006 15957
rect 3972 15923 4006 15943
rect 3972 15875 4006 15885
rect 3972 15851 4006 15875
rect 3972 15807 4006 15813
rect 3972 15779 4006 15807
rect 3972 15739 4006 15741
rect 3972 15707 4006 15739
rect 3972 15637 4006 15669
rect 3972 15635 4006 15637
rect 3972 15569 4006 15597
rect 3972 15563 4006 15569
rect 3972 15501 4006 15525
rect 3972 15491 4006 15501
rect 3972 15433 4006 15453
rect 3972 15419 4006 15433
rect 3972 15365 4006 15381
rect 3972 15347 4006 15365
rect 3972 15297 4006 15309
rect 3972 15275 4006 15297
rect 3972 15229 4006 15237
rect 3972 15203 4006 15229
rect 3972 15161 4006 15165
rect 3972 15131 4006 15161
rect 3972 15059 4006 15093
rect 3972 14991 4006 15021
rect 3972 14987 4006 14991
rect 3972 14923 4006 14949
rect 3972 14915 4006 14923
rect 3972 14855 4006 14877
rect 3972 14843 4006 14855
rect 3972 14787 4006 14805
rect 3972 14771 4006 14787
rect 3972 14719 4006 14733
rect 3972 14699 4006 14719
rect 3972 14651 4006 14661
rect 3972 14627 4006 14651
rect 3972 14583 4006 14589
rect 3972 14555 4006 14583
rect 3972 14515 4006 14517
rect 3972 14483 4006 14515
rect 3972 14413 4006 14445
rect 3972 14411 4006 14413
rect 3972 14345 4006 14373
rect 3972 14339 4006 14345
rect 3972 14277 4006 14301
rect 3972 14267 4006 14277
rect 3972 14209 4006 14229
rect 3972 14195 4006 14209
rect 3972 14141 4006 14157
rect 3972 14123 4006 14141
rect 3972 14073 4006 14085
rect 3972 14051 4006 14073
rect 3972 14005 4006 14013
rect 3972 13979 4006 14005
rect 3972 13937 4006 13941
rect 3972 13907 4006 13937
rect 3972 13835 4006 13869
rect 3972 13767 4006 13797
rect 3972 13763 4006 13767
rect 3972 13699 4006 13725
rect 3972 13691 4006 13699
rect 3972 13631 4006 13653
rect 3972 13619 4006 13631
rect 3972 13563 4006 13581
rect 3972 13547 4006 13563
rect 3972 13495 4006 13509
rect 3972 13475 4006 13495
rect 3972 13427 4006 13437
rect 3972 13403 4006 13427
rect 3972 13359 4006 13365
rect 3972 13331 4006 13359
rect 3972 13291 4006 13293
rect 3972 13259 4006 13291
rect 3972 13189 4006 13221
rect 3972 13187 4006 13189
rect 3972 13121 4006 13149
rect 3972 13115 4006 13121
rect 3972 13053 4006 13077
rect 3972 13043 4006 13053
rect 3972 12985 4006 13005
rect 3972 12971 4006 12985
rect 3972 12917 4006 12933
rect 3972 12899 4006 12917
rect 3972 12849 4006 12861
rect 3972 12827 4006 12849
rect 3972 12781 4006 12789
rect 3972 12755 4006 12781
rect 3972 12713 4006 12717
rect 3972 12683 4006 12713
rect 3972 12611 4006 12645
rect 3972 12543 4006 12573
rect 3972 12539 4006 12543
rect 3972 12475 4006 12501
rect 3972 12467 4006 12475
rect 3972 12407 4006 12429
rect 3972 12395 4006 12407
rect 3972 12339 4006 12357
rect 3972 12323 4006 12339
rect 3972 12271 4006 12285
rect 3972 12251 4006 12271
rect 3972 12203 4006 12213
rect 3972 12179 4006 12203
rect 3972 12135 4006 12141
rect 3972 12107 4006 12135
rect 3972 12067 4006 12069
rect 3972 12035 4006 12067
rect 3972 11965 4006 11997
rect 3972 11963 4006 11965
rect 3972 11897 4006 11925
rect 3972 11891 4006 11897
rect 3972 11829 4006 11853
rect 3972 11819 4006 11829
rect 3972 11761 4006 11781
rect 3972 11747 4006 11761
rect 3972 11693 4006 11709
rect 3972 11675 4006 11693
rect 3972 11625 4006 11637
rect 3972 11603 4006 11625
rect 3972 11557 4006 11565
rect 3972 11531 4006 11557
rect 3972 11489 4006 11493
rect 3972 11459 4006 11489
rect 3972 11387 4006 11421
rect 3972 11319 4006 11349
rect 3972 11315 4006 11319
rect 3972 11251 4006 11277
rect 3972 11243 4006 11251
rect 3972 11183 4006 11205
rect 3972 11171 4006 11183
rect 3972 11115 4006 11133
rect 3972 11099 4006 11115
rect 3972 11047 4006 11061
rect 3972 11027 4006 11047
rect 3972 10979 4006 10989
rect 3972 10955 4006 10979
rect 3972 10911 4006 10917
rect 3972 10883 4006 10911
rect 3972 10843 4006 10845
rect 3972 10811 4006 10843
rect 3972 10741 4006 10773
rect 3972 10739 4006 10741
rect 3972 10673 4006 10701
rect 3972 10667 4006 10673
rect 3972 10605 4006 10629
rect 3972 10595 4006 10605
rect 3972 10537 4006 10557
rect 3972 10523 4006 10537
rect 3972 10469 4006 10485
rect 3972 10451 4006 10469
rect 3972 10401 4006 10413
rect 3972 10379 4006 10401
rect 3972 10333 4006 10341
rect 3972 10307 4006 10333
rect 3972 10265 4006 10269
rect 3972 10235 4006 10265
rect 3972 10163 4006 10197
rect 3972 10095 4006 10125
rect 3972 10091 4006 10095
rect 3972 10027 4006 10053
rect 3972 10019 4006 10027
rect 3972 9959 4006 9981
rect 3972 9947 4006 9959
rect 3972 9891 4006 9909
rect 3972 9875 4006 9891
rect 3972 9823 4006 9837
rect 3972 9803 4006 9823
rect 3972 9755 4006 9765
rect 3972 9731 4006 9755
rect 3972 9687 4006 9693
rect 3972 9659 4006 9687
rect 3972 9619 4006 9621
rect 3972 9587 4006 9619
rect 3972 9517 4006 9549
rect 3972 9515 4006 9517
rect 3972 9449 4006 9477
rect 3972 9443 4006 9449
rect 3972 9381 4006 9405
rect 3972 9371 4006 9381
rect 3972 9313 4006 9333
rect 3972 9299 4006 9313
rect 3972 9245 4006 9261
rect 3972 9227 4006 9245
rect 3972 9177 4006 9189
rect 3972 9155 4006 9177
rect 3972 9109 4006 9117
rect 3972 9083 4006 9109
rect 3972 9041 4006 9045
rect 3972 9011 4006 9041
rect 3972 8939 4006 8973
rect 3972 8871 4006 8901
rect 3972 8867 4006 8871
rect 3972 8803 4006 8829
rect 3972 8795 4006 8803
rect 3972 8735 4006 8757
rect 3972 8723 4006 8735
rect 3972 8667 4006 8685
rect 3972 8651 4006 8667
rect 3972 8599 4006 8613
rect 3972 8579 4006 8599
rect 3972 8531 4006 8541
rect 3972 8507 4006 8531
rect 3972 8463 4006 8469
rect 3972 8435 4006 8463
rect 3972 8395 4006 8397
rect 3972 8363 4006 8395
rect 3972 8293 4006 8325
rect 3972 8291 4006 8293
rect 3972 8225 4006 8253
rect 3972 8219 4006 8225
rect 3972 8157 4006 8181
rect 3972 8147 4006 8157
rect 3972 8089 4006 8109
rect 3972 8075 4006 8089
rect 3972 8021 4006 8037
rect 3972 8003 4006 8021
rect 3972 7953 4006 7965
rect 3972 7931 4006 7953
rect 3972 7885 4006 7893
rect 3972 7859 4006 7885
rect 3972 7817 4006 7821
rect 3972 7787 4006 7817
rect 3972 7715 4006 7749
rect 3972 7647 4006 7677
rect 3972 7643 4006 7647
rect 3972 7579 4006 7605
rect 3972 7571 4006 7579
rect 3972 7511 4006 7533
rect 3972 7499 4006 7511
rect 3972 7443 4006 7461
rect 3972 7427 4006 7443
rect 3972 7375 4006 7389
rect 3972 7355 4006 7375
rect 3972 7307 4006 7317
rect 3972 7283 4006 7307
rect 3972 7239 4006 7245
rect 3972 7211 4006 7239
rect 3972 7171 4006 7173
rect 3972 7139 4006 7171
rect 3972 7069 4006 7101
rect 3972 7067 4006 7069
rect 3972 7001 4006 7029
rect 3972 6995 4006 7001
rect 3972 6933 4006 6957
rect 3972 6923 4006 6933
rect 3972 6865 4006 6885
rect 3972 6851 4006 6865
rect 3972 6797 4006 6813
rect 3972 6779 4006 6797
rect 3972 6729 4006 6741
rect 3972 6707 4006 6729
rect 3972 6661 4006 6669
rect 3972 6635 4006 6661
rect 3972 6593 4006 6597
rect 3972 6563 4006 6593
rect 3972 6491 4006 6525
rect 3972 6423 4006 6453
rect 3972 6419 4006 6423
rect 3972 6355 4006 6381
rect 3972 6347 4006 6355
rect 3972 6287 4006 6309
rect 3972 6275 4006 6287
rect 3972 6219 4006 6237
rect 3972 6203 4006 6219
rect 3972 6151 4006 6165
rect 3972 6131 4006 6151
rect 3972 6083 4006 6093
rect 3972 6059 4006 6083
rect 3972 6015 4006 6021
rect 3972 5987 4006 6015
rect 3972 5947 4006 5949
rect 3972 5915 4006 5947
rect 3972 5845 4006 5877
rect 3972 5843 4006 5845
rect 3972 5777 4006 5805
rect 3972 5771 4006 5777
rect 3972 5709 4006 5733
rect 3972 5699 4006 5709
rect 3972 5641 4006 5661
rect 3972 5627 4006 5641
rect 3972 5573 4006 5589
rect 3972 5555 4006 5573
rect 3972 5505 4006 5517
rect 3972 5483 4006 5505
rect 3972 5437 4006 5445
rect 3972 5411 4006 5437
rect 3972 5369 4006 5373
rect 3972 5339 4006 5369
rect 3972 5267 4006 5301
rect 3972 5199 4006 5229
rect 3972 5195 4006 5199
rect 3972 5131 4006 5157
rect 3972 5123 4006 5131
rect 3972 5063 4006 5085
rect 3972 5051 4006 5063
rect 3972 4995 4006 5013
rect 3972 4979 4006 4995
rect 3972 4927 4006 4941
rect 3972 4907 4006 4927
rect 3972 4859 4006 4869
rect 3972 4835 4006 4859
rect 3972 4791 4006 4797
rect 3972 4763 4006 4791
rect 3972 4723 4006 4725
rect 3972 4691 4006 4723
rect 3972 4621 4006 4653
rect 3972 4619 4006 4621
rect 3972 4553 4006 4581
rect 3972 4547 4006 4553
rect 3972 4485 4006 4509
rect 3972 4475 4006 4485
rect 3972 4417 4006 4437
rect 3972 4403 4006 4417
rect 3972 4349 4006 4365
rect 3972 4331 4006 4349
rect 3972 4281 4006 4293
rect 3972 4259 4006 4281
rect 3972 4213 4006 4221
rect 3972 4187 4006 4213
rect 3972 4145 4006 4149
rect 3972 4115 4006 4145
rect 3972 4043 4006 4077
rect 3972 3975 4006 4005
rect 3972 3971 4006 3975
rect 3972 3907 4006 3933
rect 3972 3899 4006 3907
rect 3972 3839 4006 3861
rect 3972 3827 4006 3839
rect 3972 3771 4006 3789
rect 3972 3755 4006 3771
rect 3972 3703 4006 3717
rect 3972 3683 4006 3703
rect 3972 3635 4006 3645
rect 3972 3611 4006 3635
rect 3972 3567 4006 3573
rect 3972 3539 4006 3567
rect 1830 3417 1864 3429
rect 1830 3395 1864 3417
rect -252 3329 -218 3357
rect -252 3323 -218 3329
rect -252 3251 -218 3285
rect 2016 3452 2050 3486
rect 2016 3394 2050 3414
rect 2016 3380 2050 3394
rect 2134 3452 2168 3486
rect 2134 3394 2168 3414
rect 2134 3380 2168 3394
rect 2252 3452 2286 3486
rect 2252 3394 2286 3414
rect 2252 3380 2286 3394
rect 2370 3452 2404 3486
rect 2370 3394 2404 3414
rect 2370 3380 2404 3394
rect 2488 3452 2522 3486
rect 2488 3394 2522 3414
rect 2488 3380 2522 3394
rect 2606 3452 2640 3486
rect 2606 3394 2640 3414
rect 2606 3380 2640 3394
rect 2724 3452 2758 3486
rect 2724 3394 2758 3414
rect 2724 3380 2758 3394
rect 2842 3452 2876 3486
rect 2842 3394 2876 3414
rect 2842 3380 2876 3394
rect 2960 3452 2994 3486
rect 2960 3394 2994 3414
rect 2960 3380 2994 3394
rect 3078 3452 3112 3486
rect 3078 3394 3112 3414
rect 3078 3380 3112 3394
rect 3196 3452 3230 3486
rect 3196 3394 3230 3414
rect 3196 3380 3230 3394
rect 3314 3452 3348 3486
rect 3314 3394 3348 3414
rect 3314 3380 3348 3394
rect 3432 3452 3466 3486
rect 3432 3394 3466 3414
rect 3432 3380 3466 3394
rect 3550 3452 3584 3486
rect 3550 3394 3584 3414
rect 3550 3380 3584 3394
rect 3668 3452 3702 3486
rect 3668 3394 3702 3414
rect 3668 3380 3702 3394
rect 3786 3452 3820 3486
rect 3786 3394 3820 3414
rect 3786 3380 3820 3394
rect 3972 3499 4006 3501
rect 3972 3467 4006 3499
rect 6114 38651 6148 38685
rect 6114 38607 6148 38613
rect 6114 38579 6148 38607
rect 6114 38539 6148 38541
rect 6114 38507 6148 38539
rect 6114 38437 6148 38469
rect 6114 38435 6148 38437
rect 6114 38369 6148 38397
rect 6114 38363 6148 38369
rect 6114 38301 6148 38325
rect 6114 38291 6148 38301
rect 6114 38233 6148 38253
rect 6114 38219 6148 38233
rect 6114 38165 6148 38181
rect 6114 38147 6148 38165
rect 6114 38097 6148 38109
rect 6114 38075 6148 38097
rect 6114 38029 6148 38037
rect 6114 38003 6148 38029
rect 6114 37961 6148 37965
rect 6114 37931 6148 37961
rect 6114 37859 6148 37893
rect 6114 37791 6148 37821
rect 6114 37787 6148 37791
rect 6114 37723 6148 37749
rect 6114 37715 6148 37723
rect 6114 37655 6148 37677
rect 6114 37643 6148 37655
rect 6114 37587 6148 37605
rect 6114 37571 6148 37587
rect 6114 37519 6148 37533
rect 6114 37499 6148 37519
rect 6114 37451 6148 37461
rect 6114 37427 6148 37451
rect 6114 37383 6148 37389
rect 6114 37355 6148 37383
rect 6114 37315 6148 37317
rect 6114 37283 6148 37315
rect 6114 37213 6148 37245
rect 6114 37211 6148 37213
rect 6114 37145 6148 37173
rect 6114 37139 6148 37145
rect 6114 37077 6148 37101
rect 6114 37067 6148 37077
rect 6114 37009 6148 37029
rect 6114 36995 6148 37009
rect 6114 36941 6148 36957
rect 6114 36923 6148 36941
rect 6114 36873 6148 36885
rect 6114 36851 6148 36873
rect 6114 36805 6148 36813
rect 6114 36779 6148 36805
rect 6114 36737 6148 36741
rect 6114 36707 6148 36737
rect 6114 36635 6148 36669
rect 6114 36567 6148 36597
rect 6114 36563 6148 36567
rect 6114 36499 6148 36525
rect 6114 36491 6148 36499
rect 6114 36431 6148 36453
rect 6114 36419 6148 36431
rect 6114 36363 6148 36381
rect 6114 36347 6148 36363
rect 6114 36295 6148 36309
rect 6114 36275 6148 36295
rect 6114 36227 6148 36237
rect 6114 36203 6148 36227
rect 6114 36159 6148 36165
rect 6114 36131 6148 36159
rect 6114 36091 6148 36093
rect 6114 36059 6148 36091
rect 6114 35989 6148 36021
rect 6114 35987 6148 35989
rect 6114 35921 6148 35949
rect 6114 35915 6148 35921
rect 6114 35853 6148 35877
rect 6114 35843 6148 35853
rect 6114 35785 6148 35805
rect 6114 35771 6148 35785
rect 6114 35717 6148 35733
rect 6114 35699 6148 35717
rect 6114 35649 6148 35661
rect 6114 35627 6148 35649
rect 6114 35581 6148 35589
rect 6114 35555 6148 35581
rect 6114 35513 6148 35517
rect 6114 35483 6148 35513
rect 6114 35411 6148 35445
rect 6114 35343 6148 35373
rect 6114 35339 6148 35343
rect 6114 35275 6148 35301
rect 6114 35267 6148 35275
rect 6114 35207 6148 35229
rect 6114 35195 6148 35207
rect 6114 35139 6148 35157
rect 6114 35123 6148 35139
rect 6114 35071 6148 35085
rect 6114 35051 6148 35071
rect 6114 35003 6148 35013
rect 6114 34979 6148 35003
rect 6114 34935 6148 34941
rect 6114 34907 6148 34935
rect 6114 34867 6148 34869
rect 6114 34835 6148 34867
rect 6114 34765 6148 34797
rect 6114 34763 6148 34765
rect 6114 34697 6148 34725
rect 6114 34691 6148 34697
rect 6114 34629 6148 34653
rect 6114 34619 6148 34629
rect 6114 34561 6148 34581
rect 6114 34547 6148 34561
rect 6114 34493 6148 34509
rect 6114 34475 6148 34493
rect 6114 34425 6148 34437
rect 6114 34403 6148 34425
rect 6114 34357 6148 34365
rect 6114 34331 6148 34357
rect 6114 34289 6148 34293
rect 6114 34259 6148 34289
rect 6114 34187 6148 34221
rect 6114 34119 6148 34149
rect 6114 34115 6148 34119
rect 6114 34051 6148 34077
rect 6114 34043 6148 34051
rect 6114 33983 6148 34005
rect 6114 33971 6148 33983
rect 6114 33915 6148 33933
rect 6114 33899 6148 33915
rect 6114 33847 6148 33861
rect 6114 33827 6148 33847
rect 6114 33779 6148 33789
rect 6114 33755 6148 33779
rect 6114 33711 6148 33717
rect 6114 33683 6148 33711
rect 6114 33643 6148 33645
rect 6114 33611 6148 33643
rect 6114 33541 6148 33573
rect 6114 33539 6148 33541
rect 6114 33473 6148 33501
rect 6114 33467 6148 33473
rect 6114 33405 6148 33429
rect 6114 33395 6148 33405
rect 6114 33337 6148 33357
rect 6114 33323 6148 33337
rect 6114 33269 6148 33285
rect 6114 33251 6148 33269
rect 6114 33201 6148 33213
rect 6114 33179 6148 33201
rect 6114 33133 6148 33141
rect 6114 33107 6148 33133
rect 6114 33065 6148 33069
rect 6114 33035 6148 33065
rect 6114 32963 6148 32997
rect 6114 32895 6148 32925
rect 6114 32891 6148 32895
rect 6114 32827 6148 32853
rect 6114 32819 6148 32827
rect 6114 32759 6148 32781
rect 6114 32747 6148 32759
rect 6114 32691 6148 32709
rect 6114 32675 6148 32691
rect 6114 32623 6148 32637
rect 6114 32603 6148 32623
rect 6114 32555 6148 32565
rect 6114 32531 6148 32555
rect 6114 32487 6148 32493
rect 6114 32459 6148 32487
rect 6114 32419 6148 32421
rect 6114 32387 6148 32419
rect 6114 32317 6148 32349
rect 6114 32315 6148 32317
rect 6114 32249 6148 32277
rect 6114 32243 6148 32249
rect 6114 32181 6148 32205
rect 6114 32171 6148 32181
rect 6114 32113 6148 32133
rect 6114 32099 6148 32113
rect 6114 32045 6148 32061
rect 6114 32027 6148 32045
rect 6114 31977 6148 31989
rect 6114 31955 6148 31977
rect 6114 31909 6148 31917
rect 6114 31883 6148 31909
rect 6114 31841 6148 31845
rect 6114 31811 6148 31841
rect 6114 31739 6148 31773
rect 6114 31671 6148 31701
rect 6114 31667 6148 31671
rect 6114 31603 6148 31629
rect 6114 31595 6148 31603
rect 6114 31535 6148 31557
rect 6114 31523 6148 31535
rect 6114 31467 6148 31485
rect 6114 31451 6148 31467
rect 6114 31399 6148 31413
rect 6114 31379 6148 31399
rect 6114 31331 6148 31341
rect 6114 31307 6148 31331
rect 6114 31263 6148 31269
rect 6114 31235 6148 31263
rect 6114 31195 6148 31197
rect 6114 31163 6148 31195
rect 6114 31093 6148 31125
rect 6114 31091 6148 31093
rect 6114 31025 6148 31053
rect 6114 31019 6148 31025
rect 6114 30957 6148 30981
rect 6114 30947 6148 30957
rect 6114 30889 6148 30909
rect 6114 30875 6148 30889
rect 6114 30821 6148 30837
rect 6114 30803 6148 30821
rect 6114 30753 6148 30765
rect 6114 30731 6148 30753
rect 6114 30685 6148 30693
rect 6114 30659 6148 30685
rect 6114 30617 6148 30621
rect 6114 30587 6148 30617
rect 6114 30515 6148 30549
rect 6114 30447 6148 30477
rect 6114 30443 6148 30447
rect 6114 30379 6148 30405
rect 6114 30371 6148 30379
rect 6114 30311 6148 30333
rect 6114 30299 6148 30311
rect 6114 30243 6148 30261
rect 6114 30227 6148 30243
rect 6114 30175 6148 30189
rect 6114 30155 6148 30175
rect 6114 30107 6148 30117
rect 6114 30083 6148 30107
rect 6114 30039 6148 30045
rect 6114 30011 6148 30039
rect 6114 29971 6148 29973
rect 6114 29939 6148 29971
rect 6114 29869 6148 29901
rect 6114 29867 6148 29869
rect 6114 29801 6148 29829
rect 6114 29795 6148 29801
rect 6114 29733 6148 29757
rect 6114 29723 6148 29733
rect 6114 29665 6148 29685
rect 6114 29651 6148 29665
rect 6114 29597 6148 29613
rect 6114 29579 6148 29597
rect 6114 29529 6148 29541
rect 6114 29507 6148 29529
rect 6114 29461 6148 29469
rect 6114 29435 6148 29461
rect 6114 29393 6148 29397
rect 6114 29363 6148 29393
rect 6114 29291 6148 29325
rect 6114 29223 6148 29253
rect 6114 29219 6148 29223
rect 6114 29155 6148 29181
rect 6114 29147 6148 29155
rect 6114 29087 6148 29109
rect 6114 29075 6148 29087
rect 6114 29019 6148 29037
rect 6114 29003 6148 29019
rect 6114 28951 6148 28965
rect 6114 28931 6148 28951
rect 6114 28883 6148 28893
rect 6114 28859 6148 28883
rect 6114 28815 6148 28821
rect 6114 28787 6148 28815
rect 6114 28747 6148 28749
rect 6114 28715 6148 28747
rect 6114 28645 6148 28677
rect 6114 28643 6148 28645
rect 6114 28577 6148 28605
rect 6114 28571 6148 28577
rect 6114 28509 6148 28533
rect 6114 28499 6148 28509
rect 6114 28441 6148 28461
rect 6114 28427 6148 28441
rect 6114 28373 6148 28389
rect 6114 28355 6148 28373
rect 6114 28305 6148 28317
rect 6114 28283 6148 28305
rect 6114 28237 6148 28245
rect 6114 28211 6148 28237
rect 6114 28169 6148 28173
rect 6114 28139 6148 28169
rect 6114 28067 6148 28101
rect 6114 27999 6148 28029
rect 6114 27995 6148 27999
rect 6114 27931 6148 27957
rect 6114 27923 6148 27931
rect 6114 27863 6148 27885
rect 6114 27851 6148 27863
rect 6114 27795 6148 27813
rect 6114 27779 6148 27795
rect 6114 27727 6148 27741
rect 6114 27707 6148 27727
rect 6114 27659 6148 27669
rect 6114 27635 6148 27659
rect 6114 27591 6148 27597
rect 6114 27563 6148 27591
rect 6114 27523 6148 27525
rect 6114 27491 6148 27523
rect 6114 27421 6148 27453
rect 6114 27419 6148 27421
rect 6114 27353 6148 27381
rect 6114 27347 6148 27353
rect 6114 27285 6148 27309
rect 6114 27275 6148 27285
rect 6114 27217 6148 27237
rect 6114 27203 6148 27217
rect 6114 27149 6148 27165
rect 6114 27131 6148 27149
rect 6114 27081 6148 27093
rect 6114 27059 6148 27081
rect 6114 27013 6148 27021
rect 6114 26987 6148 27013
rect 6114 26945 6148 26949
rect 6114 26915 6148 26945
rect 6114 26843 6148 26877
rect 6114 26775 6148 26805
rect 6114 26771 6148 26775
rect 6114 26707 6148 26733
rect 6114 26699 6148 26707
rect 6114 26639 6148 26661
rect 6114 26627 6148 26639
rect 6114 26571 6148 26589
rect 6114 26555 6148 26571
rect 6114 26503 6148 26517
rect 6114 26483 6148 26503
rect 6114 26435 6148 26445
rect 6114 26411 6148 26435
rect 6114 26367 6148 26373
rect 6114 26339 6148 26367
rect 6114 26299 6148 26301
rect 6114 26267 6148 26299
rect 6114 26197 6148 26229
rect 6114 26195 6148 26197
rect 6114 26129 6148 26157
rect 6114 26123 6148 26129
rect 6114 26061 6148 26085
rect 6114 26051 6148 26061
rect 6114 25993 6148 26013
rect 6114 25979 6148 25993
rect 6114 25925 6148 25941
rect 6114 25907 6148 25925
rect 6114 25857 6148 25869
rect 6114 25835 6148 25857
rect 6114 25789 6148 25797
rect 6114 25763 6148 25789
rect 6114 25721 6148 25725
rect 6114 25691 6148 25721
rect 6114 25619 6148 25653
rect 6114 25551 6148 25581
rect 6114 25547 6148 25551
rect 6114 25483 6148 25509
rect 6114 25475 6148 25483
rect 6114 25415 6148 25437
rect 6114 25403 6148 25415
rect 6114 25347 6148 25365
rect 6114 25331 6148 25347
rect 6114 25279 6148 25293
rect 6114 25259 6148 25279
rect 6114 25211 6148 25221
rect 6114 25187 6148 25211
rect 6114 25143 6148 25149
rect 6114 25115 6148 25143
rect 6114 25075 6148 25077
rect 6114 25043 6148 25075
rect 6114 24973 6148 25005
rect 6114 24971 6148 24973
rect 6114 24905 6148 24933
rect 6114 24899 6148 24905
rect 6114 24837 6148 24861
rect 6114 24827 6148 24837
rect 6114 24769 6148 24789
rect 6114 24755 6148 24769
rect 6114 24701 6148 24717
rect 6114 24683 6148 24701
rect 6114 24633 6148 24645
rect 6114 24611 6148 24633
rect 6114 24565 6148 24573
rect 6114 24539 6148 24565
rect 6114 24497 6148 24501
rect 6114 24467 6148 24497
rect 6114 24395 6148 24429
rect 6114 24327 6148 24357
rect 6114 24323 6148 24327
rect 6114 24259 6148 24285
rect 6114 24251 6148 24259
rect 6114 24191 6148 24213
rect 6114 24179 6148 24191
rect 6114 24123 6148 24141
rect 6114 24107 6148 24123
rect 6114 24055 6148 24069
rect 6114 24035 6148 24055
rect 6114 23987 6148 23997
rect 6114 23963 6148 23987
rect 6114 23919 6148 23925
rect 6114 23891 6148 23919
rect 6114 23851 6148 23853
rect 6114 23819 6148 23851
rect 6114 23749 6148 23781
rect 6114 23747 6148 23749
rect 6114 23681 6148 23709
rect 6114 23675 6148 23681
rect 6114 23613 6148 23637
rect 6114 23603 6148 23613
rect 6114 23545 6148 23565
rect 6114 23531 6148 23545
rect 6114 23477 6148 23493
rect 6114 23459 6148 23477
rect 6114 23409 6148 23421
rect 6114 23387 6148 23409
rect 6114 23341 6148 23349
rect 6114 23315 6148 23341
rect 6114 23273 6148 23277
rect 6114 23243 6148 23273
rect 6114 23171 6148 23205
rect 6114 23103 6148 23133
rect 6114 23099 6148 23103
rect 6114 23035 6148 23061
rect 6114 23027 6148 23035
rect 6114 22967 6148 22989
rect 6114 22955 6148 22967
rect 6114 22899 6148 22917
rect 6114 22883 6148 22899
rect 6114 22831 6148 22845
rect 6114 22811 6148 22831
rect 6114 22763 6148 22773
rect 6114 22739 6148 22763
rect 6114 22695 6148 22701
rect 6114 22667 6148 22695
rect 6114 22627 6148 22629
rect 6114 22595 6148 22627
rect 6114 22525 6148 22557
rect 6114 22523 6148 22525
rect 6114 22457 6148 22485
rect 6114 22451 6148 22457
rect 6114 22389 6148 22413
rect 6114 22379 6148 22389
rect 6114 22321 6148 22341
rect 6114 22307 6148 22321
rect 6114 22253 6148 22269
rect 6114 22235 6148 22253
rect 6114 22185 6148 22197
rect 6114 22163 6148 22185
rect 6114 22117 6148 22125
rect 6114 22091 6148 22117
rect 6114 22049 6148 22053
rect 6114 22019 6148 22049
rect 6114 21947 6148 21981
rect 6114 21879 6148 21909
rect 6114 21875 6148 21879
rect 6114 21811 6148 21837
rect 6114 21803 6148 21811
rect 6114 21743 6148 21765
rect 6114 21731 6148 21743
rect 6114 21675 6148 21693
rect 6114 21659 6148 21675
rect 6114 21607 6148 21621
rect 6114 21587 6148 21607
rect 6114 21539 6148 21549
rect 6114 21515 6148 21539
rect 6114 21471 6148 21477
rect 6114 21443 6148 21471
rect 6114 21403 6148 21405
rect 6114 21371 6148 21403
rect 6114 21301 6148 21333
rect 6114 21299 6148 21301
rect 6114 21233 6148 21261
rect 6114 21227 6148 21233
rect 6114 21165 6148 21189
rect 6114 21155 6148 21165
rect 6114 21097 6148 21117
rect 6114 21083 6148 21097
rect 6114 21029 6148 21045
rect 6114 21011 6148 21029
rect 6114 20961 6148 20973
rect 6114 20939 6148 20961
rect 6114 20893 6148 20901
rect 6114 20867 6148 20893
rect 6114 20825 6148 20829
rect 6114 20795 6148 20825
rect 6114 20723 6148 20757
rect 6114 20655 6148 20685
rect 6114 20651 6148 20655
rect 6114 20587 6148 20613
rect 6114 20579 6148 20587
rect 6114 20519 6148 20541
rect 6114 20507 6148 20519
rect 6114 20451 6148 20469
rect 6114 20435 6148 20451
rect 6114 20383 6148 20397
rect 6114 20363 6148 20383
rect 6114 20315 6148 20325
rect 6114 20291 6148 20315
rect 6114 20247 6148 20253
rect 6114 20219 6148 20247
rect 6114 20179 6148 20181
rect 6114 20147 6148 20179
rect 6114 20077 6148 20109
rect 6114 20075 6148 20077
rect 6114 20009 6148 20037
rect 6114 20003 6148 20009
rect 6114 19941 6148 19965
rect 6114 19931 6148 19941
rect 6114 19873 6148 19893
rect 6114 19859 6148 19873
rect 6114 19805 6148 19821
rect 6114 19787 6148 19805
rect 6114 19737 6148 19749
rect 6114 19715 6148 19737
rect 6114 19669 6148 19677
rect 6114 19643 6148 19669
rect 6114 19601 6148 19605
rect 6114 19571 6148 19601
rect 6114 19499 6148 19533
rect 6114 19431 6148 19461
rect 6114 19427 6148 19431
rect 6114 19363 6148 19389
rect 6114 19355 6148 19363
rect 6114 19295 6148 19317
rect 6114 19283 6148 19295
rect 6114 19227 6148 19245
rect 6114 19211 6148 19227
rect 6114 19159 6148 19173
rect 6114 19139 6148 19159
rect 6114 19091 6148 19101
rect 6114 19067 6148 19091
rect 6114 19023 6148 19029
rect 6114 18995 6148 19023
rect 6114 18955 6148 18957
rect 6114 18923 6148 18955
rect 6114 18853 6148 18885
rect 6114 18851 6148 18853
rect 6114 18785 6148 18813
rect 6114 18779 6148 18785
rect 6114 18717 6148 18741
rect 6114 18707 6148 18717
rect 6114 18649 6148 18669
rect 6114 18635 6148 18649
rect 6114 18581 6148 18597
rect 6114 18563 6148 18581
rect 6114 18513 6148 18525
rect 6114 18491 6148 18513
rect 6114 18445 6148 18453
rect 6114 18419 6148 18445
rect 6114 18377 6148 18381
rect 6114 18347 6148 18377
rect 6114 18275 6148 18309
rect 6114 18207 6148 18237
rect 6114 18203 6148 18207
rect 6114 18139 6148 18165
rect 6114 18131 6148 18139
rect 6114 18071 6148 18093
rect 6114 18059 6148 18071
rect 6114 18003 6148 18021
rect 6114 17987 6148 18003
rect 6114 17935 6148 17949
rect 6114 17915 6148 17935
rect 6114 17867 6148 17877
rect 6114 17843 6148 17867
rect 6114 17799 6148 17805
rect 6114 17771 6148 17799
rect 6114 17731 6148 17733
rect 6114 17699 6148 17731
rect 6114 17629 6148 17661
rect 6114 17627 6148 17629
rect 6114 17561 6148 17589
rect 6114 17555 6148 17561
rect 6114 17493 6148 17517
rect 6114 17483 6148 17493
rect 6114 17425 6148 17445
rect 6114 17411 6148 17425
rect 6114 17357 6148 17373
rect 6114 17339 6148 17357
rect 6114 17289 6148 17301
rect 6114 17267 6148 17289
rect 6114 17221 6148 17229
rect 6114 17195 6148 17221
rect 6114 17153 6148 17157
rect 6114 17123 6148 17153
rect 6114 17051 6148 17085
rect 6114 16983 6148 17013
rect 6114 16979 6148 16983
rect 6114 16915 6148 16941
rect 6114 16907 6148 16915
rect 6114 16847 6148 16869
rect 6114 16835 6148 16847
rect 6114 16779 6148 16797
rect 6114 16763 6148 16779
rect 6114 16711 6148 16725
rect 6114 16691 6148 16711
rect 6114 16643 6148 16653
rect 6114 16619 6148 16643
rect 6114 16575 6148 16581
rect 6114 16547 6148 16575
rect 6114 16507 6148 16509
rect 6114 16475 6148 16507
rect 6114 16405 6148 16437
rect 6114 16403 6148 16405
rect 6114 16337 6148 16365
rect 6114 16331 6148 16337
rect 6114 16269 6148 16293
rect 6114 16259 6148 16269
rect 6114 16201 6148 16221
rect 6114 16187 6148 16201
rect 6114 16133 6148 16149
rect 6114 16115 6148 16133
rect 6114 16065 6148 16077
rect 6114 16043 6148 16065
rect 6114 15997 6148 16005
rect 6114 15971 6148 15997
rect 6114 15929 6148 15933
rect 6114 15899 6148 15929
rect 6114 15827 6148 15861
rect 6114 15759 6148 15789
rect 6114 15755 6148 15759
rect 6114 15691 6148 15717
rect 6114 15683 6148 15691
rect 6114 15623 6148 15645
rect 6114 15611 6148 15623
rect 6114 15555 6148 15573
rect 6114 15539 6148 15555
rect 6114 15487 6148 15501
rect 6114 15467 6148 15487
rect 6114 15419 6148 15429
rect 6114 15395 6148 15419
rect 6114 15351 6148 15357
rect 6114 15323 6148 15351
rect 6114 15283 6148 15285
rect 6114 15251 6148 15283
rect 6114 15181 6148 15213
rect 6114 15179 6148 15181
rect 6114 15113 6148 15141
rect 6114 15107 6148 15113
rect 6114 15045 6148 15069
rect 6114 15035 6148 15045
rect 6114 14977 6148 14997
rect 6114 14963 6148 14977
rect 6114 14909 6148 14925
rect 6114 14891 6148 14909
rect 6114 14841 6148 14853
rect 6114 14819 6148 14841
rect 6114 14773 6148 14781
rect 6114 14747 6148 14773
rect 6114 14705 6148 14709
rect 6114 14675 6148 14705
rect 6114 14603 6148 14637
rect 6114 14535 6148 14565
rect 6114 14531 6148 14535
rect 6114 14467 6148 14493
rect 6114 14459 6148 14467
rect 6114 14399 6148 14421
rect 6114 14387 6148 14399
rect 6114 14331 6148 14349
rect 6114 14315 6148 14331
rect 6114 14263 6148 14277
rect 6114 14243 6148 14263
rect 6114 14195 6148 14205
rect 6114 14171 6148 14195
rect 6114 14127 6148 14133
rect 6114 14099 6148 14127
rect 6114 14059 6148 14061
rect 6114 14027 6148 14059
rect 6114 13957 6148 13989
rect 6114 13955 6148 13957
rect 6114 13889 6148 13917
rect 6114 13883 6148 13889
rect 6114 13821 6148 13845
rect 6114 13811 6148 13821
rect 6114 13753 6148 13773
rect 6114 13739 6148 13753
rect 6114 13685 6148 13701
rect 6114 13667 6148 13685
rect 6114 13617 6148 13629
rect 6114 13595 6148 13617
rect 6114 13549 6148 13557
rect 6114 13523 6148 13549
rect 6114 13481 6148 13485
rect 6114 13451 6148 13481
rect 6114 13379 6148 13413
rect 6114 13311 6148 13341
rect 6114 13307 6148 13311
rect 6114 13243 6148 13269
rect 6114 13235 6148 13243
rect 6114 13175 6148 13197
rect 6114 13163 6148 13175
rect 6114 13107 6148 13125
rect 6114 13091 6148 13107
rect 6114 13039 6148 13053
rect 6114 13019 6148 13039
rect 6114 12971 6148 12981
rect 6114 12947 6148 12971
rect 6114 12903 6148 12909
rect 6114 12875 6148 12903
rect 6114 12835 6148 12837
rect 6114 12803 6148 12835
rect 6114 12733 6148 12765
rect 6114 12731 6148 12733
rect 6114 12665 6148 12693
rect 6114 12659 6148 12665
rect 6114 12597 6148 12621
rect 6114 12587 6148 12597
rect 6114 12529 6148 12549
rect 6114 12515 6148 12529
rect 6114 12461 6148 12477
rect 6114 12443 6148 12461
rect 6114 12393 6148 12405
rect 6114 12371 6148 12393
rect 6114 12325 6148 12333
rect 6114 12299 6148 12325
rect 6114 12257 6148 12261
rect 6114 12227 6148 12257
rect 6114 12155 6148 12189
rect 6114 12087 6148 12117
rect 6114 12083 6148 12087
rect 6114 12019 6148 12045
rect 6114 12011 6148 12019
rect 6114 11951 6148 11973
rect 6114 11939 6148 11951
rect 6114 11883 6148 11901
rect 6114 11867 6148 11883
rect 6114 11815 6148 11829
rect 6114 11795 6148 11815
rect 6114 11747 6148 11757
rect 6114 11723 6148 11747
rect 6114 11679 6148 11685
rect 6114 11651 6148 11679
rect 6114 11611 6148 11613
rect 6114 11579 6148 11611
rect 6114 11509 6148 11541
rect 6114 11507 6148 11509
rect 6114 11441 6148 11469
rect 6114 11435 6148 11441
rect 6114 11373 6148 11397
rect 6114 11363 6148 11373
rect 6114 11305 6148 11325
rect 6114 11291 6148 11305
rect 6114 11237 6148 11253
rect 6114 11219 6148 11237
rect 6114 11169 6148 11181
rect 6114 11147 6148 11169
rect 6114 11101 6148 11109
rect 6114 11075 6148 11101
rect 6114 11033 6148 11037
rect 6114 11003 6148 11033
rect 6114 10931 6148 10965
rect 6114 10863 6148 10893
rect 6114 10859 6148 10863
rect 6114 10795 6148 10821
rect 6114 10787 6148 10795
rect 6114 10727 6148 10749
rect 6114 10715 6148 10727
rect 6114 10659 6148 10677
rect 6114 10643 6148 10659
rect 6114 10591 6148 10605
rect 6114 10571 6148 10591
rect 6114 10523 6148 10533
rect 6114 10499 6148 10523
rect 6114 10455 6148 10461
rect 6114 10427 6148 10455
rect 6114 10387 6148 10389
rect 6114 10355 6148 10387
rect 6114 10285 6148 10317
rect 6114 10283 6148 10285
rect 6114 10217 6148 10245
rect 6114 10211 6148 10217
rect 6114 10149 6148 10173
rect 6114 10139 6148 10149
rect 6114 10081 6148 10101
rect 6114 10067 6148 10081
rect 6114 10013 6148 10029
rect 6114 9995 6148 10013
rect 6114 9945 6148 9957
rect 6114 9923 6148 9945
rect 6114 9877 6148 9885
rect 6114 9851 6148 9877
rect 6114 9809 6148 9813
rect 6114 9779 6148 9809
rect 6114 9707 6148 9741
rect 6114 9639 6148 9669
rect 6114 9635 6148 9639
rect 6114 9571 6148 9597
rect 6114 9563 6148 9571
rect 6114 9503 6148 9525
rect 6114 9491 6148 9503
rect 6114 9435 6148 9453
rect 6114 9419 6148 9435
rect 6114 9367 6148 9381
rect 6114 9347 6148 9367
rect 6114 9299 6148 9309
rect 6114 9275 6148 9299
rect 6114 9231 6148 9237
rect 6114 9203 6148 9231
rect 6114 9163 6148 9165
rect 6114 9131 6148 9163
rect 6114 9061 6148 9093
rect 6114 9059 6148 9061
rect 6114 8993 6148 9021
rect 6114 8987 6148 8993
rect 6114 8925 6148 8949
rect 6114 8915 6148 8925
rect 6114 8857 6148 8877
rect 6114 8843 6148 8857
rect 6114 8789 6148 8805
rect 6114 8771 6148 8789
rect 6114 8721 6148 8733
rect 6114 8699 6148 8721
rect 6114 8653 6148 8661
rect 6114 8627 6148 8653
rect 6114 8585 6148 8589
rect 6114 8555 6148 8585
rect 6114 8483 6148 8517
rect 6114 8415 6148 8445
rect 6114 8411 6148 8415
rect 6114 8347 6148 8373
rect 6114 8339 6148 8347
rect 6114 8279 6148 8301
rect 6114 8267 6148 8279
rect 6114 8211 6148 8229
rect 6114 8195 6148 8211
rect 6114 8143 6148 8157
rect 6114 8123 6148 8143
rect 6114 8075 6148 8085
rect 6114 8051 6148 8075
rect 6114 8007 6148 8013
rect 6114 7979 6148 8007
rect 6114 7939 6148 7941
rect 6114 7907 6148 7939
rect 6114 7837 6148 7869
rect 6114 7835 6148 7837
rect 6114 7769 6148 7797
rect 6114 7763 6148 7769
rect 6114 7701 6148 7725
rect 6114 7691 6148 7701
rect 6114 7633 6148 7653
rect 6114 7619 6148 7633
rect 6114 7565 6148 7581
rect 6114 7547 6148 7565
rect 6114 7497 6148 7509
rect 6114 7475 6148 7497
rect 6114 7429 6148 7437
rect 6114 7403 6148 7429
rect 6114 7361 6148 7365
rect 6114 7331 6148 7361
rect 6114 7259 6148 7293
rect 6114 7191 6148 7221
rect 6114 7187 6148 7191
rect 6114 7123 6148 7149
rect 6114 7115 6148 7123
rect 6114 7055 6148 7077
rect 6114 7043 6148 7055
rect 6114 6987 6148 7005
rect 6114 6971 6148 6987
rect 6114 6919 6148 6933
rect 6114 6899 6148 6919
rect 6114 6851 6148 6861
rect 6114 6827 6148 6851
rect 6114 6783 6148 6789
rect 6114 6755 6148 6783
rect 6114 6715 6148 6716
rect 6114 6682 6148 6715
rect 6114 6613 6148 6643
rect 6114 6609 6148 6613
rect 6114 6545 6148 6570
rect 6114 6536 6148 6545
rect 6114 6477 6148 6497
rect 6114 6463 6148 6477
rect 6114 6409 6148 6424
rect 6114 6390 6148 6409
rect 6114 6341 6148 6351
rect 6114 6317 6148 6341
rect 6114 6273 6148 6278
rect 6114 6244 6148 6273
rect 6114 6171 6148 6205
rect 6114 6103 6148 6132
rect 6114 6098 6148 6103
rect 6114 6035 6148 6059
rect 6114 6025 6148 6035
rect 6114 5967 6148 5986
rect 6114 5952 6148 5967
rect 6114 5899 6148 5913
rect 6114 5879 6148 5899
rect 6114 5831 6148 5840
rect 6114 5806 6148 5831
rect 6114 5763 6148 5767
rect 6114 5733 6148 5763
rect 6114 5661 6148 5694
rect 6114 5660 6148 5661
rect 6114 5593 6148 5621
rect 6114 5587 6148 5593
rect 6114 5525 6148 5548
rect 6114 5514 6148 5525
rect 6114 5457 6148 5475
rect 6114 5441 6148 5457
rect 6114 5389 6148 5402
rect 6114 5368 6148 5389
rect 6114 5321 6148 5329
rect 6114 5295 6148 5321
rect 6114 5253 6148 5256
rect 6114 5222 6148 5253
rect 6114 5151 6148 5183
rect 6114 5149 6148 5151
rect 6114 5083 6148 5110
rect 6114 5076 6148 5083
rect 6114 5015 6148 5037
rect 6114 5003 6148 5015
rect 6114 4947 6148 4964
rect 6114 4930 6148 4947
rect 6114 4879 6148 4891
rect 6114 4857 6148 4879
rect 6114 4811 6148 4818
rect 6114 4784 6148 4811
rect 6114 4743 6148 4745
rect 6114 4711 6148 4743
rect 6114 4641 6148 4672
rect 6114 4638 6148 4641
rect 6114 4573 6148 4599
rect 6114 4565 6148 4573
rect 6114 4505 6148 4526
rect 6114 4492 6148 4505
rect 6114 4437 6148 4453
rect 6114 4419 6148 4437
rect 6114 4369 6148 4380
rect 6114 4346 6148 4369
rect 6114 4301 6148 4307
rect 6114 4273 6148 4301
rect 6114 4233 6148 4234
rect 6114 4200 6148 4233
rect 6114 4131 6148 4161
rect 6114 4127 6148 4131
rect 6114 4063 6148 4088
rect 6114 4054 6148 4063
rect 6114 3995 6148 4015
rect 6114 3981 6148 3995
rect 6114 3927 6148 3942
rect 6114 3908 6148 3927
rect 6114 3859 6148 3869
rect 6114 3835 6148 3859
rect 6114 3791 6148 3796
rect 6114 3762 6148 3791
rect 6114 3689 6148 3723
rect 6114 3621 6148 3650
rect 6114 3616 6148 3621
rect 6114 3553 6148 3577
rect 6114 3543 6148 3553
rect 3972 3397 4006 3429
rect 3972 3395 4006 3397
rect 1830 3349 1864 3357
rect 1830 3323 1864 3349
rect 1830 3281 1864 3285
rect 1830 3251 1864 3281
rect 4158 3453 4192 3487
rect 4158 3395 4192 3415
rect 4158 3381 4192 3395
rect 4276 3453 4310 3487
rect 4276 3395 4310 3415
rect 4276 3381 4310 3395
rect 4394 3453 4428 3487
rect 4394 3395 4428 3415
rect 4394 3381 4428 3395
rect 4512 3453 4546 3487
rect 4512 3395 4546 3415
rect 4512 3381 4546 3395
rect 4630 3453 4664 3487
rect 4630 3395 4664 3415
rect 4630 3381 4664 3395
rect 4748 3453 4782 3487
rect 4748 3395 4782 3415
rect 4748 3381 4782 3395
rect 4866 3453 4900 3487
rect 4866 3395 4900 3415
rect 4866 3381 4900 3395
rect 4984 3453 5018 3487
rect 4984 3395 5018 3415
rect 4984 3381 5018 3395
rect 5102 3453 5136 3487
rect 5102 3395 5136 3415
rect 5102 3381 5136 3395
rect 5220 3452 5254 3486
rect 5220 3395 5254 3414
rect 5220 3380 5254 3395
rect 5338 3452 5372 3486
rect 5338 3395 5372 3414
rect 5338 3380 5372 3395
rect 5456 3452 5490 3486
rect 5456 3395 5490 3414
rect 5456 3380 5490 3395
rect 5574 3452 5608 3486
rect 5574 3395 5608 3414
rect 5574 3380 5608 3395
rect 5692 3452 5726 3486
rect 5692 3395 5726 3414
rect 5692 3380 5726 3395
rect 5810 3452 5844 3486
rect 5810 3395 5844 3414
rect 5810 3380 5844 3395
rect 5928 3452 5962 3486
rect 5928 3395 5962 3414
rect 5928 3380 5962 3395
rect 6114 3485 6148 3504
rect 6114 3470 6148 3485
rect 6114 3417 6148 3431
rect 6114 3397 6148 3417
rect 3972 3329 4006 3357
rect 3972 3323 4006 3329
rect 3972 3251 4006 3285
rect 6114 3349 6148 3358
rect 6114 3324 6148 3349
rect 6114 3281 6148 3285
rect 6114 3251 6148 3281
rect -180 3179 -150 3213
rect -150 3179 -146 3213
rect -107 3179 -82 3213
rect -82 3179 -73 3213
rect -34 3179 -14 3213
rect -14 3179 0 3213
rect 39 3179 54 3213
rect 54 3179 73 3213
rect 112 3179 122 3213
rect 122 3179 146 3213
rect 185 3179 190 3213
rect 190 3179 219 3213
rect 258 3179 292 3213
rect 331 3179 360 3213
rect 360 3179 365 3213
rect 404 3179 428 3213
rect 428 3179 438 3213
rect 477 3179 496 3213
rect 496 3179 511 3213
rect 550 3179 564 3213
rect 564 3179 584 3213
rect 623 3179 632 3213
rect 632 3179 657 3213
rect 696 3179 700 3213
rect 700 3179 730 3213
rect 769 3179 802 3213
rect 802 3179 803 3213
rect 842 3179 870 3213
rect 870 3179 876 3213
rect 915 3179 938 3213
rect 938 3179 949 3213
rect 988 3179 1006 3213
rect 1006 3179 1022 3213
rect 1061 3179 1074 3213
rect 1074 3179 1095 3213
rect 1134 3179 1142 3213
rect 1142 3179 1168 3213
rect 1207 3179 1210 3213
rect 1210 3179 1241 3213
rect 1280 3179 1312 3213
rect 1312 3179 1314 3213
rect 1353 3179 1380 3213
rect 1380 3179 1387 3213
rect 1426 3179 1448 3213
rect 1448 3179 1460 3213
rect 1499 3179 1516 3213
rect 1516 3179 1533 3213
rect 1572 3179 1584 3213
rect 1584 3179 1606 3213
rect 1645 3179 1652 3213
rect 1652 3179 1679 3213
rect 1718 3179 1720 3213
rect 1720 3179 1752 3213
rect 1791 3179 1825 3213
rect 1864 3179 1898 3213
rect 1937 3179 1966 3213
rect 1966 3179 1971 3213
rect 2010 3179 2034 3213
rect 2034 3179 2044 3213
rect 2082 3179 2102 3213
rect 2102 3179 2116 3213
rect 2154 3179 2170 3213
rect 2170 3179 2188 3213
rect 2226 3179 2238 3213
rect 2238 3179 2260 3213
rect 2298 3179 2306 3213
rect 2306 3179 2332 3213
rect 2370 3179 2374 3213
rect 2374 3179 2404 3213
rect 2442 3179 2476 3213
rect 2514 3179 2544 3213
rect 2544 3179 2548 3213
rect 2586 3179 2612 3213
rect 2612 3179 2620 3213
rect 2658 3179 2680 3213
rect 2680 3179 2692 3213
rect 2730 3179 2748 3213
rect 2748 3179 2764 3213
rect 2802 3179 2816 3213
rect 2816 3179 2836 3213
rect 2874 3179 2884 3213
rect 2884 3179 2908 3213
rect 2946 3179 2952 3213
rect 2952 3179 2980 3213
rect 3018 3179 3020 3213
rect 3020 3179 3052 3213
rect 3090 3179 3122 3213
rect 3122 3179 3124 3213
rect 3162 3179 3190 3213
rect 3190 3179 3196 3213
rect 3234 3179 3258 3213
rect 3258 3179 3268 3213
rect 3306 3179 3326 3213
rect 3326 3179 3340 3213
rect 3378 3179 3394 3213
rect 3394 3179 3412 3213
rect 3450 3179 3462 3213
rect 3462 3179 3484 3213
rect 3522 3179 3530 3213
rect 3530 3179 3556 3213
rect 3594 3179 3598 3213
rect 3598 3179 3628 3213
rect 3666 3179 3700 3213
rect 3738 3179 3768 3213
rect 3768 3179 3772 3213
rect 3810 3179 3836 3213
rect 3836 3179 3844 3213
rect 3882 3179 3904 3213
rect 3904 3179 3916 3213
rect 3954 3179 3988 3213
rect 4026 3179 4040 3213
rect 4040 3179 4060 3213
rect 4098 3179 4108 3213
rect 4108 3179 4132 3213
rect 4170 3179 4176 3213
rect 4176 3179 4204 3213
rect 4242 3179 4244 3213
rect 4244 3179 4276 3213
rect 4314 3179 4346 3213
rect 4346 3179 4348 3213
rect 4386 3179 4414 3213
rect 4414 3179 4420 3213
rect 4458 3179 4482 3213
rect 4482 3179 4492 3213
rect 4530 3179 4550 3213
rect 4550 3179 4564 3213
rect 4602 3179 4618 3213
rect 4618 3179 4636 3213
rect 4674 3179 4686 3213
rect 4686 3179 4708 3213
rect 4746 3179 4754 3213
rect 4754 3179 4780 3213
rect 4818 3179 4822 3213
rect 4822 3179 4852 3213
rect 4890 3179 4924 3213
rect 4962 3179 4992 3213
rect 4992 3179 4996 3213
rect 5034 3179 5060 3213
rect 5060 3179 5068 3213
rect 5106 3179 5128 3213
rect 5128 3179 5140 3213
rect 5178 3179 5196 3213
rect 5196 3179 5212 3213
rect 5250 3179 5264 3213
rect 5264 3179 5284 3213
rect 5322 3179 5332 3213
rect 5332 3179 5356 3213
rect 5394 3179 5400 3213
rect 5400 3179 5428 3213
rect 5466 3179 5468 3213
rect 5468 3179 5500 3213
rect 5538 3179 5570 3213
rect 5570 3179 5572 3213
rect 5610 3179 5638 3213
rect 5638 3179 5644 3213
rect 5682 3179 5706 3213
rect 5706 3179 5716 3213
rect 5754 3179 5774 3213
rect 5774 3179 5788 3213
rect 5826 3179 5842 3213
rect 5842 3179 5860 3213
rect 5898 3179 5910 3213
rect 5910 3179 5932 3213
rect 5970 3179 5978 3213
rect 5978 3179 6004 3213
rect 6042 3179 6046 3213
rect 6046 3179 6076 3213
rect 9162 38722 9196 38756
rect 9237 38723 9240 38756
rect 9240 38723 9271 38756
rect 9312 38723 9342 38756
rect 9342 38723 9346 38756
rect 9422 38723 9444 38756
rect 9444 38723 9456 38756
rect 9494 38723 9512 38756
rect 9512 38723 9528 38756
rect 9566 38723 9580 38756
rect 9580 38723 9600 38756
rect 9638 38723 9648 38756
rect 9648 38723 9672 38756
rect 9710 38723 9716 38756
rect 9716 38723 9744 38756
rect 9782 38723 9784 38756
rect 9784 38723 9816 38756
rect 9854 38723 9886 38756
rect 9886 38723 9888 38756
rect 9926 38723 9954 38756
rect 9954 38723 9960 38756
rect 9998 38723 10022 38756
rect 10022 38723 10032 38756
rect 10070 38723 10090 38756
rect 10090 38723 10104 38756
rect 10142 38723 10158 38756
rect 10158 38723 10176 38756
rect 9237 38722 9271 38723
rect 9312 38722 9346 38723
rect 9422 38722 9456 38723
rect 9494 38722 9528 38723
rect 9566 38722 9600 38723
rect 9638 38722 9672 38723
rect 9710 38722 9744 38723
rect 9782 38722 9816 38723
rect 9854 38722 9888 38723
rect 9926 38722 9960 38723
rect 9998 38722 10032 38723
rect 10070 38722 10104 38723
rect 10142 38722 10176 38723
rect 10214 38722 10248 38756
rect 10286 38723 10294 38756
rect 10294 38723 10320 38756
rect 10358 38723 10362 38756
rect 10362 38723 10392 38756
rect 10430 38723 10464 38756
rect 10502 38723 10532 38756
rect 10532 38723 10536 38756
rect 10574 38723 10600 38756
rect 10600 38723 10608 38756
rect 10646 38723 10668 38756
rect 10668 38723 10680 38756
rect 10718 38723 10736 38756
rect 10736 38723 10752 38756
rect 10790 38723 10804 38756
rect 10804 38723 10824 38756
rect 10862 38723 10872 38756
rect 10872 38723 10896 38756
rect 10934 38723 10940 38756
rect 10940 38723 10968 38756
rect 11006 38723 11008 38756
rect 11008 38723 11040 38756
rect 11078 38723 11110 38756
rect 11110 38723 11112 38756
rect 11150 38723 11178 38756
rect 11178 38723 11184 38756
rect 11222 38723 11246 38756
rect 11246 38723 11256 38756
rect 11294 38723 11314 38756
rect 11314 38723 11328 38756
rect 10286 38722 10320 38723
rect 10358 38722 10392 38723
rect 10430 38722 10464 38723
rect 10502 38722 10536 38723
rect 10574 38722 10608 38723
rect 10646 38722 10680 38723
rect 10718 38722 10752 38723
rect 10790 38722 10824 38723
rect 10862 38722 10896 38723
rect 10934 38722 10968 38723
rect 11006 38722 11040 38723
rect 11078 38722 11112 38723
rect 11150 38722 11184 38723
rect 11222 38722 11256 38723
rect 11294 38722 11328 38723
rect 11366 38722 11400 38756
rect 11438 38722 11472 38756
rect 11510 38723 11512 38756
rect 11512 38723 11544 38756
rect 11583 38723 11614 38756
rect 11614 38723 11617 38756
rect 11656 38723 11682 38756
rect 11682 38723 11690 38756
rect 11729 38723 11750 38756
rect 11750 38723 11763 38756
rect 11802 38723 11818 38756
rect 11818 38723 11836 38756
rect 11875 38723 11886 38756
rect 11886 38723 11909 38756
rect 11948 38723 11954 38756
rect 11954 38723 11982 38756
rect 12021 38723 12022 38756
rect 12022 38723 12055 38756
rect 12094 38723 12124 38756
rect 12124 38723 12128 38756
rect 12167 38723 12192 38756
rect 12192 38723 12201 38756
rect 12240 38723 12260 38756
rect 12260 38723 12274 38756
rect 12313 38723 12328 38756
rect 12328 38723 12347 38756
rect 12386 38723 12396 38756
rect 12396 38723 12420 38756
rect 12459 38723 12464 38756
rect 12464 38723 12493 38756
rect 12532 38723 12566 38756
rect 12605 38723 12634 38756
rect 12634 38723 12639 38756
rect 12678 38723 12702 38756
rect 12702 38723 12712 38756
rect 12751 38723 12770 38756
rect 12770 38723 12785 38756
rect 12824 38723 12838 38756
rect 12838 38723 12858 38756
rect 12897 38723 12906 38756
rect 12906 38723 12931 38756
rect 12970 38723 12974 38756
rect 12974 38723 13004 38756
rect 13043 38723 13076 38756
rect 13076 38723 13077 38756
rect 13116 38723 13144 38756
rect 13144 38723 13150 38756
rect 11510 38722 11544 38723
rect 11583 38722 11617 38723
rect 11656 38722 11690 38723
rect 11729 38722 11763 38723
rect 11802 38722 11836 38723
rect 11875 38722 11909 38723
rect 11948 38722 11982 38723
rect 12021 38722 12055 38723
rect 12094 38722 12128 38723
rect 12167 38722 12201 38723
rect 12240 38722 12274 38723
rect 12313 38722 12347 38723
rect 12386 38722 12420 38723
rect 12459 38722 12493 38723
rect 12532 38722 12566 38723
rect 12605 38722 12639 38723
rect 12678 38722 12712 38723
rect 12751 38722 12785 38723
rect 12824 38722 12858 38723
rect 12897 38722 12931 38723
rect 12970 38722 13004 38723
rect 13043 38722 13077 38723
rect 13116 38722 13150 38723
rect 13189 38722 13223 38756
rect 13262 38723 13280 38756
rect 13280 38723 13296 38756
rect 13335 38723 13348 38756
rect 13348 38723 13369 38756
rect 13408 38723 13416 38756
rect 13416 38723 13442 38756
rect 13481 38723 13484 38756
rect 13484 38723 13515 38756
rect 13554 38723 13586 38756
rect 13586 38723 13588 38756
rect 13627 38723 13654 38756
rect 13654 38723 13661 38756
rect 13700 38723 13722 38756
rect 13722 38723 13734 38756
rect 13773 38723 13790 38756
rect 13790 38723 13807 38756
rect 13846 38723 13858 38756
rect 13858 38723 13880 38756
rect 13919 38723 13926 38756
rect 13926 38723 13953 38756
rect 13992 38723 13994 38756
rect 13994 38723 14026 38756
rect 14065 38723 14096 38756
rect 14096 38723 14099 38756
rect 14138 38723 14164 38756
rect 14164 38723 14172 38756
rect 14211 38723 14232 38756
rect 14232 38723 14245 38756
rect 14284 38723 14300 38756
rect 14300 38723 14318 38756
rect 14357 38723 14368 38756
rect 14368 38723 14391 38756
rect 14430 38723 14436 38756
rect 14436 38723 14464 38756
rect 14503 38723 14504 38756
rect 14504 38723 14537 38756
rect 14576 38723 14606 38756
rect 14606 38723 14610 38756
rect 14649 38723 14674 38756
rect 14674 38723 14683 38756
rect 14722 38723 14742 38756
rect 14742 38723 14756 38756
rect 14795 38723 14810 38756
rect 14810 38723 14829 38756
rect 14868 38723 14878 38756
rect 14878 38723 14902 38756
rect 13262 38722 13296 38723
rect 13335 38722 13369 38723
rect 13408 38722 13442 38723
rect 13481 38722 13515 38723
rect 13554 38722 13588 38723
rect 13627 38722 13661 38723
rect 13700 38722 13734 38723
rect 13773 38722 13807 38723
rect 13846 38722 13880 38723
rect 13919 38722 13953 38723
rect 13992 38722 14026 38723
rect 14065 38722 14099 38723
rect 14138 38722 14172 38723
rect 14211 38722 14245 38723
rect 14284 38722 14318 38723
rect 14357 38722 14391 38723
rect 14430 38722 14464 38723
rect 14503 38722 14537 38723
rect 14576 38722 14610 38723
rect 14649 38722 14683 38723
rect 14722 38722 14756 38723
rect 14795 38722 14829 38723
rect 14868 38722 14902 38723
rect 9088 38655 9122 38684
rect 9088 38650 9122 38655
rect 9088 38587 9122 38611
rect 9088 38577 9122 38587
rect 9088 38519 9122 38538
rect 9088 38504 9122 38519
rect 9088 38451 9122 38465
rect 9088 38431 9122 38451
rect 9088 38383 9122 38392
rect 9088 38358 9122 38383
rect 9088 38315 9122 38319
rect 9088 38285 9122 38315
rect 9088 38213 9122 38246
rect 9088 38212 9122 38213
rect 9088 38145 9122 38173
rect 9088 38139 9122 38145
rect 9088 38077 9122 38100
rect 9088 38066 9122 38077
rect 9088 38009 9122 38027
rect 9088 37993 9122 38009
rect 9088 37941 9122 37954
rect 9088 37920 9122 37941
rect 9088 37873 9122 37881
rect 9088 37847 9122 37873
rect 9088 37805 9122 37808
rect 9088 37774 9122 37805
rect 9088 37703 9122 37735
rect 9088 37701 9122 37703
rect 9088 37635 9122 37662
rect 9088 37628 9122 37635
rect 9088 37567 9122 37589
rect 9088 37555 9122 37567
rect 9088 37499 9122 37516
rect 9088 37482 9122 37499
rect 9088 37431 9122 37443
rect 9088 37409 9122 37431
rect 9088 37363 9122 37370
rect 9088 37336 9122 37363
rect 9088 37295 9122 37297
rect 9088 37263 9122 37295
rect 9088 37193 9122 37224
rect 9088 37190 9122 37193
rect 9088 37125 9122 37151
rect 9088 37117 9122 37125
rect 9088 37057 9122 37078
rect 9088 37044 9122 37057
rect 9088 36989 9122 37005
rect 9088 36971 9122 36989
rect 9088 36921 9122 36932
rect 9088 36898 9122 36921
rect 9088 36853 9122 36859
rect 9088 36825 9122 36853
rect 9088 36785 9122 36786
rect 9088 36752 9122 36785
rect 9088 36683 9122 36713
rect 9088 36679 9122 36683
rect 9088 36615 9122 36640
rect 9088 36606 9122 36615
rect 9088 36547 9122 36567
rect 9088 36533 9122 36547
rect 9088 36479 9122 36494
rect 9088 36460 9122 36479
rect 9088 36411 9122 36421
rect 9088 36387 9122 36411
rect 9088 36343 9122 36348
rect 9088 36314 9122 36343
rect 9088 36241 9122 36275
rect 9088 36173 9122 36202
rect 9088 36168 9122 36173
rect 9088 36105 9122 36129
rect 9088 36095 9122 36105
rect 9088 36037 9122 36056
rect 9088 36022 9122 36037
rect 9088 35969 9122 35983
rect 9088 35949 9122 35969
rect 9088 35901 9122 35910
rect 9088 35876 9122 35901
rect 9088 35833 9122 35837
rect 9088 35803 9122 35833
rect 9088 35731 9122 35764
rect 9088 35730 9122 35731
rect 9088 35663 9122 35691
rect 9088 35657 9122 35663
rect 9088 35595 9122 35618
rect 9088 35584 9122 35595
rect 9088 35527 9122 35545
rect 9088 35511 9122 35527
rect 9088 35459 9122 35472
rect 9088 35438 9122 35459
rect 9088 35391 9122 35399
rect 9088 35365 9122 35391
rect 9088 35323 9122 35326
rect 9088 35292 9122 35323
rect 9088 35221 9122 35253
rect 9088 35219 9122 35221
rect 9088 35153 9122 35180
rect 9088 35146 9122 35153
rect 9088 35085 9122 35108
rect 9088 35074 9122 35085
rect 9088 35017 9122 35036
rect 9088 35002 9122 35017
rect 9088 34949 9122 34964
rect 9088 34930 9122 34949
rect 9088 34881 9122 34892
rect 9088 34858 9122 34881
rect 9088 34813 9122 34820
rect 9088 34786 9122 34813
rect 9088 34745 9122 34748
rect 9088 34714 9122 34745
rect 9088 34643 9122 34676
rect 9088 34642 9122 34643
rect 9088 34575 9122 34604
rect 9088 34570 9122 34575
rect 9088 34507 9122 34532
rect 9088 34498 9122 34507
rect 9088 34439 9122 34460
rect 9088 34426 9122 34439
rect 9088 34371 9122 34388
rect 9088 34354 9122 34371
rect 9088 34303 9122 34316
rect 9088 34282 9122 34303
rect 9088 34235 9122 34244
rect 9088 34210 9122 34235
rect 9088 34167 9122 34172
rect 9088 34138 9122 34167
rect 9088 34099 9122 34100
rect 9088 34066 9122 34099
rect 9088 33997 9122 34028
rect 9088 33994 9122 33997
rect 9088 33929 9122 33956
rect 9088 33922 9122 33929
rect 9088 33861 9122 33884
rect 9088 33850 9122 33861
rect 9088 33793 9122 33812
rect 9088 33778 9122 33793
rect 9088 33725 9122 33740
rect 9088 33706 9122 33725
rect 9088 33657 9122 33668
rect 9088 33634 9122 33657
rect 9088 33589 9122 33596
rect 9088 33562 9122 33589
rect 9088 33521 9122 33524
rect 9088 33490 9122 33521
rect 9088 33419 9122 33452
rect 9088 33418 9122 33419
rect 9088 33351 9122 33380
rect 9088 33346 9122 33351
rect 9088 33283 9122 33308
rect 9088 33274 9122 33283
rect 9088 33215 9122 33236
rect 9088 33202 9122 33215
rect 9088 33147 9122 33164
rect 9088 33130 9122 33147
rect 9088 33079 9122 33092
rect 9088 33058 9122 33079
rect 9088 33011 9122 33020
rect 9088 32986 9122 33011
rect 9088 32943 9122 32948
rect 9088 32914 9122 32943
rect 9088 32875 9122 32876
rect 9088 32842 9122 32875
rect 9088 32773 9122 32804
rect 9088 32770 9122 32773
rect 9088 32705 9122 32732
rect 9088 32698 9122 32705
rect 9088 32637 9122 32660
rect 9088 32626 9122 32637
rect 9088 32569 9122 32588
rect 9088 32554 9122 32569
rect 9088 32501 9122 32516
rect 9088 32482 9122 32501
rect 9088 32433 9122 32444
rect 9088 32410 9122 32433
rect 9088 32365 9122 32372
rect 9088 32338 9122 32365
rect 9088 32297 9122 32300
rect 9088 32266 9122 32297
rect 9088 32195 9122 32228
rect 9088 32194 9122 32195
rect 9088 32127 9122 32156
rect 9088 32122 9122 32127
rect 9088 32059 9122 32084
rect 9088 32050 9122 32059
rect 9088 31991 9122 32012
rect 9088 31978 9122 31991
rect 9088 31923 9122 31940
rect 9088 31906 9122 31923
rect 9088 31855 9122 31868
rect 9088 31834 9122 31855
rect 9088 31787 9122 31796
rect 9088 31762 9122 31787
rect 9088 31719 9122 31724
rect 9088 31690 9122 31719
rect 9088 31651 9122 31652
rect 9088 31618 9122 31651
rect 9088 31549 9122 31580
rect 9088 31546 9122 31549
rect 9088 31481 9122 31508
rect 9088 31474 9122 31481
rect 9088 31413 9122 31436
rect 9088 31402 9122 31413
rect 9088 31345 9122 31364
rect 9088 31330 9122 31345
rect 9088 31277 9122 31292
rect 9088 31258 9122 31277
rect 9088 31209 9122 31220
rect 9088 31186 9122 31209
rect 9088 31141 9122 31148
rect 9088 31114 9122 31141
rect 9088 31073 9122 31076
rect 9088 31042 9122 31073
rect 9088 30971 9122 31004
rect 9088 30970 9122 30971
rect 9088 30903 9122 30932
rect 9088 30898 9122 30903
rect 9088 30835 9122 30860
rect 9088 30826 9122 30835
rect 9088 30767 9122 30788
rect 9088 30754 9122 30767
rect 9088 30699 9122 30716
rect 9088 30682 9122 30699
rect 9088 30631 9122 30644
rect 9088 30610 9122 30631
rect 9088 30563 9122 30572
rect 9088 30538 9122 30563
rect 9088 30495 9122 30500
rect 9088 30466 9122 30495
rect 9088 30427 9122 30428
rect 9088 30394 9122 30427
rect 9088 30325 9122 30356
rect 9088 30322 9122 30325
rect 9088 30257 9122 30284
rect 9088 30250 9122 30257
rect 9088 30189 9122 30212
rect 9088 30178 9122 30189
rect 9088 30121 9122 30140
rect 9088 30106 9122 30121
rect 9088 30053 9122 30068
rect 9088 30034 9122 30053
rect 9088 29985 9122 29996
rect 9088 29962 9122 29985
rect 9088 29917 9122 29924
rect 9088 29890 9122 29917
rect 9088 29849 9122 29852
rect 9088 29818 9122 29849
rect 9088 29747 9122 29780
rect 9088 29746 9122 29747
rect 9088 29679 9122 29708
rect 9088 29674 9122 29679
rect 9088 29611 9122 29636
rect 9088 29602 9122 29611
rect 9088 29543 9122 29564
rect 9088 29530 9122 29543
rect 9088 29475 9122 29492
rect 9088 29458 9122 29475
rect 9088 29407 9122 29420
rect 9088 29386 9122 29407
rect 9088 29339 9122 29348
rect 9088 29314 9122 29339
rect 9088 29271 9122 29276
rect 9088 29242 9122 29271
rect 9088 29203 9122 29204
rect 9088 29170 9122 29203
rect 9088 29101 9122 29132
rect 9088 29098 9122 29101
rect 9088 29033 9122 29060
rect 9088 29026 9122 29033
rect 9088 28965 9122 28988
rect 9088 28954 9122 28965
rect 9088 28897 9122 28916
rect 9088 28882 9122 28897
rect 9088 28829 9122 28844
rect 9088 28810 9122 28829
rect 9088 28761 9122 28772
rect 9088 28738 9122 28761
rect 9088 28693 9122 28700
rect 9088 28666 9122 28693
rect 9088 28625 9122 28628
rect 9088 28594 9122 28625
rect 9088 28523 9122 28556
rect 9088 28522 9122 28523
rect 9088 28455 9122 28484
rect 9088 28450 9122 28455
rect 9088 28387 9122 28412
rect 9088 28378 9122 28387
rect 9088 28319 9122 28340
rect 9088 28306 9122 28319
rect 9088 28251 9122 28268
rect 9088 28234 9122 28251
rect 9088 28183 9122 28196
rect 9088 28162 9122 28183
rect 9088 28115 9122 28124
rect 9088 28090 9122 28115
rect 9088 28047 9122 28052
rect 9088 28018 9122 28047
rect 9088 27979 9122 27980
rect 9088 27946 9122 27979
rect 9088 27877 9122 27908
rect 9088 27874 9122 27877
rect 9088 27809 9122 27836
rect 9088 27802 9122 27809
rect 9088 27741 9122 27764
rect 9088 27730 9122 27741
rect 9088 27673 9122 27692
rect 9088 27658 9122 27673
rect 9088 27605 9122 27620
rect 9088 27586 9122 27605
rect 9088 27537 9122 27548
rect 9088 27514 9122 27537
rect 9088 27469 9122 27476
rect 9088 27442 9122 27469
rect 9088 27401 9122 27404
rect 9088 27370 9122 27401
rect 9088 27299 9122 27332
rect 9088 27298 9122 27299
rect 9088 27231 9122 27260
rect 9088 27226 9122 27231
rect 9088 27163 9122 27188
rect 9088 27154 9122 27163
rect 9088 27095 9122 27116
rect 9088 27082 9122 27095
rect 9088 27027 9122 27044
rect 9088 27010 9122 27027
rect 9088 26959 9122 26972
rect 9088 26938 9122 26959
rect 9088 26891 9122 26900
rect 9088 26866 9122 26891
rect 9088 26823 9122 26828
rect 9088 26794 9122 26823
rect 9088 26755 9122 26756
rect 9088 26722 9122 26755
rect 9088 26653 9122 26684
rect 9088 26650 9122 26653
rect 9088 26585 9122 26612
rect 9088 26578 9122 26585
rect 9088 26517 9122 26540
rect 9088 26506 9122 26517
rect 9088 26449 9122 26468
rect 9088 26434 9122 26449
rect 9088 26381 9122 26396
rect 9088 26362 9122 26381
rect 9088 26313 9122 26324
rect 9088 26290 9122 26313
rect 9088 26245 9122 26252
rect 9088 26218 9122 26245
rect 9088 26177 9122 26180
rect 9088 26146 9122 26177
rect 9088 26075 9122 26108
rect 9088 26074 9122 26075
rect 9088 26007 9122 26036
rect 9088 26002 9122 26007
rect 9088 25939 9122 25964
rect 9088 25930 9122 25939
rect 9088 25871 9122 25892
rect 9088 25858 9122 25871
rect 9088 25803 9122 25820
rect 9088 25786 9122 25803
rect 9088 25735 9122 25748
rect 9088 25714 9122 25735
rect 9088 25667 9122 25676
rect 9088 25642 9122 25667
rect 9088 25599 9122 25604
rect 9088 25570 9122 25599
rect 9088 25531 9122 25532
rect 9088 25498 9122 25531
rect 9088 25429 9122 25460
rect 9088 25426 9122 25429
rect 9088 25361 9122 25388
rect 9088 25354 9122 25361
rect 9088 25293 9122 25316
rect 9088 25282 9122 25293
rect 9088 25225 9122 25244
rect 9088 25210 9122 25225
rect 9088 25157 9122 25172
rect 9088 25138 9122 25157
rect 9088 25089 9122 25100
rect 9088 25066 9122 25089
rect 9088 25021 9122 25028
rect 9088 24994 9122 25021
rect 9088 24953 9122 24956
rect 9088 24922 9122 24953
rect 9088 24851 9122 24884
rect 9088 24850 9122 24851
rect 9088 24783 9122 24812
rect 9088 24778 9122 24783
rect 9088 24715 9122 24740
rect 9088 24706 9122 24715
rect 9088 24647 9122 24668
rect 9088 24634 9122 24647
rect 9088 24579 9122 24596
rect 9088 24562 9122 24579
rect 9088 24511 9122 24524
rect 9088 24490 9122 24511
rect 9088 24443 9122 24452
rect 9088 24418 9122 24443
rect 9088 24375 9122 24380
rect 9088 24346 9122 24375
rect 9088 24307 9122 24308
rect 9088 24274 9122 24307
rect 9088 24205 9122 24236
rect 9088 24202 9122 24205
rect 9088 24137 9122 24164
rect 9088 24130 9122 24137
rect 9088 24069 9122 24092
rect 9088 24058 9122 24069
rect 9088 24001 9122 24020
rect 9088 23986 9122 24001
rect 9088 23933 9122 23948
rect 9088 23914 9122 23933
rect 9088 23865 9122 23876
rect 9088 23842 9122 23865
rect 9088 23797 9122 23804
rect 9088 23770 9122 23797
rect 9088 23729 9122 23732
rect 9088 23698 9122 23729
rect 9088 23627 9122 23660
rect 9088 23626 9122 23627
rect 9088 23559 9122 23588
rect 9088 23554 9122 23559
rect 9088 23491 9122 23516
rect 9088 23482 9122 23491
rect 9088 23423 9122 23444
rect 9088 23410 9122 23423
rect 9088 23355 9122 23372
rect 9088 23338 9122 23355
rect 9088 23287 9122 23300
rect 9088 23266 9122 23287
rect 9088 23219 9122 23228
rect 9088 23194 9122 23219
rect 9088 23151 9122 23156
rect 9088 23122 9122 23151
rect 9088 23083 9122 23084
rect 9088 23050 9122 23083
rect 9088 22981 9122 23012
rect 9088 22978 9122 22981
rect 9088 22913 9122 22940
rect 9088 22906 9122 22913
rect 9088 22845 9122 22868
rect 9088 22834 9122 22845
rect 9088 22777 9122 22796
rect 9088 22762 9122 22777
rect 9088 22709 9122 22724
rect 9088 22690 9122 22709
rect 9088 22641 9122 22652
rect 9088 22618 9122 22641
rect 9088 22573 9122 22580
rect 9088 22546 9122 22573
rect 9088 22505 9122 22508
rect 9088 22474 9122 22505
rect 9088 22403 9122 22436
rect 9088 22402 9122 22403
rect 9088 22335 9122 22364
rect 9088 22330 9122 22335
rect 9088 22267 9122 22292
rect 9088 22258 9122 22267
rect 9088 22199 9122 22220
rect 9088 22186 9122 22199
rect 9088 22131 9122 22148
rect 9088 22114 9122 22131
rect 9088 22063 9122 22076
rect 9088 22042 9122 22063
rect 9088 21995 9122 22004
rect 9088 21970 9122 21995
rect 9088 21927 9122 21932
rect 9088 21898 9122 21927
rect 9088 21859 9122 21860
rect 9088 21826 9122 21859
rect 9088 21757 9122 21788
rect 9088 21754 9122 21757
rect 9088 21689 9122 21716
rect 9088 21682 9122 21689
rect 9088 21621 9122 21644
rect 9088 21610 9122 21621
rect 9088 21553 9122 21572
rect 9088 21538 9122 21553
rect 9088 21485 9122 21500
rect 9088 21466 9122 21485
rect 9088 21417 9122 21428
rect 9088 21394 9122 21417
rect 9088 21349 9122 21356
rect 9088 21322 9122 21349
rect 9088 21281 9122 21284
rect 9088 21250 9122 21281
rect 9088 21179 9122 21212
rect 9088 21178 9122 21179
rect 9088 21111 9122 21140
rect 9088 21106 9122 21111
rect 9088 21043 9122 21068
rect 9088 21034 9122 21043
rect 9088 20975 9122 20996
rect 9088 20962 9122 20975
rect 9088 20907 9122 20924
rect 9088 20890 9122 20907
rect 9088 20839 9122 20852
rect 9088 20818 9122 20839
rect 9088 20771 9122 20780
rect 9088 20746 9122 20771
rect 9088 20703 9122 20708
rect 9088 20674 9122 20703
rect 9088 20635 9122 20636
rect 9088 20602 9122 20635
rect 9088 20533 9122 20564
rect 9088 20530 9122 20533
rect 9088 20465 9122 20492
rect 9088 20458 9122 20465
rect 9088 20397 9122 20420
rect 9088 20386 9122 20397
rect 9088 20329 9122 20348
rect 9088 20314 9122 20329
rect 9088 20261 9122 20276
rect 9088 20242 9122 20261
rect 9088 20193 9122 20204
rect 9088 20170 9122 20193
rect 9088 20125 9122 20132
rect 9088 20098 9122 20125
rect 9088 20057 9122 20060
rect 9088 20026 9122 20057
rect 9088 19955 9122 19988
rect 9088 19954 9122 19955
rect 9088 19887 9122 19916
rect 9088 19882 9122 19887
rect 9088 19819 9122 19844
rect 9088 19810 9122 19819
rect 9088 19751 9122 19772
rect 9088 19738 9122 19751
rect 9088 19683 9122 19700
rect 9088 19666 9122 19683
rect 9088 19615 9122 19628
rect 9088 19594 9122 19615
rect 9088 19547 9122 19556
rect 9088 19522 9122 19547
rect 9088 19479 9122 19484
rect 9088 19450 9122 19479
rect 9088 19411 9122 19412
rect 9088 19378 9122 19411
rect 9088 19309 9122 19340
rect 9088 19306 9122 19309
rect 9088 19241 9122 19268
rect 9088 19234 9122 19241
rect 9088 19173 9122 19196
rect 9088 19162 9122 19173
rect 9088 19105 9122 19124
rect 9088 19090 9122 19105
rect 9088 19037 9122 19052
rect 9088 19018 9122 19037
rect 9088 18969 9122 18980
rect 9088 18946 9122 18969
rect 9088 18901 9122 18908
rect 9088 18874 9122 18901
rect 9088 18833 9122 18836
rect 9088 18802 9122 18833
rect 9088 18731 9122 18764
rect 9088 18730 9122 18731
rect 9088 18663 9122 18692
rect 9088 18658 9122 18663
rect 9088 18595 9122 18620
rect 9088 18586 9122 18595
rect 9088 18527 9122 18548
rect 9088 18514 9122 18527
rect 9088 18459 9122 18476
rect 9088 18442 9122 18459
rect 9088 18391 9122 18404
rect 9088 18370 9122 18391
rect 9088 18323 9122 18332
rect 9088 18298 9122 18323
rect 9088 18255 9122 18260
rect 9088 18226 9122 18255
rect 9088 18187 9122 18188
rect 9088 18154 9122 18187
rect 9088 18085 9122 18116
rect 9088 18082 9122 18085
rect 9088 18017 9122 18044
rect 9088 18010 9122 18017
rect 9088 17949 9122 17972
rect 9088 17938 9122 17949
rect 9088 17881 9122 17900
rect 9088 17866 9122 17881
rect 9088 17813 9122 17828
rect 9088 17794 9122 17813
rect 9088 17745 9122 17756
rect 9088 17722 9122 17745
rect 9088 17677 9122 17684
rect 9088 17650 9122 17677
rect 9088 17609 9122 17612
rect 9088 17578 9122 17609
rect 9088 17507 9122 17540
rect 9088 17506 9122 17507
rect 9088 17439 9122 17468
rect 9088 17434 9122 17439
rect 9088 17371 9122 17396
rect 9088 17362 9122 17371
rect 9088 17303 9122 17324
rect 9088 17290 9122 17303
rect 9088 17235 9122 17252
rect 9088 17218 9122 17235
rect 9088 17167 9122 17180
rect 9088 17146 9122 17167
rect 9088 17099 9122 17108
rect 9088 17074 9122 17099
rect 9088 17031 9122 17036
rect 9088 17002 9122 17031
rect 9088 16963 9122 16964
rect 9088 16930 9122 16963
rect 9088 16861 9122 16892
rect 9088 16858 9122 16861
rect 9088 16793 9122 16820
rect 9088 16786 9122 16793
rect 9088 16725 9122 16748
rect 9088 16714 9122 16725
rect 9088 16657 9122 16676
rect 9088 16642 9122 16657
rect 9088 16589 9122 16604
rect 9088 16570 9122 16589
rect 9088 16521 9122 16532
rect 9088 16498 9122 16521
rect 9088 16453 9122 16460
rect 9088 16426 9122 16453
rect 9088 16385 9122 16388
rect 9088 16354 9122 16385
rect 9088 16283 9122 16316
rect 9088 16282 9122 16283
rect 9088 16215 9122 16244
rect 9088 16210 9122 16215
rect 9088 16147 9122 16172
rect 9088 16138 9122 16147
rect 9088 16079 9122 16100
rect 9088 16066 9122 16079
rect 9088 16011 9122 16028
rect 9088 15994 9122 16011
rect 9088 15943 9122 15956
rect 9088 15922 9122 15943
rect 9088 15875 9122 15884
rect 9088 15850 9122 15875
rect 9088 15807 9122 15812
rect 9088 15778 9122 15807
rect 9088 15739 9122 15740
rect 9088 15706 9122 15739
rect 9088 15637 9122 15668
rect 9088 15634 9122 15637
rect 9088 15569 9122 15596
rect 9088 15562 9122 15569
rect 9088 15501 9122 15524
rect 9088 15490 9122 15501
rect 9088 15433 9122 15452
rect 9088 15418 9122 15433
rect 9088 15365 9122 15380
rect 9088 15346 9122 15365
rect 9088 15297 9122 15308
rect 9088 15274 9122 15297
rect 9088 15229 9122 15236
rect 9088 15202 9122 15229
rect 9088 15161 9122 15164
rect 9088 15130 9122 15161
rect 9088 15059 9122 15092
rect 9088 15058 9122 15059
rect 9088 14991 9122 15020
rect 9088 14986 9122 14991
rect 9088 14923 9122 14948
rect 9088 14914 9122 14923
rect 9088 14855 9122 14876
rect 9088 14842 9122 14855
rect 9088 14787 9122 14804
rect 9088 14770 9122 14787
rect 9088 14719 9122 14732
rect 9088 14698 9122 14719
rect 9088 14651 9122 14660
rect 9088 14626 9122 14651
rect 9088 14583 9122 14588
rect 9088 14554 9122 14583
rect 9088 14515 9122 14516
rect 9088 14482 9122 14515
rect 9088 14413 9122 14444
rect 9088 14410 9122 14413
rect 9088 14345 9122 14372
rect 9088 14338 9122 14345
rect 9088 14277 9122 14300
rect 9088 14266 9122 14277
rect 9088 14209 9122 14228
rect 9088 14194 9122 14209
rect 9088 14141 9122 14156
rect 9088 14122 9122 14141
rect 9088 14073 9122 14084
rect 9088 14050 9122 14073
rect 9088 14005 9122 14012
rect 9088 13978 9122 14005
rect 9088 13937 9122 13940
rect 9088 13906 9122 13937
rect 9088 13835 9122 13868
rect 9088 13834 9122 13835
rect 9088 13767 9122 13796
rect 9088 13762 9122 13767
rect 9088 13699 9122 13724
rect 9088 13690 9122 13699
rect 9088 13631 9122 13652
rect 9088 13618 9122 13631
rect 9088 13563 9122 13580
rect 9088 13546 9122 13563
rect 9088 13495 9122 13508
rect 9088 13474 9122 13495
rect 9088 13427 9122 13436
rect 9088 13402 9122 13427
rect 9088 13359 9122 13364
rect 9088 13330 9122 13359
rect 9088 13291 9122 13292
rect 9088 13258 9122 13291
rect 9088 13189 9122 13220
rect 9088 13186 9122 13189
rect 9088 13121 9122 13148
rect 9088 13114 9122 13121
rect 9088 13053 9122 13076
rect 9088 13042 9122 13053
rect 9088 12985 9122 13004
rect 9088 12970 9122 12985
rect 9088 12917 9122 12932
rect 9088 12898 9122 12917
rect 9088 12849 9122 12860
rect 9088 12826 9122 12849
rect 9088 12781 9122 12788
rect 9088 12754 9122 12781
rect 9088 12713 9122 12716
rect 9088 12682 9122 12713
rect 9088 12611 9122 12644
rect 9088 12610 9122 12611
rect 9088 12543 9122 12572
rect 9088 12538 9122 12543
rect 9088 12475 9122 12500
rect 9088 12466 9122 12475
rect 9088 12407 9122 12428
rect 9088 12394 9122 12407
rect 9088 12339 9122 12356
rect 9088 12322 9122 12339
rect 9088 12271 9122 12284
rect 9088 12250 9122 12271
rect 9088 12203 9122 12212
rect 9088 12178 9122 12203
rect 9088 12135 9122 12140
rect 9088 12106 9122 12135
rect 9088 12067 9122 12068
rect 9088 12034 9122 12067
rect 9088 11965 9122 11996
rect 9088 11962 9122 11965
rect 9088 11897 9122 11924
rect 9088 11890 9122 11897
rect 9088 11829 9122 11852
rect 9088 11818 9122 11829
rect 9088 11761 9122 11780
rect 9088 11746 9122 11761
rect 9088 11693 9122 11708
rect 9088 11674 9122 11693
rect 9088 11625 9122 11636
rect 9088 11602 9122 11625
rect 9088 11557 9122 11564
rect 9088 11530 9122 11557
rect 9088 11489 9122 11492
rect 9088 11458 9122 11489
rect 9088 11387 9122 11420
rect 9088 11386 9122 11387
rect 9088 11319 9122 11348
rect 9088 11314 9122 11319
rect 9088 11251 9122 11276
rect 9088 11242 9122 11251
rect 9088 11183 9122 11204
rect 9088 11170 9122 11183
rect 9088 11115 9122 11132
rect 9088 11098 9122 11115
rect 9088 11047 9122 11060
rect 9088 11026 9122 11047
rect 9088 10979 9122 10988
rect 9088 10954 9122 10979
rect 9088 10911 9122 10916
rect 9088 10882 9122 10911
rect 9088 10843 9122 10844
rect 9088 10810 9122 10843
rect 9088 10741 9122 10772
rect 9088 10738 9122 10741
rect 9088 10673 9122 10700
rect 9088 10666 9122 10673
rect 9088 10605 9122 10628
rect 9088 10594 9122 10605
rect 9088 10537 9122 10556
rect 9088 10522 9122 10537
rect 9088 10469 9122 10484
rect 9088 10450 9122 10469
rect 9088 10401 9122 10412
rect 9088 10378 9122 10401
rect 9088 10333 9122 10340
rect 9088 10306 9122 10333
rect 9088 10265 9122 10268
rect 9088 10234 9122 10265
rect 9088 10163 9122 10196
rect 9088 10162 9122 10163
rect 9088 10095 9122 10124
rect 9088 10090 9122 10095
rect 9088 10027 9122 10052
rect 9088 10018 9122 10027
rect 9088 9959 9122 9980
rect 9088 9946 9122 9959
rect 9088 9891 9122 9908
rect 9088 9874 9122 9891
rect 9088 9823 9122 9836
rect 9088 9802 9122 9823
rect 9088 9755 9122 9764
rect 9088 9730 9122 9755
rect 9088 9687 9122 9692
rect 9088 9658 9122 9687
rect 9088 9619 9122 9620
rect 9088 9586 9122 9619
rect 9088 9517 9122 9548
rect 9088 9514 9122 9517
rect 9088 9449 9122 9476
rect 9088 9442 9122 9449
rect 9088 9381 9122 9404
rect 9088 9370 9122 9381
rect 9088 9313 9122 9332
rect 9088 9298 9122 9313
rect 9088 9245 9122 9260
rect 9088 9226 9122 9245
rect 9088 9177 9122 9188
rect 9088 9154 9122 9177
rect 9088 9109 9122 9116
rect 9088 9082 9122 9109
rect 9088 9041 9122 9044
rect 9088 9010 9122 9041
rect 9088 8939 9122 8972
rect 9088 8938 9122 8939
rect 9088 8871 9122 8900
rect 9088 8866 9122 8871
rect 9088 8803 9122 8828
rect 9088 8794 9122 8803
rect 9088 8735 9122 8756
rect 9088 8722 9122 8735
rect 9088 8667 9122 8684
rect 9088 8650 9122 8667
rect 9088 8599 9122 8612
rect 9088 8578 9122 8599
rect 9088 8531 9122 8540
rect 9088 8506 9122 8531
rect 9088 8463 9122 8468
rect 9088 8434 9122 8463
rect 9088 8395 9122 8396
rect 9088 8362 9122 8395
rect 9088 8293 9122 8324
rect 9088 8290 9122 8293
rect 9088 8225 9122 8252
rect 9088 8218 9122 8225
rect 9088 8157 9122 8180
rect 9088 8146 9122 8157
rect 9088 8089 9122 8108
rect 9088 8074 9122 8089
rect 9088 8021 9122 8036
rect 9088 8002 9122 8021
rect 9088 7953 9122 7964
rect 9088 7930 9122 7953
rect 9088 7885 9122 7892
rect 9088 7858 9122 7885
rect 9088 7817 9122 7820
rect 9088 7786 9122 7817
rect 9088 7715 9122 7748
rect 9088 7714 9122 7715
rect 9088 7647 9122 7676
rect 9088 7642 9122 7647
rect 9088 7579 9122 7604
rect 9088 7570 9122 7579
rect 9088 7511 9122 7532
rect 9088 7498 9122 7511
rect 9088 7443 9122 7460
rect 9088 7426 9122 7443
rect 9088 7375 9122 7388
rect 9088 7354 9122 7375
rect 9088 7307 9122 7316
rect 9088 7282 9122 7307
rect 9088 7239 9122 7244
rect 9088 7210 9122 7239
rect 9088 7171 9122 7172
rect 9088 7138 9122 7171
rect 9088 7069 9122 7100
rect 9088 7066 9122 7069
rect 9088 7001 9122 7028
rect 9088 6994 9122 7001
rect 9088 6933 9122 6956
rect 9088 6922 9122 6933
rect 9088 6865 9122 6884
rect 9088 6850 9122 6865
rect 9088 6797 9122 6812
rect 9088 6778 9122 6797
rect 9088 6729 9122 6740
rect 9088 6706 9122 6729
rect 9088 6661 9122 6668
rect 9088 6634 9122 6661
rect 9088 6593 9122 6596
rect 9088 6562 9122 6593
rect 9088 6491 9122 6524
rect 9088 6490 9122 6491
rect 9088 6423 9122 6452
rect 9088 6418 9122 6423
rect 9088 6355 9122 6380
rect 9088 6346 9122 6355
rect 9088 6287 9122 6308
rect 9088 6274 9122 6287
rect 9088 6219 9122 6236
rect 9088 6202 9122 6219
rect 9088 6151 9122 6164
rect 9088 6130 9122 6151
rect 9088 6083 9122 6092
rect 9088 6058 9122 6083
rect 9088 6015 9122 6020
rect 9088 5986 9122 6015
rect 9088 5947 9122 5948
rect 9088 5914 9122 5947
rect 9088 5845 9122 5876
rect 9088 5842 9122 5845
rect 9088 5777 9122 5804
rect 9088 5770 9122 5777
rect 9088 5709 9122 5732
rect 9088 5698 9122 5709
rect 9088 5641 9122 5660
rect 9088 5626 9122 5641
rect 9088 5573 9122 5588
rect 9088 5554 9122 5573
rect 9088 5505 9122 5516
rect 9088 5482 9122 5505
rect 9088 5437 9122 5444
rect 9088 5410 9122 5437
rect 9088 5369 9122 5372
rect 9088 5338 9122 5369
rect 9088 5267 9122 5300
rect 9088 5266 9122 5267
rect 9088 5199 9122 5228
rect 9088 5194 9122 5199
rect 9088 5131 9122 5156
rect 9088 5122 9122 5131
rect 9088 5063 9122 5084
rect 9088 5050 9122 5063
rect 9088 4995 9122 5012
rect 9088 4978 9122 4995
rect 9088 4927 9122 4940
rect 9088 4906 9122 4927
rect 9088 4859 9122 4868
rect 9088 4834 9122 4859
rect 9088 4791 9122 4796
rect 9088 4762 9122 4791
rect 9088 4723 9122 4724
rect 9088 4690 9122 4723
rect 9088 4621 9122 4652
rect 9088 4618 9122 4621
rect 9088 4553 9122 4580
rect 9088 4546 9122 4553
rect 9088 4485 9122 4508
rect 9088 4474 9122 4485
rect 9088 4417 9122 4436
rect 9088 4402 9122 4417
rect 9088 4349 9122 4364
rect 9088 4330 9122 4349
rect 9088 4281 9122 4292
rect 9088 4258 9122 4281
rect 9088 4213 9122 4220
rect 9088 4186 9122 4213
rect 9088 4145 9122 4148
rect 9088 4114 9122 4145
rect 9088 4043 9122 4076
rect 9088 4042 9122 4043
rect 9088 3975 9122 4004
rect 9088 3970 9122 3975
rect 9088 3907 9122 3932
rect 9088 3898 9122 3907
rect 9088 3839 9122 3860
rect 9088 3826 9122 3839
rect 9088 3771 9122 3788
rect 9088 3754 9122 3771
rect 9088 3703 9122 3716
rect 9088 3682 9122 3703
rect 9088 3635 9122 3644
rect 9088 3610 9122 3635
rect 9088 3567 9122 3572
rect 9088 3538 9122 3567
rect 9088 3499 9122 3500
rect 9088 3466 9122 3499
rect 10226 38650 10260 38684
rect 10226 38607 10260 38611
rect 10226 38577 10260 38607
rect 10226 38505 10260 38538
rect 10226 38504 10260 38505
rect 10226 38437 10260 38465
rect 10226 38431 10260 38437
rect 10226 38369 10260 38392
rect 10226 38358 10260 38369
rect 10226 38301 10260 38319
rect 10226 38285 10260 38301
rect 10226 38233 10260 38246
rect 10226 38212 10260 38233
rect 10226 38165 10260 38173
rect 10226 38139 10260 38165
rect 10226 38097 10260 38100
rect 10226 38066 10260 38097
rect 10226 37995 10260 38027
rect 10226 37993 10260 37995
rect 10226 37927 10260 37954
rect 10226 37920 10260 37927
rect 10226 37859 10260 37881
rect 10226 37847 10260 37859
rect 10226 37791 10260 37808
rect 10226 37774 10260 37791
rect 10226 37723 10260 37735
rect 10226 37701 10260 37723
rect 10226 37655 10260 37662
rect 10226 37628 10260 37655
rect 10226 37587 10260 37589
rect 10226 37555 10260 37587
rect 10226 37485 10260 37516
rect 10226 37482 10260 37485
rect 10226 37417 10260 37443
rect 10226 37409 10260 37417
rect 10226 37349 10260 37370
rect 10226 37336 10260 37349
rect 10226 37281 10260 37297
rect 10226 37263 10260 37281
rect 10226 37213 10260 37224
rect 10226 37190 10260 37213
rect 10226 37145 10260 37151
rect 10226 37117 10260 37145
rect 10226 37077 10260 37078
rect 10226 37044 10260 37077
rect 10226 36975 10260 37005
rect 10226 36971 10260 36975
rect 10226 36907 10260 36932
rect 10226 36898 10260 36907
rect 10226 36839 10260 36859
rect 10226 36825 10260 36839
rect 10226 36771 10260 36786
rect 10226 36752 10260 36771
rect 10226 36703 10260 36713
rect 10226 36679 10260 36703
rect 10226 36635 10260 36640
rect 10226 36606 10260 36635
rect 10226 36533 10260 36567
rect 10226 36465 10260 36494
rect 10226 36460 10260 36465
rect 10226 36397 10260 36421
rect 10226 36387 10260 36397
rect 10226 36329 10260 36348
rect 10226 36314 10260 36329
rect 10226 36261 10260 36275
rect 10226 36241 10260 36261
rect 10226 36193 10260 36202
rect 10226 36168 10260 36193
rect 10226 36125 10260 36129
rect 10226 36095 10260 36125
rect 10226 36023 10260 36056
rect 10226 36022 10260 36023
rect 10226 35955 10260 35983
rect 10226 35949 10260 35955
rect 10226 35887 10260 35910
rect 10226 35876 10260 35887
rect 10226 35819 10260 35837
rect 10226 35803 10260 35819
rect 10226 35751 10260 35764
rect 10226 35730 10260 35751
rect 10226 35683 10260 35691
rect 10226 35657 10260 35683
rect 10226 35615 10260 35618
rect 10226 35584 10260 35615
rect 10226 35513 10260 35545
rect 10226 35511 10260 35513
rect 10226 35445 10260 35472
rect 10226 35438 10260 35445
rect 10226 35377 10260 35399
rect 10226 35365 10260 35377
rect 10226 35309 10260 35326
rect 10226 35292 10260 35309
rect 10226 35241 10260 35253
rect 10226 35219 10260 35241
rect 10226 35173 10260 35180
rect 10226 35146 10260 35173
rect 10226 35105 10260 35108
rect 10226 35074 10260 35105
rect 10226 35003 10260 35036
rect 10226 35002 10260 35003
rect 10226 34935 10260 34964
rect 10226 34930 10260 34935
rect 10226 34867 10260 34892
rect 10226 34858 10260 34867
rect 10226 34799 10260 34820
rect 10226 34786 10260 34799
rect 10226 34731 10260 34748
rect 10226 34714 10260 34731
rect 10226 34663 10260 34676
rect 10226 34642 10260 34663
rect 10226 34595 10260 34604
rect 10226 34570 10260 34595
rect 10226 34527 10260 34532
rect 10226 34498 10260 34527
rect 10226 34459 10260 34460
rect 10226 34426 10260 34459
rect 10226 34357 10260 34388
rect 10226 34354 10260 34357
rect 10226 34289 10260 34316
rect 10226 34282 10260 34289
rect 10226 34221 10260 34244
rect 10226 34210 10260 34221
rect 10226 34153 10260 34172
rect 10226 34138 10260 34153
rect 10226 34085 10260 34100
rect 10226 34066 10260 34085
rect 10226 34017 10260 34028
rect 10226 33994 10260 34017
rect 10226 33949 10260 33956
rect 10226 33922 10260 33949
rect 10226 33881 10260 33884
rect 10226 33850 10260 33881
rect 10226 33779 10260 33812
rect 10226 33778 10260 33779
rect 10226 33711 10260 33740
rect 10226 33706 10260 33711
rect 10226 33643 10260 33668
rect 10226 33634 10260 33643
rect 10226 33575 10260 33596
rect 10226 33562 10260 33575
rect 10226 33507 10260 33524
rect 10226 33490 10260 33507
rect 10226 33439 10260 33452
rect 10226 33418 10260 33439
rect 10226 33371 10260 33380
rect 10226 33346 10260 33371
rect 10226 33303 10260 33308
rect 10226 33274 10260 33303
rect 10226 33235 10260 33236
rect 10226 33202 10260 33235
rect 10226 33133 10260 33164
rect 10226 33130 10260 33133
rect 10226 33065 10260 33092
rect 10226 33058 10260 33065
rect 10226 32997 10260 33020
rect 10226 32986 10260 32997
rect 10226 32929 10260 32948
rect 10226 32914 10260 32929
rect 10226 32861 10260 32876
rect 10226 32842 10260 32861
rect 10226 32793 10260 32804
rect 10226 32770 10260 32793
rect 10226 32725 10260 32732
rect 10226 32698 10260 32725
rect 10226 32657 10260 32660
rect 10226 32626 10260 32657
rect 10226 32555 10260 32588
rect 10226 32554 10260 32555
rect 10226 32487 10260 32516
rect 10226 32482 10260 32487
rect 10226 32419 10260 32444
rect 10226 32410 10260 32419
rect 10226 32351 10260 32372
rect 10226 32338 10260 32351
rect 10226 32283 10260 32300
rect 10226 32266 10260 32283
rect 10226 32215 10260 32228
rect 10226 32194 10260 32215
rect 10226 32147 10260 32156
rect 10226 32122 10260 32147
rect 10226 32079 10260 32084
rect 10226 32050 10260 32079
rect 10226 32011 10260 32012
rect 10226 31978 10260 32011
rect 10226 31909 10260 31940
rect 10226 31906 10260 31909
rect 10226 31841 10260 31868
rect 10226 31834 10260 31841
rect 10226 31773 10260 31796
rect 10226 31762 10260 31773
rect 10226 31705 10260 31724
rect 10226 31690 10260 31705
rect 10226 31637 10260 31652
rect 10226 31618 10260 31637
rect 10226 31569 10260 31580
rect 10226 31546 10260 31569
rect 10226 31501 10260 31508
rect 10226 31474 10260 31501
rect 10226 31433 10260 31436
rect 10226 31402 10260 31433
rect 10226 31331 10260 31364
rect 10226 31330 10260 31331
rect 10226 31263 10260 31292
rect 10226 31258 10260 31263
rect 10226 31195 10260 31220
rect 10226 31186 10260 31195
rect 10226 31127 10260 31148
rect 10226 31114 10260 31127
rect 10226 31059 10260 31076
rect 10226 31042 10260 31059
rect 10226 30991 10260 31004
rect 10226 30970 10260 30991
rect 10226 30923 10260 30932
rect 10226 30898 10260 30923
rect 10226 30855 10260 30860
rect 10226 30826 10260 30855
rect 10226 30787 10260 30788
rect 10226 30754 10260 30787
rect 10226 30685 10260 30716
rect 10226 30682 10260 30685
rect 10226 30617 10260 30644
rect 10226 30610 10260 30617
rect 10226 30549 10260 30572
rect 10226 30538 10260 30549
rect 10226 30481 10260 30500
rect 10226 30466 10260 30481
rect 10226 30413 10260 30428
rect 10226 30394 10260 30413
rect 10226 30345 10260 30356
rect 10226 30322 10260 30345
rect 10226 30277 10260 30284
rect 10226 30250 10260 30277
rect 10226 30209 10260 30212
rect 10226 30178 10260 30209
rect 10226 30107 10260 30140
rect 10226 30106 10260 30107
rect 10226 30039 10260 30068
rect 10226 30034 10260 30039
rect 10226 29971 10260 29996
rect 10226 29962 10260 29971
rect 10226 29903 10260 29924
rect 10226 29890 10260 29903
rect 10226 29835 10260 29852
rect 10226 29818 10260 29835
rect 10226 29767 10260 29780
rect 10226 29746 10260 29767
rect 10226 29699 10260 29708
rect 10226 29674 10260 29699
rect 10226 29631 10260 29636
rect 10226 29602 10260 29631
rect 10226 29563 10260 29564
rect 10226 29530 10260 29563
rect 10226 29461 10260 29492
rect 10226 29458 10260 29461
rect 10226 29393 10260 29420
rect 10226 29386 10260 29393
rect 10226 29325 10260 29348
rect 10226 29314 10260 29325
rect 10226 29257 10260 29276
rect 10226 29242 10260 29257
rect 10226 29189 10260 29204
rect 10226 29170 10260 29189
rect 10226 29121 10260 29132
rect 10226 29098 10260 29121
rect 10226 29053 10260 29060
rect 10226 29026 10260 29053
rect 10226 28985 10260 28988
rect 10226 28954 10260 28985
rect 10226 28883 10260 28916
rect 10226 28882 10260 28883
rect 10226 28815 10260 28844
rect 10226 28810 10260 28815
rect 10226 28747 10260 28772
rect 10226 28738 10260 28747
rect 10226 28679 10260 28700
rect 10226 28666 10260 28679
rect 10226 28611 10260 28628
rect 10226 28594 10260 28611
rect 10226 28543 10260 28556
rect 10226 28522 10260 28543
rect 10226 28475 10260 28484
rect 10226 28450 10260 28475
rect 10226 28407 10260 28412
rect 10226 28378 10260 28407
rect 10226 28339 10260 28340
rect 10226 28306 10260 28339
rect 10226 28237 10260 28268
rect 10226 28234 10260 28237
rect 10226 28169 10260 28196
rect 10226 28162 10260 28169
rect 10226 28101 10260 28124
rect 10226 28090 10260 28101
rect 10226 28033 10260 28052
rect 10226 28018 10260 28033
rect 10226 27965 10260 27980
rect 10226 27946 10260 27965
rect 10226 27897 10260 27908
rect 10226 27874 10260 27897
rect 10226 27829 10260 27836
rect 10226 27802 10260 27829
rect 10226 27761 10260 27764
rect 10226 27730 10260 27761
rect 10226 27659 10260 27692
rect 10226 27658 10260 27659
rect 10226 27591 10260 27620
rect 10226 27586 10260 27591
rect 10226 27523 10260 27548
rect 10226 27514 10260 27523
rect 10226 27455 10260 27476
rect 10226 27442 10260 27455
rect 10226 27387 10260 27404
rect 10226 27370 10260 27387
rect 10226 27319 10260 27332
rect 10226 27298 10260 27319
rect 10226 27251 10260 27260
rect 10226 27226 10260 27251
rect 10226 27183 10260 27188
rect 10226 27154 10260 27183
rect 10226 27115 10260 27116
rect 10226 27082 10260 27115
rect 10226 27013 10260 27044
rect 10226 27010 10260 27013
rect 10226 26945 10260 26972
rect 10226 26938 10260 26945
rect 10226 26877 10260 26900
rect 10226 26866 10260 26877
rect 10226 26809 10260 26828
rect 10226 26794 10260 26809
rect 10226 26741 10260 26756
rect 10226 26722 10260 26741
rect 10226 26673 10260 26684
rect 10226 26650 10260 26673
rect 10226 26605 10260 26612
rect 10226 26578 10260 26605
rect 10226 26537 10260 26540
rect 10226 26506 10260 26537
rect 10226 26435 10260 26468
rect 10226 26434 10260 26435
rect 10226 26367 10260 26396
rect 10226 26362 10260 26367
rect 10226 26299 10260 26324
rect 10226 26290 10260 26299
rect 10226 26231 10260 26252
rect 10226 26218 10260 26231
rect 10226 26163 10260 26180
rect 10226 26146 10260 26163
rect 10226 26095 10260 26108
rect 10226 26074 10260 26095
rect 10226 26027 10260 26036
rect 10226 26002 10260 26027
rect 10226 25959 10260 25964
rect 10226 25930 10260 25959
rect 10226 25891 10260 25892
rect 10226 25858 10260 25891
rect 10226 25789 10260 25820
rect 10226 25786 10260 25789
rect 10226 25721 10260 25748
rect 10226 25714 10260 25721
rect 10226 25653 10260 25676
rect 10226 25642 10260 25653
rect 10226 25585 10260 25604
rect 10226 25570 10260 25585
rect 10226 25517 10260 25532
rect 10226 25498 10260 25517
rect 10226 25449 10260 25460
rect 10226 25426 10260 25449
rect 10226 25381 10260 25388
rect 10226 25354 10260 25381
rect 10226 25313 10260 25316
rect 10226 25282 10260 25313
rect 10226 25211 10260 25244
rect 10226 25210 10260 25211
rect 10226 25143 10260 25172
rect 10226 25138 10260 25143
rect 10226 25075 10260 25100
rect 10226 25066 10260 25075
rect 10226 25007 10260 25028
rect 10226 24994 10260 25007
rect 10226 24939 10260 24956
rect 10226 24922 10260 24939
rect 10226 24871 10260 24884
rect 10226 24850 10260 24871
rect 10226 24803 10260 24812
rect 10226 24778 10260 24803
rect 10226 24735 10260 24740
rect 10226 24706 10260 24735
rect 10226 24667 10260 24668
rect 10226 24634 10260 24667
rect 10226 24565 10260 24596
rect 10226 24562 10260 24565
rect 10226 24497 10260 24524
rect 10226 24490 10260 24497
rect 10226 24429 10260 24452
rect 10226 24418 10260 24429
rect 10226 24361 10260 24380
rect 10226 24346 10260 24361
rect 10226 24293 10260 24308
rect 10226 24274 10260 24293
rect 10226 24225 10260 24236
rect 10226 24202 10260 24225
rect 10226 24157 10260 24164
rect 10226 24130 10260 24157
rect 10226 24089 10260 24092
rect 10226 24058 10260 24089
rect 10226 23987 10260 24020
rect 10226 23986 10260 23987
rect 10226 23919 10260 23948
rect 10226 23914 10260 23919
rect 10226 23851 10260 23876
rect 10226 23842 10260 23851
rect 10226 23783 10260 23804
rect 10226 23770 10260 23783
rect 10226 23715 10260 23732
rect 10226 23698 10260 23715
rect 10226 23647 10260 23660
rect 10226 23626 10260 23647
rect 10226 23579 10260 23588
rect 10226 23554 10260 23579
rect 10226 23511 10260 23516
rect 10226 23482 10260 23511
rect 10226 23443 10260 23444
rect 10226 23410 10260 23443
rect 10226 23341 10260 23372
rect 10226 23338 10260 23341
rect 10226 23273 10260 23300
rect 10226 23266 10260 23273
rect 10226 23205 10260 23228
rect 10226 23194 10260 23205
rect 10226 23137 10260 23156
rect 10226 23122 10260 23137
rect 10226 23069 10260 23084
rect 10226 23050 10260 23069
rect 10226 23001 10260 23012
rect 10226 22978 10260 23001
rect 10226 22933 10260 22940
rect 10226 22906 10260 22933
rect 10226 22865 10260 22868
rect 10226 22834 10260 22865
rect 10226 22763 10260 22796
rect 10226 22762 10260 22763
rect 10226 22695 10260 22724
rect 10226 22690 10260 22695
rect 10226 22627 10260 22652
rect 10226 22618 10260 22627
rect 10226 22559 10260 22580
rect 10226 22546 10260 22559
rect 10226 22491 10260 22508
rect 10226 22474 10260 22491
rect 10226 22423 10260 22436
rect 10226 22402 10260 22423
rect 10226 22355 10260 22364
rect 10226 22330 10260 22355
rect 10226 22287 10260 22292
rect 10226 22258 10260 22287
rect 10226 22219 10260 22220
rect 10226 22186 10260 22219
rect 10226 22117 10260 22148
rect 10226 22114 10260 22117
rect 10226 22049 10260 22076
rect 10226 22042 10260 22049
rect 10226 21981 10260 22004
rect 10226 21970 10260 21981
rect 10226 21913 10260 21932
rect 10226 21898 10260 21913
rect 10226 21845 10260 21860
rect 10226 21826 10260 21845
rect 10226 21777 10260 21788
rect 10226 21754 10260 21777
rect 10226 21709 10260 21716
rect 10226 21682 10260 21709
rect 10226 21641 10260 21644
rect 10226 21610 10260 21641
rect 10226 21539 10260 21572
rect 10226 21538 10260 21539
rect 10226 21471 10260 21500
rect 10226 21466 10260 21471
rect 10226 21403 10260 21428
rect 10226 21394 10260 21403
rect 10226 21335 10260 21356
rect 10226 21322 10260 21335
rect 10226 21267 10260 21284
rect 10226 21250 10260 21267
rect 10226 21199 10260 21212
rect 10226 21178 10260 21199
rect 10226 21131 10260 21140
rect 10226 21106 10260 21131
rect 10226 21063 10260 21068
rect 10226 21034 10260 21063
rect 10226 20995 10260 20996
rect 10226 20962 10260 20995
rect 10226 20893 10260 20924
rect 10226 20890 10260 20893
rect 10226 20825 10260 20852
rect 10226 20818 10260 20825
rect 10226 20757 10260 20780
rect 10226 20746 10260 20757
rect 10226 20689 10260 20708
rect 10226 20674 10260 20689
rect 10226 20621 10260 20636
rect 10226 20602 10260 20621
rect 10226 20553 10260 20564
rect 10226 20530 10260 20553
rect 10226 20485 10260 20492
rect 10226 20458 10260 20485
rect 10226 20417 10260 20420
rect 10226 20386 10260 20417
rect 10226 20315 10260 20348
rect 10226 20314 10260 20315
rect 10226 20247 10260 20276
rect 10226 20242 10260 20247
rect 10226 20179 10260 20204
rect 10226 20170 10260 20179
rect 10226 20111 10260 20132
rect 10226 20098 10260 20111
rect 10226 20043 10260 20060
rect 10226 20026 10260 20043
rect 10226 19975 10260 19988
rect 10226 19954 10260 19975
rect 10226 19907 10260 19916
rect 10226 19882 10260 19907
rect 10226 19839 10260 19844
rect 10226 19810 10260 19839
rect 10226 19771 10260 19772
rect 10226 19738 10260 19771
rect 10226 19669 10260 19700
rect 10226 19666 10260 19669
rect 10226 19601 10260 19628
rect 10226 19594 10260 19601
rect 10226 19533 10260 19556
rect 10226 19522 10260 19533
rect 10226 19465 10260 19484
rect 10226 19450 10260 19465
rect 10226 19397 10260 19412
rect 10226 19378 10260 19397
rect 10226 19329 10260 19340
rect 10226 19306 10260 19329
rect 10226 19261 10260 19268
rect 10226 19234 10260 19261
rect 10226 19193 10260 19196
rect 10226 19162 10260 19193
rect 10226 19091 10260 19124
rect 10226 19090 10260 19091
rect 10226 19023 10260 19052
rect 10226 19018 10260 19023
rect 10226 18955 10260 18980
rect 10226 18946 10260 18955
rect 10226 18887 10260 18908
rect 10226 18874 10260 18887
rect 10226 18819 10260 18836
rect 10226 18802 10260 18819
rect 10226 18751 10260 18764
rect 10226 18730 10260 18751
rect 10226 18683 10260 18692
rect 10226 18658 10260 18683
rect 10226 18615 10260 18620
rect 10226 18586 10260 18615
rect 10226 18547 10260 18548
rect 10226 18514 10260 18547
rect 10226 18445 10260 18476
rect 10226 18442 10260 18445
rect 10226 18377 10260 18404
rect 10226 18370 10260 18377
rect 10226 18309 10260 18332
rect 10226 18298 10260 18309
rect 10226 18241 10260 18260
rect 10226 18226 10260 18241
rect 10226 18173 10260 18188
rect 10226 18154 10260 18173
rect 10226 18105 10260 18116
rect 10226 18082 10260 18105
rect 10226 18037 10260 18044
rect 10226 18010 10260 18037
rect 10226 17969 10260 17972
rect 10226 17938 10260 17969
rect 10226 17867 10260 17900
rect 10226 17866 10260 17867
rect 10226 17799 10260 17828
rect 10226 17794 10260 17799
rect 10226 17731 10260 17756
rect 10226 17722 10260 17731
rect 10226 17663 10260 17684
rect 10226 17650 10260 17663
rect 10226 17595 10260 17612
rect 10226 17578 10260 17595
rect 10226 17527 10260 17540
rect 10226 17506 10260 17527
rect 10226 17459 10260 17468
rect 10226 17434 10260 17459
rect 10226 17391 10260 17396
rect 10226 17362 10260 17391
rect 10226 17323 10260 17324
rect 10226 17290 10260 17323
rect 10226 17221 10260 17252
rect 10226 17218 10260 17221
rect 10226 17153 10260 17180
rect 10226 17146 10260 17153
rect 10226 17085 10260 17108
rect 10226 17074 10260 17085
rect 10226 17017 10260 17036
rect 10226 17002 10260 17017
rect 10226 16949 10260 16964
rect 10226 16930 10260 16949
rect 10226 16881 10260 16892
rect 10226 16858 10260 16881
rect 10226 16813 10260 16820
rect 10226 16786 10260 16813
rect 10226 16745 10260 16748
rect 10226 16714 10260 16745
rect 10226 16643 10260 16676
rect 10226 16642 10260 16643
rect 10226 16575 10260 16604
rect 10226 16570 10260 16575
rect 10226 16507 10260 16532
rect 10226 16498 10260 16507
rect 10226 16439 10260 16460
rect 10226 16426 10260 16439
rect 10226 16371 10260 16388
rect 10226 16354 10260 16371
rect 10226 16303 10260 16316
rect 10226 16282 10260 16303
rect 10226 16235 10260 16244
rect 10226 16210 10260 16235
rect 10226 16167 10260 16172
rect 10226 16138 10260 16167
rect 10226 16099 10260 16100
rect 10226 16066 10260 16099
rect 10226 15997 10260 16028
rect 10226 15994 10260 15997
rect 10226 15929 10260 15956
rect 10226 15922 10260 15929
rect 10226 15861 10260 15884
rect 10226 15850 10260 15861
rect 10226 15793 10260 15812
rect 10226 15778 10260 15793
rect 10226 15725 10260 15740
rect 10226 15706 10260 15725
rect 10226 15657 10260 15668
rect 10226 15634 10260 15657
rect 10226 15589 10260 15596
rect 10226 15562 10260 15589
rect 10226 15521 10260 15524
rect 10226 15490 10260 15521
rect 10226 15419 10260 15452
rect 10226 15418 10260 15419
rect 10226 15351 10260 15380
rect 10226 15346 10260 15351
rect 10226 15283 10260 15308
rect 10226 15274 10260 15283
rect 10226 15215 10260 15236
rect 10226 15202 10260 15215
rect 10226 15147 10260 15164
rect 10226 15130 10260 15147
rect 10226 15079 10260 15092
rect 10226 15058 10260 15079
rect 10226 15011 10260 15020
rect 10226 14986 10260 15011
rect 10226 14943 10260 14948
rect 10226 14914 10260 14943
rect 10226 14875 10260 14876
rect 10226 14842 10260 14875
rect 10226 14773 10260 14804
rect 10226 14770 10260 14773
rect 10226 14705 10260 14732
rect 10226 14698 10260 14705
rect 10226 14637 10260 14660
rect 10226 14626 10260 14637
rect 10226 14569 10260 14588
rect 10226 14554 10260 14569
rect 10226 14501 10260 14516
rect 10226 14482 10260 14501
rect 10226 14433 10260 14444
rect 10226 14410 10260 14433
rect 10226 14365 10260 14372
rect 10226 14338 10260 14365
rect 10226 14297 10260 14300
rect 10226 14266 10260 14297
rect 10226 14195 10260 14228
rect 10226 14194 10260 14195
rect 10226 14127 10260 14156
rect 10226 14122 10260 14127
rect 10226 14059 10260 14084
rect 10226 14050 10260 14059
rect 10226 13991 10260 14012
rect 10226 13978 10260 13991
rect 10226 13923 10260 13940
rect 10226 13906 10260 13923
rect 10226 13855 10260 13868
rect 10226 13834 10260 13855
rect 10226 13787 10260 13796
rect 10226 13762 10260 13787
rect 10226 13719 10260 13724
rect 10226 13690 10260 13719
rect 10226 13651 10260 13652
rect 10226 13618 10260 13651
rect 10226 13549 10260 13580
rect 10226 13546 10260 13549
rect 10226 13481 10260 13508
rect 10226 13474 10260 13481
rect 10226 13413 10260 13436
rect 10226 13402 10260 13413
rect 10226 13345 10260 13364
rect 10226 13330 10260 13345
rect 10226 13277 10260 13292
rect 10226 13258 10260 13277
rect 10226 13209 10260 13220
rect 10226 13186 10260 13209
rect 10226 13141 10260 13148
rect 10226 13114 10260 13141
rect 10226 13073 10260 13076
rect 10226 13042 10260 13073
rect 10226 12971 10260 13004
rect 10226 12970 10260 12971
rect 10226 12903 10260 12932
rect 10226 12898 10260 12903
rect 10226 12835 10260 12860
rect 10226 12826 10260 12835
rect 10226 12767 10260 12788
rect 10226 12754 10260 12767
rect 10226 12699 10260 12716
rect 10226 12682 10260 12699
rect 10226 12631 10260 12644
rect 10226 12610 10260 12631
rect 10226 12563 10260 12572
rect 10226 12538 10260 12563
rect 10226 12495 10260 12500
rect 10226 12466 10260 12495
rect 10226 12427 10260 12428
rect 10226 12394 10260 12427
rect 10226 12325 10260 12356
rect 10226 12322 10260 12325
rect 10226 12257 10260 12284
rect 10226 12250 10260 12257
rect 10226 12189 10260 12212
rect 10226 12178 10260 12189
rect 10226 12121 10260 12140
rect 10226 12106 10260 12121
rect 10226 12053 10260 12068
rect 10226 12034 10260 12053
rect 10226 11985 10260 11996
rect 10226 11962 10260 11985
rect 10226 11917 10260 11924
rect 10226 11890 10260 11917
rect 10226 11849 10260 11852
rect 10226 11818 10260 11849
rect 10226 11747 10260 11780
rect 10226 11746 10260 11747
rect 10226 11679 10260 11708
rect 10226 11674 10260 11679
rect 10226 11611 10260 11636
rect 10226 11602 10260 11611
rect 10226 11543 10260 11564
rect 10226 11530 10260 11543
rect 10226 11475 10260 11492
rect 10226 11458 10260 11475
rect 10226 11407 10260 11420
rect 10226 11386 10260 11407
rect 10226 11339 10260 11348
rect 10226 11314 10260 11339
rect 10226 11271 10260 11276
rect 10226 11242 10260 11271
rect 10226 11203 10260 11204
rect 10226 11170 10260 11203
rect 10226 11101 10260 11132
rect 10226 11098 10260 11101
rect 10226 11033 10260 11060
rect 10226 11026 10260 11033
rect 10226 10965 10260 10988
rect 10226 10954 10260 10965
rect 10226 10897 10260 10916
rect 10226 10882 10260 10897
rect 10226 10829 10260 10844
rect 10226 10810 10260 10829
rect 10226 10761 10260 10772
rect 10226 10738 10260 10761
rect 10226 10693 10260 10700
rect 10226 10666 10260 10693
rect 10226 10625 10260 10628
rect 10226 10594 10260 10625
rect 10226 10523 10260 10556
rect 10226 10522 10260 10523
rect 10226 10455 10260 10484
rect 10226 10450 10260 10455
rect 10226 10387 10260 10412
rect 10226 10378 10260 10387
rect 10226 10319 10260 10340
rect 10226 10306 10260 10319
rect 10226 10251 10260 10268
rect 10226 10234 10260 10251
rect 10226 10183 10260 10196
rect 10226 10162 10260 10183
rect 10226 10115 10260 10124
rect 10226 10090 10260 10115
rect 10226 10047 10260 10052
rect 10226 10018 10260 10047
rect 10226 9979 10260 9980
rect 10226 9946 10260 9979
rect 10226 9877 10260 9908
rect 10226 9874 10260 9877
rect 10226 9809 10260 9836
rect 10226 9802 10260 9809
rect 10226 9741 10260 9764
rect 10226 9730 10260 9741
rect 10226 9673 10260 9692
rect 10226 9658 10260 9673
rect 10226 9605 10260 9620
rect 10226 9586 10260 9605
rect 10226 9537 10260 9548
rect 10226 9514 10260 9537
rect 10226 9469 10260 9476
rect 10226 9442 10260 9469
rect 10226 9401 10260 9404
rect 10226 9370 10260 9401
rect 10226 9299 10260 9332
rect 10226 9298 10260 9299
rect 10226 9231 10260 9260
rect 10226 9226 10260 9231
rect 10226 9163 10260 9188
rect 10226 9154 10260 9163
rect 10226 9095 10260 9116
rect 10226 9082 10260 9095
rect 10226 9027 10260 9044
rect 10226 9010 10260 9027
rect 10226 8959 10260 8972
rect 10226 8938 10260 8959
rect 10226 8891 10260 8900
rect 10226 8866 10260 8891
rect 10226 8823 10260 8828
rect 10226 8794 10260 8823
rect 10226 8755 10260 8756
rect 10226 8722 10260 8755
rect 10226 8653 10260 8684
rect 10226 8650 10260 8653
rect 10226 8585 10260 8612
rect 10226 8578 10260 8585
rect 10226 8517 10260 8540
rect 10226 8506 10260 8517
rect 10226 8449 10260 8468
rect 10226 8434 10260 8449
rect 10226 8381 10260 8396
rect 10226 8362 10260 8381
rect 10226 8313 10260 8324
rect 10226 8290 10260 8313
rect 10226 8245 10260 8252
rect 10226 8218 10260 8245
rect 10226 8177 10260 8180
rect 10226 8146 10260 8177
rect 10226 8075 10260 8108
rect 10226 8074 10260 8075
rect 10226 8007 10260 8036
rect 10226 8002 10260 8007
rect 10226 7939 10260 7964
rect 10226 7930 10260 7939
rect 10226 7871 10260 7892
rect 10226 7858 10260 7871
rect 10226 7803 10260 7820
rect 10226 7786 10260 7803
rect 10226 7735 10260 7748
rect 10226 7714 10260 7735
rect 10226 7667 10260 7676
rect 10226 7642 10260 7667
rect 10226 7599 10260 7604
rect 10226 7570 10260 7599
rect 10226 7531 10260 7532
rect 10226 7498 10260 7531
rect 10226 7429 10260 7460
rect 10226 7426 10260 7429
rect 10226 7361 10260 7388
rect 10226 7354 10260 7361
rect 10226 7293 10260 7316
rect 10226 7282 10260 7293
rect 10226 7225 10260 7244
rect 10226 7210 10260 7225
rect 10226 7157 10260 7172
rect 10226 7138 10260 7157
rect 10226 7089 10260 7100
rect 10226 7066 10260 7089
rect 10226 7021 10260 7028
rect 10226 6994 10260 7021
rect 10226 6953 10260 6956
rect 10226 6922 10260 6953
rect 10226 6851 10260 6884
rect 10226 6850 10260 6851
rect 10226 6783 10260 6812
rect 10226 6778 10260 6783
rect 10226 6715 10260 6740
rect 10226 6706 10260 6715
rect 10226 6647 10260 6668
rect 10226 6634 10260 6647
rect 10226 6579 10260 6596
rect 10226 6562 10260 6579
rect 10226 6511 10260 6524
rect 10226 6490 10260 6511
rect 10226 6443 10260 6452
rect 10226 6418 10260 6443
rect 10226 6375 10260 6380
rect 10226 6346 10260 6375
rect 10226 6307 10260 6308
rect 10226 6274 10260 6307
rect 10226 6205 10260 6236
rect 10226 6202 10260 6205
rect 10226 6137 10260 6164
rect 10226 6130 10260 6137
rect 10226 6069 10260 6092
rect 10226 6058 10260 6069
rect 10226 6001 10260 6020
rect 10226 5986 10260 6001
rect 10226 5933 10260 5948
rect 10226 5914 10260 5933
rect 10226 5865 10260 5876
rect 10226 5842 10260 5865
rect 10226 5797 10260 5804
rect 10226 5770 10260 5797
rect 10226 5729 10260 5732
rect 10226 5698 10260 5729
rect 10226 5627 10260 5660
rect 10226 5626 10260 5627
rect 10226 5559 10260 5588
rect 10226 5554 10260 5559
rect 10226 5491 10260 5516
rect 10226 5482 10260 5491
rect 10226 5423 10260 5444
rect 10226 5410 10260 5423
rect 10226 5355 10260 5372
rect 10226 5338 10260 5355
rect 10226 5287 10260 5300
rect 10226 5266 10260 5287
rect 10226 5219 10260 5228
rect 10226 5194 10260 5219
rect 10226 5151 10260 5156
rect 10226 5122 10260 5151
rect 10226 5083 10260 5084
rect 10226 5050 10260 5083
rect 10226 4981 10260 5012
rect 10226 4978 10260 4981
rect 10226 4913 10260 4940
rect 10226 4906 10260 4913
rect 10226 4845 10260 4868
rect 10226 4834 10260 4845
rect 10226 4777 10260 4796
rect 10226 4762 10260 4777
rect 10226 4709 10260 4724
rect 10226 4690 10260 4709
rect 10226 4641 10260 4652
rect 10226 4618 10260 4641
rect 10226 4573 10260 4580
rect 10226 4546 10260 4573
rect 10226 4505 10260 4508
rect 10226 4474 10260 4505
rect 10226 4403 10260 4436
rect 10226 4402 10260 4403
rect 10226 4335 10260 4364
rect 10226 4330 10260 4335
rect 10226 4267 10260 4292
rect 10226 4258 10260 4267
rect 10226 4199 10260 4220
rect 10226 4186 10260 4199
rect 10226 4131 10260 4148
rect 10226 4114 10260 4131
rect 10226 4063 10260 4076
rect 10226 4042 10260 4063
rect 10226 3995 10260 4004
rect 10226 3970 10260 3995
rect 10226 3927 10260 3932
rect 10226 3898 10260 3927
rect 10226 3859 10260 3860
rect 10226 3826 10260 3859
rect 10226 3757 10260 3788
rect 10226 3754 10260 3757
rect 10226 3689 10260 3716
rect 10226 3682 10260 3689
rect 10226 3621 10260 3644
rect 10226 3610 10260 3621
rect 10226 3553 10260 3572
rect 10226 3538 10260 3553
rect 9088 3397 9122 3428
rect 9088 3394 9122 3397
rect 9214 3453 9248 3487
rect 9214 3395 9248 3415
rect 9214 3381 9248 3395
rect 9332 3453 9366 3487
rect 9332 3395 9366 3415
rect 9332 3381 9366 3395
rect 9450 3453 9484 3487
rect 9450 3395 9484 3415
rect 9450 3381 9484 3395
rect 9568 3453 9602 3487
rect 9568 3395 9602 3415
rect 9568 3381 9602 3395
rect 9686 3453 9720 3487
rect 9686 3395 9720 3415
rect 9686 3381 9720 3395
rect 9804 3453 9838 3487
rect 9804 3395 9838 3415
rect 9804 3381 9838 3395
rect 9922 3453 9956 3487
rect 9922 3395 9956 3415
rect 9922 3381 9956 3395
rect 10040 3453 10074 3487
rect 10040 3395 10074 3415
rect 10040 3381 10074 3395
rect 10226 3485 10260 3500
rect 10226 3466 10260 3485
rect 11424 38655 11458 38684
rect 11424 38650 11458 38655
rect 11424 38587 11458 38611
rect 11424 38577 11458 38587
rect 13212 38650 13246 38684
rect 12892 38581 12908 38615
rect 12908 38581 12926 38615
rect 12964 38581 12998 38615
rect 13038 38581 13060 38612
rect 13060 38581 13072 38612
rect 11424 38519 11458 38538
rect 11424 38504 11458 38519
rect 13038 38578 13072 38581
rect 11424 38451 11458 38465
rect 11424 38431 11458 38451
rect 13038 38483 13072 38517
rect 13212 38596 13246 38611
rect 13212 38577 13246 38596
rect 14940 38655 14974 38684
rect 14940 38650 14974 38655
rect 13212 38528 13246 38538
rect 13212 38504 13246 38528
rect 13392 38581 13398 38612
rect 13398 38581 13426 38612
rect 13466 38581 13500 38615
rect 13538 38581 13550 38615
rect 13550 38581 13572 38615
rect 13392 38578 13426 38581
rect 11424 38383 11458 38392
rect 11424 38358 11458 38383
rect 11424 38315 11458 38319
rect 11424 38285 11458 38315
rect 11424 38213 11458 38246
rect 11424 38212 11458 38213
rect 11424 38145 11458 38173
rect 11424 38139 11458 38145
rect 11424 38077 11458 38100
rect 11424 38066 11458 38077
rect 11424 38009 11458 38027
rect 11424 37993 11458 38009
rect 11424 37941 11458 37954
rect 11424 37920 11458 37941
rect 11424 37873 11458 37881
rect 11424 37847 11458 37873
rect 11424 37805 11458 37808
rect 11424 37774 11458 37805
rect 11424 37703 11458 37735
rect 11424 37701 11458 37703
rect 11424 37635 11458 37662
rect 11424 37628 11458 37635
rect 11424 37567 11458 37589
rect 11424 37555 11458 37567
rect 11424 37499 11458 37516
rect 11424 37482 11458 37499
rect 11424 37431 11458 37443
rect 11424 37409 11458 37431
rect 11424 37363 11458 37370
rect 11424 37336 11458 37363
rect 11424 37295 11458 37297
rect 11424 37263 11458 37295
rect 11424 37193 11458 37224
rect 11424 37190 11458 37193
rect 11424 37125 11458 37151
rect 11424 37117 11458 37125
rect 11424 37057 11458 37078
rect 11424 37044 11458 37057
rect 11424 36989 11458 37005
rect 11424 36971 11458 36989
rect 11424 36921 11458 36932
rect 11424 36898 11458 36921
rect 11424 36853 11458 36859
rect 11424 36825 11458 36853
rect 11424 36785 11458 36786
rect 11424 36752 11458 36785
rect 11424 36683 11458 36713
rect 11424 36679 11458 36683
rect 11424 36615 11458 36640
rect 11424 36606 11458 36615
rect 11424 36547 11458 36567
rect 11424 36533 11458 36547
rect 11424 36479 11458 36494
rect 11424 36460 11458 36479
rect 11424 36411 11458 36421
rect 11424 36387 11458 36411
rect 11424 36343 11458 36348
rect 11424 36314 11458 36343
rect 11424 36241 11458 36275
rect 11424 36173 11458 36202
rect 11424 36168 11458 36173
rect 11424 36105 11458 36129
rect 11424 36095 11458 36105
rect 11424 36037 11458 36056
rect 11424 36022 11458 36037
rect 11424 35969 11458 35983
rect 11424 35949 11458 35969
rect 11424 35901 11458 35910
rect 11424 35876 11458 35901
rect 11424 35833 11458 35837
rect 11424 35803 11458 35833
rect 11424 35731 11458 35764
rect 11424 35730 11458 35731
rect 11424 35663 11458 35691
rect 11424 35657 11458 35663
rect 11424 35595 11458 35618
rect 11424 35584 11458 35595
rect 11424 35527 11458 35545
rect 11424 35511 11458 35527
rect 11424 35459 11458 35472
rect 11424 35438 11458 35459
rect 11424 35391 11458 35399
rect 11424 35365 11458 35391
rect 11424 35323 11458 35326
rect 11424 35292 11458 35323
rect 11424 35221 11458 35253
rect 11424 35219 11458 35221
rect 11424 35153 11458 35180
rect 11424 35146 11458 35153
rect 11424 35085 11458 35108
rect 11424 35074 11458 35085
rect 11424 35017 11458 35036
rect 11424 35002 11458 35017
rect 11424 34949 11458 34964
rect 11424 34930 11458 34949
rect 11424 34881 11458 34892
rect 11424 34858 11458 34881
rect 11424 34813 11458 34820
rect 11424 34786 11458 34813
rect 11424 34745 11458 34748
rect 11424 34714 11458 34745
rect 11424 34643 11458 34676
rect 11424 34642 11458 34643
rect 11424 34575 11458 34604
rect 11424 34570 11458 34575
rect 11424 34507 11458 34532
rect 11424 34498 11458 34507
rect 11424 34439 11458 34460
rect 11424 34426 11458 34439
rect 11424 34371 11458 34388
rect 11424 34354 11458 34371
rect 11424 34303 11458 34316
rect 11424 34282 11458 34303
rect 11424 34235 11458 34244
rect 11424 34210 11458 34235
rect 11424 34167 11458 34172
rect 11424 34138 11458 34167
rect 11424 34099 11458 34100
rect 11424 34066 11458 34099
rect 11424 33997 11458 34028
rect 11424 33994 11458 33997
rect 11424 33929 11458 33956
rect 11424 33922 11458 33929
rect 11424 33861 11458 33884
rect 11424 33850 11458 33861
rect 11424 33793 11458 33812
rect 11424 33778 11458 33793
rect 11424 33725 11458 33740
rect 11424 33706 11458 33725
rect 11424 33657 11458 33668
rect 11424 33634 11458 33657
rect 11424 33589 11458 33596
rect 11424 33562 11458 33589
rect 11424 33521 11458 33524
rect 11424 33490 11458 33521
rect 11424 33419 11458 33452
rect 11424 33418 11458 33419
rect 11424 33351 11458 33380
rect 11424 33346 11458 33351
rect 11424 33283 11458 33308
rect 11424 33274 11458 33283
rect 11424 33215 11458 33236
rect 11424 33202 11458 33215
rect 11424 33147 11458 33164
rect 11424 33130 11458 33147
rect 11424 33079 11458 33092
rect 11424 33058 11458 33079
rect 11424 33011 11458 33020
rect 11424 32986 11458 33011
rect 11424 32943 11458 32948
rect 11424 32914 11458 32943
rect 11424 32875 11458 32876
rect 11424 32842 11458 32875
rect 11424 32773 11458 32804
rect 11424 32770 11458 32773
rect 11424 32705 11458 32732
rect 11424 32698 11458 32705
rect 11424 32637 11458 32660
rect 11424 32626 11458 32637
rect 11424 32569 11458 32588
rect 11424 32554 11458 32569
rect 11424 32501 11458 32516
rect 11424 32482 11458 32501
rect 11424 32433 11458 32444
rect 11424 32410 11458 32433
rect 11424 32365 11458 32372
rect 11424 32338 11458 32365
rect 11424 32297 11458 32300
rect 11424 32266 11458 32297
rect 11424 32195 11458 32228
rect 11424 32194 11458 32195
rect 11424 32127 11458 32156
rect 11424 32122 11458 32127
rect 11424 32059 11458 32084
rect 11424 32050 11458 32059
rect 11424 31991 11458 32012
rect 11424 31978 11458 31991
rect 11424 31923 11458 31940
rect 11424 31906 11458 31923
rect 11424 31855 11458 31868
rect 11424 31834 11458 31855
rect 11424 31787 11458 31796
rect 11424 31762 11458 31787
rect 11424 31719 11458 31724
rect 11424 31690 11458 31719
rect 11424 31651 11458 31652
rect 11424 31618 11458 31651
rect 11424 31549 11458 31580
rect 11424 31546 11458 31549
rect 11424 31481 11458 31508
rect 11424 31474 11458 31481
rect 11424 31413 11458 31436
rect 11424 31402 11458 31413
rect 11424 31345 11458 31364
rect 11424 31330 11458 31345
rect 11424 31277 11458 31292
rect 11424 31258 11458 31277
rect 11424 31209 11458 31220
rect 11424 31186 11458 31209
rect 11424 31141 11458 31148
rect 11424 31114 11458 31141
rect 11424 31073 11458 31076
rect 11424 31042 11458 31073
rect 11424 30971 11458 31004
rect 11424 30970 11458 30971
rect 11424 30903 11458 30932
rect 11424 30898 11458 30903
rect 11424 30835 11458 30860
rect 11424 30826 11458 30835
rect 11424 30767 11458 30788
rect 11424 30754 11458 30767
rect 11424 30699 11458 30716
rect 11424 30682 11458 30699
rect 11424 30631 11458 30644
rect 11424 30610 11458 30631
rect 11424 30563 11458 30572
rect 11424 30538 11458 30563
rect 11424 30495 11458 30500
rect 11424 30466 11458 30495
rect 11424 30427 11458 30428
rect 11424 30394 11458 30427
rect 11424 30325 11458 30356
rect 11424 30322 11458 30325
rect 11424 30257 11458 30284
rect 11424 30250 11458 30257
rect 11424 30189 11458 30212
rect 11424 30178 11458 30189
rect 11424 30121 11458 30140
rect 11424 30106 11458 30121
rect 11424 30053 11458 30068
rect 11424 30034 11458 30053
rect 11424 29985 11458 29996
rect 11424 29962 11458 29985
rect 11424 29917 11458 29924
rect 11424 29890 11458 29917
rect 11424 29849 11458 29852
rect 11424 29818 11458 29849
rect 11424 29747 11458 29780
rect 11424 29746 11458 29747
rect 11424 29679 11458 29708
rect 11424 29674 11458 29679
rect 11424 29611 11458 29636
rect 11424 29602 11458 29611
rect 11424 29543 11458 29564
rect 11424 29530 11458 29543
rect 11424 29475 11458 29492
rect 11424 29458 11458 29475
rect 11424 29407 11458 29420
rect 11424 29386 11458 29407
rect 11424 29339 11458 29348
rect 11424 29314 11458 29339
rect 11424 29271 11458 29276
rect 11424 29242 11458 29271
rect 11424 29203 11458 29204
rect 11424 29170 11458 29203
rect 11424 29101 11458 29132
rect 11424 29098 11458 29101
rect 11424 29033 11458 29060
rect 11424 29026 11458 29033
rect 11424 28965 11458 28988
rect 11424 28954 11458 28965
rect 11424 28897 11458 28916
rect 11424 28882 11458 28897
rect 11424 28829 11458 28844
rect 11424 28810 11458 28829
rect 11424 28761 11458 28772
rect 11424 28738 11458 28761
rect 11424 28693 11458 28700
rect 11424 28666 11458 28693
rect 11424 28625 11458 28628
rect 11424 28594 11458 28625
rect 11424 28523 11458 28556
rect 11424 28522 11458 28523
rect 11424 28455 11458 28484
rect 11424 28450 11458 28455
rect 11424 28387 11458 28412
rect 11424 28378 11458 28387
rect 11424 28319 11458 28340
rect 11424 28306 11458 28319
rect 11424 28251 11458 28268
rect 11424 28234 11458 28251
rect 11424 28183 11458 28196
rect 11424 28162 11458 28183
rect 11424 28115 11458 28124
rect 11424 28090 11458 28115
rect 11424 28047 11458 28052
rect 11424 28018 11458 28047
rect 11424 27979 11458 27980
rect 11424 27946 11458 27979
rect 11424 27877 11458 27908
rect 11424 27874 11458 27877
rect 11424 27809 11458 27836
rect 11424 27802 11458 27809
rect 11424 27741 11458 27764
rect 11424 27730 11458 27741
rect 11424 27673 11458 27692
rect 11424 27658 11458 27673
rect 11424 27605 11458 27620
rect 11424 27586 11458 27605
rect 11424 27537 11458 27548
rect 11424 27514 11458 27537
rect 11424 27469 11458 27476
rect 11424 27442 11458 27469
rect 11424 27401 11458 27404
rect 11424 27370 11458 27401
rect 11424 27299 11458 27332
rect 11424 27298 11458 27299
rect 11424 27231 11458 27260
rect 11424 27226 11458 27231
rect 11424 27163 11458 27188
rect 11424 27154 11458 27163
rect 11424 27095 11458 27116
rect 11424 27082 11458 27095
rect 11424 27027 11458 27044
rect 11424 27010 11458 27027
rect 11424 26959 11458 26972
rect 11424 26938 11458 26959
rect 11424 26891 11458 26900
rect 11424 26866 11458 26891
rect 11424 26823 11458 26828
rect 11424 26794 11458 26823
rect 11424 26755 11458 26756
rect 11424 26722 11458 26755
rect 11424 26653 11458 26684
rect 11424 26650 11458 26653
rect 11424 26585 11458 26612
rect 11424 26578 11458 26585
rect 11424 26517 11458 26540
rect 11424 26506 11458 26517
rect 11424 26449 11458 26468
rect 11424 26434 11458 26449
rect 11424 26381 11458 26396
rect 11424 26362 11458 26381
rect 11424 26313 11458 26324
rect 11424 26290 11458 26313
rect 11424 26245 11458 26252
rect 11424 26218 11458 26245
rect 11424 26177 11458 26180
rect 11424 26146 11458 26177
rect 11424 26075 11458 26108
rect 11424 26074 11458 26075
rect 11424 26007 11458 26036
rect 11424 26002 11458 26007
rect 11424 25939 11458 25964
rect 11424 25930 11458 25939
rect 11424 25871 11458 25892
rect 11424 25858 11458 25871
rect 11424 25803 11458 25820
rect 11424 25786 11458 25803
rect 11424 25735 11458 25748
rect 11424 25714 11458 25735
rect 11424 25667 11458 25676
rect 11424 25642 11458 25667
rect 11424 25599 11458 25604
rect 11424 25570 11458 25599
rect 11424 25531 11458 25532
rect 11424 25498 11458 25531
rect 11424 25429 11458 25460
rect 11424 25426 11458 25429
rect 11424 25361 11458 25388
rect 11424 25354 11458 25361
rect 11424 25293 11458 25316
rect 11424 25282 11458 25293
rect 11424 25225 11458 25244
rect 11424 25210 11458 25225
rect 11424 25157 11458 25172
rect 11424 25138 11458 25157
rect 11424 25089 11458 25100
rect 11424 25066 11458 25089
rect 11424 25021 11458 25028
rect 11424 24994 11458 25021
rect 11424 24953 11458 24956
rect 11424 24922 11458 24953
rect 11424 24851 11458 24884
rect 11424 24850 11458 24851
rect 11424 24783 11458 24812
rect 11424 24778 11458 24783
rect 11424 24715 11458 24740
rect 11424 24706 11458 24715
rect 11424 24647 11458 24668
rect 11424 24634 11458 24647
rect 11424 24579 11458 24596
rect 11424 24562 11458 24579
rect 11424 24511 11458 24524
rect 11424 24490 11458 24511
rect 11424 24443 11458 24452
rect 11424 24418 11458 24443
rect 11424 24375 11458 24380
rect 11424 24346 11458 24375
rect 11424 24307 11458 24308
rect 11424 24274 11458 24307
rect 11424 24205 11458 24236
rect 11424 24202 11458 24205
rect 11424 24137 11458 24164
rect 11424 24130 11458 24137
rect 11424 24069 11458 24092
rect 11424 24058 11458 24069
rect 11424 24001 11458 24020
rect 11424 23986 11458 24001
rect 11424 23933 11458 23948
rect 11424 23914 11458 23933
rect 11424 23865 11458 23876
rect 11424 23842 11458 23865
rect 11424 23797 11458 23804
rect 11424 23770 11458 23797
rect 11424 23729 11458 23732
rect 11424 23698 11458 23729
rect 11424 23627 11458 23660
rect 11424 23626 11458 23627
rect 11424 23559 11458 23588
rect 11424 23554 11458 23559
rect 11424 23491 11458 23516
rect 11424 23482 11458 23491
rect 11424 23423 11458 23444
rect 11424 23410 11458 23423
rect 11424 23355 11458 23372
rect 11424 23338 11458 23355
rect 11424 23287 11458 23300
rect 11424 23266 11458 23287
rect 11424 23219 11458 23228
rect 11424 23194 11458 23219
rect 11424 23151 11458 23156
rect 11424 23122 11458 23151
rect 11424 23083 11458 23084
rect 11424 23050 11458 23083
rect 11424 22981 11458 23012
rect 11424 22978 11458 22981
rect 11424 22913 11458 22940
rect 11424 22906 11458 22913
rect 11424 22845 11458 22868
rect 11424 22834 11458 22845
rect 11424 22777 11458 22796
rect 11424 22762 11458 22777
rect 11424 22709 11458 22724
rect 11424 22690 11458 22709
rect 11424 22641 11458 22652
rect 11424 22618 11458 22641
rect 11424 22573 11458 22580
rect 11424 22546 11458 22573
rect 11424 22505 11458 22508
rect 11424 22474 11458 22505
rect 11424 22403 11458 22436
rect 11424 22402 11458 22403
rect 11424 22335 11458 22364
rect 11424 22330 11458 22335
rect 11424 22267 11458 22292
rect 11424 22258 11458 22267
rect 11424 22199 11458 22220
rect 11424 22186 11458 22199
rect 11424 22131 11458 22148
rect 11424 22114 11458 22131
rect 11424 22063 11458 22076
rect 11424 22042 11458 22063
rect 11424 21995 11458 22004
rect 11424 21970 11458 21995
rect 11424 21927 11458 21932
rect 11424 21898 11458 21927
rect 11424 21859 11458 21860
rect 11424 21826 11458 21859
rect 11424 21757 11458 21788
rect 11424 21754 11458 21757
rect 11424 21689 11458 21716
rect 11424 21682 11458 21689
rect 11424 21621 11458 21644
rect 11424 21610 11458 21621
rect 11424 21553 11458 21572
rect 11424 21538 11458 21553
rect 11424 21485 11458 21500
rect 11424 21466 11458 21485
rect 11424 21417 11458 21428
rect 11424 21394 11458 21417
rect 11424 21349 11458 21356
rect 11424 21322 11458 21349
rect 11424 21281 11458 21284
rect 11424 21250 11458 21281
rect 11424 21179 11458 21212
rect 11424 21178 11458 21179
rect 11424 21111 11458 21140
rect 11424 21106 11458 21111
rect 11424 21043 11458 21068
rect 11424 21034 11458 21043
rect 11424 20975 11458 20996
rect 11424 20962 11458 20975
rect 11424 20907 11458 20924
rect 11424 20890 11458 20907
rect 11424 20839 11458 20852
rect 11424 20818 11458 20839
rect 11424 20771 11458 20780
rect 11424 20746 11458 20771
rect 11424 20703 11458 20708
rect 11424 20674 11458 20703
rect 11424 20635 11458 20636
rect 11424 20602 11458 20635
rect 11424 20533 11458 20564
rect 11424 20530 11458 20533
rect 11424 20465 11458 20492
rect 11424 20458 11458 20465
rect 11424 20397 11458 20420
rect 11424 20386 11458 20397
rect 11424 20329 11458 20348
rect 11424 20314 11458 20329
rect 11424 20261 11458 20276
rect 11424 20242 11458 20261
rect 11424 20193 11458 20204
rect 11424 20170 11458 20193
rect 11424 20125 11458 20132
rect 11424 20098 11458 20125
rect 11424 20057 11458 20060
rect 11424 20026 11458 20057
rect 11424 19955 11458 19988
rect 11424 19954 11458 19955
rect 11424 19887 11458 19916
rect 11424 19882 11458 19887
rect 11424 19819 11458 19844
rect 11424 19810 11458 19819
rect 11424 19751 11458 19772
rect 11424 19738 11458 19751
rect 11424 19683 11458 19700
rect 11424 19666 11458 19683
rect 11424 19615 11458 19628
rect 11424 19594 11458 19615
rect 11424 19547 11458 19556
rect 11424 19522 11458 19547
rect 11424 19479 11458 19484
rect 11424 19450 11458 19479
rect 11424 19411 11458 19412
rect 11424 19378 11458 19411
rect 11424 19309 11458 19340
rect 11424 19306 11458 19309
rect 11424 19241 11458 19268
rect 11424 19234 11458 19241
rect 11424 19173 11458 19196
rect 11424 19162 11458 19173
rect 11424 19105 11458 19124
rect 11424 19090 11458 19105
rect 11424 19037 11458 19052
rect 11424 19018 11458 19037
rect 11424 18969 11458 18980
rect 11424 18946 11458 18969
rect 11424 18901 11458 18908
rect 11424 18874 11458 18901
rect 11424 18833 11458 18836
rect 11424 18802 11458 18833
rect 11424 18731 11458 18764
rect 11424 18730 11458 18731
rect 11424 18663 11458 18692
rect 11424 18658 11458 18663
rect 11424 18595 11458 18620
rect 11424 18586 11458 18595
rect 11424 18527 11458 18548
rect 11424 18514 11458 18527
rect 11424 18459 11458 18476
rect 11424 18442 11458 18459
rect 11424 18391 11458 18404
rect 11424 18370 11458 18391
rect 11424 18323 11458 18332
rect 11424 18298 11458 18323
rect 11424 18255 11458 18260
rect 11424 18226 11458 18255
rect 11424 18187 11458 18188
rect 11424 18154 11458 18187
rect 11424 18085 11458 18116
rect 11424 18082 11458 18085
rect 11424 18017 11458 18044
rect 11424 18010 11458 18017
rect 11424 17949 11458 17972
rect 11424 17938 11458 17949
rect 11424 17881 11458 17900
rect 11424 17866 11458 17881
rect 11424 17813 11458 17828
rect 11424 17794 11458 17813
rect 11424 17745 11458 17756
rect 11424 17722 11458 17745
rect 11424 17677 11458 17684
rect 11424 17650 11458 17677
rect 11424 17609 11458 17612
rect 11424 17578 11458 17609
rect 11424 17507 11458 17540
rect 11424 17506 11458 17507
rect 11424 17439 11458 17468
rect 11424 17434 11458 17439
rect 11424 17371 11458 17396
rect 11424 17362 11458 17371
rect 11424 17303 11458 17324
rect 11424 17290 11458 17303
rect 11424 17235 11458 17252
rect 11424 17218 11458 17235
rect 11424 17167 11458 17180
rect 11424 17146 11458 17167
rect 11424 17099 11458 17108
rect 11424 17074 11458 17099
rect 11424 17031 11458 17036
rect 11424 17002 11458 17031
rect 11424 16963 11458 16964
rect 11424 16930 11458 16963
rect 11424 16861 11458 16892
rect 11424 16858 11458 16861
rect 11424 16793 11458 16820
rect 11424 16786 11458 16793
rect 11424 16725 11458 16748
rect 11424 16714 11458 16725
rect 11424 16657 11458 16676
rect 11424 16642 11458 16657
rect 11424 16589 11458 16604
rect 11424 16570 11458 16589
rect 11424 16521 11458 16532
rect 11424 16498 11458 16521
rect 11424 16453 11458 16460
rect 11424 16426 11458 16453
rect 11424 16385 11458 16388
rect 11424 16354 11458 16385
rect 11424 16283 11458 16316
rect 11424 16282 11458 16283
rect 11424 16215 11458 16244
rect 11424 16210 11458 16215
rect 11424 16147 11458 16172
rect 11424 16138 11458 16147
rect 11424 16079 11458 16100
rect 11424 16066 11458 16079
rect 11424 16011 11458 16028
rect 11424 15994 11458 16011
rect 11424 15943 11458 15956
rect 11424 15922 11458 15943
rect 11424 15875 11458 15884
rect 11424 15850 11458 15875
rect 11424 15807 11458 15812
rect 11424 15778 11458 15807
rect 11424 15739 11458 15740
rect 11424 15706 11458 15739
rect 11424 15637 11458 15668
rect 11424 15634 11458 15637
rect 11424 15569 11458 15596
rect 11424 15562 11458 15569
rect 11424 15501 11458 15524
rect 11424 15490 11458 15501
rect 11424 15433 11458 15452
rect 11424 15418 11458 15433
rect 11424 15365 11458 15380
rect 11424 15346 11458 15365
rect 11424 15297 11458 15308
rect 11424 15274 11458 15297
rect 11424 15229 11458 15236
rect 11424 15202 11458 15229
rect 11424 15161 11458 15164
rect 11424 15130 11458 15161
rect 11424 15059 11458 15092
rect 11424 15058 11458 15059
rect 11424 14991 11458 15020
rect 11424 14986 11458 14991
rect 11424 14923 11458 14948
rect 11424 14914 11458 14923
rect 11424 14855 11458 14876
rect 11424 14842 11458 14855
rect 11424 14787 11458 14804
rect 11424 14770 11458 14787
rect 11424 14719 11458 14732
rect 11424 14698 11458 14719
rect 11424 14651 11458 14660
rect 11424 14626 11458 14651
rect 11424 14583 11458 14588
rect 11424 14554 11458 14583
rect 11424 14515 11458 14516
rect 11424 14482 11458 14515
rect 11424 14413 11458 14444
rect 11424 14410 11458 14413
rect 11424 14345 11458 14372
rect 11424 14338 11458 14345
rect 11424 14277 11458 14300
rect 11424 14266 11458 14277
rect 11424 14209 11458 14228
rect 11424 14194 11458 14209
rect 11424 14141 11458 14156
rect 11424 14122 11458 14141
rect 11424 14073 11458 14084
rect 11424 14050 11458 14073
rect 11424 14005 11458 14012
rect 11424 13978 11458 14005
rect 11424 13937 11458 13940
rect 11424 13906 11458 13937
rect 11424 13835 11458 13868
rect 11424 13834 11458 13835
rect 11424 13767 11458 13796
rect 11424 13762 11458 13767
rect 11424 13699 11458 13724
rect 11424 13690 11458 13699
rect 11424 13631 11458 13652
rect 11424 13618 11458 13631
rect 11424 13563 11458 13580
rect 11424 13546 11458 13563
rect 11424 13495 11458 13508
rect 11424 13474 11458 13495
rect 11424 13427 11458 13436
rect 11424 13402 11458 13427
rect 11424 13359 11458 13364
rect 11424 13330 11458 13359
rect 11424 13291 11458 13292
rect 11424 13258 11458 13291
rect 11424 13189 11458 13220
rect 11424 13186 11458 13189
rect 11424 13121 11458 13148
rect 11424 13114 11458 13121
rect 11424 13053 11458 13076
rect 11424 13042 11458 13053
rect 11424 12985 11458 13004
rect 11424 12970 11458 12985
rect 11424 12917 11458 12932
rect 11424 12898 11458 12917
rect 11424 12849 11458 12860
rect 11424 12826 11458 12849
rect 11424 12781 11458 12788
rect 11424 12754 11458 12781
rect 11424 12713 11458 12716
rect 11424 12682 11458 12713
rect 11424 12611 11458 12644
rect 11424 12610 11458 12611
rect 11424 12543 11458 12572
rect 11424 12538 11458 12543
rect 11424 12475 11458 12500
rect 11424 12466 11458 12475
rect 11424 12407 11458 12428
rect 11424 12394 11458 12407
rect 11424 12339 11458 12356
rect 11424 12322 11458 12339
rect 11424 12271 11458 12284
rect 11424 12250 11458 12271
rect 11424 12203 11458 12212
rect 11424 12178 11458 12203
rect 11424 12135 11458 12140
rect 11424 12106 11458 12135
rect 11424 12067 11458 12068
rect 11424 12034 11458 12067
rect 11424 11965 11458 11996
rect 11424 11962 11458 11965
rect 11424 11897 11458 11924
rect 11424 11890 11458 11897
rect 11424 11829 11458 11852
rect 11424 11818 11458 11829
rect 11424 11761 11458 11780
rect 11424 11746 11458 11761
rect 11424 11693 11458 11708
rect 11424 11674 11458 11693
rect 11424 11625 11458 11636
rect 11424 11602 11458 11625
rect 11424 11557 11458 11564
rect 11424 11530 11458 11557
rect 11424 11489 11458 11492
rect 11424 11458 11458 11489
rect 11424 11387 11458 11420
rect 11424 11386 11458 11387
rect 11424 11319 11458 11348
rect 11424 11314 11458 11319
rect 11424 11251 11458 11276
rect 11424 11242 11458 11251
rect 11424 11183 11458 11204
rect 11424 11170 11458 11183
rect 11424 11115 11458 11132
rect 11424 11098 11458 11115
rect 11424 11047 11458 11060
rect 11424 11026 11458 11047
rect 11424 10979 11458 10988
rect 11424 10954 11458 10979
rect 11424 10911 11458 10916
rect 11424 10882 11458 10911
rect 11424 10843 11458 10844
rect 11424 10810 11458 10843
rect 11424 10741 11458 10772
rect 11424 10738 11458 10741
rect 11424 10673 11458 10700
rect 11424 10666 11458 10673
rect 11424 10605 11458 10628
rect 11424 10594 11458 10605
rect 11424 10537 11458 10556
rect 11424 10522 11458 10537
rect 11424 10469 11458 10484
rect 11424 10450 11458 10469
rect 11424 10401 11458 10412
rect 11424 10378 11458 10401
rect 11424 10333 11458 10340
rect 11424 10306 11458 10333
rect 11424 10265 11458 10268
rect 11424 10234 11458 10265
rect 11424 10163 11458 10196
rect 11424 10162 11458 10163
rect 11424 10095 11458 10124
rect 11424 10090 11458 10095
rect 11424 10027 11458 10052
rect 11424 10018 11458 10027
rect 11424 9959 11458 9980
rect 11424 9946 11458 9959
rect 11424 9891 11458 9908
rect 11424 9874 11458 9891
rect 11424 9823 11458 9836
rect 11424 9802 11458 9823
rect 11424 9755 11458 9764
rect 11424 9730 11458 9755
rect 11424 9687 11458 9692
rect 11424 9658 11458 9687
rect 11424 9619 11458 9620
rect 11424 9586 11458 9619
rect 11424 9517 11458 9548
rect 11424 9514 11458 9517
rect 11424 9449 11458 9476
rect 11424 9442 11458 9449
rect 11424 9381 11458 9404
rect 11424 9370 11458 9381
rect 11424 9313 11458 9332
rect 11424 9298 11458 9313
rect 11424 9245 11458 9260
rect 11424 9226 11458 9245
rect 11424 9177 11458 9188
rect 11424 9154 11458 9177
rect 11424 9109 11458 9116
rect 11424 9082 11458 9109
rect 11424 9041 11458 9044
rect 11424 9010 11458 9041
rect 11424 8939 11458 8972
rect 11424 8938 11458 8939
rect 11424 8871 11458 8900
rect 11424 8866 11458 8871
rect 11424 8803 11458 8828
rect 11424 8794 11458 8803
rect 11424 8735 11458 8756
rect 11424 8722 11458 8735
rect 11424 8667 11458 8684
rect 11424 8650 11458 8667
rect 11424 8599 11458 8612
rect 11424 8578 11458 8599
rect 11424 8531 11458 8540
rect 11424 8506 11458 8531
rect 11424 8463 11458 8468
rect 11424 8434 11458 8463
rect 11424 8395 11458 8396
rect 11424 8362 11458 8395
rect 11424 8293 11458 8324
rect 11424 8290 11458 8293
rect 11424 8225 11458 8252
rect 11424 8218 11458 8225
rect 11424 8157 11458 8180
rect 11424 8146 11458 8157
rect 11424 8089 11458 8108
rect 11424 8074 11458 8089
rect 11424 8021 11458 8036
rect 11424 8002 11458 8021
rect 11424 7953 11458 7964
rect 11424 7930 11458 7953
rect 11424 7885 11458 7892
rect 11424 7858 11458 7885
rect 11424 7817 11458 7820
rect 11424 7786 11458 7817
rect 11424 7715 11458 7748
rect 11424 7714 11458 7715
rect 11424 7647 11458 7676
rect 11424 7642 11458 7647
rect 11424 7579 11458 7604
rect 11424 7570 11458 7579
rect 11424 7511 11458 7532
rect 11424 7498 11458 7511
rect 11424 7443 11458 7460
rect 11424 7426 11458 7443
rect 11424 7375 11458 7388
rect 11424 7354 11458 7375
rect 11424 7307 11458 7316
rect 11424 7282 11458 7307
rect 11424 7239 11458 7244
rect 11424 7210 11458 7239
rect 11424 7171 11458 7172
rect 11424 7138 11458 7171
rect 11424 7069 11458 7100
rect 11424 7066 11458 7069
rect 11424 7001 11458 7028
rect 11424 6994 11458 7001
rect 11424 6933 11458 6956
rect 11424 6922 11458 6933
rect 11424 6865 11458 6884
rect 11424 6850 11458 6865
rect 11424 6797 11458 6812
rect 11424 6778 11458 6797
rect 11424 6729 11458 6740
rect 11424 6706 11458 6729
rect 11424 6661 11458 6668
rect 11424 6634 11458 6661
rect 11424 6593 11458 6596
rect 11424 6562 11458 6593
rect 11424 6491 11458 6524
rect 11424 6490 11458 6491
rect 11424 6423 11458 6452
rect 11424 6418 11458 6423
rect 11424 6355 11458 6380
rect 11424 6346 11458 6355
rect 11424 6287 11458 6308
rect 11424 6274 11458 6287
rect 11424 6219 11458 6236
rect 11424 6202 11458 6219
rect 11424 6151 11458 6164
rect 11424 6130 11458 6151
rect 11424 6083 11458 6092
rect 11424 6058 11458 6083
rect 11424 6015 11458 6020
rect 11424 5986 11458 6015
rect 11424 5947 11458 5948
rect 11424 5914 11458 5947
rect 11424 5845 11458 5876
rect 11424 5842 11458 5845
rect 11424 5777 11458 5804
rect 11424 5770 11458 5777
rect 11424 5709 11458 5732
rect 11424 5698 11458 5709
rect 11424 5641 11458 5660
rect 11424 5626 11458 5641
rect 11424 5573 11458 5588
rect 11424 5554 11458 5573
rect 11424 5505 11458 5516
rect 11424 5482 11458 5505
rect 11424 5437 11458 5444
rect 11424 5410 11458 5437
rect 11424 5369 11458 5372
rect 11424 5338 11458 5369
rect 11424 5267 11458 5300
rect 11424 5266 11458 5267
rect 11424 5199 11458 5228
rect 11424 5194 11458 5199
rect 11424 5131 11458 5156
rect 11424 5122 11458 5131
rect 11424 5063 11458 5084
rect 11424 5050 11458 5063
rect 11424 4995 11458 5012
rect 11424 4978 11458 4995
rect 11424 4927 11458 4940
rect 11424 4906 11458 4927
rect 11424 4859 11458 4868
rect 11424 4834 11458 4859
rect 11424 4791 11458 4796
rect 11424 4762 11458 4791
rect 11424 4723 11458 4724
rect 11424 4690 11458 4723
rect 11424 4621 11458 4652
rect 11424 4618 11458 4621
rect 11424 4553 11458 4580
rect 11424 4546 11458 4553
rect 11424 4485 11458 4508
rect 11424 4474 11458 4485
rect 11424 4417 11458 4436
rect 11424 4402 11458 4417
rect 11424 4349 11458 4364
rect 11424 4330 11458 4349
rect 11424 4281 11458 4292
rect 11424 4258 11458 4281
rect 11424 4213 11458 4220
rect 11424 4186 11458 4213
rect 11424 4145 11458 4148
rect 11424 4114 11458 4145
rect 11424 4043 11458 4076
rect 11424 4042 11458 4043
rect 11424 3975 11458 4004
rect 11424 3970 11458 3975
rect 11424 3907 11458 3932
rect 11424 3898 11458 3907
rect 11424 3839 11458 3860
rect 11424 3826 11458 3839
rect 11424 3771 11458 3788
rect 11424 3754 11458 3771
rect 11424 3703 11458 3716
rect 11424 3682 11458 3703
rect 11424 3635 11458 3644
rect 11424 3610 11458 3635
rect 11424 3567 11458 3572
rect 11424 3538 11458 3567
rect 10226 3417 10260 3428
rect 10226 3394 10260 3417
rect 9088 3329 9122 3356
rect 9088 3322 9122 3329
rect 9088 3250 9122 3284
rect 10412 3453 10446 3487
rect 10412 3395 10446 3415
rect 10412 3381 10446 3395
rect 10530 3453 10564 3487
rect 10530 3395 10564 3415
rect 10530 3381 10564 3395
rect 10648 3453 10682 3487
rect 10648 3395 10682 3415
rect 10648 3381 10682 3395
rect 10766 3453 10800 3487
rect 10766 3395 10800 3415
rect 10766 3381 10800 3395
rect 10884 3453 10918 3487
rect 10884 3395 10918 3415
rect 10884 3381 10918 3395
rect 11002 3453 11036 3487
rect 11002 3395 11036 3415
rect 11002 3381 11036 3395
rect 11120 3453 11154 3487
rect 11120 3395 11154 3415
rect 11120 3381 11154 3395
rect 11238 3453 11272 3487
rect 11238 3395 11272 3415
rect 11238 3381 11272 3395
rect 11424 3499 11458 3500
rect 11424 3466 11458 3499
rect 11424 3397 11458 3428
rect 11424 3394 11458 3397
rect 10226 3349 10260 3356
rect 10226 3322 10260 3349
rect 10226 3281 10260 3284
rect 10226 3250 10260 3281
rect 11424 3329 11458 3356
rect 11424 3322 11458 3329
rect 11424 3250 11458 3284
rect 9160 3179 9190 3212
rect 9190 3179 9194 3212
rect 9234 3179 9258 3212
rect 9258 3179 9268 3212
rect 9307 3179 9326 3212
rect 9326 3179 9341 3212
rect 9380 3179 9394 3212
rect 9394 3179 9414 3212
rect 9453 3179 9462 3212
rect 9462 3179 9487 3212
rect 9526 3179 9530 3212
rect 9530 3179 9560 3212
rect 9599 3179 9632 3212
rect 9632 3179 9633 3212
rect 9672 3179 9700 3212
rect 9700 3179 9706 3212
rect 9745 3179 9768 3212
rect 9768 3179 9779 3212
rect 9818 3179 9836 3212
rect 9836 3179 9852 3212
rect 9891 3179 9904 3212
rect 9904 3179 9925 3212
rect 9964 3179 9972 3212
rect 9972 3179 9998 3212
rect 10037 3179 10040 3212
rect 10040 3179 10071 3212
rect 10110 3179 10142 3212
rect 10142 3179 10144 3212
rect 9160 3178 9194 3179
rect 9234 3178 9268 3179
rect 9307 3178 9341 3179
rect 9380 3178 9414 3179
rect 9453 3178 9487 3179
rect 9526 3178 9560 3179
rect 9599 3178 9633 3179
rect 9672 3178 9706 3179
rect 9745 3178 9779 3179
rect 9818 3178 9852 3179
rect 9891 3178 9925 3179
rect 9964 3178 9998 3179
rect 10037 3178 10071 3179
rect 10110 3178 10144 3179
rect 10183 3178 10217 3212
rect 10256 3178 10290 3212
rect 10329 3179 10336 3212
rect 10336 3179 10363 3212
rect 10402 3179 10404 3212
rect 10404 3179 10436 3212
rect 10475 3179 10506 3212
rect 10506 3179 10509 3212
rect 10548 3179 10574 3212
rect 10574 3179 10582 3212
rect 10621 3179 10642 3212
rect 10642 3179 10655 3212
rect 10694 3179 10710 3212
rect 10710 3179 10728 3212
rect 10767 3179 10778 3212
rect 10778 3179 10801 3212
rect 10840 3179 10846 3212
rect 10846 3179 10874 3212
rect 10913 3179 10914 3212
rect 10914 3179 10947 3212
rect 10986 3179 11016 3212
rect 11016 3179 11020 3212
rect 11059 3179 11084 3212
rect 11084 3179 11093 3212
rect 11132 3179 11152 3212
rect 11152 3179 11166 3212
rect 11205 3179 11220 3212
rect 11220 3179 11239 3212
rect 11278 3179 11288 3212
rect 11288 3179 11312 3212
rect 11351 3179 11356 3212
rect 11356 3179 11385 3212
rect 10329 3178 10363 3179
rect 10402 3178 10436 3179
rect 10475 3178 10509 3179
rect 10548 3178 10582 3179
rect 10621 3178 10655 3179
rect 10694 3178 10728 3179
rect 10767 3178 10801 3179
rect 10840 3178 10874 3179
rect 10913 3178 10947 3179
rect 10986 3178 11020 3179
rect 11059 3178 11093 3179
rect 11132 3178 11166 3179
rect 11205 3178 11239 3179
rect 11278 3178 11312 3179
rect 11351 3178 11385 3179
rect 11424 3137 11458 3140
rect 11424 3106 11458 3137
rect 11424 3035 11458 3067
rect 11424 3033 11458 3035
rect 11424 2967 11458 2994
rect 11424 2960 11458 2967
rect 11424 2899 11458 2921
rect 11424 2887 11458 2899
rect 11424 2831 11458 2848
rect 11424 2814 11458 2831
rect 11424 2763 11458 2775
rect 11424 2741 11458 2763
rect 11424 2695 11458 2702
rect 11424 2668 11458 2695
rect 5418 2561 5452 2595
rect 5500 2561 5534 2595
rect 5583 2561 5617 2595
rect 5666 2561 5700 2595
rect 5749 2561 5783 2595
rect 5832 2561 5866 2595
rect 5940 2568 5974 2589
rect 5940 2555 5974 2568
rect 5184 2534 5218 2549
rect 5184 2515 5218 2534
rect 5184 2465 5218 2476
rect 5184 2442 5218 2465
rect 5940 2500 5974 2515
rect 5940 2481 5974 2500
rect 5278 2405 5312 2439
rect 5357 2405 5391 2439
rect 5436 2405 5470 2439
rect 5515 2405 5549 2439
rect 5595 2405 5629 2439
rect 5675 2405 5709 2439
rect 5755 2405 5789 2439
rect 5940 2432 5974 2441
rect 5940 2407 5974 2432
rect 5184 2396 5218 2403
rect 5184 2369 5218 2396
rect 5184 2327 5218 2330
rect 5184 2296 5218 2327
rect 5940 2364 5974 2367
rect 5940 2333 5974 2364
rect 5184 2224 5218 2257
rect 5418 2249 5452 2283
rect 5500 2249 5534 2283
rect 5583 2249 5617 2283
rect 5666 2249 5700 2283
rect 5749 2249 5783 2283
rect 5832 2249 5866 2283
rect 5940 2262 5974 2293
rect 5940 2259 5974 2262
rect 5184 2223 5218 2224
rect 5184 2155 5218 2184
rect 5184 2150 5218 2155
rect 5940 2194 5974 2219
rect 5940 2185 5974 2194
rect 5184 2086 5218 2111
rect 5278 2093 5312 2127
rect 5357 2093 5391 2127
rect 5436 2093 5470 2127
rect 5515 2093 5549 2127
rect 5595 2093 5629 2127
rect 5675 2093 5709 2127
rect 5755 2093 5789 2127
rect 5940 2126 5974 2145
rect 5940 2111 5974 2126
rect 5184 2077 5218 2086
rect 5184 2017 5218 2038
rect 5184 2004 5218 2017
rect 5940 2058 5974 2071
rect 5940 2037 5974 2058
rect 5940 1990 5974 1997
rect 5184 1948 5218 1965
rect 5184 1931 5218 1948
rect 5418 1937 5452 1971
rect 5500 1937 5534 1971
rect 5583 1937 5617 1971
rect 5666 1937 5700 1971
rect 5749 1937 5783 1971
rect 5832 1937 5866 1971
rect 5940 1963 5974 1990
rect 5184 1879 5218 1892
rect 5184 1858 5218 1879
rect 5184 1810 5218 1819
rect 5940 1922 5974 1923
rect 5940 1889 5974 1922
rect 5940 1820 5974 1849
rect 5940 1815 5974 1820
rect 5184 1785 5218 1810
rect 5278 1781 5312 1815
rect 5357 1781 5391 1815
rect 5436 1781 5470 1815
rect 5515 1781 5549 1815
rect 5595 1781 5629 1815
rect 5675 1781 5709 1815
rect 5755 1781 5789 1815
rect 5184 1742 5218 1746
rect 5184 1712 5218 1742
rect 5184 1640 5218 1673
rect 5940 1752 5974 1775
rect 5940 1741 5974 1752
rect 5940 1684 5974 1701
rect 5940 1667 5974 1684
rect 5184 1639 5218 1640
rect 5418 1625 5452 1659
rect 5500 1625 5534 1659
rect 5583 1625 5617 1659
rect 5666 1625 5700 1659
rect 5749 1625 5783 1659
rect 5832 1625 5866 1659
rect 5184 1572 5218 1600
rect 5184 1566 5218 1572
rect 5184 1504 5218 1527
rect 5184 1493 5218 1504
rect 5940 1616 5974 1627
rect 5940 1593 5974 1616
rect 5940 1548 5974 1553
rect 5940 1519 5974 1548
rect 5278 1469 5312 1503
rect 5357 1469 5391 1503
rect 5436 1469 5470 1503
rect 5515 1469 5549 1503
rect 5595 1469 5629 1503
rect 5675 1469 5709 1503
rect 5755 1469 5789 1503
rect 5184 1436 5218 1454
rect 5184 1420 5218 1436
rect 5184 1368 5218 1381
rect 5184 1347 5218 1368
rect 5940 1446 5974 1479
rect 5940 1445 5974 1446
rect 5940 1378 5974 1406
rect 5940 1372 5974 1378
rect 5418 1313 5452 1347
rect 5500 1313 5534 1347
rect 5583 1313 5617 1347
rect 5666 1313 5700 1347
rect 5749 1313 5783 1347
rect 5832 1313 5866 1347
rect 5184 1300 5218 1308
rect 5184 1274 5218 1300
rect 5184 1232 5218 1236
rect 5184 1202 5218 1232
rect 5940 1310 5974 1333
rect 5940 1299 5974 1310
rect 5940 1242 5974 1260
rect 5940 1226 5974 1242
rect 5184 1130 5218 1164
rect 5278 1157 5312 1191
rect 5357 1157 5391 1191
rect 5436 1157 5470 1191
rect 5515 1157 5549 1191
rect 5595 1157 5629 1191
rect 5675 1157 5709 1191
rect 5755 1157 5789 1191
rect 5940 1174 5974 1187
rect 5184 1062 5218 1092
rect 5184 1058 5218 1062
rect 5940 1153 5974 1174
rect 5940 1106 5974 1114
rect 5940 1080 5974 1106
rect 5940 1038 5974 1041
rect 5418 1001 5452 1035
rect 5500 1001 5534 1035
rect 5583 1001 5617 1035
rect 5666 1001 5700 1035
rect 5749 1001 5783 1035
rect 5832 1001 5866 1035
rect 5940 1007 5974 1038
rect 11424 2627 11458 2629
rect 11424 2595 11458 2627
rect 11424 2525 11458 2556
rect 11424 2522 11458 2525
rect 11424 2457 11458 2483
rect 11424 2449 11458 2457
rect 11424 2389 11458 2410
rect 11424 2376 11458 2389
rect 11424 2321 11458 2337
rect 11424 2303 11458 2321
rect 11424 2253 11458 2264
rect 11424 2230 11458 2253
rect 11424 2185 11458 2191
rect 11424 2157 11458 2185
rect 11424 2117 11458 2118
rect 11424 2084 11458 2117
rect 11424 2015 11458 2045
rect 11424 2011 11458 2015
rect 11424 1947 11458 1972
rect 11424 1938 11458 1947
rect 11424 1879 11458 1899
rect 11424 1865 11458 1879
rect 11424 1811 11458 1826
rect 11424 1792 11458 1811
rect 11424 1743 11458 1753
rect 11424 1719 11458 1743
rect 11424 1675 11458 1680
rect 11424 1646 11458 1675
rect 11424 1573 11458 1607
rect 11424 1505 11458 1534
rect 11424 1500 11458 1505
rect 11424 1437 11458 1461
rect 11424 1427 11458 1437
rect 11424 1369 11458 1388
rect 11424 1354 11458 1369
rect 11424 1301 11458 1315
rect 11424 1281 11458 1301
rect 11424 1233 11458 1242
rect 11424 1208 11458 1233
rect 11424 1165 11458 1169
rect 11424 1135 11458 1165
rect 11424 1063 11458 1096
rect 11424 1062 11458 1063
rect 11424 995 11458 1023
rect 11424 989 11458 995
rect 11424 927 11458 950
rect 11424 916 11458 927
rect 11424 859 11458 877
rect 11424 843 11458 859
rect 11424 791 11458 804
rect 11424 770 11458 791
rect 11424 723 11458 731
rect 11424 697 11458 723
rect 11424 655 11458 658
rect 11424 624 11458 655
rect 11424 553 11458 585
rect 11424 551 11458 553
rect 11424 485 11458 512
rect 11424 478 11458 485
rect 11424 417 11458 439
rect 11424 405 11458 417
rect 13212 38460 13246 38465
rect 13212 38431 13246 38460
rect 13392 38483 13426 38517
rect 14940 38587 14974 38612
rect 14940 38578 14974 38587
rect 14940 38519 14974 38540
rect 14940 38506 14974 38519
rect 13212 38358 13246 38392
rect 13212 38290 13246 38319
rect 13212 38285 13246 38290
rect 13212 38222 13246 38246
rect 13212 38212 13246 38222
rect 13212 38154 13246 38173
rect 13212 38139 13246 38154
rect 13212 38086 13246 38100
rect 13212 38066 13246 38086
rect 13212 38018 13246 38027
rect 13212 37993 13246 38018
rect 13212 37950 13246 37954
rect 13212 37920 13246 37950
rect 13212 37848 13246 37881
rect 13212 37847 13246 37848
rect 13212 37780 13246 37808
rect 13212 37774 13246 37780
rect 13212 37712 13246 37735
rect 13212 37701 13246 37712
rect 13212 37644 13246 37662
rect 13212 37628 13246 37644
rect 13212 37576 13246 37589
rect 13212 37555 13246 37576
rect 13212 37508 13246 37516
rect 13212 37482 13246 37508
rect 13212 37440 13246 37443
rect 13212 37409 13246 37440
rect 13212 37338 13246 37370
rect 13212 37336 13246 37338
rect 13212 37270 13246 37298
rect 13212 37264 13246 37270
rect 13212 37202 13246 37226
rect 13212 37192 13246 37202
rect 13212 37134 13246 37154
rect 13212 37120 13246 37134
rect 13212 37066 13246 37082
rect 13212 37048 13246 37066
rect 13212 36998 13246 37010
rect 13212 36976 13246 36998
rect 13212 36930 13246 36938
rect 13212 36904 13246 36930
rect 13212 36862 13246 36866
rect 13212 36832 13246 36862
rect 13212 36760 13246 36794
rect 13212 36692 13246 36722
rect 13212 36688 13246 36692
rect 13212 36624 13246 36650
rect 13212 36616 13246 36624
rect 13212 36556 13246 36578
rect 13212 36544 13246 36556
rect 13212 36488 13246 36506
rect 13212 36472 13246 36488
rect 13212 36420 13246 36434
rect 13212 36400 13246 36420
rect 13212 36352 13246 36362
rect 13212 36328 13246 36352
rect 13212 36284 13246 36290
rect 13212 36256 13246 36284
rect 13212 36216 13246 36218
rect 13212 36184 13246 36216
rect 13212 36114 13246 36146
rect 13212 36112 13246 36114
rect 13212 36046 13246 36074
rect 13212 36040 13246 36046
rect 13212 35978 13246 36002
rect 13212 35968 13246 35978
rect 13212 35910 13246 35930
rect 13212 35896 13246 35910
rect 13212 35842 13246 35858
rect 13212 35824 13246 35842
rect 13212 35774 13246 35786
rect 13212 35752 13246 35774
rect 13212 35706 13246 35714
rect 13212 35680 13246 35706
rect 13212 35638 13246 35642
rect 13212 35608 13246 35638
rect 13212 35536 13246 35570
rect 13212 35468 13246 35498
rect 13212 35464 13246 35468
rect 13212 35400 13246 35426
rect 13212 35392 13246 35400
rect 13212 35332 13246 35354
rect 13212 35320 13246 35332
rect 13212 35264 13246 35282
rect 13212 35248 13246 35264
rect 13212 35196 13246 35210
rect 13212 35176 13246 35196
rect 13212 35128 13246 35138
rect 13212 35104 13246 35128
rect 13212 35060 13246 35066
rect 13212 35032 13246 35060
rect 13212 34992 13246 34994
rect 13212 34960 13246 34992
rect 13212 34890 13246 34922
rect 13212 34888 13246 34890
rect 13212 34822 13246 34850
rect 13212 34816 13246 34822
rect 13212 34754 13246 34778
rect 13212 34744 13246 34754
rect 13212 34686 13246 34706
rect 13212 34672 13246 34686
rect 13212 34618 13246 34634
rect 13212 34600 13246 34618
rect 13212 34550 13246 34562
rect 13212 34528 13246 34550
rect 13212 34482 13246 34490
rect 13212 34456 13246 34482
rect 13212 34414 13246 34418
rect 13212 34384 13246 34414
rect 13212 34312 13246 34346
rect 13212 34244 13246 34274
rect 13212 34240 13246 34244
rect 13212 34176 13246 34202
rect 13212 34168 13246 34176
rect 13212 34108 13246 34130
rect 13212 34096 13246 34108
rect 13212 34040 13246 34058
rect 13212 34024 13246 34040
rect 13212 33972 13246 33986
rect 13212 33952 13246 33972
rect 13212 33904 13246 33914
rect 13212 33880 13246 33904
rect 13212 33836 13246 33842
rect 13212 33808 13246 33836
rect 13212 33768 13246 33770
rect 13212 33736 13246 33768
rect 13212 33666 13246 33698
rect 13212 33664 13246 33666
rect 13212 33598 13246 33626
rect 13212 33592 13246 33598
rect 13212 33530 13246 33554
rect 13212 33520 13246 33530
rect 13212 33462 13246 33482
rect 13212 33448 13246 33462
rect 13212 33394 13246 33410
rect 13212 33376 13246 33394
rect 13212 33326 13246 33338
rect 13212 33304 13246 33326
rect 13212 33258 13246 33266
rect 13212 33232 13246 33258
rect 13212 33190 13246 33194
rect 13212 33160 13246 33190
rect 13212 33088 13246 33122
rect 13212 33020 13246 33050
rect 13212 33016 13246 33020
rect 13212 32952 13246 32978
rect 13212 32944 13246 32952
rect 13212 32884 13246 32906
rect 13212 32872 13246 32884
rect 13212 32816 13246 32834
rect 13212 32800 13246 32816
rect 13212 32748 13246 32762
rect 13212 32728 13246 32748
rect 13212 32680 13246 32690
rect 13212 32656 13246 32680
rect 13212 32612 13246 32618
rect 13212 32584 13246 32612
rect 13212 32544 13246 32546
rect 13212 32512 13246 32544
rect 13212 32442 13246 32474
rect 13212 32440 13246 32442
rect 13212 32374 13246 32402
rect 13212 32368 13246 32374
rect 13212 32306 13246 32330
rect 13212 32296 13246 32306
rect 13212 32238 13246 32258
rect 13212 32224 13246 32238
rect 13212 32170 13246 32186
rect 13212 32152 13246 32170
rect 13212 32102 13246 32114
rect 13212 32080 13246 32102
rect 13212 32034 13246 32042
rect 13212 32008 13246 32034
rect 13212 31966 13246 31970
rect 13212 31936 13246 31966
rect 13212 31864 13246 31898
rect 13212 31796 13246 31826
rect 13212 31792 13246 31796
rect 13212 31728 13246 31754
rect 13212 31720 13246 31728
rect 13212 31660 13246 31682
rect 13212 31648 13246 31660
rect 13212 31592 13246 31610
rect 13212 31576 13246 31592
rect 13212 31524 13246 31538
rect 13212 31504 13246 31524
rect 13212 31456 13246 31466
rect 13212 31432 13246 31456
rect 13212 31388 13246 31394
rect 13212 31360 13246 31388
rect 13212 31320 13246 31322
rect 13212 31288 13246 31320
rect 13212 31218 13246 31250
rect 13212 31216 13246 31218
rect 13212 31150 13246 31178
rect 13212 31144 13246 31150
rect 13212 31082 13246 31106
rect 13212 31072 13246 31082
rect 13212 31014 13246 31034
rect 13212 31000 13246 31014
rect 13212 30946 13246 30962
rect 13212 30928 13246 30946
rect 13212 30878 13246 30890
rect 13212 30856 13246 30878
rect 13212 30810 13246 30818
rect 13212 30784 13246 30810
rect 13212 30742 13246 30746
rect 13212 30712 13246 30742
rect 13212 30640 13246 30674
rect 13212 30572 13246 30602
rect 13212 30568 13246 30572
rect 13212 30504 13246 30530
rect 13212 30496 13246 30504
rect 13212 30436 13246 30458
rect 13212 30424 13246 30436
rect 13212 30368 13246 30386
rect 13212 30352 13246 30368
rect 13212 30300 13246 30314
rect 13212 30280 13246 30300
rect 13212 30232 13246 30242
rect 13212 30208 13246 30232
rect 13212 30164 13246 30170
rect 13212 30136 13246 30164
rect 13212 30096 13246 30098
rect 13212 30064 13246 30096
rect 13212 29994 13246 30026
rect 13212 29992 13246 29994
rect 13212 29926 13246 29954
rect 13212 29920 13246 29926
rect 13212 29858 13246 29882
rect 13212 29848 13246 29858
rect 13212 29790 13246 29810
rect 13212 29776 13246 29790
rect 13212 29722 13246 29738
rect 13212 29704 13246 29722
rect 13212 29654 13246 29666
rect 13212 29632 13246 29654
rect 13212 29586 13246 29594
rect 13212 29560 13246 29586
rect 13212 29518 13246 29522
rect 13212 29488 13246 29518
rect 13212 29416 13246 29450
rect 13212 29348 13246 29378
rect 13212 29344 13246 29348
rect 13212 29280 13246 29306
rect 13212 29272 13246 29280
rect 13212 29212 13246 29234
rect 13212 29200 13246 29212
rect 13212 29144 13246 29162
rect 13212 29128 13246 29144
rect 13212 29076 13246 29090
rect 13212 29056 13246 29076
rect 13212 29008 13246 29018
rect 13212 28984 13246 29008
rect 13212 28940 13246 28946
rect 13212 28912 13246 28940
rect 13212 28872 13246 28874
rect 13212 28840 13246 28872
rect 13212 28770 13246 28802
rect 13212 28768 13246 28770
rect 13212 28702 13246 28730
rect 13212 28696 13246 28702
rect 13212 28634 13246 28658
rect 13212 28624 13246 28634
rect 13212 28566 13246 28586
rect 13212 28552 13246 28566
rect 13212 28498 13246 28514
rect 13212 28480 13246 28498
rect 13212 28430 13246 28442
rect 13212 28408 13246 28430
rect 13212 28362 13246 28370
rect 13212 28336 13246 28362
rect 13212 28294 13246 28298
rect 13212 28264 13246 28294
rect 13212 28192 13246 28226
rect 13212 28124 13246 28154
rect 13212 28120 13246 28124
rect 13212 28056 13246 28082
rect 13212 28048 13246 28056
rect 13212 27988 13246 28010
rect 13212 27976 13246 27988
rect 13212 27920 13246 27938
rect 13212 27904 13246 27920
rect 13212 27852 13246 27866
rect 13212 27832 13246 27852
rect 13212 27784 13246 27794
rect 13212 27760 13246 27784
rect 13212 27716 13246 27722
rect 13212 27688 13246 27716
rect 13212 27648 13246 27650
rect 13212 27616 13246 27648
rect 13212 27546 13246 27578
rect 13212 27544 13246 27546
rect 13212 27478 13246 27506
rect 13212 27472 13246 27478
rect 13212 27410 13246 27434
rect 13212 27400 13246 27410
rect 13212 27342 13246 27362
rect 13212 27328 13246 27342
rect 13212 27274 13246 27290
rect 13212 27256 13246 27274
rect 13212 27206 13246 27218
rect 13212 27184 13246 27206
rect 13212 27138 13246 27146
rect 13212 27112 13246 27138
rect 13212 27070 13246 27074
rect 13212 27040 13246 27070
rect 13212 26968 13246 27002
rect 13212 26900 13246 26930
rect 13212 26896 13246 26900
rect 13212 26832 13246 26858
rect 13212 26824 13246 26832
rect 13212 26764 13246 26786
rect 13212 26752 13246 26764
rect 13212 26696 13246 26714
rect 13212 26680 13246 26696
rect 13212 26628 13246 26642
rect 13212 26608 13246 26628
rect 13212 26560 13246 26570
rect 13212 26536 13246 26560
rect 13212 26492 13246 26498
rect 13212 26464 13246 26492
rect 13212 26424 13246 26426
rect 13212 26392 13246 26424
rect 13212 26322 13246 26354
rect 13212 26320 13246 26322
rect 13212 26254 13246 26282
rect 13212 26248 13246 26254
rect 13212 26186 13246 26210
rect 13212 26176 13246 26186
rect 13212 26118 13246 26138
rect 13212 26104 13246 26118
rect 13212 26050 13246 26066
rect 13212 26032 13246 26050
rect 13212 25982 13246 25994
rect 13212 25960 13246 25982
rect 13212 25914 13246 25922
rect 13212 25888 13246 25914
rect 13212 25846 13246 25850
rect 13212 25816 13246 25846
rect 13212 25744 13246 25778
rect 13212 25676 13246 25706
rect 13212 25672 13246 25676
rect 13212 25608 13246 25634
rect 13212 25600 13246 25608
rect 13212 25540 13246 25562
rect 13212 25528 13246 25540
rect 13212 25472 13246 25490
rect 13212 25456 13246 25472
rect 13212 25404 13246 25418
rect 13212 25384 13246 25404
rect 13212 25336 13246 25346
rect 13212 25312 13246 25336
rect 13212 25268 13246 25274
rect 13212 25240 13246 25268
rect 13212 25200 13246 25202
rect 13212 25168 13246 25200
rect 13212 25098 13246 25130
rect 13212 25096 13246 25098
rect 13212 25030 13246 25058
rect 13212 25024 13246 25030
rect 13212 24962 13246 24986
rect 13212 24952 13246 24962
rect 13212 24894 13246 24914
rect 13212 24880 13246 24894
rect 13212 24826 13246 24842
rect 13212 24808 13246 24826
rect 13212 24758 13246 24770
rect 13212 24736 13246 24758
rect 13212 24690 13246 24698
rect 13212 24664 13246 24690
rect 13212 24622 13246 24626
rect 13212 24592 13246 24622
rect 13212 24520 13246 24554
rect 13212 24452 13246 24482
rect 13212 24448 13246 24452
rect 13212 24384 13246 24410
rect 13212 24376 13246 24384
rect 13212 24316 13246 24338
rect 13212 24304 13246 24316
rect 13212 24248 13246 24266
rect 13212 24232 13246 24248
rect 13212 24180 13246 24194
rect 13212 24160 13246 24180
rect 13212 24112 13246 24122
rect 13212 24088 13246 24112
rect 13212 24044 13246 24050
rect 13212 24016 13246 24044
rect 13212 23976 13246 23978
rect 13212 23944 13246 23976
rect 13212 23874 13246 23906
rect 13212 23872 13246 23874
rect 13212 23806 13246 23834
rect 13212 23800 13246 23806
rect 13212 23738 13246 23762
rect 13212 23728 13246 23738
rect 13212 23670 13246 23690
rect 13212 23656 13246 23670
rect 13212 23602 13246 23618
rect 13212 23584 13246 23602
rect 13212 23534 13246 23546
rect 13212 23512 13246 23534
rect 13212 23466 13246 23474
rect 13212 23440 13246 23466
rect 13212 23398 13246 23402
rect 13212 23368 13246 23398
rect 13212 23296 13246 23330
rect 13212 23228 13246 23258
rect 13212 23224 13246 23228
rect 13212 23160 13246 23186
rect 13212 23152 13246 23160
rect 13212 23092 13246 23114
rect 13212 23080 13246 23092
rect 13212 23024 13246 23042
rect 13212 23008 13246 23024
rect 13212 22956 13246 22970
rect 13212 22936 13246 22956
rect 13212 22888 13246 22898
rect 13212 22864 13246 22888
rect 13212 22820 13246 22826
rect 13212 22792 13246 22820
rect 13212 22752 13246 22754
rect 13212 22720 13246 22752
rect 13212 22650 13246 22682
rect 13212 22648 13246 22650
rect 13212 22582 13246 22610
rect 13212 22576 13246 22582
rect 13212 22514 13246 22538
rect 13212 22504 13246 22514
rect 13212 22446 13246 22466
rect 13212 22432 13246 22446
rect 13212 22378 13246 22394
rect 13212 22360 13246 22378
rect 13212 22310 13246 22322
rect 13212 22288 13246 22310
rect 13212 22242 13246 22250
rect 13212 22216 13246 22242
rect 13212 22174 13246 22178
rect 13212 22144 13246 22174
rect 13212 22072 13246 22106
rect 13212 22004 13246 22034
rect 13212 22000 13246 22004
rect 13212 21936 13246 21962
rect 13212 21928 13246 21936
rect 13212 21868 13246 21890
rect 13212 21856 13246 21868
rect 13212 21800 13246 21818
rect 13212 21784 13246 21800
rect 13212 21732 13246 21746
rect 13212 21712 13246 21732
rect 13212 21664 13246 21674
rect 13212 21640 13246 21664
rect 13212 21596 13246 21602
rect 13212 21568 13246 21596
rect 13212 21528 13246 21530
rect 13212 21496 13246 21528
rect 13212 21426 13246 21458
rect 13212 21424 13246 21426
rect 13212 21358 13246 21386
rect 13212 21352 13246 21358
rect 13212 21290 13246 21314
rect 13212 21280 13246 21290
rect 13212 21222 13246 21242
rect 13212 21208 13246 21222
rect 13212 21154 13246 21170
rect 13212 21136 13246 21154
rect 13212 21086 13246 21098
rect 13212 21064 13246 21086
rect 13212 21018 13246 21026
rect 13212 20992 13246 21018
rect 13212 20950 13246 20954
rect 13212 20920 13246 20950
rect 13212 20848 13246 20882
rect 13212 20780 13246 20810
rect 13212 20776 13246 20780
rect 13212 20712 13246 20738
rect 13212 20704 13246 20712
rect 13212 20644 13246 20666
rect 13212 20632 13246 20644
rect 13212 20576 13246 20594
rect 13212 20560 13246 20576
rect 13212 20508 13246 20522
rect 13212 20488 13246 20508
rect 13212 20440 13246 20450
rect 13212 20416 13246 20440
rect 13212 20372 13246 20378
rect 13212 20344 13246 20372
rect 13212 20304 13246 20306
rect 13212 20272 13246 20304
rect 13212 20202 13246 20234
rect 13212 20200 13246 20202
rect 13212 20134 13246 20162
rect 13212 20128 13246 20134
rect 13212 20066 13246 20090
rect 13212 20056 13246 20066
rect 13212 19998 13246 20018
rect 13212 19984 13246 19998
rect 13212 19930 13246 19946
rect 13212 19912 13246 19930
rect 13212 19862 13246 19874
rect 13212 19840 13246 19862
rect 13212 19794 13246 19802
rect 13212 19768 13246 19794
rect 13212 19726 13246 19730
rect 13212 19696 13246 19726
rect 13212 19624 13246 19658
rect 13212 19556 13246 19586
rect 13212 19552 13246 19556
rect 13212 19488 13246 19514
rect 13212 19480 13246 19488
rect 13212 19420 13246 19442
rect 13212 19408 13246 19420
rect 13212 19352 13246 19370
rect 13212 19336 13246 19352
rect 13212 19284 13246 19298
rect 13212 19264 13246 19284
rect 13212 19216 13246 19226
rect 13212 19192 13246 19216
rect 13212 19148 13246 19154
rect 13212 19120 13246 19148
rect 13212 19080 13246 19082
rect 13212 19048 13246 19080
rect 13212 18978 13246 19010
rect 13212 18976 13246 18978
rect 13212 18910 13246 18938
rect 13212 18904 13246 18910
rect 13212 18842 13246 18866
rect 13212 18832 13246 18842
rect 13212 18774 13246 18794
rect 13212 18760 13246 18774
rect 13212 18706 13246 18722
rect 13212 18688 13246 18706
rect 13212 18638 13246 18650
rect 13212 18616 13246 18638
rect 13212 18570 13246 18578
rect 13212 18544 13246 18570
rect 13212 18502 13246 18506
rect 13212 18472 13246 18502
rect 13212 18400 13246 18434
rect 13212 18332 13246 18362
rect 13212 18328 13246 18332
rect 13212 18264 13246 18290
rect 13212 18256 13246 18264
rect 13212 18196 13246 18218
rect 13212 18184 13246 18196
rect 13212 18128 13246 18146
rect 13212 18112 13246 18128
rect 13212 18060 13246 18074
rect 13212 18040 13246 18060
rect 13212 17992 13246 18002
rect 13212 17968 13246 17992
rect 13212 17924 13246 17930
rect 13212 17896 13246 17924
rect 13212 17856 13246 17858
rect 13212 17824 13246 17856
rect 13212 17754 13246 17786
rect 13212 17752 13246 17754
rect 13212 17686 13246 17714
rect 13212 17680 13246 17686
rect 13212 17618 13246 17642
rect 13212 17608 13246 17618
rect 13212 17550 13246 17570
rect 13212 17536 13246 17550
rect 13212 17482 13246 17498
rect 13212 17464 13246 17482
rect 13212 17414 13246 17426
rect 13212 17392 13246 17414
rect 13212 17346 13246 17354
rect 13212 17320 13246 17346
rect 13212 17278 13246 17282
rect 13212 17248 13246 17278
rect 13212 17176 13246 17210
rect 13212 17108 13246 17138
rect 13212 17104 13246 17108
rect 13212 17040 13246 17066
rect 13212 17032 13246 17040
rect 13212 16972 13246 16994
rect 13212 16960 13246 16972
rect 13212 16904 13246 16922
rect 13212 16888 13246 16904
rect 13212 16836 13246 16850
rect 13212 16816 13246 16836
rect 13212 16768 13246 16778
rect 13212 16744 13246 16768
rect 13212 16700 13246 16706
rect 13212 16672 13246 16700
rect 13212 16632 13246 16634
rect 13212 16600 13246 16632
rect 13212 16530 13246 16562
rect 13212 16528 13246 16530
rect 13212 16462 13246 16490
rect 13212 16456 13246 16462
rect 13212 16394 13246 16418
rect 13212 16384 13246 16394
rect 13212 16326 13246 16346
rect 13212 16312 13246 16326
rect 13212 16258 13246 16274
rect 13212 16240 13246 16258
rect 13212 16190 13246 16202
rect 13212 16168 13246 16190
rect 13212 16122 13246 16130
rect 13212 16096 13246 16122
rect 13212 16054 13246 16058
rect 13212 16024 13246 16054
rect 13212 15952 13246 15986
rect 13212 15884 13246 15914
rect 13212 15880 13246 15884
rect 13212 15816 13246 15842
rect 13212 15808 13246 15816
rect 13212 15748 13246 15770
rect 13212 15736 13246 15748
rect 13212 15680 13246 15698
rect 13212 15664 13246 15680
rect 13212 15612 13246 15626
rect 13212 15592 13246 15612
rect 13212 15544 13246 15554
rect 13212 15520 13246 15544
rect 13212 15476 13246 15482
rect 13212 15448 13246 15476
rect 13212 15408 13246 15410
rect 13212 15376 13246 15408
rect 13212 15306 13246 15338
rect 13212 15304 13246 15306
rect 13212 15238 13246 15266
rect 13212 15232 13246 15238
rect 13212 15170 13246 15194
rect 13212 15160 13246 15170
rect 13212 15102 13246 15122
rect 13212 15088 13246 15102
rect 13212 15034 13246 15050
rect 13212 15016 13246 15034
rect 13212 14966 13246 14978
rect 13212 14944 13246 14966
rect 13212 14898 13246 14906
rect 13212 14872 13246 14898
rect 13212 14830 13246 14834
rect 13212 14800 13246 14830
rect 13212 14728 13246 14762
rect 13212 14660 13246 14690
rect 13212 14656 13246 14660
rect 13212 14592 13246 14618
rect 13212 14584 13246 14592
rect 13212 14524 13246 14546
rect 13212 14512 13246 14524
rect 13212 14456 13246 14474
rect 13212 14440 13246 14456
rect 13212 14388 13246 14402
rect 13212 14368 13246 14388
rect 13212 14320 13246 14330
rect 13212 14296 13246 14320
rect 13212 14252 13246 14258
rect 13212 14224 13246 14252
rect 13212 14184 13246 14186
rect 13212 14152 13246 14184
rect 13212 14082 13246 14114
rect 13212 14080 13246 14082
rect 13212 14014 13246 14042
rect 13212 14008 13246 14014
rect 13212 13946 13246 13970
rect 13212 13936 13246 13946
rect 13212 13878 13246 13898
rect 13212 13864 13246 13878
rect 13212 13810 13246 13826
rect 13212 13792 13246 13810
rect 13212 13742 13246 13754
rect 13212 13720 13246 13742
rect 13212 13674 13246 13682
rect 13212 13648 13246 13674
rect 13212 13606 13246 13610
rect 13212 13576 13246 13606
rect 13212 13504 13246 13538
rect 13212 13436 13246 13466
rect 13212 13432 13246 13436
rect 13212 13368 13246 13394
rect 13212 13360 13246 13368
rect 13212 13300 13246 13322
rect 13212 13288 13246 13300
rect 13212 13232 13246 13250
rect 13212 13216 13246 13232
rect 13212 13164 13246 13178
rect 13212 13144 13246 13164
rect 13212 13096 13246 13106
rect 13212 13072 13246 13096
rect 13212 13028 13246 13034
rect 13212 13000 13246 13028
rect 13212 12960 13246 12962
rect 13212 12928 13246 12960
rect 13212 12858 13246 12890
rect 13212 12856 13246 12858
rect 13212 12790 13246 12818
rect 13212 12784 13246 12790
rect 13212 12722 13246 12746
rect 13212 12712 13246 12722
rect 13212 12654 13246 12674
rect 13212 12640 13246 12654
rect 13212 12586 13246 12602
rect 13212 12568 13246 12586
rect 13212 12518 13246 12530
rect 13212 12496 13246 12518
rect 13212 12450 13246 12458
rect 13212 12424 13246 12450
rect 13212 12382 13246 12386
rect 13212 12352 13246 12382
rect 13212 12280 13246 12314
rect 13212 12212 13246 12242
rect 13212 12208 13246 12212
rect 13212 12144 13246 12170
rect 13212 12136 13246 12144
rect 13212 12076 13246 12098
rect 13212 12064 13246 12076
rect 13212 12008 13246 12026
rect 13212 11992 13246 12008
rect 13212 11940 13246 11954
rect 13212 11920 13246 11940
rect 13212 11872 13246 11882
rect 13212 11848 13246 11872
rect 13212 11804 13246 11810
rect 13212 11776 13246 11804
rect 13212 11736 13246 11738
rect 13212 11704 13246 11736
rect 13212 11634 13246 11666
rect 13212 11632 13246 11634
rect 13212 11566 13246 11594
rect 13212 11560 13246 11566
rect 13212 11498 13246 11522
rect 13212 11488 13246 11498
rect 13212 11430 13246 11450
rect 13212 11416 13246 11430
rect 13212 11362 13246 11378
rect 13212 11344 13246 11362
rect 13212 11294 13246 11306
rect 13212 11272 13246 11294
rect 13212 11226 13246 11234
rect 13212 11200 13246 11226
rect 13212 11158 13246 11162
rect 13212 11128 13246 11158
rect 13212 11056 13246 11090
rect 13212 10988 13246 11018
rect 13212 10984 13246 10988
rect 13212 10920 13246 10946
rect 13212 10912 13246 10920
rect 13212 10852 13246 10874
rect 13212 10840 13246 10852
rect 13212 10784 13246 10802
rect 13212 10768 13246 10784
rect 13212 10716 13246 10730
rect 13212 10696 13246 10716
rect 13212 10648 13246 10658
rect 13212 10624 13246 10648
rect 13212 10580 13246 10586
rect 13212 10552 13246 10580
rect 13212 10512 13246 10514
rect 13212 10480 13246 10512
rect 13212 10410 13246 10442
rect 13212 10408 13246 10410
rect 13212 10342 13246 10370
rect 13212 10336 13246 10342
rect 13212 10274 13246 10298
rect 13212 10264 13246 10274
rect 13212 10206 13246 10226
rect 13212 10192 13246 10206
rect 13212 10138 13246 10154
rect 13212 10120 13246 10138
rect 13212 10070 13246 10082
rect 13212 10048 13246 10070
rect 13212 10002 13246 10010
rect 13212 9976 13246 10002
rect 13212 9934 13246 9938
rect 13212 9904 13246 9934
rect 13212 9832 13246 9866
rect 13212 9764 13246 9794
rect 13212 9760 13246 9764
rect 13212 9696 13246 9722
rect 13212 9688 13246 9696
rect 13212 9628 13246 9650
rect 13212 9616 13246 9628
rect 13212 9560 13246 9578
rect 13212 9544 13246 9560
rect 13212 9492 13246 9506
rect 13212 9472 13246 9492
rect 13212 9424 13246 9434
rect 13212 9400 13246 9424
rect 13212 9356 13246 9362
rect 13212 9328 13246 9356
rect 13212 9288 13246 9290
rect 13212 9256 13246 9288
rect 13212 9186 13246 9218
rect 13212 9184 13246 9186
rect 13212 9118 13246 9146
rect 13212 9112 13246 9118
rect 13212 9050 13246 9074
rect 13212 9040 13246 9050
rect 13212 8982 13246 9002
rect 13212 8968 13246 8982
rect 13212 8914 13246 8930
rect 13212 8896 13246 8914
rect 13212 8846 13246 8858
rect 13212 8824 13246 8846
rect 13212 8778 13246 8786
rect 13212 8752 13246 8778
rect 13212 8710 13246 8714
rect 13212 8680 13246 8710
rect 13212 8608 13246 8642
rect 13212 8540 13246 8570
rect 13212 8536 13246 8540
rect 13212 8472 13246 8498
rect 13212 8464 13246 8472
rect 13212 8404 13246 8426
rect 13212 8392 13246 8404
rect 13212 8336 13246 8354
rect 13212 8320 13246 8336
rect 13212 8268 13246 8282
rect 13212 8248 13246 8268
rect 13212 8200 13246 8210
rect 13212 8176 13246 8200
rect 13212 8132 13246 8138
rect 13212 8104 13246 8132
rect 13212 8064 13246 8066
rect 13212 8032 13246 8064
rect 13212 7962 13246 7994
rect 13212 7960 13246 7962
rect 13212 7894 13246 7922
rect 13212 7888 13246 7894
rect 13212 7826 13246 7850
rect 13212 7816 13246 7826
rect 13212 7758 13246 7778
rect 13212 7744 13246 7758
rect 13212 7690 13246 7706
rect 13212 7672 13246 7690
rect 13212 7622 13246 7634
rect 13212 7600 13246 7622
rect 13212 7554 13246 7562
rect 13212 7528 13246 7554
rect 13212 7486 13246 7490
rect 13212 7456 13246 7486
rect 13212 7384 13246 7418
rect 13212 7316 13246 7346
rect 13212 7312 13246 7316
rect 13212 7248 13246 7274
rect 13212 7240 13246 7248
rect 13212 7180 13246 7202
rect 13212 7168 13246 7180
rect 13212 7112 13246 7130
rect 13212 7096 13246 7112
rect 13212 7044 13246 7058
rect 13212 7024 13246 7044
rect 13212 6976 13246 6986
rect 13212 6952 13246 6976
rect 13212 6908 13246 6914
rect 13212 6880 13246 6908
rect 13212 6840 13246 6842
rect 13212 6808 13246 6840
rect 13212 6738 13246 6770
rect 13212 6736 13246 6738
rect 13212 6670 13246 6698
rect 13212 6664 13246 6670
rect 13212 6602 13246 6626
rect 13212 6592 13246 6602
rect 13212 6534 13246 6554
rect 13212 6520 13246 6534
rect 13212 6466 13246 6482
rect 13212 6448 13246 6466
rect 13212 6398 13246 6410
rect 13212 6376 13246 6398
rect 13212 6330 13246 6338
rect 13212 6304 13246 6330
rect 13212 6262 13246 6266
rect 13212 6232 13246 6262
rect 13212 6160 13246 6194
rect 13212 6092 13246 6122
rect 13212 6088 13246 6092
rect 13212 6024 13246 6050
rect 13212 6016 13246 6024
rect 13212 5956 13246 5978
rect 13212 5944 13246 5956
rect 13212 5888 13246 5906
rect 13212 5872 13246 5888
rect 13212 5820 13246 5834
rect 13212 5800 13246 5820
rect 13212 5752 13246 5762
rect 13212 5728 13246 5752
rect 13212 5684 13246 5690
rect 13212 5656 13246 5684
rect 13212 5616 13246 5618
rect 13212 5584 13246 5616
rect 13212 5514 13246 5546
rect 13212 5512 13246 5514
rect 13212 5446 13246 5474
rect 13212 5440 13246 5446
rect 13212 5378 13246 5402
rect 13212 5368 13246 5378
rect 13212 5310 13246 5330
rect 13212 5296 13246 5310
rect 13212 5242 13246 5258
rect 13212 5224 13246 5242
rect 13212 5174 13246 5186
rect 13212 5152 13246 5174
rect 13212 5106 13246 5114
rect 13212 5080 13246 5106
rect 13212 5038 13246 5042
rect 13212 5008 13246 5038
rect 13212 4936 13246 4970
rect 13212 4868 13246 4898
rect 13212 4864 13246 4868
rect 13212 4800 13246 4826
rect 13212 4792 13246 4800
rect 13212 4732 13246 4754
rect 13212 4720 13246 4732
rect 13212 4664 13246 4682
rect 13212 4648 13246 4664
rect 13212 4596 13246 4610
rect 13212 4576 13246 4596
rect 13212 4528 13246 4538
rect 13212 4504 13246 4528
rect 13212 4460 13246 4466
rect 13212 4432 13246 4460
rect 13212 4392 13246 4394
rect 13212 4360 13246 4392
rect 13212 4290 13246 4322
rect 13212 4288 13246 4290
rect 13212 4222 13246 4250
rect 13212 4216 13246 4222
rect 13212 4154 13246 4178
rect 13212 4144 13246 4154
rect 13212 4086 13246 4106
rect 13212 4072 13246 4086
rect 13212 4018 13246 4034
rect 13212 4000 13246 4018
rect 13212 3950 13246 3962
rect 13212 3928 13246 3950
rect 13212 3882 13246 3890
rect 13212 3856 13246 3882
rect 13212 3814 13246 3818
rect 13212 3784 13246 3814
rect 13212 3712 13246 3746
rect 13212 3644 13246 3674
rect 13212 3640 13246 3644
rect 13212 3576 13246 3602
rect 13212 3568 13246 3576
rect 13212 3508 13246 3530
rect 13212 3496 13246 3508
rect 13212 3440 13246 3458
rect 13212 3424 13246 3440
rect 13212 3372 13246 3386
rect 13212 3352 13246 3372
rect 13212 3304 13246 3314
rect 13212 3280 13246 3304
rect 13212 3236 13246 3242
rect 13212 3208 13246 3236
rect 13212 3168 13246 3170
rect 13212 3136 13246 3168
rect 13212 3066 13246 3098
rect 13212 3064 13246 3066
rect 13212 2998 13246 3026
rect 13212 2992 13246 2998
rect 13212 2930 13246 2954
rect 13212 2920 13246 2930
rect 13212 2862 13246 2882
rect 13212 2848 13246 2862
rect 13212 2794 13246 2810
rect 13212 2776 13246 2794
rect 13212 2726 13246 2738
rect 13212 2704 13246 2726
rect 13212 2658 13246 2666
rect 13212 2632 13246 2658
rect 13212 2590 13246 2594
rect 13212 2560 13246 2590
rect 13212 2488 13246 2522
rect 13212 2420 13246 2450
rect 13212 2416 13246 2420
rect 13212 2352 13246 2378
rect 13212 2344 13246 2352
rect 13212 2284 13246 2306
rect 13212 2272 13246 2284
rect 13212 2216 13246 2234
rect 13212 2200 13246 2216
rect 13212 2148 13246 2162
rect 13212 2128 13246 2148
rect 13212 2080 13246 2090
rect 13212 2056 13246 2080
rect 13212 2012 13246 2018
rect 13212 1984 13246 2012
rect 13212 1944 13246 1946
rect 13212 1912 13246 1944
rect 13212 1842 13246 1874
rect 13212 1840 13246 1842
rect 13212 1774 13246 1802
rect 13212 1768 13246 1774
rect 13212 1706 13246 1730
rect 13212 1696 13246 1706
rect 13212 1638 13246 1658
rect 13212 1624 13246 1638
rect 13212 1570 13246 1586
rect 13212 1552 13246 1570
rect 13212 1502 13246 1514
rect 13212 1480 13246 1502
rect 13212 1434 13246 1442
rect 13212 1408 13246 1434
rect 13212 1366 13246 1370
rect 13212 1336 13246 1366
rect 13212 1264 13246 1298
rect 13212 1196 13246 1226
rect 13212 1192 13246 1196
rect 13212 1128 13246 1154
rect 13212 1120 13246 1128
rect 13212 1060 13246 1082
rect 13212 1048 13246 1060
rect 13212 992 13246 1010
rect 13212 976 13246 992
rect 13212 924 13246 938
rect 13212 904 13246 924
rect 13212 856 13246 866
rect 13212 832 13246 856
rect 13212 788 13246 794
rect 13212 760 13246 788
rect 13212 720 13246 722
rect 13212 688 13246 720
rect 13212 618 13246 650
rect 13212 616 13246 618
rect 13212 550 13246 578
rect 13212 544 13246 550
rect 13212 482 13246 506
rect 13212 472 13246 482
rect 11424 349 11458 366
rect 11424 332 11458 349
rect 11424 281 11458 293
rect 11424 259 11458 281
rect 11610 383 11644 417
rect 11610 325 11644 345
rect 13212 414 13246 434
rect 13212 400 13246 414
rect 14940 38451 14974 38468
rect 14940 38434 14974 38451
rect 14940 38383 14974 38396
rect 14940 38362 14974 38383
rect 14940 38315 14974 38324
rect 14940 38290 14974 38315
rect 14940 38247 14974 38252
rect 14940 38218 14974 38247
rect 14940 38179 14974 38180
rect 14940 38146 14974 38179
rect 14940 38077 14974 38108
rect 14940 38074 14974 38077
rect 14940 38009 14974 38036
rect 14940 38002 14974 38009
rect 14940 37941 14974 37964
rect 14940 37930 14974 37941
rect 14940 37873 14974 37892
rect 14940 37858 14974 37873
rect 14940 37805 14974 37820
rect 14940 37786 14974 37805
rect 14940 37737 14974 37748
rect 14940 37714 14974 37737
rect 14940 37669 14974 37676
rect 14940 37642 14974 37669
rect 14940 37601 14974 37604
rect 14940 37570 14974 37601
rect 14940 37499 14974 37532
rect 14940 37498 14974 37499
rect 14940 37431 14974 37460
rect 14940 37426 14974 37431
rect 14940 37363 14974 37388
rect 14940 37354 14974 37363
rect 14940 37295 14974 37316
rect 14940 37282 14974 37295
rect 14940 37227 14974 37244
rect 14940 37210 14974 37227
rect 14940 37159 14974 37172
rect 14940 37138 14974 37159
rect 14940 37091 14974 37100
rect 14940 37066 14974 37091
rect 14940 37023 14974 37028
rect 14940 36994 14974 37023
rect 14940 36955 14974 36956
rect 14940 36922 14974 36955
rect 14940 36853 14974 36884
rect 14940 36850 14974 36853
rect 14940 36785 14974 36812
rect 14940 36778 14974 36785
rect 14940 36717 14974 36740
rect 14940 36706 14974 36717
rect 14940 36649 14974 36668
rect 14940 36634 14974 36649
rect 14940 36581 14974 36596
rect 14940 36562 14974 36581
rect 14940 36513 14974 36524
rect 14940 36490 14974 36513
rect 14940 36445 14974 36452
rect 14940 36418 14974 36445
rect 14940 36377 14974 36380
rect 14940 36346 14974 36377
rect 14940 36275 14974 36308
rect 14940 36274 14974 36275
rect 14940 36207 14974 36236
rect 14940 36202 14974 36207
rect 14940 36139 14974 36164
rect 14940 36130 14974 36139
rect 14940 36071 14974 36092
rect 14940 36058 14974 36071
rect 14940 36003 14974 36020
rect 14940 35986 14974 36003
rect 14940 35935 14974 35948
rect 14940 35914 14974 35935
rect 14940 35867 14974 35876
rect 14940 35842 14974 35867
rect 14940 35799 14974 35804
rect 14940 35770 14974 35799
rect 14940 35731 14974 35732
rect 14940 35698 14974 35731
rect 14940 35629 14974 35660
rect 14940 35626 14974 35629
rect 14940 35561 14974 35588
rect 14940 35554 14974 35561
rect 14940 35493 14974 35516
rect 14940 35482 14974 35493
rect 14940 35425 14974 35444
rect 14940 35410 14974 35425
rect 14940 35357 14974 35372
rect 14940 35338 14974 35357
rect 14940 35289 14974 35300
rect 14940 35266 14974 35289
rect 14940 35221 14974 35228
rect 14940 35194 14974 35221
rect 14940 35153 14974 35156
rect 14940 35122 14974 35153
rect 14940 35051 14974 35084
rect 14940 35050 14974 35051
rect 14940 34983 14974 35012
rect 14940 34978 14974 34983
rect 14940 34915 14974 34940
rect 14940 34906 14974 34915
rect 14940 34847 14974 34868
rect 14940 34834 14974 34847
rect 14940 34779 14974 34796
rect 14940 34762 14974 34779
rect 14940 34711 14974 34724
rect 14940 34690 14974 34711
rect 14940 34643 14974 34652
rect 14940 34618 14974 34643
rect 14940 34575 14974 34580
rect 14940 34546 14974 34575
rect 14940 34507 14974 34508
rect 14940 34474 14974 34507
rect 14940 34405 14974 34436
rect 14940 34402 14974 34405
rect 14940 34337 14974 34364
rect 14940 34330 14974 34337
rect 14940 34269 14974 34292
rect 14940 34258 14974 34269
rect 14940 34201 14974 34220
rect 14940 34186 14974 34201
rect 14940 34133 14974 34148
rect 14940 34114 14974 34133
rect 14940 34065 14974 34076
rect 14940 34042 14974 34065
rect 14940 33997 14974 34004
rect 14940 33970 14974 33997
rect 14940 33929 14974 33932
rect 14940 33898 14974 33929
rect 14940 33827 14974 33860
rect 14940 33826 14974 33827
rect 14940 33759 14974 33788
rect 14940 33754 14974 33759
rect 14940 33691 14974 33716
rect 14940 33682 14974 33691
rect 14940 33623 14974 33644
rect 14940 33610 14974 33623
rect 14940 33555 14974 33572
rect 14940 33538 14974 33555
rect 14940 33487 14974 33500
rect 14940 33466 14974 33487
rect 14940 33419 14974 33428
rect 14940 33394 14974 33419
rect 14940 33351 14974 33356
rect 14940 33322 14974 33351
rect 14940 33283 14974 33284
rect 14940 33250 14974 33283
rect 14940 33181 14974 33212
rect 14940 33178 14974 33181
rect 14940 33113 14974 33140
rect 14940 33106 14974 33113
rect 14940 33045 14974 33068
rect 14940 33034 14974 33045
rect 14940 32977 14974 32996
rect 14940 32962 14974 32977
rect 14940 32909 14974 32924
rect 14940 32890 14974 32909
rect 14940 32841 14974 32852
rect 14940 32818 14974 32841
rect 14940 32773 14974 32780
rect 14940 32746 14974 32773
rect 14940 32705 14974 32708
rect 14940 32674 14974 32705
rect 14940 32603 14974 32636
rect 14940 32602 14974 32603
rect 14940 32535 14974 32564
rect 14940 32530 14974 32535
rect 14940 32467 14974 32492
rect 14940 32458 14974 32467
rect 14940 32399 14974 32420
rect 14940 32386 14974 32399
rect 14940 32331 14974 32348
rect 14940 32314 14974 32331
rect 14940 32263 14974 32276
rect 14940 32242 14974 32263
rect 14940 32195 14974 32204
rect 14940 32170 14974 32195
rect 14940 32127 14974 32132
rect 14940 32098 14974 32127
rect 14940 32059 14974 32060
rect 14940 32026 14974 32059
rect 14940 31957 14974 31988
rect 14940 31954 14974 31957
rect 14940 31889 14974 31916
rect 14940 31882 14974 31889
rect 14940 31821 14974 31844
rect 14940 31810 14974 31821
rect 14940 31753 14974 31772
rect 14940 31738 14974 31753
rect 14940 31685 14974 31700
rect 14940 31666 14974 31685
rect 14940 31617 14974 31628
rect 14940 31594 14974 31617
rect 14940 31549 14974 31556
rect 14940 31522 14974 31549
rect 14940 31481 14974 31484
rect 14940 31450 14974 31481
rect 14940 31379 14974 31412
rect 14940 31378 14974 31379
rect 14940 31311 14974 31340
rect 14940 31306 14974 31311
rect 14940 31243 14974 31268
rect 14940 31234 14974 31243
rect 14940 31175 14974 31196
rect 14940 31162 14974 31175
rect 14940 31107 14974 31124
rect 14940 31090 14974 31107
rect 14940 31039 14974 31052
rect 14940 31018 14974 31039
rect 14940 30971 14974 30980
rect 14940 30946 14974 30971
rect 14940 30903 14974 30908
rect 14940 30874 14974 30903
rect 14940 30835 14974 30836
rect 14940 30802 14974 30835
rect 14940 30733 14974 30764
rect 14940 30730 14974 30733
rect 14940 30665 14974 30692
rect 14940 30658 14974 30665
rect 14940 30597 14974 30620
rect 14940 30586 14974 30597
rect 14940 30529 14974 30548
rect 14940 30514 14974 30529
rect 14940 30461 14974 30476
rect 14940 30442 14974 30461
rect 14940 30393 14974 30404
rect 14940 30370 14974 30393
rect 14940 30325 14974 30332
rect 14940 30298 14974 30325
rect 14940 30257 14974 30260
rect 14940 30226 14974 30257
rect 14940 30155 14974 30188
rect 14940 30154 14974 30155
rect 14940 30087 14974 30116
rect 14940 30082 14974 30087
rect 14940 30019 14974 30044
rect 14940 30010 14974 30019
rect 14940 29951 14974 29972
rect 14940 29938 14974 29951
rect 14940 29883 14974 29900
rect 14940 29866 14974 29883
rect 14940 29815 14974 29828
rect 14940 29794 14974 29815
rect 14940 29747 14974 29756
rect 14940 29722 14974 29747
rect 14940 29679 14974 29684
rect 14940 29650 14974 29679
rect 14940 29611 14974 29612
rect 14940 29578 14974 29611
rect 14940 29509 14974 29540
rect 14940 29506 14974 29509
rect 14940 29441 14974 29468
rect 14940 29434 14974 29441
rect 14940 29373 14974 29396
rect 14940 29362 14974 29373
rect 14940 29305 14974 29324
rect 14940 29290 14974 29305
rect 14940 29237 14974 29252
rect 14940 29218 14974 29237
rect 14940 29169 14974 29180
rect 14940 29146 14974 29169
rect 14940 29101 14974 29108
rect 14940 29074 14974 29101
rect 14940 29033 14974 29036
rect 14940 29002 14974 29033
rect 14940 28931 14974 28964
rect 14940 28930 14974 28931
rect 14940 28863 14974 28892
rect 14940 28858 14974 28863
rect 14940 28795 14974 28820
rect 14940 28786 14974 28795
rect 14940 28727 14974 28748
rect 14940 28714 14974 28727
rect 14940 28659 14974 28676
rect 14940 28642 14974 28659
rect 14940 28591 14974 28604
rect 14940 28570 14974 28591
rect 14940 28523 14974 28532
rect 14940 28498 14974 28523
rect 14940 28455 14974 28460
rect 14940 28426 14974 28455
rect 14940 28387 14974 28388
rect 14940 28354 14974 28387
rect 14940 28285 14974 28316
rect 14940 28282 14974 28285
rect 14940 28217 14974 28244
rect 14940 28210 14974 28217
rect 14940 28149 14974 28172
rect 14940 28138 14974 28149
rect 14940 28081 14974 28100
rect 14940 28066 14974 28081
rect 14940 28013 14974 28028
rect 14940 27994 14974 28013
rect 14940 27945 14974 27956
rect 14940 27922 14974 27945
rect 14940 27877 14974 27884
rect 14940 27850 14974 27877
rect 14940 27809 14974 27812
rect 14940 27778 14974 27809
rect 14940 27707 14974 27740
rect 14940 27706 14974 27707
rect 14940 27639 14974 27668
rect 14940 27634 14974 27639
rect 14940 27571 14974 27596
rect 14940 27562 14974 27571
rect 14940 27503 14974 27524
rect 14940 27490 14974 27503
rect 14940 27435 14974 27452
rect 14940 27418 14974 27435
rect 14940 27367 14974 27380
rect 14940 27346 14974 27367
rect 14940 27299 14974 27308
rect 14940 27274 14974 27299
rect 14940 27231 14974 27236
rect 14940 27202 14974 27231
rect 14940 27163 14974 27164
rect 14940 27130 14974 27163
rect 14940 27061 14974 27092
rect 14940 27058 14974 27061
rect 14940 26993 14974 27020
rect 14940 26986 14974 26993
rect 14940 26925 14974 26948
rect 14940 26914 14974 26925
rect 14940 26857 14974 26876
rect 14940 26842 14974 26857
rect 14940 26789 14974 26804
rect 14940 26770 14974 26789
rect 14940 26721 14974 26732
rect 14940 26698 14974 26721
rect 14940 26653 14974 26660
rect 14940 26626 14974 26653
rect 14940 26585 14974 26588
rect 14940 26554 14974 26585
rect 14940 26483 14974 26516
rect 14940 26482 14974 26483
rect 14940 26415 14974 26444
rect 14940 26410 14974 26415
rect 14940 26347 14974 26372
rect 14940 26338 14974 26347
rect 14940 26279 14974 26300
rect 14940 26266 14974 26279
rect 14940 26211 14974 26228
rect 14940 26194 14974 26211
rect 14940 26143 14974 26156
rect 14940 26122 14974 26143
rect 14940 26075 14974 26084
rect 14940 26050 14974 26075
rect 14940 26007 14974 26012
rect 14940 25978 14974 26007
rect 14940 25939 14974 25940
rect 14940 25906 14974 25939
rect 14940 25837 14974 25868
rect 14940 25834 14974 25837
rect 14940 25769 14974 25796
rect 14940 25762 14974 25769
rect 14940 25701 14974 25724
rect 14940 25690 14974 25701
rect 14940 25633 14974 25652
rect 14940 25618 14974 25633
rect 14940 25565 14974 25580
rect 14940 25546 14974 25565
rect 14940 25497 14974 25508
rect 14940 25474 14974 25497
rect 14940 25429 14974 25436
rect 14940 25402 14974 25429
rect 14940 25361 14974 25364
rect 14940 25330 14974 25361
rect 14940 25259 14974 25292
rect 14940 25258 14974 25259
rect 14940 25191 14974 25220
rect 14940 25186 14974 25191
rect 14940 25123 14974 25148
rect 14940 25114 14974 25123
rect 14940 25055 14974 25076
rect 14940 25042 14974 25055
rect 14940 24987 14974 25004
rect 14940 24970 14974 24987
rect 14940 24919 14974 24932
rect 14940 24898 14974 24919
rect 14940 24851 14974 24860
rect 14940 24826 14974 24851
rect 14940 24783 14974 24788
rect 14940 24754 14974 24783
rect 14940 24715 14974 24716
rect 14940 24682 14974 24715
rect 14940 24613 14974 24644
rect 14940 24610 14974 24613
rect 14940 24545 14974 24572
rect 14940 24538 14974 24545
rect 14940 24477 14974 24500
rect 14940 24466 14974 24477
rect 14940 24409 14974 24428
rect 14940 24394 14974 24409
rect 14940 24341 14974 24356
rect 14940 24322 14974 24341
rect 14940 24273 14974 24284
rect 14940 24250 14974 24273
rect 14940 24205 14974 24212
rect 14940 24178 14974 24205
rect 14940 24137 14974 24140
rect 14940 24106 14974 24137
rect 14940 24035 14974 24068
rect 14940 24034 14974 24035
rect 14940 23967 14974 23996
rect 14940 23962 14974 23967
rect 14940 23899 14974 23924
rect 14940 23890 14974 23899
rect 14940 23831 14974 23852
rect 14940 23818 14974 23831
rect 14940 23763 14974 23780
rect 14940 23746 14974 23763
rect 14940 23695 14974 23708
rect 14940 23674 14974 23695
rect 14940 23627 14974 23636
rect 14940 23602 14974 23627
rect 14940 23559 14974 23564
rect 14940 23530 14974 23559
rect 14940 23491 14974 23492
rect 14940 23458 14974 23491
rect 14940 23389 14974 23420
rect 14940 23386 14974 23389
rect 14940 23321 14974 23348
rect 14940 23314 14974 23321
rect 14940 23253 14974 23276
rect 14940 23242 14974 23253
rect 14940 23185 14974 23204
rect 14940 23170 14974 23185
rect 14940 23117 14974 23132
rect 14940 23098 14974 23117
rect 14940 23049 14974 23060
rect 14940 23026 14974 23049
rect 14940 22981 14974 22988
rect 14940 22954 14974 22981
rect 14940 22913 14974 22916
rect 14940 22882 14974 22913
rect 14940 22811 14974 22844
rect 14940 22810 14974 22811
rect 14940 22743 14974 22772
rect 14940 22738 14974 22743
rect 14940 22675 14974 22700
rect 14940 22666 14974 22675
rect 14940 22607 14974 22628
rect 14940 22594 14974 22607
rect 14940 22539 14974 22556
rect 14940 22522 14974 22539
rect 14940 22471 14974 22484
rect 14940 22450 14974 22471
rect 14940 22403 14974 22412
rect 14940 22378 14974 22403
rect 14940 22335 14974 22340
rect 14940 22306 14974 22335
rect 14940 22267 14974 22268
rect 14940 22234 14974 22267
rect 14940 22165 14974 22196
rect 14940 22162 14974 22165
rect 14940 22097 14974 22124
rect 14940 22090 14974 22097
rect 14940 22029 14974 22052
rect 14940 22018 14974 22029
rect 14940 21961 14974 21980
rect 14940 21946 14974 21961
rect 14940 21893 14974 21908
rect 14940 21874 14974 21893
rect 14940 21825 14974 21836
rect 14940 21802 14974 21825
rect 14940 21757 14974 21764
rect 14940 21730 14974 21757
rect 14940 21689 14974 21692
rect 14940 21658 14974 21689
rect 14940 21587 14974 21620
rect 14940 21586 14974 21587
rect 14940 21519 14974 21548
rect 14940 21514 14974 21519
rect 14940 21451 14974 21476
rect 14940 21442 14974 21451
rect 14940 21383 14974 21404
rect 14940 21370 14974 21383
rect 14940 21315 14974 21332
rect 14940 21298 14974 21315
rect 14940 21247 14974 21260
rect 14940 21226 14974 21247
rect 14940 21179 14974 21188
rect 14940 21154 14974 21179
rect 14940 21111 14974 21116
rect 14940 21082 14974 21111
rect 14940 21043 14974 21044
rect 14940 21010 14974 21043
rect 14940 20941 14974 20972
rect 14940 20938 14974 20941
rect 14940 20873 14974 20900
rect 14940 20866 14974 20873
rect 14940 20805 14974 20828
rect 14940 20794 14974 20805
rect 14940 20737 14974 20756
rect 14940 20722 14974 20737
rect 14940 20669 14974 20684
rect 14940 20650 14974 20669
rect 14940 20601 14974 20612
rect 14940 20578 14974 20601
rect 14940 20533 14974 20540
rect 14940 20506 14974 20533
rect 14940 20465 14974 20468
rect 14940 20434 14974 20465
rect 14940 20363 14974 20396
rect 14940 20362 14974 20363
rect 14940 20295 14974 20324
rect 14940 20290 14974 20295
rect 14940 20227 14974 20252
rect 14940 20218 14974 20227
rect 14940 20159 14974 20180
rect 14940 20146 14974 20159
rect 14940 20091 14974 20108
rect 14940 20074 14974 20091
rect 14940 20023 14974 20036
rect 14940 20002 14974 20023
rect 14940 19955 14974 19964
rect 14940 19930 14974 19955
rect 14940 19887 14974 19892
rect 14940 19858 14974 19887
rect 14940 19819 14974 19820
rect 14940 19786 14974 19819
rect 14940 19717 14974 19748
rect 14940 19714 14974 19717
rect 14940 19649 14974 19676
rect 14940 19642 14974 19649
rect 14940 19581 14974 19604
rect 14940 19570 14974 19581
rect 14940 19513 14974 19532
rect 14940 19498 14974 19513
rect 14940 19445 14974 19460
rect 14940 19426 14974 19445
rect 14940 19377 14974 19388
rect 14940 19354 14974 19377
rect 14940 19309 14974 19316
rect 14940 19282 14974 19309
rect 14940 19241 14974 19244
rect 14940 19210 14974 19241
rect 14940 19139 14974 19172
rect 14940 19138 14974 19139
rect 14940 19071 14974 19100
rect 14940 19066 14974 19071
rect 14940 19003 14974 19028
rect 14940 18994 14974 19003
rect 14940 18935 14974 18956
rect 14940 18922 14974 18935
rect 14940 18867 14974 18884
rect 14940 18850 14974 18867
rect 14940 18799 14974 18812
rect 14940 18778 14974 18799
rect 14940 18731 14974 18740
rect 14940 18706 14974 18731
rect 14940 18663 14974 18668
rect 14940 18634 14974 18663
rect 14940 18595 14974 18596
rect 14940 18562 14974 18595
rect 14940 18493 14974 18524
rect 14940 18490 14974 18493
rect 14940 18425 14974 18452
rect 14940 18418 14974 18425
rect 14940 18357 14974 18380
rect 14940 18346 14974 18357
rect 14940 18289 14974 18308
rect 14940 18274 14974 18289
rect 14940 18221 14974 18236
rect 14940 18202 14974 18221
rect 14940 18153 14974 18164
rect 14940 18130 14974 18153
rect 14940 18085 14974 18092
rect 14940 18058 14974 18085
rect 14940 18017 14974 18020
rect 14940 17986 14974 18017
rect 14940 17915 14974 17948
rect 14940 17914 14974 17915
rect 14940 17847 14974 17876
rect 14940 17842 14974 17847
rect 14940 17779 14974 17804
rect 14940 17770 14974 17779
rect 14940 17711 14974 17732
rect 14940 17698 14974 17711
rect 14940 17643 14974 17660
rect 14940 17626 14974 17643
rect 14940 17575 14974 17588
rect 14940 17554 14974 17575
rect 14940 17507 14974 17516
rect 14940 17482 14974 17507
rect 14940 17439 14974 17444
rect 14940 17410 14974 17439
rect 14940 17371 14974 17372
rect 14940 17338 14974 17371
rect 14940 17269 14974 17300
rect 14940 17266 14974 17269
rect 14940 17201 14974 17228
rect 14940 17194 14974 17201
rect 14940 17133 14974 17156
rect 14940 17122 14974 17133
rect 14940 17065 14974 17084
rect 14940 17050 14974 17065
rect 14940 16997 14974 17012
rect 14940 16978 14974 16997
rect 14940 16929 14974 16940
rect 14940 16906 14974 16929
rect 14940 16861 14974 16868
rect 14940 16834 14974 16861
rect 14940 16793 14974 16796
rect 14940 16762 14974 16793
rect 14940 16691 14974 16724
rect 14940 16690 14974 16691
rect 14940 16623 14974 16652
rect 14940 16618 14974 16623
rect 14940 16555 14974 16580
rect 14940 16546 14974 16555
rect 14940 16487 14974 16508
rect 14940 16474 14974 16487
rect 14940 16419 14974 16436
rect 14940 16402 14974 16419
rect 14940 16351 14974 16364
rect 14940 16330 14974 16351
rect 14940 16283 14974 16292
rect 14940 16258 14974 16283
rect 14940 16215 14974 16220
rect 14940 16186 14974 16215
rect 14940 16147 14974 16148
rect 14940 16114 14974 16147
rect 14940 16045 14974 16076
rect 14940 16042 14974 16045
rect 14940 15977 14974 16004
rect 14940 15970 14974 15977
rect 14940 15909 14974 15932
rect 14940 15898 14974 15909
rect 14940 15841 14974 15860
rect 14940 15826 14974 15841
rect 14940 15773 14974 15788
rect 14940 15754 14974 15773
rect 14940 15705 14974 15716
rect 14940 15682 14974 15705
rect 14940 15637 14974 15644
rect 14940 15610 14974 15637
rect 14940 15569 14974 15572
rect 14940 15538 14974 15569
rect 14940 15467 14974 15500
rect 14940 15466 14974 15467
rect 14940 15399 14974 15428
rect 14940 15394 14974 15399
rect 14940 15331 14974 15356
rect 14940 15322 14974 15331
rect 14940 15263 14974 15284
rect 14940 15250 14974 15263
rect 14940 15195 14974 15212
rect 14940 15178 14974 15195
rect 14940 15127 14974 15140
rect 14940 15106 14974 15127
rect 14940 15059 14974 15068
rect 14940 15034 14974 15059
rect 14940 14991 14974 14996
rect 14940 14962 14974 14991
rect 14940 14923 14974 14924
rect 14940 14890 14974 14923
rect 14940 14821 14974 14852
rect 14940 14818 14974 14821
rect 14940 14753 14974 14780
rect 14940 14746 14974 14753
rect 14940 14685 14974 14708
rect 14940 14674 14974 14685
rect 14940 14617 14974 14636
rect 14940 14602 14974 14617
rect 14940 14549 14974 14564
rect 14940 14530 14974 14549
rect 14940 14481 14974 14492
rect 14940 14458 14974 14481
rect 14940 14413 14974 14420
rect 14940 14386 14974 14413
rect 14940 14345 14974 14348
rect 14940 14314 14974 14345
rect 14940 14243 14974 14276
rect 14940 14242 14974 14243
rect 14940 14175 14974 14204
rect 14940 14170 14974 14175
rect 14940 14107 14974 14132
rect 14940 14098 14974 14107
rect 14940 14039 14974 14060
rect 14940 14026 14974 14039
rect 14940 13971 14974 13988
rect 14940 13954 14974 13971
rect 14940 13903 14974 13916
rect 14940 13882 14974 13903
rect 14940 13835 14974 13844
rect 14940 13810 14974 13835
rect 14940 13767 14974 13772
rect 14940 13738 14974 13767
rect 14940 13699 14974 13700
rect 14940 13666 14974 13699
rect 14940 13597 14974 13628
rect 14940 13594 14974 13597
rect 14940 13529 14974 13556
rect 14940 13522 14974 13529
rect 14940 13461 14974 13484
rect 14940 13450 14974 13461
rect 14940 13393 14974 13412
rect 14940 13378 14974 13393
rect 14940 13325 14974 13340
rect 14940 13306 14974 13325
rect 14940 13257 14974 13268
rect 14940 13234 14974 13257
rect 14940 13189 14974 13196
rect 14940 13162 14974 13189
rect 14940 13121 14974 13124
rect 14940 13090 14974 13121
rect 14940 13019 14974 13052
rect 14940 13018 14974 13019
rect 14940 12951 14974 12980
rect 14940 12946 14974 12951
rect 14940 12883 14974 12908
rect 14940 12874 14974 12883
rect 14940 12815 14974 12836
rect 14940 12802 14974 12815
rect 14940 12747 14974 12764
rect 14940 12730 14974 12747
rect 14940 12679 14974 12692
rect 14940 12658 14974 12679
rect 14940 12611 14974 12620
rect 14940 12586 14974 12611
rect 14940 12543 14974 12548
rect 14940 12514 14974 12543
rect 14940 12475 14974 12476
rect 14940 12442 14974 12475
rect 14940 12373 14974 12404
rect 14940 12370 14974 12373
rect 14940 12305 14974 12332
rect 14940 12298 14974 12305
rect 14940 12237 14974 12260
rect 14940 12226 14974 12237
rect 14940 12169 14974 12188
rect 14940 12154 14974 12169
rect 14940 12101 14974 12116
rect 14940 12082 14974 12101
rect 14940 12033 14974 12044
rect 14940 12010 14974 12033
rect 14940 11965 14974 11972
rect 14940 11938 14974 11965
rect 14940 11897 14974 11900
rect 14940 11866 14974 11897
rect 14940 11795 14974 11828
rect 14940 11794 14974 11795
rect 14940 11727 14974 11756
rect 14940 11722 14974 11727
rect 14940 11659 14974 11684
rect 14940 11650 14974 11659
rect 14940 11591 14974 11612
rect 14940 11578 14974 11591
rect 14940 11523 14974 11540
rect 14940 11506 14974 11523
rect 14940 11455 14974 11468
rect 14940 11434 14974 11455
rect 14940 11387 14974 11396
rect 14940 11362 14974 11387
rect 14940 11319 14974 11324
rect 14940 11290 14974 11319
rect 14940 11251 14974 11252
rect 14940 11218 14974 11251
rect 14940 11149 14974 11180
rect 14940 11146 14974 11149
rect 14940 11081 14974 11108
rect 14940 11074 14974 11081
rect 14940 11013 14974 11036
rect 14940 11002 14974 11013
rect 14940 10945 14974 10964
rect 14940 10930 14974 10945
rect 14940 10877 14974 10892
rect 14940 10858 14974 10877
rect 14940 10809 14974 10820
rect 14940 10786 14974 10809
rect 14940 10741 14974 10748
rect 14940 10714 14974 10741
rect 14940 10673 14974 10676
rect 14940 10642 14974 10673
rect 14940 10571 14974 10604
rect 14940 10570 14974 10571
rect 14940 10503 14974 10532
rect 14940 10498 14974 10503
rect 14940 10435 14974 10460
rect 14940 10426 14974 10435
rect 14940 10367 14974 10388
rect 14940 10354 14974 10367
rect 14940 10299 14974 10316
rect 14940 10282 14974 10299
rect 14940 10231 14974 10244
rect 14940 10210 14974 10231
rect 14940 10163 14974 10172
rect 14940 10138 14974 10163
rect 14940 10095 14974 10100
rect 14940 10066 14974 10095
rect 14940 10027 14974 10028
rect 14940 9994 14974 10027
rect 14940 9925 14974 9956
rect 14940 9922 14974 9925
rect 14940 9857 14974 9884
rect 14940 9850 14974 9857
rect 14940 9789 14974 9812
rect 14940 9778 14974 9789
rect 14940 9721 14974 9740
rect 14940 9706 14974 9721
rect 14940 9653 14974 9668
rect 14940 9634 14974 9653
rect 14940 9585 14974 9596
rect 14940 9562 14974 9585
rect 14940 9517 14974 9524
rect 14940 9490 14974 9517
rect 14940 9449 14974 9452
rect 14940 9418 14974 9449
rect 14940 9347 14974 9380
rect 14940 9346 14974 9347
rect 14940 9279 14974 9308
rect 14940 9274 14974 9279
rect 14940 9211 14974 9236
rect 14940 9202 14974 9211
rect 14940 9143 14974 9164
rect 14940 9130 14974 9143
rect 14940 9075 14974 9092
rect 14940 9058 14974 9075
rect 14940 9007 14974 9020
rect 14940 8986 14974 9007
rect 14940 8939 14974 8948
rect 14940 8914 14974 8939
rect 14940 8871 14974 8876
rect 14940 8842 14974 8871
rect 14940 8803 14974 8804
rect 14940 8770 14974 8803
rect 14940 8701 14974 8732
rect 14940 8698 14974 8701
rect 14940 8633 14974 8660
rect 14940 8626 14974 8633
rect 14940 8565 14974 8588
rect 14940 8554 14974 8565
rect 14940 8497 14974 8516
rect 14940 8482 14974 8497
rect 14940 8429 14974 8444
rect 14940 8410 14974 8429
rect 14940 8361 14974 8372
rect 14940 8338 14974 8361
rect 14940 8293 14974 8300
rect 14940 8266 14974 8293
rect 14940 8225 14974 8228
rect 14940 8194 14974 8225
rect 14940 8123 14974 8156
rect 14940 8122 14974 8123
rect 14940 8055 14974 8084
rect 14940 8050 14974 8055
rect 14940 7987 14974 8012
rect 14940 7978 14974 7987
rect 14940 7919 14974 7940
rect 14940 7906 14974 7919
rect 14940 7851 14974 7868
rect 14940 7834 14974 7851
rect 14940 7783 14974 7796
rect 14940 7762 14974 7783
rect 14940 7715 14974 7724
rect 14940 7690 14974 7715
rect 14940 7647 14974 7652
rect 14940 7618 14974 7647
rect 14940 7579 14974 7580
rect 14940 7546 14974 7579
rect 14940 7477 14974 7508
rect 14940 7474 14974 7477
rect 14940 7409 14974 7436
rect 14940 7402 14974 7409
rect 14940 7341 14974 7364
rect 14940 7330 14974 7341
rect 14940 7273 14974 7292
rect 14940 7258 14974 7273
rect 14940 7205 14974 7220
rect 14940 7186 14974 7205
rect 14940 7137 14974 7148
rect 14940 7114 14974 7137
rect 14940 7069 14974 7076
rect 14940 7042 14974 7069
rect 14940 7001 14974 7004
rect 14940 6970 14974 7001
rect 14940 6899 14974 6932
rect 14940 6898 14974 6899
rect 14940 6831 14974 6860
rect 14940 6826 14974 6831
rect 14940 6763 14974 6788
rect 14940 6754 14974 6763
rect 14940 6695 14974 6716
rect 14940 6682 14974 6695
rect 14940 6627 14974 6644
rect 14940 6610 14974 6627
rect 14940 6559 14974 6572
rect 14940 6538 14974 6559
rect 14940 6491 14974 6500
rect 14940 6466 14974 6491
rect 14940 6423 14974 6428
rect 14940 6394 14974 6423
rect 14940 6355 14974 6356
rect 14940 6322 14974 6355
rect 14940 6253 14974 6284
rect 14940 6250 14974 6253
rect 14940 6185 14974 6212
rect 14940 6178 14974 6185
rect 14940 6117 14974 6140
rect 14940 6106 14974 6117
rect 14940 6049 14974 6068
rect 14940 6034 14974 6049
rect 14940 5981 14974 5996
rect 14940 5962 14974 5981
rect 14940 5913 14974 5924
rect 14940 5890 14974 5913
rect 14940 5845 14974 5852
rect 14940 5818 14974 5845
rect 14940 5777 14974 5780
rect 14940 5746 14974 5777
rect 14940 5675 14974 5708
rect 14940 5674 14974 5675
rect 14940 5607 14974 5636
rect 14940 5602 14974 5607
rect 14940 5539 14974 5564
rect 14940 5530 14974 5539
rect 14940 5471 14974 5492
rect 14940 5458 14974 5471
rect 14940 5403 14974 5420
rect 14940 5386 14974 5403
rect 14940 5335 14974 5348
rect 14940 5314 14974 5335
rect 14940 5267 14974 5276
rect 14940 5242 14974 5267
rect 14940 5199 14974 5204
rect 14940 5170 14974 5199
rect 14940 5131 14974 5132
rect 14940 5098 14974 5131
rect 14940 5029 14974 5060
rect 14940 5026 14974 5029
rect 14940 4961 14974 4988
rect 14940 4954 14974 4961
rect 14940 4893 14974 4916
rect 14940 4882 14974 4893
rect 14940 4825 14974 4844
rect 14940 4810 14974 4825
rect 14940 4757 14974 4772
rect 14940 4738 14974 4757
rect 14940 4689 14974 4700
rect 14940 4666 14974 4689
rect 14940 4621 14974 4628
rect 14940 4594 14974 4621
rect 14940 4553 14974 4556
rect 14940 4522 14974 4553
rect 14940 4451 14974 4484
rect 14940 4450 14974 4451
rect 14940 4383 14974 4412
rect 14940 4378 14974 4383
rect 14940 4315 14974 4340
rect 14940 4306 14974 4315
rect 14940 4247 14974 4268
rect 14940 4234 14974 4247
rect 14940 4179 14974 4196
rect 14940 4162 14974 4179
rect 14940 4111 14974 4124
rect 14940 4090 14974 4111
rect 14940 4043 14974 4052
rect 14940 4018 14974 4043
rect 14940 3975 14974 3980
rect 14940 3946 14974 3975
rect 14940 3907 14974 3908
rect 14940 3874 14974 3907
rect 14940 3805 14974 3836
rect 14940 3802 14974 3805
rect 14940 3737 14974 3764
rect 14940 3730 14974 3737
rect 14940 3669 14974 3692
rect 14940 3658 14974 3669
rect 14940 3601 14974 3620
rect 14940 3586 14974 3601
rect 14940 3533 14974 3548
rect 14940 3514 14974 3533
rect 14940 3465 14974 3476
rect 14940 3442 14974 3465
rect 14940 3397 14974 3404
rect 14940 3370 14974 3397
rect 14940 3329 14974 3332
rect 14940 3298 14974 3329
rect 14940 3226 14974 3260
rect 14940 3171 14974 3188
rect 14940 3154 14974 3171
rect 14940 3103 14974 3116
rect 14940 3082 14974 3103
rect 14940 3035 14974 3044
rect 14940 3010 14974 3035
rect 14940 2967 14974 2972
rect 14940 2938 14974 2967
rect 14940 2899 14974 2900
rect 14940 2866 14974 2899
rect 14940 2797 14974 2828
rect 14940 2794 14974 2797
rect 14940 2729 14974 2756
rect 14940 2722 14974 2729
rect 14940 2661 14974 2684
rect 14940 2650 14974 2661
rect 14940 2593 14974 2612
rect 14940 2578 14974 2593
rect 14940 2525 14974 2540
rect 14940 2506 14974 2525
rect 14940 2457 14974 2468
rect 14940 2434 14974 2457
rect 14940 2389 14974 2396
rect 14940 2362 14974 2389
rect 14940 2321 14974 2324
rect 14940 2290 14974 2321
rect 14940 2219 14974 2252
rect 14940 2218 14974 2219
rect 14940 2151 14974 2180
rect 14940 2146 14974 2151
rect 14940 2083 14974 2108
rect 14940 2074 14974 2083
rect 14940 2015 14974 2036
rect 14940 2002 14974 2015
rect 14940 1947 14974 1964
rect 14940 1930 14974 1947
rect 14940 1879 14974 1892
rect 14940 1858 14974 1879
rect 14940 1811 14974 1820
rect 14940 1786 14974 1811
rect 14940 1743 14974 1748
rect 14940 1714 14974 1743
rect 14940 1675 14974 1676
rect 14940 1642 14974 1675
rect 14940 1573 14974 1604
rect 14940 1570 14974 1573
rect 14940 1505 14974 1532
rect 14940 1498 14974 1505
rect 14940 1437 14974 1460
rect 14940 1426 14974 1437
rect 14940 1369 14974 1387
rect 14940 1353 14974 1369
rect 14940 1301 14974 1314
rect 14940 1280 14974 1301
rect 14940 1233 14974 1241
rect 14940 1207 14974 1233
rect 14940 1165 14974 1168
rect 14940 1134 14974 1165
rect 14940 1063 14974 1095
rect 14940 1061 14974 1063
rect 14940 995 14974 1022
rect 14940 988 14974 995
rect 14940 927 14974 949
rect 14940 915 14974 927
rect 14940 859 14974 876
rect 14940 842 14974 859
rect 14940 791 14974 803
rect 14940 769 14974 791
rect 14940 723 14974 730
rect 14940 696 14974 723
rect 14940 655 14974 657
rect 14940 623 14974 655
rect 14940 553 14974 584
rect 14940 550 14974 553
rect 14940 485 14974 511
rect 14940 477 14974 485
rect 11610 311 11644 325
rect 13212 346 13246 362
rect 13212 328 13246 346
rect 14817 383 14851 417
rect 14817 325 14851 345
rect 11424 213 11458 220
rect 11424 186 11458 213
rect 11424 145 11458 147
rect 11424 113 11458 145
rect 14648 290 14682 324
rect 14720 291 14730 324
rect 14730 291 14754 324
rect 14817 311 14848 325
rect 14848 311 14851 325
rect 14940 417 14974 438
rect 14940 404 14974 417
rect 14940 349 14974 365
rect 14940 331 14974 349
rect 14720 290 14754 291
rect 13212 278 13246 290
rect 13212 256 13246 278
rect 13212 210 13246 218
rect 13212 184 13246 210
rect 13212 142 13246 146
rect 13212 112 13246 142
rect 14940 281 14974 292
rect 14940 258 14974 281
rect 14940 213 14974 219
rect 14940 185 14974 213
rect 14940 145 14974 146
rect 14940 112 14974 145
rect 11496 40 11526 74
rect 11526 40 11530 74
rect 11570 40 11594 74
rect 11594 40 11604 74
rect 11644 40 11662 74
rect 11662 40 11678 74
rect 11718 40 11730 74
rect 11730 40 11752 74
rect 11792 40 11798 74
rect 11798 40 11826 74
rect 11866 40 11900 74
rect 11940 40 11968 74
rect 11968 40 11974 74
rect 12014 40 12036 74
rect 12036 40 12048 74
rect 12088 40 12104 74
rect 12104 40 12122 74
rect 12162 40 12172 74
rect 12172 40 12196 74
rect 12236 40 12240 74
rect 12240 40 12270 74
rect 12310 40 12342 74
rect 12342 40 12344 74
rect 12384 40 12410 74
rect 12410 40 12418 74
rect 12458 40 12478 74
rect 12478 40 12492 74
rect 12531 40 12546 74
rect 12546 40 12565 74
rect 12604 40 12614 74
rect 12614 40 12638 74
rect 12677 40 12682 74
rect 12682 40 12711 74
rect 12750 40 12784 74
rect 12823 40 12852 74
rect 12852 40 12857 74
rect 12896 40 12920 74
rect 12920 40 12930 74
rect 12969 40 12988 74
rect 12988 40 13003 74
rect 13042 40 13056 74
rect 13056 40 13076 74
rect 13115 40 13124 74
rect 13124 40 13149 74
rect 13188 40 13222 74
rect 13261 40 13295 74
rect 13334 40 13342 74
rect 13342 40 13368 74
rect 13407 40 13410 74
rect 13410 40 13441 74
rect 13480 40 13512 74
rect 13512 40 13514 74
rect 13553 40 13580 74
rect 13580 40 13587 74
rect 13626 40 13648 74
rect 13648 40 13660 74
rect 13699 40 13716 74
rect 13716 40 13733 74
rect 13772 40 13784 74
rect 13784 40 13806 74
rect 13845 40 13852 74
rect 13852 40 13879 74
rect 13918 40 13920 74
rect 13920 40 13952 74
rect 13991 40 14022 74
rect 14022 40 14025 74
rect 14064 40 14090 74
rect 14090 40 14098 74
rect 14137 40 14158 74
rect 14158 40 14171 74
rect 14210 40 14226 74
rect 14226 40 14244 74
rect 14283 40 14294 74
rect 14294 40 14317 74
rect 14356 40 14362 74
rect 14362 40 14390 74
rect 14429 40 14430 74
rect 14430 40 14463 74
rect 14502 40 14532 74
rect 14532 40 14536 74
rect 14575 40 14600 74
rect 14600 40 14609 74
rect 14648 40 14668 74
rect 14668 40 14682 74
rect 14721 40 14736 74
rect 14736 40 14755 74
rect 14794 40 14804 74
rect 14804 40 14828 74
rect 14867 40 14872 74
rect 14872 40 14901 74
rect 11607 -189 11631 -155
rect 11631 -189 11641 -155
rect 11679 -189 11699 -155
rect 11699 -189 11713 -155
rect 11751 -189 11767 -155
rect 11767 -189 11785 -155
rect 11823 -189 11835 -155
rect 11835 -189 11857 -155
rect 11896 -189 11903 -155
rect 11903 -189 11930 -155
rect 11969 -189 11971 -155
rect 11971 -189 12003 -155
rect 12042 -189 12073 -155
rect 12073 -189 12076 -155
rect 12115 -189 12141 -155
rect 12141 -189 12149 -155
rect 12188 -189 12209 -155
rect 12209 -189 12222 -155
rect 12261 -189 12277 -155
rect 12277 -189 12295 -155
rect 12334 -189 12345 -155
rect 12345 -189 12368 -155
rect 12407 -189 12413 -155
rect 12413 -189 12441 -155
rect 12480 -189 12481 -155
rect 12481 -189 12514 -155
rect 12553 -189 12583 -155
rect 12583 -189 12587 -155
rect 12626 -189 12651 -155
rect 12651 -189 12660 -155
rect 12699 -189 12719 -155
rect 12719 -189 12733 -155
rect 12772 -189 12787 -155
rect 12787 -189 12806 -155
rect 12845 -189 12856 -155
rect 12856 -189 12879 -155
rect 12918 -189 12925 -155
rect 12925 -189 12952 -155
rect 12991 -189 12994 -155
rect 12994 -189 13025 -155
rect 13064 -189 13097 -155
rect 13097 -189 13098 -155
rect 13137 -189 13166 -155
rect 13166 -189 13171 -155
rect 13210 -189 13235 -155
rect 13235 -189 13244 -155
rect 13283 -189 13304 -155
rect 13304 -189 13317 -155
rect 13356 -189 13373 -155
rect 13373 -189 13390 -155
rect 13429 -189 13442 -155
rect 13442 -189 13463 -155
rect 13502 -189 13511 -155
rect 13511 -189 13536 -155
rect 13575 -189 13580 -155
rect 13580 -189 13609 -155
rect 13648 -189 13649 -155
rect 13649 -189 13682 -155
rect 13721 -189 13753 -155
rect 13753 -189 13755 -155
rect 13794 -189 13822 -155
rect 13822 -189 13828 -155
rect 13867 -189 13891 -155
rect 13891 -189 13901 -155
rect 13940 -189 13960 -155
rect 13960 -189 13974 -155
rect 14013 -189 14029 -155
rect 14029 -189 14047 -155
rect 14086 -189 14098 -155
rect 14098 -189 14120 -155
rect 14159 -189 14167 -155
rect 14167 -189 14193 -155
rect 14232 -189 14236 -155
rect 14236 -189 14266 -155
rect 14305 -189 14339 -155
rect 14378 -189 14408 -155
rect 14408 -189 14412 -155
rect 14451 -189 14477 -155
rect 14477 -189 14485 -155
rect 14524 -189 14546 -155
rect 14546 -189 14558 -155
rect 14597 -189 14615 -155
rect 14615 -189 14631 -155
rect 14670 -189 14684 -155
rect 14684 -189 14704 -155
rect 14743 -189 14753 -155
rect 14753 -189 14777 -155
rect 11771 -300 11805 -266
rect 11771 -382 11805 -348
rect 11615 -432 11649 -398
rect 11615 -507 11649 -473
rect 11615 -582 11649 -548
rect 11615 -657 11649 -623
rect 11615 -732 11649 -698
rect 12083 -300 12117 -266
rect 12083 -382 12117 -348
rect 11771 -464 11805 -430
rect 11771 -546 11805 -512
rect 11771 -628 11805 -594
rect 11771 -711 11805 -677
rect 11927 -432 11961 -398
rect 11927 -507 11961 -473
rect 11927 -582 11961 -548
rect 11927 -657 11961 -623
rect 11615 -807 11649 -773
rect 11927 -732 11961 -698
rect 12395 -300 12429 -266
rect 12395 -382 12429 -348
rect 12083 -464 12117 -430
rect 12083 -546 12117 -512
rect 12083 -628 12117 -594
rect 12083 -711 12117 -677
rect 12239 -432 12273 -398
rect 12239 -507 12273 -473
rect 12239 -582 12273 -548
rect 12239 -657 12273 -623
rect 11927 -807 11961 -773
rect 12239 -732 12273 -698
rect 12707 -300 12741 -266
rect 12707 -382 12741 -348
rect 12395 -464 12429 -430
rect 12395 -546 12429 -512
rect 12395 -628 12429 -594
rect 12395 -711 12429 -677
rect 12551 -432 12585 -398
rect 12551 -507 12585 -473
rect 12551 -582 12585 -548
rect 12551 -657 12585 -623
rect 12239 -807 12273 -773
rect 12551 -732 12585 -698
rect 13018 -300 13052 -266
rect 13018 -382 13052 -348
rect 12707 -464 12741 -430
rect 12707 -546 12741 -512
rect 12707 -628 12741 -594
rect 12707 -711 12741 -677
rect 12863 -432 12897 -398
rect 12863 -507 12897 -473
rect 12863 -582 12897 -548
rect 12863 -657 12897 -623
rect 12551 -807 12585 -773
rect 12863 -732 12897 -698
rect 13331 -300 13365 -266
rect 13331 -382 13365 -348
rect 13018 -464 13052 -430
rect 13018 -546 13052 -512
rect 13018 -628 13052 -594
rect 13018 -711 13052 -677
rect 13175 -432 13209 -398
rect 13175 -507 13209 -473
rect 13175 -582 13209 -548
rect 13175 -657 13209 -623
rect 12863 -807 12897 -773
rect 13175 -732 13209 -698
rect 13643 -300 13677 -266
rect 13643 -382 13677 -348
rect 13331 -464 13365 -430
rect 13331 -546 13365 -512
rect 13331 -628 13365 -594
rect 13331 -711 13365 -677
rect 13487 -432 13521 -398
rect 13487 -507 13521 -473
rect 13487 -582 13521 -548
rect 13487 -657 13521 -623
rect 13175 -807 13209 -773
rect 13487 -732 13521 -698
rect 13955 -300 13989 -266
rect 13955 -382 13989 -348
rect 13643 -464 13677 -430
rect 13643 -546 13677 -512
rect 13643 -628 13677 -594
rect 13643 -711 13677 -677
rect 13799 -432 13833 -398
rect 13799 -507 13833 -473
rect 13799 -582 13833 -548
rect 13799 -657 13833 -623
rect 13487 -807 13521 -773
rect 13799 -732 13833 -698
rect 14267 -300 14301 -266
rect 14267 -382 14301 -348
rect 13955 -464 13989 -430
rect 13955 -546 13989 -512
rect 13955 -628 13989 -594
rect 13955 -711 13989 -677
rect 14111 -432 14145 -398
rect 14111 -507 14145 -473
rect 14111 -582 14145 -548
rect 14111 -657 14145 -623
rect 13799 -807 13833 -773
rect 14111 -732 14145 -698
rect 14579 -300 14613 -266
rect 14579 -382 14613 -348
rect 14267 -464 14301 -430
rect 14267 -546 14301 -512
rect 14267 -628 14301 -594
rect 14267 -711 14301 -677
rect 14423 -432 14457 -398
rect 14423 -507 14457 -473
rect 14423 -582 14457 -548
rect 14423 -657 14457 -623
rect 14111 -807 14145 -773
rect 14423 -732 14457 -698
rect 14579 -464 14613 -430
rect 14579 -546 14613 -512
rect 14579 -628 14613 -594
rect 14579 -711 14613 -677
rect 14735 -396 14769 -362
rect 14735 -478 14769 -444
rect 14735 -560 14769 -526
rect 14735 -642 14769 -608
rect 14423 -807 14457 -773
rect 14735 -724 14769 -690
rect 14735 -807 14769 -773
rect 11690 -951 11710 -917
rect 11710 -951 11724 -917
rect 11762 -951 11778 -917
rect 11778 -951 11796 -917
rect 11834 -951 11846 -917
rect 11846 -951 11868 -917
rect 11906 -951 11914 -917
rect 11914 -951 11940 -917
rect 11978 -951 11982 -917
rect 11982 -951 12012 -917
rect 12050 -951 12084 -917
rect 12123 -951 12152 -917
rect 12152 -951 12157 -917
rect 12196 -951 12220 -917
rect 12220 -951 12230 -917
rect 12269 -951 12288 -917
rect 12288 -951 12303 -917
rect 12342 -951 12356 -917
rect 12356 -951 12376 -917
rect 12415 -951 12424 -917
rect 12424 -951 12449 -917
rect 12488 -951 12492 -917
rect 12492 -951 12522 -917
rect 12561 -951 12594 -917
rect 12594 -951 12595 -917
rect 12634 -951 12662 -917
rect 12662 -951 12668 -917
rect 12707 -951 12730 -917
rect 12730 -951 12741 -917
rect 12780 -951 12798 -917
rect 12798 -951 12814 -917
rect 12853 -951 12866 -917
rect 12866 -951 12887 -917
rect 12926 -951 12934 -917
rect 12934 -951 12960 -917
rect 12999 -951 13002 -917
rect 13002 -951 13033 -917
rect 13072 -951 13104 -917
rect 13104 -951 13106 -917
rect 13145 -951 13172 -917
rect 13172 -951 13179 -917
rect 13218 -951 13240 -917
rect 13240 -951 13252 -917
rect 13291 -951 13308 -917
rect 13308 -951 13325 -917
rect 13364 -951 13376 -917
rect 13376 -951 13398 -917
rect 13437 -951 13444 -917
rect 13444 -951 13471 -917
rect 13510 -951 13512 -917
rect 13512 -951 13544 -917
rect 13583 -951 13614 -917
rect 13614 -951 13617 -917
rect 13656 -951 13682 -917
rect 13682 -951 13690 -917
rect 13729 -951 13750 -917
rect 13750 -951 13763 -917
rect 13802 -951 13818 -917
rect 13818 -951 13836 -917
rect 13875 -951 13886 -917
rect 13886 -951 13909 -917
rect 13948 -951 13954 -917
rect 13954 -951 13982 -917
rect 14021 -951 14022 -917
rect 14022 -951 14055 -917
rect 14094 -951 14124 -917
rect 14124 -951 14128 -917
rect 14167 -951 14192 -917
rect 14192 -951 14201 -917
rect 14240 -951 14260 -917
rect 14260 -951 14274 -917
rect 14313 -951 14329 -917
rect 14329 -951 14347 -917
rect 14386 -951 14398 -917
rect 14398 -951 14420 -917
rect 14459 -951 14467 -917
rect 14467 -951 14493 -917
rect 14532 -951 14536 -917
rect 14536 -951 14566 -917
rect 14605 -951 14639 -917
rect 14678 -951 14708 -917
rect 14708 -951 14712 -917
<< metal1 >>
rect -258 38757 6154 38763
rect -258 38723 -176 38757
rect -142 38723 -99 38757
rect -65 38723 11 38757
rect 45 38723 83 38757
rect 117 38723 155 38757
rect 189 38723 227 38757
rect 261 38723 299 38757
rect 333 38723 371 38757
rect 405 38723 443 38757
rect 477 38723 515 38757
rect 549 38723 587 38757
rect 621 38723 659 38757
rect 693 38723 731 38757
rect 765 38723 803 38757
rect 837 38723 875 38757
rect 909 38723 947 38757
rect 981 38723 1019 38757
rect 1053 38723 1091 38757
rect 1125 38723 1163 38757
rect 1197 38723 1235 38757
rect 1269 38723 1307 38757
rect 1341 38723 1379 38757
rect 1413 38723 1451 38757
rect 1485 38723 1523 38757
rect 1557 38723 1595 38757
rect 1629 38723 1667 38757
rect 1701 38723 1739 38757
rect 1773 38723 1811 38757
rect 1845 38723 1883 38757
rect 1917 38723 1955 38757
rect 1989 38723 2027 38757
rect 2061 38723 2100 38757
rect 2134 38723 2173 38757
rect 2207 38723 2246 38757
rect 2280 38723 2319 38757
rect 2353 38723 2392 38757
rect 2426 38723 2465 38757
rect 2499 38723 2538 38757
rect 2572 38723 2611 38757
rect 2645 38723 2684 38757
rect 2718 38723 2757 38757
rect 2791 38723 2830 38757
rect 2864 38723 2903 38757
rect 2937 38723 2976 38757
rect 3010 38723 3049 38757
rect 3083 38723 3122 38757
rect 3156 38723 3195 38757
rect 3229 38723 3268 38757
rect 3302 38723 3341 38757
rect 3375 38723 3414 38757
rect 3448 38723 3487 38757
rect 3521 38723 3560 38757
rect 3594 38723 3633 38757
rect 3667 38723 3706 38757
rect 3740 38723 3779 38757
rect 3813 38723 3852 38757
rect 3886 38723 3925 38757
rect 3959 38723 3998 38757
rect 4032 38723 4071 38757
rect 4105 38723 4144 38757
rect 4178 38723 4217 38757
rect 4251 38723 4290 38757
rect 4324 38723 4363 38757
rect 4397 38723 4436 38757
rect 4470 38723 4509 38757
rect 4543 38723 4582 38757
rect 4616 38723 4655 38757
rect 4689 38723 4728 38757
rect 4762 38723 4801 38757
rect 4835 38723 4874 38757
rect 4908 38723 4947 38757
rect 4981 38723 5020 38757
rect 5054 38723 5093 38757
rect 5127 38723 5166 38757
rect 5200 38723 5239 38757
rect 5273 38723 5312 38757
rect 5346 38723 5385 38757
rect 5419 38723 5458 38757
rect 5492 38723 5531 38757
rect 5565 38723 5604 38757
rect 5638 38723 5677 38757
rect 5711 38723 5750 38757
rect 5784 38723 5823 38757
rect 5857 38723 5896 38757
rect 5930 38723 5969 38757
rect 6003 38723 6042 38757
rect 6076 38723 6154 38757
rect -258 38717 6154 38723
rect -258 38685 -210 38717
tri -210 38685 -178 38717 nw
tri 1790 38685 1822 38717 ne
rect 1822 38685 1872 38717
tri 1872 38685 1904 38717 nw
tri 3932 38685 3964 38717 ne
rect 3964 38685 4014 38717
tri 4014 38685 4046 38717 nw
tri 6074 38685 6106 38717 ne
rect 6106 38685 6154 38717
rect -258 38651 -252 38685
rect -218 38651 -212 38685
tri -212 38683 -210 38685 nw
tri 1822 38683 1824 38685 ne
rect -258 38612 -212 38651
rect -258 38578 -252 38612
rect -218 38578 -212 38612
rect -258 38539 -212 38578
rect -258 38505 -252 38539
rect -218 38505 -212 38539
rect -258 38466 -212 38505
rect -258 38432 -252 38466
rect -218 38432 -212 38466
rect -258 38393 -212 38432
rect -258 38359 -252 38393
rect -218 38359 -212 38393
rect -258 38320 -212 38359
rect -258 38286 -252 38320
rect -218 38286 -212 38320
rect -258 38247 -212 38286
rect -258 38213 -252 38247
rect -218 38213 -212 38247
rect -258 38174 -212 38213
rect -258 38140 -252 38174
rect -218 38140 -212 38174
rect -258 38101 -212 38140
rect -258 38067 -252 38101
rect -218 38067 -212 38101
rect -258 38028 -212 38067
rect -258 37994 -252 38028
rect -218 37994 -212 38028
rect -258 37955 -212 37994
rect -258 37921 -252 37955
rect -218 37921 -212 37955
rect -258 37882 -212 37921
rect -258 37848 -252 37882
rect -218 37848 -212 37882
rect -258 37809 -212 37848
rect -258 37775 -252 37809
rect -218 37775 -212 37809
rect -258 37736 -212 37775
rect -258 37702 -252 37736
rect -218 37702 -212 37736
rect -258 37663 -212 37702
rect -258 37629 -252 37663
rect -218 37629 -212 37663
rect -258 37590 -212 37629
rect -258 37556 -252 37590
rect -218 37556 -212 37590
rect -258 37517 -212 37556
rect -258 37483 -252 37517
rect -218 37483 -212 37517
rect -258 37444 -212 37483
rect -258 37410 -252 37444
rect -218 37410 -212 37444
rect -258 37371 -212 37410
rect -258 37337 -252 37371
rect -218 37337 -212 37371
rect -258 37298 -212 37337
rect -258 37264 -252 37298
rect -218 37264 -212 37298
rect -258 37225 -212 37264
rect -258 37191 -252 37225
rect -218 37191 -212 37225
rect -258 37152 -212 37191
rect -258 37118 -252 37152
rect -218 37118 -212 37152
rect -258 37079 -212 37118
rect -258 37045 -252 37079
rect -218 37045 -212 37079
rect -258 37006 -212 37045
rect -258 36972 -252 37006
rect -218 36972 -212 37006
rect -258 36933 -212 36972
rect -258 36899 -252 36933
rect -218 36899 -212 36933
rect -258 36860 -212 36899
rect -258 36826 -252 36860
rect -218 36826 -212 36860
rect -258 36787 -212 36826
rect -258 36753 -252 36787
rect -218 36753 -212 36787
rect -258 36714 -212 36753
rect -258 36680 -252 36714
rect -218 36680 -212 36714
rect -258 36641 -212 36680
rect -258 36607 -252 36641
rect -218 36607 -212 36641
rect -258 36568 -212 36607
rect -258 36534 -252 36568
rect -218 36534 -212 36568
rect -258 36495 -212 36534
rect -258 36461 -252 36495
rect -218 36461 -212 36495
rect -258 36422 -212 36461
rect -258 36388 -252 36422
rect -218 36388 -212 36422
rect -258 36349 -212 36388
rect -258 36315 -252 36349
rect -218 36315 -212 36349
rect -258 36276 -212 36315
rect -258 36242 -252 36276
rect -218 36242 -212 36276
rect -258 36203 -212 36242
rect -258 36169 -252 36203
rect -218 36169 -212 36203
rect -258 36130 -212 36169
rect -258 36096 -252 36130
rect -218 36096 -212 36130
rect -258 36057 -212 36096
rect -258 36023 -252 36057
rect -218 36023 -212 36057
rect -258 35984 -212 36023
rect -258 35950 -252 35984
rect -218 35950 -212 35984
rect -258 35911 -212 35950
rect -258 35877 -252 35911
rect -218 35877 -212 35911
rect -258 35838 -212 35877
rect -258 35804 -252 35838
rect -218 35804 -212 35838
rect -258 35765 -212 35804
rect -258 35731 -252 35765
rect -218 35731 -212 35765
rect -258 35692 -212 35731
rect -258 35658 -252 35692
rect -218 35658 -212 35692
rect -258 35619 -212 35658
rect -258 35585 -252 35619
rect -218 35585 -212 35619
rect -258 35546 -212 35585
rect -258 35512 -252 35546
rect -218 35512 -212 35546
rect -258 35473 -212 35512
rect -258 35439 -252 35473
rect -218 35439 -212 35473
rect -258 35400 -212 35439
rect -258 35366 -252 35400
rect -218 35366 -212 35400
rect -258 35327 -212 35366
rect -258 35293 -252 35327
rect -218 35293 -212 35327
rect -258 35254 -212 35293
rect -258 35220 -252 35254
rect -218 35220 -212 35254
rect -258 35181 -212 35220
rect -258 35147 -252 35181
rect -218 35147 -212 35181
rect -258 35109 -212 35147
rect -258 35075 -252 35109
rect -218 35075 -212 35109
rect -258 35037 -212 35075
rect -258 35003 -252 35037
rect -218 35003 -212 35037
rect -258 34965 -212 35003
rect -258 34931 -252 34965
rect -218 34931 -212 34965
rect -258 34893 -212 34931
rect -258 34859 -252 34893
rect -218 34859 -212 34893
rect -258 34821 -212 34859
rect -258 34787 -252 34821
rect -218 34787 -212 34821
rect -258 34749 -212 34787
rect -258 34715 -252 34749
rect -218 34715 -212 34749
rect -258 34677 -212 34715
rect -258 34643 -252 34677
rect -218 34643 -212 34677
rect -258 34605 -212 34643
rect -258 34571 -252 34605
rect -218 34571 -212 34605
rect -258 34533 -212 34571
rect -258 34499 -252 34533
rect -218 34499 -212 34533
rect -258 34461 -212 34499
rect -258 34427 -252 34461
rect -218 34427 -212 34461
rect -258 34389 -212 34427
rect -258 34355 -252 34389
rect -218 34355 -212 34389
rect -258 34317 -212 34355
rect -258 34283 -252 34317
rect -218 34283 -212 34317
rect -258 34245 -212 34283
rect -258 34211 -252 34245
rect -218 34211 -212 34245
rect -258 34173 -212 34211
rect -258 34139 -252 34173
rect -218 34139 -212 34173
rect -258 34101 -212 34139
rect -258 34067 -252 34101
rect -218 34067 -212 34101
rect -258 34029 -212 34067
rect -258 33995 -252 34029
rect -218 33995 -212 34029
rect -258 33957 -212 33995
rect -258 33923 -252 33957
rect -218 33923 -212 33957
rect -258 33885 -212 33923
rect -258 33851 -252 33885
rect -218 33851 -212 33885
rect -258 33813 -212 33851
rect -258 33779 -252 33813
rect -218 33779 -212 33813
rect -258 33741 -212 33779
rect -258 33707 -252 33741
rect -218 33707 -212 33741
rect -258 33669 -212 33707
rect -258 33635 -252 33669
rect -218 33635 -212 33669
rect -258 33597 -212 33635
rect -258 33563 -252 33597
rect -218 33563 -212 33597
rect -258 33525 -212 33563
rect -258 33491 -252 33525
rect -218 33491 -212 33525
rect -258 33453 -212 33491
rect -258 33419 -252 33453
rect -218 33419 -212 33453
rect -258 33381 -212 33419
rect -258 33347 -252 33381
rect -218 33347 -212 33381
rect -258 33309 -212 33347
rect -258 33275 -252 33309
rect -218 33275 -212 33309
rect -258 33237 -212 33275
rect -258 33203 -252 33237
rect -218 33203 -212 33237
rect -258 33165 -212 33203
rect -258 33131 -252 33165
rect -218 33131 -212 33165
rect -258 33093 -212 33131
rect -258 33059 -252 33093
rect -218 33059 -212 33093
rect -258 33021 -212 33059
rect -258 32987 -252 33021
rect -218 32987 -212 33021
rect -258 32949 -212 32987
rect -258 32915 -252 32949
rect -218 32915 -212 32949
rect -258 32877 -212 32915
rect -258 32843 -252 32877
rect -218 32843 -212 32877
rect -258 32805 -212 32843
rect -258 32771 -252 32805
rect -218 32771 -212 32805
rect -258 32733 -212 32771
rect -258 32699 -252 32733
rect -218 32699 -212 32733
rect -258 32661 -212 32699
rect -258 32627 -252 32661
rect -218 32627 -212 32661
rect -258 32589 -212 32627
rect -258 32555 -252 32589
rect -218 32555 -212 32589
rect -258 32517 -212 32555
rect -258 32483 -252 32517
rect -218 32483 -212 32517
rect -258 32445 -212 32483
rect -258 32411 -252 32445
rect -218 32411 -212 32445
rect -258 32373 -212 32411
rect -258 32339 -252 32373
rect -218 32339 -212 32373
rect -258 32301 -212 32339
rect -258 32267 -252 32301
rect -218 32267 -212 32301
rect -258 32229 -212 32267
rect -258 32195 -252 32229
rect -218 32195 -212 32229
rect -258 32157 -212 32195
rect -258 32123 -252 32157
rect -218 32123 -212 32157
rect -258 32085 -212 32123
rect -258 32051 -252 32085
rect -218 32051 -212 32085
rect -258 32013 -212 32051
rect -258 31979 -252 32013
rect -218 31979 -212 32013
rect -258 31941 -212 31979
rect -258 31907 -252 31941
rect -218 31907 -212 31941
rect -258 31869 -212 31907
rect -258 31835 -252 31869
rect -218 31835 -212 31869
rect -258 31797 -212 31835
rect -258 31763 -252 31797
rect -218 31763 -212 31797
rect -258 31725 -212 31763
rect -258 31691 -252 31725
rect -218 31691 -212 31725
rect -258 31653 -212 31691
rect -258 31619 -252 31653
rect -218 31619 -212 31653
rect -258 31581 -212 31619
rect -258 31547 -252 31581
rect -218 31547 -212 31581
rect -258 31509 -212 31547
rect -258 31475 -252 31509
rect -218 31475 -212 31509
rect -258 31437 -212 31475
rect -258 31403 -252 31437
rect -218 31403 -212 31437
rect -258 31365 -212 31403
rect -258 31331 -252 31365
rect -218 31331 -212 31365
rect -258 31293 -212 31331
rect -258 31259 -252 31293
rect -218 31259 -212 31293
rect -258 31221 -212 31259
rect -258 31187 -252 31221
rect -218 31187 -212 31221
rect -258 31149 -212 31187
rect -258 31115 -252 31149
rect -218 31115 -212 31149
rect -258 31077 -212 31115
rect -258 31043 -252 31077
rect -218 31043 -212 31077
rect -258 31005 -212 31043
rect -258 30971 -252 31005
rect -218 30971 -212 31005
rect -258 30933 -212 30971
rect -258 30899 -252 30933
rect -218 30899 -212 30933
rect -258 30861 -212 30899
rect -258 30827 -252 30861
rect -218 30827 -212 30861
rect -258 30789 -212 30827
rect -258 30755 -252 30789
rect -218 30755 -212 30789
rect -258 30717 -212 30755
rect -258 30683 -252 30717
rect -218 30683 -212 30717
rect -258 30645 -212 30683
rect -258 30611 -252 30645
rect -218 30611 -212 30645
rect -258 30573 -212 30611
rect -258 30539 -252 30573
rect -218 30539 -212 30573
rect -258 30501 -212 30539
rect -258 30467 -252 30501
rect -218 30467 -212 30501
rect -258 30429 -212 30467
rect -258 30395 -252 30429
rect -218 30395 -212 30429
rect -258 30357 -212 30395
rect -258 30323 -252 30357
rect -218 30323 -212 30357
rect -258 30285 -212 30323
rect -258 30251 -252 30285
rect -218 30251 -212 30285
rect -258 30213 -212 30251
rect -258 30179 -252 30213
rect -218 30179 -212 30213
rect -258 30141 -212 30179
rect -258 30107 -252 30141
rect -218 30107 -212 30141
rect -258 30069 -212 30107
rect -258 30035 -252 30069
rect -218 30035 -212 30069
rect -258 29997 -212 30035
rect -258 29963 -252 29997
rect -218 29963 -212 29997
rect -258 29925 -212 29963
rect -258 29891 -252 29925
rect -218 29891 -212 29925
rect -258 29853 -212 29891
rect -258 29819 -252 29853
rect -218 29819 -212 29853
rect -258 29781 -212 29819
rect -258 29747 -252 29781
rect -218 29747 -212 29781
rect -258 29709 -212 29747
rect -258 29675 -252 29709
rect -218 29675 -212 29709
rect -258 29637 -212 29675
rect -258 29603 -252 29637
rect -218 29603 -212 29637
rect -258 29565 -212 29603
rect -258 29531 -252 29565
rect -218 29531 -212 29565
rect -258 29493 -212 29531
rect -258 29459 -252 29493
rect -218 29459 -212 29493
rect -258 29421 -212 29459
rect -258 29387 -252 29421
rect -218 29387 -212 29421
rect -258 29349 -212 29387
rect -258 29315 -252 29349
rect -218 29315 -212 29349
rect -258 29277 -212 29315
rect -258 29243 -252 29277
rect -218 29243 -212 29277
rect -258 29205 -212 29243
rect -258 29171 -252 29205
rect -218 29171 -212 29205
rect -258 29133 -212 29171
rect -258 29099 -252 29133
rect -218 29099 -212 29133
rect -258 29061 -212 29099
rect -258 29027 -252 29061
rect -218 29027 -212 29061
rect -258 28989 -212 29027
rect -258 28955 -252 28989
rect -218 28955 -212 28989
rect -258 28917 -212 28955
rect -258 28883 -252 28917
rect -218 28883 -212 28917
rect -258 28845 -212 28883
rect -258 28811 -252 28845
rect -218 28811 -212 28845
rect -258 28773 -212 28811
rect -258 28739 -252 28773
rect -218 28739 -212 28773
rect -258 28701 -212 28739
rect -258 28667 -252 28701
rect -218 28667 -212 28701
rect -258 28629 -212 28667
rect -258 28595 -252 28629
rect -218 28595 -212 28629
rect -258 28557 -212 28595
rect -258 28523 -252 28557
rect -218 28523 -212 28557
rect -258 28485 -212 28523
rect -258 28451 -252 28485
rect -218 28451 -212 28485
rect -258 28413 -212 28451
rect -258 28379 -252 28413
rect -218 28379 -212 28413
rect -258 28341 -212 28379
rect -258 28307 -252 28341
rect -218 28307 -212 28341
rect -258 28269 -212 28307
rect -258 28235 -252 28269
rect -218 28235 -212 28269
rect -258 28197 -212 28235
rect -258 28163 -252 28197
rect -218 28163 -212 28197
rect -258 28125 -212 28163
rect -258 28091 -252 28125
rect -218 28091 -212 28125
rect -258 28053 -212 28091
rect -258 28019 -252 28053
rect -218 28019 -212 28053
rect -258 27981 -212 28019
rect -258 27947 -252 27981
rect -218 27947 -212 27981
rect -258 27909 -212 27947
rect -258 27875 -252 27909
rect -218 27875 -212 27909
rect -258 27837 -212 27875
rect -258 27803 -252 27837
rect -218 27803 -212 27837
rect -258 27765 -212 27803
rect -258 27731 -252 27765
rect -218 27731 -212 27765
rect -258 27693 -212 27731
rect -258 27659 -252 27693
rect -218 27659 -212 27693
rect -258 27621 -212 27659
rect -258 27587 -252 27621
rect -218 27587 -212 27621
rect -258 27549 -212 27587
rect -258 27515 -252 27549
rect -218 27515 -212 27549
rect -258 27477 -212 27515
rect -258 27443 -252 27477
rect -218 27443 -212 27477
rect -258 27405 -212 27443
rect -258 27371 -252 27405
rect -218 27371 -212 27405
rect -258 27333 -212 27371
rect -258 27299 -252 27333
rect -218 27299 -212 27333
rect -258 27261 -212 27299
rect -258 27227 -252 27261
rect -218 27227 -212 27261
rect -258 27189 -212 27227
rect -258 27155 -252 27189
rect -218 27155 -212 27189
rect -258 27117 -212 27155
rect -258 27083 -252 27117
rect -218 27083 -212 27117
rect -258 27045 -212 27083
rect -258 27011 -252 27045
rect -218 27011 -212 27045
rect -258 26973 -212 27011
rect -258 26939 -252 26973
rect -218 26939 -212 26973
rect -258 26901 -212 26939
rect -258 26867 -252 26901
rect -218 26867 -212 26901
rect -258 26829 -212 26867
rect -258 26795 -252 26829
rect -218 26795 -212 26829
rect -258 26757 -212 26795
rect -258 26723 -252 26757
rect -218 26723 -212 26757
rect -258 26685 -212 26723
rect -258 26651 -252 26685
rect -218 26651 -212 26685
rect -258 26613 -212 26651
rect -258 26579 -252 26613
rect -218 26579 -212 26613
rect -258 26541 -212 26579
rect -258 26507 -252 26541
rect -218 26507 -212 26541
rect -258 26469 -212 26507
rect -258 26435 -252 26469
rect -218 26435 -212 26469
rect -258 26397 -212 26435
rect -258 26363 -252 26397
rect -218 26363 -212 26397
rect -258 26325 -212 26363
rect -258 26291 -252 26325
rect -218 26291 -212 26325
rect -258 26253 -212 26291
rect -258 26219 -252 26253
rect -218 26219 -212 26253
rect -258 26181 -212 26219
rect -258 26147 -252 26181
rect -218 26147 -212 26181
rect -258 26109 -212 26147
rect -258 26075 -252 26109
rect -218 26075 -212 26109
rect -258 26037 -212 26075
rect -258 26003 -252 26037
rect -218 26003 -212 26037
rect -258 25965 -212 26003
rect -258 25931 -252 25965
rect -218 25931 -212 25965
rect -258 25893 -212 25931
rect -258 25859 -252 25893
rect -218 25859 -212 25893
rect -258 25821 -212 25859
rect -258 25787 -252 25821
rect -218 25787 -212 25821
rect -258 25749 -212 25787
rect -258 25715 -252 25749
rect -218 25715 -212 25749
rect -258 25677 -212 25715
rect -258 25643 -252 25677
rect -218 25643 -212 25677
rect -258 25605 -212 25643
rect -258 25571 -252 25605
rect -218 25571 -212 25605
rect -258 25533 -212 25571
rect -258 25499 -252 25533
rect -218 25499 -212 25533
rect -258 25461 -212 25499
rect -258 25427 -252 25461
rect -218 25427 -212 25461
rect -258 25389 -212 25427
rect -258 25355 -252 25389
rect -218 25355 -212 25389
rect -258 25317 -212 25355
rect -258 25283 -252 25317
rect -218 25283 -212 25317
rect -258 25245 -212 25283
rect -258 25211 -252 25245
rect -218 25211 -212 25245
rect -258 25173 -212 25211
rect -258 25139 -252 25173
rect -218 25139 -212 25173
rect -258 25101 -212 25139
rect -258 25067 -252 25101
rect -218 25067 -212 25101
rect -258 25029 -212 25067
rect -258 24995 -252 25029
rect -218 24995 -212 25029
rect -258 24957 -212 24995
rect -258 24923 -252 24957
rect -218 24923 -212 24957
rect -258 24885 -212 24923
rect -258 24851 -252 24885
rect -218 24851 -212 24885
rect -258 24813 -212 24851
rect -258 24779 -252 24813
rect -218 24779 -212 24813
rect -258 24741 -212 24779
rect -258 24707 -252 24741
rect -218 24707 -212 24741
rect -258 24669 -212 24707
rect -258 24635 -252 24669
rect -218 24635 -212 24669
rect -258 24597 -212 24635
rect -258 24563 -252 24597
rect -218 24563 -212 24597
rect -258 24525 -212 24563
rect -258 24491 -252 24525
rect -218 24491 -212 24525
rect -258 24453 -212 24491
rect -258 24419 -252 24453
rect -218 24419 -212 24453
rect -258 24381 -212 24419
rect -258 24347 -252 24381
rect -218 24347 -212 24381
rect -258 24309 -212 24347
rect -258 24275 -252 24309
rect -218 24275 -212 24309
rect -258 24237 -212 24275
rect -258 24203 -252 24237
rect -218 24203 -212 24237
rect -258 24165 -212 24203
rect -258 24131 -252 24165
rect -218 24131 -212 24165
rect -258 24093 -212 24131
rect -258 24059 -252 24093
rect -218 24059 -212 24093
rect -258 24021 -212 24059
rect -258 23987 -252 24021
rect -218 23987 -212 24021
rect -258 23949 -212 23987
rect -258 23915 -252 23949
rect -218 23915 -212 23949
rect -258 23877 -212 23915
rect -258 23843 -252 23877
rect -218 23843 -212 23877
rect -258 23805 -212 23843
rect -258 23771 -252 23805
rect -218 23771 -212 23805
rect -258 23733 -212 23771
rect -258 23699 -252 23733
rect -218 23699 -212 23733
rect -258 23661 -212 23699
rect -258 23627 -252 23661
rect -218 23627 -212 23661
rect -258 23589 -212 23627
rect -258 23555 -252 23589
rect -218 23555 -212 23589
rect -258 23517 -212 23555
rect -258 23483 -252 23517
rect -218 23483 -212 23517
rect -258 23445 -212 23483
rect -258 23411 -252 23445
rect -218 23411 -212 23445
rect -258 23373 -212 23411
rect -258 23339 -252 23373
rect -218 23339 -212 23373
rect -258 23301 -212 23339
rect -258 23267 -252 23301
rect -218 23267 -212 23301
rect -258 23229 -212 23267
rect -258 23195 -252 23229
rect -218 23195 -212 23229
rect -258 23157 -212 23195
rect -258 23123 -252 23157
rect -218 23123 -212 23157
rect -258 23085 -212 23123
rect -258 23051 -252 23085
rect -218 23051 -212 23085
rect -258 23013 -212 23051
rect -258 22979 -252 23013
rect -218 22979 -212 23013
rect -258 22941 -212 22979
rect -258 22907 -252 22941
rect -218 22907 -212 22941
rect -258 22869 -212 22907
rect -258 22835 -252 22869
rect -218 22835 -212 22869
rect -258 22797 -212 22835
rect -258 22763 -252 22797
rect -218 22763 -212 22797
rect -258 22725 -212 22763
rect -258 22691 -252 22725
rect -218 22691 -212 22725
rect -258 22653 -212 22691
rect -258 22619 -252 22653
rect -218 22619 -212 22653
rect -258 22581 -212 22619
rect -258 22547 -252 22581
rect -218 22547 -212 22581
rect -258 22509 -212 22547
rect -258 22475 -252 22509
rect -218 22475 -212 22509
rect -258 22437 -212 22475
rect -258 22403 -252 22437
rect -218 22403 -212 22437
rect -258 22365 -212 22403
rect -258 22331 -252 22365
rect -218 22331 -212 22365
rect -258 22293 -212 22331
rect -258 22259 -252 22293
rect -218 22259 -212 22293
rect -258 22221 -212 22259
rect -258 22187 -252 22221
rect -218 22187 -212 22221
rect -258 22149 -212 22187
rect -258 22115 -252 22149
rect -218 22115 -212 22149
rect -258 22077 -212 22115
rect -258 22043 -252 22077
rect -218 22043 -212 22077
rect -258 22005 -212 22043
rect -258 21971 -252 22005
rect -218 21971 -212 22005
rect -258 21933 -212 21971
rect -258 21899 -252 21933
rect -218 21899 -212 21933
rect -258 21861 -212 21899
rect -258 21827 -252 21861
rect -218 21827 -212 21861
rect -258 21789 -212 21827
rect -258 21755 -252 21789
rect -218 21755 -212 21789
rect -258 21717 -212 21755
rect -258 21683 -252 21717
rect -218 21683 -212 21717
rect -258 21645 -212 21683
rect -258 21611 -252 21645
rect -218 21611 -212 21645
rect -258 21573 -212 21611
rect -258 21539 -252 21573
rect -218 21539 -212 21573
rect -258 21501 -212 21539
rect -258 21467 -252 21501
rect -218 21467 -212 21501
rect -258 21429 -212 21467
rect -258 21395 -252 21429
rect -218 21395 -212 21429
rect -258 21357 -212 21395
rect -258 21323 -252 21357
rect -218 21323 -212 21357
rect -258 21285 -212 21323
rect -258 21251 -252 21285
rect -218 21251 -212 21285
rect -258 21213 -212 21251
rect -258 21179 -252 21213
rect -218 21179 -212 21213
rect -258 21141 -212 21179
rect -258 21107 -252 21141
rect -218 21107 -212 21141
rect -258 21069 -212 21107
rect -258 21035 -252 21069
rect -218 21035 -212 21069
rect -258 20997 -212 21035
rect -258 20963 -252 20997
rect -218 20963 -212 20997
rect -258 20925 -212 20963
rect -258 20891 -252 20925
rect -218 20891 -212 20925
rect -258 20853 -212 20891
rect -258 20819 -252 20853
rect -218 20819 -212 20853
rect -258 20781 -212 20819
rect -258 20747 -252 20781
rect -218 20747 -212 20781
rect -258 20709 -212 20747
rect -258 20675 -252 20709
rect -218 20675 -212 20709
rect -258 20637 -212 20675
rect -258 20603 -252 20637
rect -218 20603 -212 20637
rect -258 20565 -212 20603
rect -258 20531 -252 20565
rect -218 20531 -212 20565
rect -258 20493 -212 20531
rect -258 20459 -252 20493
rect -218 20459 -212 20493
rect -258 20421 -212 20459
rect -258 20387 -252 20421
rect -218 20387 -212 20421
rect -258 20349 -212 20387
rect -258 20315 -252 20349
rect -218 20315 -212 20349
rect -258 20277 -212 20315
rect -258 20243 -252 20277
rect -218 20243 -212 20277
rect -258 20205 -212 20243
rect -258 20171 -252 20205
rect -218 20171 -212 20205
rect -258 20133 -212 20171
rect -258 20099 -252 20133
rect -218 20099 -212 20133
rect -258 20061 -212 20099
rect -258 20027 -252 20061
rect -218 20027 -212 20061
rect -258 19989 -212 20027
rect -258 19955 -252 19989
rect -218 19955 -212 19989
rect -258 19917 -212 19955
rect -258 19883 -252 19917
rect -218 19883 -212 19917
rect -258 19845 -212 19883
rect -258 19811 -252 19845
rect -218 19811 -212 19845
rect -258 19773 -212 19811
rect -258 19739 -252 19773
rect -218 19739 -212 19773
rect -258 19701 -212 19739
rect -258 19667 -252 19701
rect -218 19667 -212 19701
rect -258 19629 -212 19667
rect -258 19595 -252 19629
rect -218 19595 -212 19629
rect -258 19557 -212 19595
rect -258 19523 -252 19557
rect -218 19523 -212 19557
rect -258 19485 -212 19523
rect -258 19451 -252 19485
rect -218 19451 -212 19485
rect -258 19413 -212 19451
rect -258 19379 -252 19413
rect -218 19379 -212 19413
rect -258 19341 -212 19379
rect -258 19307 -252 19341
rect -218 19307 -212 19341
rect -258 19269 -212 19307
rect -258 19235 -252 19269
rect -218 19235 -212 19269
rect -258 19197 -212 19235
rect -258 19163 -252 19197
rect -218 19163 -212 19197
rect -258 19125 -212 19163
rect -258 19091 -252 19125
rect -218 19091 -212 19125
rect -258 19053 -212 19091
rect -258 19019 -252 19053
rect -218 19019 -212 19053
rect -258 18981 -212 19019
rect -258 18947 -252 18981
rect -218 18947 -212 18981
rect -258 18909 -212 18947
rect -258 18875 -252 18909
rect -218 18875 -212 18909
rect -258 18837 -212 18875
rect -258 18803 -252 18837
rect -218 18803 -212 18837
rect -258 18765 -212 18803
rect -258 18731 -252 18765
rect -218 18731 -212 18765
rect -258 18693 -212 18731
rect -258 18659 -252 18693
rect -218 18659 -212 18693
rect -258 18621 -212 18659
rect -258 18587 -252 18621
rect -218 18587 -212 18621
rect -258 18549 -212 18587
rect -258 18515 -252 18549
rect -218 18515 -212 18549
rect -258 18477 -212 18515
rect -258 18443 -252 18477
rect -218 18443 -212 18477
rect -258 18405 -212 18443
rect -258 18371 -252 18405
rect -218 18371 -212 18405
rect -258 18333 -212 18371
rect -258 18299 -252 18333
rect -218 18299 -212 18333
rect -258 18261 -212 18299
rect -258 18227 -252 18261
rect -218 18227 -212 18261
rect -258 18189 -212 18227
rect -258 18155 -252 18189
rect -218 18155 -212 18189
rect -258 18117 -212 18155
rect -258 18083 -252 18117
rect -218 18083 -212 18117
rect -258 18045 -212 18083
rect -258 18011 -252 18045
rect -218 18011 -212 18045
rect -258 17973 -212 18011
rect -258 17939 -252 17973
rect -218 17939 -212 17973
rect -258 17901 -212 17939
rect -258 17867 -252 17901
rect -218 17867 -212 17901
rect -258 17829 -212 17867
rect -258 17795 -252 17829
rect -218 17795 -212 17829
rect -258 17757 -212 17795
rect -258 17723 -252 17757
rect -218 17723 -212 17757
rect -258 17685 -212 17723
rect -258 17651 -252 17685
rect -218 17651 -212 17685
rect -258 17613 -212 17651
rect -258 17579 -252 17613
rect -218 17579 -212 17613
rect -258 17541 -212 17579
rect -258 17507 -252 17541
rect -218 17507 -212 17541
rect -258 17469 -212 17507
rect -258 17435 -252 17469
rect -218 17435 -212 17469
rect -258 17397 -212 17435
rect -258 17363 -252 17397
rect -218 17363 -212 17397
rect -258 17325 -212 17363
rect -258 17291 -252 17325
rect -218 17291 -212 17325
rect -258 17253 -212 17291
rect -258 17219 -252 17253
rect -218 17219 -212 17253
rect -258 17181 -212 17219
rect -258 17147 -252 17181
rect -218 17147 -212 17181
rect -258 17109 -212 17147
rect -258 17075 -252 17109
rect -218 17075 -212 17109
rect -258 17037 -212 17075
rect -258 17003 -252 17037
rect -218 17003 -212 17037
rect -258 16965 -212 17003
rect -258 16931 -252 16965
rect -218 16931 -212 16965
rect -258 16893 -212 16931
rect -258 16859 -252 16893
rect -218 16859 -212 16893
rect -258 16821 -212 16859
rect -258 16787 -252 16821
rect -218 16787 -212 16821
rect -258 16749 -212 16787
rect -258 16715 -252 16749
rect -218 16715 -212 16749
rect -258 16677 -212 16715
rect -258 16643 -252 16677
rect -218 16643 -212 16677
rect -258 16605 -212 16643
rect -258 16571 -252 16605
rect -218 16571 -212 16605
rect -258 16533 -212 16571
rect -258 16499 -252 16533
rect -218 16499 -212 16533
rect -258 16461 -212 16499
rect -258 16427 -252 16461
rect -218 16427 -212 16461
rect -258 16389 -212 16427
rect -258 16355 -252 16389
rect -218 16355 -212 16389
rect -258 16317 -212 16355
rect -258 16283 -252 16317
rect -218 16283 -212 16317
rect -258 16245 -212 16283
rect -258 16211 -252 16245
rect -218 16211 -212 16245
rect -258 16173 -212 16211
rect -258 16139 -252 16173
rect -218 16139 -212 16173
rect -258 16101 -212 16139
rect -258 16067 -252 16101
rect -218 16067 -212 16101
rect -258 16029 -212 16067
rect -258 15995 -252 16029
rect -218 15995 -212 16029
rect -258 15957 -212 15995
rect -258 15923 -252 15957
rect -218 15923 -212 15957
rect -258 15885 -212 15923
rect -258 15851 -252 15885
rect -218 15851 -212 15885
rect -258 15813 -212 15851
rect -258 15779 -252 15813
rect -218 15779 -212 15813
rect -258 15741 -212 15779
rect -258 15707 -252 15741
rect -218 15707 -212 15741
rect -258 15669 -212 15707
rect -258 15635 -252 15669
rect -218 15635 -212 15669
rect -258 15597 -212 15635
rect -258 15563 -252 15597
rect -218 15563 -212 15597
rect -258 15525 -212 15563
rect -258 15491 -252 15525
rect -218 15491 -212 15525
rect -258 15453 -212 15491
rect -258 15419 -252 15453
rect -218 15419 -212 15453
rect -258 15381 -212 15419
rect -258 15347 -252 15381
rect -218 15347 -212 15381
rect -258 15309 -212 15347
rect -258 15275 -252 15309
rect -218 15275 -212 15309
rect -258 15237 -212 15275
rect -258 15203 -252 15237
rect -218 15203 -212 15237
rect -258 15165 -212 15203
rect -258 15131 -252 15165
rect -218 15131 -212 15165
rect -258 15093 -212 15131
rect -258 15059 -252 15093
rect -218 15059 -212 15093
rect -258 15021 -212 15059
rect -258 14987 -252 15021
rect -218 14987 -212 15021
rect -258 14949 -212 14987
rect -258 14915 -252 14949
rect -218 14915 -212 14949
rect -258 14877 -212 14915
rect -258 14843 -252 14877
rect -218 14843 -212 14877
rect -258 14805 -212 14843
rect -258 14771 -252 14805
rect -218 14771 -212 14805
rect -258 14733 -212 14771
rect -258 14699 -252 14733
rect -218 14699 -212 14733
rect -258 14661 -212 14699
rect -258 14627 -252 14661
rect -218 14627 -212 14661
rect -258 14589 -212 14627
rect -258 14555 -252 14589
rect -218 14555 -212 14589
rect -258 14517 -212 14555
rect -258 14483 -252 14517
rect -218 14483 -212 14517
rect -258 14445 -212 14483
rect -258 14411 -252 14445
rect -218 14411 -212 14445
rect -258 14373 -212 14411
rect -258 14339 -252 14373
rect -218 14339 -212 14373
rect -258 14301 -212 14339
rect -258 14267 -252 14301
rect -218 14267 -212 14301
rect -258 14229 -212 14267
rect -258 14195 -252 14229
rect -218 14195 -212 14229
rect -258 14157 -212 14195
rect -258 14123 -252 14157
rect -218 14123 -212 14157
rect -258 14085 -212 14123
rect -258 14051 -252 14085
rect -218 14051 -212 14085
rect -258 14013 -212 14051
rect -258 13979 -252 14013
rect -218 13979 -212 14013
rect -258 13941 -212 13979
rect -258 13907 -252 13941
rect -218 13907 -212 13941
rect -258 13869 -212 13907
rect -258 13835 -252 13869
rect -218 13835 -212 13869
rect -258 13797 -212 13835
rect -258 13763 -252 13797
rect -218 13763 -212 13797
rect -258 13725 -212 13763
rect -258 13691 -252 13725
rect -218 13691 -212 13725
rect -258 13653 -212 13691
rect -258 13619 -252 13653
rect -218 13619 -212 13653
rect -258 13581 -212 13619
rect -258 13547 -252 13581
rect -218 13547 -212 13581
rect -258 13509 -212 13547
rect -258 13475 -252 13509
rect -218 13475 -212 13509
rect -258 13437 -212 13475
rect -258 13403 -252 13437
rect -218 13403 -212 13437
rect -258 13365 -212 13403
rect -258 13331 -252 13365
rect -218 13331 -212 13365
rect -258 13293 -212 13331
rect -258 13259 -252 13293
rect -218 13259 -212 13293
rect -258 13221 -212 13259
rect -258 13187 -252 13221
rect -218 13187 -212 13221
rect -258 13149 -212 13187
rect -258 13115 -252 13149
rect -218 13115 -212 13149
rect -258 13077 -212 13115
rect -258 13043 -252 13077
rect -218 13043 -212 13077
rect -258 13005 -212 13043
rect -258 12971 -252 13005
rect -218 12971 -212 13005
rect -258 12933 -212 12971
rect -258 12899 -252 12933
rect -218 12899 -212 12933
rect -258 12861 -212 12899
rect -258 12827 -252 12861
rect -218 12827 -212 12861
rect -258 12789 -212 12827
rect -258 12755 -252 12789
rect -218 12755 -212 12789
rect -258 12717 -212 12755
rect -258 12683 -252 12717
rect -218 12683 -212 12717
rect -258 12645 -212 12683
rect -258 12611 -252 12645
rect -218 12611 -212 12645
rect -258 12573 -212 12611
rect -258 12539 -252 12573
rect -218 12539 -212 12573
rect -258 12501 -212 12539
rect -258 12467 -252 12501
rect -218 12467 -212 12501
rect -258 12429 -212 12467
rect -258 12395 -252 12429
rect -218 12395 -212 12429
rect -258 12357 -212 12395
rect -258 12323 -252 12357
rect -218 12323 -212 12357
rect -258 12285 -212 12323
rect -258 12251 -252 12285
rect -218 12251 -212 12285
rect -258 12213 -212 12251
rect -258 12179 -252 12213
rect -218 12179 -212 12213
rect -258 12141 -212 12179
rect -258 12107 -252 12141
rect -218 12107 -212 12141
rect -258 12069 -212 12107
rect -258 12035 -252 12069
rect -218 12035 -212 12069
rect -258 11997 -212 12035
rect -258 11963 -252 11997
rect -218 11963 -212 11997
rect -258 11925 -212 11963
rect -258 11891 -252 11925
rect -218 11891 -212 11925
rect -258 11853 -212 11891
rect -258 11819 -252 11853
rect -218 11819 -212 11853
rect -258 11781 -212 11819
rect -258 11747 -252 11781
rect -218 11747 -212 11781
rect -258 11709 -212 11747
rect -258 11675 -252 11709
rect -218 11675 -212 11709
rect -258 11637 -212 11675
rect -258 11603 -252 11637
rect -218 11603 -212 11637
rect -258 11565 -212 11603
rect -258 11531 -252 11565
rect -218 11531 -212 11565
rect -258 11493 -212 11531
rect -258 11459 -252 11493
rect -218 11459 -212 11493
rect -258 11421 -212 11459
rect -258 11387 -252 11421
rect -218 11387 -212 11421
rect -258 11349 -212 11387
rect -258 11315 -252 11349
rect -218 11315 -212 11349
rect -258 11277 -212 11315
rect -258 11243 -252 11277
rect -218 11243 -212 11277
rect -258 11205 -212 11243
rect -258 11171 -252 11205
rect -218 11171 -212 11205
rect -258 11133 -212 11171
rect -258 11099 -252 11133
rect -218 11099 -212 11133
rect -258 11061 -212 11099
rect -258 11027 -252 11061
rect -218 11027 -212 11061
rect -258 10989 -212 11027
rect -258 10955 -252 10989
rect -218 10955 -212 10989
rect -258 10917 -212 10955
rect -258 10883 -252 10917
rect -218 10883 -212 10917
rect -258 10845 -212 10883
rect -258 10811 -252 10845
rect -218 10811 -212 10845
rect -258 10773 -212 10811
rect -258 10739 -252 10773
rect -218 10739 -212 10773
rect -258 10701 -212 10739
rect -258 10667 -252 10701
rect -218 10667 -212 10701
rect -258 10629 -212 10667
rect -258 10595 -252 10629
rect -218 10595 -212 10629
rect -258 10557 -212 10595
rect -258 10523 -252 10557
rect -218 10523 -212 10557
rect -258 10485 -212 10523
rect -258 10451 -252 10485
rect -218 10451 -212 10485
rect -258 10413 -212 10451
rect -258 10379 -252 10413
rect -218 10379 -212 10413
rect -258 10341 -212 10379
rect -258 10307 -252 10341
rect -218 10307 -212 10341
rect -258 10269 -212 10307
rect -258 10235 -252 10269
rect -218 10235 -212 10269
rect -258 10197 -212 10235
rect -258 10163 -252 10197
rect -218 10163 -212 10197
rect -258 10125 -212 10163
rect -258 10091 -252 10125
rect -218 10091 -212 10125
rect -258 10053 -212 10091
rect -258 10019 -252 10053
rect -218 10019 -212 10053
rect -258 9981 -212 10019
rect -258 9947 -252 9981
rect -218 9947 -212 9981
rect -258 9909 -212 9947
rect -258 9875 -252 9909
rect -218 9875 -212 9909
rect -258 9837 -212 9875
rect -258 9803 -252 9837
rect -218 9803 -212 9837
rect -258 9765 -212 9803
rect -258 9731 -252 9765
rect -218 9731 -212 9765
rect -258 9693 -212 9731
rect -258 9659 -252 9693
rect -218 9659 -212 9693
rect -258 9621 -212 9659
rect -258 9587 -252 9621
rect -218 9587 -212 9621
rect -258 9549 -212 9587
rect -258 9515 -252 9549
rect -218 9515 -212 9549
rect -258 9477 -212 9515
rect -258 9443 -252 9477
rect -218 9443 -212 9477
rect -258 9405 -212 9443
rect -258 9371 -252 9405
rect -218 9371 -212 9405
rect -258 9333 -212 9371
rect -258 9299 -252 9333
rect -218 9299 -212 9333
rect -258 9261 -212 9299
rect -258 9227 -252 9261
rect -218 9227 -212 9261
rect -258 9189 -212 9227
rect -258 9155 -252 9189
rect -218 9155 -212 9189
rect -258 9117 -212 9155
rect -258 9083 -252 9117
rect -218 9083 -212 9117
rect -258 9045 -212 9083
rect -258 9011 -252 9045
rect -218 9011 -212 9045
rect -258 8973 -212 9011
rect -258 8939 -252 8973
rect -218 8939 -212 8973
rect -258 8901 -212 8939
rect -258 8867 -252 8901
rect -218 8867 -212 8901
rect -258 8829 -212 8867
rect -258 8795 -252 8829
rect -218 8795 -212 8829
rect -258 8757 -212 8795
rect -258 8723 -252 8757
rect -218 8723 -212 8757
rect -258 8685 -212 8723
rect -258 8651 -252 8685
rect -218 8651 -212 8685
rect -258 8613 -212 8651
rect -258 8579 -252 8613
rect -218 8579 -212 8613
rect -258 8541 -212 8579
rect -258 8507 -252 8541
rect -218 8507 -212 8541
rect -258 8469 -212 8507
rect -258 8435 -252 8469
rect -218 8435 -212 8469
rect -258 8397 -212 8435
rect -258 8363 -252 8397
rect -218 8363 -212 8397
rect -258 8325 -212 8363
rect -258 8291 -252 8325
rect -218 8291 -212 8325
rect -258 8253 -212 8291
rect -258 8219 -252 8253
rect -218 8219 -212 8253
rect -258 8181 -212 8219
rect -258 8147 -252 8181
rect -218 8147 -212 8181
rect -258 8109 -212 8147
rect -258 8075 -252 8109
rect -218 8075 -212 8109
rect -258 8037 -212 8075
rect -258 8003 -252 8037
rect -218 8003 -212 8037
rect -258 7965 -212 8003
rect -258 7931 -252 7965
rect -218 7931 -212 7965
rect -258 7893 -212 7931
rect -258 7859 -252 7893
rect -218 7859 -212 7893
rect -258 7821 -212 7859
rect -258 7787 -252 7821
rect -218 7787 -212 7821
rect -258 7749 -212 7787
rect -258 7715 -252 7749
rect -218 7715 -212 7749
rect -258 7677 -212 7715
rect -258 7643 -252 7677
rect -218 7643 -212 7677
rect -258 7605 -212 7643
rect -258 7571 -252 7605
rect -218 7571 -212 7605
rect -258 7533 -212 7571
rect -258 7499 -252 7533
rect -218 7499 -212 7533
rect -258 7461 -212 7499
rect -258 7427 -252 7461
rect -218 7427 -212 7461
rect -258 7389 -212 7427
rect -258 7355 -252 7389
rect -218 7355 -212 7389
rect -258 7317 -212 7355
rect -258 7283 -252 7317
rect -218 7283 -212 7317
rect -258 7245 -212 7283
rect -258 7211 -252 7245
rect -218 7211 -212 7245
rect -258 7173 -212 7211
rect -258 7139 -252 7173
rect -218 7139 -212 7173
rect -258 7101 -212 7139
rect -258 7067 -252 7101
rect -218 7067 -212 7101
rect -258 7029 -212 7067
rect -258 6995 -252 7029
rect -218 6995 -212 7029
rect -258 6957 -212 6995
rect -258 6923 -252 6957
rect -218 6923 -212 6957
rect -258 6885 -212 6923
rect -258 6851 -252 6885
rect -218 6851 -212 6885
rect -258 6813 -212 6851
rect -258 6779 -252 6813
rect -218 6779 -212 6813
rect -258 6741 -212 6779
rect -258 6707 -252 6741
rect -218 6707 -212 6741
rect -258 6669 -212 6707
rect -258 6635 -252 6669
rect -218 6635 -212 6669
rect -258 6597 -212 6635
rect -258 6563 -252 6597
rect -218 6563 -212 6597
rect -258 6525 -212 6563
rect -258 6491 -252 6525
rect -218 6491 -212 6525
rect -258 6453 -212 6491
rect -258 6419 -252 6453
rect -218 6419 -212 6453
rect -258 6381 -212 6419
rect -258 6347 -252 6381
rect -218 6347 -212 6381
rect -258 6309 -212 6347
rect -258 6275 -252 6309
rect -218 6275 -212 6309
rect -258 6237 -212 6275
rect -258 6203 -252 6237
rect -218 6203 -212 6237
rect -258 6165 -212 6203
rect -258 6131 -252 6165
rect -218 6131 -212 6165
rect -258 6093 -212 6131
rect -258 6059 -252 6093
rect -218 6059 -212 6093
rect -258 6021 -212 6059
rect -258 5987 -252 6021
rect -218 5987 -212 6021
rect -258 5949 -212 5987
rect -258 5915 -252 5949
rect -218 5915 -212 5949
rect -258 5877 -212 5915
rect -258 5843 -252 5877
rect -218 5843 -212 5877
rect -258 5805 -212 5843
rect -258 5771 -252 5805
rect -218 5771 -212 5805
rect -258 5733 -212 5771
rect -258 5699 -252 5733
rect -218 5699 -212 5733
rect -258 5661 -212 5699
rect -258 5627 -252 5661
rect -218 5627 -212 5661
rect -258 5589 -212 5627
rect -258 5555 -252 5589
rect -218 5555 -212 5589
rect -258 5517 -212 5555
rect -258 5483 -252 5517
rect -218 5483 -212 5517
rect -258 5445 -212 5483
rect -258 5411 -252 5445
rect -218 5411 -212 5445
rect -258 5373 -212 5411
rect -258 5339 -252 5373
rect -218 5339 -212 5373
rect -258 5301 -212 5339
rect -258 5267 -252 5301
rect -218 5267 -212 5301
rect -258 5229 -212 5267
rect -258 5195 -252 5229
rect -218 5195 -212 5229
rect -258 5157 -212 5195
rect -258 5123 -252 5157
rect -218 5123 -212 5157
rect -258 5085 -212 5123
rect -258 5051 -252 5085
rect -218 5051 -212 5085
rect -258 5013 -212 5051
rect -258 4979 -252 5013
rect -218 4979 -212 5013
rect -258 4941 -212 4979
rect -258 4907 -252 4941
rect -218 4907 -212 4941
rect -258 4869 -212 4907
rect -258 4835 -252 4869
rect -218 4835 -212 4869
rect -258 4797 -212 4835
rect -258 4763 -252 4797
rect -218 4763 -212 4797
rect -258 4725 -212 4763
rect -258 4691 -252 4725
rect -218 4691 -212 4725
rect -258 4653 -212 4691
rect -258 4619 -252 4653
rect -218 4619 -212 4653
rect 1824 38651 1830 38685
rect 1864 38651 1870 38685
tri 1870 38683 1872 38685 nw
tri 3964 38683 3966 38685 ne
rect 1824 38612 1870 38651
rect 1824 38578 1830 38612
rect 1864 38578 1870 38612
rect 1824 38539 1870 38578
rect 1824 38505 1830 38539
rect 1864 38505 1870 38539
rect 1824 38466 1870 38505
rect 1824 38432 1830 38466
rect 1864 38432 1870 38466
rect 1824 38393 1870 38432
rect 1824 38359 1830 38393
rect 1864 38359 1870 38393
rect 1824 38320 1870 38359
rect 1824 38286 1830 38320
rect 1864 38286 1870 38320
rect 1824 38247 1870 38286
rect 1824 38213 1830 38247
rect 1864 38213 1870 38247
rect 1824 38174 1870 38213
rect 1824 38140 1830 38174
rect 1864 38140 1870 38174
rect 1824 38101 1870 38140
rect 1824 38067 1830 38101
rect 1864 38067 1870 38101
rect 1824 38028 1870 38067
rect 1824 37994 1830 38028
rect 1864 37994 1870 38028
rect 1824 37955 1870 37994
rect 1824 37921 1830 37955
rect 1864 37921 1870 37955
rect 1824 37882 1870 37921
rect 1824 37848 1830 37882
rect 1864 37848 1870 37882
rect 1824 37809 1870 37848
rect 1824 37775 1830 37809
rect 1864 37775 1870 37809
rect 1824 37736 1870 37775
rect 1824 37702 1830 37736
rect 1864 37702 1870 37736
rect 1824 37663 1870 37702
rect 1824 37629 1830 37663
rect 1864 37629 1870 37663
rect 1824 37590 1870 37629
rect 1824 37556 1830 37590
rect 1864 37556 1870 37590
rect 1824 37517 1870 37556
rect 1824 37483 1830 37517
rect 1864 37483 1870 37517
rect 1824 37444 1870 37483
rect 1824 37410 1830 37444
rect 1864 37410 1870 37444
rect 1824 37371 1870 37410
rect 1824 37337 1830 37371
rect 1864 37337 1870 37371
rect 1824 37298 1870 37337
rect 1824 37264 1830 37298
rect 1864 37264 1870 37298
rect 1824 37225 1870 37264
rect 1824 37191 1830 37225
rect 1864 37191 1870 37225
rect 1824 37152 1870 37191
rect 1824 37118 1830 37152
rect 1864 37118 1870 37152
rect 1824 37079 1870 37118
rect 1824 37045 1830 37079
rect 1864 37045 1870 37079
rect 1824 37006 1870 37045
rect 1824 36972 1830 37006
rect 1864 36972 1870 37006
rect 1824 36933 1870 36972
rect 1824 36899 1830 36933
rect 1864 36899 1870 36933
rect 1824 36860 1870 36899
rect 1824 36826 1830 36860
rect 1864 36826 1870 36860
rect 1824 36787 1870 36826
rect 1824 36753 1830 36787
rect 1864 36753 1870 36787
rect 1824 36714 1870 36753
rect 1824 36680 1830 36714
rect 1864 36680 1870 36714
rect 1824 36641 1870 36680
rect 1824 36607 1830 36641
rect 1864 36607 1870 36641
rect 1824 36568 1870 36607
rect 1824 36534 1830 36568
rect 1864 36534 1870 36568
rect 1824 36495 1870 36534
rect 1824 36461 1830 36495
rect 1864 36461 1870 36495
rect 1824 36422 1870 36461
rect 1824 36388 1830 36422
rect 1864 36388 1870 36422
rect 1824 36349 1870 36388
rect 1824 36315 1830 36349
rect 1864 36315 1870 36349
rect 1824 36276 1870 36315
rect 1824 36242 1830 36276
rect 1864 36242 1870 36276
rect 1824 36203 1870 36242
rect 1824 36169 1830 36203
rect 1864 36169 1870 36203
rect 1824 36130 1870 36169
rect 1824 36096 1830 36130
rect 1864 36096 1870 36130
rect 1824 36057 1870 36096
rect 1824 36023 1830 36057
rect 1864 36023 1870 36057
rect 1824 35984 1870 36023
rect 1824 35950 1830 35984
rect 1864 35950 1870 35984
rect 1824 35911 1870 35950
rect 1824 35877 1830 35911
rect 1864 35877 1870 35911
rect 1824 35838 1870 35877
rect 1824 35804 1830 35838
rect 1864 35804 1870 35838
rect 1824 35765 1870 35804
rect 1824 35731 1830 35765
rect 1864 35731 1870 35765
rect 1824 35692 1870 35731
rect 1824 35658 1830 35692
rect 1864 35658 1870 35692
rect 1824 35619 1870 35658
rect 1824 35585 1830 35619
rect 1864 35585 1870 35619
rect 1824 35546 1870 35585
rect 1824 35512 1830 35546
rect 1864 35512 1870 35546
rect 1824 35473 1870 35512
rect 1824 35439 1830 35473
rect 1864 35439 1870 35473
rect 1824 35400 1870 35439
rect 1824 35366 1830 35400
rect 1864 35366 1870 35400
rect 1824 35327 1870 35366
rect 1824 35293 1830 35327
rect 1864 35293 1870 35327
rect 1824 35254 1870 35293
rect 1824 35220 1830 35254
rect 1864 35220 1870 35254
rect 1824 35181 1870 35220
rect 1824 35147 1830 35181
rect 1864 35147 1870 35181
rect 1824 35109 1870 35147
rect 1824 35075 1830 35109
rect 1864 35075 1870 35109
rect 1824 35037 1870 35075
rect 1824 35003 1830 35037
rect 1864 35003 1870 35037
rect 1824 34965 1870 35003
rect 1824 34931 1830 34965
rect 1864 34931 1870 34965
rect 1824 34893 1870 34931
rect 1824 34859 1830 34893
rect 1864 34859 1870 34893
rect 1824 34821 1870 34859
rect 1824 34787 1830 34821
rect 1864 34787 1870 34821
rect 1824 34749 1870 34787
rect 1824 34715 1830 34749
rect 1864 34715 1870 34749
rect 1824 34677 1870 34715
rect 1824 34643 1830 34677
rect 1864 34643 1870 34677
rect 1824 34605 1870 34643
rect 1824 34571 1830 34605
rect 1864 34571 1870 34605
rect 1824 34533 1870 34571
rect 1824 34499 1830 34533
rect 1864 34499 1870 34533
rect 1824 34461 1870 34499
rect 1824 34427 1830 34461
rect 1864 34427 1870 34461
rect 1824 34389 1870 34427
rect 1824 34355 1830 34389
rect 1864 34355 1870 34389
rect 1824 34317 1870 34355
rect 1824 34283 1830 34317
rect 1864 34283 1870 34317
rect 1824 34245 1870 34283
rect 1824 34211 1830 34245
rect 1864 34211 1870 34245
rect 1824 34173 1870 34211
rect 1824 34139 1830 34173
rect 1864 34139 1870 34173
rect 1824 34101 1870 34139
rect 1824 34067 1830 34101
rect 1864 34067 1870 34101
rect 1824 34029 1870 34067
rect 1824 33995 1830 34029
rect 1864 33995 1870 34029
rect 1824 33957 1870 33995
rect 1824 33923 1830 33957
rect 1864 33923 1870 33957
rect 1824 33885 1870 33923
rect 1824 33851 1830 33885
rect 1864 33851 1870 33885
rect 1824 33813 1870 33851
rect 1824 33779 1830 33813
rect 1864 33779 1870 33813
rect 1824 33741 1870 33779
rect 1824 33707 1830 33741
rect 1864 33707 1870 33741
rect 1824 33669 1870 33707
rect 1824 33635 1830 33669
rect 1864 33635 1870 33669
rect 1824 33597 1870 33635
rect 1824 33563 1830 33597
rect 1864 33563 1870 33597
rect 1824 33525 1870 33563
rect 1824 33491 1830 33525
rect 1864 33491 1870 33525
rect 1824 33453 1870 33491
rect 1824 33419 1830 33453
rect 1864 33419 1870 33453
rect 1824 33381 1870 33419
rect 1824 33347 1830 33381
rect 1864 33347 1870 33381
rect 1824 33309 1870 33347
rect 1824 33275 1830 33309
rect 1864 33275 1870 33309
rect 1824 33237 1870 33275
rect 1824 33203 1830 33237
rect 1864 33203 1870 33237
rect 1824 33165 1870 33203
rect 1824 33131 1830 33165
rect 1864 33131 1870 33165
rect 1824 33093 1870 33131
rect 1824 33059 1830 33093
rect 1864 33059 1870 33093
rect 1824 33021 1870 33059
rect 1824 32987 1830 33021
rect 1864 32987 1870 33021
rect 1824 32949 1870 32987
rect 1824 32915 1830 32949
rect 1864 32915 1870 32949
rect 1824 32877 1870 32915
rect 1824 32843 1830 32877
rect 1864 32843 1870 32877
rect 1824 32805 1870 32843
rect 1824 32771 1830 32805
rect 1864 32771 1870 32805
rect 1824 32733 1870 32771
rect 1824 32699 1830 32733
rect 1864 32699 1870 32733
rect 1824 32661 1870 32699
rect 1824 32627 1830 32661
rect 1864 32627 1870 32661
rect 1824 32589 1870 32627
rect 1824 32555 1830 32589
rect 1864 32555 1870 32589
rect 1824 32517 1870 32555
rect 1824 32483 1830 32517
rect 1864 32483 1870 32517
rect 1824 32445 1870 32483
rect 1824 32411 1830 32445
rect 1864 32411 1870 32445
rect 1824 32373 1870 32411
rect 1824 32339 1830 32373
rect 1864 32339 1870 32373
rect 1824 32301 1870 32339
rect 1824 32267 1830 32301
rect 1864 32267 1870 32301
rect 1824 32229 1870 32267
rect 1824 32195 1830 32229
rect 1864 32195 1870 32229
rect 1824 32157 1870 32195
rect 1824 32123 1830 32157
rect 1864 32123 1870 32157
rect 1824 32085 1870 32123
rect 1824 32051 1830 32085
rect 1864 32051 1870 32085
rect 1824 32013 1870 32051
rect 1824 31979 1830 32013
rect 1864 31979 1870 32013
rect 1824 31941 1870 31979
rect 1824 31907 1830 31941
rect 1864 31907 1870 31941
rect 1824 31869 1870 31907
rect 1824 31835 1830 31869
rect 1864 31835 1870 31869
rect 1824 31797 1870 31835
rect 1824 31763 1830 31797
rect 1864 31763 1870 31797
rect 1824 31725 1870 31763
rect 1824 31691 1830 31725
rect 1864 31691 1870 31725
rect 1824 31653 1870 31691
rect 1824 31619 1830 31653
rect 1864 31619 1870 31653
rect 1824 31581 1870 31619
rect 1824 31547 1830 31581
rect 1864 31547 1870 31581
rect 1824 31509 1870 31547
rect 1824 31475 1830 31509
rect 1864 31475 1870 31509
rect 1824 31437 1870 31475
rect 1824 31403 1830 31437
rect 1864 31403 1870 31437
rect 1824 31365 1870 31403
rect 1824 31331 1830 31365
rect 1864 31331 1870 31365
rect 1824 31293 1870 31331
rect 1824 31259 1830 31293
rect 1864 31259 1870 31293
rect 1824 31221 1870 31259
rect 1824 31187 1830 31221
rect 1864 31187 1870 31221
rect 1824 31149 1870 31187
rect 1824 31115 1830 31149
rect 1864 31115 1870 31149
rect 1824 31077 1870 31115
rect 1824 31043 1830 31077
rect 1864 31043 1870 31077
rect 1824 31005 1870 31043
rect 1824 30971 1830 31005
rect 1864 30971 1870 31005
rect 1824 30933 1870 30971
rect 1824 30899 1830 30933
rect 1864 30899 1870 30933
rect 1824 30861 1870 30899
rect 1824 30827 1830 30861
rect 1864 30827 1870 30861
rect 1824 30789 1870 30827
rect 1824 30755 1830 30789
rect 1864 30755 1870 30789
rect 1824 30717 1870 30755
rect 1824 30683 1830 30717
rect 1864 30683 1870 30717
rect 1824 30645 1870 30683
rect 1824 30611 1830 30645
rect 1864 30611 1870 30645
rect 1824 30573 1870 30611
rect 1824 30539 1830 30573
rect 1864 30539 1870 30573
rect 1824 30501 1870 30539
rect 1824 30467 1830 30501
rect 1864 30467 1870 30501
rect 1824 30429 1870 30467
rect 1824 30395 1830 30429
rect 1864 30395 1870 30429
rect 1824 30357 1870 30395
rect 1824 30323 1830 30357
rect 1864 30323 1870 30357
rect 1824 30285 1870 30323
rect 1824 30251 1830 30285
rect 1864 30251 1870 30285
rect 1824 30213 1870 30251
rect 1824 30179 1830 30213
rect 1864 30179 1870 30213
rect 1824 30141 1870 30179
rect 1824 30107 1830 30141
rect 1864 30107 1870 30141
rect 1824 30069 1870 30107
rect 1824 30035 1830 30069
rect 1864 30035 1870 30069
rect 1824 29997 1870 30035
rect 1824 29963 1830 29997
rect 1864 29963 1870 29997
rect 1824 29925 1870 29963
rect 1824 29891 1830 29925
rect 1864 29891 1870 29925
rect 1824 29853 1870 29891
rect 1824 29819 1830 29853
rect 1864 29819 1870 29853
rect 1824 29781 1870 29819
rect 1824 29747 1830 29781
rect 1864 29747 1870 29781
rect 1824 29709 1870 29747
rect 1824 29675 1830 29709
rect 1864 29675 1870 29709
rect 1824 29637 1870 29675
rect 1824 29603 1830 29637
rect 1864 29603 1870 29637
rect 1824 29565 1870 29603
rect 1824 29531 1830 29565
rect 1864 29531 1870 29565
rect 1824 29493 1870 29531
rect 1824 29459 1830 29493
rect 1864 29459 1870 29493
rect 1824 29421 1870 29459
rect 1824 29387 1830 29421
rect 1864 29387 1870 29421
rect 1824 29349 1870 29387
rect 1824 29315 1830 29349
rect 1864 29315 1870 29349
rect 1824 29277 1870 29315
rect 1824 29243 1830 29277
rect 1864 29243 1870 29277
rect 1824 29205 1870 29243
rect 1824 29171 1830 29205
rect 1864 29171 1870 29205
rect 1824 29133 1870 29171
rect 1824 29099 1830 29133
rect 1864 29099 1870 29133
rect 1824 29061 1870 29099
rect 1824 29027 1830 29061
rect 1864 29027 1870 29061
rect 1824 28989 1870 29027
rect 1824 28955 1830 28989
rect 1864 28955 1870 28989
rect 1824 28917 1870 28955
rect 1824 28883 1830 28917
rect 1864 28883 1870 28917
rect 1824 28845 1870 28883
rect 1824 28811 1830 28845
rect 1864 28811 1870 28845
rect 1824 28773 1870 28811
rect 1824 28739 1830 28773
rect 1864 28739 1870 28773
rect 1824 28701 1870 28739
rect 1824 28667 1830 28701
rect 1864 28667 1870 28701
rect 1824 28629 1870 28667
rect 1824 28595 1830 28629
rect 1864 28595 1870 28629
rect 1824 28557 1870 28595
rect 1824 28523 1830 28557
rect 1864 28523 1870 28557
rect 1824 28485 1870 28523
rect 1824 28451 1830 28485
rect 1864 28451 1870 28485
rect 1824 28413 1870 28451
rect 1824 28379 1830 28413
rect 1864 28379 1870 28413
rect 1824 28341 1870 28379
rect 1824 28307 1830 28341
rect 1864 28307 1870 28341
rect 1824 28269 1870 28307
rect 1824 28235 1830 28269
rect 1864 28235 1870 28269
rect 1824 28197 1870 28235
rect 1824 28163 1830 28197
rect 1864 28163 1870 28197
rect 1824 28125 1870 28163
rect 1824 28091 1830 28125
rect 1864 28091 1870 28125
rect 1824 28053 1870 28091
rect 1824 28019 1830 28053
rect 1864 28019 1870 28053
rect 1824 27981 1870 28019
rect 1824 27947 1830 27981
rect 1864 27947 1870 27981
rect 1824 27909 1870 27947
rect 1824 27875 1830 27909
rect 1864 27875 1870 27909
rect 1824 27837 1870 27875
rect 1824 27803 1830 27837
rect 1864 27803 1870 27837
rect 1824 27765 1870 27803
rect 1824 27731 1830 27765
rect 1864 27731 1870 27765
rect 1824 27693 1870 27731
rect 1824 27659 1830 27693
rect 1864 27659 1870 27693
rect 1824 27621 1870 27659
rect 1824 27587 1830 27621
rect 1864 27587 1870 27621
rect 1824 27549 1870 27587
rect 1824 27515 1830 27549
rect 1864 27515 1870 27549
rect 1824 27477 1870 27515
rect 1824 27443 1830 27477
rect 1864 27443 1870 27477
rect 1824 27405 1870 27443
rect 1824 27371 1830 27405
rect 1864 27371 1870 27405
rect 1824 27333 1870 27371
rect 1824 27299 1830 27333
rect 1864 27299 1870 27333
rect 1824 27261 1870 27299
rect 1824 27227 1830 27261
rect 1864 27227 1870 27261
rect 1824 27189 1870 27227
rect 1824 27155 1830 27189
rect 1864 27155 1870 27189
rect 1824 27117 1870 27155
rect 1824 27083 1830 27117
rect 1864 27083 1870 27117
rect 1824 27045 1870 27083
rect 1824 27011 1830 27045
rect 1864 27011 1870 27045
rect 1824 26973 1870 27011
rect 1824 26939 1830 26973
rect 1864 26939 1870 26973
rect 1824 26901 1870 26939
rect 1824 26867 1830 26901
rect 1864 26867 1870 26901
rect 1824 26829 1870 26867
rect 1824 26795 1830 26829
rect 1864 26795 1870 26829
rect 1824 26757 1870 26795
rect 1824 26723 1830 26757
rect 1864 26723 1870 26757
rect 1824 26685 1870 26723
rect 1824 26651 1830 26685
rect 1864 26651 1870 26685
rect 1824 26613 1870 26651
rect 1824 26579 1830 26613
rect 1864 26579 1870 26613
rect 1824 26541 1870 26579
rect 1824 26507 1830 26541
rect 1864 26507 1870 26541
rect 1824 26469 1870 26507
rect 1824 26435 1830 26469
rect 1864 26435 1870 26469
rect 1824 26397 1870 26435
rect 1824 26363 1830 26397
rect 1864 26363 1870 26397
rect 1824 26325 1870 26363
rect 1824 26291 1830 26325
rect 1864 26291 1870 26325
rect 1824 26253 1870 26291
rect 1824 26219 1830 26253
rect 1864 26219 1870 26253
rect 1824 26181 1870 26219
rect 1824 26147 1830 26181
rect 1864 26147 1870 26181
rect 1824 26109 1870 26147
rect 1824 26075 1830 26109
rect 1864 26075 1870 26109
rect 1824 26037 1870 26075
rect 1824 26003 1830 26037
rect 1864 26003 1870 26037
rect 1824 25965 1870 26003
rect 1824 25931 1830 25965
rect 1864 25931 1870 25965
rect 1824 25893 1870 25931
rect 1824 25859 1830 25893
rect 1864 25859 1870 25893
rect 1824 25821 1870 25859
rect 1824 25787 1830 25821
rect 1864 25787 1870 25821
rect 1824 25749 1870 25787
rect 1824 25715 1830 25749
rect 1864 25715 1870 25749
rect 1824 25677 1870 25715
rect 1824 25643 1830 25677
rect 1864 25643 1870 25677
rect 1824 25605 1870 25643
rect 1824 25571 1830 25605
rect 1864 25571 1870 25605
rect 1824 25533 1870 25571
rect 1824 25499 1830 25533
rect 1864 25499 1870 25533
rect 1824 25461 1870 25499
rect 1824 25427 1830 25461
rect 1864 25427 1870 25461
rect 1824 25389 1870 25427
rect 1824 25355 1830 25389
rect 1864 25355 1870 25389
rect 1824 25317 1870 25355
rect 1824 25283 1830 25317
rect 1864 25283 1870 25317
rect 1824 25245 1870 25283
rect 1824 25211 1830 25245
rect 1864 25211 1870 25245
rect 1824 25173 1870 25211
rect 1824 25139 1830 25173
rect 1864 25139 1870 25173
rect 1824 25101 1870 25139
rect 1824 25067 1830 25101
rect 1864 25067 1870 25101
rect 1824 25029 1870 25067
rect 1824 24995 1830 25029
rect 1864 24995 1870 25029
rect 1824 24957 1870 24995
rect 1824 24923 1830 24957
rect 1864 24923 1870 24957
rect 1824 24885 1870 24923
rect 1824 24851 1830 24885
rect 1864 24851 1870 24885
rect 1824 24813 1870 24851
rect 1824 24779 1830 24813
rect 1864 24779 1870 24813
rect 1824 24741 1870 24779
rect 1824 24707 1830 24741
rect 1864 24707 1870 24741
rect 1824 24669 1870 24707
rect 1824 24635 1830 24669
rect 1864 24635 1870 24669
rect 1824 24597 1870 24635
rect 1824 24563 1830 24597
rect 1864 24563 1870 24597
rect 1824 24525 1870 24563
rect 1824 24491 1830 24525
rect 1864 24491 1870 24525
rect 1824 24453 1870 24491
rect 1824 24419 1830 24453
rect 1864 24419 1870 24453
rect 1824 24381 1870 24419
rect 1824 24347 1830 24381
rect 1864 24347 1870 24381
rect 1824 24309 1870 24347
rect 1824 24275 1830 24309
rect 1864 24275 1870 24309
rect 1824 24237 1870 24275
rect 1824 24203 1830 24237
rect 1864 24203 1870 24237
rect 1824 24165 1870 24203
rect 1824 24131 1830 24165
rect 1864 24131 1870 24165
rect 1824 24093 1870 24131
rect 1824 24059 1830 24093
rect 1864 24059 1870 24093
rect 1824 24021 1870 24059
rect 1824 23987 1830 24021
rect 1864 23987 1870 24021
rect 1824 23949 1870 23987
rect 1824 23915 1830 23949
rect 1864 23915 1870 23949
rect 1824 23877 1870 23915
rect 1824 23843 1830 23877
rect 1864 23843 1870 23877
rect 1824 23805 1870 23843
rect 1824 23771 1830 23805
rect 1864 23771 1870 23805
rect 1824 23733 1870 23771
rect 1824 23699 1830 23733
rect 1864 23699 1870 23733
rect 1824 23661 1870 23699
rect 1824 23627 1830 23661
rect 1864 23627 1870 23661
rect 1824 23589 1870 23627
rect 1824 23555 1830 23589
rect 1864 23555 1870 23589
rect 1824 23517 1870 23555
rect 1824 23483 1830 23517
rect 1864 23483 1870 23517
rect 1824 23445 1870 23483
rect 1824 23411 1830 23445
rect 1864 23411 1870 23445
rect 1824 23373 1870 23411
rect 1824 23339 1830 23373
rect 1864 23339 1870 23373
rect 1824 23301 1870 23339
rect 1824 23267 1830 23301
rect 1864 23267 1870 23301
rect 1824 23229 1870 23267
rect 1824 23195 1830 23229
rect 1864 23195 1870 23229
rect 1824 23157 1870 23195
rect 1824 23123 1830 23157
rect 1864 23123 1870 23157
rect 1824 23085 1870 23123
rect 1824 23051 1830 23085
rect 1864 23051 1870 23085
rect 1824 23013 1870 23051
rect 1824 22979 1830 23013
rect 1864 22979 1870 23013
rect 1824 22941 1870 22979
rect 1824 22907 1830 22941
rect 1864 22907 1870 22941
rect 1824 22869 1870 22907
rect 1824 22835 1830 22869
rect 1864 22835 1870 22869
rect 1824 22797 1870 22835
rect 1824 22763 1830 22797
rect 1864 22763 1870 22797
rect 1824 22725 1870 22763
rect 1824 22691 1830 22725
rect 1864 22691 1870 22725
rect 1824 22653 1870 22691
rect 1824 22619 1830 22653
rect 1864 22619 1870 22653
rect 1824 22581 1870 22619
rect 1824 22547 1830 22581
rect 1864 22547 1870 22581
rect 1824 22509 1870 22547
rect 1824 22475 1830 22509
rect 1864 22475 1870 22509
rect 1824 22437 1870 22475
rect 1824 22403 1830 22437
rect 1864 22403 1870 22437
rect 1824 22365 1870 22403
rect 1824 22331 1830 22365
rect 1864 22331 1870 22365
rect 1824 22293 1870 22331
rect 1824 22259 1830 22293
rect 1864 22259 1870 22293
rect 1824 22221 1870 22259
rect 1824 22187 1830 22221
rect 1864 22187 1870 22221
rect 1824 22149 1870 22187
rect 1824 22115 1830 22149
rect 1864 22115 1870 22149
rect 1824 22077 1870 22115
rect 1824 22043 1830 22077
rect 1864 22043 1870 22077
rect 1824 22005 1870 22043
rect 1824 21971 1830 22005
rect 1864 21971 1870 22005
rect 1824 21933 1870 21971
rect 1824 21899 1830 21933
rect 1864 21899 1870 21933
rect 1824 21861 1870 21899
rect 1824 21827 1830 21861
rect 1864 21827 1870 21861
rect 1824 21789 1870 21827
rect 1824 21755 1830 21789
rect 1864 21755 1870 21789
rect 1824 21717 1870 21755
rect 1824 21683 1830 21717
rect 1864 21683 1870 21717
rect 1824 21645 1870 21683
rect 1824 21611 1830 21645
rect 1864 21611 1870 21645
rect 1824 21573 1870 21611
rect 1824 21539 1830 21573
rect 1864 21539 1870 21573
rect 1824 21501 1870 21539
rect 1824 21467 1830 21501
rect 1864 21467 1870 21501
rect 1824 21429 1870 21467
rect 1824 21395 1830 21429
rect 1864 21395 1870 21429
rect 1824 21357 1870 21395
rect 1824 21323 1830 21357
rect 1864 21323 1870 21357
rect 1824 21285 1870 21323
rect 1824 21251 1830 21285
rect 1864 21251 1870 21285
rect 1824 21213 1870 21251
rect 1824 21179 1830 21213
rect 1864 21179 1870 21213
rect 1824 21141 1870 21179
rect 1824 21107 1830 21141
rect 1864 21107 1870 21141
rect 1824 21069 1870 21107
rect 1824 21035 1830 21069
rect 1864 21035 1870 21069
rect 1824 20997 1870 21035
rect 1824 20963 1830 20997
rect 1864 20963 1870 20997
rect 1824 20925 1870 20963
rect 1824 20891 1830 20925
rect 1864 20891 1870 20925
rect 1824 20853 1870 20891
rect 1824 20819 1830 20853
rect 1864 20819 1870 20853
rect 1824 20781 1870 20819
rect 1824 20747 1830 20781
rect 1864 20747 1870 20781
rect 1824 20709 1870 20747
rect 1824 20675 1830 20709
rect 1864 20675 1870 20709
rect 1824 20637 1870 20675
rect 1824 20603 1830 20637
rect 1864 20603 1870 20637
rect 1824 20565 1870 20603
rect 1824 20531 1830 20565
rect 1864 20531 1870 20565
rect 1824 20493 1870 20531
rect 1824 20459 1830 20493
rect 1864 20459 1870 20493
rect 1824 20421 1870 20459
rect 1824 20387 1830 20421
rect 1864 20387 1870 20421
rect 1824 20349 1870 20387
rect 1824 20315 1830 20349
rect 1864 20315 1870 20349
rect 1824 20277 1870 20315
rect 1824 20243 1830 20277
rect 1864 20243 1870 20277
rect 1824 20205 1870 20243
rect 1824 20171 1830 20205
rect 1864 20171 1870 20205
rect 1824 20133 1870 20171
rect 1824 20099 1830 20133
rect 1864 20099 1870 20133
rect 1824 20061 1870 20099
rect 1824 20027 1830 20061
rect 1864 20027 1870 20061
rect 1824 19989 1870 20027
rect 1824 19955 1830 19989
rect 1864 19955 1870 19989
rect 1824 19917 1870 19955
rect 1824 19883 1830 19917
rect 1864 19883 1870 19917
rect 1824 19845 1870 19883
rect 1824 19811 1830 19845
rect 1864 19811 1870 19845
rect 1824 19773 1870 19811
rect 1824 19739 1830 19773
rect 1864 19739 1870 19773
rect 1824 19701 1870 19739
rect 1824 19667 1830 19701
rect 1864 19667 1870 19701
rect 1824 19629 1870 19667
rect 1824 19595 1830 19629
rect 1864 19595 1870 19629
rect 1824 19557 1870 19595
rect 1824 19523 1830 19557
rect 1864 19523 1870 19557
rect 1824 19485 1870 19523
rect 1824 19451 1830 19485
rect 1864 19451 1870 19485
rect 1824 19413 1870 19451
rect 1824 19379 1830 19413
rect 1864 19379 1870 19413
rect 1824 19341 1870 19379
rect 1824 19307 1830 19341
rect 1864 19307 1870 19341
rect 1824 19269 1870 19307
rect 1824 19235 1830 19269
rect 1864 19235 1870 19269
rect 1824 19197 1870 19235
rect 1824 19163 1830 19197
rect 1864 19163 1870 19197
rect 1824 19125 1870 19163
rect 1824 19091 1830 19125
rect 1864 19091 1870 19125
rect 1824 19053 1870 19091
rect 1824 19019 1830 19053
rect 1864 19019 1870 19053
rect 1824 18981 1870 19019
rect 1824 18947 1830 18981
rect 1864 18947 1870 18981
rect 1824 18909 1870 18947
rect 1824 18875 1830 18909
rect 1864 18875 1870 18909
rect 1824 18837 1870 18875
rect 1824 18803 1830 18837
rect 1864 18803 1870 18837
rect 1824 18765 1870 18803
rect 1824 18731 1830 18765
rect 1864 18731 1870 18765
rect 1824 18693 1870 18731
rect 1824 18659 1830 18693
rect 1864 18659 1870 18693
rect 1824 18621 1870 18659
rect 1824 18587 1830 18621
rect 1864 18587 1870 18621
rect 1824 18549 1870 18587
rect 1824 18515 1830 18549
rect 1864 18515 1870 18549
rect 1824 18477 1870 18515
rect 1824 18443 1830 18477
rect 1864 18443 1870 18477
rect 1824 18405 1870 18443
rect 1824 18371 1830 18405
rect 1864 18371 1870 18405
rect 1824 18333 1870 18371
rect 1824 18299 1830 18333
rect 1864 18299 1870 18333
rect 1824 18261 1870 18299
rect 1824 18227 1830 18261
rect 1864 18227 1870 18261
rect 1824 18189 1870 18227
rect 1824 18155 1830 18189
rect 1864 18155 1870 18189
rect 1824 18117 1870 18155
rect 1824 18083 1830 18117
rect 1864 18083 1870 18117
rect 1824 18045 1870 18083
rect 1824 18011 1830 18045
rect 1864 18011 1870 18045
rect 1824 17973 1870 18011
rect 1824 17939 1830 17973
rect 1864 17939 1870 17973
rect 1824 17901 1870 17939
rect 1824 17867 1830 17901
rect 1864 17867 1870 17901
rect 1824 17829 1870 17867
rect 1824 17795 1830 17829
rect 1864 17795 1870 17829
rect 1824 17757 1870 17795
rect 1824 17723 1830 17757
rect 1864 17723 1870 17757
rect 1824 17685 1870 17723
rect 1824 17651 1830 17685
rect 1864 17651 1870 17685
rect 1824 17613 1870 17651
rect 1824 17579 1830 17613
rect 1864 17579 1870 17613
rect 1824 17541 1870 17579
rect 1824 17507 1830 17541
rect 1864 17507 1870 17541
rect 1824 17469 1870 17507
rect 1824 17435 1830 17469
rect 1864 17435 1870 17469
rect 1824 17397 1870 17435
rect 1824 17363 1830 17397
rect 1864 17363 1870 17397
rect 1824 17325 1870 17363
rect 1824 17291 1830 17325
rect 1864 17291 1870 17325
rect 1824 17253 1870 17291
rect 1824 17219 1830 17253
rect 1864 17219 1870 17253
rect 1824 17181 1870 17219
rect 1824 17147 1830 17181
rect 1864 17147 1870 17181
rect 1824 17109 1870 17147
rect 1824 17075 1830 17109
rect 1864 17075 1870 17109
rect 1824 17037 1870 17075
rect 1824 17003 1830 17037
rect 1864 17003 1870 17037
rect 1824 16965 1870 17003
rect 1824 16931 1830 16965
rect 1864 16931 1870 16965
rect 1824 16893 1870 16931
rect 1824 16859 1830 16893
rect 1864 16859 1870 16893
rect 1824 16821 1870 16859
rect 1824 16787 1830 16821
rect 1864 16787 1870 16821
rect 1824 16749 1870 16787
rect 1824 16715 1830 16749
rect 1864 16715 1870 16749
rect 1824 16677 1870 16715
rect 1824 16643 1830 16677
rect 1864 16643 1870 16677
rect 1824 16605 1870 16643
rect 1824 16571 1830 16605
rect 1864 16571 1870 16605
rect 1824 16533 1870 16571
rect 1824 16499 1830 16533
rect 1864 16499 1870 16533
rect 1824 16461 1870 16499
rect 1824 16427 1830 16461
rect 1864 16427 1870 16461
rect 1824 16389 1870 16427
rect 1824 16355 1830 16389
rect 1864 16355 1870 16389
rect 1824 16317 1870 16355
rect 1824 16283 1830 16317
rect 1864 16283 1870 16317
rect 1824 16245 1870 16283
rect 1824 16211 1830 16245
rect 1864 16211 1870 16245
rect 1824 16173 1870 16211
rect 1824 16139 1830 16173
rect 1864 16139 1870 16173
rect 1824 16101 1870 16139
rect 1824 16067 1830 16101
rect 1864 16067 1870 16101
rect 1824 16029 1870 16067
rect 1824 15995 1830 16029
rect 1864 15995 1870 16029
rect 1824 15957 1870 15995
rect 1824 15923 1830 15957
rect 1864 15923 1870 15957
rect 1824 15885 1870 15923
rect 1824 15851 1830 15885
rect 1864 15851 1870 15885
rect 1824 15813 1870 15851
rect 1824 15779 1830 15813
rect 1864 15779 1870 15813
rect 1824 15741 1870 15779
rect 1824 15707 1830 15741
rect 1864 15707 1870 15741
rect 1824 15669 1870 15707
rect 1824 15635 1830 15669
rect 1864 15635 1870 15669
rect 1824 15597 1870 15635
rect 1824 15563 1830 15597
rect 1864 15563 1870 15597
rect 1824 15525 1870 15563
rect 1824 15491 1830 15525
rect 1864 15491 1870 15525
rect 1824 15453 1870 15491
rect 1824 15419 1830 15453
rect 1864 15419 1870 15453
rect 1824 15381 1870 15419
rect 1824 15347 1830 15381
rect 1864 15347 1870 15381
rect 1824 15309 1870 15347
rect 1824 15275 1830 15309
rect 1864 15275 1870 15309
rect 1824 15237 1870 15275
rect 1824 15203 1830 15237
rect 1864 15203 1870 15237
rect 1824 15165 1870 15203
rect 1824 15131 1830 15165
rect 1864 15131 1870 15165
rect 1824 15093 1870 15131
rect 1824 15059 1830 15093
rect 1864 15059 1870 15093
rect 1824 15021 1870 15059
rect 1824 14987 1830 15021
rect 1864 14987 1870 15021
rect 1824 14949 1870 14987
rect 1824 14915 1830 14949
rect 1864 14915 1870 14949
rect 1824 14877 1870 14915
rect 1824 14843 1830 14877
rect 1864 14843 1870 14877
rect 1824 14805 1870 14843
rect 1824 14771 1830 14805
rect 1864 14771 1870 14805
rect 1824 14733 1870 14771
rect 1824 14699 1830 14733
rect 1864 14699 1870 14733
rect 1824 14661 1870 14699
rect 1824 14627 1830 14661
rect 1864 14627 1870 14661
rect 1824 14589 1870 14627
rect 1824 14555 1830 14589
rect 1864 14555 1870 14589
rect 1824 14517 1870 14555
rect 1824 14483 1830 14517
rect 1864 14483 1870 14517
rect 1824 14445 1870 14483
rect 1824 14411 1830 14445
rect 1864 14411 1870 14445
rect 1824 14373 1870 14411
rect 1824 14339 1830 14373
rect 1864 14339 1870 14373
rect 1824 14301 1870 14339
rect 1824 14267 1830 14301
rect 1864 14267 1870 14301
rect 1824 14229 1870 14267
rect 1824 14195 1830 14229
rect 1864 14195 1870 14229
rect 1824 14157 1870 14195
rect 1824 14123 1830 14157
rect 1864 14123 1870 14157
rect 1824 14085 1870 14123
rect 1824 14051 1830 14085
rect 1864 14051 1870 14085
rect 1824 14013 1870 14051
rect 1824 13979 1830 14013
rect 1864 13979 1870 14013
rect 1824 13941 1870 13979
rect 1824 13907 1830 13941
rect 1864 13907 1870 13941
rect 1824 13869 1870 13907
rect 1824 13835 1830 13869
rect 1864 13835 1870 13869
rect 1824 13797 1870 13835
rect 1824 13763 1830 13797
rect 1864 13763 1870 13797
rect 1824 13725 1870 13763
rect 1824 13691 1830 13725
rect 1864 13691 1870 13725
rect 1824 13653 1870 13691
rect 1824 13619 1830 13653
rect 1864 13619 1870 13653
rect 1824 13581 1870 13619
rect 1824 13547 1830 13581
rect 1864 13547 1870 13581
rect 1824 13509 1870 13547
rect 1824 13475 1830 13509
rect 1864 13475 1870 13509
rect 1824 13437 1870 13475
rect 1824 13403 1830 13437
rect 1864 13403 1870 13437
rect 1824 13365 1870 13403
rect 1824 13331 1830 13365
rect 1864 13331 1870 13365
rect 1824 13293 1870 13331
rect 1824 13259 1830 13293
rect 1864 13259 1870 13293
rect 1824 13221 1870 13259
rect 1824 13187 1830 13221
rect 1864 13187 1870 13221
rect 1824 13149 1870 13187
rect 1824 13115 1830 13149
rect 1864 13115 1870 13149
rect 1824 13077 1870 13115
rect 1824 13043 1830 13077
rect 1864 13043 1870 13077
rect 1824 13005 1870 13043
rect 1824 12971 1830 13005
rect 1864 12971 1870 13005
rect 1824 12933 1870 12971
rect 1824 12899 1830 12933
rect 1864 12899 1870 12933
rect 1824 12861 1870 12899
rect 1824 12827 1830 12861
rect 1864 12827 1870 12861
rect 1824 12789 1870 12827
rect 1824 12755 1830 12789
rect 1864 12755 1870 12789
rect 1824 12717 1870 12755
rect 1824 12683 1830 12717
rect 1864 12683 1870 12717
rect 1824 12645 1870 12683
rect 1824 12611 1830 12645
rect 1864 12611 1870 12645
rect 1824 12573 1870 12611
rect 1824 12539 1830 12573
rect 1864 12539 1870 12573
rect 1824 12501 1870 12539
rect 1824 12467 1830 12501
rect 1864 12467 1870 12501
rect 1824 12429 1870 12467
rect 1824 12395 1830 12429
rect 1864 12395 1870 12429
rect 1824 12357 1870 12395
rect 1824 12323 1830 12357
rect 1864 12323 1870 12357
rect 1824 12285 1870 12323
rect 1824 12251 1830 12285
rect 1864 12251 1870 12285
rect 1824 12213 1870 12251
rect 1824 12179 1830 12213
rect 1864 12179 1870 12213
rect 1824 12141 1870 12179
rect 1824 12107 1830 12141
rect 1864 12107 1870 12141
rect 1824 12069 1870 12107
rect 1824 12035 1830 12069
rect 1864 12035 1870 12069
rect 1824 11997 1870 12035
rect 1824 11963 1830 11997
rect 1864 11963 1870 11997
rect 1824 11925 1870 11963
rect 1824 11891 1830 11925
rect 1864 11891 1870 11925
rect 1824 11853 1870 11891
rect 1824 11819 1830 11853
rect 1864 11819 1870 11853
rect 1824 11781 1870 11819
rect 1824 11747 1830 11781
rect 1864 11747 1870 11781
rect 1824 11709 1870 11747
rect 1824 11675 1830 11709
rect 1864 11675 1870 11709
rect 1824 11637 1870 11675
rect 1824 11603 1830 11637
rect 1864 11603 1870 11637
rect 1824 11565 1870 11603
rect 1824 11531 1830 11565
rect 1864 11531 1870 11565
rect 1824 11493 1870 11531
rect 1824 11459 1830 11493
rect 1864 11459 1870 11493
rect 1824 11421 1870 11459
rect 1824 11387 1830 11421
rect 1864 11387 1870 11421
rect 1824 11349 1870 11387
rect 1824 11315 1830 11349
rect 1864 11315 1870 11349
rect 1824 11277 1870 11315
rect 1824 11243 1830 11277
rect 1864 11243 1870 11277
rect 1824 11205 1870 11243
rect 1824 11171 1830 11205
rect 1864 11171 1870 11205
rect 1824 11133 1870 11171
rect 1824 11099 1830 11133
rect 1864 11099 1870 11133
rect 1824 11061 1870 11099
rect 1824 11027 1830 11061
rect 1864 11027 1870 11061
rect 1824 10989 1870 11027
rect 1824 10955 1830 10989
rect 1864 10955 1870 10989
rect 1824 10917 1870 10955
rect 1824 10883 1830 10917
rect 1864 10883 1870 10917
rect 1824 10845 1870 10883
rect 1824 10811 1830 10845
rect 1864 10811 1870 10845
rect 1824 10773 1870 10811
rect 1824 10739 1830 10773
rect 1864 10739 1870 10773
rect 1824 10701 1870 10739
rect 1824 10667 1830 10701
rect 1864 10667 1870 10701
rect 1824 10629 1870 10667
rect 1824 10595 1830 10629
rect 1864 10595 1870 10629
rect 1824 10557 1870 10595
rect 1824 10523 1830 10557
rect 1864 10523 1870 10557
rect 1824 10485 1870 10523
rect 1824 10451 1830 10485
rect 1864 10451 1870 10485
rect 1824 10413 1870 10451
rect 1824 10379 1830 10413
rect 1864 10379 1870 10413
rect 1824 10341 1870 10379
rect 1824 10307 1830 10341
rect 1864 10307 1870 10341
rect 1824 10269 1870 10307
rect 1824 10235 1830 10269
rect 1864 10235 1870 10269
rect 1824 10197 1870 10235
rect 1824 10163 1830 10197
rect 1864 10163 1870 10197
rect 1824 10125 1870 10163
rect 1824 10091 1830 10125
rect 1864 10091 1870 10125
rect 1824 10053 1870 10091
rect 1824 10019 1830 10053
rect 1864 10019 1870 10053
rect 1824 9981 1870 10019
rect 1824 9947 1830 9981
rect 1864 9947 1870 9981
rect 1824 9909 1870 9947
rect 1824 9875 1830 9909
rect 1864 9875 1870 9909
rect 1824 9837 1870 9875
rect 1824 9803 1830 9837
rect 1864 9803 1870 9837
rect 1824 9765 1870 9803
rect 1824 9731 1830 9765
rect 1864 9731 1870 9765
rect 1824 9693 1870 9731
rect 1824 9659 1830 9693
rect 1864 9659 1870 9693
rect 1824 9621 1870 9659
rect 1824 9587 1830 9621
rect 1864 9587 1870 9621
rect 1824 9549 1870 9587
rect 1824 9515 1830 9549
rect 1864 9515 1870 9549
rect 1824 9477 1870 9515
rect 1824 9443 1830 9477
rect 1864 9443 1870 9477
rect 1824 9405 1870 9443
rect 1824 9371 1830 9405
rect 1864 9371 1870 9405
rect 1824 9333 1870 9371
rect 1824 9299 1830 9333
rect 1864 9299 1870 9333
rect 1824 9261 1870 9299
rect 1824 9227 1830 9261
rect 1864 9227 1870 9261
rect 1824 9189 1870 9227
rect 1824 9155 1830 9189
rect 1864 9155 1870 9189
rect 1824 9117 1870 9155
rect 1824 9083 1830 9117
rect 1864 9083 1870 9117
rect 1824 9045 1870 9083
rect 1824 9011 1830 9045
rect 1864 9011 1870 9045
rect 1824 8973 1870 9011
rect 1824 8939 1830 8973
rect 1864 8939 1870 8973
rect 1824 8901 1870 8939
rect 1824 8867 1830 8901
rect 1864 8867 1870 8901
rect 1824 8829 1870 8867
rect 1824 8795 1830 8829
rect 1864 8795 1870 8829
rect 1824 8757 1870 8795
rect 1824 8723 1830 8757
rect 1864 8723 1870 8757
rect 1824 8685 1870 8723
rect 1824 8651 1830 8685
rect 1864 8651 1870 8685
rect 1824 8613 1870 8651
rect 1824 8579 1830 8613
rect 1864 8579 1870 8613
rect 1824 8541 1870 8579
rect 1824 8507 1830 8541
rect 1864 8507 1870 8541
rect 1824 8469 1870 8507
rect 1824 8435 1830 8469
rect 1864 8435 1870 8469
rect 1824 8397 1870 8435
rect 1824 8363 1830 8397
rect 1864 8363 1870 8397
rect 1824 8325 1870 8363
rect 1824 8291 1830 8325
rect 1864 8291 1870 8325
rect 1824 8253 1870 8291
rect 1824 8219 1830 8253
rect 1864 8219 1870 8253
rect 1824 8181 1870 8219
rect 1824 8147 1830 8181
rect 1864 8147 1870 8181
rect 1824 8109 1870 8147
rect 1824 8075 1830 8109
rect 1864 8075 1870 8109
rect 1824 8037 1870 8075
rect 1824 8003 1830 8037
rect 1864 8003 1870 8037
rect 1824 7965 1870 8003
rect 1824 7931 1830 7965
rect 1864 7931 1870 7965
rect 1824 7893 1870 7931
rect 1824 7859 1830 7893
rect 1864 7859 1870 7893
rect 1824 7821 1870 7859
rect 1824 7787 1830 7821
rect 1864 7787 1870 7821
rect 1824 7749 1870 7787
rect 1824 7715 1830 7749
rect 1864 7715 1870 7749
rect 1824 7677 1870 7715
rect 1824 7643 1830 7677
rect 1864 7643 1870 7677
rect 1824 7605 1870 7643
rect 1824 7571 1830 7605
rect 1864 7571 1870 7605
rect 1824 7533 1870 7571
rect 1824 7499 1830 7533
rect 1864 7499 1870 7533
rect 1824 7461 1870 7499
rect 1824 7427 1830 7461
rect 1864 7427 1870 7461
rect 1824 7389 1870 7427
rect 1824 7355 1830 7389
rect 1864 7355 1870 7389
rect 1824 7317 1870 7355
rect 1824 7283 1830 7317
rect 1864 7283 1870 7317
rect 1824 7245 1870 7283
rect 1824 7211 1830 7245
rect 1864 7211 1870 7245
rect 1824 7173 1870 7211
rect 1824 7139 1830 7173
rect 1864 7139 1870 7173
rect 1824 7101 1870 7139
rect 1824 7067 1830 7101
rect 1864 7067 1870 7101
rect 1824 7029 1870 7067
rect 1824 6995 1830 7029
rect 1864 6995 1870 7029
rect 1824 6957 1870 6995
rect 1824 6923 1830 6957
rect 1864 6923 1870 6957
rect 1824 6885 1870 6923
rect 1824 6851 1830 6885
rect 1864 6851 1870 6885
rect 1824 6813 1870 6851
rect 1824 6779 1830 6813
rect 1864 6779 1870 6813
rect 1824 6741 1870 6779
rect 1824 6707 1830 6741
rect 1864 6707 1870 6741
rect 1824 6669 1870 6707
rect 1824 6635 1830 6669
rect 1864 6635 1870 6669
rect 1824 6597 1870 6635
rect 1824 6563 1830 6597
rect 1864 6563 1870 6597
rect 1824 6525 1870 6563
rect 1824 6491 1830 6525
rect 1864 6491 1870 6525
rect 1824 6453 1870 6491
rect 1824 6419 1830 6453
rect 1864 6419 1870 6453
rect 1824 6381 1870 6419
rect 1824 6347 1830 6381
rect 1864 6347 1870 6381
rect 1824 6309 1870 6347
rect 1824 6275 1830 6309
rect 1864 6275 1870 6309
rect 1824 6237 1870 6275
rect 1824 6203 1830 6237
rect 1864 6203 1870 6237
rect 1824 6165 1870 6203
rect 1824 6131 1830 6165
rect 1864 6131 1870 6165
rect 1824 6093 1870 6131
rect 1824 6059 1830 6093
rect 1864 6059 1870 6093
rect 1824 6021 1870 6059
rect 1824 5987 1830 6021
rect 1864 5987 1870 6021
rect 1824 5949 1870 5987
rect 1824 5915 1830 5949
rect 1864 5915 1870 5949
rect 1824 5877 1870 5915
rect 1824 5843 1830 5877
rect 1864 5843 1870 5877
rect 1824 5805 1870 5843
rect 1824 5771 1830 5805
rect 1864 5771 1870 5805
rect 1824 5733 1870 5771
rect 1824 5699 1830 5733
rect 1864 5699 1870 5733
rect 1824 5661 1870 5699
rect 1824 5627 1830 5661
rect 1864 5627 1870 5661
rect 1824 5589 1870 5627
rect 1824 5555 1830 5589
rect 1864 5555 1870 5589
rect 1824 5517 1870 5555
rect 1824 5483 1830 5517
rect 1864 5483 1870 5517
rect 1824 5445 1870 5483
rect 1824 5411 1830 5445
rect 1864 5411 1870 5445
rect 1824 5373 1870 5411
rect 1824 5339 1830 5373
rect 1864 5339 1870 5373
rect 1824 5301 1870 5339
rect 1824 5267 1830 5301
rect 1864 5267 1870 5301
rect 1824 5229 1870 5267
rect 1824 5195 1830 5229
rect 1864 5195 1870 5229
rect 1824 5157 1870 5195
rect 1824 5123 1830 5157
rect 1864 5123 1870 5157
rect 1824 5085 1870 5123
rect 1824 5051 1830 5085
rect 1864 5051 1870 5085
rect 1824 5013 1870 5051
rect 1824 4979 1830 5013
rect 1864 4979 1870 5013
rect 1824 4941 1870 4979
rect 1824 4907 1830 4941
rect 1864 4907 1870 4941
rect 1824 4869 1870 4907
rect 1824 4835 1830 4869
rect 1864 4835 1870 4869
rect 1824 4797 1870 4835
rect 1824 4763 1830 4797
rect 1864 4763 1870 4797
rect 1824 4725 1870 4763
rect 1824 4691 1830 4725
rect 1864 4691 1870 4725
rect 1824 4653 1870 4691
rect -258 4581 -212 4619
rect -258 4547 -252 4581
rect -218 4547 -212 4581
rect -258 4509 -212 4547
rect -258 4475 -252 4509
rect -218 4475 -212 4509
rect -258 4437 -212 4475
rect -258 4403 -252 4437
rect -218 4403 -212 4437
rect -258 4365 -212 4403
rect -258 4331 -252 4365
rect -218 4331 -212 4365
rect -258 4293 -212 4331
rect -258 4259 -252 4293
rect -218 4259 -212 4293
rect -258 4221 -212 4259
rect -258 4187 -252 4221
rect -218 4187 -212 4221
rect -258 4149 -212 4187
rect -258 4115 -252 4149
rect -218 4115 -212 4149
rect -258 4077 -212 4115
rect -258 4043 -252 4077
rect -218 4043 -212 4077
rect -258 4005 -212 4043
rect -258 3971 -252 4005
rect -218 3971 -212 4005
rect -258 3933 -212 3971
rect -258 3899 -252 3933
rect -218 3899 -212 3933
rect -258 3861 -212 3899
rect -258 3827 -252 3861
rect -218 3827 -212 3861
rect -258 3789 -212 3827
rect -258 3755 -252 3789
rect -218 3755 -212 3789
rect -258 3717 -212 3755
rect -258 3683 -252 3717
rect -218 3683 -212 3717
rect -258 3645 -212 3683
rect -258 3611 -252 3645
rect -218 3611 -212 3645
rect -258 3573 -212 3611
rect -258 3539 -252 3573
rect -218 3539 -212 3573
rect -258 3501 -212 3539
rect -258 3467 -252 3501
rect -218 3467 -212 3501
rect -258 3429 -212 3467
rect -258 3395 -252 3429
rect -218 3395 -212 3429
rect -258 3357 -212 3395
rect -135 4628 -83 4644
rect -135 4564 -83 4576
rect -135 3492 -83 4512
rect 1824 4619 1830 4653
rect 1864 4619 1870 4653
rect 1824 4581 1870 4619
rect 1824 4547 1830 4581
rect 1864 4547 1870 4581
rect 1824 4509 1870 4547
rect 1824 4475 1830 4509
rect 1864 4475 1870 4509
rect 1824 4437 1870 4475
rect 1824 4403 1830 4437
rect 1864 4403 1870 4437
rect 1824 4365 1870 4403
rect 1824 4331 1830 4365
rect 1864 4331 1870 4365
rect 1824 4293 1870 4331
rect 1824 4259 1830 4293
rect 1864 4259 1870 4293
rect 1824 4221 1870 4259
rect 1824 4187 1830 4221
rect 1864 4187 1870 4221
rect 1824 4149 1870 4187
rect 1824 4115 1830 4149
rect 1864 4115 1870 4149
rect 1824 4077 1870 4115
rect 1824 4043 1830 4077
rect 1864 4043 1870 4077
rect 1824 4005 1870 4043
rect 1824 3971 1830 4005
rect 1864 3971 1870 4005
rect 1824 3933 1870 3971
rect 1824 3899 1830 3933
rect 1864 3899 1870 3933
rect 1824 3861 1870 3899
rect 1824 3827 1830 3861
rect 1864 3827 1870 3861
rect 1824 3789 1870 3827
rect 1824 3755 1830 3789
rect 1864 3755 1870 3789
rect 1824 3717 1870 3755
rect 1824 3683 1830 3717
rect 1864 3683 1870 3717
rect 1824 3645 1870 3683
rect 1824 3611 1830 3645
rect 1864 3611 1870 3645
rect 1824 3573 1870 3611
rect 1824 3539 1830 3573
rect 1864 3539 1870 3573
rect 1824 3501 1870 3539
rect -135 3428 -83 3440
rect -135 3368 -83 3376
rect -17 3486 153 3498
rect -17 3452 -8 3486
rect 26 3452 110 3486
rect 144 3452 153 3486
rect -17 3414 153 3452
rect -17 3380 -8 3414
rect 26 3380 110 3414
rect 144 3380 153 3414
rect -17 3368 153 3380
rect 219 3486 389 3498
rect 219 3452 228 3486
rect 262 3452 346 3486
rect 380 3452 389 3486
rect 219 3414 389 3452
rect 219 3380 228 3414
rect 262 3380 346 3414
rect 380 3380 389 3414
rect 219 3368 389 3380
rect 455 3486 625 3498
rect 455 3452 464 3486
rect 498 3452 582 3486
rect 616 3452 625 3486
rect 455 3414 625 3452
rect 455 3380 464 3414
rect 498 3380 582 3414
rect 616 3380 625 3414
rect 455 3368 625 3380
rect 694 3486 858 3498
rect 694 3452 700 3486
rect 734 3452 818 3486
rect 852 3452 858 3486
rect 694 3414 858 3452
rect 694 3380 700 3414
rect 734 3380 818 3414
rect 852 3380 858 3414
rect 694 3368 858 3380
rect 930 3486 1094 3498
rect 930 3452 936 3486
rect 970 3452 1054 3486
rect 1088 3452 1094 3486
rect 930 3414 1094 3452
rect 930 3380 936 3414
rect 970 3380 1054 3414
rect 1088 3380 1094 3414
rect 930 3368 1094 3380
rect 1166 3486 1330 3498
rect 1166 3452 1172 3486
rect 1206 3452 1290 3486
rect 1324 3452 1330 3486
rect 1166 3414 1330 3452
rect 1166 3380 1172 3414
rect 1206 3380 1290 3414
rect 1324 3380 1330 3414
rect 1166 3368 1330 3380
rect 1402 3486 1566 3498
rect 1402 3452 1408 3486
rect 1442 3452 1526 3486
rect 1560 3452 1566 3486
rect 1402 3414 1566 3452
rect 1402 3380 1408 3414
rect 1442 3380 1526 3414
rect 1560 3380 1566 3414
rect 1402 3368 1566 3380
rect 1635 3492 1687 3498
rect 1635 3428 1687 3440
rect 1635 3368 1687 3376
rect 1824 3467 1830 3501
rect 1864 3467 1870 3501
rect 3966 38651 3972 38685
rect 4006 38651 4012 38685
tri 4012 38683 4014 38685 nw
tri 6106 38683 6108 38685 ne
rect 3966 38612 4012 38651
rect 3966 38578 3972 38612
rect 4006 38578 4012 38612
rect 3966 38539 4012 38578
rect 3966 38505 3972 38539
rect 4006 38505 4012 38539
rect 3966 38466 4012 38505
rect 3966 38432 3972 38466
rect 4006 38432 4012 38466
rect 3966 38393 4012 38432
rect 3966 38359 3972 38393
rect 4006 38359 4012 38393
rect 3966 38320 4012 38359
rect 3966 38286 3972 38320
rect 4006 38286 4012 38320
rect 3966 38247 4012 38286
rect 3966 38213 3972 38247
rect 4006 38213 4012 38247
rect 3966 38174 4012 38213
rect 3966 38140 3972 38174
rect 4006 38140 4012 38174
rect 3966 38101 4012 38140
rect 3966 38067 3972 38101
rect 4006 38067 4012 38101
rect 3966 38028 4012 38067
rect 3966 37994 3972 38028
rect 4006 37994 4012 38028
rect 3966 37955 4012 37994
rect 3966 37921 3972 37955
rect 4006 37921 4012 37955
rect 3966 37882 4012 37921
rect 3966 37848 3972 37882
rect 4006 37848 4012 37882
rect 3966 37809 4012 37848
rect 3966 37775 3972 37809
rect 4006 37775 4012 37809
rect 3966 37736 4012 37775
rect 3966 37702 3972 37736
rect 4006 37702 4012 37736
rect 3966 37663 4012 37702
rect 3966 37629 3972 37663
rect 4006 37629 4012 37663
rect 3966 37590 4012 37629
rect 3966 37556 3972 37590
rect 4006 37556 4012 37590
rect 3966 37517 4012 37556
rect 3966 37483 3972 37517
rect 4006 37483 4012 37517
rect 3966 37444 4012 37483
rect 3966 37410 3972 37444
rect 4006 37410 4012 37444
rect 3966 37371 4012 37410
rect 3966 37337 3972 37371
rect 4006 37337 4012 37371
rect 3966 37298 4012 37337
rect 3966 37264 3972 37298
rect 4006 37264 4012 37298
rect 3966 37225 4012 37264
rect 3966 37191 3972 37225
rect 4006 37191 4012 37225
rect 3966 37152 4012 37191
rect 3966 37118 3972 37152
rect 4006 37118 4012 37152
rect 3966 37079 4012 37118
rect 3966 37045 3972 37079
rect 4006 37045 4012 37079
rect 3966 37006 4012 37045
rect 3966 36972 3972 37006
rect 4006 36972 4012 37006
rect 3966 36933 4012 36972
rect 3966 36899 3972 36933
rect 4006 36899 4012 36933
rect 3966 36860 4012 36899
rect 3966 36826 3972 36860
rect 4006 36826 4012 36860
rect 3966 36787 4012 36826
rect 3966 36753 3972 36787
rect 4006 36753 4012 36787
rect 3966 36714 4012 36753
rect 3966 36680 3972 36714
rect 4006 36680 4012 36714
rect 3966 36641 4012 36680
rect 3966 36607 3972 36641
rect 4006 36607 4012 36641
rect 3966 36568 4012 36607
rect 3966 36534 3972 36568
rect 4006 36534 4012 36568
rect 3966 36495 4012 36534
rect 3966 36461 3972 36495
rect 4006 36461 4012 36495
rect 3966 36422 4012 36461
rect 3966 36388 3972 36422
rect 4006 36388 4012 36422
rect 3966 36349 4012 36388
rect 3966 36315 3972 36349
rect 4006 36315 4012 36349
rect 3966 36276 4012 36315
rect 3966 36242 3972 36276
rect 4006 36242 4012 36276
rect 3966 36203 4012 36242
rect 3966 36169 3972 36203
rect 4006 36169 4012 36203
rect 3966 36130 4012 36169
rect 3966 36096 3972 36130
rect 4006 36096 4012 36130
rect 3966 36057 4012 36096
rect 3966 36023 3972 36057
rect 4006 36023 4012 36057
rect 3966 35984 4012 36023
rect 3966 35950 3972 35984
rect 4006 35950 4012 35984
rect 3966 35911 4012 35950
rect 3966 35877 3972 35911
rect 4006 35877 4012 35911
rect 3966 35838 4012 35877
rect 3966 35804 3972 35838
rect 4006 35804 4012 35838
rect 3966 35765 4012 35804
rect 3966 35731 3972 35765
rect 4006 35731 4012 35765
rect 3966 35692 4012 35731
rect 3966 35658 3972 35692
rect 4006 35658 4012 35692
rect 3966 35619 4012 35658
rect 3966 35585 3972 35619
rect 4006 35585 4012 35619
rect 3966 35546 4012 35585
rect 3966 35512 3972 35546
rect 4006 35512 4012 35546
rect 3966 35473 4012 35512
rect 3966 35439 3972 35473
rect 4006 35439 4012 35473
rect 3966 35400 4012 35439
rect 3966 35366 3972 35400
rect 4006 35366 4012 35400
rect 3966 35327 4012 35366
rect 3966 35293 3972 35327
rect 4006 35293 4012 35327
rect 3966 35254 4012 35293
rect 3966 35220 3972 35254
rect 4006 35220 4012 35254
rect 3966 35181 4012 35220
rect 3966 35147 3972 35181
rect 4006 35147 4012 35181
rect 3966 35109 4012 35147
rect 3966 35075 3972 35109
rect 4006 35075 4012 35109
rect 3966 35037 4012 35075
rect 3966 35003 3972 35037
rect 4006 35003 4012 35037
rect 3966 34965 4012 35003
rect 3966 34931 3972 34965
rect 4006 34931 4012 34965
rect 3966 34893 4012 34931
rect 3966 34859 3972 34893
rect 4006 34859 4012 34893
rect 3966 34821 4012 34859
rect 3966 34787 3972 34821
rect 4006 34787 4012 34821
rect 3966 34749 4012 34787
rect 3966 34715 3972 34749
rect 4006 34715 4012 34749
rect 3966 34677 4012 34715
rect 3966 34643 3972 34677
rect 4006 34643 4012 34677
rect 3966 34605 4012 34643
rect 3966 34571 3972 34605
rect 4006 34571 4012 34605
rect 3966 34533 4012 34571
rect 3966 34499 3972 34533
rect 4006 34499 4012 34533
rect 3966 34461 4012 34499
rect 3966 34427 3972 34461
rect 4006 34427 4012 34461
rect 3966 34389 4012 34427
rect 3966 34355 3972 34389
rect 4006 34355 4012 34389
rect 3966 34317 4012 34355
rect 3966 34283 3972 34317
rect 4006 34283 4012 34317
rect 3966 34245 4012 34283
rect 3966 34211 3972 34245
rect 4006 34211 4012 34245
rect 3966 34173 4012 34211
rect 3966 34139 3972 34173
rect 4006 34139 4012 34173
rect 3966 34101 4012 34139
rect 3966 34067 3972 34101
rect 4006 34067 4012 34101
rect 3966 34029 4012 34067
rect 3966 33995 3972 34029
rect 4006 33995 4012 34029
rect 3966 33957 4012 33995
rect 3966 33923 3972 33957
rect 4006 33923 4012 33957
rect 3966 33885 4012 33923
rect 3966 33851 3972 33885
rect 4006 33851 4012 33885
rect 3966 33813 4012 33851
rect 3966 33779 3972 33813
rect 4006 33779 4012 33813
rect 3966 33741 4012 33779
rect 3966 33707 3972 33741
rect 4006 33707 4012 33741
rect 3966 33669 4012 33707
rect 3966 33635 3972 33669
rect 4006 33635 4012 33669
rect 3966 33597 4012 33635
rect 3966 33563 3972 33597
rect 4006 33563 4012 33597
rect 3966 33525 4012 33563
rect 3966 33491 3972 33525
rect 4006 33491 4012 33525
rect 3966 33453 4012 33491
rect 3966 33419 3972 33453
rect 4006 33419 4012 33453
rect 3966 33381 4012 33419
rect 3966 33347 3972 33381
rect 4006 33347 4012 33381
rect 3966 33309 4012 33347
rect 3966 33275 3972 33309
rect 4006 33275 4012 33309
rect 3966 33237 4012 33275
rect 3966 33203 3972 33237
rect 4006 33203 4012 33237
rect 3966 33165 4012 33203
rect 3966 33131 3972 33165
rect 4006 33131 4012 33165
rect 3966 33093 4012 33131
rect 3966 33059 3972 33093
rect 4006 33059 4012 33093
rect 3966 33021 4012 33059
rect 3966 32987 3972 33021
rect 4006 32987 4012 33021
rect 3966 32949 4012 32987
rect 3966 32915 3972 32949
rect 4006 32915 4012 32949
rect 3966 32877 4012 32915
rect 3966 32843 3972 32877
rect 4006 32843 4012 32877
rect 3966 32805 4012 32843
rect 3966 32771 3972 32805
rect 4006 32771 4012 32805
rect 3966 32733 4012 32771
rect 3966 32699 3972 32733
rect 4006 32699 4012 32733
rect 3966 32661 4012 32699
rect 3966 32627 3972 32661
rect 4006 32627 4012 32661
rect 3966 32589 4012 32627
rect 3966 32555 3972 32589
rect 4006 32555 4012 32589
rect 3966 32517 4012 32555
rect 3966 32483 3972 32517
rect 4006 32483 4012 32517
rect 3966 32445 4012 32483
rect 3966 32411 3972 32445
rect 4006 32411 4012 32445
rect 3966 32373 4012 32411
rect 3966 32339 3972 32373
rect 4006 32339 4012 32373
rect 3966 32301 4012 32339
rect 3966 32267 3972 32301
rect 4006 32267 4012 32301
rect 3966 32229 4012 32267
rect 3966 32195 3972 32229
rect 4006 32195 4012 32229
rect 3966 32157 4012 32195
rect 3966 32123 3972 32157
rect 4006 32123 4012 32157
rect 3966 32085 4012 32123
rect 3966 32051 3972 32085
rect 4006 32051 4012 32085
rect 3966 32013 4012 32051
rect 3966 31979 3972 32013
rect 4006 31979 4012 32013
rect 3966 31941 4012 31979
rect 3966 31907 3972 31941
rect 4006 31907 4012 31941
rect 3966 31869 4012 31907
rect 3966 31835 3972 31869
rect 4006 31835 4012 31869
rect 3966 31797 4012 31835
rect 3966 31763 3972 31797
rect 4006 31763 4012 31797
rect 3966 31725 4012 31763
rect 3966 31691 3972 31725
rect 4006 31691 4012 31725
rect 3966 31653 4012 31691
rect 3966 31619 3972 31653
rect 4006 31619 4012 31653
rect 3966 31581 4012 31619
rect 3966 31547 3972 31581
rect 4006 31547 4012 31581
rect 3966 31509 4012 31547
rect 3966 31475 3972 31509
rect 4006 31475 4012 31509
rect 3966 31437 4012 31475
rect 3966 31403 3972 31437
rect 4006 31403 4012 31437
rect 3966 31365 4012 31403
rect 3966 31331 3972 31365
rect 4006 31331 4012 31365
rect 3966 31293 4012 31331
rect 3966 31259 3972 31293
rect 4006 31259 4012 31293
rect 3966 31221 4012 31259
rect 3966 31187 3972 31221
rect 4006 31187 4012 31221
rect 3966 31149 4012 31187
rect 3966 31115 3972 31149
rect 4006 31115 4012 31149
rect 3966 31077 4012 31115
rect 3966 31043 3972 31077
rect 4006 31043 4012 31077
rect 3966 31005 4012 31043
rect 3966 30971 3972 31005
rect 4006 30971 4012 31005
rect 3966 30933 4012 30971
rect 3966 30899 3972 30933
rect 4006 30899 4012 30933
rect 3966 30861 4012 30899
rect 3966 30827 3972 30861
rect 4006 30827 4012 30861
rect 3966 30789 4012 30827
rect 3966 30755 3972 30789
rect 4006 30755 4012 30789
rect 3966 30717 4012 30755
rect 3966 30683 3972 30717
rect 4006 30683 4012 30717
rect 3966 30645 4012 30683
rect 3966 30611 3972 30645
rect 4006 30611 4012 30645
rect 3966 30573 4012 30611
rect 3966 30539 3972 30573
rect 4006 30539 4012 30573
rect 3966 30501 4012 30539
rect 3966 30467 3972 30501
rect 4006 30467 4012 30501
rect 3966 30429 4012 30467
rect 3966 30395 3972 30429
rect 4006 30395 4012 30429
rect 3966 30357 4012 30395
rect 3966 30323 3972 30357
rect 4006 30323 4012 30357
rect 3966 30285 4012 30323
rect 3966 30251 3972 30285
rect 4006 30251 4012 30285
rect 3966 30213 4012 30251
rect 3966 30179 3972 30213
rect 4006 30179 4012 30213
rect 3966 30141 4012 30179
rect 3966 30107 3972 30141
rect 4006 30107 4012 30141
rect 3966 30069 4012 30107
rect 3966 30035 3972 30069
rect 4006 30035 4012 30069
rect 3966 29997 4012 30035
rect 3966 29963 3972 29997
rect 4006 29963 4012 29997
rect 3966 29925 4012 29963
rect 3966 29891 3972 29925
rect 4006 29891 4012 29925
rect 3966 29853 4012 29891
rect 3966 29819 3972 29853
rect 4006 29819 4012 29853
rect 3966 29781 4012 29819
rect 3966 29747 3972 29781
rect 4006 29747 4012 29781
rect 3966 29709 4012 29747
rect 3966 29675 3972 29709
rect 4006 29675 4012 29709
rect 3966 29637 4012 29675
rect 3966 29603 3972 29637
rect 4006 29603 4012 29637
rect 3966 29565 4012 29603
rect 3966 29531 3972 29565
rect 4006 29531 4012 29565
rect 3966 29493 4012 29531
rect 3966 29459 3972 29493
rect 4006 29459 4012 29493
rect 3966 29421 4012 29459
rect 3966 29387 3972 29421
rect 4006 29387 4012 29421
rect 3966 29349 4012 29387
rect 3966 29315 3972 29349
rect 4006 29315 4012 29349
rect 3966 29277 4012 29315
rect 3966 29243 3972 29277
rect 4006 29243 4012 29277
rect 3966 29205 4012 29243
rect 3966 29171 3972 29205
rect 4006 29171 4012 29205
rect 3966 29133 4012 29171
rect 3966 29099 3972 29133
rect 4006 29099 4012 29133
rect 3966 29061 4012 29099
rect 3966 29027 3972 29061
rect 4006 29027 4012 29061
rect 3966 28989 4012 29027
rect 3966 28955 3972 28989
rect 4006 28955 4012 28989
rect 3966 28917 4012 28955
rect 3966 28883 3972 28917
rect 4006 28883 4012 28917
rect 3966 28845 4012 28883
rect 3966 28811 3972 28845
rect 4006 28811 4012 28845
rect 3966 28773 4012 28811
rect 3966 28739 3972 28773
rect 4006 28739 4012 28773
rect 3966 28701 4012 28739
rect 3966 28667 3972 28701
rect 4006 28667 4012 28701
rect 3966 28629 4012 28667
rect 3966 28595 3972 28629
rect 4006 28595 4012 28629
rect 3966 28557 4012 28595
rect 3966 28523 3972 28557
rect 4006 28523 4012 28557
rect 3966 28485 4012 28523
rect 3966 28451 3972 28485
rect 4006 28451 4012 28485
rect 3966 28413 4012 28451
rect 3966 28379 3972 28413
rect 4006 28379 4012 28413
rect 3966 28341 4012 28379
rect 3966 28307 3972 28341
rect 4006 28307 4012 28341
rect 3966 28269 4012 28307
rect 3966 28235 3972 28269
rect 4006 28235 4012 28269
rect 3966 28197 4012 28235
rect 3966 28163 3972 28197
rect 4006 28163 4012 28197
rect 3966 28125 4012 28163
rect 3966 28091 3972 28125
rect 4006 28091 4012 28125
rect 3966 28053 4012 28091
rect 3966 28019 3972 28053
rect 4006 28019 4012 28053
rect 3966 27981 4012 28019
rect 3966 27947 3972 27981
rect 4006 27947 4012 27981
rect 3966 27909 4012 27947
rect 3966 27875 3972 27909
rect 4006 27875 4012 27909
rect 3966 27837 4012 27875
rect 3966 27803 3972 27837
rect 4006 27803 4012 27837
rect 3966 27765 4012 27803
rect 3966 27731 3972 27765
rect 4006 27731 4012 27765
rect 3966 27693 4012 27731
rect 3966 27659 3972 27693
rect 4006 27659 4012 27693
rect 3966 27621 4012 27659
rect 3966 27587 3972 27621
rect 4006 27587 4012 27621
rect 3966 27549 4012 27587
rect 3966 27515 3972 27549
rect 4006 27515 4012 27549
rect 3966 27477 4012 27515
rect 3966 27443 3972 27477
rect 4006 27443 4012 27477
rect 3966 27405 4012 27443
rect 3966 27371 3972 27405
rect 4006 27371 4012 27405
rect 3966 27333 4012 27371
rect 3966 27299 3972 27333
rect 4006 27299 4012 27333
rect 3966 27261 4012 27299
rect 3966 27227 3972 27261
rect 4006 27227 4012 27261
rect 3966 27189 4012 27227
rect 3966 27155 3972 27189
rect 4006 27155 4012 27189
rect 3966 27117 4012 27155
rect 3966 27083 3972 27117
rect 4006 27083 4012 27117
rect 3966 27045 4012 27083
rect 3966 27011 3972 27045
rect 4006 27011 4012 27045
rect 3966 26973 4012 27011
rect 3966 26939 3972 26973
rect 4006 26939 4012 26973
rect 3966 26901 4012 26939
rect 3966 26867 3972 26901
rect 4006 26867 4012 26901
rect 3966 26829 4012 26867
rect 3966 26795 3972 26829
rect 4006 26795 4012 26829
rect 3966 26757 4012 26795
rect 3966 26723 3972 26757
rect 4006 26723 4012 26757
rect 3966 26685 4012 26723
rect 3966 26651 3972 26685
rect 4006 26651 4012 26685
rect 3966 26613 4012 26651
rect 3966 26579 3972 26613
rect 4006 26579 4012 26613
rect 3966 26541 4012 26579
rect 3966 26507 3972 26541
rect 4006 26507 4012 26541
rect 3966 26469 4012 26507
rect 3966 26435 3972 26469
rect 4006 26435 4012 26469
rect 3966 26397 4012 26435
rect 3966 26363 3972 26397
rect 4006 26363 4012 26397
rect 3966 26325 4012 26363
rect 3966 26291 3972 26325
rect 4006 26291 4012 26325
rect 3966 26253 4012 26291
rect 3966 26219 3972 26253
rect 4006 26219 4012 26253
rect 3966 26181 4012 26219
rect 3966 26147 3972 26181
rect 4006 26147 4012 26181
rect 3966 26109 4012 26147
rect 3966 26075 3972 26109
rect 4006 26075 4012 26109
rect 3966 26037 4012 26075
rect 3966 26003 3972 26037
rect 4006 26003 4012 26037
rect 3966 25965 4012 26003
rect 3966 25931 3972 25965
rect 4006 25931 4012 25965
rect 3966 25893 4012 25931
rect 3966 25859 3972 25893
rect 4006 25859 4012 25893
rect 3966 25821 4012 25859
rect 3966 25787 3972 25821
rect 4006 25787 4012 25821
rect 3966 25749 4012 25787
rect 3966 25715 3972 25749
rect 4006 25715 4012 25749
rect 3966 25677 4012 25715
rect 3966 25643 3972 25677
rect 4006 25643 4012 25677
rect 3966 25605 4012 25643
rect 3966 25571 3972 25605
rect 4006 25571 4012 25605
rect 3966 25533 4012 25571
rect 3966 25499 3972 25533
rect 4006 25499 4012 25533
rect 3966 25461 4012 25499
rect 3966 25427 3972 25461
rect 4006 25427 4012 25461
rect 3966 25389 4012 25427
rect 3966 25355 3972 25389
rect 4006 25355 4012 25389
rect 3966 25317 4012 25355
rect 3966 25283 3972 25317
rect 4006 25283 4012 25317
rect 3966 25245 4012 25283
rect 3966 25211 3972 25245
rect 4006 25211 4012 25245
rect 3966 25173 4012 25211
rect 3966 25139 3972 25173
rect 4006 25139 4012 25173
rect 3966 25101 4012 25139
rect 3966 25067 3972 25101
rect 4006 25067 4012 25101
rect 3966 25029 4012 25067
rect 3966 24995 3972 25029
rect 4006 24995 4012 25029
rect 3966 24957 4012 24995
rect 3966 24923 3972 24957
rect 4006 24923 4012 24957
rect 3966 24885 4012 24923
rect 3966 24851 3972 24885
rect 4006 24851 4012 24885
rect 3966 24813 4012 24851
rect 3966 24779 3972 24813
rect 4006 24779 4012 24813
rect 3966 24741 4012 24779
rect 3966 24707 3972 24741
rect 4006 24707 4012 24741
rect 3966 24669 4012 24707
rect 3966 24635 3972 24669
rect 4006 24635 4012 24669
rect 3966 24597 4012 24635
rect 3966 24563 3972 24597
rect 4006 24563 4012 24597
rect 3966 24525 4012 24563
rect 3966 24491 3972 24525
rect 4006 24491 4012 24525
rect 3966 24453 4012 24491
rect 3966 24419 3972 24453
rect 4006 24419 4012 24453
rect 3966 24381 4012 24419
rect 3966 24347 3972 24381
rect 4006 24347 4012 24381
rect 3966 24309 4012 24347
rect 3966 24275 3972 24309
rect 4006 24275 4012 24309
rect 3966 24237 4012 24275
rect 3966 24203 3972 24237
rect 4006 24203 4012 24237
rect 3966 24165 4012 24203
rect 3966 24131 3972 24165
rect 4006 24131 4012 24165
rect 3966 24093 4012 24131
rect 3966 24059 3972 24093
rect 4006 24059 4012 24093
rect 3966 24021 4012 24059
rect 3966 23987 3972 24021
rect 4006 23987 4012 24021
rect 3966 23949 4012 23987
rect 3966 23915 3972 23949
rect 4006 23915 4012 23949
rect 3966 23877 4012 23915
rect 3966 23843 3972 23877
rect 4006 23843 4012 23877
rect 3966 23805 4012 23843
rect 3966 23771 3972 23805
rect 4006 23771 4012 23805
rect 3966 23733 4012 23771
rect 3966 23699 3972 23733
rect 4006 23699 4012 23733
rect 3966 23661 4012 23699
rect 3966 23627 3972 23661
rect 4006 23627 4012 23661
rect 3966 23589 4012 23627
rect 3966 23555 3972 23589
rect 4006 23555 4012 23589
rect 3966 23517 4012 23555
rect 3966 23483 3972 23517
rect 4006 23483 4012 23517
rect 3966 23445 4012 23483
rect 3966 23411 3972 23445
rect 4006 23411 4012 23445
rect 3966 23373 4012 23411
rect 3966 23339 3972 23373
rect 4006 23339 4012 23373
rect 3966 23301 4012 23339
rect 3966 23267 3972 23301
rect 4006 23267 4012 23301
rect 3966 23229 4012 23267
rect 3966 23195 3972 23229
rect 4006 23195 4012 23229
rect 3966 23157 4012 23195
rect 3966 23123 3972 23157
rect 4006 23123 4012 23157
rect 3966 23085 4012 23123
rect 3966 23051 3972 23085
rect 4006 23051 4012 23085
rect 3966 23013 4012 23051
rect 3966 22979 3972 23013
rect 4006 22979 4012 23013
rect 3966 22941 4012 22979
rect 3966 22907 3972 22941
rect 4006 22907 4012 22941
rect 3966 22869 4012 22907
rect 3966 22835 3972 22869
rect 4006 22835 4012 22869
rect 3966 22797 4012 22835
rect 3966 22763 3972 22797
rect 4006 22763 4012 22797
rect 3966 22725 4012 22763
rect 3966 22691 3972 22725
rect 4006 22691 4012 22725
rect 3966 22653 4012 22691
rect 3966 22619 3972 22653
rect 4006 22619 4012 22653
rect 3966 22581 4012 22619
rect 3966 22547 3972 22581
rect 4006 22547 4012 22581
rect 3966 22509 4012 22547
rect 3966 22475 3972 22509
rect 4006 22475 4012 22509
rect 3966 22437 4012 22475
rect 3966 22403 3972 22437
rect 4006 22403 4012 22437
rect 3966 22365 4012 22403
rect 3966 22331 3972 22365
rect 4006 22331 4012 22365
rect 3966 22293 4012 22331
rect 3966 22259 3972 22293
rect 4006 22259 4012 22293
rect 3966 22221 4012 22259
rect 3966 22187 3972 22221
rect 4006 22187 4012 22221
rect 3966 22149 4012 22187
rect 3966 22115 3972 22149
rect 4006 22115 4012 22149
rect 3966 22077 4012 22115
rect 3966 22043 3972 22077
rect 4006 22043 4012 22077
rect 3966 22005 4012 22043
rect 3966 21971 3972 22005
rect 4006 21971 4012 22005
rect 3966 21933 4012 21971
rect 3966 21899 3972 21933
rect 4006 21899 4012 21933
rect 3966 21861 4012 21899
rect 3966 21827 3972 21861
rect 4006 21827 4012 21861
rect 3966 21789 4012 21827
rect 3966 21755 3972 21789
rect 4006 21755 4012 21789
rect 3966 21717 4012 21755
rect 3966 21683 3972 21717
rect 4006 21683 4012 21717
rect 3966 21645 4012 21683
rect 3966 21611 3972 21645
rect 4006 21611 4012 21645
rect 3966 21573 4012 21611
rect 3966 21539 3972 21573
rect 4006 21539 4012 21573
rect 3966 21501 4012 21539
rect 3966 21467 3972 21501
rect 4006 21467 4012 21501
rect 3966 21429 4012 21467
rect 3966 21395 3972 21429
rect 4006 21395 4012 21429
rect 3966 21357 4012 21395
rect 3966 21323 3972 21357
rect 4006 21323 4012 21357
rect 3966 21285 4012 21323
rect 3966 21251 3972 21285
rect 4006 21251 4012 21285
rect 3966 21213 4012 21251
rect 3966 21179 3972 21213
rect 4006 21179 4012 21213
rect 3966 21141 4012 21179
rect 3966 21107 3972 21141
rect 4006 21107 4012 21141
rect 3966 21069 4012 21107
rect 3966 21035 3972 21069
rect 4006 21035 4012 21069
rect 3966 20997 4012 21035
rect 3966 20963 3972 20997
rect 4006 20963 4012 20997
rect 3966 20925 4012 20963
rect 3966 20891 3972 20925
rect 4006 20891 4012 20925
rect 3966 20853 4012 20891
rect 3966 20819 3972 20853
rect 4006 20819 4012 20853
rect 3966 20781 4012 20819
rect 3966 20747 3972 20781
rect 4006 20747 4012 20781
rect 3966 20709 4012 20747
rect 3966 20675 3972 20709
rect 4006 20675 4012 20709
rect 3966 20637 4012 20675
rect 3966 20603 3972 20637
rect 4006 20603 4012 20637
rect 3966 20565 4012 20603
rect 3966 20531 3972 20565
rect 4006 20531 4012 20565
rect 3966 20493 4012 20531
rect 3966 20459 3972 20493
rect 4006 20459 4012 20493
rect 3966 20421 4012 20459
rect 3966 20387 3972 20421
rect 4006 20387 4012 20421
rect 3966 20349 4012 20387
rect 3966 20315 3972 20349
rect 4006 20315 4012 20349
rect 3966 20277 4012 20315
rect 3966 20243 3972 20277
rect 4006 20243 4012 20277
rect 3966 20205 4012 20243
rect 3966 20171 3972 20205
rect 4006 20171 4012 20205
rect 3966 20133 4012 20171
rect 3966 20099 3972 20133
rect 4006 20099 4012 20133
rect 3966 20061 4012 20099
rect 3966 20027 3972 20061
rect 4006 20027 4012 20061
rect 3966 19989 4012 20027
rect 3966 19955 3972 19989
rect 4006 19955 4012 19989
rect 3966 19917 4012 19955
rect 3966 19883 3972 19917
rect 4006 19883 4012 19917
rect 3966 19845 4012 19883
rect 3966 19811 3972 19845
rect 4006 19811 4012 19845
rect 3966 19773 4012 19811
rect 3966 19739 3972 19773
rect 4006 19739 4012 19773
rect 3966 19701 4012 19739
rect 3966 19667 3972 19701
rect 4006 19667 4012 19701
rect 3966 19629 4012 19667
rect 3966 19595 3972 19629
rect 4006 19595 4012 19629
rect 3966 19557 4012 19595
rect 3966 19523 3972 19557
rect 4006 19523 4012 19557
rect 3966 19485 4012 19523
rect 3966 19451 3972 19485
rect 4006 19451 4012 19485
rect 3966 19413 4012 19451
rect 3966 19379 3972 19413
rect 4006 19379 4012 19413
rect 3966 19341 4012 19379
rect 3966 19307 3972 19341
rect 4006 19307 4012 19341
rect 3966 19269 4012 19307
rect 3966 19235 3972 19269
rect 4006 19235 4012 19269
rect 3966 19197 4012 19235
rect 3966 19163 3972 19197
rect 4006 19163 4012 19197
rect 3966 19125 4012 19163
rect 3966 19091 3972 19125
rect 4006 19091 4012 19125
rect 3966 19053 4012 19091
rect 3966 19019 3972 19053
rect 4006 19019 4012 19053
rect 3966 18981 4012 19019
rect 3966 18947 3972 18981
rect 4006 18947 4012 18981
rect 3966 18909 4012 18947
rect 3966 18875 3972 18909
rect 4006 18875 4012 18909
rect 3966 18837 4012 18875
rect 3966 18803 3972 18837
rect 4006 18803 4012 18837
rect 3966 18765 4012 18803
rect 3966 18731 3972 18765
rect 4006 18731 4012 18765
rect 3966 18693 4012 18731
rect 3966 18659 3972 18693
rect 4006 18659 4012 18693
rect 3966 18621 4012 18659
rect 3966 18587 3972 18621
rect 4006 18587 4012 18621
rect 3966 18549 4012 18587
rect 3966 18515 3972 18549
rect 4006 18515 4012 18549
rect 3966 18477 4012 18515
rect 3966 18443 3972 18477
rect 4006 18443 4012 18477
rect 3966 18405 4012 18443
rect 3966 18371 3972 18405
rect 4006 18371 4012 18405
rect 3966 18333 4012 18371
rect 3966 18299 3972 18333
rect 4006 18299 4012 18333
rect 3966 18261 4012 18299
rect 3966 18227 3972 18261
rect 4006 18227 4012 18261
rect 3966 18189 4012 18227
rect 3966 18155 3972 18189
rect 4006 18155 4012 18189
rect 3966 18117 4012 18155
rect 3966 18083 3972 18117
rect 4006 18083 4012 18117
rect 3966 18045 4012 18083
rect 3966 18011 3972 18045
rect 4006 18011 4012 18045
rect 3966 17973 4012 18011
rect 3966 17939 3972 17973
rect 4006 17939 4012 17973
rect 3966 17901 4012 17939
rect 3966 17867 3972 17901
rect 4006 17867 4012 17901
rect 3966 17829 4012 17867
rect 3966 17795 3972 17829
rect 4006 17795 4012 17829
rect 3966 17757 4012 17795
rect 3966 17723 3972 17757
rect 4006 17723 4012 17757
rect 3966 17685 4012 17723
rect 3966 17651 3972 17685
rect 4006 17651 4012 17685
rect 3966 17613 4012 17651
rect 3966 17579 3972 17613
rect 4006 17579 4012 17613
rect 3966 17541 4012 17579
rect 3966 17507 3972 17541
rect 4006 17507 4012 17541
rect 3966 17469 4012 17507
rect 3966 17435 3972 17469
rect 4006 17435 4012 17469
rect 3966 17397 4012 17435
rect 3966 17363 3972 17397
rect 4006 17363 4012 17397
rect 3966 17325 4012 17363
rect 3966 17291 3972 17325
rect 4006 17291 4012 17325
rect 3966 17253 4012 17291
rect 3966 17219 3972 17253
rect 4006 17219 4012 17253
rect 3966 17181 4012 17219
rect 3966 17147 3972 17181
rect 4006 17147 4012 17181
rect 3966 17109 4012 17147
rect 3966 17075 3972 17109
rect 4006 17075 4012 17109
rect 3966 17037 4012 17075
rect 3966 17003 3972 17037
rect 4006 17003 4012 17037
rect 3966 16965 4012 17003
rect 3966 16931 3972 16965
rect 4006 16931 4012 16965
rect 3966 16893 4012 16931
rect 3966 16859 3972 16893
rect 4006 16859 4012 16893
rect 3966 16821 4012 16859
rect 3966 16787 3972 16821
rect 4006 16787 4012 16821
rect 3966 16749 4012 16787
rect 3966 16715 3972 16749
rect 4006 16715 4012 16749
rect 3966 16677 4012 16715
rect 3966 16643 3972 16677
rect 4006 16643 4012 16677
rect 3966 16605 4012 16643
rect 3966 16571 3972 16605
rect 4006 16571 4012 16605
rect 3966 16533 4012 16571
rect 3966 16499 3972 16533
rect 4006 16499 4012 16533
rect 3966 16461 4012 16499
rect 3966 16427 3972 16461
rect 4006 16427 4012 16461
rect 3966 16389 4012 16427
rect 3966 16355 3972 16389
rect 4006 16355 4012 16389
rect 3966 16317 4012 16355
rect 3966 16283 3972 16317
rect 4006 16283 4012 16317
rect 3966 16245 4012 16283
rect 3966 16211 3972 16245
rect 4006 16211 4012 16245
rect 3966 16173 4012 16211
rect 3966 16139 3972 16173
rect 4006 16139 4012 16173
rect 3966 16101 4012 16139
rect 3966 16067 3972 16101
rect 4006 16067 4012 16101
rect 3966 16029 4012 16067
rect 3966 15995 3972 16029
rect 4006 15995 4012 16029
rect 3966 15957 4012 15995
rect 3966 15923 3972 15957
rect 4006 15923 4012 15957
rect 3966 15885 4012 15923
rect 3966 15851 3972 15885
rect 4006 15851 4012 15885
rect 3966 15813 4012 15851
rect 3966 15779 3972 15813
rect 4006 15779 4012 15813
rect 3966 15741 4012 15779
rect 3966 15707 3972 15741
rect 4006 15707 4012 15741
rect 3966 15669 4012 15707
rect 3966 15635 3972 15669
rect 4006 15635 4012 15669
rect 3966 15597 4012 15635
rect 3966 15563 3972 15597
rect 4006 15563 4012 15597
rect 3966 15525 4012 15563
rect 3966 15491 3972 15525
rect 4006 15491 4012 15525
rect 3966 15453 4012 15491
rect 3966 15419 3972 15453
rect 4006 15419 4012 15453
rect 3966 15381 4012 15419
rect 3966 15347 3972 15381
rect 4006 15347 4012 15381
rect 3966 15309 4012 15347
rect 3966 15275 3972 15309
rect 4006 15275 4012 15309
rect 3966 15237 4012 15275
rect 3966 15203 3972 15237
rect 4006 15203 4012 15237
rect 3966 15165 4012 15203
rect 3966 15131 3972 15165
rect 4006 15131 4012 15165
rect 3966 15093 4012 15131
rect 3966 15059 3972 15093
rect 4006 15059 4012 15093
rect 3966 15021 4012 15059
rect 3966 14987 3972 15021
rect 4006 14987 4012 15021
rect 3966 14949 4012 14987
rect 3966 14915 3972 14949
rect 4006 14915 4012 14949
rect 3966 14877 4012 14915
rect 3966 14843 3972 14877
rect 4006 14843 4012 14877
rect 3966 14805 4012 14843
rect 3966 14771 3972 14805
rect 4006 14771 4012 14805
rect 3966 14733 4012 14771
rect 3966 14699 3972 14733
rect 4006 14699 4012 14733
rect 3966 14661 4012 14699
rect 3966 14627 3972 14661
rect 4006 14627 4012 14661
rect 3966 14589 4012 14627
rect 3966 14555 3972 14589
rect 4006 14555 4012 14589
rect 3966 14517 4012 14555
rect 3966 14483 3972 14517
rect 4006 14483 4012 14517
rect 3966 14445 4012 14483
rect 3966 14411 3972 14445
rect 4006 14411 4012 14445
rect 3966 14373 4012 14411
rect 3966 14339 3972 14373
rect 4006 14339 4012 14373
rect 3966 14301 4012 14339
rect 3966 14267 3972 14301
rect 4006 14267 4012 14301
rect 3966 14229 4012 14267
rect 3966 14195 3972 14229
rect 4006 14195 4012 14229
rect 3966 14157 4012 14195
rect 3966 14123 3972 14157
rect 4006 14123 4012 14157
rect 3966 14085 4012 14123
rect 3966 14051 3972 14085
rect 4006 14051 4012 14085
rect 3966 14013 4012 14051
rect 3966 13979 3972 14013
rect 4006 13979 4012 14013
rect 3966 13941 4012 13979
rect 3966 13907 3972 13941
rect 4006 13907 4012 13941
rect 3966 13869 4012 13907
rect 3966 13835 3972 13869
rect 4006 13835 4012 13869
rect 3966 13797 4012 13835
rect 3966 13763 3972 13797
rect 4006 13763 4012 13797
rect 3966 13725 4012 13763
rect 3966 13691 3972 13725
rect 4006 13691 4012 13725
rect 3966 13653 4012 13691
rect 3966 13619 3972 13653
rect 4006 13619 4012 13653
rect 3966 13581 4012 13619
rect 3966 13547 3972 13581
rect 4006 13547 4012 13581
rect 3966 13509 4012 13547
rect 3966 13475 3972 13509
rect 4006 13475 4012 13509
rect 3966 13437 4012 13475
rect 3966 13403 3972 13437
rect 4006 13403 4012 13437
rect 3966 13365 4012 13403
rect 3966 13331 3972 13365
rect 4006 13331 4012 13365
rect 3966 13293 4012 13331
rect 3966 13259 3972 13293
rect 4006 13259 4012 13293
rect 3966 13221 4012 13259
rect 3966 13187 3972 13221
rect 4006 13187 4012 13221
rect 3966 13149 4012 13187
rect 3966 13115 3972 13149
rect 4006 13115 4012 13149
rect 3966 13077 4012 13115
rect 3966 13043 3972 13077
rect 4006 13043 4012 13077
rect 3966 13005 4012 13043
rect 3966 12971 3972 13005
rect 4006 12971 4012 13005
rect 3966 12933 4012 12971
rect 3966 12899 3972 12933
rect 4006 12899 4012 12933
rect 3966 12861 4012 12899
rect 3966 12827 3972 12861
rect 4006 12827 4012 12861
rect 3966 12789 4012 12827
rect 3966 12755 3972 12789
rect 4006 12755 4012 12789
rect 3966 12717 4012 12755
rect 3966 12683 3972 12717
rect 4006 12683 4012 12717
rect 3966 12645 4012 12683
rect 3966 12611 3972 12645
rect 4006 12611 4012 12645
rect 3966 12573 4012 12611
rect 3966 12539 3972 12573
rect 4006 12539 4012 12573
rect 3966 12501 4012 12539
rect 3966 12467 3972 12501
rect 4006 12467 4012 12501
rect 3966 12429 4012 12467
rect 3966 12395 3972 12429
rect 4006 12395 4012 12429
rect 3966 12357 4012 12395
rect 3966 12323 3972 12357
rect 4006 12323 4012 12357
rect 3966 12285 4012 12323
rect 3966 12251 3972 12285
rect 4006 12251 4012 12285
rect 3966 12213 4012 12251
rect 3966 12179 3972 12213
rect 4006 12179 4012 12213
rect 3966 12141 4012 12179
rect 3966 12107 3972 12141
rect 4006 12107 4012 12141
rect 3966 12069 4012 12107
rect 3966 12035 3972 12069
rect 4006 12035 4012 12069
rect 3966 11997 4012 12035
rect 3966 11963 3972 11997
rect 4006 11963 4012 11997
rect 3966 11925 4012 11963
rect 3966 11891 3972 11925
rect 4006 11891 4012 11925
rect 3966 11853 4012 11891
rect 3966 11819 3972 11853
rect 4006 11819 4012 11853
rect 3966 11781 4012 11819
rect 3966 11747 3972 11781
rect 4006 11747 4012 11781
rect 3966 11709 4012 11747
rect 3966 11675 3972 11709
rect 4006 11675 4012 11709
rect 3966 11637 4012 11675
rect 3966 11603 3972 11637
rect 4006 11603 4012 11637
rect 3966 11565 4012 11603
rect 3966 11531 3972 11565
rect 4006 11531 4012 11565
rect 3966 11493 4012 11531
rect 3966 11459 3972 11493
rect 4006 11459 4012 11493
rect 3966 11421 4012 11459
rect 3966 11387 3972 11421
rect 4006 11387 4012 11421
rect 3966 11349 4012 11387
rect 3966 11315 3972 11349
rect 4006 11315 4012 11349
rect 3966 11277 4012 11315
rect 3966 11243 3972 11277
rect 4006 11243 4012 11277
rect 3966 11205 4012 11243
rect 3966 11171 3972 11205
rect 4006 11171 4012 11205
rect 3966 11133 4012 11171
rect 3966 11099 3972 11133
rect 4006 11099 4012 11133
rect 3966 11061 4012 11099
rect 3966 11027 3972 11061
rect 4006 11027 4012 11061
rect 3966 10989 4012 11027
rect 3966 10955 3972 10989
rect 4006 10955 4012 10989
rect 3966 10917 4012 10955
rect 3966 10883 3972 10917
rect 4006 10883 4012 10917
rect 3966 10845 4012 10883
rect 3966 10811 3972 10845
rect 4006 10811 4012 10845
rect 3966 10773 4012 10811
rect 3966 10739 3972 10773
rect 4006 10739 4012 10773
rect 3966 10701 4012 10739
rect 3966 10667 3972 10701
rect 4006 10667 4012 10701
rect 3966 10629 4012 10667
rect 3966 10595 3972 10629
rect 4006 10595 4012 10629
rect 3966 10557 4012 10595
rect 3966 10523 3972 10557
rect 4006 10523 4012 10557
rect 3966 10485 4012 10523
rect 3966 10451 3972 10485
rect 4006 10451 4012 10485
rect 3966 10413 4012 10451
rect 3966 10379 3972 10413
rect 4006 10379 4012 10413
rect 3966 10341 4012 10379
rect 3966 10307 3972 10341
rect 4006 10307 4012 10341
rect 3966 10269 4012 10307
rect 3966 10235 3972 10269
rect 4006 10235 4012 10269
rect 3966 10197 4012 10235
rect 3966 10163 3972 10197
rect 4006 10163 4012 10197
rect 3966 10125 4012 10163
rect 3966 10091 3972 10125
rect 4006 10091 4012 10125
rect 3966 10053 4012 10091
rect 3966 10019 3972 10053
rect 4006 10019 4012 10053
rect 3966 9981 4012 10019
rect 3966 9947 3972 9981
rect 4006 9947 4012 9981
rect 3966 9909 4012 9947
rect 3966 9875 3972 9909
rect 4006 9875 4012 9909
rect 3966 9837 4012 9875
rect 3966 9803 3972 9837
rect 4006 9803 4012 9837
rect 3966 9765 4012 9803
rect 3966 9731 3972 9765
rect 4006 9731 4012 9765
rect 3966 9693 4012 9731
rect 3966 9659 3972 9693
rect 4006 9659 4012 9693
rect 3966 9621 4012 9659
rect 3966 9587 3972 9621
rect 4006 9587 4012 9621
rect 3966 9549 4012 9587
rect 3966 9515 3972 9549
rect 4006 9515 4012 9549
rect 3966 9477 4012 9515
rect 3966 9443 3972 9477
rect 4006 9443 4012 9477
rect 3966 9405 4012 9443
rect 3966 9371 3972 9405
rect 4006 9371 4012 9405
rect 3966 9333 4012 9371
rect 3966 9299 3972 9333
rect 4006 9299 4012 9333
rect 3966 9261 4012 9299
rect 3966 9227 3972 9261
rect 4006 9227 4012 9261
rect 3966 9189 4012 9227
rect 3966 9155 3972 9189
rect 4006 9155 4012 9189
rect 3966 9117 4012 9155
rect 3966 9083 3972 9117
rect 4006 9083 4012 9117
rect 3966 9045 4012 9083
rect 3966 9011 3972 9045
rect 4006 9011 4012 9045
rect 3966 8973 4012 9011
rect 3966 8939 3972 8973
rect 4006 8939 4012 8973
rect 3966 8901 4012 8939
rect 3966 8867 3972 8901
rect 4006 8867 4012 8901
rect 3966 8829 4012 8867
rect 3966 8795 3972 8829
rect 4006 8795 4012 8829
rect 3966 8757 4012 8795
rect 3966 8723 3972 8757
rect 4006 8723 4012 8757
rect 3966 8685 4012 8723
rect 3966 8651 3972 8685
rect 4006 8651 4012 8685
rect 3966 8613 4012 8651
rect 3966 8579 3972 8613
rect 4006 8579 4012 8613
rect 3966 8541 4012 8579
rect 3966 8507 3972 8541
rect 4006 8507 4012 8541
rect 3966 8469 4012 8507
rect 3966 8435 3972 8469
rect 4006 8435 4012 8469
rect 3966 8397 4012 8435
rect 3966 8363 3972 8397
rect 4006 8363 4012 8397
rect 3966 8325 4012 8363
rect 3966 8291 3972 8325
rect 4006 8291 4012 8325
rect 3966 8253 4012 8291
rect 3966 8219 3972 8253
rect 4006 8219 4012 8253
rect 3966 8181 4012 8219
rect 3966 8147 3972 8181
rect 4006 8147 4012 8181
rect 3966 8109 4012 8147
rect 3966 8075 3972 8109
rect 4006 8075 4012 8109
rect 3966 8037 4012 8075
rect 3966 8003 3972 8037
rect 4006 8003 4012 8037
rect 3966 7965 4012 8003
rect 3966 7931 3972 7965
rect 4006 7931 4012 7965
rect 3966 7893 4012 7931
rect 3966 7859 3972 7893
rect 4006 7859 4012 7893
rect 3966 7821 4012 7859
rect 3966 7787 3972 7821
rect 4006 7787 4012 7821
rect 3966 7749 4012 7787
rect 3966 7715 3972 7749
rect 4006 7715 4012 7749
rect 3966 7677 4012 7715
rect 3966 7643 3972 7677
rect 4006 7643 4012 7677
rect 3966 7605 4012 7643
rect 3966 7571 3972 7605
rect 4006 7571 4012 7605
rect 3966 7533 4012 7571
rect 3966 7499 3972 7533
rect 4006 7499 4012 7533
rect 3966 7461 4012 7499
rect 3966 7427 3972 7461
rect 4006 7427 4012 7461
rect 3966 7389 4012 7427
rect 3966 7355 3972 7389
rect 4006 7355 4012 7389
rect 3966 7317 4012 7355
rect 3966 7283 3972 7317
rect 4006 7283 4012 7317
rect 3966 7245 4012 7283
rect 3966 7211 3972 7245
rect 4006 7211 4012 7245
rect 3966 7173 4012 7211
rect 3966 7139 3972 7173
rect 4006 7139 4012 7173
rect 3966 7101 4012 7139
rect 3966 7067 3972 7101
rect 4006 7067 4012 7101
rect 3966 7029 4012 7067
rect 3966 6995 3972 7029
rect 4006 6995 4012 7029
rect 3966 6957 4012 6995
rect 3966 6923 3972 6957
rect 4006 6923 4012 6957
rect 3966 6885 4012 6923
rect 3966 6851 3972 6885
rect 4006 6851 4012 6885
rect 3966 6813 4012 6851
rect 3966 6779 3972 6813
rect 4006 6779 4012 6813
rect 3966 6741 4012 6779
rect 3966 6707 3972 6741
rect 4006 6707 4012 6741
rect 3966 6669 4012 6707
rect 3966 6635 3972 6669
rect 4006 6635 4012 6669
rect 3966 6597 4012 6635
rect 3966 6563 3972 6597
rect 4006 6563 4012 6597
rect 3966 6525 4012 6563
rect 3966 6491 3972 6525
rect 4006 6491 4012 6525
rect 3966 6453 4012 6491
rect 3966 6419 3972 6453
rect 4006 6419 4012 6453
rect 3966 6381 4012 6419
rect 3966 6347 3972 6381
rect 4006 6347 4012 6381
rect 3966 6309 4012 6347
rect 3966 6275 3972 6309
rect 4006 6275 4012 6309
rect 3966 6237 4012 6275
rect 3966 6203 3972 6237
rect 4006 6203 4012 6237
rect 3966 6165 4012 6203
rect 3966 6131 3972 6165
rect 4006 6131 4012 6165
rect 3966 6093 4012 6131
rect 3966 6059 3972 6093
rect 4006 6059 4012 6093
rect 3966 6021 4012 6059
rect 3966 5987 3972 6021
rect 4006 5987 4012 6021
rect 3966 5949 4012 5987
rect 3966 5915 3972 5949
rect 4006 5915 4012 5949
rect 3966 5877 4012 5915
rect 3966 5843 3972 5877
rect 4006 5843 4012 5877
rect 3966 5805 4012 5843
rect 3966 5771 3972 5805
rect 4006 5771 4012 5805
rect 3966 5733 4012 5771
rect 3966 5699 3972 5733
rect 4006 5699 4012 5733
rect 3966 5661 4012 5699
rect 3966 5627 3972 5661
rect 4006 5627 4012 5661
rect 3966 5589 4012 5627
rect 3966 5555 3972 5589
rect 4006 5555 4012 5589
rect 3966 5517 4012 5555
rect 3966 5483 3972 5517
rect 4006 5483 4012 5517
rect 3966 5445 4012 5483
rect 3966 5411 3972 5445
rect 4006 5411 4012 5445
rect 3966 5373 4012 5411
rect 3966 5339 3972 5373
rect 4006 5339 4012 5373
rect 3966 5301 4012 5339
rect 3966 5267 3972 5301
rect 4006 5267 4012 5301
rect 3966 5229 4012 5267
rect 3966 5195 3972 5229
rect 4006 5195 4012 5229
rect 3966 5157 4012 5195
rect 3966 5123 3972 5157
rect 4006 5123 4012 5157
rect 3966 5085 4012 5123
rect 3966 5051 3972 5085
rect 4006 5051 4012 5085
rect 3966 5013 4012 5051
rect 3966 4979 3972 5013
rect 4006 4979 4012 5013
rect 3966 4941 4012 4979
rect 3966 4907 3972 4941
rect 4006 4907 4012 4941
rect 3966 4869 4012 4907
rect 3966 4835 3972 4869
rect 4006 4835 4012 4869
rect 3966 4797 4012 4835
rect 3966 4763 3972 4797
rect 4006 4763 4012 4797
rect 3966 4725 4012 4763
rect 3966 4691 3972 4725
rect 4006 4691 4012 4725
rect 3966 4653 4012 4691
rect 3966 4619 3972 4653
rect 4006 4619 4012 4653
rect 3966 4581 4012 4619
rect 3966 4547 3972 4581
rect 4006 4547 4012 4581
rect 3966 4509 4012 4547
rect 3966 4475 3972 4509
rect 4006 4475 4012 4509
rect 3966 4437 4012 4475
rect 3966 4403 3972 4437
rect 4006 4403 4012 4437
rect 3966 4365 4012 4403
rect 3966 4331 3972 4365
rect 4006 4331 4012 4365
rect 3966 4293 4012 4331
rect 3966 4259 3972 4293
rect 4006 4259 4012 4293
rect 3966 4221 4012 4259
rect 3966 4187 3972 4221
rect 4006 4187 4012 4221
rect 3966 4149 4012 4187
rect 3966 4115 3972 4149
rect 4006 4115 4012 4149
rect 3966 4077 4012 4115
rect 3966 4043 3972 4077
rect 4006 4043 4012 4077
rect 3966 4005 4012 4043
rect 3966 3971 3972 4005
rect 4006 3971 4012 4005
rect 3966 3933 4012 3971
rect 3966 3899 3972 3933
rect 4006 3899 4012 3933
rect 3966 3861 4012 3899
rect 3966 3827 3972 3861
rect 4006 3827 4012 3861
rect 3966 3789 4012 3827
rect 3966 3755 3972 3789
rect 4006 3755 4012 3789
rect 3966 3717 4012 3755
rect 3966 3683 3972 3717
rect 4006 3683 4012 3717
rect 3966 3645 4012 3683
rect 3966 3611 3972 3645
rect 4006 3611 4012 3645
rect 3966 3573 4012 3611
rect 3966 3539 3972 3573
rect 4006 3539 4012 3573
rect 3966 3501 4012 3539
rect 1824 3429 1870 3467
rect 1824 3395 1830 3429
rect 1864 3395 1870 3429
rect -258 3323 -252 3357
rect -218 3323 -212 3357
rect -258 3285 -212 3323
rect -258 3251 -252 3285
rect -218 3251 -212 3285
rect 1824 3357 1870 3395
rect 2007 3492 2059 3498
rect 2007 3428 2059 3440
rect 2007 3368 2059 3376
rect 2128 3486 2292 3498
rect 2128 3452 2134 3486
rect 2168 3452 2252 3486
rect 2286 3452 2292 3486
rect 2128 3414 2292 3452
rect 2128 3380 2134 3414
rect 2168 3380 2252 3414
rect 2286 3380 2292 3414
rect 2128 3368 2292 3380
rect 2364 3486 2528 3498
rect 2364 3452 2370 3486
rect 2404 3452 2488 3486
rect 2522 3452 2528 3486
rect 2364 3414 2528 3452
rect 2364 3380 2370 3414
rect 2404 3380 2488 3414
rect 2522 3380 2528 3414
rect 2364 3368 2528 3380
rect 2600 3486 2764 3498
rect 2600 3452 2606 3486
rect 2640 3452 2724 3486
rect 2758 3452 2764 3486
rect 2600 3414 2764 3452
rect 2600 3380 2606 3414
rect 2640 3380 2724 3414
rect 2758 3380 2764 3414
rect 2600 3368 2764 3380
rect 2836 3486 3000 3498
rect 2836 3452 2842 3486
rect 2876 3452 2960 3486
rect 2994 3452 3000 3486
rect 2836 3414 3000 3452
rect 2836 3380 2842 3414
rect 2876 3380 2960 3414
rect 2994 3380 3000 3414
rect 2836 3368 3000 3380
rect 3072 3486 3236 3498
rect 3072 3452 3078 3486
rect 3112 3452 3196 3486
rect 3230 3452 3236 3486
rect 3072 3414 3236 3452
rect 3072 3380 3078 3414
rect 3112 3380 3196 3414
rect 3230 3380 3236 3414
rect 3072 3368 3236 3380
rect 3308 3486 3472 3498
rect 3308 3452 3314 3486
rect 3348 3452 3432 3486
rect 3466 3452 3472 3486
rect 3308 3414 3472 3452
rect 3308 3380 3314 3414
rect 3348 3380 3432 3414
rect 3466 3380 3472 3414
rect 3308 3368 3472 3380
rect 3544 3486 3708 3498
rect 3544 3452 3550 3486
rect 3584 3452 3668 3486
rect 3702 3452 3708 3486
rect 3544 3414 3708 3452
rect 3544 3380 3550 3414
rect 3584 3380 3668 3414
rect 3702 3380 3708 3414
rect 3544 3368 3708 3380
rect 3777 3492 3829 3498
rect 3777 3428 3829 3440
rect 3777 3368 3829 3376
rect 3966 3467 3972 3501
rect 4006 3467 4012 3501
rect 6108 38651 6114 38685
rect 6148 38651 6154 38685
rect 6108 38613 6154 38651
rect 6108 38579 6114 38613
rect 6148 38579 6154 38613
rect 6108 38541 6154 38579
rect 6108 38507 6114 38541
rect 6148 38507 6154 38541
rect 6108 38469 6154 38507
rect 6108 38435 6114 38469
rect 6148 38435 6154 38469
rect 6108 38397 6154 38435
rect 6108 38363 6114 38397
rect 6148 38363 6154 38397
rect 6108 38325 6154 38363
rect 6108 38291 6114 38325
rect 6148 38291 6154 38325
rect 6108 38253 6154 38291
rect 6108 38219 6114 38253
rect 6148 38219 6154 38253
rect 6108 38181 6154 38219
rect 6108 38147 6114 38181
rect 6148 38147 6154 38181
rect 6108 38109 6154 38147
rect 6108 38075 6114 38109
rect 6148 38075 6154 38109
rect 6108 38037 6154 38075
rect 6108 38003 6114 38037
rect 6148 38003 6154 38037
rect 6108 37965 6154 38003
rect 6108 37931 6114 37965
rect 6148 37931 6154 37965
rect 6108 37893 6154 37931
rect 6108 37859 6114 37893
rect 6148 37859 6154 37893
rect 6108 37821 6154 37859
rect 6108 37787 6114 37821
rect 6148 37787 6154 37821
rect 6108 37749 6154 37787
rect 6108 37715 6114 37749
rect 6148 37715 6154 37749
rect 6108 37677 6154 37715
rect 6108 37643 6114 37677
rect 6148 37643 6154 37677
rect 6108 37605 6154 37643
rect 6108 37571 6114 37605
rect 6148 37571 6154 37605
rect 6108 37533 6154 37571
rect 6108 37499 6114 37533
rect 6148 37499 6154 37533
rect 6108 37461 6154 37499
rect 6108 37427 6114 37461
rect 6148 37427 6154 37461
rect 6108 37389 6154 37427
rect 6108 37355 6114 37389
rect 6148 37355 6154 37389
rect 6108 37317 6154 37355
rect 6108 37283 6114 37317
rect 6148 37283 6154 37317
rect 6108 37245 6154 37283
rect 6108 37211 6114 37245
rect 6148 37211 6154 37245
rect 6108 37173 6154 37211
rect 6108 37139 6114 37173
rect 6148 37139 6154 37173
rect 6108 37101 6154 37139
rect 6108 37067 6114 37101
rect 6148 37067 6154 37101
rect 6108 37029 6154 37067
rect 6108 36995 6114 37029
rect 6148 36995 6154 37029
rect 6108 36957 6154 36995
rect 6108 36923 6114 36957
rect 6148 36923 6154 36957
rect 6108 36885 6154 36923
rect 6108 36851 6114 36885
rect 6148 36851 6154 36885
rect 6108 36813 6154 36851
rect 6108 36779 6114 36813
rect 6148 36779 6154 36813
rect 6108 36741 6154 36779
rect 6108 36707 6114 36741
rect 6148 36707 6154 36741
rect 6108 36669 6154 36707
rect 6108 36635 6114 36669
rect 6148 36635 6154 36669
rect 6108 36597 6154 36635
rect 6108 36563 6114 36597
rect 6148 36563 6154 36597
rect 6108 36525 6154 36563
rect 6108 36491 6114 36525
rect 6148 36491 6154 36525
rect 6108 36453 6154 36491
rect 6108 36419 6114 36453
rect 6148 36419 6154 36453
rect 6108 36381 6154 36419
rect 6108 36347 6114 36381
rect 6148 36347 6154 36381
rect 6108 36309 6154 36347
rect 6108 36275 6114 36309
rect 6148 36275 6154 36309
rect 6108 36237 6154 36275
rect 6108 36203 6114 36237
rect 6148 36203 6154 36237
rect 6108 36165 6154 36203
rect 6108 36131 6114 36165
rect 6148 36131 6154 36165
rect 6108 36093 6154 36131
rect 6108 36059 6114 36093
rect 6148 36059 6154 36093
rect 6108 36021 6154 36059
rect 6108 35987 6114 36021
rect 6148 35987 6154 36021
rect 6108 35949 6154 35987
rect 6108 35915 6114 35949
rect 6148 35915 6154 35949
rect 6108 35877 6154 35915
rect 6108 35843 6114 35877
rect 6148 35843 6154 35877
rect 6108 35805 6154 35843
rect 6108 35771 6114 35805
rect 6148 35771 6154 35805
rect 6108 35733 6154 35771
rect 6108 35699 6114 35733
rect 6148 35699 6154 35733
rect 6108 35661 6154 35699
rect 6108 35627 6114 35661
rect 6148 35627 6154 35661
rect 6108 35589 6154 35627
rect 6108 35555 6114 35589
rect 6148 35555 6154 35589
rect 6108 35517 6154 35555
rect 6108 35483 6114 35517
rect 6148 35483 6154 35517
rect 6108 35445 6154 35483
rect 6108 35411 6114 35445
rect 6148 35411 6154 35445
rect 6108 35373 6154 35411
rect 6108 35339 6114 35373
rect 6148 35339 6154 35373
rect 6108 35301 6154 35339
rect 6108 35267 6114 35301
rect 6148 35267 6154 35301
rect 6108 35229 6154 35267
rect 6108 35195 6114 35229
rect 6148 35195 6154 35229
rect 6108 35157 6154 35195
rect 6108 35123 6114 35157
rect 6148 35123 6154 35157
rect 6108 35085 6154 35123
rect 6108 35051 6114 35085
rect 6148 35051 6154 35085
rect 6108 35013 6154 35051
rect 6108 34979 6114 35013
rect 6148 34979 6154 35013
rect 6108 34941 6154 34979
rect 6108 34907 6114 34941
rect 6148 34907 6154 34941
rect 6108 34869 6154 34907
rect 6108 34835 6114 34869
rect 6148 34835 6154 34869
rect 6108 34797 6154 34835
rect 6108 34763 6114 34797
rect 6148 34763 6154 34797
rect 6108 34725 6154 34763
rect 6108 34691 6114 34725
rect 6148 34691 6154 34725
rect 6108 34653 6154 34691
rect 6108 34619 6114 34653
rect 6148 34619 6154 34653
rect 6108 34581 6154 34619
rect 6108 34547 6114 34581
rect 6148 34547 6154 34581
rect 6108 34509 6154 34547
rect 6108 34475 6114 34509
rect 6148 34475 6154 34509
rect 6108 34437 6154 34475
rect 6108 34403 6114 34437
rect 6148 34403 6154 34437
rect 6108 34365 6154 34403
rect 6108 34331 6114 34365
rect 6148 34331 6154 34365
rect 6108 34293 6154 34331
rect 6108 34259 6114 34293
rect 6148 34259 6154 34293
rect 6108 34221 6154 34259
rect 6108 34187 6114 34221
rect 6148 34187 6154 34221
rect 6108 34149 6154 34187
rect 6108 34115 6114 34149
rect 6148 34115 6154 34149
rect 6108 34077 6154 34115
rect 6108 34043 6114 34077
rect 6148 34043 6154 34077
rect 6108 34005 6154 34043
rect 6108 33971 6114 34005
rect 6148 33971 6154 34005
rect 6108 33933 6154 33971
rect 6108 33899 6114 33933
rect 6148 33899 6154 33933
rect 6108 33861 6154 33899
rect 6108 33827 6114 33861
rect 6148 33827 6154 33861
rect 6108 33789 6154 33827
rect 6108 33755 6114 33789
rect 6148 33755 6154 33789
rect 6108 33717 6154 33755
rect 6108 33683 6114 33717
rect 6148 33683 6154 33717
rect 6108 33645 6154 33683
rect 6108 33611 6114 33645
rect 6148 33611 6154 33645
rect 6108 33573 6154 33611
rect 6108 33539 6114 33573
rect 6148 33539 6154 33573
rect 6108 33501 6154 33539
rect 6108 33467 6114 33501
rect 6148 33467 6154 33501
rect 6108 33429 6154 33467
rect 6108 33395 6114 33429
rect 6148 33395 6154 33429
rect 6108 33357 6154 33395
rect 6108 33323 6114 33357
rect 6148 33323 6154 33357
rect 6108 33285 6154 33323
rect 6108 33251 6114 33285
rect 6148 33251 6154 33285
rect 6108 33213 6154 33251
rect 6108 33179 6114 33213
rect 6148 33179 6154 33213
rect 6108 33141 6154 33179
rect 6108 33107 6114 33141
rect 6148 33107 6154 33141
rect 6108 33069 6154 33107
rect 6108 33035 6114 33069
rect 6148 33035 6154 33069
rect 6108 32997 6154 33035
rect 6108 32963 6114 32997
rect 6148 32963 6154 32997
rect 6108 32925 6154 32963
rect 6108 32891 6114 32925
rect 6148 32891 6154 32925
rect 6108 32853 6154 32891
rect 6108 32819 6114 32853
rect 6148 32819 6154 32853
rect 6108 32781 6154 32819
rect 6108 32747 6114 32781
rect 6148 32747 6154 32781
rect 6108 32709 6154 32747
rect 6108 32675 6114 32709
rect 6148 32675 6154 32709
rect 6108 32637 6154 32675
rect 6108 32603 6114 32637
rect 6148 32603 6154 32637
rect 6108 32565 6154 32603
rect 6108 32531 6114 32565
rect 6148 32531 6154 32565
rect 6108 32493 6154 32531
rect 6108 32459 6114 32493
rect 6148 32459 6154 32493
rect 6108 32421 6154 32459
rect 6108 32387 6114 32421
rect 6148 32387 6154 32421
rect 6108 32349 6154 32387
rect 6108 32315 6114 32349
rect 6148 32315 6154 32349
rect 6108 32277 6154 32315
rect 6108 32243 6114 32277
rect 6148 32243 6154 32277
rect 6108 32205 6154 32243
rect 6108 32171 6114 32205
rect 6148 32171 6154 32205
rect 6108 32133 6154 32171
rect 6108 32099 6114 32133
rect 6148 32099 6154 32133
rect 6108 32061 6154 32099
rect 6108 32027 6114 32061
rect 6148 32027 6154 32061
rect 6108 31989 6154 32027
rect 6108 31955 6114 31989
rect 6148 31955 6154 31989
rect 6108 31917 6154 31955
rect 6108 31883 6114 31917
rect 6148 31883 6154 31917
rect 6108 31845 6154 31883
rect 6108 31811 6114 31845
rect 6148 31811 6154 31845
rect 6108 31773 6154 31811
rect 6108 31739 6114 31773
rect 6148 31739 6154 31773
rect 6108 31701 6154 31739
rect 6108 31667 6114 31701
rect 6148 31667 6154 31701
rect 6108 31629 6154 31667
rect 6108 31595 6114 31629
rect 6148 31595 6154 31629
rect 6108 31557 6154 31595
rect 6108 31523 6114 31557
rect 6148 31523 6154 31557
rect 6108 31485 6154 31523
rect 6108 31451 6114 31485
rect 6148 31451 6154 31485
rect 6108 31413 6154 31451
rect 6108 31379 6114 31413
rect 6148 31379 6154 31413
rect 6108 31341 6154 31379
rect 6108 31307 6114 31341
rect 6148 31307 6154 31341
rect 6108 31269 6154 31307
rect 6108 31235 6114 31269
rect 6148 31235 6154 31269
rect 6108 31197 6154 31235
rect 6108 31163 6114 31197
rect 6148 31163 6154 31197
rect 6108 31125 6154 31163
rect 6108 31091 6114 31125
rect 6148 31091 6154 31125
rect 6108 31053 6154 31091
rect 6108 31019 6114 31053
rect 6148 31019 6154 31053
rect 6108 30981 6154 31019
rect 6108 30947 6114 30981
rect 6148 30947 6154 30981
rect 6108 30909 6154 30947
rect 6108 30875 6114 30909
rect 6148 30875 6154 30909
rect 6108 30837 6154 30875
rect 6108 30803 6114 30837
rect 6148 30803 6154 30837
rect 6108 30765 6154 30803
rect 6108 30731 6114 30765
rect 6148 30731 6154 30765
rect 6108 30693 6154 30731
rect 6108 30659 6114 30693
rect 6148 30659 6154 30693
rect 6108 30621 6154 30659
rect 6108 30587 6114 30621
rect 6148 30587 6154 30621
rect 6108 30549 6154 30587
rect 6108 30515 6114 30549
rect 6148 30515 6154 30549
rect 6108 30477 6154 30515
rect 6108 30443 6114 30477
rect 6148 30443 6154 30477
rect 6108 30405 6154 30443
rect 6108 30371 6114 30405
rect 6148 30371 6154 30405
rect 6108 30333 6154 30371
rect 6108 30299 6114 30333
rect 6148 30299 6154 30333
rect 6108 30261 6154 30299
rect 6108 30227 6114 30261
rect 6148 30227 6154 30261
rect 6108 30189 6154 30227
rect 6108 30155 6114 30189
rect 6148 30155 6154 30189
rect 6108 30117 6154 30155
rect 6108 30083 6114 30117
rect 6148 30083 6154 30117
rect 6108 30045 6154 30083
rect 6108 30011 6114 30045
rect 6148 30011 6154 30045
rect 6108 29973 6154 30011
rect 6108 29939 6114 29973
rect 6148 29939 6154 29973
rect 6108 29901 6154 29939
rect 6108 29867 6114 29901
rect 6148 29867 6154 29901
rect 6108 29829 6154 29867
rect 6108 29795 6114 29829
rect 6148 29795 6154 29829
rect 6108 29757 6154 29795
rect 6108 29723 6114 29757
rect 6148 29723 6154 29757
rect 6108 29685 6154 29723
rect 6108 29651 6114 29685
rect 6148 29651 6154 29685
rect 6108 29613 6154 29651
rect 6108 29579 6114 29613
rect 6148 29579 6154 29613
rect 6108 29541 6154 29579
rect 6108 29507 6114 29541
rect 6148 29507 6154 29541
rect 6108 29469 6154 29507
rect 6108 29435 6114 29469
rect 6148 29435 6154 29469
rect 6108 29397 6154 29435
rect 6108 29363 6114 29397
rect 6148 29363 6154 29397
rect 6108 29325 6154 29363
rect 6108 29291 6114 29325
rect 6148 29291 6154 29325
rect 6108 29253 6154 29291
rect 6108 29219 6114 29253
rect 6148 29219 6154 29253
rect 6108 29181 6154 29219
rect 6108 29147 6114 29181
rect 6148 29147 6154 29181
rect 6108 29109 6154 29147
rect 6108 29075 6114 29109
rect 6148 29075 6154 29109
rect 6108 29037 6154 29075
rect 6108 29003 6114 29037
rect 6148 29003 6154 29037
rect 6108 28965 6154 29003
rect 6108 28931 6114 28965
rect 6148 28931 6154 28965
rect 6108 28893 6154 28931
rect 6108 28859 6114 28893
rect 6148 28859 6154 28893
rect 6108 28821 6154 28859
rect 6108 28787 6114 28821
rect 6148 28787 6154 28821
rect 6108 28749 6154 28787
rect 6108 28715 6114 28749
rect 6148 28715 6154 28749
rect 6108 28677 6154 28715
rect 6108 28643 6114 28677
rect 6148 28643 6154 28677
rect 6108 28605 6154 28643
rect 6108 28571 6114 28605
rect 6148 28571 6154 28605
rect 6108 28533 6154 28571
rect 6108 28499 6114 28533
rect 6148 28499 6154 28533
rect 6108 28461 6154 28499
rect 6108 28427 6114 28461
rect 6148 28427 6154 28461
rect 6108 28389 6154 28427
rect 6108 28355 6114 28389
rect 6148 28355 6154 28389
rect 6108 28317 6154 28355
rect 6108 28283 6114 28317
rect 6148 28283 6154 28317
rect 6108 28245 6154 28283
rect 6108 28211 6114 28245
rect 6148 28211 6154 28245
rect 6108 28173 6154 28211
rect 6108 28139 6114 28173
rect 6148 28139 6154 28173
rect 6108 28101 6154 28139
rect 6108 28067 6114 28101
rect 6148 28067 6154 28101
rect 6108 28029 6154 28067
rect 6108 27995 6114 28029
rect 6148 27995 6154 28029
rect 6108 27957 6154 27995
rect 6108 27923 6114 27957
rect 6148 27923 6154 27957
rect 6108 27885 6154 27923
rect 6108 27851 6114 27885
rect 6148 27851 6154 27885
rect 6108 27813 6154 27851
rect 6108 27779 6114 27813
rect 6148 27779 6154 27813
rect 6108 27741 6154 27779
rect 6108 27707 6114 27741
rect 6148 27707 6154 27741
rect 6108 27669 6154 27707
rect 6108 27635 6114 27669
rect 6148 27635 6154 27669
rect 6108 27597 6154 27635
rect 6108 27563 6114 27597
rect 6148 27563 6154 27597
rect 6108 27525 6154 27563
rect 6108 27491 6114 27525
rect 6148 27491 6154 27525
rect 6108 27453 6154 27491
rect 6108 27419 6114 27453
rect 6148 27419 6154 27453
rect 6108 27381 6154 27419
rect 6108 27347 6114 27381
rect 6148 27347 6154 27381
rect 6108 27309 6154 27347
rect 6108 27275 6114 27309
rect 6148 27275 6154 27309
rect 6108 27237 6154 27275
rect 6108 27203 6114 27237
rect 6148 27203 6154 27237
rect 6108 27165 6154 27203
rect 6108 27131 6114 27165
rect 6148 27131 6154 27165
rect 6108 27093 6154 27131
rect 6108 27059 6114 27093
rect 6148 27059 6154 27093
rect 6108 27021 6154 27059
rect 6108 26987 6114 27021
rect 6148 26987 6154 27021
rect 6108 26949 6154 26987
rect 6108 26915 6114 26949
rect 6148 26915 6154 26949
rect 6108 26877 6154 26915
rect 6108 26843 6114 26877
rect 6148 26843 6154 26877
rect 6108 26805 6154 26843
rect 6108 26771 6114 26805
rect 6148 26771 6154 26805
rect 6108 26733 6154 26771
rect 6108 26699 6114 26733
rect 6148 26699 6154 26733
rect 6108 26661 6154 26699
rect 6108 26627 6114 26661
rect 6148 26627 6154 26661
rect 6108 26589 6154 26627
rect 6108 26555 6114 26589
rect 6148 26555 6154 26589
rect 6108 26517 6154 26555
rect 6108 26483 6114 26517
rect 6148 26483 6154 26517
rect 6108 26445 6154 26483
rect 6108 26411 6114 26445
rect 6148 26411 6154 26445
rect 6108 26373 6154 26411
rect 6108 26339 6114 26373
rect 6148 26339 6154 26373
rect 6108 26301 6154 26339
rect 6108 26267 6114 26301
rect 6148 26267 6154 26301
rect 6108 26229 6154 26267
rect 6108 26195 6114 26229
rect 6148 26195 6154 26229
rect 6108 26157 6154 26195
rect 6108 26123 6114 26157
rect 6148 26123 6154 26157
rect 6108 26085 6154 26123
rect 6108 26051 6114 26085
rect 6148 26051 6154 26085
rect 6108 26013 6154 26051
rect 6108 25979 6114 26013
rect 6148 25979 6154 26013
rect 6108 25941 6154 25979
rect 6108 25907 6114 25941
rect 6148 25907 6154 25941
rect 6108 25869 6154 25907
rect 6108 25835 6114 25869
rect 6148 25835 6154 25869
rect 6108 25797 6154 25835
rect 6108 25763 6114 25797
rect 6148 25763 6154 25797
rect 6108 25725 6154 25763
rect 6108 25691 6114 25725
rect 6148 25691 6154 25725
rect 6108 25653 6154 25691
rect 6108 25619 6114 25653
rect 6148 25619 6154 25653
rect 6108 25581 6154 25619
rect 6108 25547 6114 25581
rect 6148 25547 6154 25581
rect 6108 25509 6154 25547
rect 6108 25475 6114 25509
rect 6148 25475 6154 25509
rect 6108 25437 6154 25475
rect 6108 25403 6114 25437
rect 6148 25403 6154 25437
rect 6108 25365 6154 25403
rect 6108 25331 6114 25365
rect 6148 25331 6154 25365
rect 6108 25293 6154 25331
rect 6108 25259 6114 25293
rect 6148 25259 6154 25293
rect 6108 25221 6154 25259
rect 6108 25187 6114 25221
rect 6148 25187 6154 25221
rect 6108 25149 6154 25187
rect 6108 25115 6114 25149
rect 6148 25115 6154 25149
rect 6108 25077 6154 25115
rect 6108 25043 6114 25077
rect 6148 25043 6154 25077
rect 6108 25005 6154 25043
rect 6108 24971 6114 25005
rect 6148 24971 6154 25005
rect 6108 24933 6154 24971
rect 6108 24899 6114 24933
rect 6148 24899 6154 24933
rect 6108 24861 6154 24899
rect 6108 24827 6114 24861
rect 6148 24827 6154 24861
rect 6108 24789 6154 24827
rect 6108 24755 6114 24789
rect 6148 24755 6154 24789
rect 6108 24717 6154 24755
rect 6108 24683 6114 24717
rect 6148 24683 6154 24717
rect 6108 24645 6154 24683
rect 6108 24611 6114 24645
rect 6148 24611 6154 24645
rect 6108 24573 6154 24611
rect 6108 24539 6114 24573
rect 6148 24539 6154 24573
rect 6108 24501 6154 24539
rect 6108 24467 6114 24501
rect 6148 24467 6154 24501
rect 6108 24429 6154 24467
rect 6108 24395 6114 24429
rect 6148 24395 6154 24429
rect 6108 24357 6154 24395
rect 6108 24323 6114 24357
rect 6148 24323 6154 24357
rect 6108 24285 6154 24323
rect 6108 24251 6114 24285
rect 6148 24251 6154 24285
rect 6108 24213 6154 24251
rect 6108 24179 6114 24213
rect 6148 24179 6154 24213
rect 6108 24141 6154 24179
rect 6108 24107 6114 24141
rect 6148 24107 6154 24141
rect 6108 24069 6154 24107
rect 6108 24035 6114 24069
rect 6148 24035 6154 24069
rect 6108 23997 6154 24035
rect 6108 23963 6114 23997
rect 6148 23963 6154 23997
rect 6108 23925 6154 23963
rect 6108 23891 6114 23925
rect 6148 23891 6154 23925
rect 6108 23853 6154 23891
rect 6108 23819 6114 23853
rect 6148 23819 6154 23853
rect 6108 23781 6154 23819
rect 6108 23747 6114 23781
rect 6148 23747 6154 23781
rect 6108 23709 6154 23747
rect 6108 23675 6114 23709
rect 6148 23675 6154 23709
rect 6108 23637 6154 23675
rect 6108 23603 6114 23637
rect 6148 23603 6154 23637
rect 6108 23565 6154 23603
rect 6108 23531 6114 23565
rect 6148 23531 6154 23565
rect 6108 23493 6154 23531
rect 6108 23459 6114 23493
rect 6148 23459 6154 23493
rect 6108 23421 6154 23459
rect 6108 23387 6114 23421
rect 6148 23387 6154 23421
rect 6108 23349 6154 23387
rect 6108 23315 6114 23349
rect 6148 23315 6154 23349
rect 6108 23277 6154 23315
rect 6108 23243 6114 23277
rect 6148 23243 6154 23277
rect 6108 23205 6154 23243
rect 6108 23171 6114 23205
rect 6148 23171 6154 23205
rect 6108 23133 6154 23171
rect 6108 23099 6114 23133
rect 6148 23099 6154 23133
rect 6108 23061 6154 23099
rect 6108 23027 6114 23061
rect 6148 23027 6154 23061
rect 6108 22989 6154 23027
rect 6108 22955 6114 22989
rect 6148 22955 6154 22989
rect 6108 22917 6154 22955
rect 6108 22883 6114 22917
rect 6148 22883 6154 22917
rect 6108 22845 6154 22883
rect 6108 22811 6114 22845
rect 6148 22811 6154 22845
rect 6108 22773 6154 22811
rect 6108 22739 6114 22773
rect 6148 22739 6154 22773
rect 6108 22701 6154 22739
rect 6108 22667 6114 22701
rect 6148 22667 6154 22701
rect 6108 22629 6154 22667
rect 6108 22595 6114 22629
rect 6148 22595 6154 22629
rect 6108 22557 6154 22595
rect 6108 22523 6114 22557
rect 6148 22523 6154 22557
rect 6108 22485 6154 22523
rect 6108 22451 6114 22485
rect 6148 22451 6154 22485
rect 6108 22413 6154 22451
rect 6108 22379 6114 22413
rect 6148 22379 6154 22413
rect 6108 22341 6154 22379
rect 6108 22307 6114 22341
rect 6148 22307 6154 22341
rect 6108 22269 6154 22307
rect 6108 22235 6114 22269
rect 6148 22235 6154 22269
rect 6108 22197 6154 22235
rect 6108 22163 6114 22197
rect 6148 22163 6154 22197
rect 6108 22125 6154 22163
rect 6108 22091 6114 22125
rect 6148 22091 6154 22125
rect 6108 22053 6154 22091
rect 6108 22019 6114 22053
rect 6148 22019 6154 22053
rect 6108 21981 6154 22019
rect 6108 21947 6114 21981
rect 6148 21947 6154 21981
rect 6108 21909 6154 21947
rect 6108 21875 6114 21909
rect 6148 21875 6154 21909
rect 6108 21837 6154 21875
rect 6108 21803 6114 21837
rect 6148 21803 6154 21837
rect 6108 21765 6154 21803
rect 6108 21731 6114 21765
rect 6148 21731 6154 21765
rect 6108 21693 6154 21731
rect 6108 21659 6114 21693
rect 6148 21659 6154 21693
rect 6108 21621 6154 21659
rect 6108 21587 6114 21621
rect 6148 21587 6154 21621
rect 6108 21549 6154 21587
rect 6108 21515 6114 21549
rect 6148 21515 6154 21549
rect 6108 21477 6154 21515
rect 6108 21443 6114 21477
rect 6148 21443 6154 21477
rect 6108 21405 6154 21443
rect 6108 21371 6114 21405
rect 6148 21371 6154 21405
rect 6108 21333 6154 21371
rect 6108 21299 6114 21333
rect 6148 21299 6154 21333
rect 6108 21261 6154 21299
rect 6108 21227 6114 21261
rect 6148 21227 6154 21261
rect 6108 21189 6154 21227
rect 6108 21155 6114 21189
rect 6148 21155 6154 21189
rect 6108 21117 6154 21155
rect 6108 21083 6114 21117
rect 6148 21083 6154 21117
rect 6108 21045 6154 21083
rect 6108 21011 6114 21045
rect 6148 21011 6154 21045
rect 6108 20973 6154 21011
rect 6108 20939 6114 20973
rect 6148 20939 6154 20973
rect 6108 20901 6154 20939
rect 6108 20867 6114 20901
rect 6148 20867 6154 20901
rect 6108 20829 6154 20867
rect 6108 20795 6114 20829
rect 6148 20795 6154 20829
rect 6108 20757 6154 20795
rect 6108 20723 6114 20757
rect 6148 20723 6154 20757
rect 6108 20685 6154 20723
rect 6108 20651 6114 20685
rect 6148 20651 6154 20685
rect 6108 20613 6154 20651
rect 6108 20579 6114 20613
rect 6148 20579 6154 20613
rect 6108 20541 6154 20579
rect 6108 20507 6114 20541
rect 6148 20507 6154 20541
rect 6108 20469 6154 20507
rect 6108 20435 6114 20469
rect 6148 20435 6154 20469
rect 6108 20397 6154 20435
rect 6108 20363 6114 20397
rect 6148 20363 6154 20397
rect 6108 20325 6154 20363
rect 6108 20291 6114 20325
rect 6148 20291 6154 20325
rect 6108 20253 6154 20291
rect 6108 20219 6114 20253
rect 6148 20219 6154 20253
rect 6108 20181 6154 20219
rect 6108 20147 6114 20181
rect 6148 20147 6154 20181
rect 6108 20109 6154 20147
rect 6108 20075 6114 20109
rect 6148 20075 6154 20109
rect 6108 20037 6154 20075
rect 6108 20003 6114 20037
rect 6148 20003 6154 20037
rect 6108 19965 6154 20003
rect 6108 19931 6114 19965
rect 6148 19931 6154 19965
rect 6108 19893 6154 19931
rect 6108 19859 6114 19893
rect 6148 19859 6154 19893
rect 6108 19821 6154 19859
rect 6108 19787 6114 19821
rect 6148 19787 6154 19821
rect 6108 19749 6154 19787
rect 6108 19715 6114 19749
rect 6148 19715 6154 19749
rect 6108 19677 6154 19715
rect 6108 19643 6114 19677
rect 6148 19643 6154 19677
rect 6108 19605 6154 19643
rect 6108 19571 6114 19605
rect 6148 19571 6154 19605
rect 6108 19533 6154 19571
rect 6108 19499 6114 19533
rect 6148 19499 6154 19533
rect 6108 19461 6154 19499
rect 6108 19427 6114 19461
rect 6148 19427 6154 19461
rect 6108 19389 6154 19427
rect 6108 19355 6114 19389
rect 6148 19355 6154 19389
rect 6108 19317 6154 19355
rect 6108 19283 6114 19317
rect 6148 19283 6154 19317
rect 6108 19245 6154 19283
rect 6108 19211 6114 19245
rect 6148 19211 6154 19245
rect 6108 19173 6154 19211
rect 6108 19139 6114 19173
rect 6148 19139 6154 19173
rect 6108 19101 6154 19139
rect 6108 19067 6114 19101
rect 6148 19067 6154 19101
rect 6108 19029 6154 19067
rect 6108 18995 6114 19029
rect 6148 18995 6154 19029
rect 6108 18957 6154 18995
rect 6108 18923 6114 18957
rect 6148 18923 6154 18957
rect 6108 18885 6154 18923
rect 6108 18851 6114 18885
rect 6148 18851 6154 18885
rect 6108 18813 6154 18851
rect 6108 18779 6114 18813
rect 6148 18779 6154 18813
rect 6108 18741 6154 18779
rect 6108 18707 6114 18741
rect 6148 18707 6154 18741
rect 6108 18669 6154 18707
rect 6108 18635 6114 18669
rect 6148 18635 6154 18669
rect 6108 18597 6154 18635
rect 6108 18563 6114 18597
rect 6148 18563 6154 18597
rect 6108 18525 6154 18563
rect 6108 18491 6114 18525
rect 6148 18491 6154 18525
rect 6108 18453 6154 18491
rect 6108 18419 6114 18453
rect 6148 18419 6154 18453
rect 6108 18381 6154 18419
rect 6108 18347 6114 18381
rect 6148 18347 6154 18381
rect 6108 18309 6154 18347
rect 6108 18275 6114 18309
rect 6148 18275 6154 18309
rect 6108 18237 6154 18275
rect 6108 18203 6114 18237
rect 6148 18203 6154 18237
rect 6108 18165 6154 18203
rect 6108 18131 6114 18165
rect 6148 18131 6154 18165
rect 6108 18093 6154 18131
rect 6108 18059 6114 18093
rect 6148 18059 6154 18093
rect 6108 18021 6154 18059
rect 6108 17987 6114 18021
rect 6148 17987 6154 18021
rect 6108 17949 6154 17987
rect 6108 17915 6114 17949
rect 6148 17915 6154 17949
rect 6108 17877 6154 17915
rect 6108 17843 6114 17877
rect 6148 17843 6154 17877
rect 6108 17805 6154 17843
rect 6108 17771 6114 17805
rect 6148 17771 6154 17805
rect 6108 17733 6154 17771
rect 6108 17699 6114 17733
rect 6148 17699 6154 17733
rect 6108 17661 6154 17699
rect 6108 17627 6114 17661
rect 6148 17627 6154 17661
rect 6108 17589 6154 17627
rect 6108 17555 6114 17589
rect 6148 17555 6154 17589
rect 6108 17517 6154 17555
rect 6108 17483 6114 17517
rect 6148 17483 6154 17517
rect 6108 17445 6154 17483
rect 6108 17411 6114 17445
rect 6148 17411 6154 17445
rect 6108 17373 6154 17411
rect 6108 17339 6114 17373
rect 6148 17339 6154 17373
rect 6108 17301 6154 17339
rect 6108 17267 6114 17301
rect 6148 17267 6154 17301
rect 6108 17229 6154 17267
rect 6108 17195 6114 17229
rect 6148 17195 6154 17229
rect 6108 17157 6154 17195
rect 6108 17123 6114 17157
rect 6148 17123 6154 17157
rect 6108 17085 6154 17123
rect 6108 17051 6114 17085
rect 6148 17051 6154 17085
rect 6108 17013 6154 17051
rect 6108 16979 6114 17013
rect 6148 16979 6154 17013
rect 6108 16941 6154 16979
rect 6108 16907 6114 16941
rect 6148 16907 6154 16941
rect 6108 16869 6154 16907
rect 6108 16835 6114 16869
rect 6148 16835 6154 16869
rect 6108 16797 6154 16835
rect 6108 16763 6114 16797
rect 6148 16763 6154 16797
rect 6108 16725 6154 16763
rect 6108 16691 6114 16725
rect 6148 16691 6154 16725
rect 6108 16653 6154 16691
rect 6108 16619 6114 16653
rect 6148 16619 6154 16653
rect 6108 16581 6154 16619
rect 6108 16547 6114 16581
rect 6148 16547 6154 16581
rect 6108 16509 6154 16547
rect 6108 16475 6114 16509
rect 6148 16475 6154 16509
rect 6108 16437 6154 16475
rect 6108 16403 6114 16437
rect 6148 16403 6154 16437
rect 6108 16365 6154 16403
rect 6108 16331 6114 16365
rect 6148 16331 6154 16365
rect 6108 16293 6154 16331
rect 6108 16259 6114 16293
rect 6148 16259 6154 16293
rect 6108 16221 6154 16259
rect 6108 16187 6114 16221
rect 6148 16187 6154 16221
rect 6108 16149 6154 16187
rect 6108 16115 6114 16149
rect 6148 16115 6154 16149
rect 6108 16077 6154 16115
rect 6108 16043 6114 16077
rect 6148 16043 6154 16077
rect 6108 16005 6154 16043
rect 6108 15971 6114 16005
rect 6148 15971 6154 16005
rect 6108 15933 6154 15971
rect 6108 15899 6114 15933
rect 6148 15899 6154 15933
rect 6108 15861 6154 15899
rect 6108 15827 6114 15861
rect 6148 15827 6154 15861
rect 6108 15789 6154 15827
rect 6108 15755 6114 15789
rect 6148 15755 6154 15789
rect 6108 15717 6154 15755
rect 6108 15683 6114 15717
rect 6148 15683 6154 15717
rect 6108 15645 6154 15683
rect 6108 15611 6114 15645
rect 6148 15611 6154 15645
rect 6108 15573 6154 15611
rect 6108 15539 6114 15573
rect 6148 15539 6154 15573
rect 6108 15501 6154 15539
rect 6108 15467 6114 15501
rect 6148 15467 6154 15501
rect 6108 15429 6154 15467
rect 6108 15395 6114 15429
rect 6148 15395 6154 15429
rect 6108 15357 6154 15395
rect 6108 15323 6114 15357
rect 6148 15323 6154 15357
rect 6108 15285 6154 15323
rect 6108 15251 6114 15285
rect 6148 15251 6154 15285
rect 6108 15213 6154 15251
rect 6108 15179 6114 15213
rect 6148 15179 6154 15213
rect 6108 15141 6154 15179
rect 6108 15107 6114 15141
rect 6148 15107 6154 15141
rect 6108 15069 6154 15107
rect 6108 15035 6114 15069
rect 6148 15035 6154 15069
rect 6108 14997 6154 15035
rect 6108 14963 6114 14997
rect 6148 14963 6154 14997
rect 6108 14925 6154 14963
rect 6108 14891 6114 14925
rect 6148 14891 6154 14925
rect 6108 14853 6154 14891
rect 6108 14819 6114 14853
rect 6148 14819 6154 14853
rect 6108 14781 6154 14819
rect 6108 14747 6114 14781
rect 6148 14747 6154 14781
rect 6108 14709 6154 14747
rect 6108 14675 6114 14709
rect 6148 14675 6154 14709
rect 6108 14637 6154 14675
rect 6108 14603 6114 14637
rect 6148 14603 6154 14637
rect 6108 14565 6154 14603
rect 6108 14531 6114 14565
rect 6148 14531 6154 14565
rect 6108 14493 6154 14531
rect 6108 14459 6114 14493
rect 6148 14459 6154 14493
rect 6108 14421 6154 14459
rect 6108 14387 6114 14421
rect 6148 14387 6154 14421
rect 6108 14349 6154 14387
rect 6108 14315 6114 14349
rect 6148 14315 6154 14349
rect 6108 14277 6154 14315
rect 6108 14243 6114 14277
rect 6148 14243 6154 14277
rect 6108 14205 6154 14243
rect 6108 14171 6114 14205
rect 6148 14171 6154 14205
rect 6108 14133 6154 14171
rect 6108 14099 6114 14133
rect 6148 14099 6154 14133
rect 6108 14061 6154 14099
rect 6108 14027 6114 14061
rect 6148 14027 6154 14061
rect 6108 13989 6154 14027
rect 6108 13955 6114 13989
rect 6148 13955 6154 13989
rect 6108 13917 6154 13955
rect 6108 13883 6114 13917
rect 6148 13883 6154 13917
rect 6108 13845 6154 13883
rect 6108 13811 6114 13845
rect 6148 13811 6154 13845
rect 6108 13773 6154 13811
rect 6108 13739 6114 13773
rect 6148 13739 6154 13773
rect 6108 13701 6154 13739
rect 6108 13667 6114 13701
rect 6148 13667 6154 13701
rect 6108 13629 6154 13667
rect 6108 13595 6114 13629
rect 6148 13595 6154 13629
rect 6108 13557 6154 13595
rect 6108 13523 6114 13557
rect 6148 13523 6154 13557
rect 6108 13485 6154 13523
rect 6108 13451 6114 13485
rect 6148 13451 6154 13485
rect 6108 13413 6154 13451
rect 6108 13379 6114 13413
rect 6148 13379 6154 13413
rect 6108 13341 6154 13379
rect 6108 13307 6114 13341
rect 6148 13307 6154 13341
rect 6108 13269 6154 13307
rect 6108 13235 6114 13269
rect 6148 13235 6154 13269
rect 6108 13197 6154 13235
rect 6108 13163 6114 13197
rect 6148 13163 6154 13197
rect 6108 13125 6154 13163
rect 6108 13091 6114 13125
rect 6148 13091 6154 13125
rect 6108 13053 6154 13091
rect 6108 13019 6114 13053
rect 6148 13019 6154 13053
rect 6108 12981 6154 13019
rect 6108 12947 6114 12981
rect 6148 12947 6154 12981
rect 6108 12909 6154 12947
rect 6108 12875 6114 12909
rect 6148 12875 6154 12909
rect 6108 12837 6154 12875
rect 6108 12803 6114 12837
rect 6148 12803 6154 12837
rect 6108 12765 6154 12803
rect 6108 12731 6114 12765
rect 6148 12731 6154 12765
rect 6108 12693 6154 12731
rect 6108 12659 6114 12693
rect 6148 12659 6154 12693
rect 6108 12621 6154 12659
rect 6108 12587 6114 12621
rect 6148 12587 6154 12621
rect 6108 12549 6154 12587
rect 6108 12515 6114 12549
rect 6148 12515 6154 12549
rect 6108 12477 6154 12515
rect 6108 12443 6114 12477
rect 6148 12443 6154 12477
rect 6108 12405 6154 12443
rect 6108 12371 6114 12405
rect 6148 12371 6154 12405
rect 6108 12333 6154 12371
rect 6108 12299 6114 12333
rect 6148 12299 6154 12333
rect 6108 12261 6154 12299
rect 6108 12227 6114 12261
rect 6148 12227 6154 12261
rect 6108 12189 6154 12227
rect 6108 12155 6114 12189
rect 6148 12155 6154 12189
rect 6108 12117 6154 12155
rect 6108 12083 6114 12117
rect 6148 12083 6154 12117
rect 6108 12045 6154 12083
rect 6108 12011 6114 12045
rect 6148 12011 6154 12045
rect 6108 11973 6154 12011
rect 6108 11939 6114 11973
rect 6148 11939 6154 11973
rect 6108 11901 6154 11939
rect 6108 11867 6114 11901
rect 6148 11867 6154 11901
rect 6108 11829 6154 11867
rect 6108 11795 6114 11829
rect 6148 11795 6154 11829
rect 6108 11757 6154 11795
rect 6108 11723 6114 11757
rect 6148 11723 6154 11757
rect 6108 11685 6154 11723
rect 6108 11651 6114 11685
rect 6148 11651 6154 11685
rect 6108 11613 6154 11651
rect 6108 11579 6114 11613
rect 6148 11579 6154 11613
rect 6108 11541 6154 11579
rect 6108 11507 6114 11541
rect 6148 11507 6154 11541
rect 6108 11469 6154 11507
rect 6108 11435 6114 11469
rect 6148 11435 6154 11469
rect 6108 11397 6154 11435
rect 6108 11363 6114 11397
rect 6148 11363 6154 11397
rect 6108 11325 6154 11363
rect 6108 11291 6114 11325
rect 6148 11291 6154 11325
rect 6108 11253 6154 11291
rect 6108 11219 6114 11253
rect 6148 11219 6154 11253
rect 6108 11181 6154 11219
rect 6108 11147 6114 11181
rect 6148 11147 6154 11181
rect 6108 11109 6154 11147
rect 6108 11075 6114 11109
rect 6148 11075 6154 11109
rect 6108 11037 6154 11075
rect 6108 11003 6114 11037
rect 6148 11003 6154 11037
rect 6108 10965 6154 11003
rect 6108 10931 6114 10965
rect 6148 10931 6154 10965
rect 6108 10893 6154 10931
rect 6108 10859 6114 10893
rect 6148 10859 6154 10893
rect 6108 10821 6154 10859
rect 6108 10787 6114 10821
rect 6148 10787 6154 10821
rect 6108 10749 6154 10787
rect 6108 10715 6114 10749
rect 6148 10715 6154 10749
rect 6108 10677 6154 10715
rect 6108 10643 6114 10677
rect 6148 10643 6154 10677
rect 6108 10605 6154 10643
rect 6108 10571 6114 10605
rect 6148 10571 6154 10605
rect 6108 10533 6154 10571
rect 6108 10499 6114 10533
rect 6148 10499 6154 10533
rect 6108 10461 6154 10499
rect 6108 10427 6114 10461
rect 6148 10427 6154 10461
rect 6108 10389 6154 10427
rect 6108 10355 6114 10389
rect 6148 10355 6154 10389
rect 6108 10317 6154 10355
rect 6108 10283 6114 10317
rect 6148 10283 6154 10317
rect 6108 10245 6154 10283
rect 6108 10211 6114 10245
rect 6148 10211 6154 10245
rect 6108 10173 6154 10211
rect 6108 10139 6114 10173
rect 6148 10139 6154 10173
rect 6108 10101 6154 10139
rect 6108 10067 6114 10101
rect 6148 10067 6154 10101
rect 6108 10029 6154 10067
rect 6108 9995 6114 10029
rect 6148 9995 6154 10029
rect 6108 9957 6154 9995
rect 6108 9923 6114 9957
rect 6148 9923 6154 9957
rect 6108 9885 6154 9923
rect 6108 9851 6114 9885
rect 6148 9851 6154 9885
rect 6108 9813 6154 9851
rect 6108 9779 6114 9813
rect 6148 9779 6154 9813
rect 6108 9741 6154 9779
rect 6108 9707 6114 9741
rect 6148 9707 6154 9741
rect 6108 9669 6154 9707
rect 6108 9635 6114 9669
rect 6148 9635 6154 9669
rect 6108 9597 6154 9635
rect 6108 9563 6114 9597
rect 6148 9563 6154 9597
rect 6108 9525 6154 9563
rect 6108 9491 6114 9525
rect 6148 9491 6154 9525
rect 6108 9453 6154 9491
rect 6108 9419 6114 9453
rect 6148 9419 6154 9453
rect 6108 9381 6154 9419
rect 6108 9347 6114 9381
rect 6148 9347 6154 9381
rect 6108 9309 6154 9347
rect 6108 9275 6114 9309
rect 6148 9275 6154 9309
rect 6108 9237 6154 9275
rect 6108 9203 6114 9237
rect 6148 9203 6154 9237
rect 6108 9165 6154 9203
rect 6108 9131 6114 9165
rect 6148 9131 6154 9165
rect 6108 9093 6154 9131
rect 6108 9059 6114 9093
rect 6148 9059 6154 9093
rect 6108 9021 6154 9059
rect 6108 8987 6114 9021
rect 6148 8987 6154 9021
rect 6108 8949 6154 8987
rect 6108 8915 6114 8949
rect 6148 8915 6154 8949
rect 6108 8877 6154 8915
rect 6108 8843 6114 8877
rect 6148 8843 6154 8877
rect 6108 8805 6154 8843
rect 6108 8771 6114 8805
rect 6148 8771 6154 8805
rect 6108 8733 6154 8771
rect 6108 8699 6114 8733
rect 6148 8699 6154 8733
rect 6108 8661 6154 8699
rect 6108 8627 6114 8661
rect 6148 8627 6154 8661
rect 6108 8589 6154 8627
rect 6108 8555 6114 8589
rect 6148 8555 6154 8589
rect 6108 8517 6154 8555
rect 6108 8483 6114 8517
rect 6148 8483 6154 8517
rect 6108 8445 6154 8483
rect 6108 8411 6114 8445
rect 6148 8411 6154 8445
rect 6108 8373 6154 8411
rect 6108 8339 6114 8373
rect 6148 8339 6154 8373
rect 6108 8301 6154 8339
rect 6108 8267 6114 8301
rect 6148 8267 6154 8301
rect 6108 8229 6154 8267
rect 6108 8195 6114 8229
rect 6148 8195 6154 8229
rect 6108 8157 6154 8195
rect 6108 8123 6114 8157
rect 6148 8123 6154 8157
rect 6108 8085 6154 8123
rect 6108 8051 6114 8085
rect 6148 8051 6154 8085
rect 6108 8013 6154 8051
rect 6108 7979 6114 8013
rect 6148 7979 6154 8013
rect 6108 7941 6154 7979
rect 6108 7907 6114 7941
rect 6148 7907 6154 7941
rect 6108 7869 6154 7907
rect 6108 7835 6114 7869
rect 6148 7835 6154 7869
rect 6108 7797 6154 7835
rect 6108 7763 6114 7797
rect 6148 7763 6154 7797
rect 6108 7725 6154 7763
rect 6108 7691 6114 7725
rect 6148 7691 6154 7725
rect 6108 7653 6154 7691
rect 6108 7619 6114 7653
rect 6148 7619 6154 7653
rect 6108 7581 6154 7619
rect 6108 7547 6114 7581
rect 6148 7547 6154 7581
rect 6108 7509 6154 7547
rect 6108 7475 6114 7509
rect 6148 7475 6154 7509
rect 6108 7437 6154 7475
rect 6108 7403 6114 7437
rect 6148 7403 6154 7437
rect 6108 7365 6154 7403
rect 6108 7331 6114 7365
rect 6148 7331 6154 7365
rect 6108 7293 6154 7331
rect 6108 7259 6114 7293
rect 6148 7259 6154 7293
rect 6108 7221 6154 7259
rect 6108 7187 6114 7221
rect 6148 7187 6154 7221
rect 6108 7149 6154 7187
rect 6108 7115 6114 7149
rect 6148 7115 6154 7149
rect 6108 7077 6154 7115
rect 6108 7043 6114 7077
rect 6148 7043 6154 7077
rect 6108 7005 6154 7043
rect 6108 6971 6114 7005
rect 6148 6971 6154 7005
rect 6108 6933 6154 6971
rect 6108 6899 6114 6933
rect 6148 6899 6154 6933
rect 6108 6861 6154 6899
rect 6108 6827 6114 6861
rect 6148 6827 6154 6861
rect 6108 6789 6154 6827
rect 6108 6755 6114 6789
rect 6148 6755 6154 6789
rect 6108 6716 6154 6755
rect 6108 6682 6114 6716
rect 6148 6682 6154 6716
rect 6108 6643 6154 6682
rect 6108 6609 6114 6643
rect 6148 6609 6154 6643
rect 6108 6570 6154 6609
rect 6108 6536 6114 6570
rect 6148 6536 6154 6570
rect 6108 6497 6154 6536
rect 6108 6463 6114 6497
rect 6148 6463 6154 6497
rect 6108 6424 6154 6463
rect 6108 6390 6114 6424
rect 6148 6390 6154 6424
rect 6108 6351 6154 6390
rect 6108 6317 6114 6351
rect 6148 6317 6154 6351
rect 6108 6278 6154 6317
rect 6108 6244 6114 6278
rect 6148 6244 6154 6278
rect 6108 6205 6154 6244
rect 6108 6171 6114 6205
rect 6148 6171 6154 6205
rect 6108 6132 6154 6171
rect 6108 6098 6114 6132
rect 6148 6098 6154 6132
rect 6108 6059 6154 6098
rect 6108 6025 6114 6059
rect 6148 6025 6154 6059
rect 6108 5986 6154 6025
rect 6108 5952 6114 5986
rect 6148 5952 6154 5986
rect 6108 5913 6154 5952
rect 6108 5879 6114 5913
rect 6148 5879 6154 5913
rect 6108 5840 6154 5879
rect 6108 5806 6114 5840
rect 6148 5806 6154 5840
rect 6108 5767 6154 5806
rect 6108 5733 6114 5767
rect 6148 5733 6154 5767
rect 6108 5694 6154 5733
rect 6108 5660 6114 5694
rect 6148 5660 6154 5694
rect 6108 5621 6154 5660
rect 6108 5587 6114 5621
rect 6148 5587 6154 5621
rect 6108 5548 6154 5587
rect 6108 5514 6114 5548
rect 6148 5514 6154 5548
rect 6108 5475 6154 5514
rect 6108 5441 6114 5475
rect 6148 5441 6154 5475
rect 6108 5402 6154 5441
rect 6108 5368 6114 5402
rect 6148 5368 6154 5402
rect 6108 5329 6154 5368
rect 6108 5295 6114 5329
rect 6148 5295 6154 5329
rect 6108 5256 6154 5295
rect 6108 5222 6114 5256
rect 6148 5222 6154 5256
rect 6108 5183 6154 5222
rect 6108 5149 6114 5183
rect 6148 5149 6154 5183
rect 6108 5110 6154 5149
rect 6108 5076 6114 5110
rect 6148 5076 6154 5110
rect 6108 5037 6154 5076
rect 6108 5003 6114 5037
rect 6148 5003 6154 5037
rect 6108 4964 6154 5003
rect 6108 4930 6114 4964
rect 6148 4930 6154 4964
rect 6108 4891 6154 4930
rect 6108 4857 6114 4891
rect 6148 4857 6154 4891
rect 6108 4818 6154 4857
rect 6108 4784 6114 4818
rect 6148 4784 6154 4818
rect 6108 4745 6154 4784
rect 6108 4711 6114 4745
rect 6148 4711 6154 4745
rect 6108 4672 6154 4711
rect 6108 4638 6114 4672
rect 6148 4638 6154 4672
rect 6108 4599 6154 4638
rect 6108 4565 6114 4599
rect 6148 4565 6154 4599
rect 6108 4526 6154 4565
rect 6108 4492 6114 4526
rect 6148 4492 6154 4526
rect 6108 4453 6154 4492
rect 6108 4419 6114 4453
rect 6148 4419 6154 4453
rect 6108 4380 6154 4419
rect 6108 4346 6114 4380
rect 6148 4346 6154 4380
rect 6108 4307 6154 4346
rect 6108 4273 6114 4307
rect 6148 4273 6154 4307
rect 6108 4234 6154 4273
rect 6108 4200 6114 4234
rect 6148 4200 6154 4234
rect 6108 4161 6154 4200
rect 6108 4127 6114 4161
rect 6148 4127 6154 4161
rect 6108 4088 6154 4127
rect 6108 4054 6114 4088
rect 6148 4054 6154 4088
rect 6108 4015 6154 4054
rect 6108 3981 6114 4015
rect 6148 3981 6154 4015
rect 6108 3942 6154 3981
rect 6108 3908 6114 3942
rect 6148 3908 6154 3942
rect 6108 3869 6154 3908
rect 6108 3835 6114 3869
rect 6148 3835 6154 3869
rect 6108 3796 6154 3835
rect 6108 3762 6114 3796
rect 6148 3762 6154 3796
rect 6108 3723 6154 3762
rect 6108 3689 6114 3723
rect 6148 3689 6154 3723
rect 6108 3650 6154 3689
rect 6108 3616 6114 3650
rect 6148 3616 6154 3650
rect 6108 3577 6154 3616
rect 6108 3543 6114 3577
rect 6148 3543 6154 3577
rect 6108 3504 6154 3543
rect 3966 3429 4012 3467
rect 3966 3395 3972 3429
rect 4006 3395 4012 3429
rect 1824 3323 1830 3357
rect 1864 3323 1870 3357
rect 1824 3285 1870 3323
tri -212 3251 -210 3253 sw
tri 1822 3251 1824 3253 se
rect 1824 3251 1830 3285
rect 1864 3251 1870 3285
rect 3966 3357 4012 3395
rect 4149 3492 4201 3499
rect 4149 3428 4201 3440
rect 4149 3369 4201 3376
rect 4267 3487 4437 3499
rect 4267 3453 4276 3487
rect 4310 3453 4394 3487
rect 4428 3453 4437 3487
rect 4267 3415 4437 3453
rect 4267 3381 4276 3415
rect 4310 3381 4394 3415
rect 4428 3381 4437 3415
rect 4267 3369 4437 3381
rect 4503 3487 4673 3499
rect 4503 3453 4512 3487
rect 4546 3453 4630 3487
rect 4664 3453 4673 3487
rect 4503 3415 4673 3453
rect 4503 3381 4512 3415
rect 4546 3381 4630 3415
rect 4664 3381 4673 3415
rect 4503 3369 4673 3381
rect 4739 3487 4909 3499
rect 4739 3453 4748 3487
rect 4782 3453 4866 3487
rect 4900 3453 4909 3487
rect 4739 3415 4909 3453
rect 4739 3381 4748 3415
rect 4782 3381 4866 3415
rect 4900 3381 4909 3415
rect 4739 3369 4909 3381
rect 4975 3487 5145 3499
rect 4975 3453 4984 3487
rect 5018 3453 5102 3487
rect 5136 3453 5145 3487
rect 4975 3415 5145 3453
rect 4975 3381 4984 3415
rect 5018 3381 5102 3415
rect 5136 3381 5145 3415
rect 4975 3369 5145 3381
rect 5211 3486 5381 3499
rect 5211 3452 5220 3486
rect 5254 3452 5338 3486
rect 5372 3452 5381 3486
rect 5211 3414 5381 3452
rect 5211 3380 5220 3414
rect 5254 3380 5338 3414
rect 5372 3380 5381 3414
rect 5211 3368 5381 3380
rect 5447 3486 5617 3499
rect 5447 3452 5456 3486
rect 5490 3452 5574 3486
rect 5608 3452 5617 3486
rect 5447 3414 5617 3452
rect 5447 3380 5456 3414
rect 5490 3380 5574 3414
rect 5608 3380 5617 3414
rect 5447 3368 5617 3380
rect 5683 3486 5853 3499
rect 5683 3452 5692 3486
rect 5726 3452 5810 3486
rect 5844 3452 5853 3486
rect 5683 3414 5853 3452
rect 5683 3380 5692 3414
rect 5726 3380 5810 3414
rect 5844 3380 5853 3414
rect 5683 3368 5853 3380
rect 5919 3492 5971 3499
rect 5919 3428 5971 3440
rect 5919 3368 5971 3376
rect 6108 3470 6114 3504
rect 6148 3470 6154 3504
rect 6108 3431 6154 3470
rect 6108 3397 6114 3431
rect 6148 3397 6154 3431
rect 3966 3323 3972 3357
rect 4006 3323 4012 3357
rect 3966 3285 4012 3323
tri 1870 3251 1872 3253 sw
tri 3964 3251 3966 3253 se
rect 3966 3251 3972 3285
rect 4006 3251 4012 3285
rect 6108 3358 6154 3397
rect 6108 3324 6114 3358
rect 6148 3324 6154 3358
rect 6108 3285 6154 3324
tri 4012 3251 4014 3253 sw
tri 6106 3251 6108 3253 se
rect 6108 3251 6114 3285
rect 6148 3251 6154 3285
rect -258 3250 -210 3251
tri -210 3250 -209 3251 sw
tri 1821 3250 1822 3251 se
rect 1822 3250 1872 3251
tri 1872 3250 1873 3251 sw
tri 3963 3250 3964 3251 se
rect 3964 3250 4014 3251
tri 4014 3250 4015 3251 sw
tri 6105 3250 6106 3251 se
rect 6106 3250 6154 3251
rect -258 3242 -209 3250
tri -209 3242 -201 3250 sw
tri 1813 3242 1821 3250 se
rect 1821 3242 1873 3250
tri 1873 3242 1881 3250 sw
tri 3955 3242 3963 3250 se
rect 3963 3242 4015 3250
tri 4015 3242 4023 3250 sw
tri 6097 3242 6105 3250 se
rect 6105 3242 6154 3250
rect -258 3219 -201 3242
tri -201 3219 -178 3242 sw
tri 1790 3219 1813 3242 se
rect 1813 3219 1881 3242
tri 1881 3219 1904 3242 sw
tri 3932 3219 3955 3242 se
rect 3955 3219 4023 3242
tri 4023 3219 4046 3242 sw
tri 6074 3219 6097 3242 se
rect 6097 3219 6154 3242
rect -258 3213 6154 3219
rect -258 3179 -180 3213
rect -146 3179 -107 3213
rect -73 3179 -34 3213
rect 0 3179 39 3213
rect 73 3179 112 3213
rect 146 3179 185 3213
rect 219 3179 258 3213
rect 292 3179 331 3213
rect 365 3179 404 3213
rect 438 3179 477 3213
rect 511 3179 550 3213
rect 584 3179 623 3213
rect 657 3179 696 3213
rect 730 3179 769 3213
rect 803 3179 842 3213
rect 876 3179 915 3213
rect 949 3179 988 3213
rect 1022 3179 1061 3213
rect 1095 3179 1134 3213
rect 1168 3179 1207 3213
rect 1241 3179 1280 3213
rect 1314 3179 1353 3213
rect 1387 3179 1426 3213
rect 1460 3179 1499 3213
rect 1533 3179 1572 3213
rect 1606 3179 1645 3213
rect 1679 3179 1718 3213
rect 1752 3179 1791 3213
rect 1825 3179 1864 3213
rect 1898 3179 1937 3213
rect 1971 3179 2010 3213
rect 2044 3179 2082 3213
rect 2116 3179 2154 3213
rect 2188 3179 2226 3213
rect 2260 3179 2298 3213
rect 2332 3179 2370 3213
rect 2404 3179 2442 3213
rect 2476 3179 2514 3213
rect 2548 3179 2586 3213
rect 2620 3179 2658 3213
rect 2692 3179 2730 3213
rect 2764 3179 2802 3213
rect 2836 3179 2874 3213
rect 2908 3179 2946 3213
rect 2980 3179 3018 3213
rect 3052 3179 3090 3213
rect 3124 3179 3162 3213
rect 3196 3179 3234 3213
rect 3268 3179 3306 3213
rect 3340 3179 3378 3213
rect 3412 3179 3450 3213
rect 3484 3179 3522 3213
rect 3556 3179 3594 3213
rect 3628 3179 3666 3213
rect 3700 3179 3738 3213
rect 3772 3179 3810 3213
rect 3844 3179 3882 3213
rect 3916 3179 3954 3213
rect 3988 3179 4026 3213
rect 4060 3179 4098 3213
rect 4132 3179 4170 3213
rect 4204 3179 4242 3213
rect 4276 3179 4314 3213
rect 4348 3179 4386 3213
rect 4420 3179 4458 3213
rect 4492 3179 4530 3213
rect 4564 3179 4602 3213
rect 4636 3179 4674 3213
rect 4708 3179 4746 3213
rect 4780 3179 4818 3213
rect 4852 3179 4890 3213
rect 4924 3179 4962 3213
rect 4996 3179 5034 3213
rect 5068 3179 5106 3213
rect 5140 3179 5178 3213
rect 5212 3179 5250 3213
rect 5284 3179 5322 3213
rect 5356 3179 5394 3213
rect 5428 3179 5466 3213
rect 5500 3179 5538 3213
rect 5572 3179 5610 3213
rect 5644 3179 5682 3213
rect 5716 3179 5754 3213
rect 5788 3179 5826 3213
rect 5860 3179 5898 3213
rect 5932 3179 5970 3213
rect 6004 3179 6042 3213
rect 6076 3179 6154 3213
rect -258 3173 6154 3179
rect 9082 38756 14980 38762
rect 9082 38722 9162 38756
rect 9196 38722 9237 38756
rect 9271 38722 9312 38756
rect 9346 38722 9422 38756
rect 9456 38722 9494 38756
rect 9528 38722 9566 38756
rect 9600 38722 9638 38756
rect 9672 38722 9710 38756
rect 9744 38722 9782 38756
rect 9816 38722 9854 38756
rect 9888 38722 9926 38756
rect 9960 38722 9998 38756
rect 10032 38722 10070 38756
rect 10104 38722 10142 38756
rect 10176 38722 10214 38756
rect 10248 38722 10286 38756
rect 10320 38722 10358 38756
rect 10392 38722 10430 38756
rect 10464 38722 10502 38756
rect 10536 38722 10574 38756
rect 10608 38722 10646 38756
rect 10680 38722 10718 38756
rect 10752 38722 10790 38756
rect 10824 38722 10862 38756
rect 10896 38722 10934 38756
rect 10968 38722 11006 38756
rect 11040 38722 11078 38756
rect 11112 38722 11150 38756
rect 11184 38722 11222 38756
rect 11256 38722 11294 38756
rect 11328 38722 11366 38756
rect 11400 38722 11438 38756
rect 11472 38722 11510 38756
rect 11544 38722 11583 38756
rect 11617 38722 11656 38756
rect 11690 38722 11729 38756
rect 11763 38722 11802 38756
rect 11836 38722 11875 38756
rect 11909 38722 11948 38756
rect 11982 38722 12021 38756
rect 12055 38722 12094 38756
rect 12128 38722 12167 38756
rect 12201 38722 12240 38756
rect 12274 38722 12313 38756
rect 12347 38722 12386 38756
rect 12420 38722 12459 38756
rect 12493 38722 12532 38756
rect 12566 38722 12605 38756
rect 12639 38722 12678 38756
rect 12712 38722 12751 38756
rect 12785 38722 12824 38756
rect 12858 38722 12897 38756
rect 12931 38722 12970 38756
rect 13004 38722 13043 38756
rect 13077 38722 13116 38756
rect 13150 38722 13189 38756
rect 13223 38722 13262 38756
rect 13296 38722 13335 38756
rect 13369 38722 13408 38756
rect 13442 38722 13481 38756
rect 13515 38722 13554 38756
rect 13588 38722 13627 38756
rect 13661 38722 13700 38756
rect 13734 38722 13773 38756
rect 13807 38722 13846 38756
rect 13880 38722 13919 38756
rect 13953 38722 13992 38756
rect 14026 38722 14065 38756
rect 14099 38722 14138 38756
rect 14172 38722 14211 38756
rect 14245 38722 14284 38756
rect 14318 38722 14357 38756
rect 14391 38722 14430 38756
rect 14464 38722 14503 38756
rect 14537 38722 14576 38756
rect 14610 38722 14649 38756
rect 14683 38722 14722 38756
rect 14756 38722 14795 38756
rect 14829 38722 14868 38756
rect 14902 38722 14980 38756
rect 9082 38716 14980 38722
rect 9082 38684 9130 38716
tri 9130 38684 9162 38716 nw
tri 10186 38684 10218 38716 ne
rect 10218 38684 10268 38716
tri 10268 38684 10300 38716 nw
tri 11384 38684 11416 38716 ne
rect 11416 38684 11466 38716
tri 11466 38684 11498 38716 nw
tri 13172 38684 13204 38716 ne
rect 13204 38684 13254 38716
tri 13254 38684 13286 38716 nw
tri 14900 38684 14932 38716 ne
rect 14932 38684 14980 38716
rect 9082 38650 9088 38684
rect 9122 38650 9128 38684
tri 9128 38682 9130 38684 nw
tri 10218 38682 10220 38684 ne
rect 9082 38611 9128 38650
rect 9082 38577 9088 38611
rect 9122 38577 9128 38611
rect 9082 38538 9128 38577
rect 9082 38504 9088 38538
rect 9122 38504 9128 38538
rect 9082 38465 9128 38504
rect 9082 38431 9088 38465
rect 9122 38431 9128 38465
rect 9082 38392 9128 38431
rect 9082 38358 9088 38392
rect 9122 38358 9128 38392
rect 9082 38319 9128 38358
rect 9082 38285 9088 38319
rect 9122 38285 9128 38319
rect 9082 38246 9128 38285
rect 9082 38212 9088 38246
rect 9122 38212 9128 38246
rect 9082 38173 9128 38212
rect 9082 38139 9088 38173
rect 9122 38139 9128 38173
rect 9082 38100 9128 38139
rect 9082 38066 9088 38100
rect 9122 38066 9128 38100
rect 9082 38027 9128 38066
rect 9082 37993 9088 38027
rect 9122 37993 9128 38027
rect 9082 37954 9128 37993
rect 9082 37920 9088 37954
rect 9122 37920 9128 37954
rect 9082 37881 9128 37920
rect 9082 37847 9088 37881
rect 9122 37847 9128 37881
rect 9082 37808 9128 37847
rect 9082 37774 9088 37808
rect 9122 37774 9128 37808
rect 9082 37735 9128 37774
rect 9082 37701 9088 37735
rect 9122 37701 9128 37735
rect 9082 37662 9128 37701
rect 9082 37628 9088 37662
rect 9122 37628 9128 37662
rect 9082 37589 9128 37628
rect 9082 37555 9088 37589
rect 9122 37555 9128 37589
rect 9082 37516 9128 37555
rect 9082 37482 9088 37516
rect 9122 37482 9128 37516
rect 9082 37443 9128 37482
rect 9082 37409 9088 37443
rect 9122 37409 9128 37443
rect 9082 37370 9128 37409
rect 9082 37336 9088 37370
rect 9122 37336 9128 37370
rect 9082 37297 9128 37336
rect 9082 37263 9088 37297
rect 9122 37263 9128 37297
rect 9082 37224 9128 37263
rect 9082 37190 9088 37224
rect 9122 37190 9128 37224
rect 9082 37151 9128 37190
rect 9082 37117 9088 37151
rect 9122 37117 9128 37151
rect 9082 37078 9128 37117
rect 9082 37044 9088 37078
rect 9122 37044 9128 37078
rect 9082 37005 9128 37044
rect 9082 36971 9088 37005
rect 9122 36971 9128 37005
rect 9082 36932 9128 36971
rect 9082 36898 9088 36932
rect 9122 36898 9128 36932
rect 9082 36859 9128 36898
rect 9082 36825 9088 36859
rect 9122 36825 9128 36859
rect 9082 36786 9128 36825
rect 9082 36752 9088 36786
rect 9122 36752 9128 36786
rect 9082 36713 9128 36752
rect 9082 36679 9088 36713
rect 9122 36679 9128 36713
rect 9082 36640 9128 36679
rect 9082 36606 9088 36640
rect 9122 36606 9128 36640
rect 9082 36567 9128 36606
rect 9082 36533 9088 36567
rect 9122 36533 9128 36567
rect 9082 36494 9128 36533
rect 9082 36460 9088 36494
rect 9122 36460 9128 36494
rect 9082 36421 9128 36460
rect 9082 36387 9088 36421
rect 9122 36387 9128 36421
rect 9082 36348 9128 36387
rect 9082 36314 9088 36348
rect 9122 36314 9128 36348
rect 9082 36275 9128 36314
rect 9082 36241 9088 36275
rect 9122 36241 9128 36275
rect 9082 36202 9128 36241
rect 9082 36168 9088 36202
rect 9122 36168 9128 36202
rect 9082 36129 9128 36168
rect 9082 36095 9088 36129
rect 9122 36095 9128 36129
rect 9082 36056 9128 36095
rect 9082 36022 9088 36056
rect 9122 36022 9128 36056
rect 9082 35983 9128 36022
rect 9082 35949 9088 35983
rect 9122 35949 9128 35983
rect 9082 35910 9128 35949
rect 9082 35876 9088 35910
rect 9122 35876 9128 35910
rect 9082 35837 9128 35876
rect 9082 35803 9088 35837
rect 9122 35803 9128 35837
rect 9082 35764 9128 35803
rect 9082 35730 9088 35764
rect 9122 35730 9128 35764
rect 9082 35691 9128 35730
rect 9082 35657 9088 35691
rect 9122 35657 9128 35691
rect 9082 35618 9128 35657
rect 9082 35584 9088 35618
rect 9122 35584 9128 35618
rect 9082 35545 9128 35584
rect 9082 35511 9088 35545
rect 9122 35511 9128 35545
rect 9082 35472 9128 35511
rect 9082 35438 9088 35472
rect 9122 35438 9128 35472
rect 9082 35399 9128 35438
rect 9082 35365 9088 35399
rect 9122 35365 9128 35399
rect 9082 35326 9128 35365
rect 9082 35292 9088 35326
rect 9122 35292 9128 35326
rect 9082 35253 9128 35292
rect 9082 35219 9088 35253
rect 9122 35219 9128 35253
rect 9082 35180 9128 35219
rect 9082 35146 9088 35180
rect 9122 35146 9128 35180
rect 9082 35108 9128 35146
rect 9082 35074 9088 35108
rect 9122 35074 9128 35108
rect 9082 35036 9128 35074
rect 9082 35002 9088 35036
rect 9122 35002 9128 35036
rect 9082 34964 9128 35002
rect 9082 34930 9088 34964
rect 9122 34930 9128 34964
rect 9082 34892 9128 34930
rect 9082 34858 9088 34892
rect 9122 34858 9128 34892
rect 9082 34820 9128 34858
rect 9082 34786 9088 34820
rect 9122 34786 9128 34820
rect 9082 34748 9128 34786
rect 9082 34714 9088 34748
rect 9122 34714 9128 34748
rect 9082 34676 9128 34714
rect 9082 34642 9088 34676
rect 9122 34642 9128 34676
rect 9082 34604 9128 34642
rect 9082 34570 9088 34604
rect 9122 34570 9128 34604
rect 9082 34532 9128 34570
rect 9082 34498 9088 34532
rect 9122 34498 9128 34532
rect 9082 34460 9128 34498
rect 9082 34426 9088 34460
rect 9122 34426 9128 34460
rect 9082 34388 9128 34426
rect 9082 34354 9088 34388
rect 9122 34354 9128 34388
rect 9082 34316 9128 34354
rect 9082 34282 9088 34316
rect 9122 34282 9128 34316
rect 9082 34244 9128 34282
rect 9082 34210 9088 34244
rect 9122 34210 9128 34244
rect 9082 34172 9128 34210
rect 9082 34138 9088 34172
rect 9122 34138 9128 34172
rect 9082 34100 9128 34138
rect 9082 34066 9088 34100
rect 9122 34066 9128 34100
rect 9082 34028 9128 34066
rect 9082 33994 9088 34028
rect 9122 33994 9128 34028
rect 9082 33956 9128 33994
rect 9082 33922 9088 33956
rect 9122 33922 9128 33956
rect 9082 33884 9128 33922
rect 9082 33850 9088 33884
rect 9122 33850 9128 33884
rect 9082 33812 9128 33850
rect 9082 33778 9088 33812
rect 9122 33778 9128 33812
rect 9082 33740 9128 33778
rect 9082 33706 9088 33740
rect 9122 33706 9128 33740
rect 9082 33668 9128 33706
rect 9082 33634 9088 33668
rect 9122 33634 9128 33668
rect 9082 33596 9128 33634
rect 9082 33562 9088 33596
rect 9122 33562 9128 33596
rect 9082 33524 9128 33562
rect 9082 33490 9088 33524
rect 9122 33490 9128 33524
rect 9082 33452 9128 33490
rect 9082 33418 9088 33452
rect 9122 33418 9128 33452
rect 9082 33380 9128 33418
rect 9082 33346 9088 33380
rect 9122 33346 9128 33380
rect 9082 33308 9128 33346
rect 9082 33274 9088 33308
rect 9122 33274 9128 33308
rect 9082 33236 9128 33274
rect 9082 33202 9088 33236
rect 9122 33202 9128 33236
rect 9082 33164 9128 33202
rect 9082 33130 9088 33164
rect 9122 33130 9128 33164
rect 9082 33092 9128 33130
rect 9082 33058 9088 33092
rect 9122 33058 9128 33092
rect 9082 33020 9128 33058
rect 9082 32986 9088 33020
rect 9122 32986 9128 33020
rect 9082 32948 9128 32986
rect 9082 32914 9088 32948
rect 9122 32914 9128 32948
rect 9082 32876 9128 32914
rect 9082 32842 9088 32876
rect 9122 32842 9128 32876
rect 9082 32804 9128 32842
rect 9082 32770 9088 32804
rect 9122 32770 9128 32804
rect 9082 32732 9128 32770
rect 9082 32698 9088 32732
rect 9122 32698 9128 32732
rect 9082 32660 9128 32698
rect 9082 32626 9088 32660
rect 9122 32626 9128 32660
rect 9082 32588 9128 32626
rect 9082 32554 9088 32588
rect 9122 32554 9128 32588
rect 9082 32516 9128 32554
rect 9082 32482 9088 32516
rect 9122 32482 9128 32516
rect 9082 32444 9128 32482
rect 9082 32410 9088 32444
rect 9122 32410 9128 32444
rect 9082 32372 9128 32410
rect 9082 32338 9088 32372
rect 9122 32338 9128 32372
rect 9082 32300 9128 32338
rect 9082 32266 9088 32300
rect 9122 32266 9128 32300
rect 9082 32228 9128 32266
rect 9082 32194 9088 32228
rect 9122 32194 9128 32228
rect 9082 32156 9128 32194
rect 9082 32122 9088 32156
rect 9122 32122 9128 32156
rect 9082 32084 9128 32122
rect 9082 32050 9088 32084
rect 9122 32050 9128 32084
rect 9082 32012 9128 32050
rect 9082 31978 9088 32012
rect 9122 31978 9128 32012
rect 9082 31940 9128 31978
rect 9082 31906 9088 31940
rect 9122 31906 9128 31940
rect 9082 31868 9128 31906
rect 9082 31834 9088 31868
rect 9122 31834 9128 31868
rect 9082 31796 9128 31834
rect 9082 31762 9088 31796
rect 9122 31762 9128 31796
rect 9082 31724 9128 31762
rect 9082 31690 9088 31724
rect 9122 31690 9128 31724
rect 9082 31652 9128 31690
rect 9082 31618 9088 31652
rect 9122 31618 9128 31652
rect 9082 31580 9128 31618
rect 9082 31546 9088 31580
rect 9122 31546 9128 31580
rect 9082 31508 9128 31546
rect 9082 31474 9088 31508
rect 9122 31474 9128 31508
rect 9082 31436 9128 31474
rect 9082 31402 9088 31436
rect 9122 31402 9128 31436
rect 9082 31364 9128 31402
rect 9082 31330 9088 31364
rect 9122 31330 9128 31364
rect 9082 31292 9128 31330
rect 9082 31258 9088 31292
rect 9122 31258 9128 31292
rect 9082 31220 9128 31258
rect 9082 31186 9088 31220
rect 9122 31186 9128 31220
rect 9082 31148 9128 31186
rect 9082 31114 9088 31148
rect 9122 31114 9128 31148
rect 9082 31076 9128 31114
rect 9082 31042 9088 31076
rect 9122 31042 9128 31076
rect 9082 31004 9128 31042
rect 9082 30970 9088 31004
rect 9122 30970 9128 31004
rect 9082 30932 9128 30970
rect 9082 30898 9088 30932
rect 9122 30898 9128 30932
rect 9082 30860 9128 30898
rect 9082 30826 9088 30860
rect 9122 30826 9128 30860
rect 9082 30788 9128 30826
rect 9082 30754 9088 30788
rect 9122 30754 9128 30788
rect 9082 30716 9128 30754
rect 9082 30682 9088 30716
rect 9122 30682 9128 30716
rect 9082 30644 9128 30682
rect 9082 30610 9088 30644
rect 9122 30610 9128 30644
rect 9082 30572 9128 30610
rect 9082 30538 9088 30572
rect 9122 30538 9128 30572
rect 9082 30500 9128 30538
rect 9082 30466 9088 30500
rect 9122 30466 9128 30500
rect 9082 30428 9128 30466
rect 9082 30394 9088 30428
rect 9122 30394 9128 30428
rect 9082 30356 9128 30394
rect 9082 30322 9088 30356
rect 9122 30322 9128 30356
rect 9082 30284 9128 30322
rect 9082 30250 9088 30284
rect 9122 30250 9128 30284
rect 9082 30212 9128 30250
rect 9082 30178 9088 30212
rect 9122 30178 9128 30212
rect 9082 30140 9128 30178
rect 9082 30106 9088 30140
rect 9122 30106 9128 30140
rect 9082 30068 9128 30106
rect 9082 30034 9088 30068
rect 9122 30034 9128 30068
rect 9082 29996 9128 30034
rect 9082 29962 9088 29996
rect 9122 29962 9128 29996
rect 9082 29924 9128 29962
rect 9082 29890 9088 29924
rect 9122 29890 9128 29924
rect 9082 29852 9128 29890
rect 9082 29818 9088 29852
rect 9122 29818 9128 29852
rect 9082 29780 9128 29818
rect 9082 29746 9088 29780
rect 9122 29746 9128 29780
rect 9082 29708 9128 29746
rect 9082 29674 9088 29708
rect 9122 29674 9128 29708
rect 9082 29636 9128 29674
rect 9082 29602 9088 29636
rect 9122 29602 9128 29636
rect 9082 29564 9128 29602
rect 9082 29530 9088 29564
rect 9122 29530 9128 29564
rect 9082 29492 9128 29530
rect 9082 29458 9088 29492
rect 9122 29458 9128 29492
rect 9082 29420 9128 29458
rect 9082 29386 9088 29420
rect 9122 29386 9128 29420
rect 9082 29348 9128 29386
rect 9082 29314 9088 29348
rect 9122 29314 9128 29348
rect 9082 29276 9128 29314
rect 9082 29242 9088 29276
rect 9122 29242 9128 29276
rect 9082 29204 9128 29242
rect 9082 29170 9088 29204
rect 9122 29170 9128 29204
rect 9082 29132 9128 29170
rect 9082 29098 9088 29132
rect 9122 29098 9128 29132
rect 9082 29060 9128 29098
rect 9082 29026 9088 29060
rect 9122 29026 9128 29060
rect 9082 28988 9128 29026
rect 9082 28954 9088 28988
rect 9122 28954 9128 28988
rect 9082 28916 9128 28954
rect 9082 28882 9088 28916
rect 9122 28882 9128 28916
rect 9082 28844 9128 28882
rect 9082 28810 9088 28844
rect 9122 28810 9128 28844
rect 9082 28772 9128 28810
rect 9082 28738 9088 28772
rect 9122 28738 9128 28772
rect 9082 28700 9128 28738
rect 9082 28666 9088 28700
rect 9122 28666 9128 28700
rect 9082 28628 9128 28666
rect 9082 28594 9088 28628
rect 9122 28594 9128 28628
rect 9082 28556 9128 28594
rect 9082 28522 9088 28556
rect 9122 28522 9128 28556
rect 9082 28484 9128 28522
rect 9082 28450 9088 28484
rect 9122 28450 9128 28484
rect 9082 28412 9128 28450
rect 9082 28378 9088 28412
rect 9122 28378 9128 28412
rect 9082 28340 9128 28378
rect 9082 28306 9088 28340
rect 9122 28306 9128 28340
rect 9082 28268 9128 28306
rect 9082 28234 9088 28268
rect 9122 28234 9128 28268
rect 9082 28196 9128 28234
rect 9082 28162 9088 28196
rect 9122 28162 9128 28196
rect 9082 28124 9128 28162
rect 9082 28090 9088 28124
rect 9122 28090 9128 28124
rect 9082 28052 9128 28090
rect 9082 28018 9088 28052
rect 9122 28018 9128 28052
rect 9082 27980 9128 28018
rect 9082 27946 9088 27980
rect 9122 27946 9128 27980
rect 9082 27908 9128 27946
rect 9082 27874 9088 27908
rect 9122 27874 9128 27908
rect 9082 27836 9128 27874
rect 9082 27802 9088 27836
rect 9122 27802 9128 27836
rect 9082 27764 9128 27802
rect 9082 27730 9088 27764
rect 9122 27730 9128 27764
rect 9082 27692 9128 27730
rect 9082 27658 9088 27692
rect 9122 27658 9128 27692
rect 9082 27620 9128 27658
rect 9082 27586 9088 27620
rect 9122 27586 9128 27620
rect 9082 27548 9128 27586
rect 9082 27514 9088 27548
rect 9122 27514 9128 27548
rect 9082 27476 9128 27514
rect 9082 27442 9088 27476
rect 9122 27442 9128 27476
rect 9082 27404 9128 27442
rect 9082 27370 9088 27404
rect 9122 27370 9128 27404
rect 9082 27332 9128 27370
rect 9082 27298 9088 27332
rect 9122 27298 9128 27332
rect 9082 27260 9128 27298
rect 9082 27226 9088 27260
rect 9122 27226 9128 27260
rect 9082 27188 9128 27226
rect 9082 27154 9088 27188
rect 9122 27154 9128 27188
rect 9082 27116 9128 27154
rect 9082 27082 9088 27116
rect 9122 27082 9128 27116
rect 9082 27044 9128 27082
rect 9082 27010 9088 27044
rect 9122 27010 9128 27044
rect 9082 26972 9128 27010
rect 9082 26938 9088 26972
rect 9122 26938 9128 26972
rect 9082 26900 9128 26938
rect 9082 26866 9088 26900
rect 9122 26866 9128 26900
rect 9082 26828 9128 26866
rect 9082 26794 9088 26828
rect 9122 26794 9128 26828
rect 9082 26756 9128 26794
rect 9082 26722 9088 26756
rect 9122 26722 9128 26756
rect 9082 26684 9128 26722
rect 9082 26650 9088 26684
rect 9122 26650 9128 26684
rect 9082 26612 9128 26650
rect 9082 26578 9088 26612
rect 9122 26578 9128 26612
rect 9082 26540 9128 26578
rect 9082 26506 9088 26540
rect 9122 26506 9128 26540
rect 9082 26468 9128 26506
rect 9082 26434 9088 26468
rect 9122 26434 9128 26468
rect 9082 26396 9128 26434
rect 9082 26362 9088 26396
rect 9122 26362 9128 26396
rect 9082 26324 9128 26362
rect 9082 26290 9088 26324
rect 9122 26290 9128 26324
rect 9082 26252 9128 26290
rect 9082 26218 9088 26252
rect 9122 26218 9128 26252
rect 9082 26180 9128 26218
rect 9082 26146 9088 26180
rect 9122 26146 9128 26180
rect 9082 26108 9128 26146
rect 9082 26074 9088 26108
rect 9122 26074 9128 26108
rect 9082 26036 9128 26074
rect 9082 26002 9088 26036
rect 9122 26002 9128 26036
rect 9082 25964 9128 26002
rect 9082 25930 9088 25964
rect 9122 25930 9128 25964
rect 9082 25892 9128 25930
rect 9082 25858 9088 25892
rect 9122 25858 9128 25892
rect 9082 25820 9128 25858
rect 9082 25786 9088 25820
rect 9122 25786 9128 25820
rect 9082 25748 9128 25786
rect 9082 25714 9088 25748
rect 9122 25714 9128 25748
rect 9082 25676 9128 25714
rect 9082 25642 9088 25676
rect 9122 25642 9128 25676
rect 9082 25604 9128 25642
rect 9082 25570 9088 25604
rect 9122 25570 9128 25604
rect 9082 25532 9128 25570
rect 9082 25498 9088 25532
rect 9122 25498 9128 25532
rect 9082 25460 9128 25498
rect 9082 25426 9088 25460
rect 9122 25426 9128 25460
rect 9082 25388 9128 25426
rect 9082 25354 9088 25388
rect 9122 25354 9128 25388
rect 9082 25316 9128 25354
rect 9082 25282 9088 25316
rect 9122 25282 9128 25316
rect 9082 25244 9128 25282
rect 9082 25210 9088 25244
rect 9122 25210 9128 25244
rect 9082 25172 9128 25210
rect 9082 25138 9088 25172
rect 9122 25138 9128 25172
rect 9082 25100 9128 25138
rect 9082 25066 9088 25100
rect 9122 25066 9128 25100
rect 9082 25028 9128 25066
rect 9082 24994 9088 25028
rect 9122 24994 9128 25028
rect 9082 24956 9128 24994
rect 9082 24922 9088 24956
rect 9122 24922 9128 24956
rect 9082 24884 9128 24922
rect 9082 24850 9088 24884
rect 9122 24850 9128 24884
rect 9082 24812 9128 24850
rect 9082 24778 9088 24812
rect 9122 24778 9128 24812
rect 9082 24740 9128 24778
rect 9082 24706 9088 24740
rect 9122 24706 9128 24740
rect 9082 24668 9128 24706
rect 9082 24634 9088 24668
rect 9122 24634 9128 24668
rect 9082 24596 9128 24634
rect 9082 24562 9088 24596
rect 9122 24562 9128 24596
rect 9082 24524 9128 24562
rect 9082 24490 9088 24524
rect 9122 24490 9128 24524
rect 9082 24452 9128 24490
rect 9082 24418 9088 24452
rect 9122 24418 9128 24452
rect 9082 24380 9128 24418
rect 9082 24346 9088 24380
rect 9122 24346 9128 24380
rect 9082 24308 9128 24346
rect 9082 24274 9088 24308
rect 9122 24274 9128 24308
rect 9082 24236 9128 24274
rect 9082 24202 9088 24236
rect 9122 24202 9128 24236
rect 9082 24164 9128 24202
rect 9082 24130 9088 24164
rect 9122 24130 9128 24164
rect 9082 24092 9128 24130
rect 9082 24058 9088 24092
rect 9122 24058 9128 24092
rect 9082 24020 9128 24058
rect 9082 23986 9088 24020
rect 9122 23986 9128 24020
rect 9082 23948 9128 23986
rect 9082 23914 9088 23948
rect 9122 23914 9128 23948
rect 9082 23876 9128 23914
rect 9082 23842 9088 23876
rect 9122 23842 9128 23876
rect 9082 23804 9128 23842
rect 9082 23770 9088 23804
rect 9122 23770 9128 23804
rect 9082 23732 9128 23770
rect 9082 23698 9088 23732
rect 9122 23698 9128 23732
rect 9082 23660 9128 23698
rect 9082 23626 9088 23660
rect 9122 23626 9128 23660
rect 9082 23588 9128 23626
rect 9082 23554 9088 23588
rect 9122 23554 9128 23588
rect 9082 23516 9128 23554
rect 9082 23482 9088 23516
rect 9122 23482 9128 23516
rect 9082 23444 9128 23482
rect 9082 23410 9088 23444
rect 9122 23410 9128 23444
rect 9082 23372 9128 23410
rect 9082 23338 9088 23372
rect 9122 23338 9128 23372
rect 9082 23300 9128 23338
rect 9082 23266 9088 23300
rect 9122 23266 9128 23300
rect 9082 23228 9128 23266
rect 9082 23194 9088 23228
rect 9122 23194 9128 23228
rect 9082 23156 9128 23194
rect 9082 23122 9088 23156
rect 9122 23122 9128 23156
rect 9082 23084 9128 23122
rect 9082 23050 9088 23084
rect 9122 23050 9128 23084
rect 9082 23012 9128 23050
rect 9082 22978 9088 23012
rect 9122 22978 9128 23012
rect 9082 22940 9128 22978
rect 9082 22906 9088 22940
rect 9122 22906 9128 22940
rect 9082 22868 9128 22906
rect 9082 22834 9088 22868
rect 9122 22834 9128 22868
rect 9082 22796 9128 22834
rect 9082 22762 9088 22796
rect 9122 22762 9128 22796
rect 9082 22724 9128 22762
rect 9082 22690 9088 22724
rect 9122 22690 9128 22724
rect 9082 22652 9128 22690
rect 9082 22618 9088 22652
rect 9122 22618 9128 22652
rect 9082 22580 9128 22618
rect 9082 22546 9088 22580
rect 9122 22546 9128 22580
rect 9082 22508 9128 22546
rect 9082 22474 9088 22508
rect 9122 22474 9128 22508
rect 9082 22436 9128 22474
rect 9082 22402 9088 22436
rect 9122 22402 9128 22436
rect 9082 22364 9128 22402
rect 9082 22330 9088 22364
rect 9122 22330 9128 22364
rect 9082 22292 9128 22330
rect 9082 22258 9088 22292
rect 9122 22258 9128 22292
rect 9082 22220 9128 22258
rect 9082 22186 9088 22220
rect 9122 22186 9128 22220
rect 9082 22148 9128 22186
rect 9082 22114 9088 22148
rect 9122 22114 9128 22148
rect 9082 22076 9128 22114
rect 9082 22042 9088 22076
rect 9122 22042 9128 22076
rect 9082 22004 9128 22042
rect 9082 21970 9088 22004
rect 9122 21970 9128 22004
rect 9082 21932 9128 21970
rect 9082 21898 9088 21932
rect 9122 21898 9128 21932
rect 9082 21860 9128 21898
rect 9082 21826 9088 21860
rect 9122 21826 9128 21860
rect 9082 21788 9128 21826
rect 9082 21754 9088 21788
rect 9122 21754 9128 21788
rect 9082 21716 9128 21754
rect 9082 21682 9088 21716
rect 9122 21682 9128 21716
rect 9082 21644 9128 21682
rect 9082 21610 9088 21644
rect 9122 21610 9128 21644
rect 9082 21572 9128 21610
rect 9082 21538 9088 21572
rect 9122 21538 9128 21572
rect 9082 21500 9128 21538
rect 9082 21466 9088 21500
rect 9122 21466 9128 21500
rect 9082 21428 9128 21466
rect 9082 21394 9088 21428
rect 9122 21394 9128 21428
rect 9082 21356 9128 21394
rect 9082 21322 9088 21356
rect 9122 21322 9128 21356
rect 9082 21284 9128 21322
rect 9082 21250 9088 21284
rect 9122 21250 9128 21284
rect 9082 21212 9128 21250
rect 9082 21178 9088 21212
rect 9122 21178 9128 21212
rect 9082 21140 9128 21178
rect 9082 21106 9088 21140
rect 9122 21106 9128 21140
rect 9082 21068 9128 21106
rect 9082 21034 9088 21068
rect 9122 21034 9128 21068
rect 9082 20996 9128 21034
rect 9082 20962 9088 20996
rect 9122 20962 9128 20996
rect 9082 20924 9128 20962
rect 9082 20890 9088 20924
rect 9122 20890 9128 20924
rect 9082 20852 9128 20890
rect 9082 20818 9088 20852
rect 9122 20818 9128 20852
rect 9082 20780 9128 20818
rect 9082 20746 9088 20780
rect 9122 20746 9128 20780
rect 9082 20708 9128 20746
rect 9082 20674 9088 20708
rect 9122 20674 9128 20708
rect 9082 20636 9128 20674
rect 9082 20602 9088 20636
rect 9122 20602 9128 20636
rect 9082 20564 9128 20602
rect 9082 20530 9088 20564
rect 9122 20530 9128 20564
rect 9082 20492 9128 20530
rect 9082 20458 9088 20492
rect 9122 20458 9128 20492
rect 9082 20420 9128 20458
rect 9082 20386 9088 20420
rect 9122 20386 9128 20420
rect 9082 20348 9128 20386
rect 9082 20314 9088 20348
rect 9122 20314 9128 20348
rect 9082 20276 9128 20314
rect 9082 20242 9088 20276
rect 9122 20242 9128 20276
rect 9082 20204 9128 20242
rect 9082 20170 9088 20204
rect 9122 20170 9128 20204
rect 9082 20132 9128 20170
rect 9082 20098 9088 20132
rect 9122 20098 9128 20132
rect 9082 20060 9128 20098
rect 9082 20026 9088 20060
rect 9122 20026 9128 20060
rect 9082 19988 9128 20026
rect 9082 19954 9088 19988
rect 9122 19954 9128 19988
rect 9082 19916 9128 19954
rect 9082 19882 9088 19916
rect 9122 19882 9128 19916
rect 9082 19844 9128 19882
rect 9082 19810 9088 19844
rect 9122 19810 9128 19844
rect 9082 19772 9128 19810
rect 9082 19738 9088 19772
rect 9122 19738 9128 19772
rect 9082 19700 9128 19738
rect 9082 19666 9088 19700
rect 9122 19666 9128 19700
rect 9082 19628 9128 19666
rect 9082 19594 9088 19628
rect 9122 19594 9128 19628
rect 9082 19556 9128 19594
rect 9082 19522 9088 19556
rect 9122 19522 9128 19556
rect 9082 19484 9128 19522
rect 9082 19450 9088 19484
rect 9122 19450 9128 19484
rect 9082 19412 9128 19450
rect 9082 19378 9088 19412
rect 9122 19378 9128 19412
rect 9082 19340 9128 19378
rect 9082 19306 9088 19340
rect 9122 19306 9128 19340
rect 9082 19268 9128 19306
rect 9082 19234 9088 19268
rect 9122 19234 9128 19268
rect 9082 19196 9128 19234
rect 9082 19162 9088 19196
rect 9122 19162 9128 19196
rect 9082 19124 9128 19162
rect 9082 19090 9088 19124
rect 9122 19090 9128 19124
rect 9082 19052 9128 19090
rect 9082 19018 9088 19052
rect 9122 19018 9128 19052
rect 9082 18980 9128 19018
rect 9082 18946 9088 18980
rect 9122 18946 9128 18980
rect 9082 18908 9128 18946
rect 9082 18874 9088 18908
rect 9122 18874 9128 18908
rect 9082 18836 9128 18874
rect 9082 18802 9088 18836
rect 9122 18802 9128 18836
rect 9082 18764 9128 18802
rect 9082 18730 9088 18764
rect 9122 18730 9128 18764
rect 9082 18692 9128 18730
rect 9082 18658 9088 18692
rect 9122 18658 9128 18692
rect 9082 18620 9128 18658
rect 9082 18586 9088 18620
rect 9122 18586 9128 18620
rect 9082 18548 9128 18586
rect 9082 18514 9088 18548
rect 9122 18514 9128 18548
rect 9082 18476 9128 18514
rect 9082 18442 9088 18476
rect 9122 18442 9128 18476
rect 9082 18404 9128 18442
rect 9082 18370 9088 18404
rect 9122 18370 9128 18404
rect 9082 18332 9128 18370
rect 9082 18298 9088 18332
rect 9122 18298 9128 18332
rect 9082 18260 9128 18298
rect 9082 18226 9088 18260
rect 9122 18226 9128 18260
rect 9082 18188 9128 18226
rect 9082 18154 9088 18188
rect 9122 18154 9128 18188
rect 9082 18116 9128 18154
rect 9082 18082 9088 18116
rect 9122 18082 9128 18116
rect 9082 18044 9128 18082
rect 9082 18010 9088 18044
rect 9122 18010 9128 18044
rect 9082 17972 9128 18010
rect 9082 17938 9088 17972
rect 9122 17938 9128 17972
rect 9082 17900 9128 17938
rect 9082 17866 9088 17900
rect 9122 17866 9128 17900
rect 9082 17828 9128 17866
rect 9082 17794 9088 17828
rect 9122 17794 9128 17828
rect 9082 17756 9128 17794
rect 9082 17722 9088 17756
rect 9122 17722 9128 17756
rect 9082 17684 9128 17722
rect 9082 17650 9088 17684
rect 9122 17650 9128 17684
rect 9082 17612 9128 17650
rect 9082 17578 9088 17612
rect 9122 17578 9128 17612
rect 9082 17540 9128 17578
rect 9082 17506 9088 17540
rect 9122 17506 9128 17540
rect 9082 17468 9128 17506
rect 9082 17434 9088 17468
rect 9122 17434 9128 17468
rect 9082 17396 9128 17434
rect 9082 17362 9088 17396
rect 9122 17362 9128 17396
rect 9082 17324 9128 17362
rect 9082 17290 9088 17324
rect 9122 17290 9128 17324
rect 9082 17252 9128 17290
rect 9082 17218 9088 17252
rect 9122 17218 9128 17252
rect 9082 17180 9128 17218
rect 9082 17146 9088 17180
rect 9122 17146 9128 17180
rect 9082 17108 9128 17146
rect 9082 17074 9088 17108
rect 9122 17074 9128 17108
rect 9082 17036 9128 17074
rect 9082 17002 9088 17036
rect 9122 17002 9128 17036
rect 9082 16964 9128 17002
rect 9082 16930 9088 16964
rect 9122 16930 9128 16964
rect 9082 16892 9128 16930
rect 9082 16858 9088 16892
rect 9122 16858 9128 16892
rect 9082 16820 9128 16858
rect 9082 16786 9088 16820
rect 9122 16786 9128 16820
rect 9082 16748 9128 16786
rect 9082 16714 9088 16748
rect 9122 16714 9128 16748
rect 9082 16676 9128 16714
rect 9082 16642 9088 16676
rect 9122 16642 9128 16676
rect 9082 16604 9128 16642
rect 9082 16570 9088 16604
rect 9122 16570 9128 16604
rect 9082 16532 9128 16570
rect 9082 16498 9088 16532
rect 9122 16498 9128 16532
rect 9082 16460 9128 16498
rect 9082 16426 9088 16460
rect 9122 16426 9128 16460
rect 9082 16388 9128 16426
rect 9082 16354 9088 16388
rect 9122 16354 9128 16388
rect 9082 16316 9128 16354
rect 9082 16282 9088 16316
rect 9122 16282 9128 16316
rect 9082 16244 9128 16282
rect 9082 16210 9088 16244
rect 9122 16210 9128 16244
rect 9082 16172 9128 16210
rect 9082 16138 9088 16172
rect 9122 16138 9128 16172
rect 9082 16100 9128 16138
rect 9082 16066 9088 16100
rect 9122 16066 9128 16100
rect 9082 16028 9128 16066
rect 9082 15994 9088 16028
rect 9122 15994 9128 16028
rect 9082 15956 9128 15994
rect 9082 15922 9088 15956
rect 9122 15922 9128 15956
rect 9082 15884 9128 15922
rect 9082 15850 9088 15884
rect 9122 15850 9128 15884
rect 9082 15812 9128 15850
rect 9082 15778 9088 15812
rect 9122 15778 9128 15812
rect 9082 15740 9128 15778
rect 9082 15706 9088 15740
rect 9122 15706 9128 15740
rect 9082 15668 9128 15706
rect 9082 15634 9088 15668
rect 9122 15634 9128 15668
rect 9082 15596 9128 15634
rect 9082 15562 9088 15596
rect 9122 15562 9128 15596
rect 9082 15524 9128 15562
rect 9082 15490 9088 15524
rect 9122 15490 9128 15524
rect 9082 15452 9128 15490
rect 9082 15418 9088 15452
rect 9122 15418 9128 15452
rect 9082 15380 9128 15418
rect 9082 15346 9088 15380
rect 9122 15346 9128 15380
rect 9082 15308 9128 15346
rect 9082 15274 9088 15308
rect 9122 15274 9128 15308
rect 9082 15236 9128 15274
rect 9082 15202 9088 15236
rect 9122 15202 9128 15236
rect 9082 15164 9128 15202
rect 9082 15130 9088 15164
rect 9122 15130 9128 15164
rect 9082 15092 9128 15130
rect 9082 15058 9088 15092
rect 9122 15058 9128 15092
rect 9082 15020 9128 15058
rect 9082 14986 9088 15020
rect 9122 14986 9128 15020
rect 9082 14948 9128 14986
rect 9082 14914 9088 14948
rect 9122 14914 9128 14948
rect 9082 14876 9128 14914
rect 9082 14842 9088 14876
rect 9122 14842 9128 14876
rect 9082 14804 9128 14842
rect 9082 14770 9088 14804
rect 9122 14770 9128 14804
rect 9082 14732 9128 14770
rect 9082 14698 9088 14732
rect 9122 14698 9128 14732
rect 9082 14660 9128 14698
rect 9082 14626 9088 14660
rect 9122 14626 9128 14660
rect 9082 14588 9128 14626
rect 9082 14554 9088 14588
rect 9122 14554 9128 14588
rect 9082 14516 9128 14554
rect 9082 14482 9088 14516
rect 9122 14482 9128 14516
rect 9082 14444 9128 14482
rect 9082 14410 9088 14444
rect 9122 14410 9128 14444
rect 9082 14372 9128 14410
rect 9082 14338 9088 14372
rect 9122 14338 9128 14372
rect 9082 14300 9128 14338
rect 9082 14266 9088 14300
rect 9122 14266 9128 14300
rect 9082 14228 9128 14266
rect 9082 14194 9088 14228
rect 9122 14194 9128 14228
rect 9082 14156 9128 14194
rect 9082 14122 9088 14156
rect 9122 14122 9128 14156
rect 9082 14084 9128 14122
rect 9082 14050 9088 14084
rect 9122 14050 9128 14084
rect 9082 14012 9128 14050
rect 9082 13978 9088 14012
rect 9122 13978 9128 14012
rect 9082 13940 9128 13978
rect 9082 13906 9088 13940
rect 9122 13906 9128 13940
rect 9082 13868 9128 13906
rect 9082 13834 9088 13868
rect 9122 13834 9128 13868
rect 9082 13796 9128 13834
rect 9082 13762 9088 13796
rect 9122 13762 9128 13796
rect 9082 13724 9128 13762
rect 9082 13690 9088 13724
rect 9122 13690 9128 13724
rect 9082 13652 9128 13690
rect 9082 13618 9088 13652
rect 9122 13618 9128 13652
rect 9082 13580 9128 13618
rect 9082 13546 9088 13580
rect 9122 13546 9128 13580
rect 9082 13508 9128 13546
rect 9082 13474 9088 13508
rect 9122 13474 9128 13508
rect 9082 13436 9128 13474
rect 9082 13402 9088 13436
rect 9122 13402 9128 13436
rect 9082 13364 9128 13402
rect 9082 13330 9088 13364
rect 9122 13330 9128 13364
rect 9082 13292 9128 13330
rect 9082 13258 9088 13292
rect 9122 13258 9128 13292
rect 9082 13220 9128 13258
rect 9082 13186 9088 13220
rect 9122 13186 9128 13220
rect 9082 13148 9128 13186
rect 9082 13114 9088 13148
rect 9122 13114 9128 13148
rect 9082 13076 9128 13114
rect 9082 13042 9088 13076
rect 9122 13042 9128 13076
rect 9082 13004 9128 13042
rect 9082 12970 9088 13004
rect 9122 12970 9128 13004
rect 9082 12932 9128 12970
rect 9082 12898 9088 12932
rect 9122 12898 9128 12932
rect 9082 12860 9128 12898
rect 9082 12826 9088 12860
rect 9122 12826 9128 12860
rect 9082 12788 9128 12826
rect 9082 12754 9088 12788
rect 9122 12754 9128 12788
rect 9082 12716 9128 12754
rect 9082 12682 9088 12716
rect 9122 12682 9128 12716
rect 9082 12644 9128 12682
rect 9082 12610 9088 12644
rect 9122 12610 9128 12644
rect 9082 12572 9128 12610
rect 9082 12538 9088 12572
rect 9122 12538 9128 12572
rect 9082 12500 9128 12538
rect 9082 12466 9088 12500
rect 9122 12466 9128 12500
rect 9082 12428 9128 12466
rect 9082 12394 9088 12428
rect 9122 12394 9128 12428
rect 9082 12356 9128 12394
rect 9082 12322 9088 12356
rect 9122 12322 9128 12356
rect 9082 12284 9128 12322
rect 9082 12250 9088 12284
rect 9122 12250 9128 12284
rect 9082 12212 9128 12250
rect 9082 12178 9088 12212
rect 9122 12178 9128 12212
rect 9082 12140 9128 12178
rect 9082 12106 9088 12140
rect 9122 12106 9128 12140
rect 9082 12068 9128 12106
rect 9082 12034 9088 12068
rect 9122 12034 9128 12068
rect 9082 11996 9128 12034
rect 9082 11962 9088 11996
rect 9122 11962 9128 11996
rect 9082 11924 9128 11962
rect 9082 11890 9088 11924
rect 9122 11890 9128 11924
rect 9082 11852 9128 11890
rect 9082 11818 9088 11852
rect 9122 11818 9128 11852
rect 9082 11780 9128 11818
rect 9082 11746 9088 11780
rect 9122 11746 9128 11780
rect 9082 11708 9128 11746
rect 9082 11674 9088 11708
rect 9122 11674 9128 11708
rect 9082 11636 9128 11674
rect 9082 11602 9088 11636
rect 9122 11602 9128 11636
rect 9082 11564 9128 11602
rect 9082 11530 9088 11564
rect 9122 11530 9128 11564
rect 9082 11492 9128 11530
rect 9082 11458 9088 11492
rect 9122 11458 9128 11492
rect 9082 11420 9128 11458
rect 9082 11386 9088 11420
rect 9122 11386 9128 11420
rect 9082 11348 9128 11386
rect 9082 11314 9088 11348
rect 9122 11314 9128 11348
rect 9082 11276 9128 11314
rect 9082 11242 9088 11276
rect 9122 11242 9128 11276
rect 9082 11204 9128 11242
rect 9082 11170 9088 11204
rect 9122 11170 9128 11204
rect 9082 11132 9128 11170
rect 9082 11098 9088 11132
rect 9122 11098 9128 11132
rect 9082 11060 9128 11098
rect 9082 11026 9088 11060
rect 9122 11026 9128 11060
rect 9082 10988 9128 11026
rect 9082 10954 9088 10988
rect 9122 10954 9128 10988
rect 9082 10916 9128 10954
rect 9082 10882 9088 10916
rect 9122 10882 9128 10916
rect 9082 10844 9128 10882
rect 9082 10810 9088 10844
rect 9122 10810 9128 10844
rect 9082 10772 9128 10810
rect 9082 10738 9088 10772
rect 9122 10738 9128 10772
rect 9082 10700 9128 10738
rect 9082 10666 9088 10700
rect 9122 10666 9128 10700
rect 9082 10628 9128 10666
rect 9082 10594 9088 10628
rect 9122 10594 9128 10628
rect 9082 10556 9128 10594
rect 9082 10522 9088 10556
rect 9122 10522 9128 10556
rect 9082 10484 9128 10522
rect 9082 10450 9088 10484
rect 9122 10450 9128 10484
rect 9082 10412 9128 10450
rect 9082 10378 9088 10412
rect 9122 10378 9128 10412
rect 9082 10340 9128 10378
rect 9082 10306 9088 10340
rect 9122 10306 9128 10340
rect 9082 10268 9128 10306
rect 9082 10234 9088 10268
rect 9122 10234 9128 10268
rect 9082 10196 9128 10234
rect 9082 10162 9088 10196
rect 9122 10162 9128 10196
rect 9082 10124 9128 10162
rect 9082 10090 9088 10124
rect 9122 10090 9128 10124
rect 9082 10052 9128 10090
rect 9082 10018 9088 10052
rect 9122 10018 9128 10052
rect 9082 9980 9128 10018
rect 9082 9946 9088 9980
rect 9122 9946 9128 9980
rect 9082 9908 9128 9946
rect 9082 9874 9088 9908
rect 9122 9874 9128 9908
rect 9082 9836 9128 9874
rect 9082 9802 9088 9836
rect 9122 9802 9128 9836
rect 9082 9764 9128 9802
rect 9082 9730 9088 9764
rect 9122 9730 9128 9764
rect 9082 9692 9128 9730
rect 9082 9658 9088 9692
rect 9122 9658 9128 9692
rect 9082 9620 9128 9658
rect 9082 9586 9088 9620
rect 9122 9586 9128 9620
rect 9082 9548 9128 9586
rect 9082 9514 9088 9548
rect 9122 9514 9128 9548
rect 9082 9476 9128 9514
rect 9082 9442 9088 9476
rect 9122 9442 9128 9476
rect 9082 9404 9128 9442
rect 9082 9370 9088 9404
rect 9122 9370 9128 9404
rect 9082 9332 9128 9370
rect 9082 9298 9088 9332
rect 9122 9298 9128 9332
rect 9082 9260 9128 9298
rect 9082 9226 9088 9260
rect 9122 9226 9128 9260
rect 9082 9188 9128 9226
rect 9082 9154 9088 9188
rect 9122 9154 9128 9188
rect 9082 9116 9128 9154
rect 9082 9082 9088 9116
rect 9122 9082 9128 9116
rect 9082 9044 9128 9082
rect 9082 9010 9088 9044
rect 9122 9010 9128 9044
rect 9082 8972 9128 9010
rect 9082 8938 9088 8972
rect 9122 8938 9128 8972
rect 9082 8900 9128 8938
rect 9082 8866 9088 8900
rect 9122 8866 9128 8900
rect 9082 8828 9128 8866
rect 9082 8794 9088 8828
rect 9122 8794 9128 8828
rect 9082 8756 9128 8794
rect 9082 8722 9088 8756
rect 9122 8722 9128 8756
rect 9082 8684 9128 8722
rect 9082 8650 9088 8684
rect 9122 8650 9128 8684
rect 9082 8612 9128 8650
rect 9082 8578 9088 8612
rect 9122 8578 9128 8612
rect 9082 8540 9128 8578
rect 9082 8506 9088 8540
rect 9122 8506 9128 8540
rect 9082 8468 9128 8506
rect 9082 8434 9088 8468
rect 9122 8434 9128 8468
rect 9082 8396 9128 8434
rect 9082 8362 9088 8396
rect 9122 8362 9128 8396
rect 9082 8324 9128 8362
rect 9082 8290 9088 8324
rect 9122 8290 9128 8324
rect 9082 8252 9128 8290
rect 9082 8218 9088 8252
rect 9122 8218 9128 8252
rect 9082 8180 9128 8218
rect 9082 8146 9088 8180
rect 9122 8146 9128 8180
rect 9082 8108 9128 8146
rect 9082 8074 9088 8108
rect 9122 8074 9128 8108
rect 9082 8036 9128 8074
rect 9082 8002 9088 8036
rect 9122 8002 9128 8036
rect 9082 7964 9128 8002
rect 9082 7930 9088 7964
rect 9122 7930 9128 7964
rect 9082 7892 9128 7930
rect 9082 7858 9088 7892
rect 9122 7858 9128 7892
rect 9082 7820 9128 7858
rect 9082 7786 9088 7820
rect 9122 7786 9128 7820
rect 9082 7748 9128 7786
rect 9082 7714 9088 7748
rect 9122 7714 9128 7748
rect 9082 7676 9128 7714
rect 9082 7642 9088 7676
rect 9122 7642 9128 7676
rect 9082 7604 9128 7642
rect 9082 7570 9088 7604
rect 9122 7570 9128 7604
rect 9082 7532 9128 7570
rect 9082 7498 9088 7532
rect 9122 7498 9128 7532
rect 9082 7460 9128 7498
rect 9082 7426 9088 7460
rect 9122 7426 9128 7460
rect 9082 7388 9128 7426
rect 9082 7354 9088 7388
rect 9122 7354 9128 7388
rect 9082 7316 9128 7354
rect 9082 7282 9088 7316
rect 9122 7282 9128 7316
rect 9082 7244 9128 7282
rect 9082 7210 9088 7244
rect 9122 7210 9128 7244
rect 9082 7172 9128 7210
rect 9082 7138 9088 7172
rect 9122 7138 9128 7172
rect 9082 7100 9128 7138
rect 9082 7066 9088 7100
rect 9122 7066 9128 7100
rect 9082 7028 9128 7066
rect 9082 6994 9088 7028
rect 9122 6994 9128 7028
rect 9082 6956 9128 6994
rect 9082 6922 9088 6956
rect 9122 6922 9128 6956
rect 9082 6884 9128 6922
rect 9082 6850 9088 6884
rect 9122 6850 9128 6884
rect 9082 6812 9128 6850
rect 9082 6778 9088 6812
rect 9122 6778 9128 6812
rect 9082 6740 9128 6778
rect 9082 6706 9088 6740
rect 9122 6706 9128 6740
rect 9082 6668 9128 6706
rect 9082 6634 9088 6668
rect 9122 6634 9128 6668
rect 9082 6596 9128 6634
rect 9082 6562 9088 6596
rect 9122 6562 9128 6596
rect 9082 6524 9128 6562
rect 9082 6490 9088 6524
rect 9122 6490 9128 6524
rect 9082 6452 9128 6490
rect 9082 6418 9088 6452
rect 9122 6418 9128 6452
rect 9082 6380 9128 6418
rect 9082 6346 9088 6380
rect 9122 6346 9128 6380
rect 9082 6308 9128 6346
rect 9082 6274 9088 6308
rect 9122 6274 9128 6308
rect 9082 6236 9128 6274
rect 9082 6202 9088 6236
rect 9122 6202 9128 6236
rect 9082 6164 9128 6202
rect 9082 6130 9088 6164
rect 9122 6130 9128 6164
rect 9082 6092 9128 6130
rect 9082 6058 9088 6092
rect 9122 6058 9128 6092
rect 9082 6020 9128 6058
rect 9082 5986 9088 6020
rect 9122 5986 9128 6020
rect 9082 5948 9128 5986
rect 9082 5914 9088 5948
rect 9122 5914 9128 5948
rect 9082 5876 9128 5914
rect 9082 5842 9088 5876
rect 9122 5842 9128 5876
rect 9082 5804 9128 5842
rect 9082 5770 9088 5804
rect 9122 5770 9128 5804
rect 9082 5732 9128 5770
rect 9082 5698 9088 5732
rect 9122 5698 9128 5732
rect 9082 5660 9128 5698
rect 9082 5626 9088 5660
rect 9122 5626 9128 5660
rect 9082 5588 9128 5626
rect 9082 5554 9088 5588
rect 9122 5554 9128 5588
rect 9082 5516 9128 5554
rect 9082 5482 9088 5516
rect 9122 5482 9128 5516
rect 9082 5444 9128 5482
rect 9082 5410 9088 5444
rect 9122 5410 9128 5444
rect 9082 5372 9128 5410
rect 9082 5338 9088 5372
rect 9122 5338 9128 5372
rect 9082 5300 9128 5338
rect 9082 5266 9088 5300
rect 9122 5266 9128 5300
rect 9082 5228 9128 5266
rect 9082 5194 9088 5228
rect 9122 5194 9128 5228
rect 9082 5156 9128 5194
rect 9082 5122 9088 5156
rect 9122 5122 9128 5156
rect 9082 5084 9128 5122
rect 9082 5050 9088 5084
rect 9122 5050 9128 5084
rect 9082 5012 9128 5050
rect 9082 4978 9088 5012
rect 9122 4978 9128 5012
rect 9082 4940 9128 4978
rect 9082 4906 9088 4940
rect 9122 4906 9128 4940
rect 9082 4868 9128 4906
rect 9082 4834 9088 4868
rect 9122 4834 9128 4868
rect 9082 4796 9128 4834
rect 9082 4762 9088 4796
rect 9122 4762 9128 4796
rect 9082 4724 9128 4762
rect 9082 4690 9088 4724
rect 9122 4690 9128 4724
rect 9082 4652 9128 4690
rect 9082 4618 9088 4652
rect 9122 4618 9128 4652
rect 9082 4580 9128 4618
rect 9082 4546 9088 4580
rect 9122 4546 9128 4580
rect 9082 4508 9128 4546
rect 9082 4474 9088 4508
rect 9122 4474 9128 4508
rect 9082 4436 9128 4474
rect 9082 4402 9088 4436
rect 9122 4402 9128 4436
rect 9082 4364 9128 4402
rect 9082 4330 9088 4364
rect 9122 4330 9128 4364
rect 9082 4292 9128 4330
rect 9082 4258 9088 4292
rect 9122 4258 9128 4292
rect 9082 4220 9128 4258
rect 9082 4186 9088 4220
rect 9122 4186 9128 4220
rect 9082 4148 9128 4186
rect 9082 4114 9088 4148
rect 9122 4114 9128 4148
rect 9082 4076 9128 4114
rect 9082 4042 9088 4076
rect 9122 4042 9128 4076
rect 9082 4004 9128 4042
rect 9082 3970 9088 4004
rect 9122 3970 9128 4004
rect 9082 3932 9128 3970
rect 9082 3898 9088 3932
rect 9122 3898 9128 3932
rect 9082 3860 9128 3898
rect 9082 3826 9088 3860
rect 9122 3826 9128 3860
rect 9082 3788 9128 3826
rect 9082 3754 9088 3788
rect 9122 3754 9128 3788
rect 9082 3716 9128 3754
rect 9082 3682 9088 3716
rect 9122 3682 9128 3716
rect 9082 3644 9128 3682
rect 9082 3610 9088 3644
rect 9122 3610 9128 3644
rect 9082 3572 9128 3610
rect 9082 3538 9088 3572
rect 9122 3538 9128 3572
rect 9082 3500 9128 3538
rect 9082 3466 9088 3500
rect 9122 3466 9128 3500
rect 10220 38650 10226 38684
rect 10260 38650 10266 38684
tri 10266 38682 10268 38684 nw
tri 11416 38682 11418 38684 ne
rect 10220 38611 10266 38650
rect 10220 38577 10226 38611
rect 10260 38577 10266 38611
rect 10220 38538 10266 38577
rect 10220 38504 10226 38538
rect 10260 38504 10266 38538
rect 10220 38465 10266 38504
rect 10220 38431 10226 38465
rect 10260 38431 10266 38465
rect 10220 38392 10266 38431
rect 10220 38358 10226 38392
rect 10260 38358 10266 38392
rect 10220 38319 10266 38358
rect 10220 38285 10226 38319
rect 10260 38285 10266 38319
rect 10220 38246 10266 38285
rect 10220 38212 10226 38246
rect 10260 38212 10266 38246
rect 10220 38173 10266 38212
rect 10220 38139 10226 38173
rect 10260 38139 10266 38173
rect 10220 38100 10266 38139
rect 10220 38066 10226 38100
rect 10260 38066 10266 38100
rect 10220 38027 10266 38066
rect 10220 37993 10226 38027
rect 10260 37993 10266 38027
rect 10220 37954 10266 37993
rect 10220 37920 10226 37954
rect 10260 37920 10266 37954
rect 10220 37881 10266 37920
rect 10220 37847 10226 37881
rect 10260 37847 10266 37881
rect 10220 37808 10266 37847
rect 10220 37774 10226 37808
rect 10260 37774 10266 37808
rect 10220 37735 10266 37774
rect 10220 37701 10226 37735
rect 10260 37701 10266 37735
rect 10220 37662 10266 37701
rect 10220 37628 10226 37662
rect 10260 37628 10266 37662
rect 10220 37589 10266 37628
rect 10220 37555 10226 37589
rect 10260 37555 10266 37589
rect 10220 37516 10266 37555
rect 10220 37482 10226 37516
rect 10260 37482 10266 37516
rect 10220 37443 10266 37482
rect 10220 37409 10226 37443
rect 10260 37409 10266 37443
rect 10220 37370 10266 37409
rect 10220 37336 10226 37370
rect 10260 37336 10266 37370
rect 10220 37297 10266 37336
rect 10220 37263 10226 37297
rect 10260 37263 10266 37297
rect 10220 37224 10266 37263
rect 10220 37190 10226 37224
rect 10260 37190 10266 37224
rect 10220 37151 10266 37190
rect 10220 37117 10226 37151
rect 10260 37117 10266 37151
rect 10220 37078 10266 37117
rect 10220 37044 10226 37078
rect 10260 37044 10266 37078
rect 10220 37005 10266 37044
rect 10220 36971 10226 37005
rect 10260 36971 10266 37005
rect 10220 36932 10266 36971
rect 10220 36898 10226 36932
rect 10260 36898 10266 36932
rect 10220 36859 10266 36898
rect 10220 36825 10226 36859
rect 10260 36825 10266 36859
rect 10220 36786 10266 36825
rect 10220 36752 10226 36786
rect 10260 36752 10266 36786
rect 10220 36713 10266 36752
rect 10220 36679 10226 36713
rect 10260 36679 10266 36713
rect 10220 36640 10266 36679
rect 10220 36606 10226 36640
rect 10260 36606 10266 36640
rect 10220 36567 10266 36606
rect 10220 36533 10226 36567
rect 10260 36533 10266 36567
rect 10220 36494 10266 36533
rect 10220 36460 10226 36494
rect 10260 36460 10266 36494
rect 10220 36421 10266 36460
rect 10220 36387 10226 36421
rect 10260 36387 10266 36421
rect 10220 36348 10266 36387
rect 10220 36314 10226 36348
rect 10260 36314 10266 36348
rect 10220 36275 10266 36314
rect 10220 36241 10226 36275
rect 10260 36241 10266 36275
rect 10220 36202 10266 36241
rect 10220 36168 10226 36202
rect 10260 36168 10266 36202
rect 10220 36129 10266 36168
rect 10220 36095 10226 36129
rect 10260 36095 10266 36129
rect 10220 36056 10266 36095
rect 10220 36022 10226 36056
rect 10260 36022 10266 36056
rect 10220 35983 10266 36022
rect 10220 35949 10226 35983
rect 10260 35949 10266 35983
rect 10220 35910 10266 35949
rect 10220 35876 10226 35910
rect 10260 35876 10266 35910
rect 10220 35837 10266 35876
rect 10220 35803 10226 35837
rect 10260 35803 10266 35837
rect 10220 35764 10266 35803
rect 10220 35730 10226 35764
rect 10260 35730 10266 35764
rect 10220 35691 10266 35730
rect 10220 35657 10226 35691
rect 10260 35657 10266 35691
rect 10220 35618 10266 35657
rect 10220 35584 10226 35618
rect 10260 35584 10266 35618
rect 10220 35545 10266 35584
rect 10220 35511 10226 35545
rect 10260 35511 10266 35545
rect 10220 35472 10266 35511
rect 10220 35438 10226 35472
rect 10260 35438 10266 35472
rect 10220 35399 10266 35438
rect 10220 35365 10226 35399
rect 10260 35365 10266 35399
rect 10220 35326 10266 35365
rect 10220 35292 10226 35326
rect 10260 35292 10266 35326
rect 10220 35253 10266 35292
rect 10220 35219 10226 35253
rect 10260 35219 10266 35253
rect 10220 35180 10266 35219
rect 10220 35146 10226 35180
rect 10260 35146 10266 35180
rect 10220 35108 10266 35146
rect 10220 35074 10226 35108
rect 10260 35074 10266 35108
rect 10220 35036 10266 35074
rect 10220 35002 10226 35036
rect 10260 35002 10266 35036
rect 10220 34964 10266 35002
rect 10220 34930 10226 34964
rect 10260 34930 10266 34964
rect 10220 34892 10266 34930
rect 10220 34858 10226 34892
rect 10260 34858 10266 34892
rect 10220 34820 10266 34858
rect 10220 34786 10226 34820
rect 10260 34786 10266 34820
rect 10220 34748 10266 34786
rect 10220 34714 10226 34748
rect 10260 34714 10266 34748
rect 10220 34676 10266 34714
rect 10220 34642 10226 34676
rect 10260 34642 10266 34676
rect 10220 34604 10266 34642
rect 10220 34570 10226 34604
rect 10260 34570 10266 34604
rect 10220 34532 10266 34570
rect 10220 34498 10226 34532
rect 10260 34498 10266 34532
rect 10220 34460 10266 34498
rect 10220 34426 10226 34460
rect 10260 34426 10266 34460
rect 10220 34388 10266 34426
rect 10220 34354 10226 34388
rect 10260 34354 10266 34388
rect 10220 34316 10266 34354
rect 10220 34282 10226 34316
rect 10260 34282 10266 34316
rect 10220 34244 10266 34282
rect 10220 34210 10226 34244
rect 10260 34210 10266 34244
rect 10220 34172 10266 34210
rect 10220 34138 10226 34172
rect 10260 34138 10266 34172
rect 10220 34100 10266 34138
rect 10220 34066 10226 34100
rect 10260 34066 10266 34100
rect 10220 34028 10266 34066
rect 10220 33994 10226 34028
rect 10260 33994 10266 34028
rect 10220 33956 10266 33994
rect 10220 33922 10226 33956
rect 10260 33922 10266 33956
rect 10220 33884 10266 33922
rect 10220 33850 10226 33884
rect 10260 33850 10266 33884
rect 10220 33812 10266 33850
rect 10220 33778 10226 33812
rect 10260 33778 10266 33812
rect 10220 33740 10266 33778
rect 10220 33706 10226 33740
rect 10260 33706 10266 33740
rect 10220 33668 10266 33706
rect 10220 33634 10226 33668
rect 10260 33634 10266 33668
rect 10220 33596 10266 33634
rect 10220 33562 10226 33596
rect 10260 33562 10266 33596
rect 10220 33524 10266 33562
rect 10220 33490 10226 33524
rect 10260 33490 10266 33524
rect 10220 33452 10266 33490
rect 10220 33418 10226 33452
rect 10260 33418 10266 33452
rect 10220 33380 10266 33418
rect 10220 33346 10226 33380
rect 10260 33346 10266 33380
rect 10220 33308 10266 33346
rect 10220 33274 10226 33308
rect 10260 33274 10266 33308
rect 10220 33236 10266 33274
rect 10220 33202 10226 33236
rect 10260 33202 10266 33236
rect 10220 33164 10266 33202
rect 10220 33130 10226 33164
rect 10260 33130 10266 33164
rect 10220 33092 10266 33130
rect 10220 33058 10226 33092
rect 10260 33058 10266 33092
rect 10220 33020 10266 33058
rect 10220 32986 10226 33020
rect 10260 32986 10266 33020
rect 10220 32948 10266 32986
rect 10220 32914 10226 32948
rect 10260 32914 10266 32948
rect 10220 32876 10266 32914
rect 10220 32842 10226 32876
rect 10260 32842 10266 32876
rect 10220 32804 10266 32842
rect 10220 32770 10226 32804
rect 10260 32770 10266 32804
rect 10220 32732 10266 32770
rect 10220 32698 10226 32732
rect 10260 32698 10266 32732
rect 10220 32660 10266 32698
rect 10220 32626 10226 32660
rect 10260 32626 10266 32660
rect 10220 32588 10266 32626
rect 10220 32554 10226 32588
rect 10260 32554 10266 32588
rect 10220 32516 10266 32554
rect 10220 32482 10226 32516
rect 10260 32482 10266 32516
rect 10220 32444 10266 32482
rect 10220 32410 10226 32444
rect 10260 32410 10266 32444
rect 10220 32372 10266 32410
rect 10220 32338 10226 32372
rect 10260 32338 10266 32372
rect 10220 32300 10266 32338
rect 10220 32266 10226 32300
rect 10260 32266 10266 32300
rect 10220 32228 10266 32266
rect 10220 32194 10226 32228
rect 10260 32194 10266 32228
rect 10220 32156 10266 32194
rect 10220 32122 10226 32156
rect 10260 32122 10266 32156
rect 10220 32084 10266 32122
rect 10220 32050 10226 32084
rect 10260 32050 10266 32084
rect 10220 32012 10266 32050
rect 10220 31978 10226 32012
rect 10260 31978 10266 32012
rect 10220 31940 10266 31978
rect 10220 31906 10226 31940
rect 10260 31906 10266 31940
rect 10220 31868 10266 31906
rect 10220 31834 10226 31868
rect 10260 31834 10266 31868
rect 10220 31796 10266 31834
rect 10220 31762 10226 31796
rect 10260 31762 10266 31796
rect 10220 31724 10266 31762
rect 10220 31690 10226 31724
rect 10260 31690 10266 31724
rect 10220 31652 10266 31690
rect 10220 31618 10226 31652
rect 10260 31618 10266 31652
rect 10220 31580 10266 31618
rect 10220 31546 10226 31580
rect 10260 31546 10266 31580
rect 10220 31508 10266 31546
rect 10220 31474 10226 31508
rect 10260 31474 10266 31508
rect 10220 31436 10266 31474
rect 10220 31402 10226 31436
rect 10260 31402 10266 31436
rect 10220 31364 10266 31402
rect 10220 31330 10226 31364
rect 10260 31330 10266 31364
rect 10220 31292 10266 31330
rect 10220 31258 10226 31292
rect 10260 31258 10266 31292
rect 10220 31220 10266 31258
rect 10220 31186 10226 31220
rect 10260 31186 10266 31220
rect 10220 31148 10266 31186
rect 10220 31114 10226 31148
rect 10260 31114 10266 31148
rect 10220 31076 10266 31114
rect 10220 31042 10226 31076
rect 10260 31042 10266 31076
rect 10220 31004 10266 31042
rect 10220 30970 10226 31004
rect 10260 30970 10266 31004
rect 10220 30932 10266 30970
rect 10220 30898 10226 30932
rect 10260 30898 10266 30932
rect 10220 30860 10266 30898
rect 10220 30826 10226 30860
rect 10260 30826 10266 30860
rect 10220 30788 10266 30826
rect 10220 30754 10226 30788
rect 10260 30754 10266 30788
rect 10220 30716 10266 30754
rect 10220 30682 10226 30716
rect 10260 30682 10266 30716
rect 10220 30644 10266 30682
rect 10220 30610 10226 30644
rect 10260 30610 10266 30644
rect 10220 30572 10266 30610
rect 10220 30538 10226 30572
rect 10260 30538 10266 30572
rect 10220 30500 10266 30538
rect 10220 30466 10226 30500
rect 10260 30466 10266 30500
rect 10220 30428 10266 30466
rect 10220 30394 10226 30428
rect 10260 30394 10266 30428
rect 10220 30356 10266 30394
rect 10220 30322 10226 30356
rect 10260 30322 10266 30356
rect 10220 30284 10266 30322
rect 10220 30250 10226 30284
rect 10260 30250 10266 30284
rect 10220 30212 10266 30250
rect 10220 30178 10226 30212
rect 10260 30178 10266 30212
rect 10220 30140 10266 30178
rect 10220 30106 10226 30140
rect 10260 30106 10266 30140
rect 10220 30068 10266 30106
rect 10220 30034 10226 30068
rect 10260 30034 10266 30068
rect 10220 29996 10266 30034
rect 10220 29962 10226 29996
rect 10260 29962 10266 29996
rect 10220 29924 10266 29962
rect 10220 29890 10226 29924
rect 10260 29890 10266 29924
rect 10220 29852 10266 29890
rect 10220 29818 10226 29852
rect 10260 29818 10266 29852
rect 10220 29780 10266 29818
rect 10220 29746 10226 29780
rect 10260 29746 10266 29780
rect 10220 29708 10266 29746
rect 10220 29674 10226 29708
rect 10260 29674 10266 29708
rect 10220 29636 10266 29674
rect 10220 29602 10226 29636
rect 10260 29602 10266 29636
rect 10220 29564 10266 29602
rect 10220 29530 10226 29564
rect 10260 29530 10266 29564
rect 10220 29492 10266 29530
rect 10220 29458 10226 29492
rect 10260 29458 10266 29492
rect 10220 29420 10266 29458
rect 10220 29386 10226 29420
rect 10260 29386 10266 29420
rect 10220 29348 10266 29386
rect 10220 29314 10226 29348
rect 10260 29314 10266 29348
rect 10220 29276 10266 29314
rect 10220 29242 10226 29276
rect 10260 29242 10266 29276
rect 10220 29204 10266 29242
rect 10220 29170 10226 29204
rect 10260 29170 10266 29204
rect 10220 29132 10266 29170
rect 10220 29098 10226 29132
rect 10260 29098 10266 29132
rect 10220 29060 10266 29098
rect 10220 29026 10226 29060
rect 10260 29026 10266 29060
rect 10220 28988 10266 29026
rect 10220 28954 10226 28988
rect 10260 28954 10266 28988
rect 10220 28916 10266 28954
rect 10220 28882 10226 28916
rect 10260 28882 10266 28916
rect 10220 28844 10266 28882
rect 10220 28810 10226 28844
rect 10260 28810 10266 28844
rect 10220 28772 10266 28810
rect 10220 28738 10226 28772
rect 10260 28738 10266 28772
rect 10220 28700 10266 28738
rect 10220 28666 10226 28700
rect 10260 28666 10266 28700
rect 10220 28628 10266 28666
rect 10220 28594 10226 28628
rect 10260 28594 10266 28628
rect 10220 28556 10266 28594
rect 10220 28522 10226 28556
rect 10260 28522 10266 28556
rect 10220 28484 10266 28522
rect 10220 28450 10226 28484
rect 10260 28450 10266 28484
rect 10220 28412 10266 28450
rect 10220 28378 10226 28412
rect 10260 28378 10266 28412
rect 10220 28340 10266 28378
rect 10220 28306 10226 28340
rect 10260 28306 10266 28340
rect 10220 28268 10266 28306
rect 10220 28234 10226 28268
rect 10260 28234 10266 28268
rect 10220 28196 10266 28234
rect 10220 28162 10226 28196
rect 10260 28162 10266 28196
rect 10220 28124 10266 28162
rect 10220 28090 10226 28124
rect 10260 28090 10266 28124
rect 10220 28052 10266 28090
rect 10220 28018 10226 28052
rect 10260 28018 10266 28052
rect 10220 27980 10266 28018
rect 10220 27946 10226 27980
rect 10260 27946 10266 27980
rect 10220 27908 10266 27946
rect 10220 27874 10226 27908
rect 10260 27874 10266 27908
rect 10220 27836 10266 27874
rect 10220 27802 10226 27836
rect 10260 27802 10266 27836
rect 10220 27764 10266 27802
rect 10220 27730 10226 27764
rect 10260 27730 10266 27764
rect 10220 27692 10266 27730
rect 10220 27658 10226 27692
rect 10260 27658 10266 27692
rect 10220 27620 10266 27658
rect 10220 27586 10226 27620
rect 10260 27586 10266 27620
rect 10220 27548 10266 27586
rect 10220 27514 10226 27548
rect 10260 27514 10266 27548
rect 10220 27476 10266 27514
rect 10220 27442 10226 27476
rect 10260 27442 10266 27476
rect 10220 27404 10266 27442
rect 10220 27370 10226 27404
rect 10260 27370 10266 27404
rect 10220 27332 10266 27370
rect 10220 27298 10226 27332
rect 10260 27298 10266 27332
rect 10220 27260 10266 27298
rect 10220 27226 10226 27260
rect 10260 27226 10266 27260
rect 10220 27188 10266 27226
rect 10220 27154 10226 27188
rect 10260 27154 10266 27188
rect 10220 27116 10266 27154
rect 10220 27082 10226 27116
rect 10260 27082 10266 27116
rect 10220 27044 10266 27082
rect 10220 27010 10226 27044
rect 10260 27010 10266 27044
rect 10220 26972 10266 27010
rect 10220 26938 10226 26972
rect 10260 26938 10266 26972
rect 10220 26900 10266 26938
rect 10220 26866 10226 26900
rect 10260 26866 10266 26900
rect 10220 26828 10266 26866
rect 10220 26794 10226 26828
rect 10260 26794 10266 26828
rect 10220 26756 10266 26794
rect 10220 26722 10226 26756
rect 10260 26722 10266 26756
rect 10220 26684 10266 26722
rect 10220 26650 10226 26684
rect 10260 26650 10266 26684
rect 10220 26612 10266 26650
rect 10220 26578 10226 26612
rect 10260 26578 10266 26612
rect 10220 26540 10266 26578
rect 10220 26506 10226 26540
rect 10260 26506 10266 26540
rect 10220 26468 10266 26506
rect 10220 26434 10226 26468
rect 10260 26434 10266 26468
rect 10220 26396 10266 26434
rect 10220 26362 10226 26396
rect 10260 26362 10266 26396
rect 10220 26324 10266 26362
rect 10220 26290 10226 26324
rect 10260 26290 10266 26324
rect 10220 26252 10266 26290
rect 10220 26218 10226 26252
rect 10260 26218 10266 26252
rect 10220 26180 10266 26218
rect 10220 26146 10226 26180
rect 10260 26146 10266 26180
rect 10220 26108 10266 26146
rect 10220 26074 10226 26108
rect 10260 26074 10266 26108
rect 10220 26036 10266 26074
rect 10220 26002 10226 26036
rect 10260 26002 10266 26036
rect 10220 25964 10266 26002
rect 10220 25930 10226 25964
rect 10260 25930 10266 25964
rect 10220 25892 10266 25930
rect 10220 25858 10226 25892
rect 10260 25858 10266 25892
rect 10220 25820 10266 25858
rect 10220 25786 10226 25820
rect 10260 25786 10266 25820
rect 10220 25748 10266 25786
rect 10220 25714 10226 25748
rect 10260 25714 10266 25748
rect 10220 25676 10266 25714
rect 10220 25642 10226 25676
rect 10260 25642 10266 25676
rect 10220 25604 10266 25642
rect 10220 25570 10226 25604
rect 10260 25570 10266 25604
rect 10220 25532 10266 25570
rect 10220 25498 10226 25532
rect 10260 25498 10266 25532
rect 10220 25460 10266 25498
rect 10220 25426 10226 25460
rect 10260 25426 10266 25460
rect 10220 25388 10266 25426
rect 10220 25354 10226 25388
rect 10260 25354 10266 25388
rect 10220 25316 10266 25354
rect 10220 25282 10226 25316
rect 10260 25282 10266 25316
rect 10220 25244 10266 25282
rect 10220 25210 10226 25244
rect 10260 25210 10266 25244
rect 10220 25172 10266 25210
rect 10220 25138 10226 25172
rect 10260 25138 10266 25172
rect 10220 25100 10266 25138
rect 10220 25066 10226 25100
rect 10260 25066 10266 25100
rect 10220 25028 10266 25066
rect 10220 24994 10226 25028
rect 10260 24994 10266 25028
rect 10220 24956 10266 24994
rect 10220 24922 10226 24956
rect 10260 24922 10266 24956
rect 10220 24884 10266 24922
rect 10220 24850 10226 24884
rect 10260 24850 10266 24884
rect 10220 24812 10266 24850
rect 10220 24778 10226 24812
rect 10260 24778 10266 24812
rect 10220 24740 10266 24778
rect 10220 24706 10226 24740
rect 10260 24706 10266 24740
rect 10220 24668 10266 24706
rect 10220 24634 10226 24668
rect 10260 24634 10266 24668
rect 10220 24596 10266 24634
rect 10220 24562 10226 24596
rect 10260 24562 10266 24596
rect 10220 24524 10266 24562
rect 10220 24490 10226 24524
rect 10260 24490 10266 24524
rect 10220 24452 10266 24490
rect 10220 24418 10226 24452
rect 10260 24418 10266 24452
rect 10220 24380 10266 24418
rect 10220 24346 10226 24380
rect 10260 24346 10266 24380
rect 10220 24308 10266 24346
rect 10220 24274 10226 24308
rect 10260 24274 10266 24308
rect 10220 24236 10266 24274
rect 10220 24202 10226 24236
rect 10260 24202 10266 24236
rect 10220 24164 10266 24202
rect 10220 24130 10226 24164
rect 10260 24130 10266 24164
rect 10220 24092 10266 24130
rect 10220 24058 10226 24092
rect 10260 24058 10266 24092
rect 10220 24020 10266 24058
rect 10220 23986 10226 24020
rect 10260 23986 10266 24020
rect 10220 23948 10266 23986
rect 10220 23914 10226 23948
rect 10260 23914 10266 23948
rect 10220 23876 10266 23914
rect 10220 23842 10226 23876
rect 10260 23842 10266 23876
rect 10220 23804 10266 23842
rect 10220 23770 10226 23804
rect 10260 23770 10266 23804
rect 10220 23732 10266 23770
rect 10220 23698 10226 23732
rect 10260 23698 10266 23732
rect 10220 23660 10266 23698
rect 10220 23626 10226 23660
rect 10260 23626 10266 23660
rect 10220 23588 10266 23626
rect 10220 23554 10226 23588
rect 10260 23554 10266 23588
rect 10220 23516 10266 23554
rect 10220 23482 10226 23516
rect 10260 23482 10266 23516
rect 10220 23444 10266 23482
rect 10220 23410 10226 23444
rect 10260 23410 10266 23444
rect 10220 23372 10266 23410
rect 10220 23338 10226 23372
rect 10260 23338 10266 23372
rect 10220 23300 10266 23338
rect 10220 23266 10226 23300
rect 10260 23266 10266 23300
rect 10220 23228 10266 23266
rect 10220 23194 10226 23228
rect 10260 23194 10266 23228
rect 10220 23156 10266 23194
rect 10220 23122 10226 23156
rect 10260 23122 10266 23156
rect 10220 23084 10266 23122
rect 10220 23050 10226 23084
rect 10260 23050 10266 23084
rect 10220 23012 10266 23050
rect 10220 22978 10226 23012
rect 10260 22978 10266 23012
rect 10220 22940 10266 22978
rect 10220 22906 10226 22940
rect 10260 22906 10266 22940
rect 10220 22868 10266 22906
rect 10220 22834 10226 22868
rect 10260 22834 10266 22868
rect 10220 22796 10266 22834
rect 10220 22762 10226 22796
rect 10260 22762 10266 22796
rect 10220 22724 10266 22762
rect 10220 22690 10226 22724
rect 10260 22690 10266 22724
rect 10220 22652 10266 22690
rect 10220 22618 10226 22652
rect 10260 22618 10266 22652
rect 10220 22580 10266 22618
rect 10220 22546 10226 22580
rect 10260 22546 10266 22580
rect 10220 22508 10266 22546
rect 10220 22474 10226 22508
rect 10260 22474 10266 22508
rect 10220 22436 10266 22474
rect 10220 22402 10226 22436
rect 10260 22402 10266 22436
rect 10220 22364 10266 22402
rect 10220 22330 10226 22364
rect 10260 22330 10266 22364
rect 10220 22292 10266 22330
rect 10220 22258 10226 22292
rect 10260 22258 10266 22292
rect 10220 22220 10266 22258
rect 10220 22186 10226 22220
rect 10260 22186 10266 22220
rect 10220 22148 10266 22186
rect 10220 22114 10226 22148
rect 10260 22114 10266 22148
rect 10220 22076 10266 22114
rect 10220 22042 10226 22076
rect 10260 22042 10266 22076
rect 10220 22004 10266 22042
rect 10220 21970 10226 22004
rect 10260 21970 10266 22004
rect 10220 21932 10266 21970
rect 10220 21898 10226 21932
rect 10260 21898 10266 21932
rect 10220 21860 10266 21898
rect 10220 21826 10226 21860
rect 10260 21826 10266 21860
rect 10220 21788 10266 21826
rect 10220 21754 10226 21788
rect 10260 21754 10266 21788
rect 10220 21716 10266 21754
rect 10220 21682 10226 21716
rect 10260 21682 10266 21716
rect 10220 21644 10266 21682
rect 10220 21610 10226 21644
rect 10260 21610 10266 21644
rect 10220 21572 10266 21610
rect 10220 21538 10226 21572
rect 10260 21538 10266 21572
rect 10220 21500 10266 21538
rect 10220 21466 10226 21500
rect 10260 21466 10266 21500
rect 10220 21428 10266 21466
rect 10220 21394 10226 21428
rect 10260 21394 10266 21428
rect 10220 21356 10266 21394
rect 10220 21322 10226 21356
rect 10260 21322 10266 21356
rect 10220 21284 10266 21322
rect 10220 21250 10226 21284
rect 10260 21250 10266 21284
rect 10220 21212 10266 21250
rect 10220 21178 10226 21212
rect 10260 21178 10266 21212
rect 10220 21140 10266 21178
rect 10220 21106 10226 21140
rect 10260 21106 10266 21140
rect 10220 21068 10266 21106
rect 10220 21034 10226 21068
rect 10260 21034 10266 21068
rect 10220 20996 10266 21034
rect 10220 20962 10226 20996
rect 10260 20962 10266 20996
rect 10220 20924 10266 20962
rect 10220 20890 10226 20924
rect 10260 20890 10266 20924
rect 10220 20852 10266 20890
rect 10220 20818 10226 20852
rect 10260 20818 10266 20852
rect 10220 20780 10266 20818
rect 10220 20746 10226 20780
rect 10260 20746 10266 20780
rect 10220 20708 10266 20746
rect 10220 20674 10226 20708
rect 10260 20674 10266 20708
rect 10220 20636 10266 20674
rect 10220 20602 10226 20636
rect 10260 20602 10266 20636
rect 10220 20564 10266 20602
rect 10220 20530 10226 20564
rect 10260 20530 10266 20564
rect 10220 20492 10266 20530
rect 10220 20458 10226 20492
rect 10260 20458 10266 20492
rect 10220 20420 10266 20458
rect 10220 20386 10226 20420
rect 10260 20386 10266 20420
rect 10220 20348 10266 20386
rect 10220 20314 10226 20348
rect 10260 20314 10266 20348
rect 10220 20276 10266 20314
rect 10220 20242 10226 20276
rect 10260 20242 10266 20276
rect 10220 20204 10266 20242
rect 10220 20170 10226 20204
rect 10260 20170 10266 20204
rect 10220 20132 10266 20170
rect 10220 20098 10226 20132
rect 10260 20098 10266 20132
rect 10220 20060 10266 20098
rect 10220 20026 10226 20060
rect 10260 20026 10266 20060
rect 10220 19988 10266 20026
rect 10220 19954 10226 19988
rect 10260 19954 10266 19988
rect 10220 19916 10266 19954
rect 10220 19882 10226 19916
rect 10260 19882 10266 19916
rect 10220 19844 10266 19882
rect 10220 19810 10226 19844
rect 10260 19810 10266 19844
rect 10220 19772 10266 19810
rect 10220 19738 10226 19772
rect 10260 19738 10266 19772
rect 10220 19700 10266 19738
rect 10220 19666 10226 19700
rect 10260 19666 10266 19700
rect 10220 19628 10266 19666
rect 10220 19594 10226 19628
rect 10260 19594 10266 19628
rect 10220 19556 10266 19594
rect 10220 19522 10226 19556
rect 10260 19522 10266 19556
rect 10220 19484 10266 19522
rect 10220 19450 10226 19484
rect 10260 19450 10266 19484
rect 10220 19412 10266 19450
rect 10220 19378 10226 19412
rect 10260 19378 10266 19412
rect 10220 19340 10266 19378
rect 10220 19306 10226 19340
rect 10260 19306 10266 19340
rect 10220 19268 10266 19306
rect 10220 19234 10226 19268
rect 10260 19234 10266 19268
rect 10220 19196 10266 19234
rect 10220 19162 10226 19196
rect 10260 19162 10266 19196
rect 10220 19124 10266 19162
rect 10220 19090 10226 19124
rect 10260 19090 10266 19124
rect 10220 19052 10266 19090
rect 10220 19018 10226 19052
rect 10260 19018 10266 19052
rect 10220 18980 10266 19018
rect 10220 18946 10226 18980
rect 10260 18946 10266 18980
rect 10220 18908 10266 18946
rect 10220 18874 10226 18908
rect 10260 18874 10266 18908
rect 10220 18836 10266 18874
rect 10220 18802 10226 18836
rect 10260 18802 10266 18836
rect 10220 18764 10266 18802
rect 10220 18730 10226 18764
rect 10260 18730 10266 18764
rect 10220 18692 10266 18730
rect 10220 18658 10226 18692
rect 10260 18658 10266 18692
rect 10220 18620 10266 18658
rect 10220 18586 10226 18620
rect 10260 18586 10266 18620
rect 10220 18548 10266 18586
rect 10220 18514 10226 18548
rect 10260 18514 10266 18548
rect 10220 18476 10266 18514
rect 10220 18442 10226 18476
rect 10260 18442 10266 18476
rect 10220 18404 10266 18442
rect 10220 18370 10226 18404
rect 10260 18370 10266 18404
rect 10220 18332 10266 18370
rect 10220 18298 10226 18332
rect 10260 18298 10266 18332
rect 10220 18260 10266 18298
rect 10220 18226 10226 18260
rect 10260 18226 10266 18260
rect 10220 18188 10266 18226
rect 10220 18154 10226 18188
rect 10260 18154 10266 18188
rect 10220 18116 10266 18154
rect 10220 18082 10226 18116
rect 10260 18082 10266 18116
rect 10220 18044 10266 18082
rect 10220 18010 10226 18044
rect 10260 18010 10266 18044
rect 10220 17972 10266 18010
rect 10220 17938 10226 17972
rect 10260 17938 10266 17972
rect 10220 17900 10266 17938
rect 10220 17866 10226 17900
rect 10260 17866 10266 17900
rect 10220 17828 10266 17866
rect 10220 17794 10226 17828
rect 10260 17794 10266 17828
rect 10220 17756 10266 17794
rect 10220 17722 10226 17756
rect 10260 17722 10266 17756
rect 10220 17684 10266 17722
rect 10220 17650 10226 17684
rect 10260 17650 10266 17684
rect 10220 17612 10266 17650
rect 10220 17578 10226 17612
rect 10260 17578 10266 17612
rect 10220 17540 10266 17578
rect 10220 17506 10226 17540
rect 10260 17506 10266 17540
rect 10220 17468 10266 17506
rect 10220 17434 10226 17468
rect 10260 17434 10266 17468
rect 10220 17396 10266 17434
rect 10220 17362 10226 17396
rect 10260 17362 10266 17396
rect 10220 17324 10266 17362
rect 10220 17290 10226 17324
rect 10260 17290 10266 17324
rect 10220 17252 10266 17290
rect 10220 17218 10226 17252
rect 10260 17218 10266 17252
rect 10220 17180 10266 17218
rect 10220 17146 10226 17180
rect 10260 17146 10266 17180
rect 10220 17108 10266 17146
rect 10220 17074 10226 17108
rect 10260 17074 10266 17108
rect 10220 17036 10266 17074
rect 10220 17002 10226 17036
rect 10260 17002 10266 17036
rect 10220 16964 10266 17002
rect 10220 16930 10226 16964
rect 10260 16930 10266 16964
rect 10220 16892 10266 16930
rect 10220 16858 10226 16892
rect 10260 16858 10266 16892
rect 10220 16820 10266 16858
rect 10220 16786 10226 16820
rect 10260 16786 10266 16820
rect 10220 16748 10266 16786
rect 10220 16714 10226 16748
rect 10260 16714 10266 16748
rect 10220 16676 10266 16714
rect 10220 16642 10226 16676
rect 10260 16642 10266 16676
rect 10220 16604 10266 16642
rect 10220 16570 10226 16604
rect 10260 16570 10266 16604
rect 10220 16532 10266 16570
rect 10220 16498 10226 16532
rect 10260 16498 10266 16532
rect 10220 16460 10266 16498
rect 10220 16426 10226 16460
rect 10260 16426 10266 16460
rect 10220 16388 10266 16426
rect 10220 16354 10226 16388
rect 10260 16354 10266 16388
rect 10220 16316 10266 16354
rect 10220 16282 10226 16316
rect 10260 16282 10266 16316
rect 10220 16244 10266 16282
rect 10220 16210 10226 16244
rect 10260 16210 10266 16244
rect 10220 16172 10266 16210
rect 10220 16138 10226 16172
rect 10260 16138 10266 16172
rect 10220 16100 10266 16138
rect 10220 16066 10226 16100
rect 10260 16066 10266 16100
rect 10220 16028 10266 16066
rect 10220 15994 10226 16028
rect 10260 15994 10266 16028
rect 10220 15956 10266 15994
rect 10220 15922 10226 15956
rect 10260 15922 10266 15956
rect 10220 15884 10266 15922
rect 10220 15850 10226 15884
rect 10260 15850 10266 15884
rect 10220 15812 10266 15850
rect 10220 15778 10226 15812
rect 10260 15778 10266 15812
rect 10220 15740 10266 15778
rect 10220 15706 10226 15740
rect 10260 15706 10266 15740
rect 10220 15668 10266 15706
rect 10220 15634 10226 15668
rect 10260 15634 10266 15668
rect 10220 15596 10266 15634
rect 10220 15562 10226 15596
rect 10260 15562 10266 15596
rect 10220 15524 10266 15562
rect 10220 15490 10226 15524
rect 10260 15490 10266 15524
rect 10220 15452 10266 15490
rect 10220 15418 10226 15452
rect 10260 15418 10266 15452
rect 10220 15380 10266 15418
rect 10220 15346 10226 15380
rect 10260 15346 10266 15380
rect 10220 15308 10266 15346
rect 10220 15274 10226 15308
rect 10260 15274 10266 15308
rect 10220 15236 10266 15274
rect 10220 15202 10226 15236
rect 10260 15202 10266 15236
rect 10220 15164 10266 15202
rect 10220 15130 10226 15164
rect 10260 15130 10266 15164
rect 10220 15092 10266 15130
rect 10220 15058 10226 15092
rect 10260 15058 10266 15092
rect 10220 15020 10266 15058
rect 10220 14986 10226 15020
rect 10260 14986 10266 15020
rect 10220 14948 10266 14986
rect 10220 14914 10226 14948
rect 10260 14914 10266 14948
rect 10220 14876 10266 14914
rect 10220 14842 10226 14876
rect 10260 14842 10266 14876
rect 10220 14804 10266 14842
rect 10220 14770 10226 14804
rect 10260 14770 10266 14804
rect 10220 14732 10266 14770
rect 10220 14698 10226 14732
rect 10260 14698 10266 14732
rect 10220 14660 10266 14698
rect 10220 14626 10226 14660
rect 10260 14626 10266 14660
rect 10220 14588 10266 14626
rect 10220 14554 10226 14588
rect 10260 14554 10266 14588
rect 10220 14516 10266 14554
rect 10220 14482 10226 14516
rect 10260 14482 10266 14516
rect 10220 14444 10266 14482
rect 10220 14410 10226 14444
rect 10260 14410 10266 14444
rect 10220 14372 10266 14410
rect 10220 14338 10226 14372
rect 10260 14338 10266 14372
rect 10220 14300 10266 14338
rect 10220 14266 10226 14300
rect 10260 14266 10266 14300
rect 10220 14228 10266 14266
rect 10220 14194 10226 14228
rect 10260 14194 10266 14228
rect 10220 14156 10266 14194
rect 10220 14122 10226 14156
rect 10260 14122 10266 14156
rect 10220 14084 10266 14122
rect 10220 14050 10226 14084
rect 10260 14050 10266 14084
rect 10220 14012 10266 14050
rect 10220 13978 10226 14012
rect 10260 13978 10266 14012
rect 10220 13940 10266 13978
rect 10220 13906 10226 13940
rect 10260 13906 10266 13940
rect 10220 13868 10266 13906
rect 10220 13834 10226 13868
rect 10260 13834 10266 13868
rect 10220 13796 10266 13834
rect 10220 13762 10226 13796
rect 10260 13762 10266 13796
rect 10220 13724 10266 13762
rect 10220 13690 10226 13724
rect 10260 13690 10266 13724
rect 10220 13652 10266 13690
rect 10220 13618 10226 13652
rect 10260 13618 10266 13652
rect 10220 13580 10266 13618
rect 10220 13546 10226 13580
rect 10260 13546 10266 13580
rect 10220 13508 10266 13546
rect 10220 13474 10226 13508
rect 10260 13474 10266 13508
rect 10220 13436 10266 13474
rect 10220 13402 10226 13436
rect 10260 13402 10266 13436
rect 10220 13364 10266 13402
rect 10220 13330 10226 13364
rect 10260 13330 10266 13364
rect 10220 13292 10266 13330
rect 10220 13258 10226 13292
rect 10260 13258 10266 13292
rect 10220 13220 10266 13258
rect 10220 13186 10226 13220
rect 10260 13186 10266 13220
rect 10220 13148 10266 13186
rect 10220 13114 10226 13148
rect 10260 13114 10266 13148
rect 10220 13076 10266 13114
rect 10220 13042 10226 13076
rect 10260 13042 10266 13076
rect 10220 13004 10266 13042
rect 10220 12970 10226 13004
rect 10260 12970 10266 13004
rect 10220 12932 10266 12970
rect 10220 12898 10226 12932
rect 10260 12898 10266 12932
rect 10220 12860 10266 12898
rect 10220 12826 10226 12860
rect 10260 12826 10266 12860
rect 10220 12788 10266 12826
rect 10220 12754 10226 12788
rect 10260 12754 10266 12788
rect 10220 12716 10266 12754
rect 10220 12682 10226 12716
rect 10260 12682 10266 12716
rect 10220 12644 10266 12682
rect 10220 12610 10226 12644
rect 10260 12610 10266 12644
rect 10220 12572 10266 12610
rect 10220 12538 10226 12572
rect 10260 12538 10266 12572
rect 10220 12500 10266 12538
rect 10220 12466 10226 12500
rect 10260 12466 10266 12500
rect 10220 12428 10266 12466
rect 10220 12394 10226 12428
rect 10260 12394 10266 12428
rect 10220 12356 10266 12394
rect 10220 12322 10226 12356
rect 10260 12322 10266 12356
rect 10220 12284 10266 12322
rect 10220 12250 10226 12284
rect 10260 12250 10266 12284
rect 10220 12212 10266 12250
rect 10220 12178 10226 12212
rect 10260 12178 10266 12212
rect 10220 12140 10266 12178
rect 10220 12106 10226 12140
rect 10260 12106 10266 12140
rect 10220 12068 10266 12106
rect 10220 12034 10226 12068
rect 10260 12034 10266 12068
rect 10220 11996 10266 12034
rect 10220 11962 10226 11996
rect 10260 11962 10266 11996
rect 10220 11924 10266 11962
rect 10220 11890 10226 11924
rect 10260 11890 10266 11924
rect 10220 11852 10266 11890
rect 10220 11818 10226 11852
rect 10260 11818 10266 11852
rect 10220 11780 10266 11818
rect 10220 11746 10226 11780
rect 10260 11746 10266 11780
rect 10220 11708 10266 11746
rect 10220 11674 10226 11708
rect 10260 11674 10266 11708
rect 10220 11636 10266 11674
rect 10220 11602 10226 11636
rect 10260 11602 10266 11636
rect 10220 11564 10266 11602
rect 10220 11530 10226 11564
rect 10260 11530 10266 11564
rect 10220 11492 10266 11530
rect 10220 11458 10226 11492
rect 10260 11458 10266 11492
rect 10220 11420 10266 11458
rect 10220 11386 10226 11420
rect 10260 11386 10266 11420
rect 10220 11348 10266 11386
rect 10220 11314 10226 11348
rect 10260 11314 10266 11348
rect 10220 11276 10266 11314
rect 10220 11242 10226 11276
rect 10260 11242 10266 11276
rect 10220 11204 10266 11242
rect 10220 11170 10226 11204
rect 10260 11170 10266 11204
rect 10220 11132 10266 11170
rect 10220 11098 10226 11132
rect 10260 11098 10266 11132
rect 10220 11060 10266 11098
rect 10220 11026 10226 11060
rect 10260 11026 10266 11060
rect 10220 10988 10266 11026
rect 10220 10954 10226 10988
rect 10260 10954 10266 10988
rect 10220 10916 10266 10954
rect 10220 10882 10226 10916
rect 10260 10882 10266 10916
rect 10220 10844 10266 10882
rect 10220 10810 10226 10844
rect 10260 10810 10266 10844
rect 10220 10772 10266 10810
rect 10220 10738 10226 10772
rect 10260 10738 10266 10772
rect 10220 10700 10266 10738
rect 10220 10666 10226 10700
rect 10260 10666 10266 10700
rect 10220 10628 10266 10666
rect 10220 10594 10226 10628
rect 10260 10594 10266 10628
rect 10220 10556 10266 10594
rect 10220 10522 10226 10556
rect 10260 10522 10266 10556
rect 10220 10484 10266 10522
rect 10220 10450 10226 10484
rect 10260 10450 10266 10484
rect 10220 10412 10266 10450
rect 10220 10378 10226 10412
rect 10260 10378 10266 10412
rect 10220 10340 10266 10378
rect 10220 10306 10226 10340
rect 10260 10306 10266 10340
rect 10220 10268 10266 10306
rect 10220 10234 10226 10268
rect 10260 10234 10266 10268
rect 10220 10196 10266 10234
rect 10220 10162 10226 10196
rect 10260 10162 10266 10196
rect 10220 10124 10266 10162
rect 10220 10090 10226 10124
rect 10260 10090 10266 10124
rect 10220 10052 10266 10090
rect 10220 10018 10226 10052
rect 10260 10018 10266 10052
rect 10220 9980 10266 10018
rect 10220 9946 10226 9980
rect 10260 9946 10266 9980
rect 10220 9908 10266 9946
rect 10220 9874 10226 9908
rect 10260 9874 10266 9908
rect 10220 9836 10266 9874
rect 10220 9802 10226 9836
rect 10260 9802 10266 9836
rect 10220 9764 10266 9802
rect 10220 9730 10226 9764
rect 10260 9730 10266 9764
rect 10220 9692 10266 9730
rect 10220 9658 10226 9692
rect 10260 9658 10266 9692
rect 10220 9620 10266 9658
rect 10220 9586 10226 9620
rect 10260 9586 10266 9620
rect 10220 9548 10266 9586
rect 10220 9514 10226 9548
rect 10260 9514 10266 9548
rect 10220 9476 10266 9514
rect 10220 9442 10226 9476
rect 10260 9442 10266 9476
rect 10220 9404 10266 9442
rect 10220 9370 10226 9404
rect 10260 9370 10266 9404
rect 10220 9332 10266 9370
rect 10220 9298 10226 9332
rect 10260 9298 10266 9332
rect 10220 9260 10266 9298
rect 10220 9226 10226 9260
rect 10260 9226 10266 9260
rect 10220 9188 10266 9226
rect 10220 9154 10226 9188
rect 10260 9154 10266 9188
rect 10220 9116 10266 9154
rect 10220 9082 10226 9116
rect 10260 9082 10266 9116
rect 10220 9044 10266 9082
rect 10220 9010 10226 9044
rect 10260 9010 10266 9044
rect 10220 8972 10266 9010
rect 10220 8938 10226 8972
rect 10260 8938 10266 8972
rect 10220 8900 10266 8938
rect 10220 8866 10226 8900
rect 10260 8866 10266 8900
rect 10220 8828 10266 8866
rect 10220 8794 10226 8828
rect 10260 8794 10266 8828
rect 10220 8756 10266 8794
rect 10220 8722 10226 8756
rect 10260 8722 10266 8756
rect 10220 8684 10266 8722
rect 10220 8650 10226 8684
rect 10260 8650 10266 8684
rect 10220 8612 10266 8650
rect 10220 8578 10226 8612
rect 10260 8578 10266 8612
rect 10220 8540 10266 8578
rect 10220 8506 10226 8540
rect 10260 8506 10266 8540
rect 10220 8468 10266 8506
rect 10220 8434 10226 8468
rect 10260 8434 10266 8468
rect 10220 8396 10266 8434
rect 10220 8362 10226 8396
rect 10260 8362 10266 8396
rect 10220 8324 10266 8362
rect 10220 8290 10226 8324
rect 10260 8290 10266 8324
rect 10220 8252 10266 8290
rect 10220 8218 10226 8252
rect 10260 8218 10266 8252
rect 10220 8180 10266 8218
rect 10220 8146 10226 8180
rect 10260 8146 10266 8180
rect 10220 8108 10266 8146
rect 10220 8074 10226 8108
rect 10260 8074 10266 8108
rect 10220 8036 10266 8074
rect 10220 8002 10226 8036
rect 10260 8002 10266 8036
rect 10220 7964 10266 8002
rect 10220 7930 10226 7964
rect 10260 7930 10266 7964
rect 10220 7892 10266 7930
rect 10220 7858 10226 7892
rect 10260 7858 10266 7892
rect 10220 7820 10266 7858
rect 10220 7786 10226 7820
rect 10260 7786 10266 7820
rect 10220 7748 10266 7786
rect 10220 7714 10226 7748
rect 10260 7714 10266 7748
rect 10220 7676 10266 7714
rect 10220 7642 10226 7676
rect 10260 7642 10266 7676
rect 10220 7604 10266 7642
rect 10220 7570 10226 7604
rect 10260 7570 10266 7604
rect 10220 7532 10266 7570
rect 10220 7498 10226 7532
rect 10260 7498 10266 7532
rect 10220 7460 10266 7498
rect 10220 7426 10226 7460
rect 10260 7426 10266 7460
rect 10220 7388 10266 7426
rect 10220 7354 10226 7388
rect 10260 7354 10266 7388
rect 10220 7316 10266 7354
rect 10220 7282 10226 7316
rect 10260 7282 10266 7316
rect 10220 7244 10266 7282
rect 10220 7210 10226 7244
rect 10260 7210 10266 7244
rect 10220 7172 10266 7210
rect 10220 7138 10226 7172
rect 10260 7138 10266 7172
rect 10220 7100 10266 7138
rect 10220 7066 10226 7100
rect 10260 7066 10266 7100
rect 10220 7028 10266 7066
rect 10220 6994 10226 7028
rect 10260 6994 10266 7028
rect 10220 6956 10266 6994
rect 10220 6922 10226 6956
rect 10260 6922 10266 6956
rect 10220 6884 10266 6922
rect 10220 6850 10226 6884
rect 10260 6850 10266 6884
rect 10220 6812 10266 6850
rect 10220 6778 10226 6812
rect 10260 6778 10266 6812
rect 10220 6740 10266 6778
rect 10220 6706 10226 6740
rect 10260 6706 10266 6740
rect 10220 6668 10266 6706
rect 10220 6634 10226 6668
rect 10260 6634 10266 6668
rect 10220 6596 10266 6634
rect 10220 6562 10226 6596
rect 10260 6562 10266 6596
rect 10220 6524 10266 6562
rect 10220 6490 10226 6524
rect 10260 6490 10266 6524
rect 10220 6452 10266 6490
rect 10220 6418 10226 6452
rect 10260 6418 10266 6452
rect 10220 6380 10266 6418
rect 10220 6346 10226 6380
rect 10260 6346 10266 6380
rect 10220 6308 10266 6346
rect 10220 6274 10226 6308
rect 10260 6274 10266 6308
rect 10220 6236 10266 6274
rect 10220 6202 10226 6236
rect 10260 6202 10266 6236
rect 10220 6164 10266 6202
rect 10220 6130 10226 6164
rect 10260 6130 10266 6164
rect 10220 6092 10266 6130
rect 10220 6058 10226 6092
rect 10260 6058 10266 6092
rect 10220 6020 10266 6058
rect 10220 5986 10226 6020
rect 10260 5986 10266 6020
rect 10220 5948 10266 5986
rect 10220 5914 10226 5948
rect 10260 5914 10266 5948
rect 10220 5876 10266 5914
rect 10220 5842 10226 5876
rect 10260 5842 10266 5876
rect 10220 5804 10266 5842
rect 10220 5770 10226 5804
rect 10260 5770 10266 5804
rect 10220 5732 10266 5770
rect 10220 5698 10226 5732
rect 10260 5698 10266 5732
rect 10220 5660 10266 5698
rect 10220 5626 10226 5660
rect 10260 5626 10266 5660
rect 10220 5588 10266 5626
rect 10220 5554 10226 5588
rect 10260 5554 10266 5588
rect 10220 5516 10266 5554
rect 10220 5482 10226 5516
rect 10260 5482 10266 5516
rect 10220 5444 10266 5482
rect 10220 5410 10226 5444
rect 10260 5410 10266 5444
rect 10220 5372 10266 5410
rect 10220 5338 10226 5372
rect 10260 5338 10266 5372
rect 10220 5300 10266 5338
rect 10220 5266 10226 5300
rect 10260 5266 10266 5300
rect 10220 5228 10266 5266
rect 10220 5194 10226 5228
rect 10260 5194 10266 5228
rect 10220 5156 10266 5194
rect 10220 5122 10226 5156
rect 10260 5122 10266 5156
rect 10220 5084 10266 5122
rect 10220 5050 10226 5084
rect 10260 5050 10266 5084
rect 10220 5012 10266 5050
rect 10220 4978 10226 5012
rect 10260 4978 10266 5012
rect 10220 4940 10266 4978
rect 10220 4906 10226 4940
rect 10260 4906 10266 4940
rect 10220 4868 10266 4906
rect 10220 4834 10226 4868
rect 10260 4834 10266 4868
rect 10220 4796 10266 4834
rect 10220 4762 10226 4796
rect 10260 4762 10266 4796
rect 10220 4724 10266 4762
rect 10220 4690 10226 4724
rect 10260 4690 10266 4724
rect 10220 4652 10266 4690
rect 10220 4618 10226 4652
rect 10260 4618 10266 4652
rect 10220 4580 10266 4618
rect 10220 4546 10226 4580
rect 10260 4546 10266 4580
rect 10220 4508 10266 4546
rect 10220 4474 10226 4508
rect 10260 4474 10266 4508
rect 10220 4436 10266 4474
rect 10220 4402 10226 4436
rect 10260 4402 10266 4436
rect 10220 4364 10266 4402
rect 10220 4330 10226 4364
rect 10260 4330 10266 4364
rect 10220 4292 10266 4330
rect 10220 4258 10226 4292
rect 10260 4258 10266 4292
rect 10220 4220 10266 4258
rect 10220 4186 10226 4220
rect 10260 4186 10266 4220
rect 10220 4148 10266 4186
rect 10220 4114 10226 4148
rect 10260 4114 10266 4148
rect 10220 4076 10266 4114
rect 10220 4042 10226 4076
rect 10260 4042 10266 4076
rect 10220 4004 10266 4042
rect 10220 3970 10226 4004
rect 10260 3970 10266 4004
rect 10220 3932 10266 3970
rect 10220 3898 10226 3932
rect 10260 3898 10266 3932
rect 10220 3860 10266 3898
rect 10220 3826 10226 3860
rect 10260 3826 10266 3860
rect 10220 3788 10266 3826
rect 10220 3754 10226 3788
rect 10260 3754 10266 3788
rect 10220 3716 10266 3754
rect 10220 3682 10226 3716
rect 10260 3682 10266 3716
rect 10220 3644 10266 3682
rect 10220 3610 10226 3644
rect 10260 3610 10266 3644
rect 10220 3572 10266 3610
rect 10220 3538 10226 3572
rect 10260 3538 10266 3572
rect 10220 3500 10266 3538
rect 9082 3428 9128 3466
rect 9082 3394 9088 3428
rect 9122 3394 9128 3428
rect 9082 3356 9128 3394
rect 9205 3493 9257 3499
rect 9205 3429 9257 3441
rect 9205 3369 9257 3377
rect 9323 3487 9493 3499
rect 9323 3453 9332 3487
rect 9366 3453 9450 3487
rect 9484 3453 9493 3487
rect 9323 3415 9493 3453
rect 9323 3381 9332 3415
rect 9366 3381 9450 3415
rect 9484 3381 9493 3415
rect 9323 3369 9493 3381
rect 9559 3487 9729 3499
rect 9559 3453 9568 3487
rect 9602 3453 9686 3487
rect 9720 3453 9729 3487
rect 9559 3415 9729 3453
rect 9559 3381 9568 3415
rect 9602 3381 9686 3415
rect 9720 3381 9729 3415
rect 9559 3369 9729 3381
rect 9795 3487 9965 3499
rect 9795 3453 9804 3487
rect 9838 3453 9922 3487
rect 9956 3453 9965 3487
rect 9795 3415 9965 3453
rect 9795 3381 9804 3415
rect 9838 3381 9922 3415
rect 9956 3381 9965 3415
rect 9795 3369 9965 3381
rect 10031 3493 10083 3499
rect 10031 3429 10083 3441
rect 10031 3369 10083 3377
rect 10220 3466 10226 3500
rect 10260 3466 10266 3500
rect 11418 38650 11424 38684
rect 11458 38650 11464 38684
tri 11464 38682 11466 38684 nw
tri 13204 38682 13206 38684 ne
rect 11418 38611 11464 38650
rect 13206 38650 13212 38684
rect 13246 38650 13252 38684
tri 13252 38682 13254 38684 nw
tri 14932 38682 14934 38684 ne
rect 11418 38577 11424 38611
rect 11458 38577 11464 38611
rect 11418 38538 11464 38577
rect 12880 38572 12886 38624
rect 12938 38615 13000 38624
rect 12938 38581 12964 38615
rect 12998 38581 13000 38615
rect 13052 38612 13078 38624
rect 12938 38572 13000 38581
rect 13072 38578 13078 38612
rect 13052 38572 13078 38578
tri 12998 38540 13030 38572 ne
rect 13030 38540 13078 38572
tri 13030 38538 13032 38540 ne
rect 11418 38504 11424 38538
rect 11458 38504 11464 38538
rect 11418 38465 11464 38504
rect 13032 38517 13078 38540
rect 13032 38483 13038 38517
rect 13072 38483 13078 38517
rect 13032 38471 13078 38483
rect 13206 38611 13252 38650
rect 14934 38650 14940 38684
rect 14974 38650 14980 38684
rect 13206 38577 13212 38611
rect 13246 38577 13252 38611
rect 13206 38538 13252 38577
rect 13206 38504 13212 38538
rect 13246 38504 13252 38538
rect 11418 38431 11424 38465
rect 11458 38431 11464 38465
rect 11418 38392 11464 38431
rect 11418 38358 11424 38392
rect 11458 38358 11464 38392
rect 11418 38319 11464 38358
rect 11418 38285 11424 38319
rect 11458 38285 11464 38319
rect 11418 38246 11464 38285
rect 11418 38212 11424 38246
rect 11458 38212 11464 38246
rect 11418 38173 11464 38212
rect 11418 38139 11424 38173
rect 11458 38139 11464 38173
rect 11418 38100 11464 38139
rect 11418 38066 11424 38100
rect 11458 38066 11464 38100
rect 11418 38027 11464 38066
rect 11418 37993 11424 38027
rect 11458 37993 11464 38027
rect 11418 37954 11464 37993
rect 11418 37920 11424 37954
rect 11458 37920 11464 37954
rect 11418 37881 11464 37920
rect 11418 37847 11424 37881
rect 11458 37847 11464 37881
rect 11418 37808 11464 37847
rect 11418 37774 11424 37808
rect 11458 37774 11464 37808
rect 11418 37735 11464 37774
rect 11418 37701 11424 37735
rect 11458 37701 11464 37735
rect 11418 37662 11464 37701
rect 11418 37628 11424 37662
rect 11458 37628 11464 37662
rect 11418 37589 11464 37628
rect 11418 37555 11424 37589
rect 11458 37555 11464 37589
rect 11418 37516 11464 37555
rect 11418 37482 11424 37516
rect 11458 37482 11464 37516
rect 11418 37443 11464 37482
rect 11418 37409 11424 37443
rect 11458 37409 11464 37443
rect 11418 37370 11464 37409
rect 11418 37336 11424 37370
rect 11458 37336 11464 37370
rect 11418 37297 11464 37336
rect 11418 37263 11424 37297
rect 11458 37263 11464 37297
rect 11418 37224 11464 37263
rect 11418 37190 11424 37224
rect 11458 37190 11464 37224
rect 11418 37151 11464 37190
rect 11418 37117 11424 37151
rect 11458 37117 11464 37151
rect 11418 37078 11464 37117
rect 11418 37044 11424 37078
rect 11458 37044 11464 37078
rect 11418 37005 11464 37044
rect 11418 36971 11424 37005
rect 11458 36971 11464 37005
rect 11418 36932 11464 36971
rect 11418 36898 11424 36932
rect 11458 36898 11464 36932
rect 11418 36859 11464 36898
rect 11418 36825 11424 36859
rect 11458 36825 11464 36859
rect 11418 36786 11464 36825
rect 11418 36752 11424 36786
rect 11458 36752 11464 36786
rect 11418 36713 11464 36752
rect 11418 36679 11424 36713
rect 11458 36679 11464 36713
rect 11418 36640 11464 36679
rect 11418 36606 11424 36640
rect 11458 36606 11464 36640
rect 11418 36567 11464 36606
rect 11418 36533 11424 36567
rect 11458 36533 11464 36567
rect 11418 36494 11464 36533
rect 11418 36460 11424 36494
rect 11458 36460 11464 36494
rect 11418 36421 11464 36460
rect 11418 36387 11424 36421
rect 11458 36387 11464 36421
rect 11418 36348 11464 36387
rect 11418 36314 11424 36348
rect 11458 36314 11464 36348
rect 11418 36275 11464 36314
rect 11418 36241 11424 36275
rect 11458 36241 11464 36275
rect 11418 36202 11464 36241
rect 11418 36168 11424 36202
rect 11458 36168 11464 36202
rect 11418 36129 11464 36168
rect 11418 36095 11424 36129
rect 11458 36095 11464 36129
rect 11418 36056 11464 36095
rect 11418 36022 11424 36056
rect 11458 36022 11464 36056
rect 11418 35983 11464 36022
rect 11418 35949 11424 35983
rect 11458 35949 11464 35983
rect 11418 35910 11464 35949
rect 11418 35876 11424 35910
rect 11458 35876 11464 35910
rect 11418 35837 11464 35876
rect 11418 35803 11424 35837
rect 11458 35803 11464 35837
rect 11418 35764 11464 35803
rect 11418 35730 11424 35764
rect 11458 35730 11464 35764
rect 11418 35691 11464 35730
rect 11418 35657 11424 35691
rect 11458 35657 11464 35691
rect 11418 35618 11464 35657
rect 11418 35584 11424 35618
rect 11458 35584 11464 35618
rect 11418 35545 11464 35584
rect 11418 35511 11424 35545
rect 11458 35511 11464 35545
rect 11418 35472 11464 35511
rect 11418 35438 11424 35472
rect 11458 35438 11464 35472
rect 11418 35399 11464 35438
rect 11418 35365 11424 35399
rect 11458 35365 11464 35399
rect 11418 35326 11464 35365
rect 11418 35292 11424 35326
rect 11458 35292 11464 35326
rect 11418 35253 11464 35292
rect 11418 35219 11424 35253
rect 11458 35219 11464 35253
rect 11418 35180 11464 35219
rect 11418 35146 11424 35180
rect 11458 35146 11464 35180
rect 11418 35108 11464 35146
rect 11418 35074 11424 35108
rect 11458 35074 11464 35108
rect 11418 35036 11464 35074
rect 11418 35002 11424 35036
rect 11458 35002 11464 35036
rect 11418 34964 11464 35002
rect 11418 34930 11424 34964
rect 11458 34930 11464 34964
rect 11418 34892 11464 34930
rect 11418 34858 11424 34892
rect 11458 34858 11464 34892
rect 11418 34820 11464 34858
rect 11418 34786 11424 34820
rect 11458 34786 11464 34820
rect 11418 34748 11464 34786
rect 11418 34714 11424 34748
rect 11458 34714 11464 34748
rect 11418 34676 11464 34714
rect 11418 34642 11424 34676
rect 11458 34642 11464 34676
rect 11418 34604 11464 34642
rect 11418 34570 11424 34604
rect 11458 34570 11464 34604
rect 11418 34532 11464 34570
rect 11418 34498 11424 34532
rect 11458 34498 11464 34532
rect 11418 34460 11464 34498
rect 11418 34426 11424 34460
rect 11458 34426 11464 34460
rect 11418 34388 11464 34426
rect 11418 34354 11424 34388
rect 11458 34354 11464 34388
rect 11418 34316 11464 34354
rect 11418 34282 11424 34316
rect 11458 34282 11464 34316
rect 11418 34244 11464 34282
rect 11418 34210 11424 34244
rect 11458 34210 11464 34244
rect 11418 34172 11464 34210
rect 11418 34138 11424 34172
rect 11458 34138 11464 34172
rect 11418 34100 11464 34138
rect 11418 34066 11424 34100
rect 11458 34066 11464 34100
rect 11418 34028 11464 34066
rect 11418 33994 11424 34028
rect 11458 33994 11464 34028
rect 11418 33956 11464 33994
rect 11418 33922 11424 33956
rect 11458 33922 11464 33956
rect 11418 33884 11464 33922
rect 11418 33850 11424 33884
rect 11458 33850 11464 33884
rect 11418 33812 11464 33850
rect 11418 33778 11424 33812
rect 11458 33778 11464 33812
rect 11418 33740 11464 33778
rect 11418 33706 11424 33740
rect 11458 33706 11464 33740
rect 11418 33668 11464 33706
rect 11418 33634 11424 33668
rect 11458 33634 11464 33668
rect 11418 33596 11464 33634
rect 11418 33562 11424 33596
rect 11458 33562 11464 33596
rect 11418 33524 11464 33562
rect 11418 33490 11424 33524
rect 11458 33490 11464 33524
rect 11418 33452 11464 33490
rect 11418 33418 11424 33452
rect 11458 33418 11464 33452
rect 11418 33380 11464 33418
rect 11418 33346 11424 33380
rect 11458 33346 11464 33380
rect 11418 33308 11464 33346
rect 11418 33274 11424 33308
rect 11458 33274 11464 33308
rect 11418 33236 11464 33274
rect 11418 33202 11424 33236
rect 11458 33202 11464 33236
rect 11418 33164 11464 33202
rect 11418 33130 11424 33164
rect 11458 33130 11464 33164
rect 11418 33092 11464 33130
rect 11418 33058 11424 33092
rect 11458 33058 11464 33092
rect 11418 33020 11464 33058
rect 11418 32986 11424 33020
rect 11458 32986 11464 33020
rect 11418 32948 11464 32986
rect 11418 32914 11424 32948
rect 11458 32914 11464 32948
rect 11418 32876 11464 32914
rect 11418 32842 11424 32876
rect 11458 32842 11464 32876
rect 11418 32804 11464 32842
rect 11418 32770 11424 32804
rect 11458 32770 11464 32804
rect 11418 32732 11464 32770
rect 11418 32698 11424 32732
rect 11458 32698 11464 32732
rect 11418 32660 11464 32698
rect 11418 32626 11424 32660
rect 11458 32626 11464 32660
rect 11418 32588 11464 32626
rect 11418 32554 11424 32588
rect 11458 32554 11464 32588
rect 11418 32516 11464 32554
rect 11418 32482 11424 32516
rect 11458 32482 11464 32516
rect 11418 32444 11464 32482
rect 11418 32410 11424 32444
rect 11458 32410 11464 32444
rect 11418 32372 11464 32410
rect 11418 32338 11424 32372
rect 11458 32338 11464 32372
rect 11418 32300 11464 32338
rect 11418 32266 11424 32300
rect 11458 32266 11464 32300
rect 11418 32228 11464 32266
rect 11418 32194 11424 32228
rect 11458 32194 11464 32228
rect 11418 32156 11464 32194
rect 11418 32122 11424 32156
rect 11458 32122 11464 32156
rect 11418 32084 11464 32122
rect 11418 32050 11424 32084
rect 11458 32050 11464 32084
rect 11418 32012 11464 32050
rect 11418 31978 11424 32012
rect 11458 31978 11464 32012
rect 11418 31940 11464 31978
rect 11418 31906 11424 31940
rect 11458 31906 11464 31940
rect 11418 31868 11464 31906
rect 11418 31834 11424 31868
rect 11458 31834 11464 31868
rect 11418 31796 11464 31834
rect 11418 31762 11424 31796
rect 11458 31762 11464 31796
rect 11418 31724 11464 31762
rect 11418 31690 11424 31724
rect 11458 31690 11464 31724
rect 11418 31652 11464 31690
rect 11418 31618 11424 31652
rect 11458 31618 11464 31652
rect 11418 31580 11464 31618
rect 11418 31546 11424 31580
rect 11458 31546 11464 31580
rect 11418 31508 11464 31546
rect 11418 31474 11424 31508
rect 11458 31474 11464 31508
rect 11418 31436 11464 31474
rect 11418 31402 11424 31436
rect 11458 31402 11464 31436
rect 11418 31364 11464 31402
rect 11418 31330 11424 31364
rect 11458 31330 11464 31364
rect 11418 31292 11464 31330
rect 11418 31258 11424 31292
rect 11458 31258 11464 31292
rect 11418 31220 11464 31258
rect 11418 31186 11424 31220
rect 11458 31186 11464 31220
rect 11418 31148 11464 31186
rect 11418 31114 11424 31148
rect 11458 31114 11464 31148
rect 11418 31076 11464 31114
rect 11418 31042 11424 31076
rect 11458 31042 11464 31076
rect 11418 31004 11464 31042
rect 11418 30970 11424 31004
rect 11458 30970 11464 31004
rect 11418 30932 11464 30970
rect 11418 30898 11424 30932
rect 11458 30898 11464 30932
rect 11418 30860 11464 30898
rect 11418 30826 11424 30860
rect 11458 30826 11464 30860
rect 11418 30788 11464 30826
rect 11418 30754 11424 30788
rect 11458 30754 11464 30788
rect 11418 30716 11464 30754
rect 11418 30682 11424 30716
rect 11458 30682 11464 30716
rect 11418 30644 11464 30682
rect 11418 30610 11424 30644
rect 11458 30610 11464 30644
rect 11418 30572 11464 30610
rect 11418 30538 11424 30572
rect 11458 30538 11464 30572
rect 11418 30500 11464 30538
rect 11418 30466 11424 30500
rect 11458 30466 11464 30500
rect 11418 30428 11464 30466
rect 11418 30394 11424 30428
rect 11458 30394 11464 30428
rect 11418 30356 11464 30394
rect 11418 30322 11424 30356
rect 11458 30322 11464 30356
rect 11418 30284 11464 30322
rect 11418 30250 11424 30284
rect 11458 30250 11464 30284
rect 11418 30212 11464 30250
rect 11418 30178 11424 30212
rect 11458 30178 11464 30212
rect 11418 30140 11464 30178
rect 11418 30106 11424 30140
rect 11458 30106 11464 30140
rect 11418 30068 11464 30106
rect 11418 30034 11424 30068
rect 11458 30034 11464 30068
rect 11418 29996 11464 30034
rect 11418 29962 11424 29996
rect 11458 29962 11464 29996
rect 11418 29924 11464 29962
rect 11418 29890 11424 29924
rect 11458 29890 11464 29924
rect 11418 29852 11464 29890
rect 11418 29818 11424 29852
rect 11458 29818 11464 29852
rect 11418 29780 11464 29818
rect 11418 29746 11424 29780
rect 11458 29746 11464 29780
rect 11418 29708 11464 29746
rect 11418 29674 11424 29708
rect 11458 29674 11464 29708
rect 11418 29636 11464 29674
rect 11418 29602 11424 29636
rect 11458 29602 11464 29636
rect 11418 29564 11464 29602
rect 11418 29530 11424 29564
rect 11458 29530 11464 29564
rect 11418 29492 11464 29530
rect 11418 29458 11424 29492
rect 11458 29458 11464 29492
rect 11418 29420 11464 29458
rect 11418 29386 11424 29420
rect 11458 29386 11464 29420
rect 11418 29348 11464 29386
rect 11418 29314 11424 29348
rect 11458 29314 11464 29348
rect 11418 29276 11464 29314
rect 11418 29242 11424 29276
rect 11458 29242 11464 29276
rect 11418 29204 11464 29242
rect 11418 29170 11424 29204
rect 11458 29170 11464 29204
rect 11418 29132 11464 29170
rect 11418 29098 11424 29132
rect 11458 29098 11464 29132
rect 11418 29060 11464 29098
rect 11418 29026 11424 29060
rect 11458 29026 11464 29060
rect 11418 28988 11464 29026
rect 11418 28954 11424 28988
rect 11458 28954 11464 28988
rect 11418 28916 11464 28954
rect 11418 28882 11424 28916
rect 11458 28882 11464 28916
rect 11418 28844 11464 28882
rect 11418 28810 11424 28844
rect 11458 28810 11464 28844
rect 11418 28772 11464 28810
rect 11418 28738 11424 28772
rect 11458 28738 11464 28772
rect 11418 28700 11464 28738
rect 11418 28666 11424 28700
rect 11458 28666 11464 28700
rect 11418 28628 11464 28666
rect 11418 28594 11424 28628
rect 11458 28594 11464 28628
rect 11418 28556 11464 28594
rect 11418 28522 11424 28556
rect 11458 28522 11464 28556
rect 11418 28484 11464 28522
rect 11418 28450 11424 28484
rect 11458 28450 11464 28484
rect 11418 28412 11464 28450
rect 11418 28378 11424 28412
rect 11458 28378 11464 28412
rect 11418 28340 11464 28378
rect 11418 28306 11424 28340
rect 11458 28306 11464 28340
rect 11418 28268 11464 28306
rect 11418 28234 11424 28268
rect 11458 28234 11464 28268
rect 11418 28196 11464 28234
rect 11418 28162 11424 28196
rect 11458 28162 11464 28196
rect 11418 28124 11464 28162
rect 11418 28090 11424 28124
rect 11458 28090 11464 28124
rect 11418 28052 11464 28090
rect 11418 28018 11424 28052
rect 11458 28018 11464 28052
rect 11418 27980 11464 28018
rect 11418 27946 11424 27980
rect 11458 27946 11464 27980
rect 11418 27908 11464 27946
rect 11418 27874 11424 27908
rect 11458 27874 11464 27908
rect 11418 27836 11464 27874
rect 11418 27802 11424 27836
rect 11458 27802 11464 27836
rect 11418 27764 11464 27802
rect 11418 27730 11424 27764
rect 11458 27730 11464 27764
rect 11418 27692 11464 27730
rect 11418 27658 11424 27692
rect 11458 27658 11464 27692
rect 11418 27620 11464 27658
rect 11418 27586 11424 27620
rect 11458 27586 11464 27620
rect 11418 27548 11464 27586
rect 11418 27514 11424 27548
rect 11458 27514 11464 27548
rect 11418 27476 11464 27514
rect 11418 27442 11424 27476
rect 11458 27442 11464 27476
rect 11418 27404 11464 27442
rect 11418 27370 11424 27404
rect 11458 27370 11464 27404
rect 11418 27332 11464 27370
rect 11418 27298 11424 27332
rect 11458 27298 11464 27332
rect 11418 27260 11464 27298
rect 11418 27226 11424 27260
rect 11458 27226 11464 27260
rect 11418 27188 11464 27226
rect 11418 27154 11424 27188
rect 11458 27154 11464 27188
rect 11418 27116 11464 27154
rect 11418 27082 11424 27116
rect 11458 27082 11464 27116
rect 11418 27044 11464 27082
rect 11418 27010 11424 27044
rect 11458 27010 11464 27044
rect 11418 26972 11464 27010
rect 11418 26938 11424 26972
rect 11458 26938 11464 26972
rect 11418 26900 11464 26938
rect 11418 26866 11424 26900
rect 11458 26866 11464 26900
rect 11418 26828 11464 26866
rect 11418 26794 11424 26828
rect 11458 26794 11464 26828
rect 11418 26756 11464 26794
rect 11418 26722 11424 26756
rect 11458 26722 11464 26756
rect 11418 26684 11464 26722
rect 11418 26650 11424 26684
rect 11458 26650 11464 26684
rect 11418 26612 11464 26650
rect 11418 26578 11424 26612
rect 11458 26578 11464 26612
rect 11418 26540 11464 26578
rect 11418 26506 11424 26540
rect 11458 26506 11464 26540
rect 11418 26468 11464 26506
rect 11418 26434 11424 26468
rect 11458 26434 11464 26468
rect 11418 26396 11464 26434
rect 11418 26362 11424 26396
rect 11458 26362 11464 26396
rect 11418 26324 11464 26362
rect 11418 26290 11424 26324
rect 11458 26290 11464 26324
rect 11418 26252 11464 26290
rect 11418 26218 11424 26252
rect 11458 26218 11464 26252
rect 11418 26180 11464 26218
rect 11418 26146 11424 26180
rect 11458 26146 11464 26180
rect 11418 26108 11464 26146
rect 11418 26074 11424 26108
rect 11458 26074 11464 26108
rect 11418 26036 11464 26074
rect 11418 26002 11424 26036
rect 11458 26002 11464 26036
rect 11418 25964 11464 26002
rect 11418 25930 11424 25964
rect 11458 25930 11464 25964
rect 11418 25892 11464 25930
rect 11418 25858 11424 25892
rect 11458 25858 11464 25892
rect 11418 25820 11464 25858
rect 11418 25786 11424 25820
rect 11458 25786 11464 25820
rect 11418 25748 11464 25786
rect 11418 25714 11424 25748
rect 11458 25714 11464 25748
rect 11418 25676 11464 25714
rect 11418 25642 11424 25676
rect 11458 25642 11464 25676
rect 11418 25604 11464 25642
rect 11418 25570 11424 25604
rect 11458 25570 11464 25604
rect 11418 25532 11464 25570
rect 11418 25498 11424 25532
rect 11458 25498 11464 25532
rect 11418 25460 11464 25498
rect 11418 25426 11424 25460
rect 11458 25426 11464 25460
rect 11418 25388 11464 25426
rect 11418 25354 11424 25388
rect 11458 25354 11464 25388
rect 11418 25316 11464 25354
rect 11418 25282 11424 25316
rect 11458 25282 11464 25316
rect 11418 25244 11464 25282
rect 11418 25210 11424 25244
rect 11458 25210 11464 25244
rect 11418 25172 11464 25210
rect 11418 25138 11424 25172
rect 11458 25138 11464 25172
rect 11418 25100 11464 25138
rect 11418 25066 11424 25100
rect 11458 25066 11464 25100
rect 11418 25028 11464 25066
rect 11418 24994 11424 25028
rect 11458 24994 11464 25028
rect 11418 24956 11464 24994
rect 11418 24922 11424 24956
rect 11458 24922 11464 24956
rect 11418 24884 11464 24922
rect 11418 24850 11424 24884
rect 11458 24850 11464 24884
rect 11418 24812 11464 24850
rect 11418 24778 11424 24812
rect 11458 24778 11464 24812
rect 11418 24740 11464 24778
rect 11418 24706 11424 24740
rect 11458 24706 11464 24740
rect 11418 24668 11464 24706
rect 11418 24634 11424 24668
rect 11458 24634 11464 24668
rect 11418 24596 11464 24634
rect 11418 24562 11424 24596
rect 11458 24562 11464 24596
rect 11418 24524 11464 24562
rect 11418 24490 11424 24524
rect 11458 24490 11464 24524
rect 11418 24452 11464 24490
rect 11418 24418 11424 24452
rect 11458 24418 11464 24452
rect 11418 24380 11464 24418
rect 11418 24346 11424 24380
rect 11458 24346 11464 24380
rect 11418 24308 11464 24346
rect 11418 24274 11424 24308
rect 11458 24274 11464 24308
rect 11418 24236 11464 24274
rect 11418 24202 11424 24236
rect 11458 24202 11464 24236
rect 11418 24164 11464 24202
rect 11418 24130 11424 24164
rect 11458 24130 11464 24164
rect 11418 24092 11464 24130
rect 11418 24058 11424 24092
rect 11458 24058 11464 24092
rect 11418 24020 11464 24058
rect 11418 23986 11424 24020
rect 11458 23986 11464 24020
rect 11418 23948 11464 23986
rect 11418 23914 11424 23948
rect 11458 23914 11464 23948
rect 11418 23876 11464 23914
rect 11418 23842 11424 23876
rect 11458 23842 11464 23876
rect 11418 23804 11464 23842
rect 11418 23770 11424 23804
rect 11458 23770 11464 23804
rect 11418 23732 11464 23770
rect 11418 23698 11424 23732
rect 11458 23698 11464 23732
rect 11418 23660 11464 23698
rect 11418 23626 11424 23660
rect 11458 23626 11464 23660
rect 11418 23588 11464 23626
rect 11418 23554 11424 23588
rect 11458 23554 11464 23588
rect 11418 23516 11464 23554
rect 11418 23482 11424 23516
rect 11458 23482 11464 23516
rect 11418 23444 11464 23482
rect 11418 23410 11424 23444
rect 11458 23410 11464 23444
rect 11418 23372 11464 23410
rect 11418 23338 11424 23372
rect 11458 23338 11464 23372
rect 11418 23300 11464 23338
rect 11418 23266 11424 23300
rect 11458 23266 11464 23300
rect 11418 23228 11464 23266
rect 11418 23194 11424 23228
rect 11458 23194 11464 23228
rect 11418 23156 11464 23194
rect 11418 23122 11424 23156
rect 11458 23122 11464 23156
rect 11418 23084 11464 23122
rect 11418 23050 11424 23084
rect 11458 23050 11464 23084
rect 11418 23012 11464 23050
rect 11418 22978 11424 23012
rect 11458 22978 11464 23012
rect 11418 22940 11464 22978
rect 11418 22906 11424 22940
rect 11458 22906 11464 22940
rect 11418 22868 11464 22906
rect 11418 22834 11424 22868
rect 11458 22834 11464 22868
rect 11418 22796 11464 22834
rect 11418 22762 11424 22796
rect 11458 22762 11464 22796
rect 11418 22724 11464 22762
rect 11418 22690 11424 22724
rect 11458 22690 11464 22724
rect 11418 22652 11464 22690
rect 11418 22618 11424 22652
rect 11458 22618 11464 22652
rect 11418 22580 11464 22618
rect 11418 22546 11424 22580
rect 11458 22546 11464 22580
rect 11418 22508 11464 22546
rect 11418 22474 11424 22508
rect 11458 22474 11464 22508
rect 11418 22436 11464 22474
rect 11418 22402 11424 22436
rect 11458 22402 11464 22436
rect 11418 22364 11464 22402
rect 11418 22330 11424 22364
rect 11458 22330 11464 22364
rect 11418 22292 11464 22330
rect 11418 22258 11424 22292
rect 11458 22258 11464 22292
rect 11418 22220 11464 22258
rect 11418 22186 11424 22220
rect 11458 22186 11464 22220
rect 11418 22148 11464 22186
rect 11418 22114 11424 22148
rect 11458 22114 11464 22148
rect 11418 22076 11464 22114
rect 11418 22042 11424 22076
rect 11458 22042 11464 22076
rect 11418 22004 11464 22042
rect 11418 21970 11424 22004
rect 11458 21970 11464 22004
rect 11418 21932 11464 21970
rect 11418 21898 11424 21932
rect 11458 21898 11464 21932
rect 11418 21860 11464 21898
rect 11418 21826 11424 21860
rect 11458 21826 11464 21860
rect 11418 21788 11464 21826
rect 11418 21754 11424 21788
rect 11458 21754 11464 21788
rect 11418 21716 11464 21754
rect 11418 21682 11424 21716
rect 11458 21682 11464 21716
rect 11418 21644 11464 21682
rect 11418 21610 11424 21644
rect 11458 21610 11464 21644
rect 11418 21572 11464 21610
rect 11418 21538 11424 21572
rect 11458 21538 11464 21572
rect 11418 21500 11464 21538
rect 11418 21466 11424 21500
rect 11458 21466 11464 21500
rect 11418 21428 11464 21466
rect 11418 21394 11424 21428
rect 11458 21394 11464 21428
rect 11418 21356 11464 21394
rect 11418 21322 11424 21356
rect 11458 21322 11464 21356
rect 11418 21284 11464 21322
rect 11418 21250 11424 21284
rect 11458 21250 11464 21284
rect 11418 21212 11464 21250
rect 11418 21178 11424 21212
rect 11458 21178 11464 21212
rect 11418 21140 11464 21178
rect 11418 21106 11424 21140
rect 11458 21106 11464 21140
rect 11418 21068 11464 21106
rect 11418 21034 11424 21068
rect 11458 21034 11464 21068
rect 11418 20996 11464 21034
rect 11418 20962 11424 20996
rect 11458 20962 11464 20996
rect 11418 20924 11464 20962
rect 11418 20890 11424 20924
rect 11458 20890 11464 20924
rect 11418 20852 11464 20890
rect 11418 20818 11424 20852
rect 11458 20818 11464 20852
rect 11418 20780 11464 20818
rect 11418 20746 11424 20780
rect 11458 20746 11464 20780
rect 11418 20708 11464 20746
rect 11418 20674 11424 20708
rect 11458 20674 11464 20708
rect 11418 20636 11464 20674
rect 11418 20602 11424 20636
rect 11458 20602 11464 20636
rect 11418 20564 11464 20602
rect 11418 20530 11424 20564
rect 11458 20530 11464 20564
rect 11418 20492 11464 20530
rect 11418 20458 11424 20492
rect 11458 20458 11464 20492
rect 11418 20420 11464 20458
rect 11418 20386 11424 20420
rect 11458 20386 11464 20420
rect 11418 20348 11464 20386
rect 11418 20314 11424 20348
rect 11458 20314 11464 20348
rect 11418 20276 11464 20314
rect 11418 20242 11424 20276
rect 11458 20242 11464 20276
rect 11418 20204 11464 20242
rect 11418 20170 11424 20204
rect 11458 20170 11464 20204
rect 11418 20132 11464 20170
rect 11418 20098 11424 20132
rect 11458 20098 11464 20132
rect 11418 20060 11464 20098
rect 11418 20026 11424 20060
rect 11458 20026 11464 20060
rect 11418 19988 11464 20026
rect 11418 19954 11424 19988
rect 11458 19954 11464 19988
rect 11418 19916 11464 19954
rect 11418 19882 11424 19916
rect 11458 19882 11464 19916
rect 11418 19844 11464 19882
rect 11418 19810 11424 19844
rect 11458 19810 11464 19844
rect 11418 19772 11464 19810
rect 11418 19738 11424 19772
rect 11458 19738 11464 19772
rect 11418 19700 11464 19738
rect 11418 19666 11424 19700
rect 11458 19666 11464 19700
rect 11418 19628 11464 19666
rect 11418 19594 11424 19628
rect 11458 19594 11464 19628
rect 11418 19556 11464 19594
rect 11418 19522 11424 19556
rect 11458 19522 11464 19556
rect 11418 19484 11464 19522
rect 11418 19450 11424 19484
rect 11458 19450 11464 19484
rect 11418 19412 11464 19450
rect 11418 19378 11424 19412
rect 11458 19378 11464 19412
rect 11418 19340 11464 19378
rect 11418 19306 11424 19340
rect 11458 19306 11464 19340
rect 11418 19268 11464 19306
rect 11418 19234 11424 19268
rect 11458 19234 11464 19268
rect 11418 19196 11464 19234
rect 11418 19162 11424 19196
rect 11458 19162 11464 19196
rect 11418 19124 11464 19162
rect 11418 19090 11424 19124
rect 11458 19090 11464 19124
rect 11418 19052 11464 19090
rect 11418 19018 11424 19052
rect 11458 19018 11464 19052
rect 11418 18980 11464 19018
rect 11418 18946 11424 18980
rect 11458 18946 11464 18980
rect 11418 18908 11464 18946
rect 11418 18874 11424 18908
rect 11458 18874 11464 18908
rect 11418 18836 11464 18874
rect 11418 18802 11424 18836
rect 11458 18802 11464 18836
rect 11418 18764 11464 18802
rect 11418 18730 11424 18764
rect 11458 18730 11464 18764
rect 11418 18692 11464 18730
rect 11418 18658 11424 18692
rect 11458 18658 11464 18692
rect 11418 18620 11464 18658
rect 11418 18586 11424 18620
rect 11458 18586 11464 18620
rect 11418 18548 11464 18586
rect 11418 18514 11424 18548
rect 11458 18514 11464 18548
rect 11418 18476 11464 18514
rect 11418 18442 11424 18476
rect 11458 18442 11464 18476
rect 11418 18404 11464 18442
rect 11418 18370 11424 18404
rect 11458 18370 11464 18404
rect 11418 18332 11464 18370
rect 11418 18298 11424 18332
rect 11458 18298 11464 18332
rect 11418 18260 11464 18298
rect 11418 18226 11424 18260
rect 11458 18226 11464 18260
rect 11418 18188 11464 18226
rect 11418 18154 11424 18188
rect 11458 18154 11464 18188
rect 11418 18116 11464 18154
rect 11418 18082 11424 18116
rect 11458 18082 11464 18116
rect 11418 18044 11464 18082
rect 11418 18010 11424 18044
rect 11458 18010 11464 18044
rect 11418 17972 11464 18010
rect 11418 17938 11424 17972
rect 11458 17938 11464 17972
rect 11418 17900 11464 17938
rect 11418 17866 11424 17900
rect 11458 17866 11464 17900
rect 11418 17828 11464 17866
rect 11418 17794 11424 17828
rect 11458 17794 11464 17828
rect 11418 17756 11464 17794
rect 11418 17722 11424 17756
rect 11458 17722 11464 17756
rect 11418 17684 11464 17722
rect 11418 17650 11424 17684
rect 11458 17650 11464 17684
rect 11418 17612 11464 17650
rect 11418 17578 11424 17612
rect 11458 17578 11464 17612
rect 11418 17540 11464 17578
rect 11418 17506 11424 17540
rect 11458 17506 11464 17540
rect 11418 17468 11464 17506
rect 11418 17434 11424 17468
rect 11458 17434 11464 17468
rect 11418 17396 11464 17434
rect 11418 17362 11424 17396
rect 11458 17362 11464 17396
rect 11418 17324 11464 17362
rect 11418 17290 11424 17324
rect 11458 17290 11464 17324
rect 11418 17252 11464 17290
rect 11418 17218 11424 17252
rect 11458 17218 11464 17252
rect 11418 17180 11464 17218
rect 11418 17146 11424 17180
rect 11458 17146 11464 17180
rect 11418 17108 11464 17146
rect 11418 17074 11424 17108
rect 11458 17074 11464 17108
rect 11418 17036 11464 17074
rect 11418 17002 11424 17036
rect 11458 17002 11464 17036
rect 11418 16964 11464 17002
rect 11418 16930 11424 16964
rect 11458 16930 11464 16964
rect 11418 16892 11464 16930
rect 11418 16858 11424 16892
rect 11458 16858 11464 16892
rect 11418 16820 11464 16858
rect 11418 16786 11424 16820
rect 11458 16786 11464 16820
rect 11418 16748 11464 16786
rect 11418 16714 11424 16748
rect 11458 16714 11464 16748
rect 11418 16676 11464 16714
rect 11418 16642 11424 16676
rect 11458 16642 11464 16676
rect 11418 16604 11464 16642
rect 11418 16570 11424 16604
rect 11458 16570 11464 16604
rect 11418 16532 11464 16570
rect 11418 16498 11424 16532
rect 11458 16498 11464 16532
rect 11418 16460 11464 16498
rect 11418 16426 11424 16460
rect 11458 16426 11464 16460
rect 11418 16388 11464 16426
rect 11418 16354 11424 16388
rect 11458 16354 11464 16388
rect 11418 16316 11464 16354
rect 11418 16282 11424 16316
rect 11458 16282 11464 16316
rect 11418 16244 11464 16282
rect 11418 16210 11424 16244
rect 11458 16210 11464 16244
rect 11418 16172 11464 16210
rect 11418 16138 11424 16172
rect 11458 16138 11464 16172
rect 11418 16100 11464 16138
rect 11418 16066 11424 16100
rect 11458 16066 11464 16100
rect 11418 16028 11464 16066
rect 11418 15994 11424 16028
rect 11458 15994 11464 16028
rect 11418 15956 11464 15994
rect 11418 15922 11424 15956
rect 11458 15922 11464 15956
rect 11418 15884 11464 15922
rect 11418 15850 11424 15884
rect 11458 15850 11464 15884
rect 11418 15812 11464 15850
rect 11418 15778 11424 15812
rect 11458 15778 11464 15812
rect 11418 15740 11464 15778
rect 11418 15706 11424 15740
rect 11458 15706 11464 15740
rect 11418 15668 11464 15706
rect 11418 15634 11424 15668
rect 11458 15634 11464 15668
rect 11418 15596 11464 15634
rect 11418 15562 11424 15596
rect 11458 15562 11464 15596
rect 11418 15524 11464 15562
rect 11418 15490 11424 15524
rect 11458 15490 11464 15524
rect 11418 15452 11464 15490
rect 11418 15418 11424 15452
rect 11458 15418 11464 15452
rect 11418 15380 11464 15418
rect 11418 15346 11424 15380
rect 11458 15346 11464 15380
rect 11418 15308 11464 15346
rect 11418 15274 11424 15308
rect 11458 15274 11464 15308
rect 11418 15236 11464 15274
rect 11418 15202 11424 15236
rect 11458 15202 11464 15236
rect 11418 15164 11464 15202
rect 11418 15130 11424 15164
rect 11458 15130 11464 15164
rect 11418 15092 11464 15130
rect 11418 15058 11424 15092
rect 11458 15058 11464 15092
rect 11418 15020 11464 15058
rect 11418 14986 11424 15020
rect 11458 14986 11464 15020
rect 11418 14948 11464 14986
rect 11418 14914 11424 14948
rect 11458 14914 11464 14948
rect 11418 14876 11464 14914
rect 11418 14842 11424 14876
rect 11458 14842 11464 14876
rect 11418 14804 11464 14842
rect 11418 14770 11424 14804
rect 11458 14770 11464 14804
rect 11418 14732 11464 14770
rect 11418 14698 11424 14732
rect 11458 14698 11464 14732
rect 11418 14660 11464 14698
rect 11418 14626 11424 14660
rect 11458 14626 11464 14660
rect 11418 14588 11464 14626
rect 11418 14554 11424 14588
rect 11458 14554 11464 14588
rect 11418 14516 11464 14554
rect 11418 14482 11424 14516
rect 11458 14482 11464 14516
rect 11418 14444 11464 14482
rect 11418 14410 11424 14444
rect 11458 14410 11464 14444
rect 11418 14372 11464 14410
rect 11418 14338 11424 14372
rect 11458 14338 11464 14372
rect 11418 14300 11464 14338
rect 11418 14266 11424 14300
rect 11458 14266 11464 14300
rect 11418 14228 11464 14266
rect 11418 14194 11424 14228
rect 11458 14194 11464 14228
rect 11418 14156 11464 14194
rect 11418 14122 11424 14156
rect 11458 14122 11464 14156
rect 11418 14084 11464 14122
rect 11418 14050 11424 14084
rect 11458 14050 11464 14084
rect 11418 14012 11464 14050
rect 11418 13978 11424 14012
rect 11458 13978 11464 14012
rect 11418 13940 11464 13978
rect 11418 13906 11424 13940
rect 11458 13906 11464 13940
rect 11418 13868 11464 13906
rect 11418 13834 11424 13868
rect 11458 13834 11464 13868
rect 11418 13796 11464 13834
rect 11418 13762 11424 13796
rect 11458 13762 11464 13796
rect 11418 13724 11464 13762
rect 11418 13690 11424 13724
rect 11458 13690 11464 13724
rect 11418 13652 11464 13690
rect 11418 13618 11424 13652
rect 11458 13618 11464 13652
rect 11418 13580 11464 13618
rect 11418 13546 11424 13580
rect 11458 13546 11464 13580
rect 11418 13508 11464 13546
rect 11418 13474 11424 13508
rect 11458 13474 11464 13508
rect 11418 13436 11464 13474
rect 11418 13402 11424 13436
rect 11458 13402 11464 13436
rect 11418 13364 11464 13402
rect 11418 13330 11424 13364
rect 11458 13330 11464 13364
rect 11418 13292 11464 13330
rect 11418 13258 11424 13292
rect 11458 13258 11464 13292
rect 11418 13220 11464 13258
rect 11418 13186 11424 13220
rect 11458 13186 11464 13220
rect 11418 13148 11464 13186
rect 11418 13114 11424 13148
rect 11458 13114 11464 13148
rect 11418 13076 11464 13114
rect 11418 13042 11424 13076
rect 11458 13042 11464 13076
rect 11418 13004 11464 13042
rect 11418 12970 11424 13004
rect 11458 12970 11464 13004
rect 11418 12932 11464 12970
rect 11418 12898 11424 12932
rect 11458 12898 11464 12932
rect 11418 12860 11464 12898
rect 11418 12826 11424 12860
rect 11458 12826 11464 12860
rect 11418 12788 11464 12826
rect 11418 12754 11424 12788
rect 11458 12754 11464 12788
rect 11418 12716 11464 12754
rect 11418 12682 11424 12716
rect 11458 12682 11464 12716
rect 11418 12644 11464 12682
rect 11418 12610 11424 12644
rect 11458 12610 11464 12644
rect 11418 12572 11464 12610
rect 11418 12538 11424 12572
rect 11458 12538 11464 12572
rect 11418 12500 11464 12538
rect 11418 12466 11424 12500
rect 11458 12466 11464 12500
rect 11418 12428 11464 12466
rect 11418 12394 11424 12428
rect 11458 12394 11464 12428
rect 11418 12356 11464 12394
rect 11418 12322 11424 12356
rect 11458 12322 11464 12356
rect 11418 12284 11464 12322
rect 11418 12250 11424 12284
rect 11458 12250 11464 12284
rect 11418 12212 11464 12250
rect 11418 12178 11424 12212
rect 11458 12178 11464 12212
rect 11418 12140 11464 12178
rect 11418 12106 11424 12140
rect 11458 12106 11464 12140
rect 11418 12068 11464 12106
rect 11418 12034 11424 12068
rect 11458 12034 11464 12068
rect 11418 11996 11464 12034
rect 11418 11962 11424 11996
rect 11458 11962 11464 11996
rect 11418 11924 11464 11962
rect 11418 11890 11424 11924
rect 11458 11890 11464 11924
rect 11418 11852 11464 11890
rect 11418 11818 11424 11852
rect 11458 11818 11464 11852
rect 11418 11780 11464 11818
rect 11418 11746 11424 11780
rect 11458 11746 11464 11780
rect 11418 11708 11464 11746
rect 11418 11674 11424 11708
rect 11458 11674 11464 11708
rect 11418 11636 11464 11674
rect 11418 11602 11424 11636
rect 11458 11602 11464 11636
rect 11418 11564 11464 11602
rect 11418 11530 11424 11564
rect 11458 11530 11464 11564
rect 11418 11492 11464 11530
rect 11418 11458 11424 11492
rect 11458 11458 11464 11492
rect 11418 11420 11464 11458
rect 11418 11386 11424 11420
rect 11458 11386 11464 11420
rect 11418 11348 11464 11386
rect 11418 11314 11424 11348
rect 11458 11314 11464 11348
rect 11418 11276 11464 11314
rect 11418 11242 11424 11276
rect 11458 11242 11464 11276
rect 11418 11204 11464 11242
rect 11418 11170 11424 11204
rect 11458 11170 11464 11204
rect 11418 11132 11464 11170
rect 11418 11098 11424 11132
rect 11458 11098 11464 11132
rect 11418 11060 11464 11098
rect 11418 11026 11424 11060
rect 11458 11026 11464 11060
rect 11418 10988 11464 11026
rect 11418 10954 11424 10988
rect 11458 10954 11464 10988
rect 11418 10916 11464 10954
rect 11418 10882 11424 10916
rect 11458 10882 11464 10916
rect 11418 10844 11464 10882
rect 11418 10810 11424 10844
rect 11458 10810 11464 10844
rect 11418 10772 11464 10810
rect 11418 10738 11424 10772
rect 11458 10738 11464 10772
rect 11418 10700 11464 10738
rect 11418 10666 11424 10700
rect 11458 10666 11464 10700
rect 11418 10628 11464 10666
rect 11418 10594 11424 10628
rect 11458 10594 11464 10628
rect 11418 10556 11464 10594
rect 11418 10522 11424 10556
rect 11458 10522 11464 10556
rect 11418 10484 11464 10522
rect 11418 10450 11424 10484
rect 11458 10450 11464 10484
rect 11418 10412 11464 10450
rect 11418 10378 11424 10412
rect 11458 10378 11464 10412
rect 11418 10340 11464 10378
rect 11418 10306 11424 10340
rect 11458 10306 11464 10340
rect 11418 10268 11464 10306
rect 11418 10234 11424 10268
rect 11458 10234 11464 10268
rect 11418 10196 11464 10234
rect 11418 10162 11424 10196
rect 11458 10162 11464 10196
rect 11418 10124 11464 10162
rect 11418 10090 11424 10124
rect 11458 10090 11464 10124
rect 11418 10052 11464 10090
rect 11418 10018 11424 10052
rect 11458 10018 11464 10052
rect 11418 9980 11464 10018
rect 11418 9946 11424 9980
rect 11458 9946 11464 9980
rect 11418 9908 11464 9946
rect 11418 9874 11424 9908
rect 11458 9874 11464 9908
rect 11418 9836 11464 9874
rect 11418 9802 11424 9836
rect 11458 9802 11464 9836
rect 11418 9764 11464 9802
rect 11418 9730 11424 9764
rect 11458 9730 11464 9764
rect 11418 9692 11464 9730
rect 11418 9658 11424 9692
rect 11458 9658 11464 9692
rect 11418 9620 11464 9658
rect 11418 9586 11424 9620
rect 11458 9586 11464 9620
rect 11418 9548 11464 9586
rect 11418 9514 11424 9548
rect 11458 9514 11464 9548
rect 11418 9476 11464 9514
rect 11418 9442 11424 9476
rect 11458 9442 11464 9476
rect 11418 9404 11464 9442
rect 11418 9370 11424 9404
rect 11458 9370 11464 9404
rect 11418 9332 11464 9370
rect 11418 9298 11424 9332
rect 11458 9298 11464 9332
rect 11418 9260 11464 9298
rect 11418 9226 11424 9260
rect 11458 9226 11464 9260
rect 11418 9188 11464 9226
rect 11418 9154 11424 9188
rect 11458 9154 11464 9188
rect 11418 9116 11464 9154
rect 11418 9082 11424 9116
rect 11458 9082 11464 9116
rect 11418 9044 11464 9082
rect 11418 9010 11424 9044
rect 11458 9010 11464 9044
rect 11418 8972 11464 9010
rect 11418 8938 11424 8972
rect 11458 8938 11464 8972
rect 11418 8900 11464 8938
rect 11418 8866 11424 8900
rect 11458 8866 11464 8900
rect 11418 8828 11464 8866
rect 11418 8794 11424 8828
rect 11458 8794 11464 8828
rect 11418 8756 11464 8794
rect 11418 8722 11424 8756
rect 11458 8722 11464 8756
rect 11418 8684 11464 8722
rect 11418 8650 11424 8684
rect 11458 8650 11464 8684
rect 11418 8612 11464 8650
rect 11418 8578 11424 8612
rect 11458 8578 11464 8612
rect 11418 8540 11464 8578
rect 11418 8506 11424 8540
rect 11458 8506 11464 8540
rect 11418 8468 11464 8506
rect 11418 8434 11424 8468
rect 11458 8434 11464 8468
rect 11418 8396 11464 8434
rect 11418 8362 11424 8396
rect 11458 8362 11464 8396
rect 11418 8324 11464 8362
rect 11418 8290 11424 8324
rect 11458 8290 11464 8324
rect 11418 8252 11464 8290
rect 11418 8218 11424 8252
rect 11458 8218 11464 8252
rect 11418 8180 11464 8218
rect 11418 8146 11424 8180
rect 11458 8146 11464 8180
rect 11418 8108 11464 8146
rect 11418 8074 11424 8108
rect 11458 8074 11464 8108
rect 11418 8036 11464 8074
rect 11418 8002 11424 8036
rect 11458 8002 11464 8036
rect 11418 7964 11464 8002
rect 11418 7930 11424 7964
rect 11458 7930 11464 7964
rect 11418 7892 11464 7930
rect 11418 7858 11424 7892
rect 11458 7858 11464 7892
rect 11418 7820 11464 7858
rect 11418 7786 11424 7820
rect 11458 7786 11464 7820
rect 11418 7748 11464 7786
rect 11418 7714 11424 7748
rect 11458 7714 11464 7748
rect 11418 7676 11464 7714
rect 11418 7642 11424 7676
rect 11458 7642 11464 7676
rect 11418 7604 11464 7642
rect 11418 7570 11424 7604
rect 11458 7570 11464 7604
rect 11418 7532 11464 7570
rect 11418 7498 11424 7532
rect 11458 7498 11464 7532
rect 11418 7460 11464 7498
rect 11418 7426 11424 7460
rect 11458 7426 11464 7460
rect 11418 7388 11464 7426
rect 11418 7354 11424 7388
rect 11458 7354 11464 7388
rect 11418 7316 11464 7354
rect 11418 7282 11424 7316
rect 11458 7282 11464 7316
rect 11418 7244 11464 7282
rect 11418 7210 11424 7244
rect 11458 7210 11464 7244
rect 11418 7172 11464 7210
rect 11418 7138 11424 7172
rect 11458 7138 11464 7172
rect 11418 7100 11464 7138
rect 11418 7066 11424 7100
rect 11458 7066 11464 7100
rect 11418 7028 11464 7066
rect 11418 6994 11424 7028
rect 11458 6994 11464 7028
rect 11418 6956 11464 6994
rect 11418 6922 11424 6956
rect 11458 6922 11464 6956
rect 11418 6884 11464 6922
rect 11418 6850 11424 6884
rect 11458 6850 11464 6884
rect 11418 6812 11464 6850
rect 11418 6778 11424 6812
rect 11458 6778 11464 6812
rect 11418 6740 11464 6778
rect 11418 6706 11424 6740
rect 11458 6706 11464 6740
rect 11418 6668 11464 6706
rect 11418 6634 11424 6668
rect 11458 6634 11464 6668
rect 11418 6596 11464 6634
rect 11418 6562 11424 6596
rect 11458 6562 11464 6596
rect 11418 6524 11464 6562
rect 11418 6490 11424 6524
rect 11458 6490 11464 6524
rect 11418 6452 11464 6490
rect 11418 6418 11424 6452
rect 11458 6418 11464 6452
rect 11418 6380 11464 6418
rect 11418 6346 11424 6380
rect 11458 6346 11464 6380
rect 11418 6308 11464 6346
rect 11418 6274 11424 6308
rect 11458 6274 11464 6308
rect 11418 6236 11464 6274
rect 11418 6202 11424 6236
rect 11458 6202 11464 6236
rect 11418 6164 11464 6202
rect 11418 6130 11424 6164
rect 11458 6130 11464 6164
rect 11418 6092 11464 6130
rect 11418 6058 11424 6092
rect 11458 6058 11464 6092
rect 11418 6020 11464 6058
rect 11418 5986 11424 6020
rect 11458 5986 11464 6020
rect 11418 5948 11464 5986
rect 11418 5914 11424 5948
rect 11458 5914 11464 5948
rect 11418 5876 11464 5914
rect 11418 5842 11424 5876
rect 11458 5842 11464 5876
rect 11418 5804 11464 5842
rect 11418 5770 11424 5804
rect 11458 5770 11464 5804
rect 11418 5732 11464 5770
rect 11418 5698 11424 5732
rect 11458 5698 11464 5732
rect 11418 5660 11464 5698
rect 11418 5626 11424 5660
rect 11458 5626 11464 5660
rect 11418 5588 11464 5626
rect 11418 5554 11424 5588
rect 11458 5554 11464 5588
rect 11418 5516 11464 5554
rect 11418 5482 11424 5516
rect 11458 5482 11464 5516
rect 11418 5444 11464 5482
rect 11418 5410 11424 5444
rect 11458 5410 11464 5444
rect 11418 5372 11464 5410
rect 11418 5338 11424 5372
rect 11458 5338 11464 5372
rect 11418 5300 11464 5338
rect 11418 5266 11424 5300
rect 11458 5266 11464 5300
rect 11418 5228 11464 5266
rect 11418 5194 11424 5228
rect 11458 5194 11464 5228
rect 11418 5156 11464 5194
rect 11418 5122 11424 5156
rect 11458 5122 11464 5156
rect 11418 5084 11464 5122
rect 11418 5050 11424 5084
rect 11458 5050 11464 5084
rect 11418 5012 11464 5050
rect 11418 4978 11424 5012
rect 11458 4978 11464 5012
rect 11418 4940 11464 4978
rect 11418 4906 11424 4940
rect 11458 4906 11464 4940
rect 11418 4868 11464 4906
rect 11418 4834 11424 4868
rect 11458 4834 11464 4868
rect 11418 4796 11464 4834
rect 11418 4762 11424 4796
rect 11458 4762 11464 4796
rect 11418 4724 11464 4762
rect 11418 4690 11424 4724
rect 11458 4690 11464 4724
rect 11418 4652 11464 4690
rect 11418 4618 11424 4652
rect 11458 4618 11464 4652
rect 11418 4580 11464 4618
rect 11418 4546 11424 4580
rect 11458 4546 11464 4580
rect 11418 4508 11464 4546
rect 11418 4474 11424 4508
rect 11458 4474 11464 4508
rect 11418 4436 11464 4474
rect 11418 4402 11424 4436
rect 11458 4402 11464 4436
rect 11418 4364 11464 4402
rect 11418 4330 11424 4364
rect 11458 4330 11464 4364
rect 11418 4292 11464 4330
rect 11418 4258 11424 4292
rect 11458 4258 11464 4292
rect 11418 4220 11464 4258
rect 11418 4186 11424 4220
rect 11458 4186 11464 4220
rect 11418 4148 11464 4186
rect 11418 4114 11424 4148
rect 11458 4114 11464 4148
rect 11418 4076 11464 4114
rect 11418 4042 11424 4076
rect 11458 4042 11464 4076
rect 11418 4004 11464 4042
rect 11418 3970 11424 4004
rect 11458 3970 11464 4004
rect 11418 3932 11464 3970
rect 11418 3898 11424 3932
rect 11458 3898 11464 3932
rect 11418 3860 11464 3898
rect 11418 3826 11424 3860
rect 11458 3826 11464 3860
rect 11418 3788 11464 3826
rect 11418 3754 11424 3788
rect 11458 3754 11464 3788
rect 11418 3716 11464 3754
rect 11418 3682 11424 3716
rect 11458 3682 11464 3716
rect 11418 3644 11464 3682
rect 11418 3610 11424 3644
rect 11458 3610 11464 3644
rect 11418 3572 11464 3610
rect 11418 3538 11424 3572
rect 11458 3538 11464 3572
rect 11418 3500 11464 3538
rect 10220 3428 10266 3466
rect 10220 3394 10226 3428
rect 10260 3394 10266 3428
rect 9082 3322 9088 3356
rect 9122 3322 9128 3356
rect 9082 3284 9128 3322
rect 9082 3250 9088 3284
rect 9122 3250 9128 3284
rect 10220 3356 10266 3394
rect 10403 3493 10455 3499
rect 10403 3429 10455 3441
rect 10403 3369 10455 3377
rect 10521 3487 10691 3499
rect 10521 3453 10530 3487
rect 10564 3453 10648 3487
rect 10682 3453 10691 3487
rect 10521 3415 10691 3453
rect 10521 3381 10530 3415
rect 10564 3381 10648 3415
rect 10682 3381 10691 3415
rect 10521 3369 10691 3381
rect 10757 3487 10927 3499
rect 10757 3453 10766 3487
rect 10800 3453 10884 3487
rect 10918 3453 10927 3487
rect 10757 3415 10927 3453
rect 10757 3381 10766 3415
rect 10800 3381 10884 3415
rect 10918 3381 10927 3415
rect 10757 3369 10927 3381
rect 10993 3487 11163 3499
rect 10993 3453 11002 3487
rect 11036 3453 11120 3487
rect 11154 3453 11163 3487
rect 10993 3415 11163 3453
rect 10993 3381 11002 3415
rect 11036 3381 11120 3415
rect 11154 3381 11163 3415
rect 10993 3369 11163 3381
rect 11229 3493 11281 3499
rect 11229 3429 11281 3441
rect 11229 3369 11281 3377
rect 11418 3466 11424 3500
rect 11458 3466 11464 3500
rect 13206 38465 13252 38504
rect 13386 38612 13412 38624
rect 13464 38615 13526 38624
rect 13386 38578 13392 38612
rect 13464 38581 13466 38615
rect 13500 38581 13526 38615
rect 13386 38572 13412 38578
rect 13464 38572 13526 38581
rect 13578 38572 13584 38624
rect 14934 38612 14980 38650
rect 14934 38578 14940 38612
rect 14974 38578 14980 38612
rect 13386 38540 13434 38572
tri 13434 38540 13466 38572 nw
rect 14934 38540 14980 38578
rect 13386 38517 13432 38540
tri 13432 38538 13434 38540 nw
rect 13386 38483 13392 38517
rect 13426 38483 13432 38517
rect 13386 38471 13432 38483
rect 14934 38506 14940 38540
rect 14974 38506 14980 38540
rect 13206 38431 13212 38465
rect 13246 38431 13252 38465
rect 13206 38392 13252 38431
rect 13206 38358 13212 38392
rect 13246 38358 13252 38392
rect 13206 38319 13252 38358
rect 13206 38285 13212 38319
rect 13246 38285 13252 38319
rect 13206 38246 13252 38285
rect 13206 38212 13212 38246
rect 13246 38212 13252 38246
rect 13206 38173 13252 38212
rect 13206 38139 13212 38173
rect 13246 38139 13252 38173
rect 13206 38100 13252 38139
rect 13206 38066 13212 38100
rect 13246 38066 13252 38100
rect 13206 38027 13252 38066
rect 13206 37993 13212 38027
rect 13246 37993 13252 38027
rect 13206 37954 13252 37993
rect 13206 37920 13212 37954
rect 13246 37920 13252 37954
rect 13206 37881 13252 37920
rect 13206 37847 13212 37881
rect 13246 37847 13252 37881
rect 13206 37808 13252 37847
rect 13206 37774 13212 37808
rect 13246 37774 13252 37808
rect 13206 37735 13252 37774
rect 13206 37701 13212 37735
rect 13246 37701 13252 37735
rect 13206 37662 13252 37701
rect 13206 37628 13212 37662
rect 13246 37628 13252 37662
rect 13206 37589 13252 37628
rect 13206 37555 13212 37589
rect 13246 37555 13252 37589
rect 13206 37516 13252 37555
rect 13206 37482 13212 37516
rect 13246 37482 13252 37516
rect 13206 37443 13252 37482
rect 13206 37409 13212 37443
rect 13246 37409 13252 37443
rect 13206 37370 13252 37409
rect 13206 37336 13212 37370
rect 13246 37336 13252 37370
rect 13206 37298 13252 37336
rect 13206 37264 13212 37298
rect 13246 37264 13252 37298
rect 13206 37226 13252 37264
rect 13206 37192 13212 37226
rect 13246 37192 13252 37226
rect 13206 37154 13252 37192
rect 13206 37120 13212 37154
rect 13246 37120 13252 37154
rect 13206 37082 13252 37120
rect 13206 37048 13212 37082
rect 13246 37048 13252 37082
rect 13206 37010 13252 37048
rect 13206 36976 13212 37010
rect 13246 36976 13252 37010
rect 13206 36938 13252 36976
rect 13206 36904 13212 36938
rect 13246 36904 13252 36938
rect 13206 36866 13252 36904
rect 13206 36832 13212 36866
rect 13246 36832 13252 36866
rect 13206 36794 13252 36832
rect 13206 36760 13212 36794
rect 13246 36760 13252 36794
rect 13206 36722 13252 36760
rect 13206 36688 13212 36722
rect 13246 36688 13252 36722
rect 13206 36650 13252 36688
rect 13206 36616 13212 36650
rect 13246 36616 13252 36650
rect 13206 36578 13252 36616
rect 13206 36544 13212 36578
rect 13246 36544 13252 36578
rect 13206 36506 13252 36544
rect 13206 36472 13212 36506
rect 13246 36472 13252 36506
rect 13206 36434 13252 36472
rect 13206 36400 13212 36434
rect 13246 36400 13252 36434
rect 13206 36362 13252 36400
rect 13206 36328 13212 36362
rect 13246 36328 13252 36362
rect 13206 36290 13252 36328
rect 13206 36256 13212 36290
rect 13246 36256 13252 36290
rect 13206 36218 13252 36256
rect 13206 36184 13212 36218
rect 13246 36184 13252 36218
rect 13206 36146 13252 36184
rect 13206 36112 13212 36146
rect 13246 36112 13252 36146
rect 13206 36074 13252 36112
rect 13206 36040 13212 36074
rect 13246 36040 13252 36074
rect 13206 36002 13252 36040
rect 13206 35968 13212 36002
rect 13246 35968 13252 36002
rect 13206 35930 13252 35968
rect 13206 35896 13212 35930
rect 13246 35896 13252 35930
rect 13206 35858 13252 35896
rect 13206 35824 13212 35858
rect 13246 35824 13252 35858
rect 13206 35786 13252 35824
rect 13206 35752 13212 35786
rect 13246 35752 13252 35786
rect 13206 35714 13252 35752
rect 13206 35680 13212 35714
rect 13246 35680 13252 35714
rect 13206 35642 13252 35680
rect 13206 35608 13212 35642
rect 13246 35608 13252 35642
rect 13206 35570 13252 35608
rect 13206 35536 13212 35570
rect 13246 35536 13252 35570
rect 13206 35498 13252 35536
rect 13206 35464 13212 35498
rect 13246 35464 13252 35498
rect 13206 35426 13252 35464
rect 13206 35392 13212 35426
rect 13246 35392 13252 35426
rect 13206 35354 13252 35392
rect 13206 35320 13212 35354
rect 13246 35320 13252 35354
rect 13206 35282 13252 35320
rect 13206 35248 13212 35282
rect 13246 35248 13252 35282
rect 13206 35210 13252 35248
rect 13206 35176 13212 35210
rect 13246 35176 13252 35210
rect 13206 35138 13252 35176
rect 13206 35104 13212 35138
rect 13246 35104 13252 35138
rect 13206 35066 13252 35104
rect 13206 35032 13212 35066
rect 13246 35032 13252 35066
rect 13206 34994 13252 35032
rect 13206 34960 13212 34994
rect 13246 34960 13252 34994
rect 13206 34922 13252 34960
rect 13206 34888 13212 34922
rect 13246 34888 13252 34922
rect 13206 34850 13252 34888
rect 13206 34816 13212 34850
rect 13246 34816 13252 34850
rect 13206 34778 13252 34816
rect 13206 34744 13212 34778
rect 13246 34744 13252 34778
rect 13206 34706 13252 34744
rect 13206 34672 13212 34706
rect 13246 34672 13252 34706
rect 13206 34634 13252 34672
rect 13206 34600 13212 34634
rect 13246 34600 13252 34634
rect 13206 34562 13252 34600
rect 13206 34528 13212 34562
rect 13246 34528 13252 34562
rect 13206 34490 13252 34528
rect 13206 34456 13212 34490
rect 13246 34456 13252 34490
rect 13206 34418 13252 34456
rect 13206 34384 13212 34418
rect 13246 34384 13252 34418
rect 13206 34346 13252 34384
rect 13206 34312 13212 34346
rect 13246 34312 13252 34346
rect 13206 34274 13252 34312
rect 13206 34240 13212 34274
rect 13246 34240 13252 34274
rect 13206 34202 13252 34240
rect 13206 34168 13212 34202
rect 13246 34168 13252 34202
rect 13206 34130 13252 34168
rect 13206 34096 13212 34130
rect 13246 34096 13252 34130
rect 13206 34058 13252 34096
rect 13206 34024 13212 34058
rect 13246 34024 13252 34058
rect 13206 33986 13252 34024
rect 13206 33952 13212 33986
rect 13246 33952 13252 33986
rect 13206 33914 13252 33952
rect 13206 33880 13212 33914
rect 13246 33880 13252 33914
rect 13206 33842 13252 33880
rect 13206 33808 13212 33842
rect 13246 33808 13252 33842
rect 13206 33770 13252 33808
rect 13206 33736 13212 33770
rect 13246 33736 13252 33770
rect 13206 33698 13252 33736
rect 13206 33664 13212 33698
rect 13246 33664 13252 33698
rect 13206 33626 13252 33664
rect 13206 33592 13212 33626
rect 13246 33592 13252 33626
rect 13206 33554 13252 33592
rect 13206 33520 13212 33554
rect 13246 33520 13252 33554
rect 13206 33482 13252 33520
rect 13206 33448 13212 33482
rect 13246 33448 13252 33482
rect 13206 33410 13252 33448
rect 13206 33376 13212 33410
rect 13246 33376 13252 33410
rect 13206 33338 13252 33376
rect 13206 33304 13212 33338
rect 13246 33304 13252 33338
rect 13206 33266 13252 33304
rect 13206 33232 13212 33266
rect 13246 33232 13252 33266
rect 13206 33194 13252 33232
rect 13206 33160 13212 33194
rect 13246 33160 13252 33194
rect 13206 33122 13252 33160
rect 13206 33088 13212 33122
rect 13246 33088 13252 33122
rect 13206 33050 13252 33088
rect 13206 33016 13212 33050
rect 13246 33016 13252 33050
rect 13206 32978 13252 33016
rect 13206 32944 13212 32978
rect 13246 32944 13252 32978
rect 13206 32906 13252 32944
rect 13206 32872 13212 32906
rect 13246 32872 13252 32906
rect 13206 32834 13252 32872
rect 13206 32800 13212 32834
rect 13246 32800 13252 32834
rect 13206 32762 13252 32800
rect 13206 32728 13212 32762
rect 13246 32728 13252 32762
rect 13206 32690 13252 32728
rect 13206 32656 13212 32690
rect 13246 32656 13252 32690
rect 13206 32618 13252 32656
rect 13206 32584 13212 32618
rect 13246 32584 13252 32618
rect 13206 32546 13252 32584
rect 13206 32512 13212 32546
rect 13246 32512 13252 32546
rect 13206 32474 13252 32512
rect 13206 32440 13212 32474
rect 13246 32440 13252 32474
rect 13206 32402 13252 32440
rect 13206 32368 13212 32402
rect 13246 32368 13252 32402
rect 13206 32330 13252 32368
rect 13206 32296 13212 32330
rect 13246 32296 13252 32330
rect 13206 32258 13252 32296
rect 13206 32224 13212 32258
rect 13246 32224 13252 32258
rect 13206 32186 13252 32224
rect 13206 32152 13212 32186
rect 13246 32152 13252 32186
rect 13206 32114 13252 32152
rect 13206 32080 13212 32114
rect 13246 32080 13252 32114
rect 13206 32042 13252 32080
rect 13206 32008 13212 32042
rect 13246 32008 13252 32042
rect 13206 31970 13252 32008
rect 13206 31936 13212 31970
rect 13246 31936 13252 31970
rect 13206 31898 13252 31936
rect 13206 31864 13212 31898
rect 13246 31864 13252 31898
rect 13206 31826 13252 31864
rect 13206 31792 13212 31826
rect 13246 31792 13252 31826
rect 13206 31754 13252 31792
rect 13206 31720 13212 31754
rect 13246 31720 13252 31754
rect 13206 31682 13252 31720
rect 13206 31648 13212 31682
rect 13246 31648 13252 31682
rect 13206 31610 13252 31648
rect 13206 31576 13212 31610
rect 13246 31576 13252 31610
rect 13206 31538 13252 31576
rect 13206 31504 13212 31538
rect 13246 31504 13252 31538
rect 13206 31466 13252 31504
rect 13206 31432 13212 31466
rect 13246 31432 13252 31466
rect 13206 31394 13252 31432
rect 13206 31360 13212 31394
rect 13246 31360 13252 31394
rect 13206 31322 13252 31360
rect 13206 31288 13212 31322
rect 13246 31288 13252 31322
rect 13206 31250 13252 31288
rect 13206 31216 13212 31250
rect 13246 31216 13252 31250
rect 13206 31178 13252 31216
rect 13206 31144 13212 31178
rect 13246 31144 13252 31178
rect 13206 31106 13252 31144
rect 13206 31072 13212 31106
rect 13246 31072 13252 31106
rect 13206 31034 13252 31072
rect 13206 31000 13212 31034
rect 13246 31000 13252 31034
rect 13206 30962 13252 31000
rect 13206 30928 13212 30962
rect 13246 30928 13252 30962
rect 13206 30890 13252 30928
rect 13206 30856 13212 30890
rect 13246 30856 13252 30890
rect 13206 30818 13252 30856
rect 13206 30784 13212 30818
rect 13246 30784 13252 30818
rect 13206 30746 13252 30784
rect 13206 30712 13212 30746
rect 13246 30712 13252 30746
rect 13206 30674 13252 30712
rect 13206 30640 13212 30674
rect 13246 30640 13252 30674
rect 13206 30602 13252 30640
rect 13206 30568 13212 30602
rect 13246 30568 13252 30602
rect 13206 30530 13252 30568
rect 13206 30496 13212 30530
rect 13246 30496 13252 30530
rect 13206 30458 13252 30496
rect 13206 30424 13212 30458
rect 13246 30424 13252 30458
rect 13206 30386 13252 30424
rect 13206 30352 13212 30386
rect 13246 30352 13252 30386
rect 13206 30314 13252 30352
rect 13206 30280 13212 30314
rect 13246 30280 13252 30314
rect 13206 30242 13252 30280
rect 13206 30208 13212 30242
rect 13246 30208 13252 30242
rect 13206 30170 13252 30208
rect 13206 30136 13212 30170
rect 13246 30136 13252 30170
rect 13206 30098 13252 30136
rect 13206 30064 13212 30098
rect 13246 30064 13252 30098
rect 13206 30026 13252 30064
rect 13206 29992 13212 30026
rect 13246 29992 13252 30026
rect 13206 29954 13252 29992
rect 13206 29920 13212 29954
rect 13246 29920 13252 29954
rect 13206 29882 13252 29920
rect 13206 29848 13212 29882
rect 13246 29848 13252 29882
rect 13206 29810 13252 29848
rect 13206 29776 13212 29810
rect 13246 29776 13252 29810
rect 13206 29738 13252 29776
rect 13206 29704 13212 29738
rect 13246 29704 13252 29738
rect 13206 29666 13252 29704
rect 13206 29632 13212 29666
rect 13246 29632 13252 29666
rect 13206 29594 13252 29632
rect 13206 29560 13212 29594
rect 13246 29560 13252 29594
rect 13206 29522 13252 29560
rect 13206 29488 13212 29522
rect 13246 29488 13252 29522
rect 13206 29450 13252 29488
rect 13206 29416 13212 29450
rect 13246 29416 13252 29450
rect 13206 29378 13252 29416
rect 13206 29344 13212 29378
rect 13246 29344 13252 29378
rect 13206 29306 13252 29344
rect 13206 29272 13212 29306
rect 13246 29272 13252 29306
rect 13206 29234 13252 29272
rect 13206 29200 13212 29234
rect 13246 29200 13252 29234
rect 13206 29162 13252 29200
rect 13206 29128 13212 29162
rect 13246 29128 13252 29162
rect 13206 29090 13252 29128
rect 13206 29056 13212 29090
rect 13246 29056 13252 29090
rect 13206 29018 13252 29056
rect 13206 28984 13212 29018
rect 13246 28984 13252 29018
rect 13206 28946 13252 28984
rect 13206 28912 13212 28946
rect 13246 28912 13252 28946
rect 13206 28874 13252 28912
rect 13206 28840 13212 28874
rect 13246 28840 13252 28874
rect 13206 28802 13252 28840
rect 13206 28768 13212 28802
rect 13246 28768 13252 28802
rect 13206 28730 13252 28768
rect 13206 28696 13212 28730
rect 13246 28696 13252 28730
rect 13206 28658 13252 28696
rect 13206 28624 13212 28658
rect 13246 28624 13252 28658
rect 13206 28586 13252 28624
rect 13206 28552 13212 28586
rect 13246 28552 13252 28586
rect 13206 28514 13252 28552
rect 13206 28480 13212 28514
rect 13246 28480 13252 28514
rect 13206 28442 13252 28480
rect 13206 28408 13212 28442
rect 13246 28408 13252 28442
rect 13206 28370 13252 28408
rect 13206 28336 13212 28370
rect 13246 28336 13252 28370
rect 13206 28298 13252 28336
rect 13206 28264 13212 28298
rect 13246 28264 13252 28298
rect 13206 28226 13252 28264
rect 13206 28192 13212 28226
rect 13246 28192 13252 28226
rect 13206 28154 13252 28192
rect 13206 28120 13212 28154
rect 13246 28120 13252 28154
rect 13206 28082 13252 28120
rect 13206 28048 13212 28082
rect 13246 28048 13252 28082
rect 13206 28010 13252 28048
rect 13206 27976 13212 28010
rect 13246 27976 13252 28010
rect 13206 27938 13252 27976
rect 13206 27904 13212 27938
rect 13246 27904 13252 27938
rect 13206 27866 13252 27904
rect 13206 27832 13212 27866
rect 13246 27832 13252 27866
rect 13206 27794 13252 27832
rect 13206 27760 13212 27794
rect 13246 27760 13252 27794
rect 13206 27722 13252 27760
rect 13206 27688 13212 27722
rect 13246 27688 13252 27722
rect 13206 27650 13252 27688
rect 13206 27616 13212 27650
rect 13246 27616 13252 27650
rect 13206 27578 13252 27616
rect 13206 27544 13212 27578
rect 13246 27544 13252 27578
rect 13206 27506 13252 27544
rect 13206 27472 13212 27506
rect 13246 27472 13252 27506
rect 13206 27434 13252 27472
rect 13206 27400 13212 27434
rect 13246 27400 13252 27434
rect 13206 27362 13252 27400
rect 13206 27328 13212 27362
rect 13246 27328 13252 27362
rect 13206 27290 13252 27328
rect 13206 27256 13212 27290
rect 13246 27256 13252 27290
rect 13206 27218 13252 27256
rect 13206 27184 13212 27218
rect 13246 27184 13252 27218
rect 13206 27146 13252 27184
rect 13206 27112 13212 27146
rect 13246 27112 13252 27146
rect 13206 27074 13252 27112
rect 13206 27040 13212 27074
rect 13246 27040 13252 27074
rect 13206 27002 13252 27040
rect 13206 26968 13212 27002
rect 13246 26968 13252 27002
rect 13206 26930 13252 26968
rect 13206 26896 13212 26930
rect 13246 26896 13252 26930
rect 13206 26858 13252 26896
rect 13206 26824 13212 26858
rect 13246 26824 13252 26858
rect 13206 26786 13252 26824
rect 13206 26752 13212 26786
rect 13246 26752 13252 26786
rect 13206 26714 13252 26752
rect 13206 26680 13212 26714
rect 13246 26680 13252 26714
rect 13206 26642 13252 26680
rect 13206 26608 13212 26642
rect 13246 26608 13252 26642
rect 13206 26570 13252 26608
rect 13206 26536 13212 26570
rect 13246 26536 13252 26570
rect 13206 26498 13252 26536
rect 13206 26464 13212 26498
rect 13246 26464 13252 26498
rect 13206 26426 13252 26464
rect 13206 26392 13212 26426
rect 13246 26392 13252 26426
rect 13206 26354 13252 26392
rect 13206 26320 13212 26354
rect 13246 26320 13252 26354
rect 13206 26282 13252 26320
rect 13206 26248 13212 26282
rect 13246 26248 13252 26282
rect 13206 26210 13252 26248
rect 13206 26176 13212 26210
rect 13246 26176 13252 26210
rect 13206 26138 13252 26176
rect 13206 26104 13212 26138
rect 13246 26104 13252 26138
rect 13206 26066 13252 26104
rect 13206 26032 13212 26066
rect 13246 26032 13252 26066
rect 13206 25994 13252 26032
rect 13206 25960 13212 25994
rect 13246 25960 13252 25994
rect 13206 25922 13252 25960
rect 13206 25888 13212 25922
rect 13246 25888 13252 25922
rect 13206 25850 13252 25888
rect 13206 25816 13212 25850
rect 13246 25816 13252 25850
rect 13206 25778 13252 25816
rect 13206 25744 13212 25778
rect 13246 25744 13252 25778
rect 13206 25706 13252 25744
rect 13206 25672 13212 25706
rect 13246 25672 13252 25706
rect 13206 25634 13252 25672
rect 13206 25600 13212 25634
rect 13246 25600 13252 25634
rect 13206 25562 13252 25600
rect 13206 25528 13212 25562
rect 13246 25528 13252 25562
rect 13206 25490 13252 25528
rect 13206 25456 13212 25490
rect 13246 25456 13252 25490
rect 13206 25418 13252 25456
rect 13206 25384 13212 25418
rect 13246 25384 13252 25418
rect 13206 25346 13252 25384
rect 13206 25312 13212 25346
rect 13246 25312 13252 25346
rect 13206 25274 13252 25312
rect 13206 25240 13212 25274
rect 13246 25240 13252 25274
rect 13206 25202 13252 25240
rect 13206 25168 13212 25202
rect 13246 25168 13252 25202
rect 13206 25130 13252 25168
rect 13206 25096 13212 25130
rect 13246 25096 13252 25130
rect 13206 25058 13252 25096
rect 13206 25024 13212 25058
rect 13246 25024 13252 25058
rect 13206 24986 13252 25024
rect 13206 24952 13212 24986
rect 13246 24952 13252 24986
rect 13206 24914 13252 24952
rect 13206 24880 13212 24914
rect 13246 24880 13252 24914
rect 13206 24842 13252 24880
rect 13206 24808 13212 24842
rect 13246 24808 13252 24842
rect 13206 24770 13252 24808
rect 13206 24736 13212 24770
rect 13246 24736 13252 24770
rect 13206 24698 13252 24736
rect 13206 24664 13212 24698
rect 13246 24664 13252 24698
rect 13206 24626 13252 24664
rect 13206 24592 13212 24626
rect 13246 24592 13252 24626
rect 13206 24554 13252 24592
rect 13206 24520 13212 24554
rect 13246 24520 13252 24554
rect 13206 24482 13252 24520
rect 13206 24448 13212 24482
rect 13246 24448 13252 24482
rect 13206 24410 13252 24448
rect 13206 24376 13212 24410
rect 13246 24376 13252 24410
rect 13206 24338 13252 24376
rect 13206 24304 13212 24338
rect 13246 24304 13252 24338
rect 13206 24266 13252 24304
rect 13206 24232 13212 24266
rect 13246 24232 13252 24266
rect 13206 24194 13252 24232
rect 13206 24160 13212 24194
rect 13246 24160 13252 24194
rect 13206 24122 13252 24160
rect 13206 24088 13212 24122
rect 13246 24088 13252 24122
rect 13206 24050 13252 24088
rect 13206 24016 13212 24050
rect 13246 24016 13252 24050
rect 13206 23978 13252 24016
rect 13206 23944 13212 23978
rect 13246 23944 13252 23978
rect 13206 23906 13252 23944
rect 13206 23872 13212 23906
rect 13246 23872 13252 23906
rect 13206 23834 13252 23872
rect 13206 23800 13212 23834
rect 13246 23800 13252 23834
rect 13206 23762 13252 23800
rect 13206 23728 13212 23762
rect 13246 23728 13252 23762
rect 13206 23690 13252 23728
rect 13206 23656 13212 23690
rect 13246 23656 13252 23690
rect 13206 23618 13252 23656
rect 13206 23584 13212 23618
rect 13246 23584 13252 23618
rect 13206 23546 13252 23584
rect 13206 23512 13212 23546
rect 13246 23512 13252 23546
rect 13206 23474 13252 23512
rect 13206 23440 13212 23474
rect 13246 23440 13252 23474
rect 13206 23402 13252 23440
rect 13206 23368 13212 23402
rect 13246 23368 13252 23402
rect 13206 23330 13252 23368
rect 13206 23296 13212 23330
rect 13246 23296 13252 23330
rect 13206 23258 13252 23296
rect 13206 23224 13212 23258
rect 13246 23224 13252 23258
rect 13206 23186 13252 23224
rect 13206 23152 13212 23186
rect 13246 23152 13252 23186
rect 13206 23114 13252 23152
rect 13206 23080 13212 23114
rect 13246 23080 13252 23114
rect 13206 23042 13252 23080
rect 13206 23008 13212 23042
rect 13246 23008 13252 23042
rect 13206 22970 13252 23008
rect 13206 22936 13212 22970
rect 13246 22936 13252 22970
rect 13206 22898 13252 22936
rect 13206 22864 13212 22898
rect 13246 22864 13252 22898
rect 13206 22826 13252 22864
rect 13206 22792 13212 22826
rect 13246 22792 13252 22826
rect 13206 22754 13252 22792
rect 13206 22720 13212 22754
rect 13246 22720 13252 22754
rect 13206 22682 13252 22720
rect 13206 22648 13212 22682
rect 13246 22648 13252 22682
rect 13206 22610 13252 22648
rect 13206 22576 13212 22610
rect 13246 22576 13252 22610
rect 13206 22538 13252 22576
rect 13206 22504 13212 22538
rect 13246 22504 13252 22538
rect 13206 22466 13252 22504
rect 13206 22432 13212 22466
rect 13246 22432 13252 22466
rect 13206 22394 13252 22432
rect 13206 22360 13212 22394
rect 13246 22360 13252 22394
rect 13206 22322 13252 22360
rect 13206 22288 13212 22322
rect 13246 22288 13252 22322
rect 13206 22250 13252 22288
rect 13206 22216 13212 22250
rect 13246 22216 13252 22250
rect 13206 22178 13252 22216
rect 13206 22144 13212 22178
rect 13246 22144 13252 22178
rect 13206 22106 13252 22144
rect 13206 22072 13212 22106
rect 13246 22072 13252 22106
rect 13206 22034 13252 22072
rect 13206 22000 13212 22034
rect 13246 22000 13252 22034
rect 13206 21962 13252 22000
rect 13206 21928 13212 21962
rect 13246 21928 13252 21962
rect 13206 21890 13252 21928
rect 13206 21856 13212 21890
rect 13246 21856 13252 21890
rect 13206 21818 13252 21856
rect 13206 21784 13212 21818
rect 13246 21784 13252 21818
rect 13206 21746 13252 21784
rect 13206 21712 13212 21746
rect 13246 21712 13252 21746
rect 13206 21674 13252 21712
rect 13206 21640 13212 21674
rect 13246 21640 13252 21674
rect 13206 21602 13252 21640
rect 13206 21568 13212 21602
rect 13246 21568 13252 21602
rect 13206 21530 13252 21568
rect 13206 21496 13212 21530
rect 13246 21496 13252 21530
rect 13206 21458 13252 21496
rect 13206 21424 13212 21458
rect 13246 21424 13252 21458
rect 13206 21386 13252 21424
rect 13206 21352 13212 21386
rect 13246 21352 13252 21386
rect 13206 21314 13252 21352
rect 13206 21280 13212 21314
rect 13246 21280 13252 21314
rect 13206 21242 13252 21280
rect 13206 21208 13212 21242
rect 13246 21208 13252 21242
rect 13206 21170 13252 21208
rect 13206 21136 13212 21170
rect 13246 21136 13252 21170
rect 13206 21098 13252 21136
rect 13206 21064 13212 21098
rect 13246 21064 13252 21098
rect 13206 21026 13252 21064
rect 13206 20992 13212 21026
rect 13246 20992 13252 21026
rect 13206 20954 13252 20992
rect 13206 20920 13212 20954
rect 13246 20920 13252 20954
rect 13206 20882 13252 20920
rect 13206 20848 13212 20882
rect 13246 20848 13252 20882
rect 13206 20810 13252 20848
rect 13206 20776 13212 20810
rect 13246 20776 13252 20810
rect 13206 20738 13252 20776
rect 13206 20704 13212 20738
rect 13246 20704 13252 20738
rect 13206 20666 13252 20704
rect 13206 20632 13212 20666
rect 13246 20632 13252 20666
rect 13206 20594 13252 20632
rect 13206 20560 13212 20594
rect 13246 20560 13252 20594
rect 13206 20522 13252 20560
rect 13206 20488 13212 20522
rect 13246 20488 13252 20522
rect 13206 20450 13252 20488
rect 13206 20416 13212 20450
rect 13246 20416 13252 20450
rect 13206 20378 13252 20416
rect 13206 20344 13212 20378
rect 13246 20344 13252 20378
rect 13206 20306 13252 20344
rect 13206 20272 13212 20306
rect 13246 20272 13252 20306
rect 13206 20234 13252 20272
rect 13206 20200 13212 20234
rect 13246 20200 13252 20234
rect 13206 20162 13252 20200
rect 13206 20128 13212 20162
rect 13246 20128 13252 20162
rect 13206 20090 13252 20128
rect 13206 20056 13212 20090
rect 13246 20056 13252 20090
rect 13206 20018 13252 20056
rect 13206 19984 13212 20018
rect 13246 19984 13252 20018
rect 13206 19946 13252 19984
rect 13206 19912 13212 19946
rect 13246 19912 13252 19946
rect 13206 19874 13252 19912
rect 13206 19840 13212 19874
rect 13246 19840 13252 19874
rect 13206 19802 13252 19840
rect 13206 19768 13212 19802
rect 13246 19768 13252 19802
rect 13206 19730 13252 19768
rect 13206 19696 13212 19730
rect 13246 19696 13252 19730
rect 13206 19658 13252 19696
rect 13206 19624 13212 19658
rect 13246 19624 13252 19658
rect 13206 19586 13252 19624
rect 13206 19552 13212 19586
rect 13246 19552 13252 19586
rect 13206 19514 13252 19552
rect 13206 19480 13212 19514
rect 13246 19480 13252 19514
rect 13206 19442 13252 19480
rect 13206 19408 13212 19442
rect 13246 19408 13252 19442
rect 13206 19370 13252 19408
rect 13206 19336 13212 19370
rect 13246 19336 13252 19370
rect 13206 19298 13252 19336
rect 13206 19264 13212 19298
rect 13246 19264 13252 19298
rect 13206 19226 13252 19264
rect 13206 19192 13212 19226
rect 13246 19192 13252 19226
rect 13206 19154 13252 19192
rect 13206 19120 13212 19154
rect 13246 19120 13252 19154
rect 13206 19082 13252 19120
rect 13206 19048 13212 19082
rect 13246 19048 13252 19082
rect 13206 19010 13252 19048
rect 13206 18976 13212 19010
rect 13246 18976 13252 19010
rect 13206 18938 13252 18976
rect 13206 18904 13212 18938
rect 13246 18904 13252 18938
rect 13206 18866 13252 18904
rect 13206 18832 13212 18866
rect 13246 18832 13252 18866
rect 13206 18794 13252 18832
rect 13206 18760 13212 18794
rect 13246 18760 13252 18794
rect 13206 18722 13252 18760
rect 13206 18688 13212 18722
rect 13246 18688 13252 18722
rect 13206 18650 13252 18688
rect 13206 18616 13212 18650
rect 13246 18616 13252 18650
rect 13206 18578 13252 18616
rect 13206 18544 13212 18578
rect 13246 18544 13252 18578
rect 13206 18506 13252 18544
rect 13206 18472 13212 18506
rect 13246 18472 13252 18506
rect 13206 18434 13252 18472
rect 13206 18400 13212 18434
rect 13246 18400 13252 18434
rect 13206 18362 13252 18400
rect 13206 18328 13212 18362
rect 13246 18328 13252 18362
rect 13206 18290 13252 18328
rect 13206 18256 13212 18290
rect 13246 18256 13252 18290
rect 13206 18218 13252 18256
rect 13206 18184 13212 18218
rect 13246 18184 13252 18218
rect 13206 18146 13252 18184
rect 13206 18112 13212 18146
rect 13246 18112 13252 18146
rect 13206 18074 13252 18112
rect 13206 18040 13212 18074
rect 13246 18040 13252 18074
rect 13206 18002 13252 18040
rect 13206 17968 13212 18002
rect 13246 17968 13252 18002
rect 13206 17930 13252 17968
rect 13206 17896 13212 17930
rect 13246 17896 13252 17930
rect 13206 17858 13252 17896
rect 13206 17824 13212 17858
rect 13246 17824 13252 17858
rect 13206 17786 13252 17824
rect 13206 17752 13212 17786
rect 13246 17752 13252 17786
rect 13206 17714 13252 17752
rect 13206 17680 13212 17714
rect 13246 17680 13252 17714
rect 13206 17642 13252 17680
rect 13206 17608 13212 17642
rect 13246 17608 13252 17642
rect 13206 17570 13252 17608
rect 13206 17536 13212 17570
rect 13246 17536 13252 17570
rect 13206 17498 13252 17536
rect 13206 17464 13212 17498
rect 13246 17464 13252 17498
rect 13206 17426 13252 17464
rect 13206 17392 13212 17426
rect 13246 17392 13252 17426
rect 13206 17354 13252 17392
rect 13206 17320 13212 17354
rect 13246 17320 13252 17354
rect 13206 17282 13252 17320
rect 13206 17248 13212 17282
rect 13246 17248 13252 17282
rect 13206 17210 13252 17248
rect 13206 17176 13212 17210
rect 13246 17176 13252 17210
rect 13206 17138 13252 17176
rect 13206 17104 13212 17138
rect 13246 17104 13252 17138
rect 13206 17066 13252 17104
rect 13206 17032 13212 17066
rect 13246 17032 13252 17066
rect 13206 16994 13252 17032
rect 13206 16960 13212 16994
rect 13246 16960 13252 16994
rect 13206 16922 13252 16960
rect 13206 16888 13212 16922
rect 13246 16888 13252 16922
rect 13206 16850 13252 16888
rect 13206 16816 13212 16850
rect 13246 16816 13252 16850
rect 13206 16778 13252 16816
rect 13206 16744 13212 16778
rect 13246 16744 13252 16778
rect 13206 16706 13252 16744
rect 13206 16672 13212 16706
rect 13246 16672 13252 16706
rect 13206 16634 13252 16672
rect 13206 16600 13212 16634
rect 13246 16600 13252 16634
rect 13206 16562 13252 16600
rect 13206 16528 13212 16562
rect 13246 16528 13252 16562
rect 13206 16490 13252 16528
rect 13206 16456 13212 16490
rect 13246 16456 13252 16490
rect 13206 16418 13252 16456
rect 13206 16384 13212 16418
rect 13246 16384 13252 16418
rect 13206 16346 13252 16384
rect 13206 16312 13212 16346
rect 13246 16312 13252 16346
rect 13206 16274 13252 16312
rect 13206 16240 13212 16274
rect 13246 16240 13252 16274
rect 13206 16202 13252 16240
rect 13206 16168 13212 16202
rect 13246 16168 13252 16202
rect 13206 16130 13252 16168
rect 13206 16096 13212 16130
rect 13246 16096 13252 16130
rect 13206 16058 13252 16096
rect 13206 16024 13212 16058
rect 13246 16024 13252 16058
rect 13206 15986 13252 16024
rect 13206 15952 13212 15986
rect 13246 15952 13252 15986
rect 13206 15914 13252 15952
rect 13206 15880 13212 15914
rect 13246 15880 13252 15914
rect 13206 15842 13252 15880
rect 13206 15808 13212 15842
rect 13246 15808 13252 15842
rect 13206 15770 13252 15808
rect 13206 15736 13212 15770
rect 13246 15736 13252 15770
rect 13206 15698 13252 15736
rect 13206 15664 13212 15698
rect 13246 15664 13252 15698
rect 13206 15626 13252 15664
rect 13206 15592 13212 15626
rect 13246 15592 13252 15626
rect 13206 15554 13252 15592
rect 13206 15520 13212 15554
rect 13246 15520 13252 15554
rect 13206 15482 13252 15520
rect 13206 15448 13212 15482
rect 13246 15448 13252 15482
rect 13206 15410 13252 15448
rect 13206 15376 13212 15410
rect 13246 15376 13252 15410
rect 13206 15338 13252 15376
rect 13206 15304 13212 15338
rect 13246 15304 13252 15338
rect 13206 15266 13252 15304
rect 13206 15232 13212 15266
rect 13246 15232 13252 15266
rect 13206 15194 13252 15232
rect 13206 15160 13212 15194
rect 13246 15160 13252 15194
rect 13206 15122 13252 15160
rect 13206 15088 13212 15122
rect 13246 15088 13252 15122
rect 13206 15050 13252 15088
rect 13206 15016 13212 15050
rect 13246 15016 13252 15050
rect 13206 14978 13252 15016
rect 13206 14944 13212 14978
rect 13246 14944 13252 14978
rect 13206 14906 13252 14944
rect 13206 14872 13212 14906
rect 13246 14872 13252 14906
rect 13206 14834 13252 14872
rect 13206 14800 13212 14834
rect 13246 14800 13252 14834
rect 13206 14762 13252 14800
rect 13206 14728 13212 14762
rect 13246 14728 13252 14762
rect 13206 14690 13252 14728
rect 13206 14656 13212 14690
rect 13246 14656 13252 14690
rect 13206 14618 13252 14656
rect 13206 14584 13212 14618
rect 13246 14584 13252 14618
rect 13206 14546 13252 14584
rect 13206 14512 13212 14546
rect 13246 14512 13252 14546
rect 13206 14474 13252 14512
rect 13206 14440 13212 14474
rect 13246 14440 13252 14474
rect 13206 14402 13252 14440
rect 13206 14368 13212 14402
rect 13246 14368 13252 14402
rect 13206 14330 13252 14368
rect 13206 14296 13212 14330
rect 13246 14296 13252 14330
rect 13206 14258 13252 14296
rect 13206 14224 13212 14258
rect 13246 14224 13252 14258
rect 13206 14186 13252 14224
rect 13206 14152 13212 14186
rect 13246 14152 13252 14186
rect 13206 14114 13252 14152
rect 13206 14080 13212 14114
rect 13246 14080 13252 14114
rect 13206 14042 13252 14080
rect 13206 14008 13212 14042
rect 13246 14008 13252 14042
rect 13206 13970 13252 14008
rect 13206 13936 13212 13970
rect 13246 13936 13252 13970
rect 13206 13898 13252 13936
rect 13206 13864 13212 13898
rect 13246 13864 13252 13898
rect 13206 13826 13252 13864
rect 13206 13792 13212 13826
rect 13246 13792 13252 13826
rect 13206 13754 13252 13792
rect 13206 13720 13212 13754
rect 13246 13720 13252 13754
rect 13206 13682 13252 13720
rect 13206 13648 13212 13682
rect 13246 13648 13252 13682
rect 13206 13610 13252 13648
rect 13206 13576 13212 13610
rect 13246 13576 13252 13610
rect 13206 13538 13252 13576
rect 13206 13504 13212 13538
rect 13246 13504 13252 13538
rect 13206 13466 13252 13504
rect 13206 13432 13212 13466
rect 13246 13432 13252 13466
rect 13206 13394 13252 13432
rect 13206 13360 13212 13394
rect 13246 13360 13252 13394
rect 13206 13322 13252 13360
rect 13206 13288 13212 13322
rect 13246 13288 13252 13322
rect 13206 13250 13252 13288
rect 13206 13216 13212 13250
rect 13246 13216 13252 13250
rect 13206 13178 13252 13216
rect 13206 13144 13212 13178
rect 13246 13144 13252 13178
rect 13206 13106 13252 13144
rect 13206 13072 13212 13106
rect 13246 13072 13252 13106
rect 13206 13034 13252 13072
rect 13206 13000 13212 13034
rect 13246 13000 13252 13034
rect 13206 12962 13252 13000
rect 13206 12928 13212 12962
rect 13246 12928 13252 12962
rect 13206 12890 13252 12928
rect 13206 12856 13212 12890
rect 13246 12856 13252 12890
rect 13206 12818 13252 12856
rect 13206 12784 13212 12818
rect 13246 12784 13252 12818
rect 13206 12746 13252 12784
rect 13206 12712 13212 12746
rect 13246 12712 13252 12746
rect 13206 12674 13252 12712
rect 13206 12640 13212 12674
rect 13246 12640 13252 12674
rect 13206 12602 13252 12640
rect 13206 12568 13212 12602
rect 13246 12568 13252 12602
rect 13206 12530 13252 12568
rect 13206 12496 13212 12530
rect 13246 12496 13252 12530
rect 13206 12458 13252 12496
rect 13206 12424 13212 12458
rect 13246 12424 13252 12458
rect 13206 12386 13252 12424
rect 13206 12352 13212 12386
rect 13246 12352 13252 12386
rect 13206 12314 13252 12352
rect 13206 12280 13212 12314
rect 13246 12280 13252 12314
rect 13206 12242 13252 12280
rect 13206 12208 13212 12242
rect 13246 12208 13252 12242
rect 13206 12170 13252 12208
rect 13206 12136 13212 12170
rect 13246 12136 13252 12170
rect 13206 12098 13252 12136
rect 13206 12064 13212 12098
rect 13246 12064 13252 12098
rect 13206 12026 13252 12064
rect 13206 11992 13212 12026
rect 13246 11992 13252 12026
rect 13206 11954 13252 11992
rect 13206 11920 13212 11954
rect 13246 11920 13252 11954
rect 13206 11882 13252 11920
rect 13206 11848 13212 11882
rect 13246 11848 13252 11882
rect 13206 11810 13252 11848
rect 13206 11776 13212 11810
rect 13246 11776 13252 11810
rect 13206 11738 13252 11776
rect 13206 11704 13212 11738
rect 13246 11704 13252 11738
rect 13206 11666 13252 11704
rect 13206 11632 13212 11666
rect 13246 11632 13252 11666
rect 13206 11594 13252 11632
rect 13206 11560 13212 11594
rect 13246 11560 13252 11594
rect 13206 11522 13252 11560
rect 13206 11488 13212 11522
rect 13246 11488 13252 11522
rect 13206 11450 13252 11488
rect 13206 11416 13212 11450
rect 13246 11416 13252 11450
rect 13206 11378 13252 11416
rect 13206 11344 13212 11378
rect 13246 11344 13252 11378
rect 13206 11306 13252 11344
rect 13206 11272 13212 11306
rect 13246 11272 13252 11306
rect 13206 11234 13252 11272
rect 13206 11200 13212 11234
rect 13246 11200 13252 11234
rect 13206 11162 13252 11200
rect 13206 11128 13212 11162
rect 13246 11128 13252 11162
rect 13206 11090 13252 11128
rect 13206 11056 13212 11090
rect 13246 11056 13252 11090
rect 13206 11018 13252 11056
rect 13206 10984 13212 11018
rect 13246 10984 13252 11018
rect 13206 10946 13252 10984
rect 13206 10912 13212 10946
rect 13246 10912 13252 10946
rect 13206 10874 13252 10912
rect 13206 10840 13212 10874
rect 13246 10840 13252 10874
rect 13206 10802 13252 10840
rect 13206 10768 13212 10802
rect 13246 10768 13252 10802
rect 13206 10730 13252 10768
rect 13206 10696 13212 10730
rect 13246 10696 13252 10730
rect 13206 10658 13252 10696
rect 13206 10624 13212 10658
rect 13246 10624 13252 10658
rect 13206 10586 13252 10624
rect 13206 10552 13212 10586
rect 13246 10552 13252 10586
rect 13206 10514 13252 10552
rect 13206 10480 13212 10514
rect 13246 10480 13252 10514
rect 13206 10442 13252 10480
rect 13206 10408 13212 10442
rect 13246 10408 13252 10442
rect 13206 10370 13252 10408
rect 13206 10336 13212 10370
rect 13246 10336 13252 10370
rect 13206 10298 13252 10336
rect 13206 10264 13212 10298
rect 13246 10264 13252 10298
rect 13206 10226 13252 10264
rect 13206 10192 13212 10226
rect 13246 10192 13252 10226
rect 13206 10154 13252 10192
rect 13206 10120 13212 10154
rect 13246 10120 13252 10154
rect 13206 10082 13252 10120
rect 13206 10048 13212 10082
rect 13246 10048 13252 10082
rect 13206 10010 13252 10048
rect 13206 9976 13212 10010
rect 13246 9976 13252 10010
rect 13206 9938 13252 9976
rect 13206 9904 13212 9938
rect 13246 9904 13252 9938
rect 13206 9866 13252 9904
rect 13206 9832 13212 9866
rect 13246 9832 13252 9866
rect 13206 9794 13252 9832
rect 13206 9760 13212 9794
rect 13246 9760 13252 9794
rect 13206 9722 13252 9760
rect 13206 9688 13212 9722
rect 13246 9688 13252 9722
rect 13206 9650 13252 9688
rect 13206 9616 13212 9650
rect 13246 9616 13252 9650
rect 13206 9578 13252 9616
rect 13206 9544 13212 9578
rect 13246 9544 13252 9578
rect 13206 9506 13252 9544
rect 13206 9472 13212 9506
rect 13246 9472 13252 9506
rect 13206 9434 13252 9472
rect 13206 9400 13212 9434
rect 13246 9400 13252 9434
rect 13206 9362 13252 9400
rect 13206 9328 13212 9362
rect 13246 9328 13252 9362
rect 13206 9290 13252 9328
rect 13206 9256 13212 9290
rect 13246 9256 13252 9290
rect 13206 9218 13252 9256
rect 13206 9184 13212 9218
rect 13246 9184 13252 9218
rect 13206 9146 13252 9184
rect 13206 9112 13212 9146
rect 13246 9112 13252 9146
rect 13206 9074 13252 9112
rect 13206 9040 13212 9074
rect 13246 9040 13252 9074
rect 13206 9002 13252 9040
rect 13206 8968 13212 9002
rect 13246 8968 13252 9002
rect 13206 8930 13252 8968
rect 13206 8896 13212 8930
rect 13246 8896 13252 8930
rect 13206 8858 13252 8896
rect 13206 8824 13212 8858
rect 13246 8824 13252 8858
rect 13206 8786 13252 8824
rect 13206 8752 13212 8786
rect 13246 8752 13252 8786
rect 13206 8714 13252 8752
rect 13206 8680 13212 8714
rect 13246 8680 13252 8714
rect 13206 8642 13252 8680
rect 13206 8608 13212 8642
rect 13246 8608 13252 8642
rect 13206 8570 13252 8608
rect 13206 8536 13212 8570
rect 13246 8536 13252 8570
rect 13206 8498 13252 8536
rect 13206 8464 13212 8498
rect 13246 8464 13252 8498
rect 13206 8426 13252 8464
rect 13206 8392 13212 8426
rect 13246 8392 13252 8426
rect 13206 8354 13252 8392
rect 13206 8320 13212 8354
rect 13246 8320 13252 8354
rect 13206 8282 13252 8320
rect 13206 8248 13212 8282
rect 13246 8248 13252 8282
rect 13206 8210 13252 8248
rect 13206 8176 13212 8210
rect 13246 8176 13252 8210
rect 13206 8138 13252 8176
rect 13206 8104 13212 8138
rect 13246 8104 13252 8138
rect 13206 8066 13252 8104
rect 13206 8032 13212 8066
rect 13246 8032 13252 8066
rect 13206 7994 13252 8032
rect 13206 7960 13212 7994
rect 13246 7960 13252 7994
rect 13206 7922 13252 7960
rect 13206 7888 13212 7922
rect 13246 7888 13252 7922
rect 13206 7850 13252 7888
rect 13206 7816 13212 7850
rect 13246 7816 13252 7850
rect 13206 7778 13252 7816
rect 13206 7744 13212 7778
rect 13246 7744 13252 7778
rect 13206 7706 13252 7744
rect 13206 7672 13212 7706
rect 13246 7672 13252 7706
rect 13206 7634 13252 7672
rect 13206 7600 13212 7634
rect 13246 7600 13252 7634
rect 13206 7562 13252 7600
rect 13206 7528 13212 7562
rect 13246 7528 13252 7562
rect 13206 7490 13252 7528
rect 13206 7456 13212 7490
rect 13246 7456 13252 7490
rect 13206 7418 13252 7456
rect 13206 7384 13212 7418
rect 13246 7384 13252 7418
rect 13206 7346 13252 7384
rect 13206 7312 13212 7346
rect 13246 7312 13252 7346
rect 13206 7274 13252 7312
rect 13206 7240 13212 7274
rect 13246 7240 13252 7274
rect 13206 7202 13252 7240
rect 13206 7168 13212 7202
rect 13246 7168 13252 7202
rect 13206 7130 13252 7168
rect 13206 7096 13212 7130
rect 13246 7096 13252 7130
rect 13206 7058 13252 7096
rect 13206 7024 13212 7058
rect 13246 7024 13252 7058
rect 13206 6986 13252 7024
rect 13206 6952 13212 6986
rect 13246 6952 13252 6986
rect 13206 6914 13252 6952
rect 13206 6880 13212 6914
rect 13246 6880 13252 6914
rect 13206 6842 13252 6880
rect 13206 6808 13212 6842
rect 13246 6808 13252 6842
rect 13206 6770 13252 6808
rect 13206 6736 13212 6770
rect 13246 6736 13252 6770
rect 13206 6698 13252 6736
rect 13206 6664 13212 6698
rect 13246 6664 13252 6698
rect 13206 6626 13252 6664
rect 13206 6592 13212 6626
rect 13246 6592 13252 6626
rect 13206 6554 13252 6592
rect 13206 6520 13212 6554
rect 13246 6520 13252 6554
rect 13206 6482 13252 6520
rect 13206 6448 13212 6482
rect 13246 6448 13252 6482
rect 13206 6410 13252 6448
rect 13206 6376 13212 6410
rect 13246 6376 13252 6410
rect 13206 6338 13252 6376
rect 13206 6304 13212 6338
rect 13246 6304 13252 6338
rect 13206 6266 13252 6304
rect 13206 6232 13212 6266
rect 13246 6232 13252 6266
rect 13206 6194 13252 6232
rect 13206 6160 13212 6194
rect 13246 6160 13252 6194
rect 13206 6122 13252 6160
rect 13206 6088 13212 6122
rect 13246 6088 13252 6122
rect 13206 6050 13252 6088
rect 13206 6016 13212 6050
rect 13246 6016 13252 6050
rect 13206 5978 13252 6016
rect 13206 5944 13212 5978
rect 13246 5944 13252 5978
rect 13206 5906 13252 5944
rect 13206 5872 13212 5906
rect 13246 5872 13252 5906
rect 13206 5834 13252 5872
rect 13206 5800 13212 5834
rect 13246 5800 13252 5834
rect 13206 5762 13252 5800
rect 13206 5728 13212 5762
rect 13246 5728 13252 5762
rect 13206 5690 13252 5728
rect 13206 5656 13212 5690
rect 13246 5656 13252 5690
rect 13206 5618 13252 5656
rect 13206 5584 13212 5618
rect 13246 5584 13252 5618
rect 13206 5546 13252 5584
rect 13206 5512 13212 5546
rect 13246 5512 13252 5546
rect 13206 5474 13252 5512
rect 13206 5440 13212 5474
rect 13246 5440 13252 5474
rect 13206 5402 13252 5440
rect 13206 5368 13212 5402
rect 13246 5368 13252 5402
rect 13206 5330 13252 5368
rect 13206 5296 13212 5330
rect 13246 5296 13252 5330
rect 13206 5258 13252 5296
rect 13206 5224 13212 5258
rect 13246 5224 13252 5258
rect 13206 5186 13252 5224
rect 13206 5152 13212 5186
rect 13246 5152 13252 5186
rect 13206 5114 13252 5152
rect 13206 5080 13212 5114
rect 13246 5080 13252 5114
rect 13206 5042 13252 5080
rect 13206 5008 13212 5042
rect 13246 5008 13252 5042
rect 13206 4970 13252 5008
rect 13206 4936 13212 4970
rect 13246 4936 13252 4970
rect 13206 4898 13252 4936
rect 13206 4864 13212 4898
rect 13246 4864 13252 4898
rect 13206 4826 13252 4864
rect 13206 4792 13212 4826
rect 13246 4792 13252 4826
rect 13206 4754 13252 4792
rect 13206 4720 13212 4754
rect 13246 4720 13252 4754
rect 13206 4682 13252 4720
rect 13206 4648 13212 4682
rect 13246 4648 13252 4682
rect 13206 4610 13252 4648
rect 13206 4576 13212 4610
rect 13246 4576 13252 4610
rect 13206 4538 13252 4576
rect 13206 4504 13212 4538
rect 13246 4504 13252 4538
rect 13206 4466 13252 4504
rect 13206 4432 13212 4466
rect 13246 4432 13252 4466
rect 13206 4394 13252 4432
rect 13206 4360 13212 4394
rect 13246 4360 13252 4394
rect 13206 4322 13252 4360
rect 13206 4288 13212 4322
rect 13246 4288 13252 4322
rect 13206 4250 13252 4288
rect 13206 4216 13212 4250
rect 13246 4216 13252 4250
rect 13206 4178 13252 4216
rect 13206 4144 13212 4178
rect 13246 4144 13252 4178
rect 13206 4106 13252 4144
rect 13206 4072 13212 4106
rect 13246 4072 13252 4106
rect 13206 4034 13252 4072
rect 13206 4000 13212 4034
rect 13246 4000 13252 4034
rect 13206 3962 13252 4000
rect 13206 3928 13212 3962
rect 13246 3928 13252 3962
rect 13206 3890 13252 3928
rect 13206 3856 13212 3890
rect 13246 3856 13252 3890
rect 13206 3818 13252 3856
rect 13206 3784 13212 3818
rect 13246 3784 13252 3818
rect 13206 3746 13252 3784
rect 13206 3712 13212 3746
rect 13246 3712 13252 3746
rect 13206 3674 13252 3712
rect 13206 3640 13212 3674
rect 13246 3640 13252 3674
rect 13206 3602 13252 3640
rect 13206 3568 13212 3602
rect 13246 3568 13252 3602
rect 13206 3530 13252 3568
rect 11418 3428 11464 3466
rect 11418 3394 11424 3428
rect 11458 3394 11464 3428
rect 10220 3322 10226 3356
rect 10260 3322 10266 3356
rect 10220 3284 10266 3322
tri 9128 3250 9130 3252 sw
tri 10218 3250 10220 3252 se
rect 10220 3250 10226 3284
rect 10260 3250 10266 3284
rect 11418 3356 11464 3394
rect 11418 3322 11424 3356
rect 11458 3322 11464 3356
rect 11418 3284 11464 3322
tri 10266 3250 10268 3252 sw
tri 11416 3250 11418 3252 se
rect 11418 3250 11424 3284
rect 11458 3250 11464 3284
rect 9082 3242 9130 3250
tri 9130 3242 9138 3250 sw
tri 10210 3242 10218 3250 se
rect 10218 3242 10268 3250
tri 10268 3242 10276 3250 sw
tri 11408 3242 11416 3250 se
rect 11416 3242 11464 3250
rect 9082 3218 9138 3242
tri 9138 3218 9162 3242 sw
tri 10186 3218 10210 3242 se
rect 10210 3218 10276 3242
tri 10276 3218 10300 3242 sw
tri 11384 3218 11408 3242 se
rect 11408 3218 11464 3242
rect 9082 3212 11464 3218
rect 9082 3178 9160 3212
rect 9194 3178 9234 3212
rect 9268 3178 9307 3212
rect 9341 3178 9380 3212
rect 9414 3178 9453 3212
rect 9487 3178 9526 3212
rect 9560 3178 9599 3212
rect 9633 3178 9672 3212
rect 9706 3178 9745 3212
rect 9779 3178 9818 3212
rect 9852 3178 9891 3212
rect 9925 3178 9964 3212
rect 9998 3178 10037 3212
rect 10071 3178 10110 3212
rect 10144 3178 10183 3212
rect 10217 3178 10256 3212
rect 10290 3178 10329 3212
rect 10363 3178 10402 3212
rect 10436 3178 10475 3212
rect 10509 3178 10548 3212
rect 10582 3178 10621 3212
rect 10655 3178 10694 3212
rect 10728 3178 10767 3212
rect 10801 3178 10840 3212
rect 10874 3178 10913 3212
rect 10947 3178 10986 3212
rect 11020 3178 11059 3212
rect 11093 3178 11132 3212
rect 11166 3178 11205 3212
rect 11239 3178 11278 3212
rect 11312 3178 11351 3212
rect 11385 3178 11464 3212
rect 9082 3172 11464 3178
tri 11384 3170 11386 3172 ne
rect 11386 3170 11464 3172
tri 11386 3140 11416 3170 ne
rect 11416 3140 11464 3170
tri 11416 3138 11418 3140 ne
rect -135 3076 -129 3128
rect -77 3076 -65 3128
rect -13 3076 5366 3128
tri 5238 3067 5247 3076 ne
rect 5247 3067 5366 3076
tri 5247 3048 5266 3067 ne
rect 5178 2549 5224 2561
rect 5178 2515 5184 2549
rect 5218 2515 5224 2549
rect 5178 2476 5224 2515
rect 5178 2442 5184 2476
rect 5218 2442 5224 2476
rect 5178 2403 5224 2442
rect 5178 2369 5184 2403
rect 5218 2369 5224 2403
rect 5178 2330 5224 2369
rect 5178 2296 5184 2330
rect 5218 2296 5224 2330
rect 5178 2257 5224 2296
rect 5178 2223 5184 2257
rect 5218 2223 5224 2257
rect 5178 2184 5224 2223
rect 5178 2150 5184 2184
rect 5218 2150 5224 2184
rect 5178 2111 5224 2150
rect 5178 2077 5184 2111
rect 5218 2077 5224 2111
rect 5178 2038 5224 2077
rect 5178 2004 5184 2038
rect 5218 2004 5224 2038
rect 5178 1965 5224 2004
rect 5178 1931 5184 1965
rect 5218 1931 5224 1965
rect 5178 1892 5224 1931
rect 5178 1858 5184 1892
rect 5218 1858 5224 1892
rect 5178 1819 5224 1858
rect 5178 1785 5184 1819
rect 5218 1785 5224 1819
rect 5178 1746 5224 1785
rect 5178 1712 5184 1746
rect 5218 1712 5224 1746
rect 5178 1673 5224 1712
rect 5178 1639 5184 1673
rect 5218 1639 5224 1673
rect 5178 1600 5224 1639
rect 5178 1566 5184 1600
rect 5218 1566 5224 1600
rect 5178 1527 5224 1566
rect 5178 1493 5184 1527
rect 5218 1493 5224 1527
rect 5178 1454 5224 1493
rect 5178 1420 5184 1454
rect 5218 1420 5224 1454
rect 5178 1381 5224 1420
rect 5178 1347 5184 1381
rect 5218 1347 5224 1381
rect 5178 1308 5224 1347
rect 5178 1274 5184 1308
rect 5218 1274 5224 1308
rect 5178 1236 5224 1274
rect 5178 1202 5184 1236
rect 5218 1202 5224 1236
rect 5178 1164 5224 1202
rect 5178 1130 5184 1164
rect 5218 1130 5224 1164
rect 5266 2449 5366 3067
rect 11418 3106 11424 3140
rect 11458 3106 11464 3140
rect 11418 3067 11464 3106
rect 11418 3033 11424 3067
rect 11458 3033 11464 3067
rect 11418 2994 11464 3033
rect 11418 2960 11424 2994
rect 11458 2960 11464 2994
rect 11418 2921 11464 2960
rect 11418 2887 11424 2921
rect 11458 2887 11464 2921
rect 11418 2848 11464 2887
rect 11418 2814 11424 2848
rect 11458 2814 11464 2848
rect 11418 2775 11464 2814
rect 11418 2741 11424 2775
rect 11458 2741 11464 2775
rect 11418 2702 11464 2741
rect 11418 2668 11424 2702
rect 11458 2668 11464 2702
rect 11418 2629 11464 2668
rect 5406 2595 6041 2601
rect 5406 2561 5418 2595
rect 5452 2561 5500 2595
rect 5534 2561 5583 2595
rect 5617 2561 5666 2595
rect 5700 2561 5749 2595
rect 5783 2561 5832 2595
rect 5866 2589 6041 2595
rect 5866 2561 5940 2589
rect 5406 2555 5940 2561
rect 5974 2555 6041 2589
tri 5807 2522 5840 2555 ne
rect 5840 2522 6041 2555
tri 5840 2521 5841 2522 ne
rect 5841 2515 6041 2522
rect 5841 2481 5940 2515
rect 5974 2481 6041 2515
tri 5366 2449 5396 2479 sw
rect 5266 2445 5396 2449
tri 5396 2445 5400 2449 sw
rect 5266 2439 5801 2445
rect 5266 2405 5278 2439
rect 5312 2405 5357 2439
rect 5391 2405 5436 2439
rect 5470 2405 5515 2439
rect 5549 2405 5595 2439
rect 5629 2405 5675 2439
rect 5709 2405 5755 2439
rect 5789 2405 5801 2439
rect 5266 2399 5801 2405
rect 5841 2441 6041 2481
rect 5841 2407 5940 2441
rect 5974 2407 6041 2441
rect 5266 2376 5377 2399
tri 5377 2376 5400 2399 nw
rect 5266 2367 5368 2376
tri 5368 2367 5377 2376 nw
rect 5841 2367 6041 2407
rect 5266 2157 5366 2367
tri 5366 2365 5368 2367 nw
rect 5841 2333 5940 2367
rect 5974 2333 6041 2367
tri 5821 2303 5841 2323 se
rect 5841 2303 6041 2333
tri 5811 2293 5821 2303 se
rect 5821 2293 6041 2303
tri 5807 2289 5811 2293 se
rect 5811 2289 5940 2293
rect 5406 2283 5940 2289
rect 5406 2249 5418 2283
rect 5452 2249 5500 2283
rect 5534 2249 5583 2283
rect 5617 2249 5666 2283
rect 5700 2249 5749 2283
rect 5783 2249 5832 2283
rect 5866 2259 5940 2283
rect 5974 2259 6041 2293
rect 5866 2249 6041 2259
rect 5406 2243 6041 2249
tri 5807 2230 5820 2243 ne
rect 5820 2230 6041 2243
tri 5820 2219 5831 2230 ne
rect 5831 2219 6041 2230
tri 5831 2209 5841 2219 ne
rect 5841 2185 5940 2219
rect 5974 2185 6041 2219
tri 5366 2157 5376 2167 sw
rect 5266 2145 5376 2157
tri 5376 2145 5388 2157 sw
rect 5841 2145 6041 2185
rect 5266 2133 5388 2145
tri 5388 2133 5400 2145 sw
rect 5266 2127 5801 2133
rect 5266 2093 5278 2127
rect 5312 2093 5357 2127
rect 5391 2093 5436 2127
rect 5470 2093 5515 2127
rect 5549 2093 5595 2127
rect 5629 2093 5675 2127
rect 5709 2093 5755 2127
rect 5789 2093 5801 2127
rect 5266 2087 5801 2093
rect 5841 2111 5940 2145
rect 5974 2111 6041 2145
rect 5266 2084 5397 2087
tri 5397 2084 5400 2087 nw
rect 5266 2071 5384 2084
tri 5384 2071 5397 2084 nw
rect 5841 2071 6041 2111
rect 5266 1849 5366 2071
tri 5366 2053 5384 2071 nw
rect 5841 2037 5940 2071
rect 5974 2037 6041 2071
tri 5827 1997 5841 2011 se
rect 5841 1997 6041 2037
tri 5807 1977 5827 1997 se
rect 5827 1977 5940 1997
rect 5406 1971 5940 1977
rect 5406 1937 5418 1971
rect 5452 1937 5500 1971
rect 5534 1937 5583 1971
rect 5617 1937 5666 1971
rect 5700 1937 5749 1971
rect 5783 1937 5832 1971
rect 5866 1963 5940 1971
rect 5974 1963 6041 1997
rect 5866 1937 6041 1963
rect 5406 1931 6041 1937
tri 5807 1923 5815 1931 ne
rect 5815 1923 6041 1931
tri 5815 1897 5841 1923 ne
rect 5841 1889 5940 1923
rect 5974 1889 6041 1923
tri 5366 1849 5372 1855 sw
rect 5841 1849 6041 1889
rect 5266 1821 5372 1849
tri 5372 1821 5400 1849 sw
rect 5266 1815 5801 1821
rect 5266 1781 5278 1815
rect 5312 1781 5357 1815
rect 5391 1781 5436 1815
rect 5470 1781 5515 1815
rect 5549 1781 5595 1815
rect 5629 1781 5675 1815
rect 5709 1781 5755 1815
rect 5789 1781 5801 1815
rect 5266 1775 5801 1781
rect 5841 1815 5940 1849
rect 5974 1815 6041 1849
rect 5841 1775 6041 1815
rect 5266 1519 5366 1775
tri 5366 1741 5400 1775 nw
rect 5841 1741 5940 1775
rect 5974 1741 6041 1775
rect 5841 1701 6041 1741
tri 5809 1667 5841 1699 se
rect 5841 1667 5940 1701
rect 5974 1667 6041 1701
tri 5807 1665 5809 1667 se
rect 5809 1665 6041 1667
rect 5406 1659 6041 1665
rect 5406 1625 5418 1659
rect 5452 1625 5500 1659
rect 5534 1625 5583 1659
rect 5617 1625 5666 1659
rect 5700 1625 5749 1659
rect 5783 1625 5832 1659
rect 5866 1627 6041 1659
rect 5866 1625 5940 1627
rect 5406 1619 5940 1625
tri 5807 1593 5833 1619 ne
rect 5833 1593 5940 1619
rect 5974 1593 6041 1627
tri 5833 1585 5841 1593 ne
rect 5841 1553 6041 1593
tri 5366 1519 5390 1543 sw
rect 5841 1519 5940 1553
rect 5974 1519 6041 1553
rect 5266 1509 5390 1519
tri 5390 1509 5400 1519 sw
rect 5266 1503 5801 1509
rect 5266 1469 5278 1503
rect 5312 1469 5357 1503
rect 5391 1469 5436 1503
rect 5470 1469 5515 1503
rect 5549 1469 5595 1503
rect 5629 1469 5675 1503
rect 5709 1469 5755 1503
rect 5789 1469 5801 1503
rect 5266 1463 5801 1469
rect 5841 1479 6041 1519
rect 5266 1445 5382 1463
tri 5382 1445 5400 1463 nw
rect 5841 1445 5940 1479
rect 5974 1445 6041 1479
rect 5266 1226 5366 1445
tri 5366 1429 5382 1445 nw
rect 5841 1406 6041 1445
tri 5826 1372 5841 1387 se
rect 5841 1372 5940 1406
rect 5974 1372 6041 1406
tri 5808 1354 5826 1372 se
rect 5826 1354 6041 1372
tri 5807 1353 5808 1354 se
rect 5808 1353 6041 1354
rect 5406 1347 6041 1353
rect 5406 1313 5418 1347
rect 5452 1313 5500 1347
rect 5534 1313 5583 1347
rect 5617 1313 5666 1347
rect 5700 1313 5749 1347
rect 5783 1313 5832 1347
rect 5866 1333 6041 1347
rect 5866 1313 5940 1333
rect 5406 1307 5940 1313
tri 5807 1299 5815 1307 ne
rect 5815 1299 5940 1307
rect 5974 1299 6041 1333
tri 5815 1281 5833 1299 ne
rect 5833 1281 6041 1299
tri 5833 1273 5841 1281 ne
rect 5841 1260 6041 1281
tri 5366 1226 5371 1231 sw
rect 5841 1226 5940 1260
rect 5974 1226 6041 1260
rect 5266 1208 5371 1226
tri 5371 1208 5389 1226 sw
rect 5266 1197 5389 1208
tri 5389 1197 5400 1208 sw
rect 5266 1191 5801 1197
rect 5266 1157 5278 1191
rect 5312 1157 5357 1191
rect 5391 1157 5436 1191
rect 5470 1157 5515 1191
rect 5549 1157 5595 1191
rect 5629 1157 5675 1191
rect 5709 1157 5755 1191
rect 5789 1157 5801 1191
rect 5266 1151 5801 1157
rect 5841 1187 6041 1226
rect 5841 1153 5940 1187
rect 5974 1153 6041 1187
rect 5178 1092 5224 1130
rect 5178 1058 5184 1092
rect 5218 1058 5224 1092
rect 5841 1114 6041 1153
rect 5841 1080 5940 1114
rect 5974 1080 6041 1114
tri 5828 1062 5841 1075 se
rect 5841 1062 6041 1080
rect 5178 1046 5224 1058
tri 5814 1048 5828 1062 se
rect 5828 1048 6041 1062
tri 5812 1046 5814 1048 se
rect 5814 1046 6041 1048
tri 5807 1041 5812 1046 se
rect 5812 1041 6041 1046
rect 5406 1035 5940 1041
rect 5406 1001 5418 1035
rect 5452 1001 5500 1035
rect 5534 1001 5583 1035
rect 5617 1001 5666 1035
rect 5700 1001 5749 1035
rect 5783 1001 5832 1035
rect 5866 1007 5940 1035
rect 5974 1007 6041 1041
rect 5866 1001 6041 1007
rect 5406 995 6041 1001
rect 11418 2595 11424 2629
rect 11458 2595 11464 2629
rect 11418 2556 11464 2595
rect 11418 2522 11424 2556
rect 11458 2522 11464 2556
rect 11418 2483 11464 2522
rect 11418 2449 11424 2483
rect 11458 2449 11464 2483
rect 11418 2410 11464 2449
rect 11418 2376 11424 2410
rect 11458 2376 11464 2410
rect 11418 2337 11464 2376
rect 11418 2303 11424 2337
rect 11458 2303 11464 2337
rect 11418 2264 11464 2303
rect 11418 2230 11424 2264
rect 11458 2230 11464 2264
rect 11418 2191 11464 2230
rect 11418 2157 11424 2191
rect 11458 2157 11464 2191
rect 11418 2118 11464 2157
rect 11418 2084 11424 2118
rect 11458 2084 11464 2118
rect 11418 2045 11464 2084
rect 11418 2011 11424 2045
rect 11458 2011 11464 2045
rect 11418 1972 11464 2011
rect 11418 1938 11424 1972
rect 11458 1938 11464 1972
rect 11418 1899 11464 1938
rect 11418 1865 11424 1899
rect 11458 1865 11464 1899
rect 11418 1826 11464 1865
rect 11418 1792 11424 1826
rect 11458 1792 11464 1826
rect 11418 1753 11464 1792
rect 11418 1719 11424 1753
rect 11458 1719 11464 1753
rect 11418 1680 11464 1719
rect 11418 1646 11424 1680
rect 11458 1646 11464 1680
rect 11418 1607 11464 1646
rect 11418 1573 11424 1607
rect 11458 1573 11464 1607
rect 11418 1534 11464 1573
rect 11418 1500 11424 1534
rect 11458 1500 11464 1534
rect 11418 1461 11464 1500
rect 11418 1427 11424 1461
rect 11458 1427 11464 1461
rect 11418 1388 11464 1427
rect 11418 1354 11424 1388
rect 11458 1354 11464 1388
rect 11418 1315 11464 1354
rect 11418 1281 11424 1315
rect 11458 1281 11464 1315
rect 11418 1242 11464 1281
rect 11418 1208 11424 1242
rect 11458 1208 11464 1242
rect 11418 1169 11464 1208
rect 11418 1135 11424 1169
rect 11458 1135 11464 1169
rect 11418 1096 11464 1135
rect 11418 1062 11424 1096
rect 11458 1062 11464 1096
rect 11418 1023 11464 1062
rect 11418 989 11424 1023
rect 11458 989 11464 1023
rect 11418 950 11464 989
rect 11418 916 11424 950
rect 11458 916 11464 950
rect 11418 877 11464 916
rect 11418 843 11424 877
rect 11458 843 11464 877
rect 11418 804 11464 843
rect 11418 770 11424 804
rect 11458 770 11464 804
rect 11418 731 11464 770
rect 11418 697 11424 731
rect 11458 697 11464 731
rect 11418 658 11464 697
rect 11418 624 11424 658
rect 11458 624 11464 658
rect 11418 585 11464 624
rect 11418 551 11424 585
rect 11458 551 11464 585
rect 11418 512 11464 551
rect 11418 478 11424 512
rect 11458 478 11464 512
rect 11418 439 11464 478
rect 11418 405 11424 439
rect 11458 405 11464 439
rect 11418 366 11464 405
rect 11418 332 11424 366
rect 11458 332 11464 366
rect 11418 293 11464 332
rect 11601 3493 11653 3499
rect 11601 3429 11653 3441
rect 11601 417 11653 3377
rect 11601 383 11610 417
rect 11644 383 11653 417
rect 11601 345 11653 383
rect 11601 311 11610 345
rect 11644 311 11653 345
rect 11601 299 11653 311
rect 13206 3496 13212 3530
rect 13246 3496 13252 3530
rect 13206 3458 13252 3496
rect 13206 3424 13212 3458
rect 13246 3424 13252 3458
rect 13206 3386 13252 3424
rect 13206 3352 13212 3386
rect 13246 3352 13252 3386
rect 13206 3314 13252 3352
rect 13206 3280 13212 3314
rect 13246 3280 13252 3314
rect 13206 3242 13252 3280
rect 13206 3208 13212 3242
rect 13246 3208 13252 3242
rect 13206 3170 13252 3208
rect 13206 3136 13212 3170
rect 13246 3136 13252 3170
rect 13206 3098 13252 3136
rect 13206 3064 13212 3098
rect 13246 3064 13252 3098
rect 13206 3026 13252 3064
rect 13206 2992 13212 3026
rect 13246 2992 13252 3026
rect 13206 2954 13252 2992
rect 13206 2920 13212 2954
rect 13246 2920 13252 2954
rect 13206 2882 13252 2920
rect 13206 2848 13212 2882
rect 13246 2848 13252 2882
rect 13206 2810 13252 2848
rect 13206 2776 13212 2810
rect 13246 2776 13252 2810
rect 13206 2738 13252 2776
rect 13206 2704 13212 2738
rect 13246 2704 13252 2738
rect 13206 2666 13252 2704
rect 13206 2632 13212 2666
rect 13246 2632 13252 2666
rect 13206 2594 13252 2632
rect 13206 2560 13212 2594
rect 13246 2560 13252 2594
rect 13206 2522 13252 2560
rect 13206 2488 13212 2522
rect 13246 2488 13252 2522
rect 13206 2450 13252 2488
rect 13206 2416 13212 2450
rect 13246 2416 13252 2450
rect 13206 2378 13252 2416
rect 13206 2344 13212 2378
rect 13246 2344 13252 2378
rect 13206 2306 13252 2344
rect 13206 2272 13212 2306
rect 13246 2272 13252 2306
rect 13206 2234 13252 2272
rect 13206 2200 13212 2234
rect 13246 2200 13252 2234
rect 13206 2162 13252 2200
rect 13206 2128 13212 2162
rect 13246 2128 13252 2162
rect 13206 2090 13252 2128
rect 13206 2056 13212 2090
rect 13246 2056 13252 2090
rect 13206 2018 13252 2056
rect 13206 1984 13212 2018
rect 13246 1984 13252 2018
rect 13206 1946 13252 1984
rect 13206 1912 13212 1946
rect 13246 1912 13252 1946
rect 13206 1874 13252 1912
rect 13206 1840 13212 1874
rect 13246 1840 13252 1874
rect 13206 1802 13252 1840
rect 13206 1768 13212 1802
rect 13246 1768 13252 1802
rect 13206 1730 13252 1768
rect 13206 1696 13212 1730
rect 13246 1696 13252 1730
rect 13206 1658 13252 1696
rect 13206 1624 13212 1658
rect 13246 1624 13252 1658
rect 13206 1586 13252 1624
rect 13206 1552 13212 1586
rect 13246 1552 13252 1586
rect 13206 1514 13252 1552
rect 13206 1480 13212 1514
rect 13246 1480 13252 1514
rect 13206 1442 13252 1480
rect 13206 1408 13212 1442
rect 13246 1408 13252 1442
rect 13206 1370 13252 1408
rect 13206 1336 13212 1370
rect 13246 1336 13252 1370
rect 13206 1298 13252 1336
rect 13206 1264 13212 1298
rect 13246 1264 13252 1298
rect 13206 1226 13252 1264
rect 13206 1192 13212 1226
rect 13246 1192 13252 1226
rect 13206 1154 13252 1192
rect 13206 1120 13212 1154
rect 13246 1120 13252 1154
rect 13206 1082 13252 1120
rect 13206 1048 13212 1082
rect 13246 1048 13252 1082
rect 13206 1010 13252 1048
rect 13206 976 13212 1010
rect 13246 976 13252 1010
rect 13206 938 13252 976
rect 13206 904 13212 938
rect 13246 904 13252 938
rect 13206 866 13252 904
rect 13206 832 13212 866
rect 13246 832 13252 866
rect 13206 794 13252 832
rect 13206 760 13212 794
rect 13246 760 13252 794
rect 13206 722 13252 760
rect 13206 688 13212 722
rect 13246 688 13252 722
rect 13206 650 13252 688
rect 13206 616 13212 650
rect 13246 616 13252 650
rect 13206 578 13252 616
rect 13206 544 13212 578
rect 13246 544 13252 578
rect 13206 506 13252 544
rect 13206 472 13212 506
rect 13246 472 13252 506
rect 13206 434 13252 472
rect 13206 400 13212 434
rect 13246 400 13252 434
rect 14934 38468 14980 38506
rect 14934 38434 14940 38468
rect 14974 38434 14980 38468
rect 14934 38396 14980 38434
rect 14934 38362 14940 38396
rect 14974 38362 14980 38396
rect 14934 38324 14980 38362
rect 14934 38290 14940 38324
rect 14974 38290 14980 38324
rect 14934 38252 14980 38290
rect 14934 38218 14940 38252
rect 14974 38218 14980 38252
rect 14934 38180 14980 38218
rect 14934 38146 14940 38180
rect 14974 38146 14980 38180
rect 14934 38108 14980 38146
rect 14934 38074 14940 38108
rect 14974 38074 14980 38108
rect 14934 38036 14980 38074
rect 14934 38002 14940 38036
rect 14974 38002 14980 38036
rect 14934 37964 14980 38002
rect 14934 37930 14940 37964
rect 14974 37930 14980 37964
rect 14934 37892 14980 37930
rect 14934 37858 14940 37892
rect 14974 37858 14980 37892
rect 14934 37820 14980 37858
rect 14934 37786 14940 37820
rect 14974 37786 14980 37820
rect 14934 37748 14980 37786
rect 14934 37714 14940 37748
rect 14974 37714 14980 37748
rect 14934 37676 14980 37714
rect 14934 37642 14940 37676
rect 14974 37642 14980 37676
rect 14934 37604 14980 37642
rect 14934 37570 14940 37604
rect 14974 37570 14980 37604
rect 14934 37532 14980 37570
rect 14934 37498 14940 37532
rect 14974 37498 14980 37532
rect 14934 37460 14980 37498
rect 14934 37426 14940 37460
rect 14974 37426 14980 37460
rect 14934 37388 14980 37426
rect 14934 37354 14940 37388
rect 14974 37354 14980 37388
rect 14934 37316 14980 37354
rect 14934 37282 14940 37316
rect 14974 37282 14980 37316
rect 14934 37244 14980 37282
rect 14934 37210 14940 37244
rect 14974 37210 14980 37244
rect 14934 37172 14980 37210
rect 14934 37138 14940 37172
rect 14974 37138 14980 37172
rect 14934 37100 14980 37138
rect 14934 37066 14940 37100
rect 14974 37066 14980 37100
rect 14934 37028 14980 37066
rect 14934 36994 14940 37028
rect 14974 36994 14980 37028
rect 14934 36956 14980 36994
rect 14934 36922 14940 36956
rect 14974 36922 14980 36956
rect 14934 36884 14980 36922
rect 14934 36850 14940 36884
rect 14974 36850 14980 36884
rect 14934 36812 14980 36850
rect 14934 36778 14940 36812
rect 14974 36778 14980 36812
rect 14934 36740 14980 36778
rect 14934 36706 14940 36740
rect 14974 36706 14980 36740
rect 14934 36668 14980 36706
rect 14934 36634 14940 36668
rect 14974 36634 14980 36668
rect 14934 36596 14980 36634
rect 14934 36562 14940 36596
rect 14974 36562 14980 36596
rect 14934 36524 14980 36562
rect 14934 36490 14940 36524
rect 14974 36490 14980 36524
rect 14934 36452 14980 36490
rect 14934 36418 14940 36452
rect 14974 36418 14980 36452
rect 14934 36380 14980 36418
rect 14934 36346 14940 36380
rect 14974 36346 14980 36380
rect 14934 36308 14980 36346
rect 14934 36274 14940 36308
rect 14974 36274 14980 36308
rect 14934 36236 14980 36274
rect 14934 36202 14940 36236
rect 14974 36202 14980 36236
rect 14934 36164 14980 36202
rect 14934 36130 14940 36164
rect 14974 36130 14980 36164
rect 14934 36092 14980 36130
rect 14934 36058 14940 36092
rect 14974 36058 14980 36092
rect 14934 36020 14980 36058
rect 14934 35986 14940 36020
rect 14974 35986 14980 36020
rect 14934 35948 14980 35986
rect 14934 35914 14940 35948
rect 14974 35914 14980 35948
rect 14934 35876 14980 35914
rect 14934 35842 14940 35876
rect 14974 35842 14980 35876
rect 14934 35804 14980 35842
rect 14934 35770 14940 35804
rect 14974 35770 14980 35804
rect 14934 35732 14980 35770
rect 14934 35698 14940 35732
rect 14974 35698 14980 35732
rect 14934 35660 14980 35698
rect 14934 35626 14940 35660
rect 14974 35626 14980 35660
rect 14934 35588 14980 35626
rect 14934 35554 14940 35588
rect 14974 35554 14980 35588
rect 14934 35516 14980 35554
rect 14934 35482 14940 35516
rect 14974 35482 14980 35516
rect 14934 35444 14980 35482
rect 14934 35410 14940 35444
rect 14974 35410 14980 35444
rect 14934 35372 14980 35410
rect 14934 35338 14940 35372
rect 14974 35338 14980 35372
rect 14934 35300 14980 35338
rect 14934 35266 14940 35300
rect 14974 35266 14980 35300
rect 14934 35228 14980 35266
rect 14934 35194 14940 35228
rect 14974 35194 14980 35228
rect 14934 35156 14980 35194
rect 14934 35122 14940 35156
rect 14974 35122 14980 35156
rect 14934 35084 14980 35122
rect 14934 35050 14940 35084
rect 14974 35050 14980 35084
rect 14934 35012 14980 35050
rect 14934 34978 14940 35012
rect 14974 34978 14980 35012
rect 14934 34940 14980 34978
rect 14934 34906 14940 34940
rect 14974 34906 14980 34940
rect 14934 34868 14980 34906
rect 14934 34834 14940 34868
rect 14974 34834 14980 34868
rect 14934 34796 14980 34834
rect 14934 34762 14940 34796
rect 14974 34762 14980 34796
rect 14934 34724 14980 34762
rect 14934 34690 14940 34724
rect 14974 34690 14980 34724
rect 14934 34652 14980 34690
rect 14934 34618 14940 34652
rect 14974 34618 14980 34652
rect 14934 34580 14980 34618
rect 14934 34546 14940 34580
rect 14974 34546 14980 34580
rect 14934 34508 14980 34546
rect 14934 34474 14940 34508
rect 14974 34474 14980 34508
rect 14934 34436 14980 34474
rect 14934 34402 14940 34436
rect 14974 34402 14980 34436
rect 14934 34364 14980 34402
rect 14934 34330 14940 34364
rect 14974 34330 14980 34364
rect 14934 34292 14980 34330
rect 14934 34258 14940 34292
rect 14974 34258 14980 34292
rect 14934 34220 14980 34258
rect 14934 34186 14940 34220
rect 14974 34186 14980 34220
rect 14934 34148 14980 34186
rect 14934 34114 14940 34148
rect 14974 34114 14980 34148
rect 14934 34076 14980 34114
rect 14934 34042 14940 34076
rect 14974 34042 14980 34076
rect 14934 34004 14980 34042
rect 14934 33970 14940 34004
rect 14974 33970 14980 34004
rect 14934 33932 14980 33970
rect 14934 33898 14940 33932
rect 14974 33898 14980 33932
rect 14934 33860 14980 33898
rect 14934 33826 14940 33860
rect 14974 33826 14980 33860
rect 14934 33788 14980 33826
rect 14934 33754 14940 33788
rect 14974 33754 14980 33788
rect 14934 33716 14980 33754
rect 14934 33682 14940 33716
rect 14974 33682 14980 33716
rect 14934 33644 14980 33682
rect 14934 33610 14940 33644
rect 14974 33610 14980 33644
rect 14934 33572 14980 33610
rect 14934 33538 14940 33572
rect 14974 33538 14980 33572
rect 14934 33500 14980 33538
rect 14934 33466 14940 33500
rect 14974 33466 14980 33500
rect 14934 33428 14980 33466
rect 14934 33394 14940 33428
rect 14974 33394 14980 33428
rect 14934 33356 14980 33394
rect 14934 33322 14940 33356
rect 14974 33322 14980 33356
rect 14934 33284 14980 33322
rect 14934 33250 14940 33284
rect 14974 33250 14980 33284
rect 14934 33212 14980 33250
rect 14934 33178 14940 33212
rect 14974 33178 14980 33212
rect 14934 33140 14980 33178
rect 14934 33106 14940 33140
rect 14974 33106 14980 33140
rect 14934 33068 14980 33106
rect 14934 33034 14940 33068
rect 14974 33034 14980 33068
rect 14934 32996 14980 33034
rect 14934 32962 14940 32996
rect 14974 32962 14980 32996
rect 14934 32924 14980 32962
rect 14934 32890 14940 32924
rect 14974 32890 14980 32924
rect 14934 32852 14980 32890
rect 14934 32818 14940 32852
rect 14974 32818 14980 32852
rect 14934 32780 14980 32818
rect 14934 32746 14940 32780
rect 14974 32746 14980 32780
rect 14934 32708 14980 32746
rect 14934 32674 14940 32708
rect 14974 32674 14980 32708
rect 14934 32636 14980 32674
rect 14934 32602 14940 32636
rect 14974 32602 14980 32636
rect 14934 32564 14980 32602
rect 14934 32530 14940 32564
rect 14974 32530 14980 32564
rect 14934 32492 14980 32530
rect 14934 32458 14940 32492
rect 14974 32458 14980 32492
rect 14934 32420 14980 32458
rect 14934 32386 14940 32420
rect 14974 32386 14980 32420
rect 14934 32348 14980 32386
rect 14934 32314 14940 32348
rect 14974 32314 14980 32348
rect 14934 32276 14980 32314
rect 14934 32242 14940 32276
rect 14974 32242 14980 32276
rect 14934 32204 14980 32242
rect 14934 32170 14940 32204
rect 14974 32170 14980 32204
rect 14934 32132 14980 32170
rect 14934 32098 14940 32132
rect 14974 32098 14980 32132
rect 14934 32060 14980 32098
rect 14934 32026 14940 32060
rect 14974 32026 14980 32060
rect 14934 31988 14980 32026
rect 14934 31954 14940 31988
rect 14974 31954 14980 31988
rect 14934 31916 14980 31954
rect 14934 31882 14940 31916
rect 14974 31882 14980 31916
rect 14934 31844 14980 31882
rect 14934 31810 14940 31844
rect 14974 31810 14980 31844
rect 14934 31772 14980 31810
rect 14934 31738 14940 31772
rect 14974 31738 14980 31772
rect 14934 31700 14980 31738
rect 14934 31666 14940 31700
rect 14974 31666 14980 31700
rect 14934 31628 14980 31666
rect 14934 31594 14940 31628
rect 14974 31594 14980 31628
rect 14934 31556 14980 31594
rect 14934 31522 14940 31556
rect 14974 31522 14980 31556
rect 14934 31484 14980 31522
rect 14934 31450 14940 31484
rect 14974 31450 14980 31484
rect 14934 31412 14980 31450
rect 14934 31378 14940 31412
rect 14974 31378 14980 31412
rect 14934 31340 14980 31378
rect 14934 31306 14940 31340
rect 14974 31306 14980 31340
rect 14934 31268 14980 31306
rect 14934 31234 14940 31268
rect 14974 31234 14980 31268
rect 14934 31196 14980 31234
rect 14934 31162 14940 31196
rect 14974 31162 14980 31196
rect 14934 31124 14980 31162
rect 14934 31090 14940 31124
rect 14974 31090 14980 31124
rect 14934 31052 14980 31090
rect 14934 31018 14940 31052
rect 14974 31018 14980 31052
rect 14934 30980 14980 31018
rect 14934 30946 14940 30980
rect 14974 30946 14980 30980
rect 14934 30908 14980 30946
rect 14934 30874 14940 30908
rect 14974 30874 14980 30908
rect 14934 30836 14980 30874
rect 14934 30802 14940 30836
rect 14974 30802 14980 30836
rect 14934 30764 14980 30802
rect 14934 30730 14940 30764
rect 14974 30730 14980 30764
rect 14934 30692 14980 30730
rect 14934 30658 14940 30692
rect 14974 30658 14980 30692
rect 14934 30620 14980 30658
rect 14934 30586 14940 30620
rect 14974 30586 14980 30620
rect 14934 30548 14980 30586
rect 14934 30514 14940 30548
rect 14974 30514 14980 30548
rect 14934 30476 14980 30514
rect 14934 30442 14940 30476
rect 14974 30442 14980 30476
rect 14934 30404 14980 30442
rect 14934 30370 14940 30404
rect 14974 30370 14980 30404
rect 14934 30332 14980 30370
rect 14934 30298 14940 30332
rect 14974 30298 14980 30332
rect 14934 30260 14980 30298
rect 14934 30226 14940 30260
rect 14974 30226 14980 30260
rect 14934 30188 14980 30226
rect 14934 30154 14940 30188
rect 14974 30154 14980 30188
rect 14934 30116 14980 30154
rect 14934 30082 14940 30116
rect 14974 30082 14980 30116
rect 14934 30044 14980 30082
rect 14934 30010 14940 30044
rect 14974 30010 14980 30044
rect 14934 29972 14980 30010
rect 14934 29938 14940 29972
rect 14974 29938 14980 29972
rect 14934 29900 14980 29938
rect 14934 29866 14940 29900
rect 14974 29866 14980 29900
rect 14934 29828 14980 29866
rect 14934 29794 14940 29828
rect 14974 29794 14980 29828
rect 14934 29756 14980 29794
rect 14934 29722 14940 29756
rect 14974 29722 14980 29756
rect 14934 29684 14980 29722
rect 14934 29650 14940 29684
rect 14974 29650 14980 29684
rect 14934 29612 14980 29650
rect 14934 29578 14940 29612
rect 14974 29578 14980 29612
rect 14934 29540 14980 29578
rect 14934 29506 14940 29540
rect 14974 29506 14980 29540
rect 14934 29468 14980 29506
rect 14934 29434 14940 29468
rect 14974 29434 14980 29468
rect 14934 29396 14980 29434
rect 14934 29362 14940 29396
rect 14974 29362 14980 29396
rect 14934 29324 14980 29362
rect 14934 29290 14940 29324
rect 14974 29290 14980 29324
rect 14934 29252 14980 29290
rect 14934 29218 14940 29252
rect 14974 29218 14980 29252
rect 14934 29180 14980 29218
rect 14934 29146 14940 29180
rect 14974 29146 14980 29180
rect 14934 29108 14980 29146
rect 14934 29074 14940 29108
rect 14974 29074 14980 29108
rect 14934 29036 14980 29074
rect 14934 29002 14940 29036
rect 14974 29002 14980 29036
rect 14934 28964 14980 29002
rect 14934 28930 14940 28964
rect 14974 28930 14980 28964
rect 14934 28892 14980 28930
rect 14934 28858 14940 28892
rect 14974 28858 14980 28892
rect 14934 28820 14980 28858
rect 14934 28786 14940 28820
rect 14974 28786 14980 28820
rect 14934 28748 14980 28786
rect 14934 28714 14940 28748
rect 14974 28714 14980 28748
rect 14934 28676 14980 28714
rect 14934 28642 14940 28676
rect 14974 28642 14980 28676
rect 14934 28604 14980 28642
rect 14934 28570 14940 28604
rect 14974 28570 14980 28604
rect 14934 28532 14980 28570
rect 14934 28498 14940 28532
rect 14974 28498 14980 28532
rect 14934 28460 14980 28498
rect 14934 28426 14940 28460
rect 14974 28426 14980 28460
rect 14934 28388 14980 28426
rect 14934 28354 14940 28388
rect 14974 28354 14980 28388
rect 14934 28316 14980 28354
rect 14934 28282 14940 28316
rect 14974 28282 14980 28316
rect 14934 28244 14980 28282
rect 14934 28210 14940 28244
rect 14974 28210 14980 28244
rect 14934 28172 14980 28210
rect 14934 28138 14940 28172
rect 14974 28138 14980 28172
rect 14934 28100 14980 28138
rect 14934 28066 14940 28100
rect 14974 28066 14980 28100
rect 14934 28028 14980 28066
rect 14934 27994 14940 28028
rect 14974 27994 14980 28028
rect 14934 27956 14980 27994
rect 14934 27922 14940 27956
rect 14974 27922 14980 27956
rect 14934 27884 14980 27922
rect 14934 27850 14940 27884
rect 14974 27850 14980 27884
rect 14934 27812 14980 27850
rect 14934 27778 14940 27812
rect 14974 27778 14980 27812
rect 14934 27740 14980 27778
rect 14934 27706 14940 27740
rect 14974 27706 14980 27740
rect 14934 27668 14980 27706
rect 14934 27634 14940 27668
rect 14974 27634 14980 27668
rect 14934 27596 14980 27634
rect 14934 27562 14940 27596
rect 14974 27562 14980 27596
rect 14934 27524 14980 27562
rect 14934 27490 14940 27524
rect 14974 27490 14980 27524
rect 14934 27452 14980 27490
rect 14934 27418 14940 27452
rect 14974 27418 14980 27452
rect 14934 27380 14980 27418
rect 14934 27346 14940 27380
rect 14974 27346 14980 27380
rect 14934 27308 14980 27346
rect 14934 27274 14940 27308
rect 14974 27274 14980 27308
rect 14934 27236 14980 27274
rect 14934 27202 14940 27236
rect 14974 27202 14980 27236
rect 14934 27164 14980 27202
rect 14934 27130 14940 27164
rect 14974 27130 14980 27164
rect 14934 27092 14980 27130
rect 14934 27058 14940 27092
rect 14974 27058 14980 27092
rect 14934 27020 14980 27058
rect 14934 26986 14940 27020
rect 14974 26986 14980 27020
rect 14934 26948 14980 26986
rect 14934 26914 14940 26948
rect 14974 26914 14980 26948
rect 14934 26876 14980 26914
rect 14934 26842 14940 26876
rect 14974 26842 14980 26876
rect 14934 26804 14980 26842
rect 14934 26770 14940 26804
rect 14974 26770 14980 26804
rect 14934 26732 14980 26770
rect 14934 26698 14940 26732
rect 14974 26698 14980 26732
rect 14934 26660 14980 26698
rect 14934 26626 14940 26660
rect 14974 26626 14980 26660
rect 14934 26588 14980 26626
rect 14934 26554 14940 26588
rect 14974 26554 14980 26588
rect 14934 26516 14980 26554
rect 14934 26482 14940 26516
rect 14974 26482 14980 26516
rect 14934 26444 14980 26482
rect 14934 26410 14940 26444
rect 14974 26410 14980 26444
rect 14934 26372 14980 26410
rect 14934 26338 14940 26372
rect 14974 26338 14980 26372
rect 14934 26300 14980 26338
rect 14934 26266 14940 26300
rect 14974 26266 14980 26300
rect 14934 26228 14980 26266
rect 14934 26194 14940 26228
rect 14974 26194 14980 26228
rect 14934 26156 14980 26194
rect 14934 26122 14940 26156
rect 14974 26122 14980 26156
rect 14934 26084 14980 26122
rect 14934 26050 14940 26084
rect 14974 26050 14980 26084
rect 14934 26012 14980 26050
rect 14934 25978 14940 26012
rect 14974 25978 14980 26012
rect 14934 25940 14980 25978
rect 14934 25906 14940 25940
rect 14974 25906 14980 25940
rect 14934 25868 14980 25906
rect 14934 25834 14940 25868
rect 14974 25834 14980 25868
rect 14934 25796 14980 25834
rect 14934 25762 14940 25796
rect 14974 25762 14980 25796
rect 14934 25724 14980 25762
rect 14934 25690 14940 25724
rect 14974 25690 14980 25724
rect 14934 25652 14980 25690
rect 14934 25618 14940 25652
rect 14974 25618 14980 25652
rect 14934 25580 14980 25618
rect 14934 25546 14940 25580
rect 14974 25546 14980 25580
rect 14934 25508 14980 25546
rect 14934 25474 14940 25508
rect 14974 25474 14980 25508
rect 14934 25436 14980 25474
rect 14934 25402 14940 25436
rect 14974 25402 14980 25436
rect 14934 25364 14980 25402
rect 14934 25330 14940 25364
rect 14974 25330 14980 25364
rect 14934 25292 14980 25330
rect 14934 25258 14940 25292
rect 14974 25258 14980 25292
rect 14934 25220 14980 25258
rect 14934 25186 14940 25220
rect 14974 25186 14980 25220
rect 14934 25148 14980 25186
rect 14934 25114 14940 25148
rect 14974 25114 14980 25148
rect 14934 25076 14980 25114
rect 14934 25042 14940 25076
rect 14974 25042 14980 25076
rect 14934 25004 14980 25042
rect 14934 24970 14940 25004
rect 14974 24970 14980 25004
rect 14934 24932 14980 24970
rect 14934 24898 14940 24932
rect 14974 24898 14980 24932
rect 14934 24860 14980 24898
rect 14934 24826 14940 24860
rect 14974 24826 14980 24860
rect 14934 24788 14980 24826
rect 14934 24754 14940 24788
rect 14974 24754 14980 24788
rect 14934 24716 14980 24754
rect 14934 24682 14940 24716
rect 14974 24682 14980 24716
rect 14934 24644 14980 24682
rect 14934 24610 14940 24644
rect 14974 24610 14980 24644
rect 14934 24572 14980 24610
rect 14934 24538 14940 24572
rect 14974 24538 14980 24572
rect 14934 24500 14980 24538
rect 14934 24466 14940 24500
rect 14974 24466 14980 24500
rect 14934 24428 14980 24466
rect 14934 24394 14940 24428
rect 14974 24394 14980 24428
rect 14934 24356 14980 24394
rect 14934 24322 14940 24356
rect 14974 24322 14980 24356
rect 14934 24284 14980 24322
rect 14934 24250 14940 24284
rect 14974 24250 14980 24284
rect 14934 24212 14980 24250
rect 14934 24178 14940 24212
rect 14974 24178 14980 24212
rect 14934 24140 14980 24178
rect 14934 24106 14940 24140
rect 14974 24106 14980 24140
rect 14934 24068 14980 24106
rect 14934 24034 14940 24068
rect 14974 24034 14980 24068
rect 14934 23996 14980 24034
rect 14934 23962 14940 23996
rect 14974 23962 14980 23996
rect 14934 23924 14980 23962
rect 14934 23890 14940 23924
rect 14974 23890 14980 23924
rect 14934 23852 14980 23890
rect 14934 23818 14940 23852
rect 14974 23818 14980 23852
rect 14934 23780 14980 23818
rect 14934 23746 14940 23780
rect 14974 23746 14980 23780
rect 14934 23708 14980 23746
rect 14934 23674 14940 23708
rect 14974 23674 14980 23708
rect 14934 23636 14980 23674
rect 14934 23602 14940 23636
rect 14974 23602 14980 23636
rect 14934 23564 14980 23602
rect 14934 23530 14940 23564
rect 14974 23530 14980 23564
rect 14934 23492 14980 23530
rect 14934 23458 14940 23492
rect 14974 23458 14980 23492
rect 14934 23420 14980 23458
rect 14934 23386 14940 23420
rect 14974 23386 14980 23420
rect 14934 23348 14980 23386
rect 14934 23314 14940 23348
rect 14974 23314 14980 23348
rect 14934 23276 14980 23314
rect 14934 23242 14940 23276
rect 14974 23242 14980 23276
rect 14934 23204 14980 23242
rect 14934 23170 14940 23204
rect 14974 23170 14980 23204
rect 14934 23132 14980 23170
rect 14934 23098 14940 23132
rect 14974 23098 14980 23132
rect 14934 23060 14980 23098
rect 14934 23026 14940 23060
rect 14974 23026 14980 23060
rect 14934 22988 14980 23026
rect 14934 22954 14940 22988
rect 14974 22954 14980 22988
rect 14934 22916 14980 22954
rect 14934 22882 14940 22916
rect 14974 22882 14980 22916
rect 14934 22844 14980 22882
rect 14934 22810 14940 22844
rect 14974 22810 14980 22844
rect 14934 22772 14980 22810
rect 14934 22738 14940 22772
rect 14974 22738 14980 22772
rect 14934 22700 14980 22738
rect 14934 22666 14940 22700
rect 14974 22666 14980 22700
rect 14934 22628 14980 22666
rect 14934 22594 14940 22628
rect 14974 22594 14980 22628
rect 14934 22556 14980 22594
rect 14934 22522 14940 22556
rect 14974 22522 14980 22556
rect 14934 22484 14980 22522
rect 14934 22450 14940 22484
rect 14974 22450 14980 22484
rect 14934 22412 14980 22450
rect 14934 22378 14940 22412
rect 14974 22378 14980 22412
rect 14934 22340 14980 22378
rect 14934 22306 14940 22340
rect 14974 22306 14980 22340
rect 14934 22268 14980 22306
rect 14934 22234 14940 22268
rect 14974 22234 14980 22268
rect 14934 22196 14980 22234
rect 14934 22162 14940 22196
rect 14974 22162 14980 22196
rect 14934 22124 14980 22162
rect 14934 22090 14940 22124
rect 14974 22090 14980 22124
rect 14934 22052 14980 22090
rect 14934 22018 14940 22052
rect 14974 22018 14980 22052
rect 14934 21980 14980 22018
rect 14934 21946 14940 21980
rect 14974 21946 14980 21980
rect 14934 21908 14980 21946
rect 14934 21874 14940 21908
rect 14974 21874 14980 21908
rect 14934 21836 14980 21874
rect 14934 21802 14940 21836
rect 14974 21802 14980 21836
rect 14934 21764 14980 21802
rect 14934 21730 14940 21764
rect 14974 21730 14980 21764
rect 14934 21692 14980 21730
rect 14934 21658 14940 21692
rect 14974 21658 14980 21692
rect 14934 21620 14980 21658
rect 14934 21586 14940 21620
rect 14974 21586 14980 21620
rect 14934 21548 14980 21586
rect 14934 21514 14940 21548
rect 14974 21514 14980 21548
rect 14934 21476 14980 21514
rect 14934 21442 14940 21476
rect 14974 21442 14980 21476
rect 14934 21404 14980 21442
rect 14934 21370 14940 21404
rect 14974 21370 14980 21404
rect 14934 21332 14980 21370
rect 14934 21298 14940 21332
rect 14974 21298 14980 21332
rect 14934 21260 14980 21298
rect 14934 21226 14940 21260
rect 14974 21226 14980 21260
rect 14934 21188 14980 21226
rect 14934 21154 14940 21188
rect 14974 21154 14980 21188
rect 14934 21116 14980 21154
rect 14934 21082 14940 21116
rect 14974 21082 14980 21116
rect 14934 21044 14980 21082
rect 14934 21010 14940 21044
rect 14974 21010 14980 21044
rect 14934 20972 14980 21010
rect 14934 20938 14940 20972
rect 14974 20938 14980 20972
rect 14934 20900 14980 20938
rect 14934 20866 14940 20900
rect 14974 20866 14980 20900
rect 14934 20828 14980 20866
rect 14934 20794 14940 20828
rect 14974 20794 14980 20828
rect 14934 20756 14980 20794
rect 14934 20722 14940 20756
rect 14974 20722 14980 20756
rect 14934 20684 14980 20722
rect 14934 20650 14940 20684
rect 14974 20650 14980 20684
rect 14934 20612 14980 20650
rect 14934 20578 14940 20612
rect 14974 20578 14980 20612
rect 14934 20540 14980 20578
rect 14934 20506 14940 20540
rect 14974 20506 14980 20540
rect 14934 20468 14980 20506
rect 14934 20434 14940 20468
rect 14974 20434 14980 20468
rect 14934 20396 14980 20434
rect 14934 20362 14940 20396
rect 14974 20362 14980 20396
rect 14934 20324 14980 20362
rect 14934 20290 14940 20324
rect 14974 20290 14980 20324
rect 14934 20252 14980 20290
rect 14934 20218 14940 20252
rect 14974 20218 14980 20252
rect 14934 20180 14980 20218
rect 14934 20146 14940 20180
rect 14974 20146 14980 20180
rect 14934 20108 14980 20146
rect 14934 20074 14940 20108
rect 14974 20074 14980 20108
rect 14934 20036 14980 20074
rect 14934 20002 14940 20036
rect 14974 20002 14980 20036
rect 14934 19964 14980 20002
rect 14934 19930 14940 19964
rect 14974 19930 14980 19964
rect 14934 19892 14980 19930
rect 14934 19858 14940 19892
rect 14974 19858 14980 19892
rect 14934 19820 14980 19858
rect 14934 19786 14940 19820
rect 14974 19786 14980 19820
rect 14934 19748 14980 19786
rect 14934 19714 14940 19748
rect 14974 19714 14980 19748
rect 14934 19676 14980 19714
rect 14934 19642 14940 19676
rect 14974 19642 14980 19676
rect 14934 19604 14980 19642
rect 14934 19570 14940 19604
rect 14974 19570 14980 19604
rect 14934 19532 14980 19570
rect 14934 19498 14940 19532
rect 14974 19498 14980 19532
rect 14934 19460 14980 19498
rect 14934 19426 14940 19460
rect 14974 19426 14980 19460
rect 14934 19388 14980 19426
rect 14934 19354 14940 19388
rect 14974 19354 14980 19388
rect 14934 19316 14980 19354
rect 14934 19282 14940 19316
rect 14974 19282 14980 19316
rect 14934 19244 14980 19282
rect 14934 19210 14940 19244
rect 14974 19210 14980 19244
rect 14934 19172 14980 19210
rect 14934 19138 14940 19172
rect 14974 19138 14980 19172
rect 14934 19100 14980 19138
rect 14934 19066 14940 19100
rect 14974 19066 14980 19100
rect 14934 19028 14980 19066
rect 14934 18994 14940 19028
rect 14974 18994 14980 19028
rect 14934 18956 14980 18994
rect 14934 18922 14940 18956
rect 14974 18922 14980 18956
rect 14934 18884 14980 18922
rect 14934 18850 14940 18884
rect 14974 18850 14980 18884
rect 14934 18812 14980 18850
rect 14934 18778 14940 18812
rect 14974 18778 14980 18812
rect 14934 18740 14980 18778
rect 14934 18706 14940 18740
rect 14974 18706 14980 18740
rect 14934 18668 14980 18706
rect 14934 18634 14940 18668
rect 14974 18634 14980 18668
rect 14934 18596 14980 18634
rect 14934 18562 14940 18596
rect 14974 18562 14980 18596
rect 14934 18524 14980 18562
rect 14934 18490 14940 18524
rect 14974 18490 14980 18524
rect 14934 18452 14980 18490
rect 14934 18418 14940 18452
rect 14974 18418 14980 18452
rect 14934 18380 14980 18418
rect 14934 18346 14940 18380
rect 14974 18346 14980 18380
rect 14934 18308 14980 18346
rect 14934 18274 14940 18308
rect 14974 18274 14980 18308
rect 14934 18236 14980 18274
rect 14934 18202 14940 18236
rect 14974 18202 14980 18236
rect 14934 18164 14980 18202
rect 14934 18130 14940 18164
rect 14974 18130 14980 18164
rect 14934 18092 14980 18130
rect 14934 18058 14940 18092
rect 14974 18058 14980 18092
rect 14934 18020 14980 18058
rect 14934 17986 14940 18020
rect 14974 17986 14980 18020
rect 14934 17948 14980 17986
rect 14934 17914 14940 17948
rect 14974 17914 14980 17948
rect 14934 17876 14980 17914
rect 14934 17842 14940 17876
rect 14974 17842 14980 17876
rect 14934 17804 14980 17842
rect 14934 17770 14940 17804
rect 14974 17770 14980 17804
rect 14934 17732 14980 17770
rect 14934 17698 14940 17732
rect 14974 17698 14980 17732
rect 14934 17660 14980 17698
rect 14934 17626 14940 17660
rect 14974 17626 14980 17660
rect 14934 17588 14980 17626
rect 14934 17554 14940 17588
rect 14974 17554 14980 17588
rect 14934 17516 14980 17554
rect 14934 17482 14940 17516
rect 14974 17482 14980 17516
rect 14934 17444 14980 17482
rect 14934 17410 14940 17444
rect 14974 17410 14980 17444
rect 14934 17372 14980 17410
rect 14934 17338 14940 17372
rect 14974 17338 14980 17372
rect 14934 17300 14980 17338
rect 14934 17266 14940 17300
rect 14974 17266 14980 17300
rect 14934 17228 14980 17266
rect 14934 17194 14940 17228
rect 14974 17194 14980 17228
rect 14934 17156 14980 17194
rect 14934 17122 14940 17156
rect 14974 17122 14980 17156
rect 14934 17084 14980 17122
rect 14934 17050 14940 17084
rect 14974 17050 14980 17084
rect 14934 17012 14980 17050
rect 14934 16978 14940 17012
rect 14974 16978 14980 17012
rect 14934 16940 14980 16978
rect 14934 16906 14940 16940
rect 14974 16906 14980 16940
rect 14934 16868 14980 16906
rect 14934 16834 14940 16868
rect 14974 16834 14980 16868
rect 14934 16796 14980 16834
rect 14934 16762 14940 16796
rect 14974 16762 14980 16796
rect 14934 16724 14980 16762
rect 14934 16690 14940 16724
rect 14974 16690 14980 16724
rect 14934 16652 14980 16690
rect 14934 16618 14940 16652
rect 14974 16618 14980 16652
rect 14934 16580 14980 16618
rect 14934 16546 14940 16580
rect 14974 16546 14980 16580
rect 14934 16508 14980 16546
rect 14934 16474 14940 16508
rect 14974 16474 14980 16508
rect 14934 16436 14980 16474
rect 14934 16402 14940 16436
rect 14974 16402 14980 16436
rect 14934 16364 14980 16402
rect 14934 16330 14940 16364
rect 14974 16330 14980 16364
rect 14934 16292 14980 16330
rect 14934 16258 14940 16292
rect 14974 16258 14980 16292
rect 14934 16220 14980 16258
rect 14934 16186 14940 16220
rect 14974 16186 14980 16220
rect 14934 16148 14980 16186
rect 14934 16114 14940 16148
rect 14974 16114 14980 16148
rect 14934 16076 14980 16114
rect 14934 16042 14940 16076
rect 14974 16042 14980 16076
rect 14934 16004 14980 16042
rect 14934 15970 14940 16004
rect 14974 15970 14980 16004
rect 14934 15932 14980 15970
rect 14934 15898 14940 15932
rect 14974 15898 14980 15932
rect 14934 15860 14980 15898
rect 14934 15826 14940 15860
rect 14974 15826 14980 15860
rect 14934 15788 14980 15826
rect 14934 15754 14940 15788
rect 14974 15754 14980 15788
rect 14934 15716 14980 15754
rect 14934 15682 14940 15716
rect 14974 15682 14980 15716
rect 14934 15644 14980 15682
rect 14934 15610 14940 15644
rect 14974 15610 14980 15644
rect 14934 15572 14980 15610
rect 14934 15538 14940 15572
rect 14974 15538 14980 15572
rect 14934 15500 14980 15538
rect 14934 15466 14940 15500
rect 14974 15466 14980 15500
rect 14934 15428 14980 15466
rect 14934 15394 14940 15428
rect 14974 15394 14980 15428
rect 14934 15356 14980 15394
rect 14934 15322 14940 15356
rect 14974 15322 14980 15356
rect 14934 15284 14980 15322
rect 14934 15250 14940 15284
rect 14974 15250 14980 15284
rect 14934 15212 14980 15250
rect 14934 15178 14940 15212
rect 14974 15178 14980 15212
rect 14934 15140 14980 15178
rect 14934 15106 14940 15140
rect 14974 15106 14980 15140
rect 14934 15068 14980 15106
rect 14934 15034 14940 15068
rect 14974 15034 14980 15068
rect 14934 14996 14980 15034
rect 14934 14962 14940 14996
rect 14974 14962 14980 14996
rect 14934 14924 14980 14962
rect 14934 14890 14940 14924
rect 14974 14890 14980 14924
rect 14934 14852 14980 14890
rect 14934 14818 14940 14852
rect 14974 14818 14980 14852
rect 14934 14780 14980 14818
rect 14934 14746 14940 14780
rect 14974 14746 14980 14780
rect 14934 14708 14980 14746
rect 14934 14674 14940 14708
rect 14974 14674 14980 14708
rect 14934 14636 14980 14674
rect 14934 14602 14940 14636
rect 14974 14602 14980 14636
rect 14934 14564 14980 14602
rect 14934 14530 14940 14564
rect 14974 14530 14980 14564
rect 14934 14492 14980 14530
rect 14934 14458 14940 14492
rect 14974 14458 14980 14492
rect 14934 14420 14980 14458
rect 14934 14386 14940 14420
rect 14974 14386 14980 14420
rect 14934 14348 14980 14386
rect 14934 14314 14940 14348
rect 14974 14314 14980 14348
rect 14934 14276 14980 14314
rect 14934 14242 14940 14276
rect 14974 14242 14980 14276
rect 14934 14204 14980 14242
rect 14934 14170 14940 14204
rect 14974 14170 14980 14204
rect 14934 14132 14980 14170
rect 14934 14098 14940 14132
rect 14974 14098 14980 14132
rect 14934 14060 14980 14098
rect 14934 14026 14940 14060
rect 14974 14026 14980 14060
rect 14934 13988 14980 14026
rect 14934 13954 14940 13988
rect 14974 13954 14980 13988
rect 14934 13916 14980 13954
rect 14934 13882 14940 13916
rect 14974 13882 14980 13916
rect 14934 13844 14980 13882
rect 14934 13810 14940 13844
rect 14974 13810 14980 13844
rect 14934 13772 14980 13810
rect 14934 13738 14940 13772
rect 14974 13738 14980 13772
rect 14934 13700 14980 13738
rect 14934 13666 14940 13700
rect 14974 13666 14980 13700
rect 14934 13628 14980 13666
rect 14934 13594 14940 13628
rect 14974 13594 14980 13628
rect 14934 13556 14980 13594
rect 14934 13522 14940 13556
rect 14974 13522 14980 13556
rect 14934 13484 14980 13522
rect 14934 13450 14940 13484
rect 14974 13450 14980 13484
rect 14934 13412 14980 13450
rect 14934 13378 14940 13412
rect 14974 13378 14980 13412
rect 14934 13340 14980 13378
rect 14934 13306 14940 13340
rect 14974 13306 14980 13340
rect 14934 13268 14980 13306
rect 14934 13234 14940 13268
rect 14974 13234 14980 13268
rect 14934 13196 14980 13234
rect 14934 13162 14940 13196
rect 14974 13162 14980 13196
rect 14934 13124 14980 13162
rect 14934 13090 14940 13124
rect 14974 13090 14980 13124
rect 14934 13052 14980 13090
rect 14934 13018 14940 13052
rect 14974 13018 14980 13052
rect 14934 12980 14980 13018
rect 14934 12946 14940 12980
rect 14974 12946 14980 12980
rect 14934 12908 14980 12946
rect 14934 12874 14940 12908
rect 14974 12874 14980 12908
rect 14934 12836 14980 12874
rect 14934 12802 14940 12836
rect 14974 12802 14980 12836
rect 14934 12764 14980 12802
rect 14934 12730 14940 12764
rect 14974 12730 14980 12764
rect 14934 12692 14980 12730
rect 14934 12658 14940 12692
rect 14974 12658 14980 12692
rect 14934 12620 14980 12658
rect 14934 12586 14940 12620
rect 14974 12586 14980 12620
rect 14934 12548 14980 12586
rect 14934 12514 14940 12548
rect 14974 12514 14980 12548
rect 14934 12476 14980 12514
rect 14934 12442 14940 12476
rect 14974 12442 14980 12476
rect 14934 12404 14980 12442
rect 14934 12370 14940 12404
rect 14974 12370 14980 12404
rect 14934 12332 14980 12370
rect 14934 12298 14940 12332
rect 14974 12298 14980 12332
rect 14934 12260 14980 12298
rect 14934 12226 14940 12260
rect 14974 12226 14980 12260
rect 14934 12188 14980 12226
rect 14934 12154 14940 12188
rect 14974 12154 14980 12188
rect 14934 12116 14980 12154
rect 14934 12082 14940 12116
rect 14974 12082 14980 12116
rect 14934 12044 14980 12082
rect 14934 12010 14940 12044
rect 14974 12010 14980 12044
rect 14934 11972 14980 12010
rect 14934 11938 14940 11972
rect 14974 11938 14980 11972
rect 14934 11900 14980 11938
rect 14934 11866 14940 11900
rect 14974 11866 14980 11900
rect 14934 11828 14980 11866
rect 14934 11794 14940 11828
rect 14974 11794 14980 11828
rect 14934 11756 14980 11794
rect 14934 11722 14940 11756
rect 14974 11722 14980 11756
rect 14934 11684 14980 11722
rect 14934 11650 14940 11684
rect 14974 11650 14980 11684
rect 14934 11612 14980 11650
rect 14934 11578 14940 11612
rect 14974 11578 14980 11612
rect 14934 11540 14980 11578
rect 14934 11506 14940 11540
rect 14974 11506 14980 11540
rect 14934 11468 14980 11506
rect 14934 11434 14940 11468
rect 14974 11434 14980 11468
rect 14934 11396 14980 11434
rect 14934 11362 14940 11396
rect 14974 11362 14980 11396
rect 14934 11324 14980 11362
rect 14934 11290 14940 11324
rect 14974 11290 14980 11324
rect 14934 11252 14980 11290
rect 14934 11218 14940 11252
rect 14974 11218 14980 11252
rect 14934 11180 14980 11218
rect 14934 11146 14940 11180
rect 14974 11146 14980 11180
rect 14934 11108 14980 11146
rect 14934 11074 14940 11108
rect 14974 11074 14980 11108
rect 14934 11036 14980 11074
rect 14934 11002 14940 11036
rect 14974 11002 14980 11036
rect 14934 10964 14980 11002
rect 14934 10930 14940 10964
rect 14974 10930 14980 10964
rect 14934 10892 14980 10930
rect 14934 10858 14940 10892
rect 14974 10858 14980 10892
rect 14934 10820 14980 10858
rect 14934 10786 14940 10820
rect 14974 10786 14980 10820
rect 14934 10748 14980 10786
rect 14934 10714 14940 10748
rect 14974 10714 14980 10748
rect 14934 10676 14980 10714
rect 14934 10642 14940 10676
rect 14974 10642 14980 10676
rect 14934 10604 14980 10642
rect 14934 10570 14940 10604
rect 14974 10570 14980 10604
rect 14934 10532 14980 10570
rect 14934 10498 14940 10532
rect 14974 10498 14980 10532
rect 14934 10460 14980 10498
rect 14934 10426 14940 10460
rect 14974 10426 14980 10460
rect 14934 10388 14980 10426
rect 14934 10354 14940 10388
rect 14974 10354 14980 10388
rect 14934 10316 14980 10354
rect 14934 10282 14940 10316
rect 14974 10282 14980 10316
rect 14934 10244 14980 10282
rect 14934 10210 14940 10244
rect 14974 10210 14980 10244
rect 14934 10172 14980 10210
rect 14934 10138 14940 10172
rect 14974 10138 14980 10172
rect 14934 10100 14980 10138
rect 14934 10066 14940 10100
rect 14974 10066 14980 10100
rect 14934 10028 14980 10066
rect 14934 9994 14940 10028
rect 14974 9994 14980 10028
rect 14934 9956 14980 9994
rect 14934 9922 14940 9956
rect 14974 9922 14980 9956
rect 14934 9884 14980 9922
rect 14934 9850 14940 9884
rect 14974 9850 14980 9884
rect 14934 9812 14980 9850
rect 14934 9778 14940 9812
rect 14974 9778 14980 9812
rect 14934 9740 14980 9778
rect 14934 9706 14940 9740
rect 14974 9706 14980 9740
rect 14934 9668 14980 9706
rect 14934 9634 14940 9668
rect 14974 9634 14980 9668
rect 14934 9596 14980 9634
rect 14934 9562 14940 9596
rect 14974 9562 14980 9596
rect 14934 9524 14980 9562
rect 14934 9490 14940 9524
rect 14974 9490 14980 9524
rect 14934 9452 14980 9490
rect 14934 9418 14940 9452
rect 14974 9418 14980 9452
rect 14934 9380 14980 9418
rect 14934 9346 14940 9380
rect 14974 9346 14980 9380
rect 14934 9308 14980 9346
rect 14934 9274 14940 9308
rect 14974 9274 14980 9308
rect 14934 9236 14980 9274
rect 14934 9202 14940 9236
rect 14974 9202 14980 9236
rect 14934 9164 14980 9202
rect 14934 9130 14940 9164
rect 14974 9130 14980 9164
rect 14934 9092 14980 9130
rect 14934 9058 14940 9092
rect 14974 9058 14980 9092
rect 14934 9020 14980 9058
rect 14934 8986 14940 9020
rect 14974 8986 14980 9020
rect 14934 8948 14980 8986
rect 14934 8914 14940 8948
rect 14974 8914 14980 8948
rect 14934 8876 14980 8914
rect 14934 8842 14940 8876
rect 14974 8842 14980 8876
rect 14934 8804 14980 8842
rect 14934 8770 14940 8804
rect 14974 8770 14980 8804
rect 14934 8732 14980 8770
rect 14934 8698 14940 8732
rect 14974 8698 14980 8732
rect 14934 8660 14980 8698
rect 14934 8626 14940 8660
rect 14974 8626 14980 8660
rect 14934 8588 14980 8626
rect 14934 8554 14940 8588
rect 14974 8554 14980 8588
rect 14934 8516 14980 8554
rect 14934 8482 14940 8516
rect 14974 8482 14980 8516
rect 14934 8444 14980 8482
rect 14934 8410 14940 8444
rect 14974 8410 14980 8444
rect 14934 8372 14980 8410
rect 14934 8338 14940 8372
rect 14974 8338 14980 8372
rect 14934 8300 14980 8338
rect 14934 8266 14940 8300
rect 14974 8266 14980 8300
rect 14934 8228 14980 8266
rect 14934 8194 14940 8228
rect 14974 8194 14980 8228
rect 14934 8156 14980 8194
rect 14934 8122 14940 8156
rect 14974 8122 14980 8156
rect 14934 8084 14980 8122
rect 14934 8050 14940 8084
rect 14974 8050 14980 8084
rect 14934 8012 14980 8050
rect 14934 7978 14940 8012
rect 14974 7978 14980 8012
rect 14934 7940 14980 7978
rect 14934 7906 14940 7940
rect 14974 7906 14980 7940
rect 14934 7868 14980 7906
rect 14934 7834 14940 7868
rect 14974 7834 14980 7868
rect 14934 7796 14980 7834
rect 14934 7762 14940 7796
rect 14974 7762 14980 7796
rect 14934 7724 14980 7762
rect 14934 7690 14940 7724
rect 14974 7690 14980 7724
rect 14934 7652 14980 7690
rect 14934 7618 14940 7652
rect 14974 7618 14980 7652
rect 14934 7580 14980 7618
rect 14934 7546 14940 7580
rect 14974 7546 14980 7580
rect 14934 7508 14980 7546
rect 14934 7474 14940 7508
rect 14974 7474 14980 7508
rect 14934 7436 14980 7474
rect 14934 7402 14940 7436
rect 14974 7402 14980 7436
rect 14934 7364 14980 7402
rect 14934 7330 14940 7364
rect 14974 7330 14980 7364
rect 14934 7292 14980 7330
rect 14934 7258 14940 7292
rect 14974 7258 14980 7292
rect 14934 7220 14980 7258
rect 14934 7186 14940 7220
rect 14974 7186 14980 7220
rect 14934 7148 14980 7186
rect 14934 7114 14940 7148
rect 14974 7114 14980 7148
rect 14934 7076 14980 7114
rect 14934 7042 14940 7076
rect 14974 7042 14980 7076
rect 14934 7004 14980 7042
rect 14934 6970 14940 7004
rect 14974 6970 14980 7004
rect 14934 6932 14980 6970
rect 14934 6898 14940 6932
rect 14974 6898 14980 6932
rect 14934 6860 14980 6898
rect 14934 6826 14940 6860
rect 14974 6826 14980 6860
rect 14934 6788 14980 6826
rect 14934 6754 14940 6788
rect 14974 6754 14980 6788
rect 14934 6716 14980 6754
rect 14934 6682 14940 6716
rect 14974 6682 14980 6716
rect 14934 6644 14980 6682
rect 14934 6610 14940 6644
rect 14974 6610 14980 6644
rect 14934 6572 14980 6610
rect 14934 6538 14940 6572
rect 14974 6538 14980 6572
rect 14934 6500 14980 6538
rect 14934 6466 14940 6500
rect 14974 6466 14980 6500
rect 14934 6428 14980 6466
rect 14934 6394 14940 6428
rect 14974 6394 14980 6428
rect 14934 6356 14980 6394
rect 14934 6322 14940 6356
rect 14974 6322 14980 6356
rect 14934 6284 14980 6322
rect 14934 6250 14940 6284
rect 14974 6250 14980 6284
rect 14934 6212 14980 6250
rect 14934 6178 14940 6212
rect 14974 6178 14980 6212
rect 14934 6140 14980 6178
rect 14934 6106 14940 6140
rect 14974 6106 14980 6140
rect 14934 6068 14980 6106
rect 14934 6034 14940 6068
rect 14974 6034 14980 6068
rect 14934 5996 14980 6034
rect 14934 5962 14940 5996
rect 14974 5962 14980 5996
rect 14934 5924 14980 5962
rect 14934 5890 14940 5924
rect 14974 5890 14980 5924
rect 14934 5852 14980 5890
rect 14934 5818 14940 5852
rect 14974 5818 14980 5852
rect 14934 5780 14980 5818
rect 14934 5746 14940 5780
rect 14974 5746 14980 5780
rect 14934 5708 14980 5746
rect 14934 5674 14940 5708
rect 14974 5674 14980 5708
rect 14934 5636 14980 5674
rect 14934 5602 14940 5636
rect 14974 5602 14980 5636
rect 14934 5564 14980 5602
rect 14934 5530 14940 5564
rect 14974 5530 14980 5564
rect 14934 5492 14980 5530
rect 14934 5458 14940 5492
rect 14974 5458 14980 5492
rect 14934 5420 14980 5458
rect 14934 5386 14940 5420
rect 14974 5386 14980 5420
rect 14934 5348 14980 5386
rect 14934 5314 14940 5348
rect 14974 5314 14980 5348
rect 14934 5276 14980 5314
rect 14934 5242 14940 5276
rect 14974 5242 14980 5276
rect 14934 5204 14980 5242
rect 14934 5170 14940 5204
rect 14974 5170 14980 5204
rect 14934 5132 14980 5170
rect 14934 5098 14940 5132
rect 14974 5098 14980 5132
rect 14934 5060 14980 5098
rect 14934 5026 14940 5060
rect 14974 5026 14980 5060
rect 14934 4988 14980 5026
rect 14934 4954 14940 4988
rect 14974 4954 14980 4988
rect 14934 4916 14980 4954
rect 14934 4882 14940 4916
rect 14974 4882 14980 4916
rect 14934 4844 14980 4882
rect 14934 4810 14940 4844
rect 14974 4810 14980 4844
rect 14934 4772 14980 4810
rect 14934 4738 14940 4772
rect 14974 4738 14980 4772
rect 14934 4700 14980 4738
rect 14934 4666 14940 4700
rect 14974 4666 14980 4700
rect 14934 4628 14980 4666
rect 14934 4594 14940 4628
rect 14974 4594 14980 4628
rect 14934 4556 14980 4594
rect 14934 4522 14940 4556
rect 14974 4522 14980 4556
rect 14934 4484 14980 4522
rect 14934 4450 14940 4484
rect 14974 4450 14980 4484
rect 14934 4412 14980 4450
rect 14934 4378 14940 4412
rect 14974 4378 14980 4412
rect 14934 4340 14980 4378
rect 14934 4306 14940 4340
rect 14974 4306 14980 4340
rect 14934 4268 14980 4306
rect 14934 4234 14940 4268
rect 14974 4234 14980 4268
rect 14934 4196 14980 4234
rect 14934 4162 14940 4196
rect 14974 4162 14980 4196
rect 14934 4124 14980 4162
rect 14934 4090 14940 4124
rect 14974 4090 14980 4124
rect 14934 4052 14980 4090
rect 14934 4018 14940 4052
rect 14974 4018 14980 4052
rect 14934 3980 14980 4018
rect 14934 3946 14940 3980
rect 14974 3946 14980 3980
rect 14934 3908 14980 3946
rect 14934 3874 14940 3908
rect 14974 3874 14980 3908
rect 14934 3836 14980 3874
rect 14934 3802 14940 3836
rect 14974 3802 14980 3836
rect 14934 3764 14980 3802
rect 14934 3730 14940 3764
rect 14974 3730 14980 3764
rect 14934 3692 14980 3730
rect 14934 3658 14940 3692
rect 14974 3658 14980 3692
rect 14934 3620 14980 3658
rect 14934 3586 14940 3620
rect 14974 3586 14980 3620
rect 14934 3548 14980 3586
rect 14934 3514 14940 3548
rect 14974 3514 14980 3548
rect 14934 3476 14980 3514
rect 14934 3442 14940 3476
rect 14974 3442 14980 3476
rect 14934 3404 14980 3442
rect 14934 3370 14940 3404
rect 14974 3370 14980 3404
rect 14934 3332 14980 3370
rect 14934 3298 14940 3332
rect 14974 3298 14980 3332
rect 14934 3260 14980 3298
rect 14934 3226 14940 3260
rect 14974 3226 14980 3260
rect 14934 3188 14980 3226
rect 14934 3154 14940 3188
rect 14974 3154 14980 3188
rect 14934 3116 14980 3154
rect 14934 3082 14940 3116
rect 14974 3082 14980 3116
rect 14934 3044 14980 3082
rect 14934 3010 14940 3044
rect 14974 3010 14980 3044
rect 14934 2972 14980 3010
rect 14934 2938 14940 2972
rect 14974 2938 14980 2972
rect 14934 2900 14980 2938
rect 14934 2866 14940 2900
rect 14974 2866 14980 2900
rect 14934 2828 14980 2866
rect 14934 2794 14940 2828
rect 14974 2794 14980 2828
rect 14934 2756 14980 2794
rect 14934 2722 14940 2756
rect 14974 2722 14980 2756
rect 14934 2684 14980 2722
rect 14934 2650 14940 2684
rect 14974 2650 14980 2684
rect 14934 2612 14980 2650
rect 14934 2578 14940 2612
rect 14974 2578 14980 2612
rect 14934 2540 14980 2578
rect 14934 2506 14940 2540
rect 14974 2506 14980 2540
rect 14934 2468 14980 2506
rect 14934 2434 14940 2468
rect 14974 2434 14980 2468
rect 14934 2396 14980 2434
rect 14934 2362 14940 2396
rect 14974 2362 14980 2396
rect 14934 2324 14980 2362
rect 14934 2290 14940 2324
rect 14974 2290 14980 2324
rect 14934 2252 14980 2290
rect 14934 2218 14940 2252
rect 14974 2218 14980 2252
rect 14934 2180 14980 2218
rect 14934 2146 14940 2180
rect 14974 2146 14980 2180
rect 14934 2108 14980 2146
rect 14934 2074 14940 2108
rect 14974 2074 14980 2108
rect 14934 2036 14980 2074
rect 14934 2002 14940 2036
rect 14974 2002 14980 2036
rect 14934 1964 14980 2002
rect 14934 1930 14940 1964
rect 14974 1930 14980 1964
rect 14934 1892 14980 1930
rect 14934 1858 14940 1892
rect 14974 1858 14980 1892
rect 14934 1820 14980 1858
rect 14934 1786 14940 1820
rect 14974 1786 14980 1820
rect 14934 1748 14980 1786
rect 14934 1714 14940 1748
rect 14974 1714 14980 1748
rect 14934 1676 14980 1714
rect 14934 1642 14940 1676
rect 14974 1642 14980 1676
rect 14934 1604 14980 1642
rect 14934 1570 14940 1604
rect 14974 1570 14980 1604
rect 14934 1532 14980 1570
rect 14934 1498 14940 1532
rect 14974 1498 14980 1532
rect 14934 1460 14980 1498
rect 14934 1426 14940 1460
rect 14974 1426 14980 1460
rect 14934 1387 14980 1426
rect 14934 1353 14940 1387
rect 14974 1353 14980 1387
rect 14934 1314 14980 1353
rect 14934 1280 14940 1314
rect 14974 1280 14980 1314
rect 14934 1241 14980 1280
rect 14934 1207 14940 1241
rect 14974 1207 14980 1241
rect 14934 1168 14980 1207
rect 14934 1134 14940 1168
rect 14974 1134 14980 1168
rect 14934 1095 14980 1134
rect 14934 1061 14940 1095
rect 14974 1061 14980 1095
rect 14934 1022 14980 1061
rect 14934 988 14940 1022
rect 14974 988 14980 1022
rect 14934 949 14980 988
rect 14934 915 14940 949
rect 14974 915 14980 949
rect 14934 876 14980 915
rect 14934 842 14940 876
rect 14974 842 14980 876
rect 14934 803 14980 842
rect 14934 769 14940 803
rect 14974 769 14980 803
rect 14934 730 14980 769
rect 14934 696 14940 730
rect 14974 696 14980 730
rect 14934 657 14980 696
rect 14934 623 14940 657
rect 14974 623 14980 657
rect 14934 584 14980 623
rect 14934 550 14940 584
rect 14974 550 14980 584
rect 14934 511 14980 550
rect 14934 477 14940 511
rect 14974 477 14980 511
rect 14934 438 14980 477
rect 13206 362 13252 400
rect 14811 417 14857 429
rect 14811 383 14817 417
rect 14851 383 14857 417
rect 13206 328 13212 362
rect 13246 328 13252 362
tri 14792 345 14811 364 se
rect 14811 345 14857 383
tri 14777 330 14792 345 se
rect 14792 330 14817 345
rect 11418 259 11424 293
rect 11458 259 11464 293
rect 11418 220 11464 259
rect 11418 186 11424 220
rect 11458 186 11464 220
rect 11418 147 11464 186
rect 11418 113 11424 147
rect 11458 113 11464 147
rect 13206 290 13252 328
rect 13206 256 13212 290
rect 13246 256 13252 290
rect 13976 326 14817 330
rect 13976 274 13982 326
rect 14034 274 14046 326
rect 14098 324 14817 326
rect 14098 290 14648 324
rect 14682 290 14720 324
rect 14754 311 14817 324
rect 14851 311 14857 345
rect 14754 290 14857 311
rect 14098 274 14857 290
rect 13976 270 14857 274
rect 14934 404 14940 438
rect 14974 404 14980 438
rect 14934 365 14980 404
rect 14934 331 14940 365
rect 14974 331 14980 365
rect 14934 292 14980 331
rect 13206 218 13252 256
rect 13206 184 13212 218
rect 13246 184 13252 218
rect 13206 146 13252 184
rect 11418 112 11464 113
tri 11464 112 11466 114 sw
tri 13204 112 13206 114 se
rect 13206 112 13212 146
rect 13246 112 13252 146
rect 14934 258 14940 292
rect 14974 258 14980 292
rect 14934 219 14980 258
rect 14934 185 14940 219
rect 14974 185 14980 219
rect 14934 146 14980 185
tri 13252 112 13254 114 sw
tri 14932 112 14934 114 se
rect 14934 112 14940 146
rect 14974 112 14980 146
rect 11418 80 11466 112
tri 11466 80 11498 112 sw
tri 13172 80 13204 112 se
rect 13204 80 13254 112
tri 13254 80 13286 112 sw
tri 14900 80 14932 112 se
rect 14932 80 14980 112
rect 11418 74 14980 80
rect 11418 40 11496 74
rect 11530 40 11570 74
rect 11604 40 11644 74
rect 11678 40 11718 74
rect 11752 40 11792 74
rect 11826 40 11866 74
rect 11900 40 11940 74
rect 11974 40 12014 74
rect 12048 40 12088 74
rect 12122 40 12162 74
rect 12196 40 12236 74
rect 12270 40 12310 74
rect 12344 40 12384 74
rect 12418 40 12458 74
rect 12492 40 12531 74
rect 12565 40 12604 74
rect 12638 40 12677 74
rect 12711 40 12750 74
rect 12784 40 12823 74
rect 12857 40 12896 74
rect 12930 40 12969 74
rect 13003 40 13042 74
rect 13076 40 13115 74
rect 13149 40 13188 74
rect 13222 40 13261 74
rect 13295 40 13334 74
rect 13368 40 13407 74
rect 13441 40 13480 74
rect 13514 40 13553 74
rect 13587 40 13626 74
rect 13660 40 13699 74
rect 13733 40 13772 74
rect 13806 40 13845 74
rect 13879 40 13918 74
rect 13952 40 13991 74
rect 14025 40 14064 74
rect 14098 40 14137 74
rect 14171 40 14210 74
rect 14244 40 14283 74
rect 14317 40 14356 74
rect 14390 40 14429 74
rect 14463 40 14502 74
rect 14536 40 14575 74
rect 14609 40 14648 74
rect 14682 40 14721 74
rect 14755 40 14794 74
rect 14828 40 14867 74
rect 14901 40 14980 74
rect 11418 34 14980 40
rect 11595 -149 13058 -129
tri 13058 -149 13078 -129 sw
rect 11595 -155 14789 -149
rect 11595 -189 11607 -155
rect 11641 -189 11679 -155
rect 11713 -189 11751 -155
rect 11785 -189 11823 -155
rect 11857 -189 11896 -155
rect 11930 -189 11969 -155
rect 12003 -189 12042 -155
rect 12076 -189 12115 -155
rect 12149 -189 12188 -155
rect 12222 -189 12261 -155
rect 12295 -189 12334 -155
rect 12368 -189 12407 -155
rect 12441 -189 12480 -155
rect 12514 -189 12553 -155
rect 12587 -189 12626 -155
rect 12660 -189 12699 -155
rect 12733 -189 12772 -155
rect 12806 -189 12845 -155
rect 12879 -189 12918 -155
rect 12952 -189 12991 -155
rect 13025 -189 13064 -155
rect 13098 -189 13137 -155
rect 13171 -189 13210 -155
rect 13244 -189 13283 -155
rect 13317 -189 13356 -155
rect 13390 -189 13429 -155
rect 13463 -189 13502 -155
rect 13536 -189 13575 -155
rect 13609 -189 13648 -155
rect 13682 -189 13721 -155
rect 13755 -189 13794 -155
rect 13828 -189 13867 -155
rect 13901 -189 13940 -155
rect 13974 -189 14013 -155
rect 14047 -189 14086 -155
rect 14120 -189 14159 -155
rect 14193 -189 14232 -155
rect 14266 -189 14305 -155
rect 14339 -189 14378 -155
rect 14412 -189 14451 -155
rect 14485 -189 14524 -155
rect 14558 -189 14597 -155
rect 14631 -189 14670 -155
rect 14704 -189 14743 -155
rect 14777 -189 14789 -155
rect 11595 -195 14789 -189
rect 11595 -266 13058 -195
tri 13058 -229 13092 -195 nw
rect 11595 -300 11771 -266
rect 11805 -300 12083 -266
rect 12117 -300 12395 -266
rect 12429 -300 12707 -266
rect 12741 -300 13018 -266
rect 13052 -300 13058 -266
rect 11595 -348 13058 -300
rect 11595 -354 11771 -348
tri 11731 -382 11759 -354 ne
rect 11759 -382 11771 -354
rect 11805 -354 12083 -348
rect 11805 -382 11817 -354
tri 11817 -382 11845 -354 nw
tri 12043 -382 12071 -354 ne
rect 12071 -382 12083 -354
rect 12117 -354 12395 -348
rect 12117 -382 12129 -354
tri 12129 -382 12157 -354 nw
tri 12355 -382 12383 -354 ne
rect 12383 -382 12395 -354
rect 12429 -354 12707 -348
rect 12429 -382 12441 -354
tri 12441 -382 12469 -354 nw
tri 12667 -382 12695 -354 ne
rect 12695 -382 12707 -354
rect 12741 -354 13018 -348
rect 12741 -382 12753 -354
tri 12753 -382 12781 -354 nw
tri 12978 -382 13006 -354 ne
rect 13006 -382 13018 -354
rect 13052 -382 13058 -348
tri 11759 -386 11763 -382 ne
rect 11763 -386 11813 -382
tri 11813 -386 11817 -382 nw
tri 12071 -386 12075 -382 ne
rect 12075 -386 12125 -382
tri 12125 -386 12129 -382 nw
tri 12383 -386 12387 -382 ne
rect 12387 -386 12437 -382
tri 12437 -386 12441 -382 nw
tri 12695 -386 12699 -382 ne
rect 12699 -386 12749 -382
tri 12749 -386 12753 -382 nw
tri 13006 -386 13010 -382 ne
rect 13010 -386 13058 -382
rect 13325 -266 14619 -254
rect 13325 -300 13331 -266
rect 13365 -300 13643 -266
rect 13677 -300 13955 -266
rect 13989 -278 14267 -266
rect 13325 -330 13982 -300
rect 14034 -330 14046 -278
rect 14098 -300 14267 -278
rect 14301 -300 14579 -266
rect 14613 -300 14619 -266
rect 14098 -330 14619 -300
rect 13325 -348 14619 -330
rect 13325 -382 13331 -348
rect 13365 -354 13643 -348
rect 13365 -382 13377 -354
tri 13377 -382 13405 -354 nw
tri 13603 -382 13631 -354 ne
rect 13631 -382 13643 -354
rect 13677 -354 13955 -348
rect 13677 -382 13689 -354
tri 13689 -382 13717 -354 nw
tri 13915 -382 13943 -354 ne
rect 13943 -382 13955 -354
rect 13989 -354 14267 -348
rect 13989 -382 14001 -354
tri 14001 -382 14029 -354 nw
tri 14227 -382 14255 -354 ne
rect 14255 -382 14267 -354
rect 14301 -354 14579 -348
rect 14301 -382 14313 -354
tri 14313 -382 14341 -354 nw
tri 14539 -382 14567 -354 ne
rect 14567 -382 14579 -354
rect 14613 -382 14619 -348
rect 13325 -386 13373 -382
tri 13373 -386 13377 -382 nw
tri 13631 -386 13635 -382 ne
rect 13635 -386 13685 -382
tri 13685 -386 13689 -382 nw
tri 13943 -386 13947 -382 ne
rect 13947 -386 13997 -382
tri 13997 -386 14001 -382 nw
tri 14255 -386 14259 -382 ne
rect 14259 -386 14309 -382
tri 14309 -386 14313 -382 nw
tri 14567 -386 14571 -382 ne
rect 14571 -386 14619 -382
rect 11609 -398 11655 -386
tri 11763 -388 11765 -386 ne
rect 11609 -432 11615 -398
rect 11649 -432 11655 -398
rect 11609 -473 11655 -432
rect 11609 -507 11615 -473
rect 11649 -507 11655 -473
rect 11609 -548 11655 -507
rect 11609 -582 11615 -548
rect 11649 -582 11655 -548
rect 11609 -623 11655 -582
rect 11609 -657 11615 -623
rect 11649 -657 11655 -623
rect 11609 -698 11655 -657
rect 11609 -732 11615 -698
rect 11649 -732 11655 -698
rect 11765 -430 11811 -386
tri 11811 -388 11813 -386 nw
rect 11765 -464 11771 -430
rect 11805 -464 11811 -430
rect 11765 -512 11811 -464
rect 11765 -546 11771 -512
rect 11805 -546 11811 -512
rect 11765 -594 11811 -546
rect 11765 -628 11771 -594
rect 11805 -628 11811 -594
rect 11765 -677 11811 -628
rect 11765 -711 11771 -677
rect 11805 -711 11811 -677
rect 11765 -723 11811 -711
rect 11921 -398 11967 -386
tri 12075 -388 12077 -386 ne
rect 11921 -432 11927 -398
rect 11961 -432 11967 -398
rect 11921 -473 11967 -432
rect 11921 -507 11927 -473
rect 11961 -507 11967 -473
rect 11921 -548 11967 -507
rect 11921 -582 11927 -548
rect 11961 -582 11967 -548
rect 11921 -623 11967 -582
rect 11921 -657 11927 -623
rect 11961 -657 11967 -623
rect 11921 -698 11967 -657
rect 11609 -771 11655 -732
rect 11921 -732 11927 -698
rect 11961 -732 11967 -698
rect 12077 -430 12123 -386
tri 12123 -388 12125 -386 nw
rect 12077 -464 12083 -430
rect 12117 -464 12123 -430
rect 12077 -512 12123 -464
rect 12077 -546 12083 -512
rect 12117 -546 12123 -512
rect 12077 -594 12123 -546
rect 12077 -628 12083 -594
rect 12117 -628 12123 -594
rect 12077 -677 12123 -628
rect 12077 -711 12083 -677
rect 12117 -711 12123 -677
rect 12077 -723 12123 -711
rect 12233 -398 12279 -386
tri 12387 -388 12389 -386 ne
rect 12233 -432 12239 -398
rect 12273 -432 12279 -398
rect 12233 -473 12279 -432
rect 12233 -507 12239 -473
rect 12273 -507 12279 -473
rect 12233 -548 12279 -507
rect 12233 -582 12239 -548
rect 12273 -582 12279 -548
rect 12233 -623 12279 -582
rect 12233 -657 12239 -623
rect 12273 -657 12279 -623
rect 12233 -698 12279 -657
tri 11655 -771 11689 -737 sw
tri 11887 -771 11921 -737 se
rect 11921 -771 11967 -732
rect 12233 -732 12239 -698
rect 12273 -732 12279 -698
rect 12389 -430 12435 -386
tri 12435 -388 12437 -386 nw
rect 12389 -464 12395 -430
rect 12429 -464 12435 -430
rect 12389 -512 12435 -464
rect 12389 -546 12395 -512
rect 12429 -546 12435 -512
rect 12389 -594 12435 -546
rect 12389 -628 12395 -594
rect 12429 -628 12435 -594
rect 12389 -677 12435 -628
rect 12389 -711 12395 -677
rect 12429 -711 12435 -677
rect 12389 -723 12435 -711
rect 12545 -398 12591 -386
tri 12699 -388 12701 -386 ne
rect 12545 -432 12551 -398
rect 12585 -432 12591 -398
rect 12545 -473 12591 -432
rect 12545 -507 12551 -473
rect 12585 -507 12591 -473
rect 12545 -548 12591 -507
rect 12545 -582 12551 -548
rect 12585 -582 12591 -548
rect 12545 -623 12591 -582
rect 12545 -657 12551 -623
rect 12585 -657 12591 -623
rect 12545 -698 12591 -657
tri 11967 -771 12001 -737 sw
tri 12199 -771 12233 -737 se
rect 12233 -771 12279 -732
rect 12545 -732 12551 -698
rect 12585 -732 12591 -698
rect 12701 -430 12747 -386
tri 12747 -388 12749 -386 nw
rect 12701 -464 12707 -430
rect 12741 -464 12747 -430
rect 12701 -512 12747 -464
rect 12701 -546 12707 -512
rect 12741 -546 12747 -512
rect 12701 -594 12747 -546
rect 12701 -628 12707 -594
rect 12741 -628 12747 -594
rect 12701 -677 12747 -628
rect 12701 -711 12707 -677
rect 12741 -711 12747 -677
rect 12701 -723 12747 -711
rect 12857 -398 12903 -386
tri 13010 -388 13012 -386 ne
rect 12857 -432 12863 -398
rect 12897 -432 12903 -398
rect 12857 -473 12903 -432
rect 12857 -507 12863 -473
rect 12897 -507 12903 -473
rect 12857 -548 12903 -507
rect 12857 -582 12863 -548
rect 12897 -582 12903 -548
rect 12857 -623 12903 -582
rect 12857 -657 12863 -623
rect 12897 -657 12903 -623
rect 12857 -698 12903 -657
tri 12279 -771 12313 -737 sw
tri 12511 -771 12545 -737 se
rect 12545 -771 12591 -732
rect 12857 -732 12863 -698
rect 12897 -732 12903 -698
rect 13012 -430 13058 -386
rect 13012 -464 13018 -430
rect 13052 -464 13058 -430
rect 13012 -512 13058 -464
rect 13012 -546 13018 -512
rect 13052 -546 13058 -512
rect 13012 -594 13058 -546
rect 13012 -628 13018 -594
rect 13052 -628 13058 -594
rect 13012 -677 13058 -628
rect 13012 -711 13018 -677
rect 13052 -711 13058 -677
rect 13012 -723 13058 -711
rect 13169 -398 13215 -386
rect 13169 -432 13175 -398
rect 13209 -432 13215 -398
rect 13169 -473 13215 -432
rect 13169 -507 13175 -473
rect 13209 -507 13215 -473
rect 13169 -548 13215 -507
rect 13169 -582 13175 -548
rect 13209 -582 13215 -548
rect 13169 -623 13215 -582
rect 13169 -657 13175 -623
rect 13209 -657 13215 -623
rect 13169 -698 13215 -657
tri 12591 -771 12625 -737 sw
tri 12823 -771 12857 -737 se
rect 12857 -771 12903 -732
rect 13169 -732 13175 -698
rect 13209 -732 13215 -698
rect 13325 -430 13371 -386
tri 13371 -388 13373 -386 nw
rect 13325 -464 13331 -430
rect 13365 -464 13371 -430
rect 13325 -512 13371 -464
rect 13325 -546 13331 -512
rect 13365 -546 13371 -512
rect 13325 -594 13371 -546
rect 13325 -628 13331 -594
rect 13365 -628 13371 -594
rect 13325 -677 13371 -628
rect 13325 -711 13331 -677
rect 13365 -711 13371 -677
rect 13325 -723 13371 -711
rect 13481 -398 13527 -386
tri 13635 -388 13637 -386 ne
rect 13481 -432 13487 -398
rect 13521 -432 13527 -398
rect 13481 -473 13527 -432
rect 13481 -507 13487 -473
rect 13521 -507 13527 -473
rect 13481 -548 13527 -507
rect 13481 -582 13487 -548
rect 13521 -582 13527 -548
rect 13481 -623 13527 -582
rect 13481 -657 13487 -623
rect 13521 -657 13527 -623
rect 13481 -698 13527 -657
tri 12903 -771 12937 -737 sw
tri 13135 -771 13169 -737 se
rect 13169 -771 13215 -732
rect 13481 -732 13487 -698
rect 13521 -732 13527 -698
rect 13637 -430 13683 -386
tri 13683 -388 13685 -386 nw
rect 13637 -464 13643 -430
rect 13677 -464 13683 -430
rect 13637 -512 13683 -464
rect 13637 -546 13643 -512
rect 13677 -546 13683 -512
rect 13637 -594 13683 -546
rect 13637 -628 13643 -594
rect 13677 -628 13683 -594
rect 13637 -677 13683 -628
rect 13637 -711 13643 -677
rect 13677 -711 13683 -677
rect 13637 -723 13683 -711
rect 13793 -398 13839 -386
tri 13947 -388 13949 -386 ne
rect 13793 -432 13799 -398
rect 13833 -432 13839 -398
rect 13793 -473 13839 -432
rect 13793 -507 13799 -473
rect 13833 -507 13839 -473
rect 13793 -548 13839 -507
rect 13793 -582 13799 -548
rect 13833 -582 13839 -548
rect 13793 -623 13839 -582
rect 13793 -657 13799 -623
rect 13833 -657 13839 -623
rect 13793 -698 13839 -657
tri 13215 -771 13249 -737 sw
tri 13447 -771 13481 -737 se
rect 13481 -771 13527 -732
rect 13793 -732 13799 -698
rect 13833 -732 13839 -698
rect 13949 -430 13995 -386
tri 13995 -388 13997 -386 nw
rect 13949 -464 13955 -430
rect 13989 -464 13995 -430
rect 13949 -512 13995 -464
rect 13949 -546 13955 -512
rect 13989 -546 13995 -512
rect 13949 -594 13995 -546
rect 13949 -628 13955 -594
rect 13989 -628 13995 -594
rect 13949 -677 13995 -628
rect 13949 -711 13955 -677
rect 13989 -711 13995 -677
rect 13949 -723 13995 -711
rect 14105 -398 14151 -386
tri 14259 -388 14261 -386 ne
rect 14105 -432 14111 -398
rect 14145 -432 14151 -398
rect 14105 -473 14151 -432
rect 14105 -507 14111 -473
rect 14145 -507 14151 -473
rect 14105 -548 14151 -507
rect 14105 -582 14111 -548
rect 14145 -582 14151 -548
rect 14105 -623 14151 -582
rect 14105 -657 14111 -623
rect 14145 -657 14151 -623
rect 14105 -698 14151 -657
tri 13527 -771 13561 -737 sw
tri 13759 -771 13793 -737 se
rect 13793 -771 13839 -732
rect 14105 -732 14111 -698
rect 14145 -732 14151 -698
rect 14261 -430 14307 -386
tri 14307 -388 14309 -386 nw
rect 14261 -464 14267 -430
rect 14301 -464 14307 -430
rect 14261 -512 14307 -464
rect 14261 -546 14267 -512
rect 14301 -546 14307 -512
rect 14261 -594 14307 -546
rect 14261 -628 14267 -594
rect 14301 -628 14307 -594
rect 14261 -677 14307 -628
rect 14261 -711 14267 -677
rect 14301 -711 14307 -677
rect 14261 -723 14307 -711
rect 14417 -398 14463 -386
tri 14571 -388 14573 -386 ne
rect 14417 -432 14423 -398
rect 14457 -432 14463 -398
rect 14417 -473 14463 -432
rect 14417 -507 14423 -473
rect 14457 -507 14463 -473
rect 14417 -548 14463 -507
rect 14417 -582 14423 -548
rect 14457 -582 14463 -548
rect 14417 -623 14463 -582
rect 14417 -657 14423 -623
rect 14457 -657 14463 -623
rect 14417 -698 14463 -657
tri 13839 -771 13873 -737 sw
tri 14071 -771 14105 -737 se
rect 14105 -771 14151 -732
rect 14417 -732 14423 -698
rect 14457 -732 14463 -698
rect 14573 -430 14619 -386
rect 14573 -464 14579 -430
rect 14613 -464 14619 -430
rect 14573 -512 14619 -464
rect 14573 -546 14579 -512
rect 14613 -546 14619 -512
rect 14573 -594 14619 -546
rect 14573 -628 14579 -594
rect 14613 -628 14619 -594
rect 14573 -677 14619 -628
rect 14573 -711 14579 -677
rect 14613 -711 14619 -677
rect 14573 -723 14619 -711
rect 14729 -362 14775 -350
rect 14729 -396 14735 -362
rect 14769 -396 14775 -362
rect 14729 -444 14775 -396
rect 14729 -478 14735 -444
rect 14769 -478 14775 -444
rect 14729 -526 14775 -478
rect 14729 -560 14735 -526
rect 14769 -560 14775 -526
rect 14729 -608 14775 -560
rect 14729 -642 14735 -608
rect 14769 -642 14775 -608
rect 14729 -690 14775 -642
tri 14151 -771 14185 -737 sw
tri 14383 -771 14417 -737 se
rect 14417 -771 14463 -732
rect 14729 -724 14735 -690
rect 14769 -724 14775 -690
tri 14463 -771 14497 -737 sw
tri 14695 -771 14729 -737 se
rect 14729 -771 14775 -724
rect 11609 -773 14775 -771
rect 11609 -807 11615 -773
rect 11649 -807 11927 -773
rect 11961 -807 12239 -773
rect 12273 -807 12551 -773
rect 12585 -807 12863 -773
rect 12897 -807 13175 -773
rect 13209 -807 13487 -773
rect 13521 -807 13799 -773
rect 13833 -807 14111 -773
rect 14145 -807 14423 -773
rect 14457 -807 14735 -773
rect 14769 -807 14775 -773
rect 11609 -871 14775 -807
rect 11678 -917 14724 -911
rect 11678 -951 11690 -917
rect 11724 -951 11762 -917
rect 11796 -951 11834 -917
rect 11868 -951 11906 -917
rect 11940 -951 11978 -917
rect 12012 -951 12050 -917
rect 12084 -951 12123 -917
rect 12157 -951 12196 -917
rect 12230 -951 12269 -917
rect 12303 -951 12342 -917
rect 12376 -951 12415 -917
rect 12449 -951 12488 -917
rect 12522 -951 12561 -917
rect 12595 -951 12634 -917
rect 12668 -951 12707 -917
rect 12741 -951 12780 -917
rect 12814 -951 12853 -917
rect 12887 -951 12926 -917
rect 12960 -951 12999 -917
rect 13033 -951 13072 -917
rect 13106 -951 13145 -917
rect 13179 -951 13218 -917
rect 13252 -951 13291 -917
rect 13325 -951 13364 -917
rect 13398 -951 13437 -917
rect 13471 -951 13510 -917
rect 13544 -951 13583 -917
rect 13617 -951 13656 -917
rect 13690 -951 13729 -917
rect 13763 -951 13802 -917
rect 13836 -951 13875 -917
rect 13909 -951 13948 -917
rect 13982 -951 14021 -917
rect 14055 -951 14094 -917
rect 14128 -951 14167 -917
rect 14201 -951 14240 -917
rect 14274 -951 14313 -917
rect 14347 -951 14386 -917
rect 14420 -951 14459 -917
rect 14493 -951 14532 -917
rect 14566 -951 14605 -917
rect 14639 -951 14678 -917
rect 14712 -951 14724 -917
rect 11678 -957 14724 -951
<< via1 >>
rect -135 4576 -83 4628
rect -135 4512 -83 4564
rect -135 3486 -83 3492
rect -135 3452 -126 3486
rect -126 3452 -92 3486
rect -92 3452 -83 3486
rect -135 3440 -83 3452
rect -135 3414 -83 3428
rect -135 3380 -126 3414
rect -126 3380 -92 3414
rect -92 3380 -83 3414
rect -135 3376 -83 3380
rect 1635 3486 1687 3492
rect 1635 3452 1644 3486
rect 1644 3452 1678 3486
rect 1678 3452 1687 3486
rect 1635 3440 1687 3452
rect 1635 3414 1687 3428
rect 1635 3380 1644 3414
rect 1644 3380 1678 3414
rect 1678 3380 1687 3414
rect 1635 3376 1687 3380
rect 2007 3486 2059 3492
rect 2007 3452 2016 3486
rect 2016 3452 2050 3486
rect 2050 3452 2059 3486
rect 2007 3440 2059 3452
rect 2007 3414 2059 3428
rect 2007 3380 2016 3414
rect 2016 3380 2050 3414
rect 2050 3380 2059 3414
rect 2007 3376 2059 3380
rect 3777 3486 3829 3492
rect 3777 3452 3786 3486
rect 3786 3452 3820 3486
rect 3820 3452 3829 3486
rect 3777 3440 3829 3452
rect 3777 3414 3829 3428
rect 3777 3380 3786 3414
rect 3786 3380 3820 3414
rect 3820 3380 3829 3414
rect 3777 3376 3829 3380
rect 4149 3487 4201 3492
rect 4149 3453 4158 3487
rect 4158 3453 4192 3487
rect 4192 3453 4201 3487
rect 4149 3440 4201 3453
rect 4149 3415 4201 3428
rect 4149 3381 4158 3415
rect 4158 3381 4192 3415
rect 4192 3381 4201 3415
rect 4149 3376 4201 3381
rect 5919 3486 5971 3492
rect 5919 3452 5928 3486
rect 5928 3452 5962 3486
rect 5962 3452 5971 3486
rect 5919 3440 5971 3452
rect 5919 3414 5971 3428
rect 5919 3380 5928 3414
rect 5928 3380 5962 3414
rect 5962 3380 5971 3414
rect 5919 3376 5971 3380
rect 9205 3487 9257 3493
rect 9205 3453 9214 3487
rect 9214 3453 9248 3487
rect 9248 3453 9257 3487
rect 9205 3441 9257 3453
rect 9205 3415 9257 3429
rect 9205 3381 9214 3415
rect 9214 3381 9248 3415
rect 9248 3381 9257 3415
rect 9205 3377 9257 3381
rect 10031 3487 10083 3493
rect 10031 3453 10040 3487
rect 10040 3453 10074 3487
rect 10074 3453 10083 3487
rect 10031 3441 10083 3453
rect 10031 3415 10083 3429
rect 10031 3381 10040 3415
rect 10040 3381 10074 3415
rect 10074 3381 10083 3415
rect 10031 3377 10083 3381
rect 12886 38615 12938 38624
rect 12886 38581 12892 38615
rect 12892 38581 12926 38615
rect 12926 38581 12938 38615
rect 13000 38612 13052 38624
rect 12886 38572 12938 38581
rect 13000 38578 13038 38612
rect 13038 38578 13052 38612
rect 13000 38572 13052 38578
rect 10403 3487 10455 3493
rect 10403 3453 10412 3487
rect 10412 3453 10446 3487
rect 10446 3453 10455 3487
rect 10403 3441 10455 3453
rect 10403 3415 10455 3429
rect 10403 3381 10412 3415
rect 10412 3381 10446 3415
rect 10446 3381 10455 3415
rect 10403 3377 10455 3381
rect 11229 3487 11281 3493
rect 11229 3453 11238 3487
rect 11238 3453 11272 3487
rect 11272 3453 11281 3487
rect 11229 3441 11281 3453
rect 11229 3415 11281 3429
rect 11229 3381 11238 3415
rect 11238 3381 11272 3415
rect 11272 3381 11281 3415
rect 11229 3377 11281 3381
rect 13412 38612 13464 38624
rect 13526 38615 13578 38624
rect 13412 38578 13426 38612
rect 13426 38578 13464 38612
rect 13526 38581 13538 38615
rect 13538 38581 13572 38615
rect 13572 38581 13578 38615
rect 13412 38572 13464 38578
rect 13526 38572 13578 38581
rect -129 3076 -77 3128
rect -65 3076 -13 3128
rect 11601 3441 11653 3493
rect 11601 3377 11653 3429
rect 13982 274 14034 326
rect 14046 274 14098 326
rect 13982 -300 13989 -278
rect 13989 -300 14034 -278
rect 13982 -330 14034 -300
rect 14046 -330 14098 -278
<< metal2 >>
rect 12880 38572 12886 38624
rect 12938 38572 13000 38624
rect 13052 38572 13412 38624
rect 13464 38572 13526 38624
rect 13578 38572 13584 38624
rect -135 4628 -83 4634
rect -135 4564 -83 4576
rect -135 4506 -83 4512
rect -135 3492 -83 3498
rect -135 3428 -83 3440
rect -135 3128 -83 3376
rect 1635 3492 2076 3498
rect 1687 3440 2007 3492
rect 2059 3440 2076 3492
rect 1635 3428 2076 3440
rect 1687 3376 2007 3428
rect 2059 3376 2076 3428
rect 1635 3370 2076 3376
rect 3777 3492 4201 3498
rect 3829 3440 4149 3492
rect 3777 3428 4201 3440
rect 3829 3376 4149 3428
rect 3777 3370 4201 3376
rect 5919 3492 5971 3498
rect 9205 3493 9257 3499
tri 5971 3441 5986 3456 sw
tri 9190 3441 9205 3456 se
rect 5971 3440 5986 3441
rect 5919 3429 5986 3440
tri 5986 3429 5998 3441 sw
tri 9178 3429 9190 3441 se
rect 9190 3429 9257 3441
rect 5919 3428 5998 3429
rect 5971 3422 5998 3428
tri 5998 3422 6005 3429 sw
tri 9171 3422 9178 3429 se
rect 9178 3422 9205 3429
rect 5971 3377 9205 3422
rect 5971 3376 9257 3377
rect 5919 3370 9257 3376
rect 10031 3493 10455 3499
rect 10083 3441 10403 3493
rect 10031 3429 10455 3441
rect 10083 3377 10403 3429
rect 10031 3371 10455 3377
rect 11229 3493 11653 3499
rect 11281 3441 11601 3493
rect 11229 3429 11653 3441
rect 11281 3377 11601 3429
rect 11229 3371 11653 3377
tri -83 3128 -49 3162 sw
rect -135 3076 -129 3128
rect -77 3076 -65 3128
rect -13 3076 -7 3128
rect 13976 326 14104 330
rect 13976 274 13982 326
rect 14034 274 14046 326
rect 14098 274 14104 326
rect 13976 -278 14104 274
rect 13976 -330 13982 -278
rect 14034 -330 14046 -278
rect 14098 -330 14104 -278
rect 13976 -354 14104 -330
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_0
timestamp 1701704242
transform 0 -1 3124 -1 0 3402
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_1
timestamp 1701704242
transform 0 -1 3006 -1 0 3402
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_2
timestamp 1701704242
transform 0 -1 3360 -1 0 3402
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_3
timestamp 1701704242
transform 0 -1 3242 -1 0 3402
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_4
timestamp 1701704242
transform 0 -1 3596 -1 0 3402
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_5
timestamp 1701704242
transform 0 -1 3478 -1 0 3402
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_6
timestamp 1701704242
transform 0 -1 3714 -1 0 3402
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_7
timestamp 1701704242
transform 0 -1 3832 -1 0 3402
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_8
timestamp 1701704242
transform 0 -1 982 -1 0 3402
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_9
timestamp 1701704242
transform 0 -1 864 -1 0 3402
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_10
timestamp 1701704242
transform 0 -1 1218 -1 0 3402
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_11
timestamp 1701704242
transform 0 -1 1100 -1 0 3402
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_12
timestamp 1701704242
transform 0 -1 1454 -1 0 3402
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_13
timestamp 1701704242
transform 0 -1 1336 -1 0 3402
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_14
timestamp 1701704242
transform 0 -1 5974 -1 0 3403
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_15
timestamp 1701704242
transform 0 -1 5856 -1 0 3403
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_16
timestamp 1701704242
transform 0 -1 5620 -1 0 3403
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_17
timestamp 1701704242
transform 0 -1 5738 -1 0 3403
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_18
timestamp 1701704242
transform 0 -1 5384 -1 0 3403
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_19
timestamp 1701704242
transform 0 -1 5502 -1 0 3403
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_20
timestamp 1701704242
transform 0 -1 5148 -1 0 3403
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_21
timestamp 1701704242
transform 0 -1 5266 -1 0 3403
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_22
timestamp 1701704242
transform 0 -1 11770 -1 0 333
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_23
timestamp 1701704242
transform 0 -1 13562 -1 0 38623
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_24
timestamp 1701704242
transform 0 -1 12954 -1 0 38623
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_25
timestamp 1701704242
transform 0 -1 14742 -1 0 333
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_26
timestamp 1701704242
transform 0 -1 13444 -1 0 38623
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_27
timestamp 1701704242
transform 0 -1 13072 -1 0 38623
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_28
timestamp 1701704242
transform 0 -1 1572 -1 0 3402
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_29
timestamp 1701704242
transform 0 -1 1690 -1 0 3402
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_30
timestamp 1701704242
transform 0 -1 11284 -1 0 3403
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_31
timestamp 1701704242
transform 0 -1 10576 -1 0 3403
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_32
timestamp 1701704242
transform 0 -1 10458 -1 0 3403
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_33
timestamp 1701704242
transform 0 -1 10812 -1 0 3403
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_34
timestamp 1701704242
transform 0 -1 10694 -1 0 3403
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_35
timestamp 1701704242
transform 0 -1 11048 -1 0 3403
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_36
timestamp 1701704242
transform 0 -1 10930 -1 0 3403
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_37
timestamp 1701704242
transform 0 -1 11166 -1 0 3403
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_38
timestamp 1701704242
transform 0 -1 14860 -1 0 333
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_39
timestamp 1701704242
transform 0 -1 11656 -1 0 333
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_40
timestamp 1701704242
transform 0 1 2004 -1 0 3402
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_41
timestamp 1701704242
transform 0 1 2122 -1 0 3402
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_42
timestamp 1701704242
transform 0 1 2358 -1 0 3402
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_43
timestamp 1701704242
transform 0 1 2240 -1 0 3402
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_44
timestamp 1701704242
transform 0 1 2594 -1 0 3402
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_45
timestamp 1701704242
transform 0 1 2476 -1 0 3402
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_46
timestamp 1701704242
transform 0 1 2830 -1 0 3402
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_47
timestamp 1701704242
transform 0 1 2712 -1 0 3402
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_48
timestamp 1701704242
transform 0 1 570 -1 0 3402
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_49
timestamp 1701704242
transform 0 1 688 -1 0 3402
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_50
timestamp 1701704242
transform 0 1 4854 -1 0 3403
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_51
timestamp 1701704242
transform 0 1 4972 -1 0 3403
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_52
timestamp 1701704242
transform 0 1 4618 -1 0 3403
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_53
timestamp 1701704242
transform 0 1 4736 -1 0 3403
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_54
timestamp 1701704242
transform 0 1 4382 -1 0 3403
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_55
timestamp 1701704242
transform 0 1 4500 -1 0 3403
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_56
timestamp 1701704242
transform 0 1 4264 -1 0 3403
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_57
timestamp 1701704242
transform 0 1 4146 -1 0 3403
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_58
timestamp 1701704242
transform 0 1 334 -1 0 3402
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_59
timestamp 1701704242
transform 0 1 452 -1 0 3402
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_60
timestamp 1701704242
transform 0 1 98 -1 0 3402
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_61
timestamp 1701704242
transform 0 1 -20 -1 0 3402
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_62
timestamp 1701704242
transform 0 1 9202 -1 0 3403
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_63
timestamp 1701704242
transform 0 1 9320 -1 0 3403
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_64
timestamp 1701704242
transform 0 1 9556 -1 0 3403
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_65
timestamp 1701704242
transform 0 1 9438 -1 0 3403
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_66
timestamp 1701704242
transform 0 1 9792 -1 0 3403
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_67
timestamp 1701704242
transform 0 1 9674 -1 0 3403
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_68
timestamp 1701704242
transform 0 1 10028 -1 0 3403
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_69
timestamp 1701704242
transform 0 1 9910 -1 0 3403
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_70
timestamp 1701704242
transform 0 1 216 -1 0 3402
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_71
timestamp 1701704242
transform 0 1 -138 -1 0 3402
box 0 0 1 1
use nDFbentRes_CDNS_52468879185818  nDFbentRes_CDNS_52468879185818_0
timestamp 1701704242
transform 0 -1 13444 -1 0 38471
box -68 -1442 38104 84
use nDFbentRes_CDNS_52468879185818  nDFbentRes_CDNS_52468879185818_1
timestamp 1701704242
transform 0 -1 11656 1 0 435
box -68 -1442 38104 84
use nDFbentRes_CDNS_52468879185819  nDFbentRes_CDNS_52468879185819_0
timestamp 1701704242
transform 0 1 2594 1 0 3504
box -68 -144 35034 84
use nDFbentRes_CDNS_52468879185819  nDFbentRes_CDNS_52468879185819_1
timestamp 1701704242
transform 0 1 2830 1 0 3504
box -68 -144 35034 84
use nDFbentRes_CDNS_52468879185819  nDFbentRes_CDNS_52468879185819_2
timestamp 1701704242
transform 0 1 2122 1 0 3504
box -68 -144 35034 84
use nDFbentRes_CDNS_52468879185819  nDFbentRes_CDNS_52468879185819_3
timestamp 1701704242
transform 0 1 2358 1 0 3504
box -68 -144 35034 84
use nDFbentRes_CDNS_52468879185819  nDFbentRes_CDNS_52468879185819_4
timestamp 1701704242
transform 0 1 4500 1 0 3505
box -68 -144 35034 84
use nDFbentRes_CDNS_52468879185819  nDFbentRes_CDNS_52468879185819_5
timestamp 1701704242
transform 0 1 4264 1 0 3505
box -68 -144 35034 84
use nDFbentRes_CDNS_52468879185819  nDFbentRes_CDNS_52468879185819_6
timestamp 1701704242
transform 0 1 4972 1 0 3505
box -68 -144 35034 84
use nDFbentRes_CDNS_52468879185819  nDFbentRes_CDNS_52468879185819_7
timestamp 1701704242
transform 0 1 4736 1 0 3505
box -68 -144 35034 84
use nDFbentRes_CDNS_52468879185819  nDFbentRes_CDNS_52468879185819_8
timestamp 1701704242
transform 0 1 -20 1 0 3504
box -68 -144 35034 84
use nDFbentRes_CDNS_52468879185819  nDFbentRes_CDNS_52468879185819_9
timestamp 1701704242
transform 0 1 216 1 0 3504
box -68 -144 35034 84
use nDFbentRes_CDNS_52468879185819  nDFbentRes_CDNS_52468879185819_10
timestamp 1701704242
transform 0 1 688 1 0 3504
box -68 -144 35034 84
use nDFbentRes_CDNS_52468879185819  nDFbentRes_CDNS_52468879185819_11
timestamp 1701704242
transform 0 1 452 1 0 3504
box -68 -144 35034 84
use nDFbentRes_CDNS_52468879185819  nDFbentRes_CDNS_52468879185819_12
timestamp 1701704242
transform 0 1 9792 1 0 3505
box -68 -144 35034 84
use nDFbentRes_CDNS_52468879185819  nDFbentRes_CDNS_52468879185819_13
timestamp 1701704242
transform 0 1 10028 1 0 3505
box -68 -144 35034 84
use nDFbentRes_CDNS_52468879185819  nDFbentRes_CDNS_52468879185819_14
timestamp 1701704242
transform 0 1 9320 1 0 3505
box -68 -144 35034 84
use nDFbentRes_CDNS_52468879185819  nDFbentRes_CDNS_52468879185819_15
timestamp 1701704242
transform 0 1 9556 1 0 3505
box -68 -144 35034 84
use nDFbentRes_CDNS_52468879185819  nDFbentRes_CDNS_52468879185819_16
timestamp 1701704242
transform 0 -1 3478 1 0 3504
box -68 -144 35034 84
use nDFbentRes_CDNS_52468879185819  nDFbentRes_CDNS_52468879185819_17
timestamp 1701704242
transform 0 -1 3714 1 0 3504
box -68 -144 35034 84
use nDFbentRes_CDNS_52468879185819  nDFbentRes_CDNS_52468879185819_18
timestamp 1701704242
transform 0 -1 3006 1 0 3504
box -68 -144 35034 84
use nDFbentRes_CDNS_52468879185819  nDFbentRes_CDNS_52468879185819_19
timestamp 1701704242
transform 0 -1 3242 1 0 3504
box -68 -144 35034 84
use nDFbentRes_CDNS_52468879185819  nDFbentRes_CDNS_52468879185819_20
timestamp 1701704242
transform 0 -1 1100 1 0 3504
box -68 -144 35034 84
use nDFbentRes_CDNS_52468879185819  nDFbentRes_CDNS_52468879185819_21
timestamp 1701704242
transform 0 -1 864 1 0 3504
box -68 -144 35034 84
use nDFbentRes_CDNS_52468879185819  nDFbentRes_CDNS_52468879185819_22
timestamp 1701704242
transform 0 -1 5384 1 0 3505
box -68 -144 35034 84
use nDFbentRes_CDNS_52468879185819  nDFbentRes_CDNS_52468879185819_23
timestamp 1701704242
transform 0 -1 5148 1 0 3505
box -68 -144 35034 84
use nDFbentRes_CDNS_52468879185819  nDFbentRes_CDNS_52468879185819_24
timestamp 1701704242
transform 0 -1 5856 1 0 3505
box -68 -144 35034 84
use nDFbentRes_CDNS_52468879185819  nDFbentRes_CDNS_52468879185819_25
timestamp 1701704242
transform 0 -1 5620 1 0 3505
box -68 -144 35034 84
use nDFbentRes_CDNS_52468879185819  nDFbentRes_CDNS_52468879185819_26
timestamp 1701704242
transform 0 -1 10930 1 0 3505
box -68 -144 35034 84
use nDFbentRes_CDNS_52468879185819  nDFbentRes_CDNS_52468879185819_27
timestamp 1701704242
transform 0 -1 11166 1 0 3505
box -68 -144 35034 84
use nDFbentRes_CDNS_52468879185819  nDFbentRes_CDNS_52468879185819_28
timestamp 1701704242
transform 0 -1 10458 1 0 3505
box -68 -144 35034 84
use nDFbentRes_CDNS_52468879185819  nDFbentRes_CDNS_52468879185819_29
timestamp 1701704242
transform 0 -1 10694 1 0 3505
box -68 -144 35034 84
use nDFbentRes_CDNS_52468879185819  nDFbentRes_CDNS_52468879185819_30
timestamp 1701704242
transform 0 -1 1336 1 0 3504
box -68 -144 35034 84
use nDFbentRes_CDNS_52468879185819  nDFbentRes_CDNS_52468879185819_31
timestamp 1701704242
transform 0 -1 1572 1 0 3504
box -68 -144 35034 84
use nfet_CDNS_52468879185820  nfet_CDNS_52468879185820_0
timestamp 1701704242
transform -1 0 14724 0 -1 -269
box -79 -32 1583 632
use nfet_CDNS_52468879185820  nfet_CDNS_52468879185820_1
timestamp 1701704242
transform -1 0 13164 0 -1 -269
box -79 -32 1583 632
use pfet_CDNS_52468879185817  pfet_CDNS_52468879185817_0
timestamp 1701704242
transform 0 -1 5866 -1 0 2550
box -119 -66 1623 666
<< labels >>
flabel metal1 s 12724 -946 12875 -915 3 FreeSans 200 0 0 0 vrefgen_en_h
port 1 nsew
flabel metal1 s 5188 1817 5213 1971 3 FreeSans 200 0 0 0 vrefgen_en_h_n
port 2 nsew
flabel metal1 s -3 3384 37 3473 3 FreeSans 200 0 0 0 vref<31>
port 3 nsew
flabel metal1 s 224 3389 266 3486 3 FreeSans 200 0 0 0 vref<30>
port 4 nsew
flabel metal1 s 462 3381 505 3486 3 FreeSans 200 0 0 0 vref<29>
port 5 nsew
flabel metal1 s 699 3387 740 3486 3 FreeSans 200 0 0 0 vref<28>
port 6 nsew
flabel metal1 s 936 3389 974 3485 3 FreeSans 200 0 0 0 vref<27>
port 7 nsew
flabel metal1 s 1172 3388 1209 3484 3 FreeSans 200 0 0 0 vref<26>
port 8 nsew
flabel metal1 s 1409 3385 1447 3485 3 FreeSans 200 0 0 0 vref<25>
port 9 nsew
flabel metal1 s 1644 3386 1680 3483 3 FreeSans 200 0 0 0 vref<24>
port 10 nsew
flabel metal1 s 2138 3386 2178 3482 3 FreeSans 200 0 0 0 vref<23>
port 11 nsew
flabel metal1 s 2369 3394 2409 3483 3 FreeSans 200 0 0 0 vref<22>
port 12 nsew
flabel metal1 s 2608 3385 2636 3479 3 FreeSans 200 0 0 0 vref<21>
port 13 nsew
flabel metal1 s 2838 3388 2880 3488 3 FreeSans 200 0 0 0 vref<20>
port 14 nsew
flabel metal1 s 3077 3388 3115 3485 3 FreeSans 200 0 0 0 vref<19>
port 15 nsew
flabel metal1 s 3311 3385 3349 3488 3 FreeSans 200 0 0 0 vref<18>
port 16 nsew
flabel metal1 s 3546 3379 3584 3485 3 FreeSans 200 0 0 0 vref<17>
port 17 nsew
flabel metal1 s 3784 3389 3822 3487 3 FreeSans 200 0 0 0 vref<16>
port 18 nsew
flabel metal1 s 4275 3387 4312 3486 3 FreeSans 200 0 0 0 vref<15>
port 19 nsew
flabel metal1 s 4509 3390 4550 3484 3 FreeSans 200 0 0 0 vref<14>
port 20 nsew
flabel metal1 s 4749 3378 4788 3482 3 FreeSans 200 0 0 0 vref<13>
port 21 nsew
flabel metal1 s 4988 3383 5022 3488 3 FreeSans 200 0 0 0 vref<12>
port 22 nsew
flabel metal1 s 5217 3382 5258 3487 3 FreeSans 200 0 0 0 vref<11>
port 23 nsew
flabel metal1 s 5463 3382 5496 3482 3 FreeSans 200 0 0 0 vref<10>
port 24 nsew
flabel metal1 s 5693 3379 5727 3478 3 FreeSans 200 0 0 0 vref<9>
port 25 nsew
flabel metal1 s 5932 3390 5962 3477 3 FreeSans 200 0 0 0 vref<8>
port 26 nsew
flabel metal1 s 9334 3393 9367 3485 3 FreeSans 200 0 0 0 vref<7>
port 27 nsew
flabel metal1 s 9569 3381 9604 3480 3 FreeSans 200 0 0 0 vref<6>
port 28 nsew
flabel metal1 s 9800 3393 9841 3483 3 FreeSans 200 0 0 0 vref<5>
port 29 nsew
flabel metal1 s 10040 3390 10077 3480 3 FreeSans 200 0 0 0 vref<4>
port 30 nsew
flabel metal1 s 10529 3393 10564 3480 3 FreeSans 200 0 0 0 vref<3>
port 31 nsew
flabel metal1 s 10769 3393 10797 3479 3 FreeSans 200 0 0 0 vref<2>
port 32 nsew
flabel metal1 s 11011 3387 11033 3472 3 FreeSans 200 0 0 0 vref<1>
port 33 nsew
flabel metal1 s 11237 3398 11270 3484 3 FreeSans 200 0 0 0 vref<0>
port 34 nsew
flabel metal1 s 12117 -260 12751 -175 3 FreeSans 200 90 0 0 vssd
port 35 nsew
flabel metal1 s 5906 1374 6012 1596 3 FreeSans 200 180 0 0 vddio_q
port 36 nsew
<< properties >>
string GDS_END 25716498
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 24813098
string path -3.375 77.550 -0.175 77.550 
<< end >>
