magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< pwell >>
rect -191 -26 8021 1026
<< nmos >>
rect 0 0 36 1000
rect 270 0 306 1000
rect 836 0 872 1000
rect 1106 0 1142 1000
rect 1672 0 1708 1000
rect 1942 0 1978 1000
rect 2508 0 2544 1000
rect 2778 0 2814 1000
rect 3344 0 3380 1000
rect 3614 0 3650 1000
rect 4180 0 4216 1000
rect 4450 0 4486 1000
rect 5016 0 5052 1000
rect 5286 0 5322 1000
rect 5852 0 5888 1000
rect 6122 0 6158 1000
rect 6688 0 6724 1000
rect 6958 0 6994 1000
rect 7524 0 7560 1000
rect 7794 0 7830 1000
<< ndiff >>
rect -165 0 0 1000
rect 36 0 270 1000
rect 306 0 471 1000
rect 671 0 836 1000
rect 872 0 1106 1000
rect 1142 0 1307 1000
rect 1507 0 1672 1000
rect 1708 0 1942 1000
rect 1978 0 2143 1000
rect 2343 0 2508 1000
rect 2544 0 2778 1000
rect 2814 0 2979 1000
rect 3179 0 3344 1000
rect 3380 0 3614 1000
rect 3650 0 3815 1000
rect 4015 0 4180 1000
rect 4216 0 4450 1000
rect 4486 0 4651 1000
rect 4851 0 5016 1000
rect 5052 0 5286 1000
rect 5322 0 5487 1000
rect 5687 0 5852 1000
rect 5888 0 6122 1000
rect 6158 0 6323 1000
rect 6523 0 6688 1000
rect 6724 0 6958 1000
rect 6994 0 7159 1000
rect 7359 0 7524 1000
rect 7560 0 7794 1000
rect 7830 0 7995 1000
<< poly >>
rect 0 1000 36 1032
rect 270 1000 306 1032
rect 836 1000 872 1032
rect 1106 1000 1142 1032
rect 1672 1000 1708 1032
rect 1942 1000 1978 1032
rect 2508 1000 2544 1032
rect 2778 1000 2814 1032
rect 3344 1000 3380 1032
rect 3614 1000 3650 1032
rect 4180 1000 4216 1032
rect 4450 1000 4486 1032
rect 5016 1000 5052 1032
rect 5286 1000 5322 1032
rect 5852 1000 5888 1032
rect 6122 1000 6158 1032
rect 6688 1000 6724 1032
rect 6958 1000 6994 1032
rect 7524 1000 7560 1032
rect 7794 1000 7830 1032
rect 0 -32 36 0
rect 270 -32 306 0
rect 836 -32 872 0
rect 1106 -32 1142 0
rect 1672 -32 1708 0
rect 1942 -32 1978 0
rect 2508 -32 2544 0
rect 2778 -32 2814 0
rect 3344 -32 3380 0
rect 3614 -32 3650 0
rect 4180 -32 4216 0
rect 4450 -32 4486 0
rect 5016 -32 5052 0
rect 5286 -32 5322 0
rect 5852 -32 5888 0
rect 6122 -32 6158 0
rect 6688 -32 6724 0
rect 6958 -32 6994 0
rect 7524 -32 7560 0
rect 7794 -32 7830 0
<< locali >>
rect -354 -4 -176 946
rect 482 -4 660 946
rect 1318 -4 1496 946
rect 2154 -4 2332 946
rect 2990 -4 3168 946
rect 3826 -4 4004 946
rect 4662 -4 4840 946
rect 5498 -4 5676 946
rect 6334 -4 6512 946
rect 7170 -4 7348 946
rect 8006 -4 8184 946
use DFTPL1s2_CDNS_55959141808694  DFTPL1s2_CDNS_55959141808694_0
timestamp 1701704242
transform -1 0 -165 0 1 0
box -26 -26 226 1026
use DFTPL1s2_CDNS_55959141808694  DFTPL1s2_CDNS_55959141808694_1
timestamp 1701704242
transform 1 0 471 0 1 0
box -26 -26 226 1026
use DFTPL1s2_CDNS_55959141808694  DFTPL1s2_CDNS_55959141808694_2
timestamp 1701704242
transform 1 0 1307 0 1 0
box -26 -26 226 1026
use DFTPL1s2_CDNS_55959141808694  DFTPL1s2_CDNS_55959141808694_3
timestamp 1701704242
transform 1 0 2143 0 1 0
box -26 -26 226 1026
use DFTPL1s2_CDNS_55959141808694  DFTPL1s2_CDNS_55959141808694_4
timestamp 1701704242
transform 1 0 2979 0 1 0
box -26 -26 226 1026
use DFTPL1s2_CDNS_55959141808694  DFTPL1s2_CDNS_55959141808694_5
timestamp 1701704242
transform 1 0 3815 0 1 0
box -26 -26 226 1026
use DFTPL1s2_CDNS_55959141808694  DFTPL1s2_CDNS_55959141808694_6
timestamp 1701704242
transform 1 0 4651 0 1 0
box -26 -26 226 1026
use DFTPL1s2_CDNS_55959141808694  DFTPL1s2_CDNS_55959141808694_7
timestamp 1701704242
transform 1 0 5487 0 1 0
box -26 -26 226 1026
use DFTPL1s2_CDNS_55959141808694  DFTPL1s2_CDNS_55959141808694_8
timestamp 1701704242
transform 1 0 6323 0 1 0
box -26 -26 226 1026
use DFTPL1s2_CDNS_55959141808694  DFTPL1s2_CDNS_55959141808694_9
timestamp 1701704242
transform 1 0 7159 0 1 0
box -26 -26 226 1026
use DFTPL1s2_CDNS_55959141808694  DFTPL1s2_CDNS_55959141808694_10
timestamp 1701704242
transform 1 0 7995 0 1 0
box -26 -26 226 1026
<< labels >>
flabel comment s 8095 471 8095 471 0 FreeSans 300 0 0 0 S
flabel comment s 7677 500 7677 500 0 FreeSans 300 0 0 0 D
flabel comment s 7259 471 7259 471 0 FreeSans 300 0 0 0 S
flabel comment s 6841 500 6841 500 0 FreeSans 300 0 0 0 D
flabel comment s 6423 471 6423 471 0 FreeSans 300 0 0 0 S
flabel comment s 6005 500 6005 500 0 FreeSans 300 0 0 0 D
flabel comment s 5587 471 5587 471 0 FreeSans 300 0 0 0 S
flabel comment s 5169 500 5169 500 0 FreeSans 300 0 0 0 D
flabel comment s 4751 471 4751 471 0 FreeSans 300 0 0 0 S
flabel comment s 4333 500 4333 500 0 FreeSans 300 0 0 0 D
flabel comment s 3915 471 3915 471 0 FreeSans 300 0 0 0 S
flabel comment s 3497 500 3497 500 0 FreeSans 300 0 0 0 D
flabel comment s 3079 471 3079 471 0 FreeSans 300 0 0 0 S
flabel comment s 2661 500 2661 500 0 FreeSans 300 0 0 0 D
flabel comment s 2243 471 2243 471 0 FreeSans 300 0 0 0 S
flabel comment s 1825 500 1825 500 0 FreeSans 300 0 0 0 D
flabel comment s 1407 471 1407 471 0 FreeSans 300 0 0 0 S
flabel comment s 989 500 989 500 0 FreeSans 300 0 0 0 D
flabel comment s 571 471 571 471 0 FreeSans 300 0 0 0 S
flabel comment s 153 500 153 500 0 FreeSans 300 0 0 0 D
flabel comment s -265 471 -265 471 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 43008856
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 42998448
<< end >>
