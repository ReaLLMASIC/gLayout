magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< locali >>
rect 513 11329 547 11345
rect 1873 11329 1907 11345
rect 0 11295 513 11329
rect 547 11295 1873 11329
rect 1907 11295 2826 11329
rect 513 11279 547 11295
rect 1873 11279 1907 11295
rect 121 11059 155 11075
rect 1481 11059 1515 11075
rect 155 11025 1481 11059
rect 1515 11025 2093 11059
rect 121 11009 155 11025
rect 1481 11009 1515 11025
rect 245 10935 279 10951
rect 1605 10935 1639 10951
rect 279 10901 1605 10935
rect 1639 10901 2226 10935
rect 245 10885 279 10901
rect 1605 10885 1639 10901
rect 369 10811 403 10827
rect 1729 10811 1763 10827
rect 403 10777 1729 10811
rect 1763 10777 2359 10811
rect 369 10761 403 10777
rect 1729 10761 1763 10777
rect 2637 10626 2671 10660
rect 513 9915 547 9931
rect 1873 9915 1907 9931
rect 0 9881 513 9915
rect 547 9881 1873 9915
rect 1907 9881 2826 9915
rect 513 9865 547 9881
rect 1873 9865 1907 9881
rect 2637 9136 2671 9170
rect 1713 8985 1729 9019
rect 1763 8985 2359 9019
rect 1589 8861 1605 8895
rect 1639 8861 2226 8895
rect 1093 8737 1109 8771
rect 1143 8737 2093 8771
rect 513 8501 547 8517
rect 1873 8501 1907 8517
rect 0 8467 513 8501
rect 547 8467 1873 8501
rect 1907 8467 2826 8501
rect 513 8451 547 8467
rect 1873 8451 1907 8467
rect 1465 8197 1481 8231
rect 1515 8197 2093 8231
rect 1217 8073 1233 8107
rect 1267 8073 2226 8107
rect 1713 7949 1729 7983
rect 1763 7949 2359 7983
rect 2637 7798 2671 7832
rect 513 7087 547 7103
rect 1873 7087 1907 7103
rect 0 7053 513 7087
rect 547 7053 1873 7087
rect 1907 7053 2826 7087
rect 513 7037 547 7053
rect 1873 7037 1907 7053
rect 2637 6308 2671 6342
rect 1713 6157 1729 6191
rect 1763 6157 2359 6191
rect 1217 6033 1233 6067
rect 1267 6033 2226 6067
rect 1093 5909 1109 5943
rect 1143 5909 2093 5943
rect 513 5673 547 5689
rect 1873 5673 1907 5689
rect 0 5639 513 5673
rect 547 5639 1873 5673
rect 1907 5639 2826 5673
rect 513 5623 547 5639
rect 1873 5623 1907 5639
rect 1465 5369 1481 5403
rect 1515 5369 2093 5403
rect 1589 5245 1605 5279
rect 1639 5245 2226 5279
rect 1341 5121 1357 5155
rect 1391 5121 2359 5155
rect 2637 4970 2671 5004
rect 513 4259 547 4275
rect 1873 4259 1907 4275
rect 0 4225 513 4259
rect 547 4225 1873 4259
rect 1907 4225 2826 4259
rect 513 4209 547 4225
rect 1873 4209 1907 4225
rect 816 3514 850 3530
rect 353 3480 369 3514
rect 403 3480 718 3514
rect 2637 3480 2671 3514
rect 816 3464 850 3480
rect 1341 3329 1357 3363
rect 1391 3329 2359 3363
rect 1589 3205 1605 3239
rect 1639 3205 2226 3239
rect 1093 3081 1109 3115
rect 1143 3081 2093 3115
rect 513 2845 547 2861
rect 1873 2845 1907 2861
rect 0 2811 513 2845
rect 547 2811 1873 2845
rect 1907 2811 2826 2845
rect 513 2795 547 2811
rect 1873 2795 1907 2811
rect 1465 2541 1481 2575
rect 1515 2541 2093 2575
rect 1217 2417 1233 2451
rect 1267 2417 2226 2451
rect 1341 2293 1357 2327
rect 1391 2293 2359 2327
rect 816 2176 850 2192
rect 229 2142 245 2176
rect 279 2142 718 2176
rect 2637 2142 2671 2176
rect 816 2126 850 2142
rect 513 1431 547 1447
rect 1873 1431 1907 1447
rect 0 1397 513 1431
rect 547 1397 1873 1431
rect 1907 1397 2826 1431
rect 513 1381 547 1397
rect 1873 1381 1907 1397
rect 816 686 850 702
rect 105 652 121 686
rect 155 652 718 686
rect 2637 652 2671 686
rect 816 636 850 652
rect 1341 501 1357 535
rect 1391 501 2359 535
rect 1217 377 1233 411
rect 1267 377 2226 411
rect 1093 253 1109 287
rect 1143 253 2093 287
rect 513 17 547 33
rect 1873 17 1907 33
rect 0 -17 513 17
rect 547 -17 1873 17
rect 1907 -17 2826 17
rect 513 -33 547 -17
rect 1873 -33 1907 -17
<< viali >>
rect 513 11295 547 11329
rect 1873 11295 1907 11329
rect 121 11025 155 11059
rect 1481 11025 1515 11059
rect 245 10901 279 10935
rect 1605 10901 1639 10935
rect 369 10777 403 10811
rect 1729 10777 1763 10811
rect 513 9881 547 9915
rect 1873 9881 1907 9915
rect 1729 8985 1763 9019
rect 1605 8861 1639 8895
rect 1109 8737 1143 8771
rect 513 8467 547 8501
rect 1873 8467 1907 8501
rect 1481 8197 1515 8231
rect 1233 8073 1267 8107
rect 1729 7949 1763 7983
rect 513 7053 547 7087
rect 1873 7053 1907 7087
rect 1729 6157 1763 6191
rect 1233 6033 1267 6067
rect 1109 5909 1143 5943
rect 513 5639 547 5673
rect 1873 5639 1907 5673
rect 1481 5369 1515 5403
rect 1605 5245 1639 5279
rect 1357 5121 1391 5155
rect 513 4225 547 4259
rect 1873 4225 1907 4259
rect 369 3480 403 3514
rect 816 3480 850 3514
rect 1357 3329 1391 3363
rect 1605 3205 1639 3239
rect 1109 3081 1143 3115
rect 513 2811 547 2845
rect 1873 2811 1907 2845
rect 1481 2541 1515 2575
rect 1233 2417 1267 2451
rect 1357 2293 1391 2327
rect 245 2142 279 2176
rect 816 2142 850 2176
rect 513 1397 547 1431
rect 1873 1397 1907 1431
rect 121 652 155 686
rect 816 652 850 686
rect 1357 501 1391 535
rect 1233 377 1267 411
rect 1109 253 1143 287
rect 513 -17 547 17
rect 1873 -17 1907 17
<< metal1 >>
rect 498 11286 504 11338
rect 556 11286 562 11338
rect 1858 11286 1864 11338
rect 1916 11286 1922 11338
rect 124 11065 152 11188
rect 109 11059 167 11065
rect 109 11025 121 11059
rect 155 11025 167 11059
rect 109 11019 167 11025
rect 124 698 152 11019
rect 248 10941 276 11188
rect 233 10935 291 10941
rect 233 10901 245 10935
rect 279 10901 291 10935
rect 233 10895 291 10901
rect 248 2188 276 10895
rect 372 10817 400 11188
rect 357 10811 415 10817
rect 357 10777 369 10811
rect 403 10777 415 10811
rect 357 10771 415 10777
rect 372 3526 400 10771
rect 498 9872 504 9924
rect 556 9872 562 9924
rect 1112 8783 1140 11188
rect 1103 8771 1149 8783
rect 1103 8737 1109 8771
rect 1143 8737 1149 8771
rect 1103 8725 1149 8737
rect 498 8458 504 8510
rect 556 8458 562 8510
rect 498 7044 504 7096
rect 556 7044 562 7096
rect 1112 5955 1140 8725
rect 1236 8119 1264 11188
rect 1227 8107 1273 8119
rect 1227 8073 1233 8107
rect 1267 8073 1273 8107
rect 1227 8061 1273 8073
rect 1236 6079 1264 8061
rect 1227 6067 1273 6079
rect 1227 6033 1233 6067
rect 1267 6033 1273 6067
rect 1227 6021 1273 6033
rect 1103 5943 1149 5955
rect 1103 5909 1109 5943
rect 1143 5909 1149 5943
rect 1103 5897 1149 5909
rect 498 5630 504 5682
rect 556 5630 562 5682
rect 498 4216 504 4268
rect 556 4216 562 4268
rect 363 3514 409 3526
rect 363 3480 369 3514
rect 403 3480 409 3514
rect 363 3468 409 3480
rect 801 3471 807 3523
rect 859 3471 865 3523
rect 239 2176 285 2188
rect 239 2142 245 2176
rect 279 2142 285 2176
rect 239 2130 285 2142
rect 115 686 161 698
rect 115 652 121 686
rect 155 652 161 686
rect 115 640 161 652
rect 124 124 152 640
rect 248 124 276 2130
rect 372 124 400 3468
rect 1112 3127 1140 5897
rect 1103 3115 1149 3127
rect 1103 3081 1109 3115
rect 1143 3081 1149 3115
rect 1103 3069 1149 3081
rect 498 2802 504 2854
rect 556 2802 562 2854
rect 801 2133 807 2185
rect 859 2133 865 2185
rect 498 1388 504 1440
rect 556 1388 562 1440
rect 1112 1362 1140 3069
rect 1236 2776 1264 6021
rect 1360 5167 1388 11188
rect 1484 11071 1512 11188
rect 1475 11065 1521 11071
rect 1469 11059 1527 11065
rect 1469 11025 1481 11059
rect 1515 11025 1527 11059
rect 1469 11019 1527 11025
rect 1475 11013 1521 11019
rect 1484 8243 1512 11013
rect 1608 10947 1636 11188
rect 1599 10941 1645 10947
rect 1593 10935 1651 10941
rect 1593 10901 1605 10935
rect 1639 10901 1651 10935
rect 1593 10895 1651 10901
rect 1599 10889 1645 10895
rect 1608 8907 1636 10889
rect 1732 10823 1760 11188
rect 1723 10817 1769 10823
rect 1717 10811 1775 10817
rect 1717 10777 1729 10811
rect 1763 10777 1775 10811
rect 1717 10771 1775 10777
rect 1723 10765 1769 10771
rect 1732 9031 1760 10765
rect 1858 9872 1864 9924
rect 1916 9872 1922 9924
rect 1723 9019 1769 9031
rect 1723 8985 1729 9019
rect 1763 8985 1769 9019
rect 1723 8973 1769 8985
rect 1599 8895 1645 8907
rect 1599 8861 1605 8895
rect 1639 8861 1645 8895
rect 1599 8849 1645 8861
rect 1475 8231 1521 8243
rect 1475 8197 1481 8231
rect 1515 8197 1521 8231
rect 1475 8185 1521 8197
rect 1484 5415 1512 8185
rect 1475 5403 1521 5415
rect 1475 5369 1481 5403
rect 1515 5369 1521 5403
rect 1475 5357 1521 5369
rect 1351 5155 1397 5167
rect 1351 5121 1357 5155
rect 1391 5121 1397 5155
rect 1351 5109 1397 5121
rect 1360 4190 1388 5109
rect 1348 4184 1400 4190
rect 1348 4126 1400 4132
rect 1360 3375 1388 4126
rect 1351 3363 1397 3375
rect 1351 3329 1357 3363
rect 1391 3329 1397 3363
rect 1351 3317 1397 3329
rect 1224 2770 1276 2776
rect 1224 2712 1276 2718
rect 1236 2463 1264 2712
rect 1227 2451 1273 2463
rect 1227 2417 1233 2451
rect 1267 2417 1273 2451
rect 1227 2405 1273 2417
rect 1100 1356 1152 1362
rect 1100 1298 1152 1304
rect 801 643 807 695
rect 859 643 865 695
rect 1112 299 1140 1298
rect 1236 423 1264 2405
rect 1360 2339 1388 3317
rect 1484 2587 1512 5357
rect 1608 5291 1636 8849
rect 1732 7995 1760 8973
rect 1858 8458 1864 8510
rect 1916 8458 1922 8510
rect 1723 7983 1769 7995
rect 1723 7949 1729 7983
rect 1763 7949 1769 7983
rect 1723 7937 1769 7949
rect 1732 6203 1760 7937
rect 1858 7044 1864 7096
rect 1916 7044 1922 7096
rect 1723 6191 1769 6203
rect 1723 6157 1729 6191
rect 1763 6157 1769 6191
rect 1723 6145 1769 6157
rect 1599 5279 1645 5291
rect 1599 5245 1605 5279
rect 1639 5245 1645 5279
rect 1599 5233 1645 5245
rect 1608 3251 1636 5233
rect 1599 3239 1645 3251
rect 1599 3205 1605 3239
rect 1639 3205 1645 3239
rect 1599 3193 1645 3205
rect 1475 2575 1521 2587
rect 1475 2541 1481 2575
rect 1515 2541 1521 2575
rect 1475 2529 1521 2541
rect 1351 2327 1397 2339
rect 1351 2293 1357 2327
rect 1391 2293 1397 2327
rect 1351 2281 1397 2293
rect 1360 547 1388 2281
rect 1351 535 1397 547
rect 1351 501 1357 535
rect 1391 501 1397 535
rect 1351 489 1397 501
rect 1227 411 1273 423
rect 1227 377 1233 411
rect 1267 377 1273 411
rect 1227 365 1273 377
rect 1103 287 1149 299
rect 1103 253 1109 287
rect 1143 253 1149 287
rect 1103 241 1149 253
rect 1112 124 1140 241
rect 1236 124 1264 365
rect 1360 124 1388 489
rect 1484 124 1512 2529
rect 1608 124 1636 3193
rect 1732 124 1760 6145
rect 1858 5630 1864 5682
rect 1916 5630 1922 5682
rect 1858 4216 1864 4268
rect 1916 4216 1922 4268
rect 1858 2802 1864 2854
rect 1916 2802 1922 2854
rect 1858 1388 1864 1440
rect 1916 1388 1922 1440
rect 498 -26 504 26
rect 556 -26 562 26
rect 1858 -26 1864 26
rect 1916 -26 1922 26
<< via1 >>
rect 504 11329 556 11338
rect 504 11295 513 11329
rect 513 11295 547 11329
rect 547 11295 556 11329
rect 504 11286 556 11295
rect 1864 11329 1916 11338
rect 1864 11295 1873 11329
rect 1873 11295 1907 11329
rect 1907 11295 1916 11329
rect 1864 11286 1916 11295
rect 504 9915 556 9924
rect 504 9881 513 9915
rect 513 9881 547 9915
rect 547 9881 556 9915
rect 504 9872 556 9881
rect 504 8501 556 8510
rect 504 8467 513 8501
rect 513 8467 547 8501
rect 547 8467 556 8501
rect 504 8458 556 8467
rect 504 7087 556 7096
rect 504 7053 513 7087
rect 513 7053 547 7087
rect 547 7053 556 7087
rect 504 7044 556 7053
rect 504 5673 556 5682
rect 504 5639 513 5673
rect 513 5639 547 5673
rect 547 5639 556 5673
rect 504 5630 556 5639
rect 504 4259 556 4268
rect 504 4225 513 4259
rect 513 4225 547 4259
rect 547 4225 556 4259
rect 504 4216 556 4225
rect 807 3514 859 3523
rect 807 3480 816 3514
rect 816 3480 850 3514
rect 850 3480 859 3514
rect 807 3471 859 3480
rect 504 2845 556 2854
rect 504 2811 513 2845
rect 513 2811 547 2845
rect 547 2811 556 2845
rect 504 2802 556 2811
rect 807 2176 859 2185
rect 807 2142 816 2176
rect 816 2142 850 2176
rect 850 2142 859 2176
rect 807 2133 859 2142
rect 504 1431 556 1440
rect 504 1397 513 1431
rect 513 1397 547 1431
rect 547 1397 556 1431
rect 504 1388 556 1397
rect 1864 9915 1916 9924
rect 1864 9881 1873 9915
rect 1873 9881 1907 9915
rect 1907 9881 1916 9915
rect 1864 9872 1916 9881
rect 1348 4132 1400 4184
rect 1224 2718 1276 2770
rect 1100 1304 1152 1356
rect 807 686 859 695
rect 807 652 816 686
rect 816 652 850 686
rect 850 652 859 686
rect 807 643 859 652
rect 1864 8501 1916 8510
rect 1864 8467 1873 8501
rect 1873 8467 1907 8501
rect 1907 8467 1916 8501
rect 1864 8458 1916 8467
rect 1864 7087 1916 7096
rect 1864 7053 1873 7087
rect 1873 7053 1907 7087
rect 1907 7053 1916 7087
rect 1864 7044 1916 7053
rect 1864 5673 1916 5682
rect 1864 5639 1873 5673
rect 1873 5639 1907 5673
rect 1907 5639 1916 5673
rect 1864 5630 1916 5639
rect 1864 4259 1916 4268
rect 1864 4225 1873 4259
rect 1873 4225 1907 4259
rect 1907 4225 1916 4259
rect 1864 4216 1916 4225
rect 1864 2845 1916 2854
rect 1864 2811 1873 2845
rect 1873 2811 1907 2845
rect 1907 2811 1916 2845
rect 1864 2802 1916 2811
rect 1864 1431 1916 1440
rect 1864 1397 1873 1431
rect 1873 1397 1907 1431
rect 1907 1397 1916 1431
rect 1864 1388 1916 1397
rect 504 17 556 26
rect 504 -17 513 17
rect 513 -17 547 17
rect 547 -17 556 17
rect 504 -26 556 -17
rect 1864 17 1916 26
rect 1864 -17 1873 17
rect 1873 -17 1907 17
rect 1907 -17 1916 17
rect 1864 -26 1916 -17
<< metal2 >>
rect 502 11340 558 11349
rect 502 11275 558 11284
rect 1862 11340 1918 11349
rect 1862 11275 1918 11284
rect 502 9926 558 9935
rect 502 9861 558 9870
rect 1862 9926 1918 9935
rect 1862 9861 1918 9870
rect 502 8512 558 8521
rect 502 8447 558 8456
rect 1862 8512 1918 8521
rect 1862 8447 1918 8456
rect 502 7098 558 7107
rect 502 7033 558 7042
rect 1862 7098 1918 7107
rect 1862 7033 1918 7042
rect 502 5684 558 5693
rect 502 5619 558 5628
rect 1862 5684 1918 5693
rect 1862 5619 1918 5628
rect 502 4270 558 4279
rect 502 4205 558 4214
rect 1862 4270 1918 4279
rect 1862 4205 1918 4214
rect 1342 4172 1348 4184
rect 974 4144 1348 4172
rect 807 3523 859 3529
rect 974 3511 1002 4144
rect 1342 4132 1348 4144
rect 1400 4132 1406 4184
rect 859 3483 1002 3511
rect 807 3465 859 3471
rect 502 2856 558 2865
rect 502 2791 558 2800
rect 1862 2856 1918 2865
rect 1862 2791 1918 2800
rect 1218 2758 1224 2770
rect 974 2730 1224 2758
rect 807 2185 859 2191
rect 974 2173 1002 2730
rect 1218 2718 1224 2730
rect 1276 2718 1282 2770
rect 859 2145 1002 2173
rect 807 2127 859 2133
rect 502 1442 558 1451
rect 502 1377 558 1386
rect 1862 1442 1918 1451
rect 1862 1377 1918 1386
rect 1094 1344 1100 1356
rect 974 1316 1100 1344
rect 807 695 859 701
rect 974 683 1002 1316
rect 1094 1304 1100 1316
rect 1152 1304 1158 1356
rect 859 655 1002 683
rect 807 637 859 643
rect 502 28 558 37
rect 502 -37 558 -28
rect 1862 28 1918 37
rect 1862 -37 1918 -28
<< via2 >>
rect 502 11338 558 11340
rect 502 11286 504 11338
rect 504 11286 556 11338
rect 556 11286 558 11338
rect 502 11284 558 11286
rect 1862 11338 1918 11340
rect 1862 11286 1864 11338
rect 1864 11286 1916 11338
rect 1916 11286 1918 11338
rect 1862 11284 1918 11286
rect 502 9924 558 9926
rect 502 9872 504 9924
rect 504 9872 556 9924
rect 556 9872 558 9924
rect 502 9870 558 9872
rect 1862 9924 1918 9926
rect 1862 9872 1864 9924
rect 1864 9872 1916 9924
rect 1916 9872 1918 9924
rect 1862 9870 1918 9872
rect 502 8510 558 8512
rect 502 8458 504 8510
rect 504 8458 556 8510
rect 556 8458 558 8510
rect 502 8456 558 8458
rect 1862 8510 1918 8512
rect 1862 8458 1864 8510
rect 1864 8458 1916 8510
rect 1916 8458 1918 8510
rect 1862 8456 1918 8458
rect 502 7096 558 7098
rect 502 7044 504 7096
rect 504 7044 556 7096
rect 556 7044 558 7096
rect 502 7042 558 7044
rect 1862 7096 1918 7098
rect 1862 7044 1864 7096
rect 1864 7044 1916 7096
rect 1916 7044 1918 7096
rect 1862 7042 1918 7044
rect 502 5682 558 5684
rect 502 5630 504 5682
rect 504 5630 556 5682
rect 556 5630 558 5682
rect 502 5628 558 5630
rect 1862 5682 1918 5684
rect 1862 5630 1864 5682
rect 1864 5630 1916 5682
rect 1916 5630 1918 5682
rect 1862 5628 1918 5630
rect 502 4268 558 4270
rect 502 4216 504 4268
rect 504 4216 556 4268
rect 556 4216 558 4268
rect 502 4214 558 4216
rect 1862 4268 1918 4270
rect 1862 4216 1864 4268
rect 1864 4216 1916 4268
rect 1916 4216 1918 4268
rect 1862 4214 1918 4216
rect 502 2854 558 2856
rect 502 2802 504 2854
rect 504 2802 556 2854
rect 556 2802 558 2854
rect 502 2800 558 2802
rect 1862 2854 1918 2856
rect 1862 2802 1864 2854
rect 1864 2802 1916 2854
rect 1916 2802 1918 2854
rect 1862 2800 1918 2802
rect 502 1440 558 1442
rect 502 1388 504 1440
rect 504 1388 556 1440
rect 556 1388 558 1440
rect 502 1386 558 1388
rect 1862 1440 1918 1442
rect 1862 1388 1864 1440
rect 1864 1388 1916 1440
rect 1916 1388 1918 1440
rect 1862 1386 1918 1388
rect 502 26 558 28
rect 502 -26 504 26
rect 504 -26 556 26
rect 556 -26 558 26
rect 502 -28 558 -26
rect 1862 26 1918 28
rect 1862 -26 1864 26
rect 1864 -26 1916 26
rect 1916 -26 1918 26
rect 1862 -28 1918 -26
<< metal3 >>
rect 481 11340 579 11361
rect 481 11284 502 11340
rect 558 11284 579 11340
rect 481 11263 579 11284
rect 1841 11340 1939 11361
rect 1841 11284 1862 11340
rect 1918 11284 1939 11340
rect 1841 11263 1939 11284
rect 481 9926 579 9947
rect 481 9870 502 9926
rect 558 9870 579 9926
rect 481 9849 579 9870
rect 1841 9926 1939 9947
rect 1841 9870 1862 9926
rect 1918 9870 1939 9926
rect 1841 9849 1939 9870
rect 481 8512 579 8533
rect 481 8456 502 8512
rect 558 8456 579 8512
rect 481 8435 579 8456
rect 1841 8512 1939 8533
rect 1841 8456 1862 8512
rect 1918 8456 1939 8512
rect 1841 8435 1939 8456
rect 481 7098 579 7119
rect 481 7042 502 7098
rect 558 7042 579 7098
rect 481 7021 579 7042
rect 1841 7098 1939 7119
rect 1841 7042 1862 7098
rect 1918 7042 1939 7098
rect 1841 7021 1939 7042
rect 481 5684 579 5705
rect 481 5628 502 5684
rect 558 5628 579 5684
rect 481 5607 579 5628
rect 1841 5684 1939 5705
rect 1841 5628 1862 5684
rect 1918 5628 1939 5684
rect 1841 5607 1939 5628
rect 481 4270 579 4291
rect 481 4214 502 4270
rect 558 4214 579 4270
rect 481 4193 579 4214
rect 1841 4270 1939 4291
rect 1841 4214 1862 4270
rect 1918 4214 1939 4270
rect 1841 4193 1939 4214
rect 481 2856 579 2877
rect 481 2800 502 2856
rect 558 2800 579 2856
rect 481 2779 579 2800
rect 1841 2856 1939 2877
rect 1841 2800 1862 2856
rect 1918 2800 1939 2856
rect 1841 2779 1939 2800
rect 481 1442 579 1463
rect 481 1386 502 1442
rect 558 1386 579 1442
rect 481 1365 579 1386
rect 1841 1442 1939 1463
rect 1841 1386 1862 1442
rect 1918 1386 1939 1442
rect 1841 1365 1939 1386
rect 481 28 579 49
rect 481 -28 502 28
rect 558 -28 579 28
rect 481 -49 579 -28
rect 1841 28 1939 49
rect 1841 -28 1862 28
rect 1918 -28 1939 28
rect 1841 -49 1939 -28
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_0
timestamp 1701704242
transform 1 0 1857 0 1 -37
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_1
timestamp 1701704242
transform 1 0 497 0 1 -37
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_2
timestamp 1701704242
transform 1 0 1857 0 1 1377
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_3
timestamp 1701704242
transform 1 0 497 0 1 1377
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_4
timestamp 1701704242
transform 1 0 1857 0 1 2791
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_5
timestamp 1701704242
transform 1 0 497 0 1 2791
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_6
timestamp 1701704242
transform 1 0 1857 0 1 4205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_7
timestamp 1701704242
transform 1 0 497 0 1 4205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_8
timestamp 1701704242
transform 1 0 1857 0 1 11275
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_9
timestamp 1701704242
transform 1 0 497 0 1 11275
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_10
timestamp 1701704242
transform 1 0 1857 0 1 9861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_11
timestamp 1701704242
transform 1 0 497 0 1 9861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_12
timestamp 1701704242
transform 1 0 1857 0 1 8447
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_13
timestamp 1701704242
transform 1 0 497 0 1 8447
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_14
timestamp 1701704242
transform 1 0 1857 0 1 7033
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_15
timestamp 1701704242
transform 1 0 497 0 1 7033
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_16
timestamp 1701704242
transform 1 0 1857 0 1 5619
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_17
timestamp 1701704242
transform 1 0 497 0 1 5619
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_0
timestamp 1701704242
transform 1 0 1861 0 1 -33
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_1
timestamp 1701704242
transform 1 0 501 0 1 -33
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_2
timestamp 1701704242
transform 1 0 1861 0 1 1381
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_3
timestamp 1701704242
transform 1 0 501 0 1 1381
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_4
timestamp 1701704242
transform 1 0 804 0 1 3464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_5
timestamp 1701704242
transform 1 0 804 0 1 2126
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_6
timestamp 1701704242
transform 1 0 804 0 1 636
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_7
timestamp 1701704242
transform 1 0 1861 0 1 2795
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_8
timestamp 1701704242
transform 1 0 501 0 1 2795
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_9
timestamp 1701704242
transform 1 0 1861 0 1 4209
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_10
timestamp 1701704242
transform 1 0 501 0 1 4209
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_11
timestamp 1701704242
transform 1 0 1861 0 1 11279
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_12
timestamp 1701704242
transform 1 0 501 0 1 11279
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_13
timestamp 1701704242
transform 1 0 1861 0 1 9865
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_14
timestamp 1701704242
transform 1 0 501 0 1 9865
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_15
timestamp 1701704242
transform 1 0 1861 0 1 8451
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_16
timestamp 1701704242
transform 1 0 501 0 1 8451
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_17
timestamp 1701704242
transform 1 0 1861 0 1 7037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_18
timestamp 1701704242
transform 1 0 501 0 1 7037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_19
timestamp 1701704242
transform 1 0 1717 0 1 10761
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_20
timestamp 1701704242
transform 1 0 357 0 1 10761
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_21
timestamp 1701704242
transform 1 0 1593 0 1 10885
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_22
timestamp 1701704242
transform 1 0 233 0 1 10885
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_23
timestamp 1701704242
transform 1 0 1469 0 1 11009
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_24
timestamp 1701704242
transform 1 0 109 0 1 11009
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_25
timestamp 1701704242
transform 1 0 1861 0 1 5623
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_26
timestamp 1701704242
transform 1 0 501 0 1 5623
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17_0
timestamp 1701704242
transform 1 0 1341 0 1 3317
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17_1
timestamp 1701704242
transform 1 0 1589 0 1 3193
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17_2
timestamp 1701704242
transform 1 0 1093 0 1 3069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17_3
timestamp 1701704242
transform 1 0 1341 0 1 2281
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17_4
timestamp 1701704242
transform 1 0 1217 0 1 2405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17_5
timestamp 1701704242
transform 1 0 1465 0 1 2529
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17_6
timestamp 1701704242
transform 1 0 1341 0 1 489
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17_7
timestamp 1701704242
transform 1 0 1217 0 1 365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17_8
timestamp 1701704242
transform 1 0 1093 0 1 241
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17_9
timestamp 1701704242
transform 1 0 353 0 1 3468
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17_10
timestamp 1701704242
transform 1 0 229 0 1 2130
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17_11
timestamp 1701704242
transform 1 0 105 0 1 640
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17_12
timestamp 1701704242
transform 1 0 1341 0 1 5109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17_13
timestamp 1701704242
transform 1 0 1589 0 1 5233
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17_14
timestamp 1701704242
transform 1 0 1465 0 1 5357
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17_15
timestamp 1701704242
transform 1 0 1713 0 1 8973
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17_16
timestamp 1701704242
transform 1 0 1589 0 1 8849
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17_17
timestamp 1701704242
transform 1 0 1093 0 1 8725
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17_18
timestamp 1701704242
transform 1 0 1713 0 1 7937
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17_19
timestamp 1701704242
transform 1 0 1217 0 1 8061
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17_20
timestamp 1701704242
transform 1 0 1465 0 1 8185
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17_21
timestamp 1701704242
transform 1 0 1713 0 1 6145
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17_22
timestamp 1701704242
transform 1 0 1217 0 1 6021
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17_23
timestamp 1701704242
transform 1 0 1093 0 1 5897
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17_24
timestamp 1701704242
transform 1 0 1713 0 1 10765
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17_25
timestamp 1701704242
transform 1 0 1589 0 1 10889
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_17_26
timestamp 1701704242
transform 1 0 1465 0 1 11013
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_0
timestamp 1701704242
transform 1 0 1858 0 1 -32
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_1
timestamp 1701704242
transform 1 0 498 0 1 -32
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_2
timestamp 1701704242
transform 1 0 1858 0 1 1382
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_3
timestamp 1701704242
transform 1 0 498 0 1 1382
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_4
timestamp 1701704242
transform 1 0 801 0 1 3465
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_5
timestamp 1701704242
transform 1 0 801 0 1 2127
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_6
timestamp 1701704242
transform 1 0 801 0 1 637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_7
timestamp 1701704242
transform 1 0 1858 0 1 2796
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_8
timestamp 1701704242
transform 1 0 498 0 1 2796
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_9
timestamp 1701704242
transform 1 0 1858 0 1 4210
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_10
timestamp 1701704242
transform 1 0 498 0 1 4210
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_11
timestamp 1701704242
transform 1 0 1858 0 1 11280
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_12
timestamp 1701704242
transform 1 0 498 0 1 11280
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_13
timestamp 1701704242
transform 1 0 1858 0 1 9866
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_14
timestamp 1701704242
transform 1 0 498 0 1 9866
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_15
timestamp 1701704242
transform 1 0 1858 0 1 8452
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_16
timestamp 1701704242
transform 1 0 498 0 1 8452
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_17
timestamp 1701704242
transform 1 0 1858 0 1 7038
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_18
timestamp 1701704242
transform 1 0 498 0 1 7038
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_19
timestamp 1701704242
transform 1 0 1858 0 1 5624
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_20
timestamp 1701704242
transform 1 0 498 0 1 5624
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_20  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_20_0
timestamp 1701704242
transform 1 0 1342 0 1 4126
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_20  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_20_1
timestamp 1701704242
transform 1 0 1218 0 1 2712
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_20  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_20_2
timestamp 1701704242
transform 1 0 1094 0 1 1298
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_pand3  sky130_sram_1kbyte_1rw1r_8x1024_8_pand3_0
timestamp 1701704242
transform 1 0 1980 0 -1 2828
box -36 -17 882 1471
use sky130_sram_1kbyte_1rw1r_8x1024_8_pand3  sky130_sram_1kbyte_1rw1r_8x1024_8_pand3_1
timestamp 1701704242
transform 1 0 1980 0 1 0
box -36 -17 882 1471
use sky130_sram_1kbyte_1rw1r_8x1024_8_pand3  sky130_sram_1kbyte_1rw1r_8x1024_8_pand3_2
timestamp 1701704242
transform 1 0 1980 0 1 2828
box -36 -17 882 1471
use sky130_sram_1kbyte_1rw1r_8x1024_8_pand3  sky130_sram_1kbyte_1rw1r_8x1024_8_pand3_3
timestamp 1701704242
transform 1 0 1980 0 -1 11312
box -36 -17 882 1471
use sky130_sram_1kbyte_1rw1r_8x1024_8_pand3  sky130_sram_1kbyte_1rw1r_8x1024_8_pand3_4
timestamp 1701704242
transform 1 0 1980 0 1 8484
box -36 -17 882 1471
use sky130_sram_1kbyte_1rw1r_8x1024_8_pand3  sky130_sram_1kbyte_1rw1r_8x1024_8_pand3_5
timestamp 1701704242
transform 1 0 1980 0 -1 8484
box -36 -17 882 1471
use sky130_sram_1kbyte_1rw1r_8x1024_8_pand3  sky130_sram_1kbyte_1rw1r_8x1024_8_pand3_6
timestamp 1701704242
transform 1 0 1980 0 1 5656
box -36 -17 882 1471
use sky130_sram_1kbyte_1rw1r_8x1024_8_pand3  sky130_sram_1kbyte_1rw1r_8x1024_8_pand3_7
timestamp 1701704242
transform 1 0 1980 0 -1 5656
box -36 -17 882 1471
use sky130_sram_1kbyte_1rw1r_8x1024_8_pinv_1  sky130_sram_1kbyte_1rw1r_8x1024_8_pinv_1_0
timestamp 1701704242
transform 1 0 620 0 1 2828
box -36 -17 404 1471
use sky130_sram_1kbyte_1rw1r_8x1024_8_pinv_1  sky130_sram_1kbyte_1rw1r_8x1024_8_pinv_1_1
timestamp 1701704242
transform 1 0 620 0 -1 2828
box -36 -17 404 1471
use sky130_sram_1kbyte_1rw1r_8x1024_8_pinv_1  sky130_sram_1kbyte_1rw1r_8x1024_8_pinv_1_2
timestamp 1701704242
transform 1 0 620 0 1 0
box -36 -17 404 1471
<< labels >>
rlabel metal3 s 1841 1365 1939 1463 4 vdd
port 1 nsew
rlabel metal3 s 481 4193 579 4291 4 vdd
port 1 nsew
rlabel metal3 s 1841 4193 1939 4291 4 vdd
port 1 nsew
rlabel metal3 s 481 1365 579 1463 4 vdd
port 1 nsew
rlabel metal3 s 1841 9849 1939 9947 4 vdd
port 1 nsew
rlabel metal3 s 481 7021 579 7119 4 vdd
port 1 nsew
rlabel metal3 s 1841 7021 1939 7119 4 vdd
port 1 nsew
rlabel metal3 s 481 9849 579 9947 4 vdd
port 1 nsew
rlabel metal3 s 1841 5607 1939 5705 4 gnd
port 2 nsew
rlabel metal3 s 481 11263 579 11361 4 gnd
port 2 nsew
rlabel metal3 s 1841 8435 1939 8533 4 gnd
port 2 nsew
rlabel metal3 s 1841 -49 1939 49 4 gnd
port 2 nsew
rlabel metal3 s 1841 11263 1939 11361 4 gnd
port 2 nsew
rlabel metal3 s 481 5607 579 5705 4 gnd
port 2 nsew
rlabel metal3 s 1841 2779 1939 2877 4 gnd
port 2 nsew
rlabel metal3 s 481 -49 579 49 4 gnd
port 2 nsew
rlabel metal3 s 481 8435 579 8533 4 gnd
port 2 nsew
rlabel metal3 s 481 2779 579 2877 4 gnd
port 2 nsew
rlabel metal1 s 115 640 161 698 4 in_0
port 3 nsew
rlabel metal1 s 239 2130 285 2188 4 in_1
port 4 nsew
rlabel metal1 s 363 3468 409 3526 4 in_2
port 5 nsew
rlabel locali s 2654 669 2654 669 4 out_0
rlabel locali s 2654 2159 2654 2159 4 out_1
rlabel locali s 2654 3497 2654 3497 4 out_2
rlabel locali s 2654 4987 2654 4987 4 out_3
rlabel locali s 2654 6325 2654 6325 4 out_4
rlabel locali s 2654 7815 2654 7815 4 out_5
rlabel locali s 2654 9153 2654 9153 4 out_6
rlabel locali s 2654 10643 2654 10643 4 out_7
<< properties >>
string FIXED_BBOX 1857 -37 1923 0
string GDS_END 6125892
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_8x1024_8.gds
string GDS_START 6099732
<< end >>
