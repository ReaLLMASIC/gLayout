magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< pwell >>
rect -79 -26 1431 226
<< mvnmos >>
rect 0 0 120 200
rect 176 0 296 200
rect 352 0 472 200
rect 528 0 648 200
rect 704 0 824 200
rect 880 0 1000 200
rect 1056 0 1176 200
rect 1232 0 1352 200
<< mvndiff >>
rect -53 182 0 200
rect -53 148 -45 182
rect -11 148 0 182
rect -53 114 0 148
rect -53 80 -45 114
rect -11 80 0 114
rect -53 46 0 80
rect -53 12 -45 46
rect -11 12 0 46
rect -53 0 0 12
rect 120 182 176 200
rect 120 148 131 182
rect 165 148 176 182
rect 120 114 176 148
rect 120 80 131 114
rect 165 80 176 114
rect 120 46 176 80
rect 120 12 131 46
rect 165 12 176 46
rect 120 0 176 12
rect 296 182 352 200
rect 296 148 307 182
rect 341 148 352 182
rect 296 114 352 148
rect 296 80 307 114
rect 341 80 352 114
rect 296 46 352 80
rect 296 12 307 46
rect 341 12 352 46
rect 296 0 352 12
rect 472 182 528 200
rect 472 148 483 182
rect 517 148 528 182
rect 472 114 528 148
rect 472 80 483 114
rect 517 80 528 114
rect 472 46 528 80
rect 472 12 483 46
rect 517 12 528 46
rect 472 0 528 12
rect 648 182 704 200
rect 648 148 659 182
rect 693 148 704 182
rect 648 114 704 148
rect 648 80 659 114
rect 693 80 704 114
rect 648 46 704 80
rect 648 12 659 46
rect 693 12 704 46
rect 648 0 704 12
rect 824 182 880 200
rect 824 148 835 182
rect 869 148 880 182
rect 824 114 880 148
rect 824 80 835 114
rect 869 80 880 114
rect 824 46 880 80
rect 824 12 835 46
rect 869 12 880 46
rect 824 0 880 12
rect 1000 182 1056 200
rect 1000 148 1011 182
rect 1045 148 1056 182
rect 1000 114 1056 148
rect 1000 80 1011 114
rect 1045 80 1056 114
rect 1000 46 1056 80
rect 1000 12 1011 46
rect 1045 12 1056 46
rect 1000 0 1056 12
rect 1176 182 1232 200
rect 1176 148 1187 182
rect 1221 148 1232 182
rect 1176 114 1232 148
rect 1176 80 1187 114
rect 1221 80 1232 114
rect 1176 46 1232 80
rect 1176 12 1187 46
rect 1221 12 1232 46
rect 1176 0 1232 12
rect 1352 182 1405 200
rect 1352 148 1363 182
rect 1397 148 1405 182
rect 1352 114 1405 148
rect 1352 80 1363 114
rect 1397 80 1405 114
rect 1352 46 1405 80
rect 1352 12 1363 46
rect 1397 12 1405 46
rect 1352 0 1405 12
<< mvndiffc >>
rect -45 148 -11 182
rect -45 80 -11 114
rect -45 12 -11 46
rect 131 148 165 182
rect 131 80 165 114
rect 131 12 165 46
rect 307 148 341 182
rect 307 80 341 114
rect 307 12 341 46
rect 483 148 517 182
rect 483 80 517 114
rect 483 12 517 46
rect 659 148 693 182
rect 659 80 693 114
rect 659 12 693 46
rect 835 148 869 182
rect 835 80 869 114
rect 835 12 869 46
rect 1011 148 1045 182
rect 1011 80 1045 114
rect 1011 12 1045 46
rect 1187 148 1221 182
rect 1187 80 1221 114
rect 1187 12 1221 46
rect 1363 148 1397 182
rect 1363 80 1397 114
rect 1363 12 1397 46
<< poly >>
rect 0 200 120 226
rect 176 200 296 226
rect 352 200 472 226
rect 528 200 648 226
rect 704 200 824 226
rect 880 200 1000 226
rect 1056 200 1176 226
rect 1232 200 1352 226
rect 0 -26 120 0
rect 176 -26 296 0
rect 352 -26 472 0
rect 528 -26 648 0
rect 704 -26 824 0
rect 880 -26 1000 0
rect 1056 -26 1176 0
rect 1232 -26 1352 0
<< locali >>
rect -45 182 -11 198
rect -45 114 -11 148
rect -45 46 -11 80
rect -45 -4 -11 12
rect 131 182 165 198
rect 131 114 165 148
rect 131 46 165 80
rect 131 -4 165 12
rect 307 182 341 198
rect 307 114 341 148
rect 307 46 341 80
rect 307 -4 341 12
rect 483 182 517 198
rect 483 114 517 148
rect 483 46 517 80
rect 483 -4 517 12
rect 659 182 693 198
rect 659 114 693 148
rect 659 46 693 80
rect 659 -4 693 12
rect 835 182 869 198
rect 835 114 869 148
rect 835 46 869 80
rect 835 -4 869 12
rect 1011 182 1045 198
rect 1011 114 1045 148
rect 1011 46 1045 80
rect 1011 -4 1045 12
rect 1187 182 1221 198
rect 1187 114 1221 148
rect 1187 46 1221 80
rect 1187 -4 1221 12
rect 1363 182 1397 198
rect 1363 114 1397 148
rect 1363 46 1397 80
rect 1363 -4 1397 12
use hvDFL1sd2_CDNS_52468879185133  hvDFL1sd2_CDNS_52468879185133_0
timestamp 1701704242
transform 1 0 1176 0 1 0
box 0 0 1 1
use hvDFL1sd2_CDNS_52468879185133  hvDFL1sd2_CDNS_52468879185133_1
timestamp 1701704242
transform 1 0 1000 0 1 0
box 0 0 1 1
use hvDFL1sd2_CDNS_52468879185133  hvDFL1sd2_CDNS_52468879185133_2
timestamp 1701704242
transform 1 0 824 0 1 0
box 0 0 1 1
use hvDFL1sd2_CDNS_52468879185133  hvDFL1sd2_CDNS_52468879185133_3
timestamp 1701704242
transform 1 0 648 0 1 0
box 0 0 1 1
use hvDFL1sd2_CDNS_52468879185133  hvDFL1sd2_CDNS_52468879185133_4
timestamp 1701704242
transform 1 0 472 0 1 0
box 0 0 1 1
use hvDFL1sd2_CDNS_52468879185133  hvDFL1sd2_CDNS_52468879185133_5
timestamp 1701704242
transform 1 0 296 0 1 0
box 0 0 1 1
use hvDFL1sd2_CDNS_52468879185133  hvDFL1sd2_CDNS_52468879185133_6
timestamp 1701704242
transform 1 0 120 0 1 0
box 0 0 1 1
use hvDFL1sd_CDNS_52468879185132  hvDFL1sd_CDNS_52468879185132_0
timestamp 1701704242
transform -1 0 0 0 1 0
box 0 0 1 1
use hvDFL1sd_CDNS_52468879185132  hvDFL1sd_CDNS_52468879185132_1
timestamp 1701704242
transform 1 0 1352 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s -28 97 -28 97 0 FreeSans 300 0 0 0 S
flabel comment s 148 97 148 97 0 FreeSans 300 0 0 0 D
flabel comment s 324 97 324 97 0 FreeSans 300 0 0 0 S
flabel comment s 500 97 500 97 0 FreeSans 300 0 0 0 D
flabel comment s 676 97 676 97 0 FreeSans 300 0 0 0 S
flabel comment s 852 97 852 97 0 FreeSans 300 0 0 0 D
flabel comment s 1028 97 1028 97 0 FreeSans 300 0 0 0 S
flabel comment s 1204 97 1204 97 0 FreeSans 300 0 0 0 D
flabel comment s 1380 97 1380 97 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 79666294
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 79661328
<< end >>
