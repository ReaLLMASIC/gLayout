magic
tech sky130B
timestamp 1701704242
<< metal1 >>
rect 0 0 3 218
rect 61 0 64 218
<< via1 >>
rect 3 0 61 218
<< metal2 >>
rect 0 0 3 218
rect 61 0 64 218
<< properties >>
string GDS_END 86906544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86905516
<< end >>
