magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 417 157 735 203
rect 1 21 735 157
rect 30 -17 64 21
<< locali >>
rect 25 151 66 415
rect 547 299 614 493
rect 178 84 249 265
rect 284 261 318 265
rect 284 83 344 261
rect 380 83 432 265
rect 579 161 614 299
rect 547 68 614 161
rect 547 59 613 68
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 19 451 85 527
rect 120 333 170 493
rect 214 383 280 527
rect 317 333 367 493
rect 447 367 513 527
rect 100 299 511 333
rect 649 367 715 527
rect 100 117 134 299
rect 35 51 134 117
rect 466 263 511 299
rect 466 215 545 263
rect 466 17 513 178
rect 651 17 717 162
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
rlabel locali s 25 151 66 415 6 A
port 1 nsew signal input
rlabel locali s 178 84 249 265 6 B
port 2 nsew signal input
rlabel locali s 284 83 344 261 6 C
port 3 nsew signal input
rlabel locali s 284 261 318 265 6 C
port 3 nsew signal input
rlabel locali s 380 83 432 265 6 D
port 4 nsew signal input
rlabel metal1 s 0 -48 736 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1 21 735 157 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 417 157 735 203 6 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 774 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 736 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 547 59 613 68 6 X
port 9 nsew signal output
rlabel locali s 547 68 614 161 6 X
port 9 nsew signal output
rlabel locali s 579 161 614 299 6 X
port 9 nsew signal output
rlabel locali s 547 299 614 493 6 X
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 736 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 3892210
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3884992
<< end >>
