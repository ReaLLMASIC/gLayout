magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< metal3 >>
rect 0 12361 1000 13599
rect 0 11003 1000 12241
rect 0 9645 1000 10883
rect 0 8287 1000 9525
rect 0 6929 1000 8167
rect 0 5492 1000 6809
rect 0 4134 1000 5372
rect 0 2776 1000 4014
rect 0 1418 1000 2656
rect 0 250 1000 1298
<< properties >>
string GDS_END 78395150
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 78394506
<< end >>
