magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< nwell >>
rect 3981 -8 4257 557
<< pwell >>
rect 12694 2702 12871 2790
rect 13253 2702 13333 2790
rect 4161 1248 4247 2211
rect 4161 617 4247 896
<< psubdiff >>
rect 4187 820 4221 870
rect 4187 701 4221 786
rect 4187 643 4221 667
<< nsubdiff >>
rect 4187 497 4221 521
rect 4187 428 4221 463
rect 4187 359 4221 394
rect 4187 290 4221 325
rect 4187 222 4221 256
rect 4187 154 4221 188
rect 4187 86 4221 120
rect 4187 28 4221 52
<< mvpsubdiff >>
rect 12720 2728 12845 2764
rect 13279 2728 13307 2764
rect 4187 2161 4221 2185
rect 4187 2091 4221 2127
rect 4187 2022 4221 2057
rect 4187 1953 4221 1988
rect 4187 1884 4221 1919
rect 4187 1815 4221 1850
rect 4187 1746 4221 1781
rect 4187 1677 4221 1712
rect 4187 1608 4221 1643
rect 4187 1539 4221 1574
rect 4187 1470 4221 1505
rect 4187 1401 4221 1436
rect 4187 1332 4221 1367
rect 4187 1274 4221 1298
<< mvnsubdiff >>
rect 12714 2916 12845 2952
rect 13279 2916 13307 2952
<< psubdiffcont >>
rect 4187 786 4221 820
rect 4187 667 4221 701
<< nsubdiffcont >>
rect 4187 463 4221 497
rect 4187 394 4221 428
rect 4187 325 4221 359
rect 4187 256 4221 290
rect 4187 188 4221 222
rect 4187 120 4221 154
rect 4187 52 4221 86
<< mvpsubdiffcont >>
rect 4187 2127 4221 2161
rect 4187 2057 4221 2091
rect 4187 1988 4221 2022
rect 4187 1919 4221 1953
rect 4187 1850 4221 1884
rect 4187 1781 4221 1815
rect 4187 1712 4221 1746
rect 4187 1643 4221 1677
rect 4187 1574 4221 1608
rect 4187 1505 4221 1539
rect 4187 1436 4221 1470
rect 4187 1367 4221 1401
rect 4187 1298 4221 1332
<< locali >>
rect 11654 3639 11932 3705
rect 13133 3654 13167 3704
rect 11424 3555 11458 3604
rect 7277 3510 7311 3550
rect 11086 3192 11282 3544
rect 12713 3192 12903 3544
rect 13971 3396 14009 3430
rect 13045 3358 13079 3396
rect 13793 3278 13827 3316
rect 14269 3278 14303 3316
rect 11192 3014 11282 3192
rect 12741 3158 12790 3192
rect 12824 3158 12903 3192
rect 12707 3120 12903 3158
rect 12741 3086 12790 3120
rect 12824 3086 12903 3120
rect 12707 3048 12903 3086
rect 12741 3014 12790 3048
rect 12824 3014 12903 3048
rect 11086 2968 11282 3014
rect 12713 2968 12903 3014
rect 14729 3192 14902 3544
rect 14729 3158 14868 3192
rect 14729 3120 14902 3158
rect 14729 3086 14868 3120
rect 14729 3048 14902 3086
rect 14729 3014 14868 3048
rect 13221 2968 13255 3002
rect 9429 2902 9524 2968
rect 11086 2934 11176 2968
rect 11210 2934 11248 2968
rect 11086 2902 11282 2934
rect 11895 2926 12085 2968
rect 12713 2934 12790 2968
rect 12824 2934 12903 2968
rect 12713 2902 12903 2934
rect 13255 2902 13348 2968
rect 14729 2902 14902 3014
rect 11520 2820 11554 2858
rect 11776 2820 11810 2858
rect 11952 2820 11986 2858
rect 12158 2820 12192 2858
rect 14201 2820 14235 2858
rect 14465 2820 14499 2858
rect 14641 2820 14675 2858
rect 9429 2712 9514 2778
rect 11118 2746 11248 2778
rect 12707 2746 12869 2778
rect 11118 2712 11176 2746
rect 11210 2712 11248 2746
rect 12707 2712 12788 2746
rect 12822 2712 12869 2746
rect 13255 2712 13345 2778
rect 14763 2712 14902 2778
rect 8839 2548 8873 2592
rect 5473 2456 5507 2506
rect 9395 2456 9539 2666
rect 10061 2511 10095 2555
rect 10413 2508 10447 2550
rect 13221 2456 13365 2666
rect 14553 2506 14587 2556
rect 12340 2408 12378 2442
rect 6179 2370 6213 2408
rect 6342 2356 6380 2390
rect 12489 2334 12527 2368
rect 13605 2356 13643 2390
rect 233 2254 271 2288
rect 739 2254 777 2288
rect 811 2254 849 2288
rect 883 2254 921 2288
rect 3283 2254 3321 2288
rect 3355 2254 3393 2288
rect 3427 2254 3465 2288
rect 3499 2254 3537 2288
rect 3571 2254 3609 2288
rect 3744 2254 3782 2288
rect 3985 2254 4387 2288
rect 4628 2254 4666 2288
rect 4799 2254 4837 2288
rect 4871 2254 4909 2288
rect 4943 2254 4981 2288
rect 5015 2254 5053 2288
rect 5087 2254 5125 2288
rect 4187 2161 4221 2185
rect 4187 2091 4221 2127
rect 4187 2022 4221 2057
rect 4187 1972 4221 1988
rect 4187 1953 4190 1972
rect 4221 1919 4224 1938
rect 4187 1900 4224 1919
rect 4187 1884 4190 1900
rect 4187 1815 4221 1850
rect 4187 1746 4221 1781
rect 4187 1677 4221 1712
rect 4187 1608 4221 1643
rect 4187 1539 4221 1574
rect 4187 1470 4221 1505
rect 4187 1401 4221 1436
rect 4187 1332 4221 1367
rect 2495 646 2529 1032
rect 4187 820 4221 870
rect 4187 701 4221 786
rect 4187 643 4221 665
rect 2495 574 2529 612
rect 4187 497 4221 521
rect 4187 428 4221 463
rect 4187 359 4221 394
rect 4187 290 4221 325
rect 4187 222 4221 256
rect 4187 154 4221 188
rect 4187 86 4221 120
rect 4187 28 4221 52
<< viali >>
rect 13045 3396 13079 3430
rect 13937 3396 13971 3430
rect 14009 3396 14043 3430
rect 13045 3324 13079 3358
rect 13793 3316 13827 3350
rect 13793 3244 13827 3278
rect 14269 3316 14303 3350
rect 14269 3244 14303 3278
rect 11086 3014 11192 3192
rect 12707 3158 12741 3192
rect 12790 3158 12824 3192
rect 12707 3086 12741 3120
rect 12790 3086 12824 3120
rect 12707 3014 12741 3048
rect 12790 3014 12824 3048
rect 14868 3158 14902 3192
rect 14868 3086 14902 3120
rect 14868 3014 14902 3048
rect 11176 2934 11210 2968
rect 11248 2934 11282 2968
rect 12790 2934 12824 2968
rect 11520 2858 11554 2892
rect 11520 2786 11554 2820
rect 11776 2858 11810 2892
rect 11776 2786 11810 2820
rect 11952 2858 11986 2892
rect 11952 2786 11986 2820
rect 12158 2858 12192 2892
rect 12158 2786 12192 2820
rect 14201 2858 14235 2892
rect 14201 2786 14235 2820
rect 14465 2858 14499 2892
rect 14465 2786 14499 2820
rect 14641 2858 14675 2892
rect 14641 2786 14675 2820
rect 11176 2712 11210 2746
rect 11248 2712 11282 2746
rect 12788 2712 12822 2746
rect 6179 2408 6213 2442
rect 12306 2408 12340 2442
rect 12378 2408 12412 2442
rect 13432 2403 13466 2437
rect 6179 2336 6213 2370
rect 6308 2356 6342 2390
rect 6380 2356 6414 2390
rect 12455 2334 12489 2368
rect 12527 2334 12561 2368
rect 13571 2356 13605 2390
rect 13643 2356 13677 2390
rect 199 2254 233 2288
rect 271 2254 305 2288
rect 705 2254 739 2288
rect 777 2254 811 2288
rect 849 2254 883 2288
rect 921 2254 955 2288
rect 3249 2254 3283 2288
rect 3321 2254 3355 2288
rect 3393 2254 3427 2288
rect 3465 2254 3499 2288
rect 3537 2254 3571 2288
rect 3609 2254 3643 2288
rect 3710 2254 3744 2288
rect 3782 2254 3816 2288
rect 4594 2254 4628 2288
rect 4666 2254 4700 2288
rect 4765 2254 4799 2288
rect 4837 2254 4871 2288
rect 4909 2254 4943 2288
rect 4981 2254 5015 2288
rect 5053 2254 5087 2288
rect 5125 2254 5159 2288
rect 4190 1953 4224 1972
rect 4190 1938 4221 1953
rect 4221 1938 4224 1953
rect 4190 1884 4224 1900
rect 4190 1866 4221 1884
rect 4221 1866 4224 1884
rect 4187 1298 4221 1306
rect 4187 1272 4221 1298
rect 2495 612 2529 646
rect 4187 667 4221 699
rect 4187 665 4221 667
rect 2495 540 2529 574
<< metal1 >>
rect 2402 3618 2436 3652
rect 223 3501 257 3535
rect 13033 3430 14055 3436
rect 2869 3396 2903 3430
rect 13033 3396 13045 3430
rect 13079 3396 13937 3430
rect 13971 3396 14009 3430
rect 14043 3396 14055 3430
rect 13033 3390 14055 3396
rect 13033 3358 13091 3390
tri 13091 3365 13116 3390 nw
rect 563 3310 597 3344
rect 13033 3324 13045 3358
rect 13079 3324 13091 3358
rect 13033 3318 13091 3324
rect 13561 3350 13833 3362
rect 13561 3316 13793 3350
rect 13827 3316 13833 3350
rect 13561 3278 13833 3316
rect 13561 3244 13793 3278
rect 13827 3244 13833 3278
rect 13561 3232 13833 3244
rect 13861 3361 13901 3362
rect 13861 3355 13913 3361
rect 13861 3291 13913 3303
rect 13861 3233 13913 3239
rect 14131 3350 14309 3362
rect 14131 3316 14269 3350
rect 14303 3316 14309 3350
rect 14131 3278 14309 3316
rect 14131 3244 14269 3278
rect 14303 3244 14309 3278
rect 13861 3232 13901 3233
rect 14131 3232 14309 3244
rect 117 3002 129 3204
rect 11080 3192 11258 3204
rect 11080 3014 11086 3192
rect 11192 3014 11258 3192
rect 11080 3002 11258 3014
rect 11969 3002 12079 3204
rect 12693 3192 12979 3204
rect 12693 3158 12707 3192
rect 12741 3158 12790 3192
rect 12824 3158 12979 3192
rect 12693 3120 12979 3158
rect 12693 3086 12707 3120
rect 12741 3086 12790 3120
rect 12824 3086 12979 3120
rect 12693 3048 12979 3086
rect 12693 3014 12707 3048
rect 12741 3014 12790 3048
rect 12824 3014 12979 3048
rect 12693 3002 12979 3014
rect 13238 3002 13348 3204
rect 14108 3002 14218 3204
rect 14862 3192 14908 3204
rect 14862 3158 14868 3192
rect 14902 3158 14908 3192
rect 14862 3120 14908 3158
rect 14862 3086 14868 3120
rect 14902 3086 14908 3120
rect 14862 3048 14908 3086
rect 14862 3014 14868 3048
rect 14902 3014 14908 3048
rect 14862 3002 14908 3014
rect 11117 2968 14914 3002
rect 11117 2934 11176 2968
rect 11210 2934 11248 2968
rect 11282 2934 12790 2968
rect 12824 2934 14914 2968
rect 11117 2928 14914 2934
tri 5642 2848 5648 2854 ne
rect 5648 2848 5654 2900
rect 5706 2848 5718 2900
rect 5770 2848 5776 2900
rect 11508 2892 11998 2898
rect 11508 2858 11520 2892
rect 11554 2858 11776 2892
rect 11810 2858 11952 2892
rect 11986 2858 11998 2892
tri 5776 2848 5782 2854 nw
rect 11508 2820 11998 2858
rect 11508 2786 11520 2820
rect 11554 2786 11776 2820
rect 11810 2786 11952 2820
rect 11986 2786 11998 2820
rect 11508 2780 11998 2786
rect 12146 2892 12204 2898
rect 12146 2858 12158 2892
rect 12192 2858 12204 2892
rect 12146 2826 12204 2858
rect 13439 2896 14687 2898
tri 12204 2826 12229 2851 sw
rect 13439 2844 13445 2896
rect 13497 2892 14687 2896
rect 13497 2858 14201 2892
rect 14235 2858 14465 2892
rect 14499 2858 14641 2892
rect 14675 2858 14687 2892
rect 13497 2844 14687 2858
rect 13439 2832 14687 2844
rect 12146 2820 12402 2826
rect 12146 2786 12158 2820
rect 12192 2786 12402 2820
rect 12146 2780 12402 2786
rect 13439 2780 13445 2832
rect 13497 2820 14687 2832
rect 13497 2786 14201 2820
rect 14235 2786 14465 2820
rect 14499 2786 14641 2820
rect 14675 2786 14687 2820
rect 13497 2780 14687 2786
rect 117 2706 129 2752
rect 11117 2746 11294 2752
rect 11117 2712 11176 2746
rect 11210 2712 11248 2746
rect 11282 2712 11294 2746
rect 11117 2706 11294 2712
rect 11969 2706 12079 2752
rect 12693 2746 12979 2752
rect 12693 2712 12788 2746
rect 12822 2712 12979 2746
rect 12693 2706 12979 2712
rect 13238 2706 13348 2752
rect 14108 2706 14218 2752
rect 117 2476 129 2678
rect 3698 2662 3814 2668
rect 3698 2476 3814 2482
rect 4596 2662 4712 2668
rect 4596 2476 4712 2482
rect 11117 2476 11258 2678
rect 11969 2476 12079 2678
rect 12693 2476 13142 2678
rect 13238 2476 13348 2678
rect 14108 2476 14218 2678
rect 6167 2442 6264 2448
tri 10919 2442 10925 2448 se
rect 10925 2443 13331 2448
tri 13331 2443 13336 2448 sw
rect 10925 2442 13478 2443
rect 363 2404 397 2438
rect 3399 2378 3434 2412
rect 6219 2390 6264 2442
tri 10885 2408 10919 2442 se
rect 10919 2408 12306 2442
rect 12340 2408 12378 2442
rect 12412 2437 13478 2442
rect 12412 2408 13432 2437
tri 10880 2403 10885 2408 se
rect 10885 2403 13432 2408
rect 13466 2403 13478 2437
tri 10879 2402 10880 2403 se
rect 10880 2402 13478 2403
tri 10874 2397 10879 2402 se
rect 10879 2397 10940 2402
tri 10940 2397 10945 2402 nw
tri 13311 2397 13316 2402 ne
rect 13316 2397 13478 2402
tri 10873 2396 10874 2397 se
rect 10874 2396 10939 2397
tri 10939 2396 10940 2397 nw
rect 6167 2378 6264 2390
rect 295 2364 347 2370
tri 270 2294 295 2319 se
rect 6219 2326 6264 2378
rect 6296 2394 6601 2396
tri 6601 2394 6603 2396 sw
tri 10871 2394 10873 2396 se
rect 10873 2394 10937 2396
tri 10937 2394 10939 2396 nw
rect 6296 2390 6603 2394
tri 6603 2390 6607 2394 sw
tri 10867 2390 10871 2394 se
rect 10871 2390 10933 2394
tri 10933 2390 10937 2394 nw
tri 13555 2390 13559 2394 se
rect 13559 2390 13689 2402
rect 6296 2356 6308 2390
rect 6342 2356 6380 2390
rect 6414 2382 6607 2390
tri 6607 2382 6615 2390 sw
tri 10859 2382 10867 2390 se
rect 10867 2382 10925 2390
tri 10925 2382 10933 2390 nw
tri 13547 2382 13555 2390 se
rect 13555 2382 13571 2390
rect 6414 2378 6615 2382
tri 6615 2378 6619 2382 sw
tri 10855 2378 10859 2382 se
rect 10859 2378 10917 2382
rect 6414 2374 6619 2378
tri 6619 2374 6623 2378 sw
tri 10851 2374 10855 2378 se
rect 10855 2374 10917 2378
tri 10917 2374 10925 2382 nw
tri 13539 2374 13547 2382 se
rect 13547 2374 13571 2382
rect 6414 2368 6623 2374
tri 6623 2368 6629 2374 sw
tri 10845 2368 10851 2374 se
rect 10851 2368 10911 2374
tri 10911 2368 10917 2374 nw
rect 6414 2356 6629 2368
rect 6296 2350 6629 2356
tri 6629 2350 6647 2368 sw
tri 10827 2350 10845 2368 se
rect 10845 2350 10877 2368
tri 6581 2334 6597 2350 ne
rect 6597 2334 6647 2350
tri 6647 2334 6663 2350 sw
tri 10811 2334 10827 2350 se
rect 10827 2334 10877 2350
tri 10877 2334 10911 2368 nw
rect 6167 2320 6264 2326
tri 6597 2320 6611 2334 ne
rect 6611 2322 6663 2334
tri 6663 2322 6675 2334 sw
tri 10799 2322 10811 2334 se
rect 10811 2322 10865 2334
tri 10865 2322 10877 2334 nw
rect 12095 2322 12101 2374
rect 12153 2322 12165 2374
rect 12217 2368 12573 2374
tri 13534 2369 13539 2374 se
rect 13539 2369 13571 2374
rect 12217 2334 12455 2368
rect 12489 2334 12527 2368
rect 12561 2334 12573 2368
rect 12217 2322 12573 2334
rect 6611 2320 6675 2322
tri 6675 2320 6677 2322 sw
tri 10797 2320 10799 2322 se
rect 10799 2320 10860 2322
tri 6611 2312 6619 2320 ne
rect 6619 2317 6677 2320
tri 6677 2317 6680 2320 sw
tri 10794 2317 10797 2320 se
rect 10797 2317 10860 2320
tri 10860 2317 10865 2322 nw
rect 13295 2317 13301 2369
rect 13353 2317 13365 2369
rect 13417 2356 13571 2369
rect 13605 2356 13643 2390
rect 13677 2356 13689 2390
rect 13417 2317 13689 2356
rect 6619 2316 6680 2317
tri 6680 2316 6681 2317 sw
tri 10793 2316 10794 2317 se
rect 10794 2316 10859 2317
tri 10859 2316 10860 2317 nw
rect 6619 2312 6681 2316
tri 6681 2312 6685 2316 sw
tri 10789 2312 10793 2316 se
rect 10793 2312 10855 2316
tri 10855 2312 10859 2316 nw
rect 295 2300 347 2312
tri 6619 2306 6625 2312 ne
rect 6625 2306 10809 2312
rect 187 2288 295 2294
rect 3698 2300 3828 2306
rect 187 2254 199 2288
rect 233 2254 271 2288
rect 187 2248 295 2254
rect 187 2242 347 2248
rect 693 2288 3396 2294
rect 693 2254 705 2288
rect 739 2254 777 2288
rect 811 2254 849 2288
rect 883 2254 921 2288
rect 955 2254 3249 2288
rect 3283 2254 3321 2288
rect 3355 2254 3393 2288
rect 693 2242 3396 2254
rect 3448 2242 3460 2294
rect 3512 2288 3655 2294
rect 3512 2254 3537 2288
rect 3571 2254 3609 2288
rect 3643 2254 3655 2288
rect 3512 2242 3655 2254
rect 3750 2248 3762 2300
rect 3814 2288 3828 2300
rect 4582 2300 4712 2306
rect 3816 2254 3828 2288
rect 3814 2248 3828 2254
rect 3698 2242 3828 2248
rect 3856 2242 3862 2294
rect 3914 2242 3926 2294
rect 3978 2242 4521 2294
rect 4582 2288 4596 2300
rect 4582 2254 4594 2288
rect 4582 2248 4596 2254
rect 4648 2248 4660 2300
tri 6625 2294 6637 2306 ne
rect 6637 2294 10809 2306
rect 4582 2242 4712 2248
rect 4740 2242 4746 2294
rect 4798 2288 4810 2294
rect 4862 2288 5171 2294
rect 4799 2254 4810 2288
rect 4871 2254 4909 2288
rect 4943 2254 4981 2288
rect 5015 2254 5053 2288
rect 5087 2254 5125 2288
rect 5159 2254 5171 2288
tri 6637 2266 6665 2294 ne
rect 6665 2266 10809 2294
tri 10809 2266 10855 2312 nw
rect 4798 2242 4810 2254
rect 4862 2242 5171 2254
rect -11 2034 -5 2214
rect 111 2034 117 2214
rect 4165 2012 16040 2214
rect 4165 1976 16040 1984
rect 4165 1924 4178 1976
rect 4230 1924 16040 1976
rect 4165 1912 16040 1924
rect 4165 1860 4178 1912
rect 4230 1860 16040 1912
rect 4165 1854 16040 1860
rect 295 1774 301 1826
rect 353 1774 365 1826
rect 417 1774 3862 1826
rect 3914 1774 3926 1826
rect 3978 1774 3984 1826
rect 5648 1774 5654 1826
rect 5706 1774 5718 1826
rect 5770 1774 13301 1826
rect 13353 1774 13365 1826
rect 13417 1774 13423 1826
rect 3390 1694 3396 1746
rect 3448 1694 3460 1746
rect 3512 1694 4746 1746
rect 4798 1694 4810 1746
rect 4862 1694 4868 1746
rect 13343 1737 13503 1746
rect 6216 1648 12101 1654
rect 2373 1641 2524 1647
rect 1747 1607 1781 1641
rect 2373 1589 2472 1641
rect 2373 1577 2524 1589
rect 2373 1525 2472 1577
rect 6268 1602 12101 1648
rect 12153 1602 12165 1654
rect 12217 1602 12434 1654
rect 13343 1621 13381 1737
rect 13497 1621 13503 1737
rect 13941 1624 16041 1826
rect 13343 1616 13503 1621
rect 6216 1584 6268 1596
tri 6268 1577 6293 1602 nw
rect 6216 1526 6268 1532
rect 2373 1519 2524 1525
rect 4178 1471 4230 1493
tri 4153 1415 4178 1440 se
rect 4178 1407 4230 1419
tri 4230 1415 4255 1440 sw
tri 4153 1338 4178 1363 ne
rect 4178 1343 4230 1355
tri 4230 1338 4255 1363 nw
rect 4178 1279 4187 1291
rect 4221 1279 4230 1291
rect 98 1221 132 1255
rect 4071 1221 4106 1255
rect 4178 1215 4230 1227
tri 4153 1145 4178 1170 se
rect 13343 1215 13837 1223
rect 4178 1151 4230 1163
tri 4230 1145 4255 1170 sw
rect 13343 1163 13599 1215
rect 13651 1163 13837 1215
rect 13343 1151 13837 1163
rect 4178 1093 4230 1099
rect 13343 1099 13599 1151
rect 13651 1099 13837 1151
rect 13343 1093 13837 1099
rect 14035 1093 16041 1295
rect 4171 863 16041 1065
tri 15761 838 15786 863 ne
rect 1990 789 2214 835
rect 4023 789 5440 835
tri 4072 764 4097 789 nw
rect 13905 783 15094 835
rect 15146 783 15158 835
rect 15210 783 15222 835
rect 15274 783 15286 835
rect 15338 783 15350 835
rect 15402 783 15408 835
rect 13905 729 15408 783
rect 4172 711 4300 717
rect 4172 659 4178 711
rect 4230 659 4242 711
rect 4294 659 4300 711
rect 2472 650 2535 658
rect 4172 653 4300 659
rect 6216 713 6268 719
rect 2524 646 2535 650
rect 2529 612 2535 646
tri 6209 643 6216 650 se
rect 6216 649 6268 661
rect 2524 598 2535 612
rect 2472 586 2535 598
rect 2632 591 2638 643
rect 2690 591 2702 643
rect 2754 625 2760 643
tri 2760 625 2778 643 sw
tri 6191 625 6209 643 se
rect 6209 625 6216 643
rect 2754 597 6216 625
rect 2754 591 6268 597
tri 15774 591 15786 603 se
rect 15786 591 15916 863
tri 15916 838 15941 863 nw
tri 15770 587 15774 591 se
rect 15774 587 15916 591
rect 2524 578 2535 586
tri 2535 578 2544 587 sw
tri 15761 578 15770 587 se
rect 15770 578 15916 587
rect 2524 576 2544 578
tri 2544 576 2546 578 sw
rect 2524 574 2546 576
rect 2529 562 2546 574
tri 2546 562 2560 576 sw
tri 15074 562 15088 576 se
rect 15088 570 15204 576
rect 2529 554 6256 562
tri 6256 554 6264 562 sw
tri 15066 554 15074 562 se
rect 15074 554 15088 562
rect 2529 540 6142 554
rect 2524 534 6142 540
rect 2472 528 6142 534
tri 5726 502 5752 528 ne
rect 5752 502 6142 528
rect 6194 502 6206 554
rect 6258 502 6264 554
tri 15062 550 15066 554 se
rect 15066 550 15088 554
rect 13899 454 15088 550
rect 13899 448 15204 454
rect 15238 448 15916 578
rect 2078 218 2127 420
rect 9540 395 9907 420
tri 9907 395 9932 420 sw
tri 10210 395 10235 420 se
rect 10235 395 16041 420
rect -2 72 16 190
rect 9540 72 16041 395
<< via1 >>
rect 13861 3303 13913 3355
rect 13861 3239 13913 3291
rect 5654 2848 5706 2900
rect 5718 2848 5770 2900
rect 13445 2844 13497 2896
rect 13445 2780 13497 2832
rect 3698 2482 3814 2662
rect 4596 2482 4712 2662
rect 6167 2408 6179 2442
rect 6179 2408 6213 2442
rect 6213 2408 6219 2442
rect 6167 2390 6219 2408
rect 6167 2370 6219 2378
rect 295 2312 347 2364
rect 6167 2336 6179 2370
rect 6179 2336 6213 2370
rect 6213 2336 6219 2370
rect 6167 2326 6219 2336
rect 12101 2322 12153 2374
rect 12165 2322 12217 2374
rect 13301 2317 13353 2369
rect 13365 2317 13417 2369
rect 295 2288 347 2300
rect 295 2254 305 2288
rect 305 2254 347 2288
rect 295 2248 347 2254
rect 3396 2288 3448 2294
rect 3396 2254 3427 2288
rect 3427 2254 3448 2288
rect 3396 2242 3448 2254
rect 3460 2288 3512 2294
rect 3460 2254 3465 2288
rect 3465 2254 3499 2288
rect 3499 2254 3512 2288
rect 3460 2242 3512 2254
rect 3698 2288 3750 2300
rect 3698 2254 3710 2288
rect 3710 2254 3744 2288
rect 3744 2254 3750 2288
rect 3698 2248 3750 2254
rect 3762 2288 3814 2300
rect 3762 2254 3782 2288
rect 3782 2254 3814 2288
rect 3762 2248 3814 2254
rect 3862 2242 3914 2294
rect 3926 2242 3978 2294
rect 4596 2288 4648 2300
rect 4596 2254 4628 2288
rect 4628 2254 4648 2288
rect 4596 2248 4648 2254
rect 4660 2288 4712 2300
rect 4660 2254 4666 2288
rect 4666 2254 4700 2288
rect 4700 2254 4712 2288
rect 4660 2248 4712 2254
rect 4746 2288 4798 2294
rect 4810 2288 4862 2294
rect 4746 2254 4765 2288
rect 4765 2254 4798 2288
rect 4810 2254 4837 2288
rect 4837 2254 4862 2288
rect 4746 2242 4798 2254
rect 4810 2242 4862 2254
rect -5 2034 111 2214
rect 4178 1972 4230 1976
rect 4178 1938 4190 1972
rect 4190 1938 4224 1972
rect 4224 1938 4230 1972
rect 4178 1924 4230 1938
rect 4178 1900 4230 1912
rect 4178 1866 4190 1900
rect 4190 1866 4224 1900
rect 4224 1866 4230 1900
rect 4178 1860 4230 1866
rect 301 1774 353 1826
rect 365 1774 417 1826
rect 3862 1774 3914 1826
rect 3926 1774 3978 1826
rect 5654 1774 5706 1826
rect 5718 1774 5770 1826
rect 13301 1774 13353 1826
rect 13365 1774 13417 1826
rect 3396 1694 3448 1746
rect 3460 1694 3512 1746
rect 4746 1694 4798 1746
rect 4810 1694 4862 1746
rect 2472 1589 2524 1641
rect 2472 1525 2524 1577
rect 6216 1596 6268 1648
rect 12101 1602 12153 1654
rect 12165 1602 12217 1654
rect 13381 1621 13497 1737
rect 6216 1532 6268 1584
rect 4178 1419 4230 1471
rect 4178 1355 4230 1407
rect 4178 1306 4230 1343
rect 4178 1291 4187 1306
rect 4187 1291 4221 1306
rect 4221 1291 4230 1306
rect 4178 1272 4187 1279
rect 4187 1272 4221 1279
rect 4221 1272 4230 1279
rect 4178 1227 4230 1272
rect 4178 1163 4230 1215
rect 4178 1099 4230 1151
rect 13599 1163 13651 1215
rect 13599 1099 13651 1151
rect 15094 783 15146 835
rect 15158 783 15210 835
rect 15222 783 15274 835
rect 15286 783 15338 835
rect 15350 783 15402 835
rect 4178 699 4230 711
rect 4178 665 4187 699
rect 4187 665 4221 699
rect 4221 665 4230 699
rect 4178 659 4230 665
rect 4242 659 4294 711
rect 6216 661 6268 713
rect 2472 646 2524 650
rect 2472 612 2495 646
rect 2495 612 2524 646
rect 2472 598 2524 612
rect 2638 591 2690 643
rect 2702 591 2754 643
rect 6216 597 6268 649
rect 2472 574 2524 586
rect 2472 540 2495 574
rect 2495 540 2524 574
rect 2472 534 2524 540
rect 6142 502 6194 554
rect 6206 502 6258 554
rect 15088 454 15204 570
<< metal2 >>
rect 13599 3355 13913 3361
rect 13599 3303 13861 3355
rect 13599 3291 13913 3303
rect 13599 3239 13861 3291
rect 13599 3233 13913 3239
rect -11 2214 117 2960
rect 5648 2848 5654 2900
rect 5706 2848 5718 2900
rect 5770 2848 5776 2900
tri 5699 2844 5703 2848 ne
rect 5703 2844 5776 2848
tri 5703 2832 5715 2844 ne
rect 5715 2832 5776 2844
tri 5715 2823 5724 2832 ne
rect 3698 2662 3814 2668
rect -11 2034 -5 2214
rect 111 2034 117 2214
rect 295 2364 347 2370
rect 295 2300 347 2312
rect 3698 2300 3814 2482
rect 295 1826 347 2248
rect 3390 2242 3396 2294
rect 3448 2242 3460 2294
rect 3512 2242 3518 2294
rect 3750 2248 3762 2300
rect 4596 2662 4712 2668
rect 4596 2300 4712 2482
rect 3698 2242 3814 2248
rect 3856 2242 3862 2294
rect 3914 2242 3926 2294
rect 3978 2242 3984 2294
rect 4648 2248 4660 2300
rect 4596 2242 4712 2248
rect 4740 2242 4746 2294
rect 4798 2242 4810 2294
rect 4862 2242 4868 2294
tri 347 1826 372 1851 sw
rect 295 1774 301 1826
rect 353 1774 365 1826
rect 417 1774 423 1826
rect 3390 1746 3518 2242
rect 3856 1826 3984 2242
rect 3856 1774 3862 1826
rect 3914 1774 3926 1826
rect 3978 1774 3984 1826
rect 4178 1976 4230 1984
rect 4178 1912 4230 1924
rect 3390 1694 3396 1746
rect 3448 1694 3460 1746
rect 3512 1694 3518 1746
rect 2472 1641 2524 1647
rect 2472 1577 2524 1589
rect 1461 1220 1491 1250
rect 2472 650 2524 1525
rect 4178 1471 4230 1860
rect 4740 1746 4868 2242
tri 5699 1826 5724 1851 se
rect 5724 1826 5776 2832
rect 13439 2844 13445 2896
rect 13497 2844 13503 2896
rect 13439 2832 13503 2844
rect 13439 2780 13445 2832
rect 13497 2780 13503 2832
rect 13439 2777 13503 2780
tri 13439 2765 13451 2777 ne
rect 6167 2442 6219 2448
rect 6167 2378 6219 2390
rect 5648 1774 5654 1826
rect 5706 1774 5718 1826
rect 5770 1774 5776 1826
tri 6136 2261 6167 2292 se
rect 6167 2270 6219 2326
rect 12095 2322 12101 2374
rect 12153 2322 12165 2374
rect 12217 2322 12223 2374
tri 12146 2320 12148 2322 ne
rect 12148 2320 12223 2322
tri 12148 2317 12151 2320 ne
rect 12151 2317 12223 2320
tri 12151 2297 12171 2317 ne
rect 6167 2261 6210 2270
tri 6210 2261 6219 2270 nw
rect 4740 1694 4746 1746
rect 4798 1694 4810 1746
rect 4862 1694 4868 1746
rect 4178 1407 4230 1419
rect 4178 1343 4230 1355
rect 4178 1279 4230 1291
rect 4178 1215 4230 1227
tri 2683 1184 2708 1209 ne
tri 2699 659 2708 668 se
rect 2708 659 2760 1214
rect 4178 1151 4230 1163
tri 2689 649 2699 659 se
rect 2699 649 2760 659
tri 4172 711 4174 713 se
rect 4178 711 4230 1099
rect 4172 659 4178 711
rect 4230 659 4242 711
rect 4294 659 4300 711
tri 4172 657 4174 659 ne
rect 4178 653 4230 659
tri 2683 643 2689 649 se
rect 2689 643 2760 649
rect 2472 586 2524 598
rect 2632 591 2638 643
rect 2690 591 2702 643
rect 2754 591 2760 643
rect 2472 528 2524 534
rect 6136 570 6188 2261
tri 6188 2239 6210 2261 nw
tri 12146 1654 12171 1679 se
rect 12171 1654 12223 2317
rect 13295 2317 13301 2369
rect 13353 2317 13365 2369
rect 13417 2317 13423 2369
rect 13295 1826 13423 2317
rect 13295 1774 13301 1826
rect 13353 1774 13365 1826
rect 13417 1774 13423 1826
tri 13426 1737 13451 1762 se
rect 13451 1737 13503 2777
rect 6216 1648 6268 1654
rect 12095 1602 12101 1654
rect 12153 1602 12165 1654
rect 12217 1602 12223 1654
rect 13375 1621 13381 1737
rect 13497 1621 13503 1737
rect 6216 1584 6268 1596
rect 6216 713 6268 1532
rect 13599 1215 13651 3233
tri 13651 3208 13676 3233 nw
rect 13599 1151 13651 1163
rect 13599 1093 13651 1099
rect 6216 649 6268 661
rect 6216 591 6268 597
rect 15088 835 15408 1644
rect 15088 783 15094 835
rect 15146 783 15158 835
rect 15210 783 15222 835
rect 15274 783 15286 835
rect 15338 783 15350 835
rect 15402 783 15408 835
tri 6188 570 6197 579 sw
rect 15088 570 15408 783
rect 6136 554 6197 570
tri 6197 554 6213 570 sw
rect 6136 502 6142 554
rect 6194 502 6206 554
rect 6258 502 6264 554
rect 15204 454 15408 570
rect 15088 -146 15408 454
rect 15596 -146 15916 1292
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_0
timestamp 1701704242
transform -1 0 12192 0 -1 2892
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_1
timestamp 1701704242
transform -1 0 11554 0 -1 2892
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_2
timestamp 1701704242
transform 1 0 13045 0 -1 3430
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_3
timestamp 1701704242
transform 1 0 14201 0 1 2786
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_4
timestamp 1701704242
transform 1 0 14465 0 1 2786
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_5
timestamp 1701704242
transform 1 0 14641 0 1 2786
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_6
timestamp 1701704242
transform 1 0 6179 0 1 2336
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_7
timestamp 1701704242
transform 1 0 11776 0 1 2786
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_8
timestamp 1701704242
transform 1 0 11952 0 1 2786
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1701704242
transform 0 -1 4224 -1 0 1972
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1701704242
transform -1 0 3816 0 1 2254
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1701704242
transform -1 0 11282 0 1 2712
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_3
timestamp 1701704242
transform -1 0 11282 0 1 2934
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_4
timestamp 1701704242
transform -1 0 4700 0 1 2254
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_5
timestamp 1701704242
transform 0 1 14269 1 0 3244
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_6
timestamp 1701704242
transform 0 -1 13827 1 0 3244
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_7
timestamp 1701704242
transform 0 -1 2529 1 0 540
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_8
timestamp 1701704242
transform 1 0 13937 0 -1 3430
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_9
timestamp 1701704242
transform 1 0 6308 0 1 2356
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_10
timestamp 1701704242
transform 1 0 13571 0 1 2356
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_11
timestamp 1701704242
transform 1 0 12306 0 1 2408
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_12
timestamp 1701704242
transform 1 0 12455 0 1 2334
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_13
timestamp 1701704242
transform 1 0 199 0 1 2254
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_0
timestamp 1701704242
transform 0 -1 14902 -1 0 3192
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_1
timestamp 1701704242
transform 0 -1 12824 -1 0 3192
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_2
timestamp 1701704242
transform 0 -1 12741 -1 0 3192
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_0
timestamp 1701704242
transform -1 0 955 0 -1 2288
box 0 0 1 1
use L1M1_CDNS_52468879185308  L1M1_CDNS_52468879185308_0
timestamp 1701704242
transform 1 0 3249 0 1 2254
box 0 0 1 1
use L1M1_CDNS_52468879185308  L1M1_CDNS_52468879185308_1
timestamp 1701704242
transform 1 0 4765 0 1 2254
box 0 0 1 1
use L1M1_CDNS_52468879185316  L1M1_CDNS_52468879185316_0
timestamp 1701704242
transform 1 0 3899 0 1 2254
box -12 -6 622 40
use L1M1_CDNS_52468879185334  L1M1_CDNS_52468879185334_0
timestamp 1701704242
transform 0 1 11086 -1 0 3192
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_0
timestamp 1701704242
transform 0 -1 4221 1 0 1272
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_1
timestamp 1701704242
transform 0 -1 4221 1 0 665
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_2
timestamp 1701704242
transform 1 0 12790 0 -1 2968
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_3
timestamp 1701704242
transform 1 0 13432 0 1 2403
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_4
timestamp 1701704242
transform 1 0 12788 0 1 2712
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_0
timestamp 1701704242
transform 0 -1 6268 -1 0 1654
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_1
timestamp 1701704242
transform 0 -1 6268 -1 0 719
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_2
timestamp 1701704242
transform 0 -1 2524 -1 0 1647
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_3
timestamp 1701704242
transform 0 -1 347 -1 0 2370
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_4
timestamp 1701704242
transform 0 1 4178 -1 0 1982
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_5
timestamp 1701704242
transform -1 0 12223 0 1 1602
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_6
timestamp 1701704242
transform -1 0 3518 0 1 1694
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_7
timestamp 1701704242
transform -1 0 3518 0 1 2242
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_8
timestamp 1701704242
transform -1 0 5776 0 -1 2900
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_9
timestamp 1701704242
transform -1 0 3984 0 -1 1826
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_10
timestamp 1701704242
transform -1 0 2760 0 -1 643
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_11
timestamp 1701704242
transform 0 -1 13913 1 0 3233
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_12
timestamp 1701704242
transform 0 -1 6219 1 0 2320
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_13
timestamp 1701704242
transform 0 -1 2524 1 0 528
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_14
timestamp 1701704242
transform 0 -1 13651 1 0 1093
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_15
timestamp 1701704242
transform 1 0 295 0 -1 1826
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_16
timestamp 1701704242
transform 1 0 5648 0 1 1774
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_17
timestamp 1701704242
transform 1 0 13295 0 1 1774
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_18
timestamp 1701704242
transform 1 0 6136 0 1 502
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_19
timestamp 1701704242
transform 1 0 12095 0 1 2322
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_20
timestamp 1701704242
transform 1 0 3856 0 1 2242
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_21
timestamp 1701704242
transform 1 0 13295 0 1 2317
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_22
timestamp 1701704242
transform 1 0 4740 0 1 1694
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_23
timestamp 1701704242
transform 1 0 4740 0 1 2242
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_0
timestamp 1701704242
transform 0 1 3698 1 0 2476
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_1
timestamp 1701704242
transform 0 1 4596 1 0 2476
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_0
timestamp 1701704242
transform -1 0 13503 0 -1 1737
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_1
timestamp 1701704242
transform 0 1 15088 1 0 448
box 0 0 1 1
use M1M2_CDNS_52468879185200  M1M2_CDNS_52468879185200_0
timestamp 1701704242
transform 1 0 -11 0 -1 2214
box 0 0 1 1
use M1M2_CDNS_52468879185202  M1M2_CDNS_52468879185202_0
timestamp 1701704242
transform 1 0 15088 0 -1 835
box 0 0 1 1
use M1M2_CDNS_52468879185204  M1M2_CDNS_52468879185204_0
timestamp 1701704242
transform 0 -1 4230 1 0 1093
box 0 0 1 1
use M1M2_CDNS_52468879185209  M1M2_CDNS_52468879185209_0
timestamp 1701704242
transform 1 0 -11 0 -1 3204
box 0 0 128 244
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_0
timestamp 1701704242
transform 0 1 3698 1 0 2242
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_1
timestamp 1701704242
transform 0 1 4596 1 0 2242
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_2
timestamp 1701704242
transform 1 0 13439 0 1 2780
box 0 0 1 1
use M1M2_CDNS_52468879185970  M1M2_CDNS_52468879185970_0
timestamp 1701704242
transform 0 1 4178 1 0 653
box 0 0 1 1
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_0
timestamp 1701704242
transform 1 0 13679 0 1 876
box 0 0 192 180
use M1M2_CDNS_524688791851077  M1M2_CDNS_524688791851077_0
timestamp 1701704242
transform 1 0 15596 0 -1 1278
box 0 0 320 180
use M1M2_CDNS_524688791851077  M1M2_CDNS_524688791851077_1
timestamp 1701704242
transform 1 0 15088 0 -1 1824
box 0 0 320 180
use sky130_fd_io__sio_com_ctl_ls  sky130_fd_io__sio_com_ctl_ls_0
timestamp 1701704242
transform 1 0 2102 0 -1 2304
box -91 0 2150 2319
use sky130_fd_io__sio_com_octl_tsg4  sky130_fd_io__sio_com_octl_tsg4_0
timestamp 1701704242
transform 1 0 0 0 1 0
box -84 -15 11187 3738
use sky130_fd_io__sio_hvsbt_diff_space  sky130_fd_io__sio_hvsbt_diff_space_0
timestamp 1701704242
transform 1 0 11969 0 1 2335
box 0 0 1 1
use sky130_fd_io__sio_hvsbt_diff_space  sky130_fd_io__sio_hvsbt_diff_space_1
timestamp 1701704242
transform 1 0 14108 0 1 2335
box 0 0 1 1
use sky130_fd_io__sio_hvsbt_diff_space  sky130_fd_io__sio_hvsbt_diff_space_2
timestamp 1701704242
transform 1 0 13238 0 1 2335
box 0 0 1 1
use sky130_fd_io__sio_hvsbt_endcap  sky130_fd_io__sio_hvsbt_endcap_0
timestamp 1701704242
transform -1 0 14885 0 1 2335
box -84 93 164 1337
use sky130_fd_io__sio_hvsbt_endcap  sky130_fd_io__sio_hvsbt_endcap_1
timestamp 1701704242
transform -1 0 12724 0 1 2335
box -84 93 164 1337
use sky130_fd_io__sio_hvsbt_inv_x1  sky130_fd_io__sio_hvsbt_inv_x1_0
timestamp 1701704242
transform -1 0 12255 0 1 2335
box -107 21 267 1369
use sky130_fd_io__sio_hvsbt_inv_x1  sky130_fd_io__sio_hvsbt_inv_x1_1
timestamp 1701704242
transform -1 0 14394 0 1 2335
box -107 21 267 1369
use sky130_fd_io__sio_hvsbt_inv_x2  sky130_fd_io__sio_hvsbt_inv_x2_0
timestamp 1701704242
transform -1 0 14746 0 1 2335
box -107 21 459 1369
use sky130_fd_io__sio_hvsbt_inv_x2  sky130_fd_io__sio_hvsbt_inv_x2_1
timestamp 1701704242
transform 1 0 12886 0 1 2335
box -107 21 459 1369
use sky130_fd_io__sio_hvsbt_inv_x2  sky130_fd_io__sio_hvsbt_inv_x2_2
timestamp 1701704242
transform 1 0 11265 0 1 2335
box -107 21 459 1369
use sky130_fd_io__sio_hvsbt_nand2  sky130_fd_io__sio_hvsbt_nand2_0
timestamp 1701704242
transform 1 0 11617 0 1 2335
box -107 21 459 1369
use sky130_fd_io__sio_hvsbt_nand2  sky130_fd_io__sio_hvsbt_nand2_1
timestamp 1701704242
transform 1 0 12255 0 1 2335
box -107 21 459 1369
use sky130_fd_io__sio_hvsbt_nor  sky130_fd_io__sio_hvsbt_nor_0
timestamp 1701704242
transform -1 0 13728 0 1 2335
box -107 21 487 1369
use sky130_fd_io__sio_hvsbt_nor  sky130_fd_io__sio_hvsbt_nor_1
timestamp 1701704242
transform 1 0 13728 0 1 2335
box -107 21 487 1369
<< labels >>
flabel comment s 5798 1800 5798 1800 0 FreeSans 400 0 0 0 vreg_en_h_n
flabel comment s 11940 2879 11940 2879 0 FreeSans 400 0 0 0 vreg_puen2_n
flabel comment s 11608 2809 11608 2809 0 FreeSans 200 0 0 0 puen_h2_n
flabel comment s 12816 2428 12816 2428 0 FreeSans 200 0 0 0 puen_2or1_h
flabel comment s 13065 3717 13065 3717 0 FreeSans 200 0 0 0 oe_h
flabel metal1 s 4156 2254 4190 2288 3 FreeSans 400 0 0 0 od_h
port 3 nsew
flabel metal1 s 3208 2248 3249 2294 7 FreeSans 400 0 0 0 hld_i_h_n
port 4 nsew
flabel metal1 s 12263 2807 12263 2807 0 FreeSans 200 0 0 0 vreg_puen2
flabel metal1 s 12003 2427 12003 2427 0 FreeSans 400 0 0 0 puen_2or1_h
flabel metal1 s 13296 3418 13296 3418 0 FreeSans 200 0 0 0 oe_i_h_n
flabel metal1 s 14368 2837 14368 2837 0 FreeSans 200 0 0 0 oe_hs_i_h_n
flabel metal1 s 13688 3332 13688 3332 0 FreeSans 200 0 0 0 n<1>
flabel metal1 s 12390 1602 12434 1654 7 FreeSans 400 0 0 0 vreg_en_h
port 20 nsew
flabel metal1 s 16030 1093 16040 1295 7 FreeSans 200 0 0 0 vpb_ka
port 6 nsew
flabel metal1 s 16030 1624 16040 1826 7 FreeSans 200 0 0 0 vpwr_ka
port 2 nsew
flabel metal1 s 117 2706 129 2752 0 FreeSans 200 0 0 0 vgnd
port 10 nsew
flabel metal1 s 4071 1221 4106 1255 0 FreeSans 200 0 0 0 vreg_en
port 7 nsew
flabel metal1 s 2078 218 2127 420 0 FreeSans 200 0 0 0 vpwr
port 8 nsew
flabel metal1 s -2 72 16 190 0 FreeSans 200 0 0 0 vpb
port 9 nsew
flabel metal1 s 117 2476 129 2678 0 FreeSans 200 0 0 0 vgnd
port 10 nsew
flabel metal1 s 117 3002 129 3204 0 FreeSans 200 0 0 0 vcc_io
port 11 nsew
flabel metal1 s 1747 1607 1781 1641 0 FreeSans 400 0 0 0 slow_h_n
port 5 nsew
flabel metal1 s 98 1221 132 1255 0 FreeSans 200 0 0 0 slow
port 12 nsew
flabel metal1 s 5399 795 5433 829 0 FreeSans 400 0 0 0 hld_i_vpwr
port 13 nsew
flabel metal1 s 363 2404 397 2438 0 FreeSans 400 0 0 0 dm_h_n<2>
port 14 nsew
flabel metal1 s 223 3501 257 3535 3 FreeSans 400 0 0 0 dm_h_n<1>
port 15 nsew
flabel metal1 s 563 3310 597 3344 0 FreeSans 400 0 0 0 dm_h_n<0>
port 16 nsew
flabel metal1 s 3399 2378 3434 2412 0 FreeSans 400 0 0 0 dm_h<2>
port 17 nsew
flabel metal1 s 2869 3396 2903 3430 3 FreeSans 400 0 0 0 dm_h<1>
port 18 nsew
flabel metal1 s 2402 3618 2436 3652 0 FreeSans 400 0 0 0 dm_h<0>
port 19 nsew
flabel locali s 8839 2548 8873 2592 0 FreeSans 200 0 0 0 pden_h_n<2>
port 21 nsew
flabel locali s 11424 3555 11458 3604 0 FreeSans 200 0 0 0 puen_h<2>
port 22 nsew
flabel locali s 7277 3510 7311 3550 0 FreeSans 200 0 0 0 puen_h<1>
port 23 nsew
flabel locali s 5473 2456 5507 2506 0 FreeSans 200 0 0 0 puen_h<0>
port 24 nsew
flabel locali s 10061 2511 10095 2555 0 FreeSans 200 0 0 0 pden_h_n<1>
port 25 nsew
flabel locali s 10413 2508 10447 2550 0 FreeSans 200 0 0 0 pden_h_n<0>
port 26 nsew
flabel locali s 14553 2506 14587 2556 0 FreeSans 200 0 0 0 oe_hs_h
port 27 nsew
flabel locali s 13133 3654 13167 3704 0 FreeSans 200 0 0 0 oe_h
port 28 nsew
flabel metal2 s 1461 1220 1491 1250 0 FreeSans 200 0 0 0 slow_h
port 29 nsew
<< properties >>
string GDS_END 87723272
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 87702264
string path 104.300 17.125 107.500 17.125 
<< end >>
