magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -266 -66 914 666
<< mvpmos >>
rect 0 0 120 600
rect 176 0 296 600
rect 352 0 472 600
rect 528 0 648 600
<< mvpdiff >>
rect -50 0 0 600
rect 648 0 698 600
<< poly >>
rect 0 600 120 632
rect 0 -32 120 0
rect 176 600 296 632
rect 176 -32 296 0
rect 352 600 472 632
rect 352 -32 472 0
rect 528 600 648 632
rect 528 -32 648 0
<< locali >>
rect -113 -4 -11 550
rect 131 -4 165 538
rect 307 -4 341 538
rect 483 -4 517 538
rect 659 -4 761 550
use DFL1sd2_CDNS_5246887918535  DFL1sd2_CDNS_5246887918535_0
timestamp 1701704242
transform 1 0 472 0 1 0
box -36 -36 92 636
use DFL1sd2_CDNS_5246887918535  DFL1sd2_CDNS_5246887918535_1
timestamp 1701704242
transform 1 0 296 0 1 0
box -36 -36 92 636
use DFL1sd2_CDNS_5246887918535  DFL1sd2_CDNS_5246887918535_2
timestamp 1701704242
transform 1 0 120 0 1 0
box -36 -36 92 636
use hvDFTPL1s_CDNS_52468879185914  hvDFTPL1s_CDNS_52468879185914_0
timestamp 1701704242
transform -1 0 0 0 1 0
box -36 -36 236 636
use hvDFTPL1s_CDNS_52468879185914  hvDFTPL1s_CDNS_52468879185914_1
timestamp 1701704242
transform 1 0 648 0 1 0
box -36 -36 236 636
<< labels >>
flabel comment s -62 273 -62 273 0 FreeSans 300 0 0 0 S
flabel comment s 148 267 148 267 0 FreeSans 300 0 0 0 D
flabel comment s 324 267 324 267 0 FreeSans 300 0 0 0 S
flabel comment s 500 267 500 267 0 FreeSans 300 0 0 0 D
flabel comment s 710 273 710 273 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 80821178
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 80818668
<< end >>
