magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< metal2 >>
rect 0 8385 376 8394
rect 0 0 376 9
<< via2 >>
rect 0 9 376 8385
<< metal3 >>
rect -5 8385 381 8390
rect -5 9 0 8385
rect 376 9 381 8385
rect -5 4 381 9
<< properties >>
string GDS_END 93527990
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 93494258
<< end >>
