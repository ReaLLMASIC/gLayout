magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< nwell >>
rect 0 1464 92 2596
<< pwell >>
rect 20 10 110 1386
<< mvpsubdiff >>
rect 46 1323 84 1360
rect 46 1289 48 1323
rect 82 1289 84 1323
rect 46 1255 84 1289
rect 46 1221 48 1255
rect 82 1221 84 1255
rect 46 1187 84 1221
rect 46 1153 48 1187
rect 82 1153 84 1187
rect 46 1119 84 1153
rect 46 1085 48 1119
rect 82 1085 84 1119
rect 46 1051 84 1085
rect 46 1017 48 1051
rect 82 1017 84 1051
rect 46 983 84 1017
rect 46 949 48 983
rect 82 949 84 983
rect 46 915 84 949
rect 46 881 48 915
rect 82 881 84 915
rect 46 847 84 881
rect 46 813 48 847
rect 82 813 84 847
rect 46 779 84 813
rect 46 745 48 779
rect 82 745 84 779
rect 46 711 84 745
rect 46 677 48 711
rect 82 677 84 711
rect 46 643 84 677
rect 46 609 48 643
rect 82 609 84 643
rect 46 575 84 609
rect 46 541 48 575
rect 82 541 84 575
rect 46 507 84 541
rect 46 473 48 507
rect 82 473 84 507
rect 46 439 84 473
rect 46 405 48 439
rect 82 405 84 439
rect 46 371 84 405
rect 46 337 48 371
rect 82 337 84 371
rect 46 303 84 337
rect 46 269 48 303
rect 82 269 84 303
rect 46 235 84 269
rect 46 201 48 235
rect 82 201 84 235
rect 46 167 84 201
rect 46 133 48 167
rect 82 133 84 167
rect 46 99 84 133
rect 46 65 48 99
rect 82 65 84 99
rect 46 36 84 65
<< mvnsubdiff >>
rect 66 2485 104 2530
rect 66 2451 68 2485
rect 102 2451 104 2485
rect 66 2417 104 2451
rect 66 2383 68 2417
rect 102 2383 104 2417
rect 66 2349 104 2383
rect 66 2315 68 2349
rect 102 2315 104 2349
rect 66 2281 104 2315
rect 66 2247 68 2281
rect 102 2247 104 2281
rect 66 2213 104 2247
rect 66 2179 68 2213
rect 102 2179 104 2213
rect 66 2145 104 2179
rect 66 2111 68 2145
rect 102 2111 104 2145
rect 66 2077 104 2111
rect 66 2043 68 2077
rect 102 2043 104 2077
rect 66 2009 104 2043
rect 66 1975 68 2009
rect 102 1975 104 2009
rect 66 1941 104 1975
rect 66 1907 68 1941
rect 102 1907 104 1941
rect 66 1873 104 1907
rect 66 1839 68 1873
rect 102 1839 104 1873
rect 66 1798 104 1839
rect 66 1764 68 1798
rect 102 1764 104 1798
rect 66 1730 104 1764
rect 66 1696 68 1730
rect 102 1696 104 1730
rect 66 1662 104 1696
rect 66 1628 68 1662
rect 102 1628 104 1662
rect 66 1594 104 1628
rect 66 1560 68 1594
rect 102 1560 104 1594
rect 66 1530 104 1560
<< mvpsubdiffcont >>
rect 48 1289 82 1323
rect 48 1221 82 1255
rect 48 1153 82 1187
rect 48 1085 82 1119
rect 48 1017 82 1051
rect 48 949 82 983
rect 48 881 82 915
rect 48 813 82 847
rect 48 745 82 779
rect 48 677 82 711
rect 48 609 82 643
rect 48 541 82 575
rect 48 473 82 507
rect 48 405 82 439
rect 48 337 82 371
rect 48 269 82 303
rect 48 201 82 235
rect 48 133 82 167
rect 48 65 82 99
<< mvnsubdiffcont >>
rect 68 2451 102 2485
rect 68 2383 102 2417
rect 68 2315 102 2349
rect 68 2247 102 2281
rect 68 2179 102 2213
rect 68 2111 102 2145
rect 68 2043 102 2077
rect 68 1975 102 2009
rect 68 1907 102 1941
rect 68 1839 102 1873
rect 68 1764 102 1798
rect 68 1696 102 1730
rect 68 1628 102 1662
rect 68 1560 102 1594
<< poly >>
rect 211 2612 683 2632
rect 211 2578 240 2612
rect 274 2578 308 2612
rect 342 2578 376 2612
rect 410 2578 444 2612
rect 478 2578 512 2612
rect 546 2578 580 2612
rect 614 2578 683 2612
rect 211 2556 683 2578
rect 739 2612 881 2632
rect 739 2578 759 2612
rect 793 2578 827 2612
rect 861 2578 881 2612
rect 739 2556 881 2578
rect 1008 2536 1074 2552
rect 1008 2502 1024 2536
rect 1058 2502 1074 2536
rect 1008 2468 1074 2502
rect 1008 2434 1024 2468
rect 1058 2434 1074 2468
rect 1008 2418 1074 2434
rect 1170 2536 1236 2552
rect 1170 2502 1186 2536
rect 1220 2502 1236 2536
rect 1170 2468 1236 2502
rect 1170 2434 1186 2468
rect 1220 2434 1236 2468
rect 1170 2418 1236 2434
rect 1008 1634 1074 1650
rect 1008 1600 1024 1634
rect 1058 1600 1074 1634
rect 1008 1566 1074 1600
rect 1008 1532 1024 1566
rect 1058 1532 1074 1566
rect 1008 1516 1074 1532
rect 211 1386 311 1504
rect 353 1442 555 1462
rect 353 1408 369 1442
rect 403 1408 437 1442
rect 471 1408 505 1442
rect 539 1408 555 1442
rect 353 1386 555 1408
rect 609 1442 811 1462
rect 609 1408 625 1442
rect 659 1408 693 1442
rect 727 1408 761 1442
rect 795 1408 811 1442
rect 609 1386 811 1408
rect 211 1029 311 1034
rect 177 1013 311 1029
rect 177 979 193 1013
rect 227 979 261 1013
rect 295 979 311 1013
rect 177 963 311 979
rect 211 958 311 963
rect 853 1013 995 1034
rect 853 979 869 1013
rect 903 979 937 1013
rect 971 979 995 1013
rect 853 958 995 979
rect 211 476 311 606
rect 353 584 555 606
rect 353 550 369 584
rect 403 550 437 584
rect 471 550 505 584
rect 539 550 555 584
rect 353 530 555 550
rect 609 584 811 606
rect 609 550 625 584
rect 659 550 693 584
rect 727 550 761 584
rect 795 550 811 584
rect 609 530 811 550
rect 853 476 953 606
rect 211 400 1011 476
rect 1170 234 1236 250
rect 211 146 1011 222
rect 1170 200 1186 234
rect 1220 200 1236 234
rect 1170 166 1236 200
rect 1170 132 1186 166
rect 1220 132 1236 166
rect 1170 116 1236 132
<< polycont >>
rect 240 2578 274 2612
rect 308 2578 342 2612
rect 376 2578 410 2612
rect 444 2578 478 2612
rect 512 2578 546 2612
rect 580 2578 614 2612
rect 759 2578 793 2612
rect 827 2578 861 2612
rect 1024 2502 1058 2536
rect 1024 2434 1058 2468
rect 1186 2502 1220 2536
rect 1186 2434 1220 2468
rect 1024 1600 1058 1634
rect 1024 1532 1058 1566
rect 369 1408 403 1442
rect 437 1408 471 1442
rect 505 1408 539 1442
rect 625 1408 659 1442
rect 693 1408 727 1442
rect 761 1408 795 1442
rect 193 979 227 1013
rect 261 979 295 1013
rect 869 979 903 1013
rect 937 979 971 1013
rect 369 550 403 584
rect 437 550 471 584
rect 505 550 539 584
rect 625 550 659 584
rect 693 550 727 584
rect 761 550 795 584
rect 1186 200 1220 234
rect 1186 132 1220 166
<< locali >>
rect 224 2578 240 2612
rect 274 2578 308 2612
rect 346 2578 376 2612
rect 410 2578 444 2612
rect 478 2578 512 2612
rect 546 2578 580 2612
rect 614 2578 630 2612
rect 743 2578 759 2612
rect 803 2578 827 2612
rect 875 2578 877 2612
rect 1008 2502 1024 2536
rect 1058 2502 1186 2536
rect 1220 2502 1240 2536
rect 68 2485 102 2501
rect 68 2417 102 2451
rect 1008 2468 1240 2502
rect 1008 2434 1024 2468
rect 1058 2434 1186 2468
rect 1220 2434 1240 2468
rect 68 2349 102 2383
rect 68 2281 102 2315
rect 68 2213 102 2247
rect 68 2145 102 2179
rect 68 2077 102 2111
rect 68 2009 102 2043
rect 68 1941 102 1975
rect 68 1873 102 1907
rect 1170 1840 1236 1914
rect 68 1798 102 1839
rect 200 1806 238 1840
rect 518 1806 556 1840
rect 828 1806 866 1840
rect 1024 1806 1062 1840
rect 1096 1806 1236 1840
rect 68 1754 102 1764
rect 68 1682 102 1696
rect 68 1610 102 1628
rect 342 1688 376 1726
rect 342 1616 376 1654
rect 694 1688 728 1726
rect 694 1616 728 1654
rect 1008 1634 1074 1806
rect 1008 1600 1024 1634
rect 1058 1600 1074 1634
rect 68 1538 102 1560
rect 1008 1566 1074 1600
rect 1008 1532 1024 1566
rect 1058 1532 1074 1566
rect 353 1408 369 1442
rect 403 1408 437 1442
rect 471 1408 505 1442
rect 539 1408 555 1442
rect 609 1408 625 1442
rect 659 1408 693 1442
rect 727 1408 761 1442
rect 795 1408 811 1442
rect 48 1323 82 1352
rect 48 1255 82 1289
rect 48 1187 82 1206
rect 48 1119 82 1134
rect 48 1051 82 1062
rect 48 983 82 1017
rect 48 915 82 949
rect 48 847 82 881
rect 48 779 82 813
rect 48 711 82 716
rect 48 643 82 644
rect 116 1094 200 1364
rect 564 1162 598 1200
rect 116 898 150 1094
rect 564 1090 598 1128
rect 964 1094 1059 1364
rect 193 1013 295 1029
rect 227 1006 261 1013
rect 869 1013 971 1029
rect 234 979 261 1006
rect 193 972 200 979
rect 234 972 272 979
rect 903 979 937 1013
rect 193 963 295 972
rect 901 970 939 979
rect 869 963 971 970
rect 1025 898 1059 1094
rect 1170 972 1236 1806
rect 1152 938 1190 972
rect 1224 938 1236 972
rect 116 830 200 898
rect 964 830 1059 898
rect 1170 830 1236 836
rect 116 796 178 830
rect 212 796 250 830
rect 912 796 950 830
rect 984 796 1059 830
rect 1152 796 1190 830
rect 1224 796 1236 830
rect 116 628 200 796
rect 564 678 598 716
rect 964 628 1059 796
rect 48 575 82 609
rect 353 550 369 584
rect 403 550 437 584
rect 471 550 505 584
rect 539 550 555 584
rect 609 550 625 584
rect 659 550 693 584
rect 727 550 761 584
rect 795 550 811 584
rect 48 507 82 541
rect 48 439 82 473
rect 257 422 295 456
rect 48 371 82 405
rect 48 303 82 337
rect 48 235 82 269
rect 48 167 82 201
rect 48 99 82 100
rect 166 98 200 286
rect 1022 268 1056 306
rect 1170 234 1236 796
rect 901 180 939 214
rect 1170 200 1186 234
rect 1220 200 1236 234
rect 1170 166 1236 200
rect 1170 132 1186 166
rect 1220 132 1236 166
rect 48 62 82 65
rect 1022 62 1056 100
<< viali >>
rect 240 2578 274 2612
rect 312 2578 342 2612
rect 342 2578 346 2612
rect 769 2578 793 2612
rect 793 2578 803 2612
rect 841 2578 861 2612
rect 861 2578 875 2612
rect 166 1806 200 1840
rect 238 1806 272 1840
rect 484 1806 518 1840
rect 556 1806 590 1840
rect 794 1806 828 1840
rect 866 1806 900 1840
rect 990 1806 1024 1840
rect 1062 1806 1096 1840
rect 68 1730 102 1754
rect 68 1720 102 1730
rect 68 1662 102 1682
rect 68 1648 102 1662
rect 68 1594 102 1610
rect 68 1576 102 1594
rect 342 1726 376 1760
rect 342 1654 376 1688
rect 342 1582 376 1616
rect 694 1726 728 1760
rect 694 1654 728 1688
rect 694 1582 728 1616
rect 48 1221 82 1240
rect 48 1206 82 1221
rect 48 1153 82 1168
rect 48 1134 82 1153
rect 48 1085 82 1096
rect 48 1062 82 1085
rect 48 745 82 750
rect 48 716 82 745
rect 48 677 82 678
rect 48 644 82 677
rect 564 1200 598 1234
rect 564 1128 598 1162
rect 564 1056 598 1090
rect 200 979 227 1006
rect 227 979 234 1006
rect 272 979 295 1006
rect 295 979 306 1006
rect 200 972 234 979
rect 272 972 306 979
rect 867 979 869 1004
rect 869 979 901 1004
rect 939 979 971 1004
rect 971 979 973 1004
rect 867 970 901 979
rect 939 970 973 979
rect 1118 938 1152 972
rect 1190 938 1224 972
rect 178 796 212 830
rect 250 796 284 830
rect 878 796 912 830
rect 950 796 984 830
rect 1118 796 1152 830
rect 1190 796 1224 830
rect 564 716 598 750
rect 564 644 598 678
rect 223 422 257 456
rect 295 422 329 456
rect 1022 306 1056 340
rect 48 133 82 134
rect 48 100 82 133
rect 1022 234 1056 268
rect 867 180 901 214
rect 939 180 973 214
rect 1022 100 1056 134
rect 48 28 82 62
rect 1022 28 1056 62
<< metal1 >>
rect 211 2616 391 2622
rect 263 2612 275 2616
rect 327 2612 339 2616
rect 274 2578 275 2612
rect 263 2564 275 2578
rect 327 2564 339 2578
rect 211 2558 391 2564
rect 757 2616 933 2622
rect 757 2612 817 2616
rect 869 2612 881 2616
rect 757 2578 769 2612
rect 803 2578 817 2612
rect 875 2578 881 2612
rect 757 2564 817 2578
rect 869 2564 881 2578
rect 757 2558 933 2564
rect 1013 1922 1065 1928
tri 985 1846 1013 1874 se
rect 1013 1858 1065 1870
rect 0 1840 1013 1846
tri 1065 1846 1093 1874 sw
rect 1065 1840 1236 1846
rect 0 1806 166 1840
rect 200 1806 238 1840
rect 272 1806 484 1840
rect 518 1806 556 1840
rect 590 1806 794 1840
rect 828 1806 866 1840
rect 900 1806 990 1840
rect 1096 1806 1236 1840
rect 0 1800 1236 1806
rect 0 1760 1284 1772
rect 0 1754 342 1760
rect 0 1720 68 1754
rect 102 1726 342 1754
rect 376 1726 694 1760
rect 728 1726 1284 1760
rect 102 1720 1284 1726
rect 0 1688 1284 1720
rect 0 1682 342 1688
rect 0 1648 68 1682
rect 102 1654 342 1682
rect 376 1654 694 1688
rect 728 1654 1284 1688
rect 102 1648 1284 1654
rect 0 1616 1284 1648
rect 0 1610 342 1616
rect 0 1576 68 1610
rect 102 1582 342 1610
rect 376 1582 694 1616
rect 728 1582 1284 1616
rect 102 1576 1284 1582
rect 0 1570 1284 1576
rect 0 1240 1284 1246
rect 0 1206 48 1240
rect 82 1234 1284 1240
rect 82 1206 564 1234
rect 0 1200 564 1206
rect 598 1200 1111 1234
rect 0 1182 1111 1200
rect 1163 1182 1284 1234
rect 0 1170 1284 1182
rect 0 1168 1111 1170
rect 0 1134 48 1168
rect 82 1162 1111 1168
rect 82 1134 564 1162
rect 0 1128 564 1134
rect 598 1128 1111 1162
rect 0 1118 1111 1128
rect 1163 1118 1284 1170
rect 0 1106 1284 1118
rect 0 1096 1111 1106
rect 0 1062 48 1096
rect 82 1090 1111 1096
rect 82 1062 564 1090
rect 0 1056 564 1062
rect 598 1056 1111 1090
rect 0 1054 1111 1056
rect 1163 1054 1284 1106
rect 0 1044 1284 1054
rect 188 1006 217 1016
rect 269 1006 281 1016
rect 188 972 200 1006
rect 269 972 272 1006
rect 333 1004 985 1016
rect 188 964 217 972
rect 269 964 281 972
rect 333 970 867 1004
rect 901 970 939 1004
rect 973 970 985 1004
rect 333 964 985 970
rect 1106 972 1236 978
rect 1106 938 1118 972
rect 1152 938 1190 972
rect 1224 938 1236 972
rect 1106 932 1236 938
tri 1156 904 1184 932 ne
rect 1184 904 1236 932
rect 1185 902 1235 903
rect 1184 866 1236 902
rect 1185 865 1235 866
tri 1156 836 1184 864 se
rect 1184 836 1236 864
rect 166 830 1236 836
rect 166 796 178 830
rect 212 796 250 830
rect 284 796 878 830
rect 912 796 950 830
rect 984 796 1118 830
rect 1152 796 1190 830
rect 1224 796 1236 830
rect 166 790 1236 796
rect 0 754 1284 762
rect 0 750 1111 754
rect 0 716 48 750
rect 82 716 564 750
rect 598 716 1111 750
rect 0 702 1111 716
rect 1163 702 1284 754
rect 0 690 1284 702
rect 0 678 1111 690
rect 0 644 48 678
rect 82 644 564 678
rect 598 644 1111 678
rect 0 638 1111 644
rect 1163 638 1284 690
rect 0 632 1284 638
rect 211 418 217 470
rect 269 418 281 470
rect 333 418 341 470
rect 211 416 341 418
rect 1013 340 1065 352
rect 933 296 985 302
tri 919 234 933 248 se
rect 933 234 985 244
tri 905 220 919 234 se
rect 919 232 985 234
rect 919 220 933 232
rect 855 214 933 220
rect 1013 276 1065 288
rect 1013 218 1065 224
rect 855 180 867 214
rect 901 180 933 214
rect 855 174 985 180
rect 42 140 1169 146
rect 42 134 1111 140
rect 42 100 48 134
rect 82 100 1022 134
rect 1056 100 1111 134
rect 42 88 1111 100
rect 1163 88 1169 140
rect 42 76 1169 88
rect 42 62 1111 76
rect 42 28 48 62
rect 82 28 1022 62
rect 1056 28 1111 62
rect 42 24 1111 28
rect 1163 24 1169 76
rect 42 16 1169 24
<< rmetal1 >>
rect 1184 903 1236 904
rect 1184 902 1185 903
rect 1235 902 1236 903
rect 1184 865 1185 866
rect 1235 865 1236 866
rect 1184 864 1236 865
<< via1 >>
rect 211 2612 263 2616
rect 275 2612 327 2616
rect 339 2612 391 2616
rect 211 2578 240 2612
rect 240 2578 263 2612
rect 275 2578 312 2612
rect 312 2578 327 2612
rect 339 2578 346 2612
rect 346 2578 391 2612
rect 211 2564 263 2578
rect 275 2564 327 2578
rect 339 2564 391 2578
rect 817 2612 869 2616
rect 817 2578 841 2612
rect 841 2578 869 2612
rect 817 2564 869 2578
rect 881 2564 933 2616
rect 1013 1870 1065 1922
rect 1013 1840 1065 1858
rect 1013 1806 1024 1840
rect 1024 1806 1062 1840
rect 1062 1806 1065 1840
rect 1111 1182 1163 1234
rect 1111 1118 1163 1170
rect 1111 1054 1163 1106
rect 217 1006 269 1016
rect 281 1006 333 1016
rect 217 972 234 1006
rect 234 972 269 1006
rect 281 972 306 1006
rect 306 972 333 1006
rect 217 964 269 972
rect 281 964 333 972
rect 1111 702 1163 754
rect 1111 638 1163 690
rect 217 456 269 470
rect 217 422 223 456
rect 223 422 257 456
rect 257 422 269 456
rect 217 418 269 422
rect 281 456 333 470
rect 281 422 295 456
rect 295 422 329 456
rect 329 422 333 456
rect 281 418 333 422
rect 1013 306 1022 340
rect 1022 306 1056 340
rect 1056 306 1065 340
rect 933 244 985 296
rect 933 214 985 232
rect 1013 288 1065 306
rect 1013 268 1065 276
rect 1013 234 1022 268
rect 1022 234 1056 268
rect 1056 234 1065 268
rect 1013 224 1065 234
rect 933 180 939 214
rect 939 180 973 214
rect 973 180 985 214
rect 1111 88 1163 140
rect 1111 24 1163 76
<< metal2 >>
rect 211 2616 391 2622
rect 263 2564 275 2616
rect 327 2564 339 2616
rect 211 2558 391 2564
rect 817 2616 985 2622
rect 869 2564 881 2616
rect 933 2564 985 2616
rect 817 2558 985 2564
rect 211 1016 263 2558
tri 263 2530 291 2558 nw
tri 905 2530 933 2558 ne
tri 263 1016 291 1044 sw
rect 211 964 217 1016
rect 269 964 281 1016
rect 333 964 339 1016
rect 211 470 263 964
tri 263 936 291 964 nw
tri 263 470 291 498 sw
rect 211 418 217 470
rect 269 418 281 470
rect 333 418 339 470
rect 933 296 985 2558
rect 933 232 985 244
rect 1013 1922 1065 1928
rect 1013 1858 1065 1870
rect 1013 340 1065 1806
rect 1013 276 1065 288
rect 1013 218 1065 224
rect 1105 1234 1169 1246
rect 1105 1182 1111 1234
rect 1163 1182 1169 1234
rect 1105 1170 1169 1182
rect 1105 1118 1111 1170
rect 1163 1118 1169 1170
rect 1105 1106 1169 1118
rect 1105 1054 1111 1106
rect 1163 1054 1169 1106
rect 1105 754 1169 1054
rect 1105 702 1111 754
rect 1163 702 1169 754
rect 1105 690 1169 702
rect 1105 638 1111 690
rect 1163 638 1169 690
rect 933 174 985 180
rect 1105 140 1169 638
rect 1105 88 1111 140
rect 1163 88 1169 140
rect 1105 76 1169 88
rect 1105 24 1111 76
rect 1163 24 1169 76
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1701704242
transform -1 0 984 0 1 796
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1701704242
transform -1 0 284 0 1 796
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1701704242
transform -1 0 875 0 -1 2612
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_3
timestamp 1701704242
transform -1 0 973 0 -1 214
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_4
timestamp 1701704242
transform 0 1 48 1 0 644
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_5
timestamp 1701704242
transform 0 1 564 1 0 644
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_6
timestamp 1701704242
transform 0 1 1022 1 0 234
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_7
timestamp 1701704242
transform 0 1 48 1 0 28
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_8
timestamp 1701704242
transform 0 -1 1056 1 0 28
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_9
timestamp 1701704242
transform 1 0 223 0 -1 456
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_10
timestamp 1701704242
transform 1 0 1118 0 -1 830
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_11
timestamp 1701704242
transform 1 0 990 0 -1 1840
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_12
timestamp 1701704242
transform 1 0 1118 0 -1 972
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_13
timestamp 1701704242
transform 1 0 240 0 1 2578
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_14
timestamp 1701704242
transform 1 0 867 0 1 970
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_15
timestamp 1701704242
transform 1 0 166 0 1 1806
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_16
timestamp 1701704242
transform 1 0 484 0 1 1806
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_17
timestamp 1701704242
transform 1 0 794 0 1 1806
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_18
timestamp 1701704242
transform 1 0 200 0 1 972
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_0
timestamp 1701704242
transform 0 -1 376 -1 0 1760
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_1
timestamp 1701704242
transform 0 -1 728 -1 0 1760
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_2
timestamp 1701704242
transform 0 1 564 -1 0 1234
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_0
timestamp 1701704242
transform -1 0 82 0 1 1062
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_1
timestamp 1701704242
transform 1 0 68 0 1 1576
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_0
timestamp 1701704242
transform 0 1 1013 1 0 1800
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_1
timestamp 1701704242
transform 0 1 933 1 0 174
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_2
timestamp 1701704242
transform 0 -1 1065 1 0 218
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_3
timestamp 1701704242
transform 1 0 211 0 1 964
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_4
timestamp 1701704242
transform 1 0 211 0 1 418
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_0
timestamp 1701704242
transform 0 -1 933 1 0 2558
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_1
timestamp 1701704242
transform 1 0 1105 0 -1 754
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_2
timestamp 1701704242
transform 1 0 1105 0 -1 140
box 0 0 1 1
use M1M2_CDNS_52468879185371  M1M2_CDNS_52468879185371_0
timestamp 1701704242
transform 0 -1 391 1 0 2558
box 0 0 1 1
use M1M2_CDNS_52468879185371  M1M2_CDNS_52468879185371_1
timestamp 1701704242
transform 1 0 1105 0 -1 1234
box 0 0 1 1
use nfet_CDNS_52468879185374  nfet_CDNS_52468879185374_0
timestamp 1701704242
transform -1 0 1011 0 1 36
box -79 -26 879 110
use nfet_CDNS_52468879185374  nfet_CDNS_52468879185374_1
timestamp 1701704242
transform 1 0 211 0 1 290
box -79 -26 879 110
use nfet_CDNS_52468879185375  nfet_CDNS_52468879185375_0
timestamp 1701704242
transform -1 0 953 0 1 632
box -79 -26 176 326
use nfet_CDNS_52468879185375  nfet_CDNS_52468879185375_1
timestamp 1701704242
transform -1 0 953 0 -1 1360
box -79 -26 176 326
use nfet_CDNS_52468879185375  nfet_CDNS_52468879185375_2
timestamp 1701704242
transform 1 0 211 0 -1 1360
box -79 -26 176 326
use nfet_CDNS_52468879185375  nfet_CDNS_52468879185375_3
timestamp 1701704242
transform 1 0 211 0 1 632
box -79 -26 176 326
use nfet_CDNS_52468879185377  nfet_CDNS_52468879185377_0
timestamp 1701704242
transform -1 0 553 0 1 632
box -79 -26 276 326
use nfet_CDNS_52468879185377  nfet_CDNS_52468879185377_1
timestamp 1701704242
transform -1 0 553 0 -1 1360
box -79 -26 276 326
use nfet_CDNS_52468879185377  nfet_CDNS_52468879185377_2
timestamp 1701704242
transform 1 0 609 0 -1 1360
box -79 -26 276 326
use nfet_CDNS_52468879185377  nfet_CDNS_52468879185377_3
timestamp 1701704242
transform 1 0 609 0 1 632
box -79 -26 276 326
use pfet_CDNS_52468879185313  pfet_CDNS_52468879185313_0
timestamp 1701704242
transform 1 0 739 0 1 1530
box -119 -66 239 1066
use pfet_CDNS_52468879185378  pfet_CDNS_52468879185378_0
timestamp 1701704242
transform -1 0 683 0 1 1530
box -119 -66 591 1066
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_0
timestamp 1701704242
transform 0 1 1170 -1 0 2552
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_1
timestamp 1701704242
transform 0 1 1008 -1 0 1650
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_2
timestamp 1701704242
transform 0 1 1008 -1 0 2552
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_3
timestamp 1701704242
transform 0 1 1170 -1 0 250
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_4
timestamp 1701704242
transform -1 0 311 0 -1 1029
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_5
timestamp 1701704242
transform -1 0 987 0 -1 1029
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_0
timestamp 1701704242
transform 0 1 743 1 0 2562
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_0
timestamp 1701704242
transform 0 1 353 1 0 534
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_1
timestamp 1701704242
transform 0 1 609 1 0 1392
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_2
timestamp 1701704242
transform 0 1 609 1 0 534
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_3
timestamp 1701704242
transform 0 1 353 1 0 1392
box 0 0 1 1
use PYL1_CDNS_52468879185317  PYL1_CDNS_52468879185317_0
timestamp 1701704242
transform 0 -1 961 1 0 406
box 0 0 66 746
use PYL1_CDNS_52468879185327  PYL1_CDNS_52468879185327_0
timestamp 1701704242
transform 0 1 224 1 0 2562
box 0 0 1 1
use PYL1_CDNS_52468879185370  PYL1_CDNS_52468879185370_0
timestamp 1701704242
transform 0 -1 982 1 0 152
box 0 0 66 678
use PYres_CDNS_52468879185379  PYres_CDNS_52468879185379_0
timestamp 1701704242
transform 0 -1 1074 -1 0 2434
box -50 0 850 66
use PYres_CDNS_52468879185380  PYres_CDNS_52468879185380_0
timestamp 1701704242
transform 0 -1 1236 -1 0 2434
box -50 0 2250 66
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851255  sky130_fd_io__sio_tk_em1s_CDNS_524688791851255_0
timestamp 1701704242
transform 0 1 1184 1 0 812
box 0 0 1 1
<< labels >>
flabel comment s 1190 2501 1190 2501 0 FreeSans 300 0 0 0 int_res
flabel comment s 180 210 180 210 0 FreeSans 300 90 0 0 n<2>
flabel metal1 s 0 632 36 762 7 FreeSans 300 0 0 0 vgnd_io
port 2 nsew
flabel metal1 s 1242 632 1284 762 7 FreeSans 300 180 0 0 vgnd_io
port 2 nsew
flabel metal1 s 0 1800 36 1846 3 FreeSans 300 180 0 0 pu_h_n
port 3 nsew
flabel metal1 s 0 1570 36 1772 6 FreeSans 300 0 0 0 vcc_io
port 4 nsew
flabel metal1 s 0 1044 36 1246 7 FreeSans 300 0 0 0 vgnd_io
port 2 nsew
flabel metal1 s 1196 1800 1236 1846 7 FreeSans 300 0 0 0 pu_h_n
port 3 nsew
flabel metal1 s 1247 1570 1284 1772 6 FreeSans 300 180 0 0 vcc_io
port 4 nsew
flabel metal1 s 1242 1044 1284 1246 7 FreeSans 300 180 0 0 vgnd_io
port 2 nsew
flabel locali s 357 550 407 584 3 FreeSans 300 270 0 0 en_fast<3>
port 5 nsew
flabel locali s 613 550 663 584 3 FreeSans 300 270 0 0 en_fast<2>
port 6 nsew
flabel locali s 761 1408 811 1442 3 FreeSans 300 270 0 0 en_fast<1>
port 7 nsew
flabel locali s 357 1408 407 1442 3 FreeSans 300 270 0 0 en_fast<0>
port 8 nsew
flabel metal2 s 919 2558 985 2622 3 FreeSans 300 0 0 0 puen_h
port 9 nsew
flabel metal2 s 211 1402 263 1454 7 FreeSans 300 0 0 0 drvhi_h
port 10 nsew
<< properties >>
string GDS_END 87744916
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 87733112
<< end >>
