magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< nwell >>
rect 12135 10039 15401 10207
rect 15233 7872 15401 10039
rect 14811 7859 15401 7872
rect 14811 7706 15399 7859
rect 14811 7358 14985 7706
rect 14536 6991 14985 7358
rect 11603 6232 14985 6991
rect 11603 5530 14827 6232
<< pwell >>
rect 5528 11155 15803 11951
rect 5528 10547 5808 11155
rect -102 10267 5808 10547
rect 11586 8307 11689 9128
rect 11586 8206 14660 8307
rect 11586 7498 11710 8206
rect 15523 5081 15803 11155
rect 12399 2498 12564 2584
<< pdiff >>
rect 12769 2740 12816 3287
rect 16125 3208 16148 3557
rect 16105 3206 16148 3208
<< psubdiff >>
rect 5554 11896 15777 11925
rect 5554 11891 5656 11896
rect 5554 11857 5583 11891
rect 5617 11857 5656 11891
rect 11062 11862 11096 11896
rect 11130 11862 11164 11896
rect 11198 11862 11232 11896
rect 11266 11862 11300 11896
rect 11334 11862 11368 11896
rect 11402 11862 11436 11896
rect 11470 11862 11504 11896
rect 11538 11862 11572 11896
rect 11606 11862 11640 11896
rect 11674 11862 11708 11896
rect 11742 11862 11776 11896
rect 11810 11862 11845 11896
rect 11879 11862 11914 11896
rect 11948 11862 11983 11896
rect 12017 11862 12052 11896
rect 12086 11862 12121 11896
rect 12155 11862 12190 11896
rect 12224 11862 12259 11896
rect 12293 11862 12328 11896
rect 12362 11862 12397 11896
rect 12431 11862 12466 11896
rect 12500 11862 12535 11896
rect 12569 11862 12604 11896
rect 12638 11862 12673 11896
rect 12707 11862 12742 11896
rect 12776 11862 12811 11896
rect 12845 11862 12880 11896
rect 12914 11862 12949 11896
rect 12983 11862 13018 11896
rect 13052 11862 13087 11896
rect 13121 11862 13156 11896
rect 13190 11862 13225 11896
rect 13259 11862 13294 11896
rect 13328 11862 13363 11896
rect 13397 11862 13432 11896
rect 13466 11862 13501 11896
rect 13535 11862 13570 11896
rect 13604 11862 13639 11896
rect 13673 11862 13708 11896
rect 13742 11862 13777 11896
rect 13811 11862 13846 11896
rect 13880 11862 13915 11896
rect 13949 11862 13984 11896
rect 14018 11862 14053 11896
rect 14087 11862 14122 11896
rect 14156 11862 14191 11896
rect 14225 11862 14260 11896
rect 14294 11862 14329 11896
rect 14363 11862 14398 11896
rect 14432 11862 14467 11896
rect 14501 11862 14536 11896
rect 14570 11862 14605 11896
rect 14639 11862 14674 11896
rect 14708 11862 14743 11896
rect 14777 11862 14812 11896
rect 14846 11862 14881 11896
rect 14915 11862 14950 11896
rect 14984 11862 15019 11896
rect 15053 11862 15088 11896
rect 15122 11862 15157 11896
rect 15191 11862 15226 11896
rect 15260 11862 15295 11896
rect 15329 11862 15364 11896
rect 15398 11862 15433 11896
rect 15467 11862 15502 11896
rect 15536 11862 15571 11896
rect 15605 11862 15640 11896
rect 15674 11862 15709 11896
rect 15743 11862 15777 11896
rect 5554 11828 5656 11857
rect 11057 11828 15777 11862
rect 5554 11821 5651 11828
rect 5554 11787 5583 11821
rect 5617 11794 5651 11821
rect 11057 11794 11092 11828
rect 11126 11794 11161 11828
rect 11195 11794 11230 11828
rect 11264 11794 11299 11828
rect 11333 11794 11368 11828
rect 11402 11794 11437 11828
rect 11471 11794 11506 11828
rect 11540 11794 11575 11828
rect 11609 11794 11644 11828
rect 11678 11794 11713 11828
rect 11747 11794 11782 11828
rect 11816 11794 11851 11828
rect 11885 11794 11920 11828
rect 11954 11794 11989 11828
rect 12023 11794 12058 11828
rect 12092 11794 12127 11828
rect 12161 11794 12196 11828
rect 12230 11794 12265 11828
rect 12299 11794 12334 11828
rect 12368 11794 12403 11828
rect 12437 11794 12472 11828
rect 12506 11794 12541 11828
rect 12575 11794 12610 11828
rect 12644 11794 12679 11828
rect 12713 11794 12748 11828
rect 12782 11794 12817 11828
rect 12851 11794 12886 11828
rect 12920 11794 12955 11828
rect 12989 11794 13024 11828
rect 13058 11794 13093 11828
rect 13127 11794 13162 11828
rect 13196 11794 13231 11828
rect 13265 11794 13300 11828
rect 13334 11794 13369 11828
rect 13403 11794 13438 11828
rect 13472 11794 13507 11828
rect 13541 11794 13576 11828
rect 13610 11794 13645 11828
rect 13679 11794 13714 11828
rect 13748 11794 13783 11828
rect 13817 11794 13852 11828
rect 13886 11794 13921 11828
rect 13955 11794 13990 11828
rect 14024 11794 14059 11828
rect 14093 11794 14128 11828
rect 14162 11794 14197 11828
rect 14231 11794 14266 11828
rect 14300 11794 14335 11828
rect 14369 11794 14404 11828
rect 14438 11794 14473 11828
rect 14507 11794 14542 11828
rect 14576 11794 14611 11828
rect 14645 11794 14680 11828
rect 14714 11794 14749 11828
rect 14783 11794 14818 11828
rect 14852 11794 14887 11828
rect 14921 11794 14956 11828
rect 14990 11794 15025 11828
rect 15059 11794 15094 11828
rect 15128 11794 15163 11828
rect 15197 11794 15232 11828
rect 15266 11794 15301 11828
rect 15335 11794 15370 11828
rect 15404 11794 15439 11828
rect 15473 11794 15508 11828
rect 15542 11794 15577 11828
rect 15611 11794 15646 11828
rect 15680 11823 15777 11828
rect 5617 11787 5719 11794
rect 5554 11757 5719 11787
rect 5554 11751 5651 11757
rect 5554 11717 5583 11751
rect 5617 11723 5651 11751
rect 5685 11726 5719 11757
rect 10989 11760 15646 11794
rect 10989 11726 11024 11760
rect 11058 11726 11093 11760
rect 11127 11726 11162 11760
rect 11196 11726 11231 11760
rect 11265 11726 11300 11760
rect 11334 11726 11369 11760
rect 11403 11726 11438 11760
rect 11472 11726 11507 11760
rect 11541 11726 11576 11760
rect 11610 11726 11645 11760
rect 11679 11726 11714 11760
rect 11748 11726 11783 11760
rect 11817 11726 11852 11760
rect 11886 11726 11921 11760
rect 11955 11726 11990 11760
rect 12024 11726 12059 11760
rect 12093 11726 12128 11760
rect 12162 11726 12197 11760
rect 12231 11726 12266 11760
rect 12300 11726 12335 11760
rect 12369 11726 12404 11760
rect 12438 11726 12473 11760
rect 12507 11726 12542 11760
rect 12576 11726 12611 11760
rect 12645 11726 12680 11760
rect 12714 11726 12749 11760
rect 12783 11726 12818 11760
rect 12852 11726 12887 11760
rect 12921 11726 12956 11760
rect 12990 11726 13025 11760
rect 13059 11726 13094 11760
rect 13128 11726 13163 11760
rect 13197 11726 13232 11760
rect 13266 11726 13301 11760
rect 13335 11726 13370 11760
rect 13404 11726 13439 11760
rect 13473 11726 13508 11760
rect 13542 11726 13577 11760
rect 13611 11726 13646 11760
rect 13680 11726 13715 11760
rect 13749 11726 13784 11760
rect 13818 11726 13853 11760
rect 13887 11726 13922 11760
rect 13956 11726 13991 11760
rect 14025 11726 14060 11760
rect 14094 11726 14129 11760
rect 14163 11726 14198 11760
rect 14232 11726 14267 11760
rect 14301 11726 14336 11760
rect 14370 11726 14405 11760
rect 14439 11726 14474 11760
rect 14508 11726 14543 11760
rect 14577 11726 14612 11760
rect 14646 11726 14681 11760
rect 14715 11726 14750 11760
rect 14784 11726 14819 11760
rect 14853 11726 14888 11760
rect 14922 11726 14957 11760
rect 14991 11726 15026 11760
rect 15060 11726 15095 11760
rect 15129 11726 15164 11760
rect 15198 11726 15233 11760
rect 15267 11726 15302 11760
rect 15336 11726 15371 11760
rect 15405 11726 15440 11760
rect 15474 11726 15509 11760
rect 15543 11726 15578 11760
rect 5685 11723 15578 11726
rect 5617 11717 15578 11723
rect 5554 11690 15578 11717
rect 5554 11686 5719 11690
rect 5554 11681 5651 11686
rect 5554 11647 5583 11681
rect 5617 11652 5651 11681
rect 5685 11656 5719 11686
rect 5753 11656 15578 11690
rect 5685 11652 15578 11656
rect 5617 11651 15578 11652
rect 5617 11647 5806 11651
rect 5554 11620 5806 11647
rect 5554 11615 5719 11620
rect 5554 11611 5651 11615
rect 5554 11577 5583 11611
rect 5617 11581 5651 11611
rect 5685 11586 5719 11615
rect 5753 11617 5806 11620
rect 5840 11617 5875 11651
rect 5909 11617 5944 11651
rect 5978 11617 6013 11651
rect 6047 11617 6082 11651
rect 6116 11617 6151 11651
rect 6185 11617 6220 11651
rect 6254 11617 6289 11651
rect 6323 11617 6358 11651
rect 6392 11617 6427 11651
rect 6461 11617 6496 11651
rect 6530 11617 6565 11651
rect 6599 11617 6634 11651
rect 6668 11617 6703 11651
rect 6737 11617 6772 11651
rect 6806 11617 6841 11651
rect 6875 11617 6910 11651
rect 6944 11617 6979 11651
rect 7013 11617 7048 11651
rect 7082 11617 7117 11651
rect 7151 11617 7186 11651
rect 7220 11617 7255 11651
rect 7289 11617 7324 11651
rect 7358 11617 7393 11651
rect 7427 11617 7462 11651
rect 7496 11617 7531 11651
rect 7565 11617 7600 11651
rect 7634 11617 7669 11651
rect 7703 11617 7738 11651
rect 7772 11617 7807 11651
rect 7841 11617 7875 11651
rect 7909 11617 7943 11651
rect 7977 11617 8011 11651
rect 8045 11617 8079 11651
rect 8113 11617 8147 11651
rect 8181 11617 8215 11651
rect 8249 11617 8283 11651
rect 8317 11617 8351 11651
rect 8385 11617 8419 11651
rect 8453 11617 8487 11651
rect 8521 11617 8555 11651
rect 8589 11617 8623 11651
rect 8657 11617 8691 11651
rect 8725 11617 8759 11651
rect 8793 11617 8827 11651
rect 8861 11617 8895 11651
rect 8929 11617 8963 11651
rect 8997 11617 9031 11651
rect 9065 11617 9099 11651
rect 9133 11617 9167 11651
rect 9201 11617 9235 11651
rect 9269 11617 9303 11651
rect 9337 11617 9371 11651
rect 9405 11617 9439 11651
rect 9473 11617 9507 11651
rect 9541 11617 9575 11651
rect 9609 11617 9643 11651
rect 9677 11617 9711 11651
rect 9745 11617 9779 11651
rect 9813 11617 9847 11651
rect 9881 11617 9915 11651
rect 9949 11617 9983 11651
rect 10017 11617 10051 11651
rect 10085 11617 10119 11651
rect 10153 11617 10187 11651
rect 10221 11617 10255 11651
rect 10289 11617 10323 11651
rect 10357 11617 10391 11651
rect 10425 11617 10459 11651
rect 10493 11617 10527 11651
rect 10561 11617 10595 11651
rect 10629 11617 10663 11651
rect 10697 11617 10731 11651
rect 10765 11617 10799 11651
rect 10833 11617 10867 11651
rect 10901 11617 10935 11651
rect 10969 11617 11003 11651
rect 11037 11617 11071 11651
rect 11105 11617 11139 11651
rect 11173 11617 11207 11651
rect 11241 11617 11275 11651
rect 11309 11617 11343 11651
rect 11377 11617 11411 11651
rect 11445 11617 11479 11651
rect 11513 11617 11547 11651
rect 11581 11617 11615 11651
rect 11649 11617 11683 11651
rect 11717 11617 11751 11651
rect 11785 11617 11819 11651
rect 11853 11617 11887 11651
rect 11921 11617 11955 11651
rect 11989 11617 12023 11651
rect 12057 11617 12091 11651
rect 12125 11617 12159 11651
rect 12193 11617 12227 11651
rect 12261 11617 12295 11651
rect 12329 11617 12363 11651
rect 12397 11617 12431 11651
rect 12465 11617 12499 11651
rect 12533 11617 12567 11651
rect 12601 11617 12635 11651
rect 12669 11617 12703 11651
rect 12737 11617 12771 11651
rect 12805 11617 12839 11651
rect 12873 11617 12907 11651
rect 12941 11617 12975 11651
rect 13009 11617 13043 11651
rect 13077 11617 13111 11651
rect 13145 11617 13179 11651
rect 13213 11617 13247 11651
rect 13281 11617 13315 11651
rect 13349 11617 13383 11651
rect 13417 11617 13451 11651
rect 13485 11617 13519 11651
rect 13553 11617 13587 11651
rect 13621 11617 13655 11651
rect 13689 11617 13723 11651
rect 13757 11617 13791 11651
rect 13825 11617 13859 11651
rect 13893 11617 13927 11651
rect 13961 11617 13995 11651
rect 14029 11617 14063 11651
rect 14097 11617 14131 11651
rect 14165 11617 14199 11651
rect 14233 11617 14267 11651
rect 14301 11617 14335 11651
rect 14369 11617 14403 11651
rect 14437 11617 14471 11651
rect 14505 11617 14539 11651
rect 14573 11617 14607 11651
rect 14641 11617 14675 11651
rect 14709 11617 14743 11651
rect 14777 11617 14811 11651
rect 14845 11617 14879 11651
rect 14913 11617 14947 11651
rect 14981 11617 15015 11651
rect 15049 11617 15083 11651
rect 15117 11617 15151 11651
rect 15185 11617 15219 11651
rect 15253 11617 15287 11651
rect 15321 11617 15355 11651
rect 15389 11617 15423 11651
rect 15457 11617 15491 11651
rect 15525 11617 15578 11651
rect 5753 11586 15578 11617
rect 5685 11581 15578 11586
rect 5617 11579 15578 11581
rect 5617 11577 5806 11579
rect 5554 11550 5806 11577
rect 5554 11544 5719 11550
rect 5554 11541 5651 11544
rect 5554 11507 5583 11541
rect 5617 11510 5651 11541
rect 5685 11516 5719 11544
rect 5753 11545 5806 11550
rect 5840 11545 5875 11579
rect 5909 11545 5944 11579
rect 5978 11545 6013 11579
rect 6047 11545 6082 11579
rect 6116 11545 6151 11579
rect 6185 11545 6220 11579
rect 6254 11545 6289 11579
rect 6323 11545 6358 11579
rect 6392 11545 6427 11579
rect 6461 11545 6496 11579
rect 6530 11545 6565 11579
rect 6599 11545 6634 11579
rect 6668 11545 6703 11579
rect 6737 11545 6772 11579
rect 6806 11545 6841 11579
rect 6875 11545 6910 11579
rect 6944 11545 6979 11579
rect 7013 11545 7048 11579
rect 7082 11545 7117 11579
rect 7151 11545 7186 11579
rect 7220 11545 7255 11579
rect 7289 11545 7324 11579
rect 7358 11545 7393 11579
rect 7427 11545 7462 11579
rect 7496 11545 7531 11579
rect 7565 11545 7600 11579
rect 7634 11545 7669 11579
rect 7703 11545 7738 11579
rect 7772 11545 7807 11579
rect 7841 11545 7875 11579
rect 7909 11545 7943 11579
rect 7977 11545 8011 11579
rect 8045 11545 8079 11579
rect 8113 11545 8147 11579
rect 8181 11545 8215 11579
rect 8249 11545 8283 11579
rect 8317 11545 8351 11579
rect 8385 11545 8419 11579
rect 8453 11545 8487 11579
rect 8521 11545 8555 11579
rect 8589 11545 8623 11579
rect 8657 11545 8691 11579
rect 8725 11545 8759 11579
rect 8793 11545 8827 11579
rect 8861 11545 8895 11579
rect 8929 11545 8963 11579
rect 8997 11545 9031 11579
rect 9065 11545 9099 11579
rect 9133 11545 9167 11579
rect 9201 11545 9235 11579
rect 9269 11545 9303 11579
rect 9337 11545 9371 11579
rect 9405 11545 9439 11579
rect 9473 11545 9507 11579
rect 9541 11545 9575 11579
rect 9609 11545 9643 11579
rect 9677 11545 9711 11579
rect 9745 11545 9779 11579
rect 9813 11545 9847 11579
rect 9881 11545 9915 11579
rect 9949 11545 9983 11579
rect 10017 11545 10051 11579
rect 10085 11545 10119 11579
rect 10153 11545 10187 11579
rect 10221 11545 10255 11579
rect 10289 11545 10323 11579
rect 10357 11545 10391 11579
rect 10425 11545 10459 11579
rect 10493 11545 10527 11579
rect 10561 11545 10595 11579
rect 10629 11545 10663 11579
rect 10697 11545 10731 11579
rect 10765 11545 10799 11579
rect 10833 11545 10867 11579
rect 10901 11545 10935 11579
rect 10969 11545 11003 11579
rect 11037 11545 11071 11579
rect 11105 11545 11139 11579
rect 11173 11545 11207 11579
rect 11241 11545 11275 11579
rect 11309 11545 11343 11579
rect 11377 11545 11411 11579
rect 11445 11545 11479 11579
rect 11513 11545 11547 11579
rect 11581 11545 11615 11579
rect 11649 11545 11683 11579
rect 11717 11545 11751 11579
rect 11785 11545 11819 11579
rect 11853 11545 11887 11579
rect 11921 11545 11955 11579
rect 11989 11545 12023 11579
rect 12057 11545 12091 11579
rect 12125 11545 12159 11579
rect 12193 11545 12227 11579
rect 12261 11545 12295 11579
rect 12329 11545 12363 11579
rect 12397 11545 12431 11579
rect 12465 11545 12499 11579
rect 12533 11545 12567 11579
rect 12601 11545 12635 11579
rect 12669 11545 12703 11579
rect 12737 11545 12771 11579
rect 12805 11545 12839 11579
rect 12873 11545 12907 11579
rect 12941 11545 12975 11579
rect 13009 11545 13043 11579
rect 13077 11545 13111 11579
rect 13145 11545 13179 11579
rect 13213 11545 13247 11579
rect 13281 11545 13315 11579
rect 13349 11545 13383 11579
rect 13417 11545 13451 11579
rect 13485 11545 13519 11579
rect 13553 11545 13587 11579
rect 13621 11545 13655 11579
rect 13689 11545 13723 11579
rect 13757 11545 13791 11579
rect 13825 11545 13859 11579
rect 13893 11545 13927 11579
rect 13961 11545 13995 11579
rect 14029 11545 14063 11579
rect 14097 11545 14131 11579
rect 14165 11545 14199 11579
rect 14233 11545 14267 11579
rect 14301 11545 14335 11579
rect 14369 11545 14403 11579
rect 14437 11545 14471 11579
rect 14505 11545 14539 11579
rect 14573 11545 14607 11579
rect 14641 11545 14675 11579
rect 14709 11545 14743 11579
rect 14777 11545 14811 11579
rect 14845 11545 14879 11579
rect 14913 11545 14947 11579
rect 14981 11545 15015 11579
rect 15049 11545 15083 11579
rect 15117 11545 15151 11579
rect 15185 11545 15219 11579
rect 15253 11545 15287 11579
rect 15321 11545 15355 11579
rect 15389 11545 15423 11579
rect 15457 11545 15491 11579
rect 15525 11545 15578 11579
rect 5753 11516 15578 11545
rect 5685 11510 15578 11516
rect 5617 11507 15578 11510
rect 5554 11480 5806 11507
rect 5554 11474 5719 11480
rect 5554 11471 5651 11474
rect 5554 11437 5583 11471
rect 5617 11440 5651 11471
rect 5685 11446 5719 11474
rect 5753 11473 5806 11480
rect 5840 11473 5875 11507
rect 5909 11473 5944 11507
rect 5978 11473 6013 11507
rect 6047 11473 6082 11507
rect 6116 11473 6151 11507
rect 6185 11473 6220 11507
rect 6254 11473 6289 11507
rect 6323 11473 6358 11507
rect 6392 11473 6427 11507
rect 6461 11473 6496 11507
rect 6530 11473 6565 11507
rect 6599 11473 6634 11507
rect 6668 11473 6703 11507
rect 6737 11473 6772 11507
rect 6806 11473 6841 11507
rect 6875 11473 6910 11507
rect 6944 11473 6979 11507
rect 7013 11473 7048 11507
rect 7082 11473 7117 11507
rect 7151 11473 7186 11507
rect 7220 11473 7255 11507
rect 7289 11473 7324 11507
rect 7358 11473 7393 11507
rect 7427 11473 7462 11507
rect 7496 11473 7531 11507
rect 7565 11473 7600 11507
rect 7634 11473 7669 11507
rect 7703 11473 7738 11507
rect 7772 11473 7807 11507
rect 7841 11473 7875 11507
rect 7909 11473 7943 11507
rect 7977 11473 8011 11507
rect 8045 11473 8079 11507
rect 8113 11473 8147 11507
rect 8181 11473 8215 11507
rect 8249 11473 8283 11507
rect 8317 11473 8351 11507
rect 8385 11473 8419 11507
rect 8453 11473 8487 11507
rect 8521 11473 8555 11507
rect 8589 11473 8623 11507
rect 8657 11473 8691 11507
rect 8725 11473 8759 11507
rect 8793 11473 8827 11507
rect 8861 11473 8895 11507
rect 8929 11473 8963 11507
rect 8997 11473 9031 11507
rect 9065 11473 9099 11507
rect 9133 11473 9167 11507
rect 9201 11473 9235 11507
rect 9269 11473 9303 11507
rect 9337 11473 9371 11507
rect 9405 11473 9439 11507
rect 9473 11473 9507 11507
rect 9541 11473 9575 11507
rect 9609 11473 9643 11507
rect 9677 11473 9711 11507
rect 9745 11473 9779 11507
rect 9813 11473 9847 11507
rect 9881 11473 9915 11507
rect 9949 11473 9983 11507
rect 10017 11473 10051 11507
rect 10085 11473 10119 11507
rect 10153 11473 10187 11507
rect 10221 11473 10255 11507
rect 10289 11473 10323 11507
rect 10357 11473 10391 11507
rect 10425 11473 10459 11507
rect 10493 11473 10527 11507
rect 10561 11473 10595 11507
rect 10629 11473 10663 11507
rect 10697 11473 10731 11507
rect 10765 11473 10799 11507
rect 10833 11473 10867 11507
rect 10901 11473 10935 11507
rect 10969 11473 11003 11507
rect 11037 11473 11071 11507
rect 11105 11473 11139 11507
rect 11173 11473 11207 11507
rect 11241 11473 11275 11507
rect 11309 11473 11343 11507
rect 11377 11473 11411 11507
rect 11445 11473 11479 11507
rect 11513 11473 11547 11507
rect 11581 11473 11615 11507
rect 11649 11473 11683 11507
rect 11717 11473 11751 11507
rect 11785 11473 11819 11507
rect 11853 11473 11887 11507
rect 11921 11473 11955 11507
rect 11989 11473 12023 11507
rect 12057 11473 12091 11507
rect 12125 11473 12159 11507
rect 12193 11473 12227 11507
rect 12261 11473 12295 11507
rect 12329 11473 12363 11507
rect 12397 11473 12431 11507
rect 12465 11473 12499 11507
rect 12533 11473 12567 11507
rect 12601 11473 12635 11507
rect 12669 11473 12703 11507
rect 12737 11473 12771 11507
rect 12805 11473 12839 11507
rect 12873 11473 12907 11507
rect 12941 11473 12975 11507
rect 13009 11473 13043 11507
rect 13077 11473 13111 11507
rect 13145 11473 13179 11507
rect 13213 11473 13247 11507
rect 13281 11473 13315 11507
rect 13349 11473 13383 11507
rect 13417 11473 13451 11507
rect 13485 11473 13519 11507
rect 13553 11473 13587 11507
rect 13621 11473 13655 11507
rect 13689 11473 13723 11507
rect 13757 11473 13791 11507
rect 13825 11473 13859 11507
rect 13893 11473 13927 11507
rect 13961 11473 13995 11507
rect 14029 11473 14063 11507
rect 14097 11473 14131 11507
rect 14165 11473 14199 11507
rect 14233 11473 14267 11507
rect 14301 11473 14335 11507
rect 14369 11473 14403 11507
rect 14437 11473 14471 11507
rect 14505 11473 14539 11507
rect 14573 11473 14607 11507
rect 14641 11473 14675 11507
rect 14709 11473 14743 11507
rect 14777 11473 14811 11507
rect 14845 11473 14879 11507
rect 14913 11473 14947 11507
rect 14981 11473 15015 11507
rect 15049 11473 15083 11507
rect 15117 11473 15151 11507
rect 15185 11473 15219 11507
rect 15253 11473 15287 11507
rect 15321 11473 15355 11507
rect 15389 11473 15423 11507
rect 15457 11473 15491 11507
rect 15525 11473 15578 11507
rect 5753 11446 15578 11473
rect 5685 11440 15578 11446
rect 5617 11437 15578 11440
rect 5554 11435 15578 11437
rect 5554 11410 5806 11435
rect 5554 11404 5719 11410
rect 5554 11401 5651 11404
rect 5554 11367 5583 11401
rect 5617 11370 5651 11401
rect 5685 11376 5719 11404
rect 5753 11401 5806 11410
rect 5840 11401 5875 11435
rect 5909 11401 5944 11435
rect 5978 11401 6013 11435
rect 6047 11401 6082 11435
rect 6116 11401 6151 11435
rect 6185 11401 6220 11435
rect 6254 11401 6289 11435
rect 6323 11401 6358 11435
rect 6392 11401 6427 11435
rect 6461 11401 6496 11435
rect 6530 11401 6565 11435
rect 6599 11401 6634 11435
rect 6668 11401 6703 11435
rect 6737 11401 6772 11435
rect 6806 11401 6841 11435
rect 6875 11401 6910 11435
rect 6944 11401 6979 11435
rect 7013 11401 7048 11435
rect 7082 11401 7117 11435
rect 7151 11401 7186 11435
rect 7220 11401 7255 11435
rect 7289 11401 7324 11435
rect 7358 11401 7393 11435
rect 7427 11401 7462 11435
rect 7496 11401 7531 11435
rect 7565 11401 7600 11435
rect 7634 11401 7669 11435
rect 7703 11401 7738 11435
rect 7772 11401 7807 11435
rect 7841 11401 7875 11435
rect 7909 11401 7943 11435
rect 7977 11401 8011 11435
rect 8045 11401 8079 11435
rect 8113 11401 8147 11435
rect 8181 11401 8215 11435
rect 8249 11401 8283 11435
rect 8317 11401 8351 11435
rect 8385 11401 8419 11435
rect 8453 11401 8487 11435
rect 8521 11401 8555 11435
rect 8589 11401 8623 11435
rect 8657 11401 8691 11435
rect 8725 11401 8759 11435
rect 8793 11401 8827 11435
rect 8861 11401 8895 11435
rect 8929 11401 8963 11435
rect 8997 11401 9031 11435
rect 9065 11401 9099 11435
rect 9133 11401 9167 11435
rect 9201 11401 9235 11435
rect 9269 11401 9303 11435
rect 9337 11401 9371 11435
rect 9405 11401 9439 11435
rect 9473 11401 9507 11435
rect 9541 11401 9575 11435
rect 9609 11401 9643 11435
rect 9677 11401 9711 11435
rect 9745 11401 9779 11435
rect 9813 11401 9847 11435
rect 9881 11401 9915 11435
rect 9949 11401 9983 11435
rect 10017 11401 10051 11435
rect 10085 11401 10119 11435
rect 10153 11401 10187 11435
rect 10221 11401 10255 11435
rect 10289 11401 10323 11435
rect 10357 11401 10391 11435
rect 10425 11401 10459 11435
rect 10493 11401 10527 11435
rect 10561 11401 10595 11435
rect 10629 11401 10663 11435
rect 10697 11401 10731 11435
rect 10765 11401 10799 11435
rect 10833 11401 10867 11435
rect 10901 11401 10935 11435
rect 10969 11401 11003 11435
rect 11037 11401 11071 11435
rect 11105 11401 11139 11435
rect 11173 11401 11207 11435
rect 11241 11401 11275 11435
rect 11309 11401 11343 11435
rect 11377 11401 11411 11435
rect 11445 11401 11479 11435
rect 11513 11401 11547 11435
rect 11581 11401 11615 11435
rect 11649 11401 11683 11435
rect 11717 11401 11751 11435
rect 11785 11401 11819 11435
rect 11853 11401 11887 11435
rect 11921 11401 11955 11435
rect 11989 11401 12023 11435
rect 12057 11401 12091 11435
rect 12125 11401 12159 11435
rect 12193 11401 12227 11435
rect 12261 11401 12295 11435
rect 12329 11401 12363 11435
rect 12397 11401 12431 11435
rect 12465 11401 12499 11435
rect 12533 11401 12567 11435
rect 12601 11401 12635 11435
rect 12669 11401 12703 11435
rect 12737 11401 12771 11435
rect 12805 11401 12839 11435
rect 12873 11401 12907 11435
rect 12941 11401 12975 11435
rect 13009 11401 13043 11435
rect 13077 11401 13111 11435
rect 13145 11401 13179 11435
rect 13213 11401 13247 11435
rect 13281 11401 13315 11435
rect 13349 11401 13383 11435
rect 13417 11401 13451 11435
rect 13485 11401 13519 11435
rect 13553 11401 13587 11435
rect 13621 11401 13655 11435
rect 13689 11401 13723 11435
rect 13757 11401 13791 11435
rect 13825 11401 13859 11435
rect 13893 11401 13927 11435
rect 13961 11401 13995 11435
rect 14029 11401 14063 11435
rect 14097 11401 14131 11435
rect 14165 11401 14199 11435
rect 14233 11401 14267 11435
rect 14301 11401 14335 11435
rect 14369 11401 14403 11435
rect 14437 11401 14471 11435
rect 14505 11401 14539 11435
rect 14573 11401 14607 11435
rect 14641 11401 14675 11435
rect 14709 11401 14743 11435
rect 14777 11401 14811 11435
rect 14845 11401 14879 11435
rect 14913 11401 14947 11435
rect 14981 11401 15015 11435
rect 15049 11401 15083 11435
rect 15117 11401 15151 11435
rect 15185 11401 15219 11435
rect 15253 11401 15287 11435
rect 15321 11401 15355 11435
rect 15389 11401 15423 11435
rect 15457 11401 15491 11435
rect 15525 11401 15578 11435
rect 5753 11376 15578 11401
rect 5685 11370 15578 11376
rect 5617 11367 15578 11370
rect 5554 11363 15578 11367
rect 5554 11340 5806 11363
rect 5554 11334 5719 11340
rect 5554 11331 5651 11334
rect 5554 11297 5583 11331
rect 5617 11300 5651 11331
rect 5685 11306 5719 11334
rect 5753 11329 5806 11340
rect 5840 11329 5875 11363
rect 5909 11329 5944 11363
rect 5978 11329 6013 11363
rect 6047 11329 6082 11363
rect 6116 11329 6151 11363
rect 6185 11329 6220 11363
rect 6254 11329 6289 11363
rect 6323 11329 6358 11363
rect 6392 11329 6427 11363
rect 6461 11329 6496 11363
rect 6530 11329 6565 11363
rect 6599 11329 6634 11363
rect 6668 11329 6703 11363
rect 6737 11329 6772 11363
rect 6806 11329 6841 11363
rect 6875 11329 6910 11363
rect 6944 11329 6979 11363
rect 7013 11329 7048 11363
rect 7082 11329 7117 11363
rect 7151 11329 7186 11363
rect 7220 11329 7255 11363
rect 7289 11329 7324 11363
rect 7358 11329 7393 11363
rect 7427 11329 7462 11363
rect 7496 11329 7531 11363
rect 7565 11329 7600 11363
rect 7634 11329 7669 11363
rect 7703 11329 7738 11363
rect 7772 11329 7807 11363
rect 7841 11329 7875 11363
rect 7909 11329 7943 11363
rect 7977 11329 8011 11363
rect 8045 11329 8079 11363
rect 8113 11329 8147 11363
rect 8181 11329 8215 11363
rect 8249 11329 8283 11363
rect 8317 11329 8351 11363
rect 8385 11329 8419 11363
rect 8453 11329 8487 11363
rect 8521 11329 8555 11363
rect 8589 11329 8623 11363
rect 8657 11329 8691 11363
rect 8725 11329 8759 11363
rect 8793 11329 8827 11363
rect 8861 11329 8895 11363
rect 8929 11329 8963 11363
rect 8997 11329 9031 11363
rect 9065 11329 9099 11363
rect 9133 11329 9167 11363
rect 9201 11329 9235 11363
rect 9269 11329 9303 11363
rect 9337 11329 9371 11363
rect 9405 11329 9439 11363
rect 9473 11329 9507 11363
rect 9541 11329 9575 11363
rect 9609 11329 9643 11363
rect 9677 11329 9711 11363
rect 9745 11329 9779 11363
rect 9813 11329 9847 11363
rect 9881 11329 9915 11363
rect 9949 11329 9983 11363
rect 10017 11329 10051 11363
rect 10085 11329 10119 11363
rect 10153 11329 10187 11363
rect 10221 11329 10255 11363
rect 10289 11329 10323 11363
rect 10357 11329 10391 11363
rect 10425 11329 10459 11363
rect 10493 11329 10527 11363
rect 10561 11329 10595 11363
rect 10629 11329 10663 11363
rect 10697 11329 10731 11363
rect 10765 11329 10799 11363
rect 10833 11329 10867 11363
rect 10901 11329 10935 11363
rect 10969 11329 11003 11363
rect 11037 11329 11071 11363
rect 11105 11329 11139 11363
rect 11173 11329 11207 11363
rect 11241 11329 11275 11363
rect 11309 11329 11343 11363
rect 11377 11329 11411 11363
rect 11445 11329 11479 11363
rect 11513 11329 11547 11363
rect 11581 11329 11615 11363
rect 11649 11329 11683 11363
rect 11717 11329 11751 11363
rect 11785 11329 11819 11363
rect 11853 11329 11887 11363
rect 11921 11329 11955 11363
rect 11989 11329 12023 11363
rect 12057 11329 12091 11363
rect 12125 11329 12159 11363
rect 12193 11329 12227 11363
rect 12261 11329 12295 11363
rect 12329 11329 12363 11363
rect 12397 11329 12431 11363
rect 12465 11329 12499 11363
rect 12533 11329 12567 11363
rect 12601 11329 12635 11363
rect 12669 11329 12703 11363
rect 12737 11329 12771 11363
rect 12805 11329 12839 11363
rect 12873 11329 12907 11363
rect 12941 11329 12975 11363
rect 13009 11329 13043 11363
rect 13077 11329 13111 11363
rect 13145 11329 13179 11363
rect 13213 11329 13247 11363
rect 13281 11329 13315 11363
rect 13349 11329 13383 11363
rect 13417 11329 13451 11363
rect 13485 11329 13519 11363
rect 13553 11329 13587 11363
rect 13621 11329 13655 11363
rect 13689 11329 13723 11363
rect 13757 11329 13791 11363
rect 13825 11329 13859 11363
rect 13893 11329 13927 11363
rect 13961 11329 13995 11363
rect 14029 11329 14063 11363
rect 14097 11329 14131 11363
rect 14165 11329 14199 11363
rect 14233 11329 14267 11363
rect 14301 11329 14335 11363
rect 14369 11329 14403 11363
rect 14437 11329 14471 11363
rect 14505 11329 14539 11363
rect 14573 11329 14607 11363
rect 14641 11329 14675 11363
rect 14709 11329 14743 11363
rect 14777 11329 14811 11363
rect 14845 11329 14879 11363
rect 14913 11329 14947 11363
rect 14981 11329 15015 11363
rect 15049 11329 15083 11363
rect 15117 11329 15151 11363
rect 15185 11329 15219 11363
rect 15253 11329 15287 11363
rect 15321 11329 15355 11363
rect 15389 11329 15423 11363
rect 15457 11329 15491 11363
rect 15525 11329 15578 11363
rect 5753 11306 15578 11329
rect 5685 11300 15578 11306
rect 5617 11297 15578 11300
rect 5554 11291 15578 11297
rect 5554 11270 5806 11291
rect 5554 11264 5719 11270
rect 5554 11261 5651 11264
rect 5554 11227 5583 11261
rect 5617 11230 5651 11261
rect 5685 11236 5719 11264
rect 5753 11257 5806 11270
rect 5840 11257 5875 11291
rect 5909 11257 5944 11291
rect 5978 11257 6013 11291
rect 6047 11257 6082 11291
rect 6116 11257 6151 11291
rect 6185 11257 6220 11291
rect 6254 11257 6289 11291
rect 6323 11257 6358 11291
rect 6392 11257 6427 11291
rect 6461 11257 6496 11291
rect 6530 11257 6565 11291
rect 6599 11257 6634 11291
rect 6668 11257 6703 11291
rect 6737 11257 6772 11291
rect 6806 11257 6841 11291
rect 6875 11257 6910 11291
rect 6944 11257 6979 11291
rect 7013 11257 7048 11291
rect 7082 11257 7117 11291
rect 7151 11257 7186 11291
rect 7220 11257 7255 11291
rect 7289 11257 7324 11291
rect 7358 11257 7393 11291
rect 7427 11257 7462 11291
rect 7496 11257 7531 11291
rect 7565 11257 7600 11291
rect 7634 11257 7669 11291
rect 7703 11257 7738 11291
rect 7772 11257 7807 11291
rect 7841 11257 7875 11291
rect 7909 11257 7943 11291
rect 7977 11257 8011 11291
rect 8045 11257 8079 11291
rect 8113 11257 8147 11291
rect 8181 11257 8215 11291
rect 8249 11257 8283 11291
rect 8317 11257 8351 11291
rect 8385 11257 8419 11291
rect 8453 11257 8487 11291
rect 8521 11257 8555 11291
rect 8589 11257 8623 11291
rect 8657 11257 8691 11291
rect 8725 11257 8759 11291
rect 8793 11257 8827 11291
rect 8861 11257 8895 11291
rect 8929 11257 8963 11291
rect 8997 11257 9031 11291
rect 9065 11257 9099 11291
rect 9133 11257 9167 11291
rect 9201 11257 9235 11291
rect 9269 11257 9303 11291
rect 9337 11257 9371 11291
rect 9405 11257 9439 11291
rect 9473 11257 9507 11291
rect 9541 11257 9575 11291
rect 9609 11257 9643 11291
rect 9677 11257 9711 11291
rect 9745 11257 9779 11291
rect 9813 11257 9847 11291
rect 9881 11257 9915 11291
rect 9949 11257 9983 11291
rect 10017 11257 10051 11291
rect 10085 11257 10119 11291
rect 10153 11257 10187 11291
rect 10221 11257 10255 11291
rect 10289 11257 10323 11291
rect 10357 11257 10391 11291
rect 10425 11257 10459 11291
rect 10493 11257 10527 11291
rect 10561 11257 10595 11291
rect 10629 11257 10663 11291
rect 10697 11257 10731 11291
rect 10765 11257 10799 11291
rect 10833 11257 10867 11291
rect 10901 11257 10935 11291
rect 10969 11257 11003 11291
rect 11037 11257 11071 11291
rect 11105 11257 11139 11291
rect 11173 11257 11207 11291
rect 11241 11257 11275 11291
rect 11309 11257 11343 11291
rect 11377 11257 11411 11291
rect 11445 11257 11479 11291
rect 11513 11257 11547 11291
rect 11581 11257 11615 11291
rect 11649 11257 11683 11291
rect 11717 11257 11751 11291
rect 11785 11257 11819 11291
rect 11853 11257 11887 11291
rect 11921 11257 11955 11291
rect 11989 11257 12023 11291
rect 12057 11257 12091 11291
rect 12125 11257 12159 11291
rect 12193 11257 12227 11291
rect 12261 11257 12295 11291
rect 12329 11257 12363 11291
rect 12397 11257 12431 11291
rect 12465 11257 12499 11291
rect 12533 11257 12567 11291
rect 12601 11257 12635 11291
rect 12669 11257 12703 11291
rect 12737 11257 12771 11291
rect 12805 11257 12839 11291
rect 12873 11257 12907 11291
rect 12941 11257 12975 11291
rect 13009 11257 13043 11291
rect 13077 11257 13111 11291
rect 13145 11257 13179 11291
rect 13213 11257 13247 11291
rect 13281 11257 13315 11291
rect 13349 11257 13383 11291
rect 13417 11257 13451 11291
rect 13485 11257 13519 11291
rect 13553 11257 13587 11291
rect 13621 11257 13655 11291
rect 13689 11257 13723 11291
rect 13757 11257 13791 11291
rect 13825 11257 13859 11291
rect 13893 11257 13927 11291
rect 13961 11257 13995 11291
rect 14029 11257 14063 11291
rect 14097 11257 14131 11291
rect 14165 11257 14199 11291
rect 14233 11257 14267 11291
rect 14301 11257 14335 11291
rect 14369 11257 14403 11291
rect 14437 11257 14471 11291
rect 14505 11257 14539 11291
rect 14573 11257 14607 11291
rect 14641 11257 14675 11291
rect 14709 11257 14743 11291
rect 14777 11257 14811 11291
rect 14845 11257 14879 11291
rect 14913 11257 14947 11291
rect 14981 11257 15015 11291
rect 15049 11257 15083 11291
rect 15117 11257 15151 11291
rect 15185 11257 15219 11291
rect 15253 11257 15287 11291
rect 15321 11257 15355 11291
rect 15389 11257 15423 11291
rect 15457 11257 15491 11291
rect 15525 11257 15578 11291
rect 5753 11236 15578 11257
rect 5685 11230 15578 11236
rect 5617 11227 15578 11230
rect 5554 11219 15578 11227
rect 5554 11200 5806 11219
rect 5554 11194 5719 11200
rect 5554 11191 5651 11194
rect 5554 11157 5583 11191
rect 5617 11160 5651 11191
rect 5685 11166 5719 11194
rect 5753 11185 5806 11200
rect 5840 11185 5875 11219
rect 5909 11185 5944 11219
rect 5978 11185 6013 11219
rect 6047 11185 6082 11219
rect 6116 11185 6151 11219
rect 6185 11185 6220 11219
rect 6254 11185 6289 11219
rect 6323 11185 6358 11219
rect 6392 11185 6427 11219
rect 6461 11185 6496 11219
rect 6530 11185 6565 11219
rect 6599 11185 6634 11219
rect 6668 11185 6703 11219
rect 6737 11185 6772 11219
rect 6806 11185 6841 11219
rect 6875 11185 6910 11219
rect 6944 11185 6979 11219
rect 7013 11185 7048 11219
rect 7082 11185 7117 11219
rect 7151 11185 7186 11219
rect 7220 11185 7255 11219
rect 7289 11185 7324 11219
rect 7358 11185 7393 11219
rect 7427 11185 7462 11219
rect 7496 11185 7531 11219
rect 7565 11185 7600 11219
rect 7634 11185 7669 11219
rect 7703 11185 7738 11219
rect 7772 11185 7807 11219
rect 7841 11185 7875 11219
rect 7909 11185 7943 11219
rect 7977 11185 8011 11219
rect 8045 11185 8079 11219
rect 8113 11185 8147 11219
rect 8181 11185 8215 11219
rect 8249 11185 8283 11219
rect 8317 11185 8351 11219
rect 8385 11185 8419 11219
rect 8453 11185 8487 11219
rect 8521 11185 8555 11219
rect 8589 11185 8623 11219
rect 8657 11185 8691 11219
rect 8725 11185 8759 11219
rect 8793 11185 8827 11219
rect 8861 11185 8895 11219
rect 8929 11185 8963 11219
rect 8997 11185 9031 11219
rect 9065 11185 9099 11219
rect 9133 11185 9167 11219
rect 9201 11185 9235 11219
rect 9269 11185 9303 11219
rect 9337 11185 9371 11219
rect 9405 11185 9439 11219
rect 9473 11185 9507 11219
rect 9541 11185 9575 11219
rect 9609 11185 9643 11219
rect 9677 11185 9711 11219
rect 9745 11185 9779 11219
rect 9813 11185 9847 11219
rect 9881 11185 9915 11219
rect 9949 11185 9983 11219
rect 10017 11185 10051 11219
rect 10085 11185 10119 11219
rect 10153 11185 10187 11219
rect 10221 11185 10255 11219
rect 10289 11185 10323 11219
rect 10357 11185 10391 11219
rect 10425 11185 10459 11219
rect 10493 11185 10527 11219
rect 10561 11185 10595 11219
rect 10629 11185 10663 11219
rect 10697 11185 10731 11219
rect 10765 11185 10799 11219
rect 10833 11185 10867 11219
rect 10901 11185 10935 11219
rect 10969 11185 11003 11219
rect 11037 11185 11071 11219
rect 11105 11185 11139 11219
rect 11173 11185 11207 11219
rect 11241 11185 11275 11219
rect 11309 11185 11343 11219
rect 11377 11185 11411 11219
rect 11445 11185 11479 11219
rect 11513 11185 11547 11219
rect 11581 11185 11615 11219
rect 11649 11185 11683 11219
rect 11717 11185 11751 11219
rect 11785 11185 11819 11219
rect 11853 11185 11887 11219
rect 11921 11185 11955 11219
rect 11989 11185 12023 11219
rect 12057 11185 12091 11219
rect 12125 11185 12159 11219
rect 12193 11185 12227 11219
rect 12261 11185 12295 11219
rect 12329 11185 12363 11219
rect 12397 11185 12431 11219
rect 12465 11185 12499 11219
rect 12533 11185 12567 11219
rect 12601 11185 12635 11219
rect 12669 11185 12703 11219
rect 12737 11185 12771 11219
rect 12805 11185 12839 11219
rect 12873 11185 12907 11219
rect 12941 11185 12975 11219
rect 13009 11185 13043 11219
rect 13077 11185 13111 11219
rect 13145 11185 13179 11219
rect 13213 11185 13247 11219
rect 13281 11185 13315 11219
rect 13349 11185 13383 11219
rect 13417 11185 13451 11219
rect 13485 11185 13519 11219
rect 13553 11185 13587 11219
rect 13621 11185 13655 11219
rect 13689 11185 13723 11219
rect 13757 11185 13791 11219
rect 13825 11185 13859 11219
rect 13893 11185 13927 11219
rect 13961 11185 13995 11219
rect 14029 11185 14063 11219
rect 14097 11185 14131 11219
rect 14165 11185 14199 11219
rect 14233 11185 14267 11219
rect 14301 11185 14335 11219
rect 14369 11185 14403 11219
rect 14437 11185 14471 11219
rect 14505 11185 14539 11219
rect 14573 11185 14607 11219
rect 14641 11185 14675 11219
rect 14709 11185 14743 11219
rect 14777 11185 14811 11219
rect 14845 11185 14879 11219
rect 14913 11185 14947 11219
rect 14981 11185 15015 11219
rect 15049 11185 15083 11219
rect 15117 11185 15151 11219
rect 15185 11185 15219 11219
rect 15253 11185 15287 11219
rect 15321 11185 15355 11219
rect 15389 11185 15423 11219
rect 15457 11185 15491 11219
rect 15525 11185 15578 11219
rect 5753 11181 15578 11185
rect 5753 11166 5782 11181
rect 5685 11160 5782 11166
rect 5617 11157 5782 11160
rect 5554 11130 5782 11157
rect 5554 11124 5719 11130
rect 5554 11121 5651 11124
rect 5554 11087 5583 11121
rect 5617 11090 5651 11121
rect 5685 11096 5719 11124
rect 5753 11096 5782 11130
rect 5685 11090 5782 11096
rect 5617 11087 5782 11090
rect 5554 11060 5782 11087
rect 5554 11054 5719 11060
rect 5554 11051 5651 11054
rect 5554 11017 5583 11051
rect 5617 11020 5651 11051
rect 5685 11026 5719 11054
rect 5753 11026 5782 11060
rect 5685 11020 5782 11026
rect 5617 11017 5782 11020
rect 5554 10990 5782 11017
rect 5554 10984 5719 10990
rect 5554 10981 5651 10984
rect 5554 10947 5583 10981
rect 5617 10950 5651 10981
rect 5685 10956 5719 10984
rect 5753 10956 5782 10990
rect 5685 10950 5782 10956
rect 5617 10947 5782 10950
rect 5554 10920 5782 10947
rect 5554 10914 5719 10920
rect 5554 10911 5651 10914
rect 5554 10877 5583 10911
rect 5617 10880 5651 10911
rect 5685 10886 5719 10914
rect 5753 10886 5782 10920
rect 5685 10880 5782 10886
rect 5617 10877 5782 10880
rect 5554 10850 5782 10877
rect 5554 10844 5719 10850
rect 5554 10841 5651 10844
rect 5554 10807 5583 10841
rect 5617 10810 5651 10841
rect 5685 10816 5719 10844
rect 5753 10816 5782 10850
rect 5685 10810 5782 10816
rect 5617 10807 5782 10810
rect 5554 10780 5782 10807
rect 5554 10774 5719 10780
rect 5554 10771 5651 10774
rect 5554 10737 5583 10771
rect 5617 10740 5651 10771
rect 5685 10746 5719 10774
rect 5753 10746 5782 10780
rect 5685 10740 5782 10746
rect 5617 10737 5782 10740
rect 5554 10710 5782 10737
rect 5554 10704 5719 10710
rect 5554 10701 5651 10704
rect 5554 10667 5583 10701
rect 5617 10670 5651 10701
rect 5685 10676 5719 10704
rect 5753 10676 5782 10710
rect 5685 10670 5782 10676
rect 5617 10667 5782 10670
rect 5554 10640 5782 10667
rect 5554 10634 5719 10640
rect 5554 10631 5651 10634
rect 5554 10597 5583 10631
rect 5617 10600 5651 10631
rect 5685 10606 5719 10634
rect 5753 10606 5782 10640
rect 5685 10600 5782 10606
rect 5617 10597 5782 10600
rect 5554 10570 5782 10597
rect 5554 10568 5719 10570
rect 5753 10568 5782 10570
rect 15549 9754 15578 11181
rect 15549 9749 15714 9754
rect 15748 9749 15777 11823
rect 15549 9719 15777 9749
rect 15549 9685 15578 9719
rect 15612 9685 15646 9719
rect 15680 9715 15777 9719
rect 15680 9685 15714 9715
rect 15549 9681 15714 9685
rect 15748 9681 15777 9715
rect 15549 9650 15777 9681
rect 15549 9616 15578 9650
rect 15612 9616 15646 9650
rect 15680 9647 15777 9650
rect 15680 9616 15714 9647
rect 15549 9613 15714 9616
rect 15748 9613 15777 9647
rect 15549 9581 15777 9613
rect 15549 9547 15578 9581
rect 15612 9547 15646 9581
rect 15680 9579 15777 9581
rect 15680 9547 15714 9579
rect 15549 9545 15714 9547
rect 15748 9545 15777 9579
rect 15549 9512 15777 9545
rect 15549 9478 15578 9512
rect 15612 9478 15646 9512
rect 15680 9511 15777 9512
rect 15680 9478 15714 9511
rect 15549 9477 15714 9478
rect 15748 9477 15777 9511
rect 15549 9443 15777 9477
rect 15549 9409 15578 9443
rect 15612 9409 15646 9443
rect 15680 9409 15714 9443
rect 15748 9409 15777 9443
rect 15549 9374 15777 9409
rect 15549 9340 15578 9374
rect 15612 9340 15646 9374
rect 15680 9340 15714 9374
rect 15748 9340 15777 9374
rect 15549 9305 15777 9340
rect 15549 9271 15578 9305
rect 15612 9271 15646 9305
rect 15680 9271 15714 9305
rect 15748 9271 15777 9305
rect 15549 9236 15777 9271
rect 15549 9202 15578 9236
rect 15612 9202 15646 9236
rect 15680 9202 15714 9236
rect 15748 9202 15777 9236
rect 15549 9167 15777 9202
rect 15549 9133 15578 9167
rect 15612 9133 15646 9167
rect 15680 9133 15714 9167
rect 15748 9133 15777 9167
rect 15549 9098 15777 9133
rect 15549 9064 15578 9098
rect 15612 9064 15646 9098
rect 15680 9064 15714 9098
rect 15748 9064 15777 9098
rect 15549 9029 15777 9064
rect 15549 8995 15578 9029
rect 15612 8995 15646 9029
rect 15680 8995 15714 9029
rect 15748 8995 15777 9029
rect 15549 8960 15777 8995
rect 15549 8926 15578 8960
rect 15612 8926 15646 8960
rect 15680 8926 15714 8960
rect 15748 8926 15777 8960
rect 15549 8891 15777 8926
rect 15549 8857 15578 8891
rect 15612 8857 15646 8891
rect 15680 8857 15714 8891
rect 15748 8857 15777 8891
rect 15549 8822 15777 8857
rect 15549 8788 15578 8822
rect 15612 8788 15646 8822
rect 15680 8788 15714 8822
rect 15748 8788 15777 8822
rect 15549 8753 15777 8788
rect 15549 8719 15578 8753
rect 15612 8719 15646 8753
rect 15680 8719 15714 8753
rect 15748 8719 15777 8753
rect 15549 8684 15777 8719
rect 15549 8650 15578 8684
rect 15612 8650 15646 8684
rect 15680 8650 15714 8684
rect 15748 8650 15777 8684
rect 15549 8615 15777 8650
rect 15549 8581 15578 8615
rect 15612 8581 15646 8615
rect 15680 8581 15714 8615
rect 15748 8581 15777 8615
rect 15549 8546 15777 8581
rect 15549 8512 15578 8546
rect 15612 8512 15646 8546
rect 15680 8512 15714 8546
rect 15748 8512 15777 8546
rect 15549 8477 15777 8512
rect 15549 8443 15578 8477
rect 15612 8443 15646 8477
rect 15680 8443 15714 8477
rect 15748 8443 15777 8477
rect 15549 8408 15777 8443
rect 15549 8374 15578 8408
rect 15612 8374 15646 8408
rect 15680 8374 15714 8408
rect 15748 8374 15777 8408
rect 15549 8339 15777 8374
rect 15549 8305 15578 8339
rect 15612 8305 15646 8339
rect 15680 8305 15714 8339
rect 15748 8305 15777 8339
rect 15549 8270 15777 8305
rect 15549 8236 15578 8270
rect 15612 8236 15646 8270
rect 15680 8236 15714 8270
rect 15748 8236 15777 8270
rect 15549 8201 15777 8236
rect 15549 8167 15578 8201
rect 15612 8167 15646 8201
rect 15680 8167 15714 8201
rect 15748 8167 15777 8201
rect 15549 8132 15777 8167
rect 15549 8098 15578 8132
rect 15612 8098 15646 8132
rect 15680 8098 15714 8132
rect 15748 8098 15777 8132
rect 15549 8063 15777 8098
rect 15549 8029 15578 8063
rect 15612 8029 15646 8063
rect 15680 8029 15714 8063
rect 15748 8029 15777 8063
rect 15549 7994 15777 8029
rect 15549 7960 15578 7994
rect 15612 7960 15646 7994
rect 15680 7960 15714 7994
rect 15748 7960 15777 7994
rect 15549 7925 15777 7960
rect 15549 7891 15578 7925
rect 15612 7891 15646 7925
rect 15680 7891 15714 7925
rect 15748 7891 15777 7925
rect 15549 7856 15777 7891
rect 15549 7822 15578 7856
rect 15612 7822 15646 7856
rect 15680 7822 15714 7856
rect 15748 7822 15777 7856
rect 15549 7787 15777 7822
rect 15549 7753 15578 7787
rect 15612 7753 15646 7787
rect 15680 7753 15714 7787
rect 15748 7753 15777 7787
rect 15549 7718 15777 7753
rect 15549 7684 15578 7718
rect 15612 7684 15646 7718
rect 15680 7684 15714 7718
rect 15748 7684 15777 7718
rect 15549 7649 15777 7684
rect 15549 7615 15578 7649
rect 15612 7615 15646 7649
rect 15680 7615 15714 7649
rect 15748 7615 15777 7649
rect 15549 7580 15777 7615
rect 15549 7546 15578 7580
rect 15612 7546 15646 7580
rect 15680 7546 15714 7580
rect 15748 7546 15777 7580
rect 15549 7511 15777 7546
rect 15549 7477 15578 7511
rect 15612 7477 15646 7511
rect 15680 7477 15714 7511
rect 15748 7477 15777 7511
rect 15549 7442 15777 7477
rect 15549 7408 15578 7442
rect 15612 7408 15646 7442
rect 15680 7408 15714 7442
rect 15748 7408 15777 7442
rect 15549 7373 15777 7408
rect 15549 7339 15578 7373
rect 15612 7339 15646 7373
rect 15680 7339 15714 7373
rect 15748 7339 15777 7373
rect 15549 7304 15777 7339
rect 15549 7270 15578 7304
rect 15612 7270 15646 7304
rect 15680 7270 15714 7304
rect 15748 7270 15777 7304
rect 15549 7235 15777 7270
rect 15549 7201 15578 7235
rect 15612 7201 15646 7235
rect 15680 7201 15714 7235
rect 15748 7201 15777 7235
rect 15549 7166 15777 7201
rect 15549 7132 15578 7166
rect 15612 7132 15646 7166
rect 15680 7132 15714 7166
rect 15748 7132 15777 7166
rect 15549 7097 15777 7132
rect 15549 7063 15578 7097
rect 15612 7063 15646 7097
rect 15680 7063 15714 7097
rect 15748 7063 15777 7097
rect 15549 7028 15777 7063
rect 15549 6994 15578 7028
rect 15612 6994 15646 7028
rect 15680 6994 15714 7028
rect 15748 6994 15777 7028
rect 15549 6959 15777 6994
rect 15549 6925 15578 6959
rect 15612 6925 15646 6959
rect 15680 6925 15714 6959
rect 15748 6925 15777 6959
rect 15549 6890 15777 6925
rect 15549 6856 15578 6890
rect 15612 6856 15646 6890
rect 15680 6856 15714 6890
rect 15748 6856 15777 6890
rect 15549 6821 15777 6856
rect 15549 6787 15578 6821
rect 15612 6787 15646 6821
rect 15680 6787 15714 6821
rect 15748 6787 15777 6821
rect 15549 6752 15777 6787
rect 15549 6718 15578 6752
rect 15612 6718 15646 6752
rect 15680 6718 15714 6752
rect 15748 6718 15777 6752
rect 15549 6683 15777 6718
rect 15549 6649 15578 6683
rect 15612 6649 15646 6683
rect 15680 6649 15714 6683
rect 15748 6649 15777 6683
rect 15549 6614 15777 6649
rect 15549 6580 15578 6614
rect 15612 6580 15646 6614
rect 15680 6580 15714 6614
rect 15748 6580 15777 6614
rect 15549 6545 15777 6580
rect 15549 6511 15578 6545
rect 15612 6511 15646 6545
rect 15680 6511 15714 6545
rect 15748 6511 15777 6545
rect 15549 6476 15777 6511
rect 15549 6442 15578 6476
rect 15612 6442 15646 6476
rect 15680 6442 15714 6476
rect 15748 6442 15777 6476
rect 15549 6407 15777 6442
rect 15549 6373 15578 6407
rect 15612 6373 15646 6407
rect 15680 6373 15714 6407
rect 15748 6373 15777 6407
rect 15549 6338 15777 6373
rect 15549 6304 15578 6338
rect 15612 6304 15646 6338
rect 15680 6304 15714 6338
rect 15748 6304 15777 6338
rect 15549 6269 15777 6304
rect 15549 6235 15578 6269
rect 15612 6235 15646 6269
rect 15680 6235 15714 6269
rect 15748 6235 15777 6269
rect 15549 6200 15777 6235
rect 15549 6166 15578 6200
rect 15612 6166 15646 6200
rect 15680 6166 15714 6200
rect 15748 6166 15777 6200
rect 15549 6131 15777 6166
rect 15549 6097 15578 6131
rect 15612 6097 15646 6131
rect 15680 6097 15714 6131
rect 15748 6097 15777 6131
rect 15549 6062 15777 6097
rect 15549 6028 15578 6062
rect 15612 6028 15646 6062
rect 15680 6028 15714 6062
rect 15748 6028 15777 6062
rect 15549 5993 15777 6028
rect 15549 5959 15578 5993
rect 15612 5959 15646 5993
rect 15680 5959 15714 5993
rect 15748 5959 15777 5993
rect 15549 5924 15777 5959
rect 15549 5890 15578 5924
rect 15612 5890 15646 5924
rect 15680 5890 15714 5924
rect 15748 5890 15777 5924
rect 15549 5855 15777 5890
rect 15549 5821 15578 5855
rect 15612 5821 15646 5855
rect 15680 5821 15714 5855
rect 15748 5821 15777 5855
rect 15549 5786 15777 5821
rect 15549 5752 15578 5786
rect 15612 5752 15646 5786
rect 15680 5752 15714 5786
rect 15748 5752 15777 5786
rect 15549 5717 15777 5752
rect 15549 5683 15578 5717
rect 15612 5683 15646 5717
rect 15680 5683 15714 5717
rect 15748 5683 15777 5717
rect 15549 5648 15777 5683
rect 15549 5614 15578 5648
rect 15612 5614 15646 5648
rect 15680 5614 15714 5648
rect 15748 5614 15777 5648
rect 15549 5579 15777 5614
rect 15549 5545 15578 5579
rect 15612 5545 15646 5579
rect 15680 5545 15714 5579
rect 15748 5545 15777 5579
rect 15549 5510 15777 5545
rect 15549 5476 15578 5510
rect 15612 5476 15646 5510
rect 15680 5476 15714 5510
rect 15748 5476 15777 5510
rect 15549 5441 15777 5476
rect 15549 5407 15578 5441
rect 15612 5407 15646 5441
rect 15680 5407 15714 5441
rect 15748 5407 15777 5441
rect 15549 5372 15777 5407
rect 15549 5338 15578 5372
rect 15612 5338 15646 5372
rect 15680 5338 15714 5372
rect 15748 5338 15777 5372
rect 15549 5303 15777 5338
rect 15549 5269 15578 5303
rect 15612 5269 15646 5303
rect 15680 5269 15714 5303
rect 15748 5269 15777 5303
rect 15549 5234 15777 5269
rect 15549 5200 15578 5234
rect 15612 5200 15646 5234
rect 15680 5200 15714 5234
rect 15748 5200 15777 5234
rect 15549 5165 15777 5200
rect 15549 5131 15578 5165
rect 15612 5131 15646 5165
rect 15680 5131 15714 5165
rect 15748 5131 15777 5165
rect 15549 5107 15777 5131
rect 12425 2524 12538 2558
<< mvpsubdiff >>
rect 5554 10564 5719 10568
rect 5554 10561 5651 10564
rect 5554 10527 5583 10561
rect 5617 10530 5651 10561
rect 5685 10536 5719 10564
rect 5753 10536 5782 10568
rect 5685 10530 5782 10536
rect 5617 10527 5782 10530
rect 5554 10521 5782 10527
rect -76 10500 5782 10521
rect -76 10494 5719 10500
rect -76 10492 5651 10494
rect -76 10322 -52 10492
rect 1546 10458 1581 10492
rect 1615 10458 1650 10492
rect 1684 10458 1719 10492
rect 1753 10458 1788 10492
rect 1822 10458 1857 10492
rect 1891 10458 1926 10492
rect 1960 10458 1995 10492
rect 2029 10458 2064 10492
rect 2098 10458 2133 10492
rect 2167 10458 2202 10492
rect 2236 10458 2271 10492
rect 2305 10458 2340 10492
rect 2374 10458 2409 10492
rect 2443 10458 2478 10492
rect 2512 10458 2547 10492
rect 2581 10458 2616 10492
rect 2650 10458 2685 10492
rect 2719 10458 2754 10492
rect 2788 10458 2823 10492
rect 2857 10458 2892 10492
rect 2926 10458 2961 10492
rect 2995 10458 3030 10492
rect 3064 10458 3099 10492
rect 3133 10458 3168 10492
rect 3202 10458 3237 10492
rect 3271 10458 3306 10492
rect 3340 10458 3375 10492
rect 3409 10458 3444 10492
rect 3478 10458 3513 10492
rect 3547 10458 3582 10492
rect 3616 10458 3651 10492
rect 3685 10458 3720 10492
rect 3754 10458 3789 10492
rect 3823 10458 3858 10492
rect 3892 10458 3927 10492
rect 3961 10458 3996 10492
rect 4030 10458 4065 10492
rect 4099 10458 4134 10492
rect 4168 10458 4203 10492
rect 4237 10458 4272 10492
rect 4306 10458 4341 10492
rect 4375 10458 4410 10492
rect 4444 10458 4479 10492
rect 4513 10458 4548 10492
rect 4582 10458 4617 10492
rect 4651 10458 4686 10492
rect 4720 10458 4755 10492
rect 4789 10458 4824 10492
rect 4858 10458 4893 10492
rect 4927 10458 4962 10492
rect 4996 10458 5031 10492
rect 5065 10458 5100 10492
rect 5134 10458 5169 10492
rect 5203 10458 5238 10492
rect 5272 10458 5307 10492
rect 5341 10458 5376 10492
rect 5410 10458 5445 10492
rect 5479 10458 5514 10492
rect 5548 10458 5583 10492
rect 5617 10460 5651 10492
rect 5685 10466 5719 10494
rect 5753 10466 5782 10500
rect 5685 10460 5782 10466
rect 5617 10458 5782 10460
rect 1546 10431 5782 10458
rect 1546 10424 5719 10431
rect 1614 10390 1649 10424
rect 1683 10390 1718 10424
rect 1752 10390 1787 10424
rect 1821 10390 1856 10424
rect 1890 10390 1925 10424
rect 1959 10390 1994 10424
rect 2028 10390 2063 10424
rect 2097 10390 2132 10424
rect 2166 10390 2201 10424
rect 2235 10390 2270 10424
rect 2304 10390 2339 10424
rect 2373 10390 2408 10424
rect 2442 10390 2477 10424
rect 2511 10390 2546 10424
rect 2580 10390 2615 10424
rect 2649 10390 2684 10424
rect 2718 10390 2753 10424
rect 2787 10390 2822 10424
rect 2856 10390 2891 10424
rect 2925 10390 2960 10424
rect 2994 10390 3029 10424
rect 3063 10390 3098 10424
rect 3132 10390 3167 10424
rect 3201 10390 3236 10424
rect 3270 10390 3305 10424
rect 3339 10390 3374 10424
rect 3408 10390 3443 10424
rect 3477 10390 3512 10424
rect 3546 10390 3581 10424
rect 3615 10390 3650 10424
rect 3684 10390 3719 10424
rect 3753 10390 3788 10424
rect 3822 10390 3857 10424
rect 3891 10390 3926 10424
rect 3960 10390 3995 10424
rect 4029 10390 4064 10424
rect 4098 10390 4133 10424
rect 4167 10390 4202 10424
rect 4236 10390 4271 10424
rect 4305 10390 4340 10424
rect 4374 10390 4409 10424
rect 4443 10390 4478 10424
rect 4512 10390 4547 10424
rect 4581 10390 4616 10424
rect 4650 10390 4685 10424
rect 4719 10390 4754 10424
rect 4788 10390 4823 10424
rect 4857 10390 4892 10424
rect 4926 10390 4961 10424
rect 4995 10390 5030 10424
rect 5064 10390 5099 10424
rect 5133 10390 5168 10424
rect 5202 10390 5237 10424
rect 5271 10390 5306 10424
rect 5340 10390 5375 10424
rect 5409 10390 5444 10424
rect 5478 10390 5513 10424
rect 5547 10390 5582 10424
rect 5616 10390 5651 10424
rect 5685 10397 5719 10424
rect 5753 10397 5782 10431
rect 5685 10390 5782 10397
rect 1614 10356 5782 10390
rect 1614 10322 1648 10356
rect 1682 10322 1716 10356
rect 1750 10322 1784 10356
rect 1818 10322 1852 10356
rect 1886 10322 1920 10356
rect 1954 10322 1988 10356
rect 2022 10322 2057 10356
rect 2091 10322 2126 10356
rect 2160 10322 2195 10356
rect 2229 10322 2264 10356
rect 2298 10322 2333 10356
rect 2367 10322 2402 10356
rect 2436 10322 2471 10356
rect 2505 10322 2540 10356
rect 2574 10322 2609 10356
rect 2643 10322 2678 10356
rect 2712 10322 2747 10356
rect 2781 10322 2816 10356
rect 2850 10322 2885 10356
rect 2919 10322 2954 10356
rect 2988 10322 3023 10356
rect 3057 10322 3092 10356
rect 3126 10322 3161 10356
rect 3195 10322 3230 10356
rect 3264 10322 3299 10356
rect 3333 10322 3368 10356
rect 3402 10322 3437 10356
rect 3471 10322 3506 10356
rect 3540 10322 3575 10356
rect 3609 10322 3644 10356
rect 3678 10322 3713 10356
rect 3747 10322 3782 10356
rect 3816 10322 3851 10356
rect 3885 10322 3920 10356
rect 3954 10322 3989 10356
rect 4023 10322 4058 10356
rect 4092 10322 4127 10356
rect 4161 10322 4196 10356
rect 4230 10322 4265 10356
rect 4299 10322 4334 10356
rect 4368 10322 4403 10356
rect 4437 10322 4472 10356
rect 4506 10322 4541 10356
rect 4575 10322 4610 10356
rect 4644 10322 4679 10356
rect 4713 10322 4748 10356
rect 4782 10322 4817 10356
rect 4851 10322 4886 10356
rect 4920 10322 4955 10356
rect 4989 10322 5024 10356
rect 5058 10322 5093 10356
rect 5127 10322 5162 10356
rect 5196 10322 5231 10356
rect 5265 10322 5300 10356
rect 5334 10322 5369 10356
rect 5403 10322 5438 10356
rect 5472 10322 5507 10356
rect 5541 10322 5576 10356
rect 5610 10322 5645 10356
rect 5679 10322 5714 10356
rect 5748 10322 5782 10356
rect -76 10293 5782 10322
rect 11612 8281 11663 9102
rect 11612 8232 14634 8281
rect 11612 7524 11684 8232
<< mvnsubdiff >>
rect 12201 10107 12225 10141
rect 12259 10107 12295 10141
rect 12329 10107 12365 10141
rect 12399 10107 12435 10141
rect 12469 10107 12504 10141
rect 12538 10107 12573 10141
rect 12607 10107 12642 10141
rect 12676 10107 12711 10141
rect 12745 10107 12780 10141
rect 12814 10107 12849 10141
rect 12883 10107 12918 10141
rect 12952 10107 12987 10141
rect 13021 10107 13056 10141
rect 13090 10107 13125 10141
rect 13159 10107 13194 10141
rect 13228 10107 13263 10141
rect 13297 10107 13332 10141
rect 13366 10107 13401 10141
rect 13435 10107 13470 10141
rect 13504 10107 13539 10141
rect 13573 10107 13608 10141
rect 13642 10107 13677 10141
rect 13711 10107 13746 10141
rect 13780 10107 13815 10141
rect 13849 10107 13884 10141
rect 13918 10107 13953 10141
rect 13987 10107 14022 10141
rect 14056 10107 14091 10141
rect 14125 10107 14160 10141
rect 14194 10107 14229 10141
rect 14263 10107 14298 10141
rect 14332 10107 14367 10141
rect 14401 10107 14436 10141
rect 14470 10107 14505 10141
rect 14539 10107 14574 10141
rect 14608 10107 14643 10141
rect 14677 10107 14712 10141
rect 14746 10107 14781 10141
rect 14815 10107 14850 10141
rect 14884 10107 14919 10141
rect 14953 10107 14988 10141
rect 15022 10107 15057 10141
rect 15091 10107 15126 10141
rect 15160 10107 15195 10141
rect 15229 10107 15333 10141
rect 15299 10038 15333 10073
rect 15299 9969 15333 10004
rect 15299 9900 15333 9935
rect 15299 9831 15333 9866
rect 15299 9762 15333 9797
rect 15299 9693 15333 9728
rect 15299 9624 15333 9659
rect 15299 9555 15333 9590
rect 15299 9486 15333 9521
rect 15299 9417 15333 9452
rect 15299 9348 15333 9383
rect 15299 9279 15333 9314
rect 15299 9210 15333 9245
rect 15299 9141 15333 9176
rect 15299 9072 15333 9107
rect 15299 9003 15333 9038
rect 15299 8934 15333 8969
rect 15299 8865 15333 8900
rect 15299 8796 15333 8831
rect 15299 8727 15333 8762
rect 15299 8658 15333 8693
rect 15299 8589 15333 8624
rect 15299 8520 15333 8555
rect 15299 8452 15333 8486
rect 15299 8384 15333 8418
rect 15299 8316 15333 8350
rect 15299 8248 15333 8282
rect 15299 8180 15333 8214
rect 15299 8112 15333 8146
rect 15299 8044 15333 8078
rect 15299 7976 15333 8010
rect 15299 7908 15333 7942
rect 14847 7812 14949 7836
rect 14881 7778 14915 7812
rect 14949 7778 15006 7806
rect 14847 7742 15006 7778
rect 15038 7772 15062 7806
rect 15096 7772 15163 7806
rect 15197 7772 15265 7806
rect 15299 7772 15333 7874
rect 14881 7708 14915 7742
rect 14949 7708 15006 7742
rect 14847 7672 15006 7708
rect 14881 7638 14915 7672
rect 14949 7638 15006 7672
rect 14847 7602 15006 7638
rect 14881 7568 14915 7602
rect 14949 7568 15006 7602
rect 14847 7532 15006 7568
rect 14881 7498 14915 7532
rect 14949 7498 15006 7532
rect 14847 7462 15006 7498
rect 14881 7428 14915 7462
rect 14949 7428 15006 7462
rect 14847 7391 15006 7428
rect 14881 7357 14915 7391
rect 14949 7357 15006 7391
rect 14847 7320 15006 7357
rect 14881 7286 14915 7320
rect 14949 7286 15006 7320
rect 14847 7249 15006 7286
rect 14881 7215 14915 7249
rect 14949 7215 15006 7249
rect 14847 7178 15006 7215
rect 14881 7144 14915 7178
rect 14949 7144 15006 7178
rect 14847 7107 15006 7144
rect 14881 7073 14915 7107
rect 14949 7073 15006 7107
rect 14847 7036 15006 7073
rect 14881 7002 14915 7036
rect 14949 7002 15006 7036
rect 14847 6965 15006 7002
rect 14881 6931 14915 6965
rect 14949 6931 15006 6965
rect 14847 6894 15006 6931
rect 14881 6860 14915 6894
rect 14949 6860 15006 6894
rect 14847 6823 15006 6860
rect 14881 6789 14915 6823
rect 14949 6789 15006 6823
rect 14847 6752 15006 6789
rect 14881 6718 14915 6752
rect 14949 6718 15006 6752
rect 14847 6681 15006 6718
rect 14881 6647 14915 6681
rect 14949 6647 15006 6681
rect 14847 6610 15006 6647
rect 14881 6576 14915 6610
rect 14949 6576 15006 6610
rect 14847 6539 15006 6576
rect 14881 6505 14915 6539
rect 14949 6505 15006 6539
rect 14847 6468 15006 6505
rect 14881 6434 14915 6468
rect 14949 6434 15006 6468
rect 14847 6397 15006 6434
rect 14881 6363 14915 6397
rect 14949 6363 15006 6397
rect 14847 6326 15006 6363
rect 14881 6292 14915 6326
rect 14949 6292 15006 6326
rect 14847 6268 15006 6292
rect 14868 6030 15006 6268
<< psubdiffcont >>
rect 5583 11857 5617 11891
rect 5656 11862 11062 11896
rect 11096 11862 11130 11896
rect 11164 11862 11198 11896
rect 11232 11862 11266 11896
rect 11300 11862 11334 11896
rect 11368 11862 11402 11896
rect 11436 11862 11470 11896
rect 11504 11862 11538 11896
rect 11572 11862 11606 11896
rect 11640 11862 11674 11896
rect 11708 11862 11742 11896
rect 11776 11862 11810 11896
rect 11845 11862 11879 11896
rect 11914 11862 11948 11896
rect 11983 11862 12017 11896
rect 12052 11862 12086 11896
rect 12121 11862 12155 11896
rect 12190 11862 12224 11896
rect 12259 11862 12293 11896
rect 12328 11862 12362 11896
rect 12397 11862 12431 11896
rect 12466 11862 12500 11896
rect 12535 11862 12569 11896
rect 12604 11862 12638 11896
rect 12673 11862 12707 11896
rect 12742 11862 12776 11896
rect 12811 11862 12845 11896
rect 12880 11862 12914 11896
rect 12949 11862 12983 11896
rect 13018 11862 13052 11896
rect 13087 11862 13121 11896
rect 13156 11862 13190 11896
rect 13225 11862 13259 11896
rect 13294 11862 13328 11896
rect 13363 11862 13397 11896
rect 13432 11862 13466 11896
rect 13501 11862 13535 11896
rect 13570 11862 13604 11896
rect 13639 11862 13673 11896
rect 13708 11862 13742 11896
rect 13777 11862 13811 11896
rect 13846 11862 13880 11896
rect 13915 11862 13949 11896
rect 13984 11862 14018 11896
rect 14053 11862 14087 11896
rect 14122 11862 14156 11896
rect 14191 11862 14225 11896
rect 14260 11862 14294 11896
rect 14329 11862 14363 11896
rect 14398 11862 14432 11896
rect 14467 11862 14501 11896
rect 14536 11862 14570 11896
rect 14605 11862 14639 11896
rect 14674 11862 14708 11896
rect 14743 11862 14777 11896
rect 14812 11862 14846 11896
rect 14881 11862 14915 11896
rect 14950 11862 14984 11896
rect 15019 11862 15053 11896
rect 15088 11862 15122 11896
rect 15157 11862 15191 11896
rect 15226 11862 15260 11896
rect 15295 11862 15329 11896
rect 15364 11862 15398 11896
rect 15433 11862 15467 11896
rect 15502 11862 15536 11896
rect 15571 11862 15605 11896
rect 15640 11862 15674 11896
rect 15709 11862 15743 11896
rect 5656 11828 11057 11862
rect 5583 11787 5617 11821
rect 5651 11794 11057 11828
rect 11092 11794 11126 11828
rect 11161 11794 11195 11828
rect 11230 11794 11264 11828
rect 11299 11794 11333 11828
rect 11368 11794 11402 11828
rect 11437 11794 11471 11828
rect 11506 11794 11540 11828
rect 11575 11794 11609 11828
rect 11644 11794 11678 11828
rect 11713 11794 11747 11828
rect 11782 11794 11816 11828
rect 11851 11794 11885 11828
rect 11920 11794 11954 11828
rect 11989 11794 12023 11828
rect 12058 11794 12092 11828
rect 12127 11794 12161 11828
rect 12196 11794 12230 11828
rect 12265 11794 12299 11828
rect 12334 11794 12368 11828
rect 12403 11794 12437 11828
rect 12472 11794 12506 11828
rect 12541 11794 12575 11828
rect 12610 11794 12644 11828
rect 12679 11794 12713 11828
rect 12748 11794 12782 11828
rect 12817 11794 12851 11828
rect 12886 11794 12920 11828
rect 12955 11794 12989 11828
rect 13024 11794 13058 11828
rect 13093 11794 13127 11828
rect 13162 11794 13196 11828
rect 13231 11794 13265 11828
rect 13300 11794 13334 11828
rect 13369 11794 13403 11828
rect 13438 11794 13472 11828
rect 13507 11794 13541 11828
rect 13576 11794 13610 11828
rect 13645 11794 13679 11828
rect 13714 11794 13748 11828
rect 13783 11794 13817 11828
rect 13852 11794 13886 11828
rect 13921 11794 13955 11828
rect 13990 11794 14024 11828
rect 14059 11794 14093 11828
rect 14128 11794 14162 11828
rect 14197 11794 14231 11828
rect 14266 11794 14300 11828
rect 14335 11794 14369 11828
rect 14404 11794 14438 11828
rect 14473 11794 14507 11828
rect 14542 11794 14576 11828
rect 14611 11794 14645 11828
rect 14680 11794 14714 11828
rect 14749 11794 14783 11828
rect 14818 11794 14852 11828
rect 14887 11794 14921 11828
rect 14956 11794 14990 11828
rect 15025 11794 15059 11828
rect 15094 11794 15128 11828
rect 15163 11794 15197 11828
rect 15232 11794 15266 11828
rect 15301 11794 15335 11828
rect 15370 11794 15404 11828
rect 15439 11794 15473 11828
rect 15508 11794 15542 11828
rect 15577 11794 15611 11828
rect 15646 11823 15680 11828
rect 5583 11717 5617 11751
rect 5651 11723 5685 11757
rect 5719 11726 10989 11794
rect 15646 11760 15748 11823
rect 11024 11726 11058 11760
rect 11093 11726 11127 11760
rect 11162 11726 11196 11760
rect 11231 11726 11265 11760
rect 11300 11726 11334 11760
rect 11369 11726 11403 11760
rect 11438 11726 11472 11760
rect 11507 11726 11541 11760
rect 11576 11726 11610 11760
rect 11645 11726 11679 11760
rect 11714 11726 11748 11760
rect 11783 11726 11817 11760
rect 11852 11726 11886 11760
rect 11921 11726 11955 11760
rect 11990 11726 12024 11760
rect 12059 11726 12093 11760
rect 12128 11726 12162 11760
rect 12197 11726 12231 11760
rect 12266 11726 12300 11760
rect 12335 11726 12369 11760
rect 12404 11726 12438 11760
rect 12473 11726 12507 11760
rect 12542 11726 12576 11760
rect 12611 11726 12645 11760
rect 12680 11726 12714 11760
rect 12749 11726 12783 11760
rect 12818 11726 12852 11760
rect 12887 11726 12921 11760
rect 12956 11726 12990 11760
rect 13025 11726 13059 11760
rect 13094 11726 13128 11760
rect 13163 11726 13197 11760
rect 13232 11726 13266 11760
rect 13301 11726 13335 11760
rect 13370 11726 13404 11760
rect 13439 11726 13473 11760
rect 13508 11726 13542 11760
rect 13577 11726 13611 11760
rect 13646 11726 13680 11760
rect 13715 11726 13749 11760
rect 13784 11726 13818 11760
rect 13853 11726 13887 11760
rect 13922 11726 13956 11760
rect 13991 11726 14025 11760
rect 14060 11726 14094 11760
rect 14129 11726 14163 11760
rect 14198 11726 14232 11760
rect 14267 11726 14301 11760
rect 14336 11726 14370 11760
rect 14405 11726 14439 11760
rect 14474 11726 14508 11760
rect 14543 11726 14577 11760
rect 14612 11726 14646 11760
rect 14681 11726 14715 11760
rect 14750 11726 14784 11760
rect 14819 11726 14853 11760
rect 14888 11726 14922 11760
rect 14957 11726 14991 11760
rect 15026 11726 15060 11760
rect 15095 11726 15129 11760
rect 15164 11726 15198 11760
rect 15233 11726 15267 11760
rect 15302 11726 15336 11760
rect 15371 11726 15405 11760
rect 15440 11726 15474 11760
rect 15509 11726 15543 11760
rect 5583 11647 5617 11681
rect 5651 11652 5685 11686
rect 5719 11656 5753 11690
rect 5583 11577 5617 11611
rect 5651 11581 5685 11615
rect 5719 11586 5753 11620
rect 5806 11617 5840 11651
rect 5875 11617 5909 11651
rect 5944 11617 5978 11651
rect 6013 11617 6047 11651
rect 6082 11617 6116 11651
rect 6151 11617 6185 11651
rect 6220 11617 6254 11651
rect 6289 11617 6323 11651
rect 6358 11617 6392 11651
rect 6427 11617 6461 11651
rect 6496 11617 6530 11651
rect 6565 11617 6599 11651
rect 6634 11617 6668 11651
rect 6703 11617 6737 11651
rect 6772 11617 6806 11651
rect 6841 11617 6875 11651
rect 6910 11617 6944 11651
rect 6979 11617 7013 11651
rect 7048 11617 7082 11651
rect 7117 11617 7151 11651
rect 7186 11617 7220 11651
rect 7255 11617 7289 11651
rect 7324 11617 7358 11651
rect 7393 11617 7427 11651
rect 7462 11617 7496 11651
rect 7531 11617 7565 11651
rect 7600 11617 7634 11651
rect 7669 11617 7703 11651
rect 7738 11617 7772 11651
rect 7807 11617 7841 11651
rect 7875 11617 7909 11651
rect 7943 11617 7977 11651
rect 8011 11617 8045 11651
rect 8079 11617 8113 11651
rect 8147 11617 8181 11651
rect 8215 11617 8249 11651
rect 8283 11617 8317 11651
rect 8351 11617 8385 11651
rect 8419 11617 8453 11651
rect 8487 11617 8521 11651
rect 8555 11617 8589 11651
rect 8623 11617 8657 11651
rect 8691 11617 8725 11651
rect 8759 11617 8793 11651
rect 8827 11617 8861 11651
rect 8895 11617 8929 11651
rect 8963 11617 8997 11651
rect 9031 11617 9065 11651
rect 9099 11617 9133 11651
rect 9167 11617 9201 11651
rect 9235 11617 9269 11651
rect 9303 11617 9337 11651
rect 9371 11617 9405 11651
rect 9439 11617 9473 11651
rect 9507 11617 9541 11651
rect 9575 11617 9609 11651
rect 9643 11617 9677 11651
rect 9711 11617 9745 11651
rect 9779 11617 9813 11651
rect 9847 11617 9881 11651
rect 9915 11617 9949 11651
rect 9983 11617 10017 11651
rect 10051 11617 10085 11651
rect 10119 11617 10153 11651
rect 10187 11617 10221 11651
rect 10255 11617 10289 11651
rect 10323 11617 10357 11651
rect 10391 11617 10425 11651
rect 10459 11617 10493 11651
rect 10527 11617 10561 11651
rect 10595 11617 10629 11651
rect 10663 11617 10697 11651
rect 10731 11617 10765 11651
rect 10799 11617 10833 11651
rect 10867 11617 10901 11651
rect 10935 11617 10969 11651
rect 11003 11617 11037 11651
rect 11071 11617 11105 11651
rect 11139 11617 11173 11651
rect 11207 11617 11241 11651
rect 11275 11617 11309 11651
rect 11343 11617 11377 11651
rect 11411 11617 11445 11651
rect 11479 11617 11513 11651
rect 11547 11617 11581 11651
rect 11615 11617 11649 11651
rect 11683 11617 11717 11651
rect 11751 11617 11785 11651
rect 11819 11617 11853 11651
rect 11887 11617 11921 11651
rect 11955 11617 11989 11651
rect 12023 11617 12057 11651
rect 12091 11617 12125 11651
rect 12159 11617 12193 11651
rect 12227 11617 12261 11651
rect 12295 11617 12329 11651
rect 12363 11617 12397 11651
rect 12431 11617 12465 11651
rect 12499 11617 12533 11651
rect 12567 11617 12601 11651
rect 12635 11617 12669 11651
rect 12703 11617 12737 11651
rect 12771 11617 12805 11651
rect 12839 11617 12873 11651
rect 12907 11617 12941 11651
rect 12975 11617 13009 11651
rect 13043 11617 13077 11651
rect 13111 11617 13145 11651
rect 13179 11617 13213 11651
rect 13247 11617 13281 11651
rect 13315 11617 13349 11651
rect 13383 11617 13417 11651
rect 13451 11617 13485 11651
rect 13519 11617 13553 11651
rect 13587 11617 13621 11651
rect 13655 11617 13689 11651
rect 13723 11617 13757 11651
rect 13791 11617 13825 11651
rect 13859 11617 13893 11651
rect 13927 11617 13961 11651
rect 13995 11617 14029 11651
rect 14063 11617 14097 11651
rect 14131 11617 14165 11651
rect 14199 11617 14233 11651
rect 14267 11617 14301 11651
rect 14335 11617 14369 11651
rect 14403 11617 14437 11651
rect 14471 11617 14505 11651
rect 14539 11617 14573 11651
rect 14607 11617 14641 11651
rect 14675 11617 14709 11651
rect 14743 11617 14777 11651
rect 14811 11617 14845 11651
rect 14879 11617 14913 11651
rect 14947 11617 14981 11651
rect 15015 11617 15049 11651
rect 15083 11617 15117 11651
rect 15151 11617 15185 11651
rect 15219 11617 15253 11651
rect 15287 11617 15321 11651
rect 15355 11617 15389 11651
rect 15423 11617 15457 11651
rect 15491 11617 15525 11651
rect 5583 11507 5617 11541
rect 5651 11510 5685 11544
rect 5719 11516 5753 11550
rect 5806 11545 5840 11579
rect 5875 11545 5909 11579
rect 5944 11545 5978 11579
rect 6013 11545 6047 11579
rect 6082 11545 6116 11579
rect 6151 11545 6185 11579
rect 6220 11545 6254 11579
rect 6289 11545 6323 11579
rect 6358 11545 6392 11579
rect 6427 11545 6461 11579
rect 6496 11545 6530 11579
rect 6565 11545 6599 11579
rect 6634 11545 6668 11579
rect 6703 11545 6737 11579
rect 6772 11545 6806 11579
rect 6841 11545 6875 11579
rect 6910 11545 6944 11579
rect 6979 11545 7013 11579
rect 7048 11545 7082 11579
rect 7117 11545 7151 11579
rect 7186 11545 7220 11579
rect 7255 11545 7289 11579
rect 7324 11545 7358 11579
rect 7393 11545 7427 11579
rect 7462 11545 7496 11579
rect 7531 11545 7565 11579
rect 7600 11545 7634 11579
rect 7669 11545 7703 11579
rect 7738 11545 7772 11579
rect 7807 11545 7841 11579
rect 7875 11545 7909 11579
rect 7943 11545 7977 11579
rect 8011 11545 8045 11579
rect 8079 11545 8113 11579
rect 8147 11545 8181 11579
rect 8215 11545 8249 11579
rect 8283 11545 8317 11579
rect 8351 11545 8385 11579
rect 8419 11545 8453 11579
rect 8487 11545 8521 11579
rect 8555 11545 8589 11579
rect 8623 11545 8657 11579
rect 8691 11545 8725 11579
rect 8759 11545 8793 11579
rect 8827 11545 8861 11579
rect 8895 11545 8929 11579
rect 8963 11545 8997 11579
rect 9031 11545 9065 11579
rect 9099 11545 9133 11579
rect 9167 11545 9201 11579
rect 9235 11545 9269 11579
rect 9303 11545 9337 11579
rect 9371 11545 9405 11579
rect 9439 11545 9473 11579
rect 9507 11545 9541 11579
rect 9575 11545 9609 11579
rect 9643 11545 9677 11579
rect 9711 11545 9745 11579
rect 9779 11545 9813 11579
rect 9847 11545 9881 11579
rect 9915 11545 9949 11579
rect 9983 11545 10017 11579
rect 10051 11545 10085 11579
rect 10119 11545 10153 11579
rect 10187 11545 10221 11579
rect 10255 11545 10289 11579
rect 10323 11545 10357 11579
rect 10391 11545 10425 11579
rect 10459 11545 10493 11579
rect 10527 11545 10561 11579
rect 10595 11545 10629 11579
rect 10663 11545 10697 11579
rect 10731 11545 10765 11579
rect 10799 11545 10833 11579
rect 10867 11545 10901 11579
rect 10935 11545 10969 11579
rect 11003 11545 11037 11579
rect 11071 11545 11105 11579
rect 11139 11545 11173 11579
rect 11207 11545 11241 11579
rect 11275 11545 11309 11579
rect 11343 11545 11377 11579
rect 11411 11545 11445 11579
rect 11479 11545 11513 11579
rect 11547 11545 11581 11579
rect 11615 11545 11649 11579
rect 11683 11545 11717 11579
rect 11751 11545 11785 11579
rect 11819 11545 11853 11579
rect 11887 11545 11921 11579
rect 11955 11545 11989 11579
rect 12023 11545 12057 11579
rect 12091 11545 12125 11579
rect 12159 11545 12193 11579
rect 12227 11545 12261 11579
rect 12295 11545 12329 11579
rect 12363 11545 12397 11579
rect 12431 11545 12465 11579
rect 12499 11545 12533 11579
rect 12567 11545 12601 11579
rect 12635 11545 12669 11579
rect 12703 11545 12737 11579
rect 12771 11545 12805 11579
rect 12839 11545 12873 11579
rect 12907 11545 12941 11579
rect 12975 11545 13009 11579
rect 13043 11545 13077 11579
rect 13111 11545 13145 11579
rect 13179 11545 13213 11579
rect 13247 11545 13281 11579
rect 13315 11545 13349 11579
rect 13383 11545 13417 11579
rect 13451 11545 13485 11579
rect 13519 11545 13553 11579
rect 13587 11545 13621 11579
rect 13655 11545 13689 11579
rect 13723 11545 13757 11579
rect 13791 11545 13825 11579
rect 13859 11545 13893 11579
rect 13927 11545 13961 11579
rect 13995 11545 14029 11579
rect 14063 11545 14097 11579
rect 14131 11545 14165 11579
rect 14199 11545 14233 11579
rect 14267 11545 14301 11579
rect 14335 11545 14369 11579
rect 14403 11545 14437 11579
rect 14471 11545 14505 11579
rect 14539 11545 14573 11579
rect 14607 11545 14641 11579
rect 14675 11545 14709 11579
rect 14743 11545 14777 11579
rect 14811 11545 14845 11579
rect 14879 11545 14913 11579
rect 14947 11545 14981 11579
rect 15015 11545 15049 11579
rect 15083 11545 15117 11579
rect 15151 11545 15185 11579
rect 15219 11545 15253 11579
rect 15287 11545 15321 11579
rect 15355 11545 15389 11579
rect 15423 11545 15457 11579
rect 15491 11545 15525 11579
rect 5583 11437 5617 11471
rect 5651 11440 5685 11474
rect 5719 11446 5753 11480
rect 5806 11473 5840 11507
rect 5875 11473 5909 11507
rect 5944 11473 5978 11507
rect 6013 11473 6047 11507
rect 6082 11473 6116 11507
rect 6151 11473 6185 11507
rect 6220 11473 6254 11507
rect 6289 11473 6323 11507
rect 6358 11473 6392 11507
rect 6427 11473 6461 11507
rect 6496 11473 6530 11507
rect 6565 11473 6599 11507
rect 6634 11473 6668 11507
rect 6703 11473 6737 11507
rect 6772 11473 6806 11507
rect 6841 11473 6875 11507
rect 6910 11473 6944 11507
rect 6979 11473 7013 11507
rect 7048 11473 7082 11507
rect 7117 11473 7151 11507
rect 7186 11473 7220 11507
rect 7255 11473 7289 11507
rect 7324 11473 7358 11507
rect 7393 11473 7427 11507
rect 7462 11473 7496 11507
rect 7531 11473 7565 11507
rect 7600 11473 7634 11507
rect 7669 11473 7703 11507
rect 7738 11473 7772 11507
rect 7807 11473 7841 11507
rect 7875 11473 7909 11507
rect 7943 11473 7977 11507
rect 8011 11473 8045 11507
rect 8079 11473 8113 11507
rect 8147 11473 8181 11507
rect 8215 11473 8249 11507
rect 8283 11473 8317 11507
rect 8351 11473 8385 11507
rect 8419 11473 8453 11507
rect 8487 11473 8521 11507
rect 8555 11473 8589 11507
rect 8623 11473 8657 11507
rect 8691 11473 8725 11507
rect 8759 11473 8793 11507
rect 8827 11473 8861 11507
rect 8895 11473 8929 11507
rect 8963 11473 8997 11507
rect 9031 11473 9065 11507
rect 9099 11473 9133 11507
rect 9167 11473 9201 11507
rect 9235 11473 9269 11507
rect 9303 11473 9337 11507
rect 9371 11473 9405 11507
rect 9439 11473 9473 11507
rect 9507 11473 9541 11507
rect 9575 11473 9609 11507
rect 9643 11473 9677 11507
rect 9711 11473 9745 11507
rect 9779 11473 9813 11507
rect 9847 11473 9881 11507
rect 9915 11473 9949 11507
rect 9983 11473 10017 11507
rect 10051 11473 10085 11507
rect 10119 11473 10153 11507
rect 10187 11473 10221 11507
rect 10255 11473 10289 11507
rect 10323 11473 10357 11507
rect 10391 11473 10425 11507
rect 10459 11473 10493 11507
rect 10527 11473 10561 11507
rect 10595 11473 10629 11507
rect 10663 11473 10697 11507
rect 10731 11473 10765 11507
rect 10799 11473 10833 11507
rect 10867 11473 10901 11507
rect 10935 11473 10969 11507
rect 11003 11473 11037 11507
rect 11071 11473 11105 11507
rect 11139 11473 11173 11507
rect 11207 11473 11241 11507
rect 11275 11473 11309 11507
rect 11343 11473 11377 11507
rect 11411 11473 11445 11507
rect 11479 11473 11513 11507
rect 11547 11473 11581 11507
rect 11615 11473 11649 11507
rect 11683 11473 11717 11507
rect 11751 11473 11785 11507
rect 11819 11473 11853 11507
rect 11887 11473 11921 11507
rect 11955 11473 11989 11507
rect 12023 11473 12057 11507
rect 12091 11473 12125 11507
rect 12159 11473 12193 11507
rect 12227 11473 12261 11507
rect 12295 11473 12329 11507
rect 12363 11473 12397 11507
rect 12431 11473 12465 11507
rect 12499 11473 12533 11507
rect 12567 11473 12601 11507
rect 12635 11473 12669 11507
rect 12703 11473 12737 11507
rect 12771 11473 12805 11507
rect 12839 11473 12873 11507
rect 12907 11473 12941 11507
rect 12975 11473 13009 11507
rect 13043 11473 13077 11507
rect 13111 11473 13145 11507
rect 13179 11473 13213 11507
rect 13247 11473 13281 11507
rect 13315 11473 13349 11507
rect 13383 11473 13417 11507
rect 13451 11473 13485 11507
rect 13519 11473 13553 11507
rect 13587 11473 13621 11507
rect 13655 11473 13689 11507
rect 13723 11473 13757 11507
rect 13791 11473 13825 11507
rect 13859 11473 13893 11507
rect 13927 11473 13961 11507
rect 13995 11473 14029 11507
rect 14063 11473 14097 11507
rect 14131 11473 14165 11507
rect 14199 11473 14233 11507
rect 14267 11473 14301 11507
rect 14335 11473 14369 11507
rect 14403 11473 14437 11507
rect 14471 11473 14505 11507
rect 14539 11473 14573 11507
rect 14607 11473 14641 11507
rect 14675 11473 14709 11507
rect 14743 11473 14777 11507
rect 14811 11473 14845 11507
rect 14879 11473 14913 11507
rect 14947 11473 14981 11507
rect 15015 11473 15049 11507
rect 15083 11473 15117 11507
rect 15151 11473 15185 11507
rect 15219 11473 15253 11507
rect 15287 11473 15321 11507
rect 15355 11473 15389 11507
rect 15423 11473 15457 11507
rect 15491 11473 15525 11507
rect 5583 11367 5617 11401
rect 5651 11370 5685 11404
rect 5719 11376 5753 11410
rect 5806 11401 5840 11435
rect 5875 11401 5909 11435
rect 5944 11401 5978 11435
rect 6013 11401 6047 11435
rect 6082 11401 6116 11435
rect 6151 11401 6185 11435
rect 6220 11401 6254 11435
rect 6289 11401 6323 11435
rect 6358 11401 6392 11435
rect 6427 11401 6461 11435
rect 6496 11401 6530 11435
rect 6565 11401 6599 11435
rect 6634 11401 6668 11435
rect 6703 11401 6737 11435
rect 6772 11401 6806 11435
rect 6841 11401 6875 11435
rect 6910 11401 6944 11435
rect 6979 11401 7013 11435
rect 7048 11401 7082 11435
rect 7117 11401 7151 11435
rect 7186 11401 7220 11435
rect 7255 11401 7289 11435
rect 7324 11401 7358 11435
rect 7393 11401 7427 11435
rect 7462 11401 7496 11435
rect 7531 11401 7565 11435
rect 7600 11401 7634 11435
rect 7669 11401 7703 11435
rect 7738 11401 7772 11435
rect 7807 11401 7841 11435
rect 7875 11401 7909 11435
rect 7943 11401 7977 11435
rect 8011 11401 8045 11435
rect 8079 11401 8113 11435
rect 8147 11401 8181 11435
rect 8215 11401 8249 11435
rect 8283 11401 8317 11435
rect 8351 11401 8385 11435
rect 8419 11401 8453 11435
rect 8487 11401 8521 11435
rect 8555 11401 8589 11435
rect 8623 11401 8657 11435
rect 8691 11401 8725 11435
rect 8759 11401 8793 11435
rect 8827 11401 8861 11435
rect 8895 11401 8929 11435
rect 8963 11401 8997 11435
rect 9031 11401 9065 11435
rect 9099 11401 9133 11435
rect 9167 11401 9201 11435
rect 9235 11401 9269 11435
rect 9303 11401 9337 11435
rect 9371 11401 9405 11435
rect 9439 11401 9473 11435
rect 9507 11401 9541 11435
rect 9575 11401 9609 11435
rect 9643 11401 9677 11435
rect 9711 11401 9745 11435
rect 9779 11401 9813 11435
rect 9847 11401 9881 11435
rect 9915 11401 9949 11435
rect 9983 11401 10017 11435
rect 10051 11401 10085 11435
rect 10119 11401 10153 11435
rect 10187 11401 10221 11435
rect 10255 11401 10289 11435
rect 10323 11401 10357 11435
rect 10391 11401 10425 11435
rect 10459 11401 10493 11435
rect 10527 11401 10561 11435
rect 10595 11401 10629 11435
rect 10663 11401 10697 11435
rect 10731 11401 10765 11435
rect 10799 11401 10833 11435
rect 10867 11401 10901 11435
rect 10935 11401 10969 11435
rect 11003 11401 11037 11435
rect 11071 11401 11105 11435
rect 11139 11401 11173 11435
rect 11207 11401 11241 11435
rect 11275 11401 11309 11435
rect 11343 11401 11377 11435
rect 11411 11401 11445 11435
rect 11479 11401 11513 11435
rect 11547 11401 11581 11435
rect 11615 11401 11649 11435
rect 11683 11401 11717 11435
rect 11751 11401 11785 11435
rect 11819 11401 11853 11435
rect 11887 11401 11921 11435
rect 11955 11401 11989 11435
rect 12023 11401 12057 11435
rect 12091 11401 12125 11435
rect 12159 11401 12193 11435
rect 12227 11401 12261 11435
rect 12295 11401 12329 11435
rect 12363 11401 12397 11435
rect 12431 11401 12465 11435
rect 12499 11401 12533 11435
rect 12567 11401 12601 11435
rect 12635 11401 12669 11435
rect 12703 11401 12737 11435
rect 12771 11401 12805 11435
rect 12839 11401 12873 11435
rect 12907 11401 12941 11435
rect 12975 11401 13009 11435
rect 13043 11401 13077 11435
rect 13111 11401 13145 11435
rect 13179 11401 13213 11435
rect 13247 11401 13281 11435
rect 13315 11401 13349 11435
rect 13383 11401 13417 11435
rect 13451 11401 13485 11435
rect 13519 11401 13553 11435
rect 13587 11401 13621 11435
rect 13655 11401 13689 11435
rect 13723 11401 13757 11435
rect 13791 11401 13825 11435
rect 13859 11401 13893 11435
rect 13927 11401 13961 11435
rect 13995 11401 14029 11435
rect 14063 11401 14097 11435
rect 14131 11401 14165 11435
rect 14199 11401 14233 11435
rect 14267 11401 14301 11435
rect 14335 11401 14369 11435
rect 14403 11401 14437 11435
rect 14471 11401 14505 11435
rect 14539 11401 14573 11435
rect 14607 11401 14641 11435
rect 14675 11401 14709 11435
rect 14743 11401 14777 11435
rect 14811 11401 14845 11435
rect 14879 11401 14913 11435
rect 14947 11401 14981 11435
rect 15015 11401 15049 11435
rect 15083 11401 15117 11435
rect 15151 11401 15185 11435
rect 15219 11401 15253 11435
rect 15287 11401 15321 11435
rect 15355 11401 15389 11435
rect 15423 11401 15457 11435
rect 15491 11401 15525 11435
rect 5583 11297 5617 11331
rect 5651 11300 5685 11334
rect 5719 11306 5753 11340
rect 5806 11329 5840 11363
rect 5875 11329 5909 11363
rect 5944 11329 5978 11363
rect 6013 11329 6047 11363
rect 6082 11329 6116 11363
rect 6151 11329 6185 11363
rect 6220 11329 6254 11363
rect 6289 11329 6323 11363
rect 6358 11329 6392 11363
rect 6427 11329 6461 11363
rect 6496 11329 6530 11363
rect 6565 11329 6599 11363
rect 6634 11329 6668 11363
rect 6703 11329 6737 11363
rect 6772 11329 6806 11363
rect 6841 11329 6875 11363
rect 6910 11329 6944 11363
rect 6979 11329 7013 11363
rect 7048 11329 7082 11363
rect 7117 11329 7151 11363
rect 7186 11329 7220 11363
rect 7255 11329 7289 11363
rect 7324 11329 7358 11363
rect 7393 11329 7427 11363
rect 7462 11329 7496 11363
rect 7531 11329 7565 11363
rect 7600 11329 7634 11363
rect 7669 11329 7703 11363
rect 7738 11329 7772 11363
rect 7807 11329 7841 11363
rect 7875 11329 7909 11363
rect 7943 11329 7977 11363
rect 8011 11329 8045 11363
rect 8079 11329 8113 11363
rect 8147 11329 8181 11363
rect 8215 11329 8249 11363
rect 8283 11329 8317 11363
rect 8351 11329 8385 11363
rect 8419 11329 8453 11363
rect 8487 11329 8521 11363
rect 8555 11329 8589 11363
rect 8623 11329 8657 11363
rect 8691 11329 8725 11363
rect 8759 11329 8793 11363
rect 8827 11329 8861 11363
rect 8895 11329 8929 11363
rect 8963 11329 8997 11363
rect 9031 11329 9065 11363
rect 9099 11329 9133 11363
rect 9167 11329 9201 11363
rect 9235 11329 9269 11363
rect 9303 11329 9337 11363
rect 9371 11329 9405 11363
rect 9439 11329 9473 11363
rect 9507 11329 9541 11363
rect 9575 11329 9609 11363
rect 9643 11329 9677 11363
rect 9711 11329 9745 11363
rect 9779 11329 9813 11363
rect 9847 11329 9881 11363
rect 9915 11329 9949 11363
rect 9983 11329 10017 11363
rect 10051 11329 10085 11363
rect 10119 11329 10153 11363
rect 10187 11329 10221 11363
rect 10255 11329 10289 11363
rect 10323 11329 10357 11363
rect 10391 11329 10425 11363
rect 10459 11329 10493 11363
rect 10527 11329 10561 11363
rect 10595 11329 10629 11363
rect 10663 11329 10697 11363
rect 10731 11329 10765 11363
rect 10799 11329 10833 11363
rect 10867 11329 10901 11363
rect 10935 11329 10969 11363
rect 11003 11329 11037 11363
rect 11071 11329 11105 11363
rect 11139 11329 11173 11363
rect 11207 11329 11241 11363
rect 11275 11329 11309 11363
rect 11343 11329 11377 11363
rect 11411 11329 11445 11363
rect 11479 11329 11513 11363
rect 11547 11329 11581 11363
rect 11615 11329 11649 11363
rect 11683 11329 11717 11363
rect 11751 11329 11785 11363
rect 11819 11329 11853 11363
rect 11887 11329 11921 11363
rect 11955 11329 11989 11363
rect 12023 11329 12057 11363
rect 12091 11329 12125 11363
rect 12159 11329 12193 11363
rect 12227 11329 12261 11363
rect 12295 11329 12329 11363
rect 12363 11329 12397 11363
rect 12431 11329 12465 11363
rect 12499 11329 12533 11363
rect 12567 11329 12601 11363
rect 12635 11329 12669 11363
rect 12703 11329 12737 11363
rect 12771 11329 12805 11363
rect 12839 11329 12873 11363
rect 12907 11329 12941 11363
rect 12975 11329 13009 11363
rect 13043 11329 13077 11363
rect 13111 11329 13145 11363
rect 13179 11329 13213 11363
rect 13247 11329 13281 11363
rect 13315 11329 13349 11363
rect 13383 11329 13417 11363
rect 13451 11329 13485 11363
rect 13519 11329 13553 11363
rect 13587 11329 13621 11363
rect 13655 11329 13689 11363
rect 13723 11329 13757 11363
rect 13791 11329 13825 11363
rect 13859 11329 13893 11363
rect 13927 11329 13961 11363
rect 13995 11329 14029 11363
rect 14063 11329 14097 11363
rect 14131 11329 14165 11363
rect 14199 11329 14233 11363
rect 14267 11329 14301 11363
rect 14335 11329 14369 11363
rect 14403 11329 14437 11363
rect 14471 11329 14505 11363
rect 14539 11329 14573 11363
rect 14607 11329 14641 11363
rect 14675 11329 14709 11363
rect 14743 11329 14777 11363
rect 14811 11329 14845 11363
rect 14879 11329 14913 11363
rect 14947 11329 14981 11363
rect 15015 11329 15049 11363
rect 15083 11329 15117 11363
rect 15151 11329 15185 11363
rect 15219 11329 15253 11363
rect 15287 11329 15321 11363
rect 15355 11329 15389 11363
rect 15423 11329 15457 11363
rect 15491 11329 15525 11363
rect 5583 11227 5617 11261
rect 5651 11230 5685 11264
rect 5719 11236 5753 11270
rect 5806 11257 5840 11291
rect 5875 11257 5909 11291
rect 5944 11257 5978 11291
rect 6013 11257 6047 11291
rect 6082 11257 6116 11291
rect 6151 11257 6185 11291
rect 6220 11257 6254 11291
rect 6289 11257 6323 11291
rect 6358 11257 6392 11291
rect 6427 11257 6461 11291
rect 6496 11257 6530 11291
rect 6565 11257 6599 11291
rect 6634 11257 6668 11291
rect 6703 11257 6737 11291
rect 6772 11257 6806 11291
rect 6841 11257 6875 11291
rect 6910 11257 6944 11291
rect 6979 11257 7013 11291
rect 7048 11257 7082 11291
rect 7117 11257 7151 11291
rect 7186 11257 7220 11291
rect 7255 11257 7289 11291
rect 7324 11257 7358 11291
rect 7393 11257 7427 11291
rect 7462 11257 7496 11291
rect 7531 11257 7565 11291
rect 7600 11257 7634 11291
rect 7669 11257 7703 11291
rect 7738 11257 7772 11291
rect 7807 11257 7841 11291
rect 7875 11257 7909 11291
rect 7943 11257 7977 11291
rect 8011 11257 8045 11291
rect 8079 11257 8113 11291
rect 8147 11257 8181 11291
rect 8215 11257 8249 11291
rect 8283 11257 8317 11291
rect 8351 11257 8385 11291
rect 8419 11257 8453 11291
rect 8487 11257 8521 11291
rect 8555 11257 8589 11291
rect 8623 11257 8657 11291
rect 8691 11257 8725 11291
rect 8759 11257 8793 11291
rect 8827 11257 8861 11291
rect 8895 11257 8929 11291
rect 8963 11257 8997 11291
rect 9031 11257 9065 11291
rect 9099 11257 9133 11291
rect 9167 11257 9201 11291
rect 9235 11257 9269 11291
rect 9303 11257 9337 11291
rect 9371 11257 9405 11291
rect 9439 11257 9473 11291
rect 9507 11257 9541 11291
rect 9575 11257 9609 11291
rect 9643 11257 9677 11291
rect 9711 11257 9745 11291
rect 9779 11257 9813 11291
rect 9847 11257 9881 11291
rect 9915 11257 9949 11291
rect 9983 11257 10017 11291
rect 10051 11257 10085 11291
rect 10119 11257 10153 11291
rect 10187 11257 10221 11291
rect 10255 11257 10289 11291
rect 10323 11257 10357 11291
rect 10391 11257 10425 11291
rect 10459 11257 10493 11291
rect 10527 11257 10561 11291
rect 10595 11257 10629 11291
rect 10663 11257 10697 11291
rect 10731 11257 10765 11291
rect 10799 11257 10833 11291
rect 10867 11257 10901 11291
rect 10935 11257 10969 11291
rect 11003 11257 11037 11291
rect 11071 11257 11105 11291
rect 11139 11257 11173 11291
rect 11207 11257 11241 11291
rect 11275 11257 11309 11291
rect 11343 11257 11377 11291
rect 11411 11257 11445 11291
rect 11479 11257 11513 11291
rect 11547 11257 11581 11291
rect 11615 11257 11649 11291
rect 11683 11257 11717 11291
rect 11751 11257 11785 11291
rect 11819 11257 11853 11291
rect 11887 11257 11921 11291
rect 11955 11257 11989 11291
rect 12023 11257 12057 11291
rect 12091 11257 12125 11291
rect 12159 11257 12193 11291
rect 12227 11257 12261 11291
rect 12295 11257 12329 11291
rect 12363 11257 12397 11291
rect 12431 11257 12465 11291
rect 12499 11257 12533 11291
rect 12567 11257 12601 11291
rect 12635 11257 12669 11291
rect 12703 11257 12737 11291
rect 12771 11257 12805 11291
rect 12839 11257 12873 11291
rect 12907 11257 12941 11291
rect 12975 11257 13009 11291
rect 13043 11257 13077 11291
rect 13111 11257 13145 11291
rect 13179 11257 13213 11291
rect 13247 11257 13281 11291
rect 13315 11257 13349 11291
rect 13383 11257 13417 11291
rect 13451 11257 13485 11291
rect 13519 11257 13553 11291
rect 13587 11257 13621 11291
rect 13655 11257 13689 11291
rect 13723 11257 13757 11291
rect 13791 11257 13825 11291
rect 13859 11257 13893 11291
rect 13927 11257 13961 11291
rect 13995 11257 14029 11291
rect 14063 11257 14097 11291
rect 14131 11257 14165 11291
rect 14199 11257 14233 11291
rect 14267 11257 14301 11291
rect 14335 11257 14369 11291
rect 14403 11257 14437 11291
rect 14471 11257 14505 11291
rect 14539 11257 14573 11291
rect 14607 11257 14641 11291
rect 14675 11257 14709 11291
rect 14743 11257 14777 11291
rect 14811 11257 14845 11291
rect 14879 11257 14913 11291
rect 14947 11257 14981 11291
rect 15015 11257 15049 11291
rect 15083 11257 15117 11291
rect 15151 11257 15185 11291
rect 15219 11257 15253 11291
rect 15287 11257 15321 11291
rect 15355 11257 15389 11291
rect 15423 11257 15457 11291
rect 15491 11257 15525 11291
rect 5583 11157 5617 11191
rect 5651 11160 5685 11194
rect 5719 11166 5753 11200
rect 5806 11185 5840 11219
rect 5875 11185 5909 11219
rect 5944 11185 5978 11219
rect 6013 11185 6047 11219
rect 6082 11185 6116 11219
rect 6151 11185 6185 11219
rect 6220 11185 6254 11219
rect 6289 11185 6323 11219
rect 6358 11185 6392 11219
rect 6427 11185 6461 11219
rect 6496 11185 6530 11219
rect 6565 11185 6599 11219
rect 6634 11185 6668 11219
rect 6703 11185 6737 11219
rect 6772 11185 6806 11219
rect 6841 11185 6875 11219
rect 6910 11185 6944 11219
rect 6979 11185 7013 11219
rect 7048 11185 7082 11219
rect 7117 11185 7151 11219
rect 7186 11185 7220 11219
rect 7255 11185 7289 11219
rect 7324 11185 7358 11219
rect 7393 11185 7427 11219
rect 7462 11185 7496 11219
rect 7531 11185 7565 11219
rect 7600 11185 7634 11219
rect 7669 11185 7703 11219
rect 7738 11185 7772 11219
rect 7807 11185 7841 11219
rect 7875 11185 7909 11219
rect 7943 11185 7977 11219
rect 8011 11185 8045 11219
rect 8079 11185 8113 11219
rect 8147 11185 8181 11219
rect 8215 11185 8249 11219
rect 8283 11185 8317 11219
rect 8351 11185 8385 11219
rect 8419 11185 8453 11219
rect 8487 11185 8521 11219
rect 8555 11185 8589 11219
rect 8623 11185 8657 11219
rect 8691 11185 8725 11219
rect 8759 11185 8793 11219
rect 8827 11185 8861 11219
rect 8895 11185 8929 11219
rect 8963 11185 8997 11219
rect 9031 11185 9065 11219
rect 9099 11185 9133 11219
rect 9167 11185 9201 11219
rect 9235 11185 9269 11219
rect 9303 11185 9337 11219
rect 9371 11185 9405 11219
rect 9439 11185 9473 11219
rect 9507 11185 9541 11219
rect 9575 11185 9609 11219
rect 9643 11185 9677 11219
rect 9711 11185 9745 11219
rect 9779 11185 9813 11219
rect 9847 11185 9881 11219
rect 9915 11185 9949 11219
rect 9983 11185 10017 11219
rect 10051 11185 10085 11219
rect 10119 11185 10153 11219
rect 10187 11185 10221 11219
rect 10255 11185 10289 11219
rect 10323 11185 10357 11219
rect 10391 11185 10425 11219
rect 10459 11185 10493 11219
rect 10527 11185 10561 11219
rect 10595 11185 10629 11219
rect 10663 11185 10697 11219
rect 10731 11185 10765 11219
rect 10799 11185 10833 11219
rect 10867 11185 10901 11219
rect 10935 11185 10969 11219
rect 11003 11185 11037 11219
rect 11071 11185 11105 11219
rect 11139 11185 11173 11219
rect 11207 11185 11241 11219
rect 11275 11185 11309 11219
rect 11343 11185 11377 11219
rect 11411 11185 11445 11219
rect 11479 11185 11513 11219
rect 11547 11185 11581 11219
rect 11615 11185 11649 11219
rect 11683 11185 11717 11219
rect 11751 11185 11785 11219
rect 11819 11185 11853 11219
rect 11887 11185 11921 11219
rect 11955 11185 11989 11219
rect 12023 11185 12057 11219
rect 12091 11185 12125 11219
rect 12159 11185 12193 11219
rect 12227 11185 12261 11219
rect 12295 11185 12329 11219
rect 12363 11185 12397 11219
rect 12431 11185 12465 11219
rect 12499 11185 12533 11219
rect 12567 11185 12601 11219
rect 12635 11185 12669 11219
rect 12703 11185 12737 11219
rect 12771 11185 12805 11219
rect 12839 11185 12873 11219
rect 12907 11185 12941 11219
rect 12975 11185 13009 11219
rect 13043 11185 13077 11219
rect 13111 11185 13145 11219
rect 13179 11185 13213 11219
rect 13247 11185 13281 11219
rect 13315 11185 13349 11219
rect 13383 11185 13417 11219
rect 13451 11185 13485 11219
rect 13519 11185 13553 11219
rect 13587 11185 13621 11219
rect 13655 11185 13689 11219
rect 13723 11185 13757 11219
rect 13791 11185 13825 11219
rect 13859 11185 13893 11219
rect 13927 11185 13961 11219
rect 13995 11185 14029 11219
rect 14063 11185 14097 11219
rect 14131 11185 14165 11219
rect 14199 11185 14233 11219
rect 14267 11185 14301 11219
rect 14335 11185 14369 11219
rect 14403 11185 14437 11219
rect 14471 11185 14505 11219
rect 14539 11185 14573 11219
rect 14607 11185 14641 11219
rect 14675 11185 14709 11219
rect 14743 11185 14777 11219
rect 14811 11185 14845 11219
rect 14879 11185 14913 11219
rect 14947 11185 14981 11219
rect 15015 11185 15049 11219
rect 15083 11185 15117 11219
rect 15151 11185 15185 11219
rect 15219 11185 15253 11219
rect 15287 11185 15321 11219
rect 15355 11185 15389 11219
rect 15423 11185 15457 11219
rect 15491 11185 15525 11219
rect 5583 11087 5617 11121
rect 5651 11090 5685 11124
rect 5719 11096 5753 11130
rect 5583 11017 5617 11051
rect 5651 11020 5685 11054
rect 5719 11026 5753 11060
rect 5583 10947 5617 10981
rect 5651 10950 5685 10984
rect 5719 10956 5753 10990
rect 5583 10877 5617 10911
rect 5651 10880 5685 10914
rect 5719 10886 5753 10920
rect 5583 10807 5617 10841
rect 5651 10810 5685 10844
rect 5719 10816 5753 10850
rect 5583 10737 5617 10771
rect 5651 10740 5685 10774
rect 5719 10746 5753 10780
rect 5583 10667 5617 10701
rect 5651 10670 5685 10704
rect 5719 10676 5753 10710
rect 5583 10597 5617 10631
rect 5651 10600 5685 10634
rect 5719 10606 5753 10640
rect 5719 10568 5753 10570
rect 15578 9754 15748 11760
rect 15714 9749 15748 9754
rect 15578 9685 15612 9719
rect 15646 9685 15680 9719
rect 15714 9681 15748 9715
rect 15578 9616 15612 9650
rect 15646 9616 15680 9650
rect 15714 9613 15748 9647
rect 15578 9547 15612 9581
rect 15646 9547 15680 9581
rect 15714 9545 15748 9579
rect 15578 9478 15612 9512
rect 15646 9478 15680 9512
rect 15714 9477 15748 9511
rect 15578 9409 15612 9443
rect 15646 9409 15680 9443
rect 15714 9409 15748 9443
rect 15578 9340 15612 9374
rect 15646 9340 15680 9374
rect 15714 9340 15748 9374
rect 15578 9271 15612 9305
rect 15646 9271 15680 9305
rect 15714 9271 15748 9305
rect 15578 9202 15612 9236
rect 15646 9202 15680 9236
rect 15714 9202 15748 9236
rect 15578 9133 15612 9167
rect 15646 9133 15680 9167
rect 15714 9133 15748 9167
rect 15578 9064 15612 9098
rect 15646 9064 15680 9098
rect 15714 9064 15748 9098
rect 15578 8995 15612 9029
rect 15646 8995 15680 9029
rect 15714 8995 15748 9029
rect 15578 8926 15612 8960
rect 15646 8926 15680 8960
rect 15714 8926 15748 8960
rect 15578 8857 15612 8891
rect 15646 8857 15680 8891
rect 15714 8857 15748 8891
rect 15578 8788 15612 8822
rect 15646 8788 15680 8822
rect 15714 8788 15748 8822
rect 15578 8719 15612 8753
rect 15646 8719 15680 8753
rect 15714 8719 15748 8753
rect 15578 8650 15612 8684
rect 15646 8650 15680 8684
rect 15714 8650 15748 8684
rect 15578 8581 15612 8615
rect 15646 8581 15680 8615
rect 15714 8581 15748 8615
rect 15578 8512 15612 8546
rect 15646 8512 15680 8546
rect 15714 8512 15748 8546
rect 15578 8443 15612 8477
rect 15646 8443 15680 8477
rect 15714 8443 15748 8477
rect 15578 8374 15612 8408
rect 15646 8374 15680 8408
rect 15714 8374 15748 8408
rect 15578 8305 15612 8339
rect 15646 8305 15680 8339
rect 15714 8305 15748 8339
rect 15578 8236 15612 8270
rect 15646 8236 15680 8270
rect 15714 8236 15748 8270
rect 15578 8167 15612 8201
rect 15646 8167 15680 8201
rect 15714 8167 15748 8201
rect 15578 8098 15612 8132
rect 15646 8098 15680 8132
rect 15714 8098 15748 8132
rect 15578 8029 15612 8063
rect 15646 8029 15680 8063
rect 15714 8029 15748 8063
rect 15578 7960 15612 7994
rect 15646 7960 15680 7994
rect 15714 7960 15748 7994
rect 15578 7891 15612 7925
rect 15646 7891 15680 7925
rect 15714 7891 15748 7925
rect 15578 7822 15612 7856
rect 15646 7822 15680 7856
rect 15714 7822 15748 7856
rect 15578 7753 15612 7787
rect 15646 7753 15680 7787
rect 15714 7753 15748 7787
rect 15578 7684 15612 7718
rect 15646 7684 15680 7718
rect 15714 7684 15748 7718
rect 15578 7615 15612 7649
rect 15646 7615 15680 7649
rect 15714 7615 15748 7649
rect 15578 7546 15612 7580
rect 15646 7546 15680 7580
rect 15714 7546 15748 7580
rect 15578 7477 15612 7511
rect 15646 7477 15680 7511
rect 15714 7477 15748 7511
rect 15578 7408 15612 7442
rect 15646 7408 15680 7442
rect 15714 7408 15748 7442
rect 15578 7339 15612 7373
rect 15646 7339 15680 7373
rect 15714 7339 15748 7373
rect 15578 7270 15612 7304
rect 15646 7270 15680 7304
rect 15714 7270 15748 7304
rect 15578 7201 15612 7235
rect 15646 7201 15680 7235
rect 15714 7201 15748 7235
rect 15578 7132 15612 7166
rect 15646 7132 15680 7166
rect 15714 7132 15748 7166
rect 15578 7063 15612 7097
rect 15646 7063 15680 7097
rect 15714 7063 15748 7097
rect 15578 6994 15612 7028
rect 15646 6994 15680 7028
rect 15714 6994 15748 7028
rect 15578 6925 15612 6959
rect 15646 6925 15680 6959
rect 15714 6925 15748 6959
rect 15578 6856 15612 6890
rect 15646 6856 15680 6890
rect 15714 6856 15748 6890
rect 15578 6787 15612 6821
rect 15646 6787 15680 6821
rect 15714 6787 15748 6821
rect 15578 6718 15612 6752
rect 15646 6718 15680 6752
rect 15714 6718 15748 6752
rect 15578 6649 15612 6683
rect 15646 6649 15680 6683
rect 15714 6649 15748 6683
rect 15578 6580 15612 6614
rect 15646 6580 15680 6614
rect 15714 6580 15748 6614
rect 15578 6511 15612 6545
rect 15646 6511 15680 6545
rect 15714 6511 15748 6545
rect 15578 6442 15612 6476
rect 15646 6442 15680 6476
rect 15714 6442 15748 6476
rect 15578 6373 15612 6407
rect 15646 6373 15680 6407
rect 15714 6373 15748 6407
rect 15578 6304 15612 6338
rect 15646 6304 15680 6338
rect 15714 6304 15748 6338
rect 15578 6235 15612 6269
rect 15646 6235 15680 6269
rect 15714 6235 15748 6269
rect 15578 6166 15612 6200
rect 15646 6166 15680 6200
rect 15714 6166 15748 6200
rect 15578 6097 15612 6131
rect 15646 6097 15680 6131
rect 15714 6097 15748 6131
rect 15578 6028 15612 6062
rect 15646 6028 15680 6062
rect 15714 6028 15748 6062
rect 15578 5959 15612 5993
rect 15646 5959 15680 5993
rect 15714 5959 15748 5993
rect 15578 5890 15612 5924
rect 15646 5890 15680 5924
rect 15714 5890 15748 5924
rect 15578 5821 15612 5855
rect 15646 5821 15680 5855
rect 15714 5821 15748 5855
rect 15578 5752 15612 5786
rect 15646 5752 15680 5786
rect 15714 5752 15748 5786
rect 15578 5683 15612 5717
rect 15646 5683 15680 5717
rect 15714 5683 15748 5717
rect 15578 5614 15612 5648
rect 15646 5614 15680 5648
rect 15714 5614 15748 5648
rect 15578 5545 15612 5579
rect 15646 5545 15680 5579
rect 15714 5545 15748 5579
rect 15578 5476 15612 5510
rect 15646 5476 15680 5510
rect 15714 5476 15748 5510
rect 15578 5407 15612 5441
rect 15646 5407 15680 5441
rect 15714 5407 15748 5441
rect 15578 5338 15612 5372
rect 15646 5338 15680 5372
rect 15714 5338 15748 5372
rect 15578 5269 15612 5303
rect 15646 5269 15680 5303
rect 15714 5269 15748 5303
rect 15578 5200 15612 5234
rect 15646 5200 15680 5234
rect 15714 5200 15748 5234
rect 15578 5131 15612 5165
rect 15646 5131 15680 5165
rect 15714 5131 15748 5165
<< mvpsubdiffcont >>
rect 5583 10527 5617 10561
rect 5651 10530 5685 10564
rect 5719 10536 5753 10568
rect -52 10424 1546 10492
rect 1581 10458 1615 10492
rect 1650 10458 1684 10492
rect 1719 10458 1753 10492
rect 1788 10458 1822 10492
rect 1857 10458 1891 10492
rect 1926 10458 1960 10492
rect 1995 10458 2029 10492
rect 2064 10458 2098 10492
rect 2133 10458 2167 10492
rect 2202 10458 2236 10492
rect 2271 10458 2305 10492
rect 2340 10458 2374 10492
rect 2409 10458 2443 10492
rect 2478 10458 2512 10492
rect 2547 10458 2581 10492
rect 2616 10458 2650 10492
rect 2685 10458 2719 10492
rect 2754 10458 2788 10492
rect 2823 10458 2857 10492
rect 2892 10458 2926 10492
rect 2961 10458 2995 10492
rect 3030 10458 3064 10492
rect 3099 10458 3133 10492
rect 3168 10458 3202 10492
rect 3237 10458 3271 10492
rect 3306 10458 3340 10492
rect 3375 10458 3409 10492
rect 3444 10458 3478 10492
rect 3513 10458 3547 10492
rect 3582 10458 3616 10492
rect 3651 10458 3685 10492
rect 3720 10458 3754 10492
rect 3789 10458 3823 10492
rect 3858 10458 3892 10492
rect 3927 10458 3961 10492
rect 3996 10458 4030 10492
rect 4065 10458 4099 10492
rect 4134 10458 4168 10492
rect 4203 10458 4237 10492
rect 4272 10458 4306 10492
rect 4341 10458 4375 10492
rect 4410 10458 4444 10492
rect 4479 10458 4513 10492
rect 4548 10458 4582 10492
rect 4617 10458 4651 10492
rect 4686 10458 4720 10492
rect 4755 10458 4789 10492
rect 4824 10458 4858 10492
rect 4893 10458 4927 10492
rect 4962 10458 4996 10492
rect 5031 10458 5065 10492
rect 5100 10458 5134 10492
rect 5169 10458 5203 10492
rect 5238 10458 5272 10492
rect 5307 10458 5341 10492
rect 5376 10458 5410 10492
rect 5445 10458 5479 10492
rect 5514 10458 5548 10492
rect 5583 10458 5617 10492
rect 5651 10460 5685 10494
rect 5719 10466 5753 10500
rect -52 10322 1614 10424
rect 1649 10390 1683 10424
rect 1718 10390 1752 10424
rect 1787 10390 1821 10424
rect 1856 10390 1890 10424
rect 1925 10390 1959 10424
rect 1994 10390 2028 10424
rect 2063 10390 2097 10424
rect 2132 10390 2166 10424
rect 2201 10390 2235 10424
rect 2270 10390 2304 10424
rect 2339 10390 2373 10424
rect 2408 10390 2442 10424
rect 2477 10390 2511 10424
rect 2546 10390 2580 10424
rect 2615 10390 2649 10424
rect 2684 10390 2718 10424
rect 2753 10390 2787 10424
rect 2822 10390 2856 10424
rect 2891 10390 2925 10424
rect 2960 10390 2994 10424
rect 3029 10390 3063 10424
rect 3098 10390 3132 10424
rect 3167 10390 3201 10424
rect 3236 10390 3270 10424
rect 3305 10390 3339 10424
rect 3374 10390 3408 10424
rect 3443 10390 3477 10424
rect 3512 10390 3546 10424
rect 3581 10390 3615 10424
rect 3650 10390 3684 10424
rect 3719 10390 3753 10424
rect 3788 10390 3822 10424
rect 3857 10390 3891 10424
rect 3926 10390 3960 10424
rect 3995 10390 4029 10424
rect 4064 10390 4098 10424
rect 4133 10390 4167 10424
rect 4202 10390 4236 10424
rect 4271 10390 4305 10424
rect 4340 10390 4374 10424
rect 4409 10390 4443 10424
rect 4478 10390 4512 10424
rect 4547 10390 4581 10424
rect 4616 10390 4650 10424
rect 4685 10390 4719 10424
rect 4754 10390 4788 10424
rect 4823 10390 4857 10424
rect 4892 10390 4926 10424
rect 4961 10390 4995 10424
rect 5030 10390 5064 10424
rect 5099 10390 5133 10424
rect 5168 10390 5202 10424
rect 5237 10390 5271 10424
rect 5306 10390 5340 10424
rect 5375 10390 5409 10424
rect 5444 10390 5478 10424
rect 5513 10390 5547 10424
rect 5582 10390 5616 10424
rect 5651 10390 5685 10424
rect 5719 10397 5753 10431
rect 1648 10322 1682 10356
rect 1716 10322 1750 10356
rect 1784 10322 1818 10356
rect 1852 10322 1886 10356
rect 1920 10322 1954 10356
rect 1988 10322 2022 10356
rect 2057 10322 2091 10356
rect 2126 10322 2160 10356
rect 2195 10322 2229 10356
rect 2264 10322 2298 10356
rect 2333 10322 2367 10356
rect 2402 10322 2436 10356
rect 2471 10322 2505 10356
rect 2540 10322 2574 10356
rect 2609 10322 2643 10356
rect 2678 10322 2712 10356
rect 2747 10322 2781 10356
rect 2816 10322 2850 10356
rect 2885 10322 2919 10356
rect 2954 10322 2988 10356
rect 3023 10322 3057 10356
rect 3092 10322 3126 10356
rect 3161 10322 3195 10356
rect 3230 10322 3264 10356
rect 3299 10322 3333 10356
rect 3368 10322 3402 10356
rect 3437 10322 3471 10356
rect 3506 10322 3540 10356
rect 3575 10322 3609 10356
rect 3644 10322 3678 10356
rect 3713 10322 3747 10356
rect 3782 10322 3816 10356
rect 3851 10322 3885 10356
rect 3920 10322 3954 10356
rect 3989 10322 4023 10356
rect 4058 10322 4092 10356
rect 4127 10322 4161 10356
rect 4196 10322 4230 10356
rect 4265 10322 4299 10356
rect 4334 10322 4368 10356
rect 4403 10322 4437 10356
rect 4472 10322 4506 10356
rect 4541 10322 4575 10356
rect 4610 10322 4644 10356
rect 4679 10322 4713 10356
rect 4748 10322 4782 10356
rect 4817 10322 4851 10356
rect 4886 10322 4920 10356
rect 4955 10322 4989 10356
rect 5024 10322 5058 10356
rect 5093 10322 5127 10356
rect 5162 10322 5196 10356
rect 5231 10322 5265 10356
rect 5300 10322 5334 10356
rect 5369 10322 5403 10356
rect 5438 10322 5472 10356
rect 5507 10322 5541 10356
rect 5576 10322 5610 10356
rect 5645 10322 5679 10356
rect 5714 10322 5748 10356
<< mvnsubdiffcont >>
rect 12225 10107 12259 10141
rect 12295 10107 12329 10141
rect 12365 10107 12399 10141
rect 12435 10107 12469 10141
rect 12504 10107 12538 10141
rect 12573 10107 12607 10141
rect 12642 10107 12676 10141
rect 12711 10107 12745 10141
rect 12780 10107 12814 10141
rect 12849 10107 12883 10141
rect 12918 10107 12952 10141
rect 12987 10107 13021 10141
rect 13056 10107 13090 10141
rect 13125 10107 13159 10141
rect 13194 10107 13228 10141
rect 13263 10107 13297 10141
rect 13332 10107 13366 10141
rect 13401 10107 13435 10141
rect 13470 10107 13504 10141
rect 13539 10107 13573 10141
rect 13608 10107 13642 10141
rect 13677 10107 13711 10141
rect 13746 10107 13780 10141
rect 13815 10107 13849 10141
rect 13884 10107 13918 10141
rect 13953 10107 13987 10141
rect 14022 10107 14056 10141
rect 14091 10107 14125 10141
rect 14160 10107 14194 10141
rect 14229 10107 14263 10141
rect 14298 10107 14332 10141
rect 14367 10107 14401 10141
rect 14436 10107 14470 10141
rect 14505 10107 14539 10141
rect 14574 10107 14608 10141
rect 14643 10107 14677 10141
rect 14712 10107 14746 10141
rect 14781 10107 14815 10141
rect 14850 10107 14884 10141
rect 14919 10107 14953 10141
rect 14988 10107 15022 10141
rect 15057 10107 15091 10141
rect 15126 10107 15160 10141
rect 15195 10107 15229 10141
rect 15299 10073 15333 10107
rect 15299 10004 15333 10038
rect 15299 9935 15333 9969
rect 15299 9866 15333 9900
rect 15299 9797 15333 9831
rect 15299 9728 15333 9762
rect 15299 9659 15333 9693
rect 15299 9590 15333 9624
rect 15299 9521 15333 9555
rect 15299 9452 15333 9486
rect 15299 9383 15333 9417
rect 15299 9314 15333 9348
rect 15299 9245 15333 9279
rect 15299 9176 15333 9210
rect 15299 9107 15333 9141
rect 15299 9038 15333 9072
rect 15299 8969 15333 9003
rect 15299 8900 15333 8934
rect 15299 8831 15333 8865
rect 15299 8762 15333 8796
rect 15299 8693 15333 8727
rect 15299 8624 15333 8658
rect 15299 8555 15333 8589
rect 15299 8486 15333 8520
rect 15299 8418 15333 8452
rect 15299 8350 15333 8384
rect 15299 8282 15333 8316
rect 15299 8214 15333 8248
rect 15299 8146 15333 8180
rect 15299 8078 15333 8112
rect 15299 8010 15333 8044
rect 15299 7942 15333 7976
rect 15299 7874 15333 7908
rect 14847 7778 14881 7812
rect 14915 7778 14949 7812
rect 15062 7772 15096 7806
rect 15163 7772 15197 7806
rect 15265 7772 15299 7806
rect 14847 7708 14881 7742
rect 14915 7708 14949 7742
rect 14847 7638 14881 7672
rect 14915 7638 14949 7672
rect 14847 7568 14881 7602
rect 14915 7568 14949 7602
rect 14847 7498 14881 7532
rect 14915 7498 14949 7532
rect 14847 7428 14881 7462
rect 14915 7428 14949 7462
rect 14847 7357 14881 7391
rect 14915 7357 14949 7391
rect 14847 7286 14881 7320
rect 14915 7286 14949 7320
rect 14847 7215 14881 7249
rect 14915 7215 14949 7249
rect 14847 7144 14881 7178
rect 14915 7144 14949 7178
rect 14847 7073 14881 7107
rect 14915 7073 14949 7107
rect 14847 7002 14881 7036
rect 14915 7002 14949 7036
rect 14847 6931 14881 6965
rect 14915 6931 14949 6965
rect 14847 6860 14881 6894
rect 14915 6860 14949 6894
rect 14847 6789 14881 6823
rect 14915 6789 14949 6823
rect 14847 6718 14881 6752
rect 14915 6718 14949 6752
rect 14847 6647 14881 6681
rect 14915 6647 14949 6681
rect 14847 6576 14881 6610
rect 14915 6576 14949 6610
rect 14847 6505 14881 6539
rect 14915 6505 14949 6539
rect 14847 6434 14881 6468
rect 14915 6434 14949 6468
rect 14847 6363 14881 6397
rect 14915 6363 14949 6397
rect 14847 6292 14881 6326
rect 14915 6292 14949 6326
<< locali >>
rect 1988 13572 2032 13606
rect 2066 13572 2110 13606
rect 2144 13572 2188 13606
rect 2222 13572 2266 13606
rect 2300 13572 2344 13606
rect 2378 13572 2422 13606
rect 2456 13572 2500 13606
rect 2534 13572 2578 13606
rect 1954 13532 2612 13572
rect 1988 13498 2032 13532
rect 2066 13498 2110 13532
rect 2144 13498 2188 13532
rect 2222 13498 2266 13532
rect 2300 13498 2344 13532
rect 2378 13498 2422 13532
rect 2456 13498 2500 13532
rect 2534 13498 2578 13532
rect 1954 13458 2612 13498
rect 1988 13424 2032 13458
rect 2066 13424 2110 13458
rect 2144 13424 2188 13458
rect 2222 13424 2266 13458
rect 2300 13424 2344 13458
rect 2378 13424 2422 13458
rect 2456 13424 2500 13458
rect 2534 13424 2578 13458
rect 1954 13383 2612 13424
rect 1988 13349 2032 13383
rect 2066 13349 2110 13383
rect 2144 13349 2188 13383
rect 2222 13349 2266 13383
rect 2300 13349 2344 13383
rect 2378 13349 2422 13383
rect 2456 13349 2500 13383
rect 2534 13349 2578 13383
rect 1954 13308 2612 13349
rect 1988 13274 2032 13308
rect 2066 13274 2110 13308
rect 2144 13274 2188 13308
rect 2222 13274 2266 13308
rect 2300 13274 2344 13308
rect 2378 13274 2422 13308
rect 2456 13274 2500 13308
rect 2534 13274 2578 13308
rect 1954 13233 2612 13274
rect 1988 13199 2032 13233
rect 2066 13199 2110 13233
rect 2144 13199 2188 13233
rect 2222 13199 2266 13233
rect 2300 13199 2344 13233
rect 2378 13199 2422 13233
rect 2456 13199 2500 13233
rect 2534 13199 2578 13233
rect 1954 13158 2612 13199
rect 1988 13124 2032 13158
rect 2066 13124 2110 13158
rect 2144 13124 2188 13158
rect 2222 13124 2266 13158
rect 2300 13124 2344 13158
rect 2378 13124 2422 13158
rect 2456 13124 2500 13158
rect 2534 13124 2578 13158
rect 1954 13083 2612 13124
rect 1988 13049 2032 13083
rect 2066 13049 2110 13083
rect 2144 13049 2188 13083
rect 2222 13049 2266 13083
rect 2300 13049 2344 13083
rect 2378 13049 2422 13083
rect 2456 13049 2500 13083
rect 2534 13049 2578 13083
rect 1954 13008 2612 13049
rect 1988 12974 2032 13008
rect 2066 12974 2110 13008
rect 2144 12974 2188 13008
rect 2222 12974 2266 13008
rect 2300 12974 2344 13008
rect 2378 12974 2422 13008
rect 2456 12974 2500 13008
rect 2534 12974 2578 13008
rect 1954 12933 2612 12974
rect 1988 12899 2032 12933
rect 2066 12899 2110 12933
rect 2144 12899 2188 12933
rect 2222 12899 2266 12933
rect 2300 12899 2344 12933
rect 2378 12899 2422 12933
rect 2456 12899 2500 12933
rect 2534 12899 2578 12933
rect 1934 12364 4257 12367
rect 1968 12330 2008 12364
rect 2042 12330 2082 12364
rect 2116 12330 2156 12364
rect 2190 12330 2230 12364
rect 2264 12330 2304 12364
rect 2338 12330 2378 12364
rect 2412 12330 2452 12364
rect 2486 12330 2526 12364
rect 2560 12330 2600 12364
rect 2634 12330 2674 12364
rect 2708 12330 2748 12364
rect 2782 12330 2822 12364
rect 2856 12330 2896 12364
rect 2930 12330 2970 12364
rect 3004 12330 3044 12364
rect 3078 12330 3118 12364
rect 3152 12330 3192 12364
rect 3226 12330 3266 12364
rect 3300 12330 3340 12364
rect 3374 12330 3414 12364
rect 3448 12330 3488 12364
rect 3522 12330 3562 12364
rect 3596 12330 3636 12364
rect 3670 12330 3710 12364
rect 3744 12330 3784 12364
rect 3818 12330 3858 12364
rect 3892 12330 3931 12364
rect 3965 12330 4004 12364
rect 4038 12330 4077 12364
rect 4111 12330 4150 12364
rect 4184 12330 4223 12364
rect 1934 12282 4257 12330
rect 1968 12248 2008 12282
rect 2042 12248 2082 12282
rect 2116 12248 2156 12282
rect 2190 12248 2230 12282
rect 2264 12248 2304 12282
rect 2338 12248 2378 12282
rect 2412 12248 2452 12282
rect 2486 12248 2526 12282
rect 2560 12248 2600 12282
rect 2634 12248 2674 12282
rect 2708 12248 2748 12282
rect 2782 12248 2822 12282
rect 2856 12248 2896 12282
rect 2930 12248 2970 12282
rect 3004 12248 3044 12282
rect 3078 12248 3118 12282
rect 3152 12248 3192 12282
rect 3226 12248 3266 12282
rect 3300 12248 3340 12282
rect 3374 12248 3414 12282
rect 3448 12248 3488 12282
rect 3522 12248 3562 12282
rect 3596 12248 3636 12282
rect 3670 12248 3710 12282
rect 3744 12248 3784 12282
rect 3818 12248 3858 12282
rect 3892 12248 3931 12282
rect 3965 12248 4004 12282
rect 4038 12248 4077 12282
rect 4111 12248 4150 12282
rect 4184 12248 4223 12282
rect -2911 12237 307 12242
rect -2877 12203 -2838 12237
rect -2804 12203 -2765 12237
rect -2731 12203 -2692 12237
rect -2658 12203 -2619 12237
rect -2585 12203 -2546 12237
rect -2512 12203 -2473 12237
rect -2439 12203 -2400 12237
rect -2366 12203 -2327 12237
rect -2293 12203 -2254 12237
rect -2220 12203 -2181 12237
rect -2147 12203 -2108 12237
rect -2074 12203 -2035 12237
rect -2001 12203 -1962 12237
rect -1928 12203 -1889 12237
rect -1855 12203 -1816 12237
rect -1782 12203 -1743 12237
rect -2911 12165 -1743 12203
rect -2877 12131 -2838 12165
rect -2804 12131 -2765 12165
rect -2731 12131 -2692 12165
rect -2658 12131 -2619 12165
rect -2585 12131 -2546 12165
rect -2512 12131 -2473 12165
rect -2439 12131 -2400 12165
rect -2366 12131 -2327 12165
rect -2293 12131 -2254 12165
rect -2220 12131 -2181 12165
rect -2147 12131 -2108 12165
rect -2074 12131 -2035 12165
rect -2001 12131 -1962 12165
rect -1928 12131 -1889 12165
rect -1855 12131 -1816 12165
rect -1782 12131 -1743 12165
rect -2911 12093 -1743 12131
rect -2877 12059 -2838 12093
rect -2804 12059 -2765 12093
rect -2731 12059 -2692 12093
rect -2658 12059 -2619 12093
rect -2585 12059 -2546 12093
rect -2512 12059 -2473 12093
rect -2439 12059 -2400 12093
rect -2366 12059 -2327 12093
rect -2293 12059 -2254 12093
rect -2220 12059 -2181 12093
rect -2147 12059 -2108 12093
rect -2074 12059 -2035 12093
rect -2001 12059 -1962 12093
rect -1928 12059 -1889 12093
rect -1855 12059 -1816 12093
rect -1782 12059 -1743 12093
rect -2911 12021 -1743 12059
rect -2877 11987 -2838 12021
rect -2804 11987 -2765 12021
rect -2731 11987 -2692 12021
rect -2658 11987 -2619 12021
rect -2585 11987 -2546 12021
rect -2512 11987 -2473 12021
rect -2439 11987 -2400 12021
rect -2366 11987 -2327 12021
rect -2293 11987 -2254 12021
rect -2220 11987 -2181 12021
rect -2147 11987 -2108 12021
rect -2074 11987 -2035 12021
rect -2001 11987 -1962 12021
rect -1928 11987 -1889 12021
rect -1855 11987 -1816 12021
rect -1782 11987 -1743 12021
rect -2911 11949 -1743 11987
rect -2877 11915 -2838 11949
rect -2804 11915 -2765 11949
rect -2731 11915 -2692 11949
rect -2658 11915 -2619 11949
rect -2585 11915 -2546 11949
rect -2512 11915 -2473 11949
rect -2439 11915 -2400 11949
rect -2366 11915 -2327 11949
rect -2293 11915 -2254 11949
rect -2220 11915 -2181 11949
rect -2147 11915 -2108 11949
rect -2074 11915 -2035 11949
rect -2001 11915 -1962 11949
rect -1928 11915 -1889 11949
rect -1855 11915 -1816 11949
rect -1782 11915 -1743 11949
rect -2911 11877 -1743 11915
rect -2877 11843 -2838 11877
rect -2804 11843 -2765 11877
rect -2731 11843 -2692 11877
rect -2658 11843 -2619 11877
rect -2585 11843 -2546 11877
rect -2512 11843 -2473 11877
rect -2439 11843 -2400 11877
rect -2366 11843 -2327 11877
rect -2293 11843 -2254 11877
rect -2220 11843 -2181 11877
rect -2147 11843 -2108 11877
rect -2074 11843 -2035 11877
rect -2001 11843 -1962 11877
rect -1928 11843 -1889 11877
rect -1855 11843 -1816 11877
rect -1782 11843 -1743 11877
rect -2911 11805 -1743 11843
rect -2877 11771 -2838 11805
rect -2804 11771 -2765 11805
rect -2731 11771 -2692 11805
rect -2658 11771 -2619 11805
rect -2585 11771 -2546 11805
rect -2512 11771 -2473 11805
rect -2439 11771 -2400 11805
rect -2366 11771 -2327 11805
rect -2293 11771 -2254 11805
rect -2220 11771 -2181 11805
rect -2147 11771 -2108 11805
rect -2074 11771 -2035 11805
rect -2001 11771 -1962 11805
rect -1928 11771 -1889 11805
rect -1855 11771 -1816 11805
rect -1782 11771 -1743 11805
rect 1934 12200 4257 12248
rect 1968 12166 2008 12200
rect 2042 12166 2082 12200
rect 2116 12166 2156 12200
rect 2190 12166 2230 12200
rect 2264 12166 2304 12200
rect 2338 12166 2378 12200
rect 2412 12166 2452 12200
rect 2486 12166 2526 12200
rect 2560 12166 2600 12200
rect 2634 12166 2674 12200
rect 2708 12166 2748 12200
rect 2782 12166 2822 12200
rect 2856 12166 2896 12200
rect 2930 12166 2970 12200
rect 3004 12166 3044 12200
rect 3078 12166 3118 12200
rect 3152 12166 3192 12200
rect 3226 12166 3266 12200
rect 3300 12166 3340 12200
rect 3374 12166 3414 12200
rect 3448 12166 3488 12200
rect 3522 12166 3562 12200
rect 3596 12166 3636 12200
rect 3670 12166 3710 12200
rect 3744 12166 3784 12200
rect 3818 12166 3858 12200
rect 3892 12166 3931 12200
rect 3965 12166 4004 12200
rect 4038 12166 4077 12200
rect 4111 12166 4150 12200
rect 4184 12166 4223 12200
rect 1934 12118 4257 12166
rect 1968 12084 2008 12118
rect 2042 12084 2082 12118
rect 2116 12084 2156 12118
rect 2190 12084 2230 12118
rect 2264 12084 2304 12118
rect 2338 12084 2378 12118
rect 2412 12084 2452 12118
rect 2486 12084 2526 12118
rect 2560 12084 2600 12118
rect 2634 12084 2674 12118
rect 2708 12084 2748 12118
rect 2782 12084 2822 12118
rect 2856 12084 2896 12118
rect 2930 12084 2970 12118
rect 3004 12084 3044 12118
rect 3078 12084 3118 12118
rect 3152 12084 3192 12118
rect 3226 12084 3266 12118
rect 3300 12084 3340 12118
rect 3374 12084 3414 12118
rect 3448 12084 3488 12118
rect 3522 12084 3562 12118
rect 3596 12084 3636 12118
rect 3670 12084 3710 12118
rect 3744 12084 3784 12118
rect 3818 12084 3858 12118
rect 3892 12084 3931 12118
rect 3965 12084 4004 12118
rect 4038 12084 4077 12118
rect 4111 12084 4150 12118
rect 4184 12084 4223 12118
rect 1934 12036 4257 12084
rect 1968 12002 2008 12036
rect 2042 12002 2082 12036
rect 2116 12002 2156 12036
rect 2190 12002 2230 12036
rect 2264 12002 2304 12036
rect 2338 12002 2378 12036
rect 2412 12002 2452 12036
rect 2486 12002 2526 12036
rect 2560 12002 2600 12036
rect 2634 12002 2674 12036
rect 2708 12002 2748 12036
rect 2782 12002 2822 12036
rect 2856 12002 2896 12036
rect 2930 12002 2970 12036
rect 3004 12002 3044 12036
rect 3078 12002 3118 12036
rect 3152 12002 3192 12036
rect 3226 12002 3266 12036
rect 3300 12002 3340 12036
rect 3374 12002 3414 12036
rect 3448 12002 3488 12036
rect 3522 12002 3562 12036
rect 3596 12002 3636 12036
rect 3670 12002 3710 12036
rect 3744 12002 3784 12036
rect 3818 12002 3858 12036
rect 3892 12002 3931 12036
rect 3965 12002 4004 12036
rect 4038 12002 4077 12036
rect 4111 12002 4150 12036
rect 4184 12002 4223 12036
rect 1934 11999 4257 12002
rect -2911 11766 307 11771
rect 401 11942 441 11976
rect 475 11942 515 11976
rect 549 11942 588 11976
rect 622 11942 661 11976
rect 695 11942 734 11976
rect 768 11942 807 11976
rect 841 11942 880 11976
rect 914 11942 953 11976
rect 987 11942 1026 11976
rect 1060 11942 1099 11976
rect 1133 11942 1172 11976
rect 1206 11942 1245 11976
rect 1279 11942 1318 11976
rect 1352 11942 1391 11976
rect 1425 11942 1464 11976
rect 1498 11942 1537 11976
rect 1571 11942 1610 11976
rect 1644 11942 1683 11976
rect 367 11888 1717 11942
rect 401 11854 441 11888
rect 475 11854 515 11888
rect 549 11854 588 11888
rect 622 11854 661 11888
rect 695 11854 734 11888
rect 768 11854 807 11888
rect 841 11854 880 11888
rect 914 11854 953 11888
rect 987 11854 1026 11888
rect 1060 11854 1099 11888
rect 1133 11854 1172 11888
rect 1206 11854 1245 11888
rect 1279 11854 1318 11888
rect 1352 11854 1391 11888
rect 1425 11854 1464 11888
rect 1498 11854 1537 11888
rect 1571 11854 1610 11888
rect 1644 11854 1683 11888
rect 367 11800 1717 11854
rect 401 11766 441 11800
rect 475 11766 515 11800
rect 549 11766 588 11800
rect 622 11766 661 11800
rect 695 11766 734 11800
rect 768 11766 807 11800
rect 841 11766 880 11800
rect 914 11766 953 11800
rect 987 11766 1026 11800
rect 1060 11766 1099 11800
rect 1133 11766 1172 11800
rect 1206 11766 1245 11800
rect 1279 11766 1318 11800
rect 1352 11766 1391 11800
rect 1425 11766 1464 11800
rect 1498 11766 1537 11800
rect 1571 11766 1610 11800
rect 1644 11766 1683 11800
rect 5554 11896 15777 11925
rect 5554 11891 5656 11896
rect 5554 11857 5583 11891
rect 5617 11857 5656 11891
rect 11062 11862 11096 11896
rect 11130 11862 11164 11896
rect 11198 11862 11232 11896
rect 11266 11862 11300 11896
rect 11334 11862 11368 11896
rect 11402 11862 11436 11896
rect 11470 11862 11504 11896
rect 11538 11862 11572 11896
rect 11606 11862 11640 11896
rect 11674 11862 11708 11896
rect 11742 11862 11776 11896
rect 11810 11862 11845 11896
rect 11879 11862 11914 11896
rect 11948 11862 11983 11896
rect 12017 11862 12052 11896
rect 12086 11862 12121 11896
rect 12155 11862 12190 11896
rect 12224 11862 12259 11896
rect 12293 11862 12328 11896
rect 12362 11862 12397 11896
rect 12431 11862 12466 11896
rect 12500 11862 12535 11896
rect 12569 11862 12604 11896
rect 12638 11862 12673 11896
rect 12707 11862 12742 11896
rect 12776 11862 12811 11896
rect 12845 11862 12880 11896
rect 12914 11862 12949 11896
rect 12983 11862 13018 11896
rect 13052 11862 13087 11896
rect 13121 11862 13156 11896
rect 13190 11862 13225 11896
rect 13259 11862 13294 11896
rect 13328 11862 13363 11896
rect 13397 11862 13432 11896
rect 13466 11862 13501 11896
rect 13535 11862 13570 11896
rect 13604 11862 13639 11896
rect 13673 11862 13708 11896
rect 13742 11862 13777 11896
rect 13811 11862 13846 11896
rect 13880 11862 13915 11896
rect 13949 11862 13984 11896
rect 14018 11862 14053 11896
rect 14087 11862 14122 11896
rect 14156 11862 14191 11896
rect 14225 11862 14260 11896
rect 14294 11862 14329 11896
rect 14363 11862 14398 11896
rect 14432 11862 14467 11896
rect 14501 11862 14536 11896
rect 14570 11862 14605 11896
rect 14639 11862 14674 11896
rect 14708 11862 14743 11896
rect 14777 11862 14812 11896
rect 14846 11862 14881 11896
rect 14915 11862 14950 11896
rect 14984 11862 15019 11896
rect 15053 11862 15088 11896
rect 15122 11862 15157 11896
rect 15191 11862 15226 11896
rect 15260 11862 15295 11896
rect 15329 11862 15364 11896
rect 15398 11862 15433 11896
rect 15467 11862 15502 11896
rect 15536 11862 15571 11896
rect 15605 11862 15640 11896
rect 15674 11862 15709 11896
rect 15743 11862 15777 11896
rect 5554 11828 5656 11857
rect 11057 11828 15777 11862
rect 5554 11821 5651 11828
rect 5554 11787 5583 11821
rect 5617 11794 5651 11821
rect 11057 11794 11092 11828
rect 11126 11794 11161 11828
rect 11195 11794 11230 11828
rect 11264 11794 11299 11828
rect 11333 11794 11368 11828
rect 11402 11794 11437 11828
rect 11471 11794 11506 11828
rect 11540 11794 11575 11828
rect 11609 11794 11644 11828
rect 11678 11794 11713 11828
rect 11747 11794 11782 11828
rect 11816 11794 11851 11828
rect 11885 11794 11920 11828
rect 11954 11794 11989 11828
rect 12023 11794 12058 11828
rect 12092 11794 12127 11828
rect 12161 11794 12196 11828
rect 12230 11794 12265 11828
rect 12299 11794 12334 11828
rect 12368 11794 12403 11828
rect 12437 11794 12472 11828
rect 12506 11794 12541 11828
rect 12575 11794 12610 11828
rect 12644 11794 12679 11828
rect 12713 11794 12748 11828
rect 12782 11794 12817 11828
rect 12851 11794 12886 11828
rect 12920 11794 12955 11828
rect 12989 11794 13024 11828
rect 13058 11794 13093 11828
rect 13127 11794 13162 11828
rect 13196 11794 13231 11828
rect 13265 11794 13300 11828
rect 13334 11794 13369 11828
rect 13403 11794 13438 11828
rect 13472 11794 13507 11828
rect 13541 11794 13576 11828
rect 13610 11794 13645 11828
rect 13679 11794 13714 11828
rect 13748 11794 13783 11828
rect 13817 11794 13852 11828
rect 13886 11794 13921 11828
rect 13955 11794 13990 11828
rect 14024 11794 14059 11828
rect 14093 11794 14128 11828
rect 14162 11794 14197 11828
rect 14231 11794 14266 11828
rect 14300 11794 14335 11828
rect 14369 11794 14404 11828
rect 14438 11794 14473 11828
rect 14507 11794 14542 11828
rect 14576 11794 14611 11828
rect 14645 11794 14680 11828
rect 14714 11794 14749 11828
rect 14783 11794 14818 11828
rect 14852 11794 14887 11828
rect 14921 11794 14956 11828
rect 14990 11794 15025 11828
rect 15059 11794 15094 11828
rect 15128 11794 15163 11828
rect 15197 11794 15232 11828
rect 15266 11794 15301 11828
rect 15335 11794 15370 11828
rect 15404 11794 15439 11828
rect 15473 11794 15508 11828
rect 15542 11794 15577 11828
rect 15611 11794 15646 11828
rect 15680 11823 15777 11828
rect 5617 11787 5719 11794
rect 5554 11757 5719 11787
rect 5554 11751 5651 11757
rect 5554 11717 5583 11751
rect 5617 11723 5651 11751
rect 5685 11726 5719 11757
rect 10989 11760 15646 11794
rect 10989 11726 11024 11760
rect 11058 11726 11093 11760
rect 11127 11726 11162 11760
rect 11196 11726 11231 11760
rect 11265 11726 11300 11760
rect 11334 11726 11369 11760
rect 11403 11726 11438 11760
rect 11472 11726 11507 11760
rect 11541 11726 11576 11760
rect 11610 11726 11645 11760
rect 11679 11726 11714 11760
rect 11748 11726 11783 11760
rect 11817 11726 11852 11760
rect 11886 11726 11921 11760
rect 11955 11726 11990 11760
rect 12024 11726 12059 11760
rect 12093 11726 12128 11760
rect 12162 11726 12197 11760
rect 12231 11726 12266 11760
rect 12300 11726 12335 11760
rect 12369 11726 12404 11760
rect 12438 11726 12473 11760
rect 12507 11726 12542 11760
rect 12576 11726 12611 11760
rect 12645 11726 12680 11760
rect 12714 11726 12749 11760
rect 12783 11726 12818 11760
rect 12852 11726 12887 11760
rect 12921 11726 12956 11760
rect 12990 11726 13025 11760
rect 13059 11726 13094 11760
rect 13128 11726 13163 11760
rect 13197 11726 13232 11760
rect 13266 11726 13301 11760
rect 13335 11726 13370 11760
rect 13404 11726 13439 11760
rect 13473 11726 13508 11760
rect 13542 11726 13577 11760
rect 13611 11726 13646 11760
rect 13680 11726 13715 11760
rect 13749 11726 13784 11760
rect 13818 11726 13853 11760
rect 13887 11726 13922 11760
rect 13956 11726 13991 11760
rect 14025 11726 14060 11760
rect 14094 11726 14129 11760
rect 14163 11726 14198 11760
rect 14232 11726 14267 11760
rect 14301 11726 14336 11760
rect 14370 11726 14405 11760
rect 14439 11726 14474 11760
rect 14508 11726 14543 11760
rect 14577 11726 14612 11760
rect 14646 11726 14681 11760
rect 14715 11726 14750 11760
rect 14784 11726 14819 11760
rect 14853 11726 14888 11760
rect 14922 11726 14957 11760
rect 14991 11726 15026 11760
rect 15060 11726 15095 11760
rect 15129 11726 15164 11760
rect 15198 11726 15233 11760
rect 15267 11726 15302 11760
rect 15336 11726 15371 11760
rect 15405 11726 15440 11760
rect 15474 11726 15509 11760
rect 15543 11726 15578 11760
rect 5685 11723 15578 11726
rect 5617 11717 15578 11723
rect 5554 11690 15578 11717
rect 5554 11686 5719 11690
rect 5554 11681 5651 11686
rect 5554 11647 5583 11681
rect 5617 11652 5651 11681
rect 5685 11656 5719 11686
rect 5753 11656 15578 11690
rect 5685 11652 15578 11656
rect 5617 11651 15578 11652
rect 5617 11647 5806 11651
rect 5554 11620 5806 11647
rect 5554 11615 5719 11620
rect 5554 11611 5651 11615
rect 5554 11577 5583 11611
rect 5617 11581 5651 11611
rect 5685 11586 5719 11615
rect 5753 11617 5806 11620
rect 5840 11617 5875 11651
rect 5909 11617 5944 11651
rect 5978 11617 6013 11651
rect 6047 11617 6082 11651
rect 6116 11617 6151 11651
rect 6185 11617 6220 11651
rect 6254 11617 6289 11651
rect 6323 11617 6358 11651
rect 6392 11617 6427 11651
rect 6461 11617 6496 11651
rect 6530 11617 6565 11651
rect 6599 11617 6634 11651
rect 6668 11617 6703 11651
rect 6737 11617 6772 11651
rect 6806 11617 6841 11651
rect 6875 11617 6910 11651
rect 6944 11617 6979 11651
rect 7013 11617 7048 11651
rect 7082 11617 7117 11651
rect 7151 11617 7186 11651
rect 7220 11617 7255 11651
rect 7289 11617 7324 11651
rect 7358 11617 7393 11651
rect 7427 11617 7462 11651
rect 7496 11617 7531 11651
rect 7565 11617 7600 11651
rect 7634 11617 7669 11651
rect 7703 11617 7738 11651
rect 7772 11617 7807 11651
rect 7841 11617 7875 11651
rect 7909 11617 7943 11651
rect 7977 11617 8011 11651
rect 8045 11617 8079 11651
rect 8113 11617 8147 11651
rect 8181 11617 8215 11651
rect 8249 11617 8283 11651
rect 8317 11617 8351 11651
rect 8385 11617 8419 11651
rect 8453 11617 8487 11651
rect 8521 11617 8555 11651
rect 8589 11617 8623 11651
rect 8657 11617 8691 11651
rect 8725 11617 8759 11651
rect 8793 11617 8827 11651
rect 8861 11617 8895 11651
rect 8929 11617 8963 11651
rect 8997 11617 9031 11651
rect 9065 11617 9099 11651
rect 9133 11617 9167 11651
rect 9201 11617 9235 11651
rect 9269 11617 9303 11651
rect 9337 11617 9371 11651
rect 9405 11617 9439 11651
rect 9473 11617 9507 11651
rect 9541 11617 9575 11651
rect 9609 11617 9643 11651
rect 9677 11617 9711 11651
rect 9745 11617 9779 11651
rect 9813 11617 9847 11651
rect 9881 11617 9915 11651
rect 9949 11617 9983 11651
rect 10017 11617 10051 11651
rect 10085 11617 10119 11651
rect 10153 11617 10187 11651
rect 10221 11617 10255 11651
rect 10289 11617 10323 11651
rect 10357 11617 10391 11651
rect 10425 11617 10459 11651
rect 10493 11617 10527 11651
rect 10561 11617 10595 11651
rect 10629 11617 10663 11651
rect 10697 11617 10731 11651
rect 10765 11617 10799 11651
rect 10833 11617 10867 11651
rect 10901 11617 10935 11651
rect 10969 11617 11003 11651
rect 11037 11617 11071 11651
rect 11105 11617 11139 11651
rect 11173 11617 11207 11651
rect 11241 11617 11275 11651
rect 11309 11617 11343 11651
rect 11377 11617 11411 11651
rect 11445 11617 11479 11651
rect 11513 11617 11547 11651
rect 11581 11617 11615 11651
rect 11649 11617 11683 11651
rect 11717 11617 11751 11651
rect 11785 11617 11819 11651
rect 11853 11617 11887 11651
rect 11921 11617 11955 11651
rect 11989 11617 12023 11651
rect 12057 11617 12091 11651
rect 12125 11617 12159 11651
rect 12193 11617 12227 11651
rect 12261 11617 12295 11651
rect 12329 11617 12363 11651
rect 12397 11617 12431 11651
rect 12465 11617 12499 11651
rect 12533 11617 12567 11651
rect 12601 11617 12635 11651
rect 12669 11617 12703 11651
rect 12737 11617 12771 11651
rect 12805 11617 12839 11651
rect 12873 11617 12907 11651
rect 12941 11617 12975 11651
rect 13009 11617 13043 11651
rect 13077 11617 13111 11651
rect 13145 11617 13179 11651
rect 13213 11617 13247 11651
rect 13281 11617 13315 11651
rect 13349 11617 13383 11651
rect 13417 11617 13451 11651
rect 13485 11617 13519 11651
rect 13553 11617 13587 11651
rect 13621 11617 13655 11651
rect 13689 11617 13723 11651
rect 13757 11617 13791 11651
rect 13825 11617 13859 11651
rect 13893 11617 13927 11651
rect 13961 11617 13995 11651
rect 14029 11617 14063 11651
rect 14097 11617 14131 11651
rect 14165 11617 14199 11651
rect 14233 11617 14267 11651
rect 14301 11617 14335 11651
rect 14369 11617 14403 11651
rect 14437 11617 14471 11651
rect 14505 11617 14539 11651
rect 14573 11617 14607 11651
rect 14641 11617 14675 11651
rect 14709 11617 14743 11651
rect 14777 11617 14811 11651
rect 14845 11617 14879 11651
rect 14913 11617 14947 11651
rect 14981 11617 15015 11651
rect 15049 11617 15083 11651
rect 15117 11617 15151 11651
rect 15185 11617 15219 11651
rect 15253 11617 15287 11651
rect 15321 11617 15355 11651
rect 15389 11617 15423 11651
rect 15457 11617 15491 11651
rect 15525 11617 15578 11651
rect 5753 11586 15578 11617
rect 5685 11581 15578 11586
rect 5617 11579 15578 11581
rect 5617 11577 5806 11579
rect 5554 11550 5806 11577
rect 5554 11544 5719 11550
rect 5554 11541 5651 11544
rect 5554 11507 5583 11541
rect 5617 11510 5651 11541
rect 5685 11516 5719 11544
rect 5753 11545 5806 11550
rect 5840 11545 5875 11579
rect 5909 11545 5944 11579
rect 5978 11545 6013 11579
rect 6047 11545 6082 11579
rect 6116 11545 6151 11579
rect 6185 11545 6220 11579
rect 6254 11545 6289 11579
rect 6323 11545 6358 11579
rect 6392 11545 6427 11579
rect 6461 11545 6496 11579
rect 6530 11545 6565 11579
rect 6599 11545 6634 11579
rect 6668 11545 6703 11579
rect 6737 11545 6772 11579
rect 6806 11545 6841 11579
rect 6875 11545 6910 11579
rect 6944 11545 6979 11579
rect 7013 11545 7048 11579
rect 7082 11545 7117 11579
rect 7151 11545 7186 11579
rect 7220 11545 7255 11579
rect 7289 11545 7324 11579
rect 7358 11545 7393 11579
rect 7427 11545 7462 11579
rect 7496 11545 7531 11579
rect 7565 11545 7600 11579
rect 7634 11545 7669 11579
rect 7703 11545 7738 11579
rect 7772 11545 7807 11579
rect 7841 11545 7875 11579
rect 7909 11545 7943 11579
rect 7977 11545 8011 11579
rect 8045 11545 8079 11579
rect 8113 11545 8147 11579
rect 8181 11545 8215 11579
rect 8249 11545 8283 11579
rect 8317 11545 8351 11579
rect 8385 11545 8419 11579
rect 8453 11545 8487 11579
rect 8521 11545 8555 11579
rect 8589 11545 8623 11579
rect 8657 11545 8691 11579
rect 8725 11545 8759 11579
rect 8793 11545 8827 11579
rect 8861 11545 8895 11579
rect 8929 11545 8963 11579
rect 8997 11545 9031 11579
rect 9065 11545 9099 11579
rect 9133 11545 9167 11579
rect 9201 11545 9235 11579
rect 9269 11545 9303 11579
rect 9337 11545 9371 11579
rect 9405 11545 9439 11579
rect 9473 11545 9507 11579
rect 9541 11545 9575 11579
rect 9609 11545 9643 11579
rect 9677 11545 9711 11579
rect 9745 11545 9779 11579
rect 9813 11545 9847 11579
rect 9881 11545 9915 11579
rect 9949 11545 9983 11579
rect 10017 11545 10051 11579
rect 10085 11545 10119 11579
rect 10153 11545 10187 11579
rect 10221 11545 10255 11579
rect 10289 11545 10323 11579
rect 10357 11545 10391 11579
rect 10425 11545 10459 11579
rect 10493 11545 10527 11579
rect 10561 11545 10595 11579
rect 10629 11545 10663 11579
rect 10697 11545 10731 11579
rect 10765 11545 10799 11579
rect 10833 11545 10867 11579
rect 10901 11545 10935 11579
rect 10969 11545 11003 11579
rect 11037 11545 11071 11579
rect 11105 11545 11139 11579
rect 11173 11545 11207 11579
rect 11241 11545 11275 11579
rect 11309 11545 11343 11579
rect 11377 11545 11411 11579
rect 11445 11545 11479 11579
rect 11513 11545 11547 11579
rect 11581 11545 11615 11579
rect 11649 11545 11683 11579
rect 11717 11545 11751 11579
rect 11785 11545 11819 11579
rect 11853 11545 11887 11579
rect 11921 11545 11955 11579
rect 11989 11545 12023 11579
rect 12057 11545 12091 11579
rect 12125 11545 12159 11579
rect 12193 11545 12227 11579
rect 12261 11545 12295 11579
rect 12329 11545 12363 11579
rect 12397 11545 12431 11579
rect 12465 11545 12499 11579
rect 12533 11545 12567 11579
rect 12601 11545 12635 11579
rect 12669 11545 12703 11579
rect 12737 11545 12771 11579
rect 12805 11545 12839 11579
rect 12873 11545 12907 11579
rect 12941 11545 12975 11579
rect 13009 11545 13043 11579
rect 13077 11545 13111 11579
rect 13145 11545 13179 11579
rect 13213 11545 13247 11579
rect 13281 11545 13315 11579
rect 13349 11545 13383 11579
rect 13417 11545 13451 11579
rect 13485 11545 13519 11579
rect 13553 11545 13587 11579
rect 13621 11545 13655 11579
rect 13689 11545 13723 11579
rect 13757 11545 13791 11579
rect 13825 11545 13859 11579
rect 13893 11545 13927 11579
rect 13961 11545 13995 11579
rect 14029 11545 14063 11579
rect 14097 11545 14131 11579
rect 14165 11545 14199 11579
rect 14233 11545 14267 11579
rect 14301 11545 14335 11579
rect 14369 11545 14403 11579
rect 14437 11545 14471 11579
rect 14505 11545 14539 11579
rect 14573 11545 14607 11579
rect 14641 11545 14675 11579
rect 14709 11545 14743 11579
rect 14777 11545 14811 11579
rect 14845 11545 14879 11579
rect 14913 11545 14947 11579
rect 14981 11545 15015 11579
rect 15049 11545 15083 11579
rect 15117 11545 15151 11579
rect 15185 11545 15219 11579
rect 15253 11545 15287 11579
rect 15321 11545 15355 11579
rect 15389 11545 15423 11579
rect 15457 11545 15491 11579
rect 15525 11545 15578 11579
rect 5753 11516 15578 11545
rect 5685 11510 15578 11516
rect 5617 11507 15578 11510
rect 5554 11480 5806 11507
rect 5554 11474 5719 11480
rect 5554 11471 5651 11474
rect 5554 11437 5583 11471
rect 5617 11440 5651 11471
rect 5685 11446 5719 11474
rect 5753 11473 5806 11480
rect 5840 11473 5875 11507
rect 5909 11473 5944 11507
rect 5978 11473 6013 11507
rect 6047 11473 6082 11507
rect 6116 11473 6151 11507
rect 6185 11473 6220 11507
rect 6254 11473 6289 11507
rect 6323 11473 6358 11507
rect 6392 11473 6427 11507
rect 6461 11473 6496 11507
rect 6530 11473 6565 11507
rect 6599 11473 6634 11507
rect 6668 11473 6703 11507
rect 6737 11473 6772 11507
rect 6806 11473 6841 11507
rect 6875 11473 6910 11507
rect 6944 11473 6979 11507
rect 7013 11473 7048 11507
rect 7082 11473 7117 11507
rect 7151 11473 7186 11507
rect 7220 11473 7255 11507
rect 7289 11473 7324 11507
rect 7358 11473 7393 11507
rect 7427 11473 7462 11507
rect 7496 11473 7531 11507
rect 7565 11473 7600 11507
rect 7634 11473 7669 11507
rect 7703 11473 7738 11507
rect 7772 11473 7807 11507
rect 7841 11473 7875 11507
rect 7909 11473 7943 11507
rect 7977 11473 8011 11507
rect 8045 11473 8079 11507
rect 8113 11473 8147 11507
rect 8181 11473 8215 11507
rect 8249 11473 8283 11507
rect 8317 11473 8351 11507
rect 8385 11473 8419 11507
rect 8453 11473 8487 11507
rect 8521 11473 8555 11507
rect 8589 11473 8623 11507
rect 8657 11473 8691 11507
rect 8725 11473 8759 11507
rect 8793 11473 8827 11507
rect 8861 11473 8895 11507
rect 8929 11473 8963 11507
rect 8997 11473 9031 11507
rect 9065 11473 9099 11507
rect 9133 11473 9167 11507
rect 9201 11473 9235 11507
rect 9269 11473 9303 11507
rect 9337 11473 9371 11507
rect 9405 11473 9439 11507
rect 9473 11473 9507 11507
rect 9541 11473 9575 11507
rect 9609 11473 9643 11507
rect 9677 11473 9711 11507
rect 9745 11473 9779 11507
rect 9813 11473 9847 11507
rect 9881 11473 9915 11507
rect 9949 11473 9983 11507
rect 10017 11473 10051 11507
rect 10085 11473 10119 11507
rect 10153 11473 10187 11507
rect 10221 11473 10255 11507
rect 10289 11473 10323 11507
rect 10357 11473 10391 11507
rect 10425 11473 10459 11507
rect 10493 11473 10527 11507
rect 10561 11473 10595 11507
rect 10629 11473 10663 11507
rect 10697 11473 10731 11507
rect 10765 11473 10799 11507
rect 10833 11473 10867 11507
rect 10901 11473 10935 11507
rect 10969 11473 11003 11507
rect 11037 11473 11071 11507
rect 11105 11473 11139 11507
rect 11173 11473 11207 11507
rect 11241 11473 11275 11507
rect 11309 11473 11343 11507
rect 11377 11473 11411 11507
rect 11445 11473 11479 11507
rect 11513 11473 11547 11507
rect 11581 11473 11615 11507
rect 11649 11473 11683 11507
rect 11717 11473 11751 11507
rect 11785 11473 11819 11507
rect 11853 11473 11887 11507
rect 11921 11473 11955 11507
rect 11989 11473 12023 11507
rect 12057 11473 12091 11507
rect 12125 11473 12159 11507
rect 12193 11473 12227 11507
rect 12261 11473 12295 11507
rect 12329 11473 12363 11507
rect 12397 11473 12431 11507
rect 12465 11473 12499 11507
rect 12533 11473 12567 11507
rect 12601 11473 12635 11507
rect 12669 11473 12703 11507
rect 12737 11473 12771 11507
rect 12805 11473 12839 11507
rect 12873 11473 12907 11507
rect 12941 11473 12975 11507
rect 13009 11473 13043 11507
rect 13077 11473 13111 11507
rect 13145 11473 13179 11507
rect 13213 11473 13247 11507
rect 13281 11473 13315 11507
rect 13349 11473 13383 11507
rect 13417 11473 13451 11507
rect 13485 11473 13519 11507
rect 13553 11473 13587 11507
rect 13621 11473 13655 11507
rect 13689 11473 13723 11507
rect 13757 11473 13791 11507
rect 13825 11473 13859 11507
rect 13893 11473 13927 11507
rect 13961 11473 13995 11507
rect 14029 11473 14063 11507
rect 14097 11473 14131 11507
rect 14165 11473 14199 11507
rect 14233 11473 14267 11507
rect 14301 11473 14335 11507
rect 14369 11473 14403 11507
rect 14437 11473 14471 11507
rect 14505 11473 14539 11507
rect 14573 11473 14607 11507
rect 14641 11473 14675 11507
rect 14709 11473 14743 11507
rect 14777 11473 14811 11507
rect 14845 11473 14879 11507
rect 14913 11473 14947 11507
rect 14981 11473 15015 11507
rect 15049 11473 15083 11507
rect 15117 11473 15151 11507
rect 15185 11473 15219 11507
rect 15253 11473 15287 11507
rect 15321 11473 15355 11507
rect 15389 11473 15423 11507
rect 15457 11473 15491 11507
rect 15525 11473 15578 11507
rect 5753 11446 15578 11473
rect 5685 11440 15578 11446
rect 5617 11437 15578 11440
rect 5554 11435 15578 11437
rect 5554 11410 5806 11435
rect 5554 11404 5719 11410
rect 5554 11401 5651 11404
rect 5554 11367 5583 11401
rect 5617 11370 5651 11401
rect 5685 11376 5719 11404
rect 5753 11401 5806 11410
rect 5840 11401 5875 11435
rect 5909 11401 5944 11435
rect 5978 11401 6013 11435
rect 6047 11401 6082 11435
rect 6116 11401 6151 11435
rect 6185 11401 6220 11435
rect 6254 11401 6289 11435
rect 6323 11401 6358 11435
rect 6392 11401 6427 11435
rect 6461 11401 6496 11435
rect 6530 11401 6565 11435
rect 6599 11401 6634 11435
rect 6668 11401 6703 11435
rect 6737 11401 6772 11435
rect 6806 11401 6841 11435
rect 6875 11401 6910 11435
rect 6944 11401 6979 11435
rect 7013 11401 7048 11435
rect 7082 11401 7117 11435
rect 7151 11401 7186 11435
rect 7220 11401 7255 11435
rect 7289 11401 7324 11435
rect 7358 11401 7393 11435
rect 7427 11401 7462 11435
rect 7496 11401 7531 11435
rect 7565 11401 7600 11435
rect 7634 11401 7669 11435
rect 7703 11401 7738 11435
rect 7772 11401 7807 11435
rect 7841 11401 7875 11435
rect 7909 11401 7943 11435
rect 7977 11401 8011 11435
rect 8045 11401 8079 11435
rect 8113 11401 8147 11435
rect 8181 11401 8215 11435
rect 8249 11401 8283 11435
rect 8317 11401 8351 11435
rect 8385 11401 8419 11435
rect 8453 11401 8487 11435
rect 8521 11401 8555 11435
rect 8589 11401 8623 11435
rect 8657 11401 8691 11435
rect 8725 11401 8759 11435
rect 8793 11401 8827 11435
rect 8861 11401 8895 11435
rect 8929 11401 8963 11435
rect 8997 11401 9031 11435
rect 9065 11401 9099 11435
rect 9133 11401 9167 11435
rect 9201 11401 9235 11435
rect 9269 11401 9303 11435
rect 9337 11401 9371 11435
rect 9405 11401 9439 11435
rect 9473 11401 9507 11435
rect 9541 11401 9575 11435
rect 9609 11401 9643 11435
rect 9677 11401 9711 11435
rect 9745 11401 9779 11435
rect 9813 11401 9847 11435
rect 9881 11401 9915 11435
rect 9949 11401 9983 11435
rect 10017 11401 10051 11435
rect 10085 11401 10119 11435
rect 10153 11401 10187 11435
rect 10221 11401 10255 11435
rect 10289 11401 10323 11435
rect 10357 11401 10391 11435
rect 10425 11401 10459 11435
rect 10493 11401 10527 11435
rect 10561 11401 10595 11435
rect 10629 11401 10663 11435
rect 10697 11401 10731 11435
rect 10765 11401 10799 11435
rect 10833 11401 10867 11435
rect 10901 11401 10935 11435
rect 10969 11401 11003 11435
rect 11037 11401 11071 11435
rect 11105 11401 11139 11435
rect 11173 11401 11207 11435
rect 11241 11401 11275 11435
rect 11309 11401 11343 11435
rect 11377 11401 11411 11435
rect 11445 11401 11479 11435
rect 11513 11401 11547 11435
rect 11581 11401 11615 11435
rect 11649 11401 11683 11435
rect 11717 11401 11751 11435
rect 11785 11401 11819 11435
rect 11853 11401 11887 11435
rect 11921 11401 11955 11435
rect 11989 11401 12023 11435
rect 12057 11401 12091 11435
rect 12125 11401 12159 11435
rect 12193 11401 12227 11435
rect 12261 11401 12295 11435
rect 12329 11401 12363 11435
rect 12397 11401 12431 11435
rect 12465 11401 12499 11435
rect 12533 11401 12567 11435
rect 12601 11401 12635 11435
rect 12669 11401 12703 11435
rect 12737 11401 12771 11435
rect 12805 11401 12839 11435
rect 12873 11401 12907 11435
rect 12941 11401 12975 11435
rect 13009 11401 13043 11435
rect 13077 11401 13111 11435
rect 13145 11401 13179 11435
rect 13213 11401 13247 11435
rect 13281 11401 13315 11435
rect 13349 11401 13383 11435
rect 13417 11401 13451 11435
rect 13485 11401 13519 11435
rect 13553 11401 13587 11435
rect 13621 11401 13655 11435
rect 13689 11401 13723 11435
rect 13757 11401 13791 11435
rect 13825 11401 13859 11435
rect 13893 11401 13927 11435
rect 13961 11401 13995 11435
rect 14029 11401 14063 11435
rect 14097 11401 14131 11435
rect 14165 11401 14199 11435
rect 14233 11401 14267 11435
rect 14301 11401 14335 11435
rect 14369 11401 14403 11435
rect 14437 11401 14471 11435
rect 14505 11401 14539 11435
rect 14573 11401 14607 11435
rect 14641 11401 14675 11435
rect 14709 11401 14743 11435
rect 14777 11401 14811 11435
rect 14845 11401 14879 11435
rect 14913 11401 14947 11435
rect 14981 11401 15015 11435
rect 15049 11401 15083 11435
rect 15117 11401 15151 11435
rect 15185 11401 15219 11435
rect 15253 11401 15287 11435
rect 15321 11401 15355 11435
rect 15389 11401 15423 11435
rect 15457 11401 15491 11435
rect 15525 11401 15578 11435
rect 5753 11376 15578 11401
rect 5685 11370 15578 11376
rect 5617 11367 15578 11370
rect 5554 11363 15578 11367
rect 5554 11340 5806 11363
rect 5554 11334 5719 11340
rect 5554 11331 5651 11334
rect 5554 11297 5583 11331
rect 5617 11300 5651 11331
rect 5685 11306 5719 11334
rect 5753 11329 5806 11340
rect 5840 11329 5875 11363
rect 5909 11329 5944 11363
rect 5978 11329 6013 11363
rect 6047 11329 6082 11363
rect 6116 11329 6151 11363
rect 6185 11329 6220 11363
rect 6254 11329 6289 11363
rect 6323 11329 6358 11363
rect 6392 11329 6427 11363
rect 6461 11329 6496 11363
rect 6530 11329 6565 11363
rect 6599 11329 6634 11363
rect 6668 11329 6703 11363
rect 6737 11329 6772 11363
rect 6806 11329 6841 11363
rect 6875 11329 6910 11363
rect 6944 11329 6979 11363
rect 7013 11329 7048 11363
rect 7082 11329 7117 11363
rect 7151 11329 7186 11363
rect 7220 11329 7255 11363
rect 7289 11329 7324 11363
rect 7358 11329 7393 11363
rect 7427 11329 7462 11363
rect 7496 11329 7531 11363
rect 7565 11329 7600 11363
rect 7634 11329 7669 11363
rect 7703 11329 7738 11363
rect 7772 11329 7807 11363
rect 7841 11329 7875 11363
rect 7909 11329 7943 11363
rect 7977 11329 8011 11363
rect 8045 11329 8079 11363
rect 8113 11329 8147 11363
rect 8181 11329 8215 11363
rect 8249 11329 8283 11363
rect 8317 11329 8351 11363
rect 8385 11329 8419 11363
rect 8453 11329 8487 11363
rect 8521 11329 8555 11363
rect 8589 11329 8623 11363
rect 8657 11329 8691 11363
rect 8725 11329 8759 11363
rect 8793 11329 8827 11363
rect 8861 11329 8895 11363
rect 8929 11329 8963 11363
rect 8997 11329 9031 11363
rect 9065 11329 9099 11363
rect 9133 11329 9167 11363
rect 9201 11329 9235 11363
rect 9269 11329 9303 11363
rect 9337 11329 9371 11363
rect 9405 11329 9439 11363
rect 9473 11329 9507 11363
rect 9541 11329 9575 11363
rect 9609 11329 9643 11363
rect 9677 11329 9711 11363
rect 9745 11329 9779 11363
rect 9813 11329 9847 11363
rect 9881 11329 9915 11363
rect 9949 11329 9983 11363
rect 10017 11329 10051 11363
rect 10085 11329 10119 11363
rect 10153 11329 10187 11363
rect 10221 11329 10255 11363
rect 10289 11329 10323 11363
rect 10357 11329 10391 11363
rect 10425 11329 10459 11363
rect 10493 11329 10527 11363
rect 10561 11329 10595 11363
rect 10629 11329 10663 11363
rect 10697 11329 10731 11363
rect 10765 11329 10799 11363
rect 10833 11329 10867 11363
rect 10901 11329 10935 11363
rect 10969 11329 11003 11363
rect 11037 11329 11071 11363
rect 11105 11329 11139 11363
rect 11173 11329 11207 11363
rect 11241 11329 11275 11363
rect 11309 11329 11343 11363
rect 11377 11329 11411 11363
rect 11445 11329 11479 11363
rect 11513 11329 11547 11363
rect 11581 11329 11615 11363
rect 11649 11329 11683 11363
rect 11717 11329 11751 11363
rect 11785 11329 11819 11363
rect 11853 11329 11887 11363
rect 11921 11329 11955 11363
rect 11989 11329 12023 11363
rect 12057 11329 12091 11363
rect 12125 11329 12159 11363
rect 12193 11329 12227 11363
rect 12261 11329 12295 11363
rect 12329 11329 12363 11363
rect 12397 11329 12431 11363
rect 12465 11329 12499 11363
rect 12533 11329 12567 11363
rect 12601 11329 12635 11363
rect 12669 11329 12703 11363
rect 12737 11329 12771 11363
rect 12805 11329 12839 11363
rect 12873 11329 12907 11363
rect 12941 11329 12975 11363
rect 13009 11329 13043 11363
rect 13077 11329 13111 11363
rect 13145 11329 13179 11363
rect 13213 11329 13247 11363
rect 13281 11329 13315 11363
rect 13349 11329 13383 11363
rect 13417 11329 13451 11363
rect 13485 11329 13519 11363
rect 13553 11329 13587 11363
rect 13621 11329 13655 11363
rect 13689 11329 13723 11363
rect 13757 11329 13791 11363
rect 13825 11329 13859 11363
rect 13893 11329 13927 11363
rect 13961 11329 13995 11363
rect 14029 11329 14063 11363
rect 14097 11329 14131 11363
rect 14165 11329 14199 11363
rect 14233 11329 14267 11363
rect 14301 11329 14335 11363
rect 14369 11329 14403 11363
rect 14437 11329 14471 11363
rect 14505 11329 14539 11363
rect 14573 11329 14607 11363
rect 14641 11329 14675 11363
rect 14709 11329 14743 11363
rect 14777 11329 14811 11363
rect 14845 11329 14879 11363
rect 14913 11329 14947 11363
rect 14981 11329 15015 11363
rect 15049 11329 15083 11363
rect 15117 11329 15151 11363
rect 15185 11329 15219 11363
rect 15253 11329 15287 11363
rect 15321 11329 15355 11363
rect 15389 11329 15423 11363
rect 15457 11329 15491 11363
rect 15525 11329 15578 11363
rect 5753 11306 15578 11329
rect 5685 11300 15578 11306
rect 5617 11297 15578 11300
rect 5554 11291 15578 11297
rect 5554 11270 5806 11291
rect 5554 11264 5719 11270
rect 5554 11261 5651 11264
rect 5554 11227 5583 11261
rect 5617 11230 5651 11261
rect 5685 11236 5719 11264
rect 5753 11257 5806 11270
rect 5840 11257 5875 11291
rect 5909 11257 5944 11291
rect 5978 11257 6013 11291
rect 6047 11257 6082 11291
rect 6116 11257 6151 11291
rect 6185 11257 6220 11291
rect 6254 11257 6289 11291
rect 6323 11257 6358 11291
rect 6392 11257 6427 11291
rect 6461 11257 6496 11291
rect 6530 11257 6565 11291
rect 6599 11257 6634 11291
rect 6668 11257 6703 11291
rect 6737 11257 6772 11291
rect 6806 11257 6841 11291
rect 6875 11257 6910 11291
rect 6944 11257 6979 11291
rect 7013 11257 7048 11291
rect 7082 11257 7117 11291
rect 7151 11257 7186 11291
rect 7220 11257 7255 11291
rect 7289 11257 7324 11291
rect 7358 11257 7393 11291
rect 7427 11257 7462 11291
rect 7496 11257 7531 11291
rect 7565 11257 7600 11291
rect 7634 11257 7669 11291
rect 7703 11257 7738 11291
rect 7772 11257 7807 11291
rect 7841 11257 7875 11291
rect 7909 11257 7943 11291
rect 7977 11257 8011 11291
rect 8045 11257 8079 11291
rect 8113 11257 8147 11291
rect 8181 11257 8215 11291
rect 8249 11257 8283 11291
rect 8317 11257 8351 11291
rect 8385 11257 8419 11291
rect 8453 11257 8487 11291
rect 8521 11257 8555 11291
rect 8589 11257 8623 11291
rect 8657 11257 8691 11291
rect 8725 11257 8759 11291
rect 8793 11257 8827 11291
rect 8861 11257 8895 11291
rect 8929 11257 8963 11291
rect 8997 11257 9031 11291
rect 9065 11257 9099 11291
rect 9133 11257 9167 11291
rect 9201 11257 9235 11291
rect 9269 11257 9303 11291
rect 9337 11257 9371 11291
rect 9405 11257 9439 11291
rect 9473 11257 9507 11291
rect 9541 11257 9575 11291
rect 9609 11257 9643 11291
rect 9677 11257 9711 11291
rect 9745 11257 9779 11291
rect 9813 11257 9847 11291
rect 9881 11257 9915 11291
rect 9949 11257 9983 11291
rect 10017 11257 10051 11291
rect 10085 11257 10119 11291
rect 10153 11257 10187 11291
rect 10221 11257 10255 11291
rect 10289 11257 10323 11291
rect 10357 11257 10391 11291
rect 10425 11257 10459 11291
rect 10493 11257 10527 11291
rect 10561 11257 10595 11291
rect 10629 11257 10663 11291
rect 10697 11257 10731 11291
rect 10765 11257 10799 11291
rect 10833 11257 10867 11291
rect 10901 11257 10935 11291
rect 10969 11257 11003 11291
rect 11037 11257 11071 11291
rect 11105 11257 11139 11291
rect 11173 11257 11207 11291
rect 11241 11257 11275 11291
rect 11309 11257 11343 11291
rect 11377 11257 11411 11291
rect 11445 11257 11479 11291
rect 11513 11257 11547 11291
rect 11581 11257 11615 11291
rect 11649 11257 11683 11291
rect 11717 11257 11751 11291
rect 11785 11257 11819 11291
rect 11853 11257 11887 11291
rect 11921 11257 11955 11291
rect 11989 11257 12023 11291
rect 12057 11257 12091 11291
rect 12125 11257 12159 11291
rect 12193 11257 12227 11291
rect 12261 11257 12295 11291
rect 12329 11257 12363 11291
rect 12397 11257 12431 11291
rect 12465 11257 12499 11291
rect 12533 11257 12567 11291
rect 12601 11257 12635 11291
rect 12669 11257 12703 11291
rect 12737 11257 12771 11291
rect 12805 11257 12839 11291
rect 12873 11257 12907 11291
rect 12941 11257 12975 11291
rect 13009 11257 13043 11291
rect 13077 11257 13111 11291
rect 13145 11257 13179 11291
rect 13213 11257 13247 11291
rect 13281 11257 13315 11291
rect 13349 11257 13383 11291
rect 13417 11257 13451 11291
rect 13485 11257 13519 11291
rect 13553 11257 13587 11291
rect 13621 11257 13655 11291
rect 13689 11257 13723 11291
rect 13757 11257 13791 11291
rect 13825 11257 13859 11291
rect 13893 11257 13927 11291
rect 13961 11257 13995 11291
rect 14029 11257 14063 11291
rect 14097 11257 14131 11291
rect 14165 11257 14199 11291
rect 14233 11257 14267 11291
rect 14301 11257 14335 11291
rect 14369 11257 14403 11291
rect 14437 11257 14471 11291
rect 14505 11257 14539 11291
rect 14573 11257 14607 11291
rect 14641 11257 14675 11291
rect 14709 11257 14743 11291
rect 14777 11257 14811 11291
rect 14845 11257 14879 11291
rect 14913 11257 14947 11291
rect 14981 11257 15015 11291
rect 15049 11257 15083 11291
rect 15117 11257 15151 11291
rect 15185 11257 15219 11291
rect 15253 11257 15287 11291
rect 15321 11257 15355 11291
rect 15389 11257 15423 11291
rect 15457 11257 15491 11291
rect 15525 11257 15578 11291
rect 5753 11236 15578 11257
rect 5685 11230 15578 11236
rect 5617 11227 15578 11230
rect 5554 11219 15578 11227
rect 5554 11200 5806 11219
rect 5554 11194 5719 11200
rect 5554 11191 5651 11194
rect 5554 11157 5583 11191
rect 5617 11160 5651 11191
rect 5685 11166 5719 11194
rect 5753 11185 5806 11200
rect 5840 11185 5875 11219
rect 5909 11185 5944 11219
rect 5978 11185 6013 11219
rect 6047 11185 6082 11219
rect 6116 11185 6151 11219
rect 6185 11185 6220 11219
rect 6254 11185 6289 11219
rect 6323 11185 6358 11219
rect 6392 11185 6427 11219
rect 6461 11185 6496 11219
rect 6530 11185 6565 11219
rect 6599 11185 6634 11219
rect 6668 11185 6703 11219
rect 6737 11185 6772 11219
rect 6806 11185 6841 11219
rect 6875 11185 6910 11219
rect 6944 11185 6979 11219
rect 7013 11185 7048 11219
rect 7082 11185 7117 11219
rect 7151 11185 7186 11219
rect 7220 11185 7255 11219
rect 7289 11185 7324 11219
rect 7358 11185 7393 11219
rect 7427 11185 7462 11219
rect 7496 11185 7531 11219
rect 7565 11185 7600 11219
rect 7634 11185 7669 11219
rect 7703 11185 7738 11219
rect 7772 11185 7807 11219
rect 7841 11185 7875 11219
rect 7909 11185 7943 11219
rect 7977 11185 8011 11219
rect 8045 11185 8079 11219
rect 8113 11185 8147 11219
rect 8181 11185 8215 11219
rect 8249 11185 8283 11219
rect 8317 11185 8351 11219
rect 8385 11185 8419 11219
rect 8453 11185 8487 11219
rect 8521 11185 8555 11219
rect 8589 11185 8623 11219
rect 8657 11185 8691 11219
rect 8725 11185 8759 11219
rect 8793 11185 8827 11219
rect 8861 11185 8895 11219
rect 8929 11185 8963 11219
rect 8997 11185 9031 11219
rect 9065 11185 9099 11219
rect 9133 11185 9167 11219
rect 9201 11185 9235 11219
rect 9269 11185 9303 11219
rect 9337 11185 9371 11219
rect 9405 11185 9439 11219
rect 9473 11185 9507 11219
rect 9541 11185 9575 11219
rect 9609 11185 9643 11219
rect 9677 11185 9711 11219
rect 9745 11185 9779 11219
rect 9813 11185 9847 11219
rect 9881 11185 9915 11219
rect 9949 11185 9983 11219
rect 10017 11185 10051 11219
rect 10085 11185 10119 11219
rect 10153 11185 10187 11219
rect 10221 11185 10255 11219
rect 10289 11185 10323 11219
rect 10357 11185 10391 11219
rect 10425 11185 10459 11219
rect 10493 11185 10527 11219
rect 10561 11185 10595 11219
rect 10629 11185 10663 11219
rect 10697 11185 10731 11219
rect 10765 11185 10799 11219
rect 10833 11185 10867 11219
rect 10901 11185 10935 11219
rect 10969 11185 11003 11219
rect 11037 11185 11071 11219
rect 11105 11185 11139 11219
rect 11173 11185 11207 11219
rect 11241 11185 11275 11219
rect 11309 11185 11343 11219
rect 11377 11185 11411 11219
rect 11445 11185 11479 11219
rect 11513 11185 11547 11219
rect 11581 11185 11615 11219
rect 11649 11185 11683 11219
rect 11717 11185 11751 11219
rect 11785 11185 11819 11219
rect 11853 11185 11887 11219
rect 11921 11185 11955 11219
rect 11989 11185 12023 11219
rect 12057 11185 12091 11219
rect 12125 11185 12159 11219
rect 12193 11185 12227 11219
rect 12261 11185 12295 11219
rect 12329 11185 12363 11219
rect 12397 11185 12431 11219
rect 12465 11185 12499 11219
rect 12533 11185 12567 11219
rect 12601 11185 12635 11219
rect 12669 11185 12703 11219
rect 12737 11185 12771 11219
rect 12805 11185 12839 11219
rect 12873 11185 12907 11219
rect 12941 11185 12975 11219
rect 13009 11185 13043 11219
rect 13077 11185 13111 11219
rect 13145 11185 13179 11219
rect 13213 11185 13247 11219
rect 13281 11185 13315 11219
rect 13349 11185 13383 11219
rect 13417 11185 13451 11219
rect 13485 11185 13519 11219
rect 13553 11185 13587 11219
rect 13621 11185 13655 11219
rect 13689 11185 13723 11219
rect 13757 11185 13791 11219
rect 13825 11185 13859 11219
rect 13893 11185 13927 11219
rect 13961 11185 13995 11219
rect 14029 11185 14063 11219
rect 14097 11185 14131 11219
rect 14165 11185 14199 11219
rect 14233 11185 14267 11219
rect 14301 11185 14335 11219
rect 14369 11185 14403 11219
rect 14437 11185 14471 11219
rect 14505 11185 14539 11219
rect 14573 11185 14607 11219
rect 14641 11185 14675 11219
rect 14709 11185 14743 11219
rect 14777 11185 14811 11219
rect 14845 11185 14879 11219
rect 14913 11185 14947 11219
rect 14981 11185 15015 11219
rect 15049 11185 15083 11219
rect 15117 11185 15151 11219
rect 15185 11185 15219 11219
rect 15253 11185 15287 11219
rect 15321 11185 15355 11219
rect 15389 11185 15423 11219
rect 15457 11185 15491 11219
rect 15525 11185 15578 11219
rect 5753 11181 15578 11185
rect 5753 11166 5782 11181
rect 5685 11160 5782 11166
rect 5617 11157 5782 11160
rect 5554 11130 5782 11157
rect 5554 11124 5719 11130
rect 5554 11121 5651 11124
rect 5554 11087 5583 11121
rect 5617 11090 5651 11121
rect 5685 11096 5719 11124
rect 5753 11096 5782 11130
rect 5685 11090 5782 11096
rect 5617 11087 5782 11090
rect 5554 11060 5782 11087
rect 5554 11054 5719 11060
rect 5554 11051 5651 11054
rect 5554 11017 5583 11051
rect 5617 11020 5651 11051
rect 5685 11026 5719 11054
rect 5753 11026 5782 11060
rect 5685 11020 5782 11026
rect 5617 11017 5782 11020
rect 5554 10990 5782 11017
rect 5554 10984 5719 10990
rect 5554 10981 5651 10984
rect 5554 10947 5583 10981
rect 5617 10950 5651 10981
rect 5685 10956 5719 10984
rect 5753 10956 5782 10990
rect 5685 10950 5782 10956
rect 5617 10947 5782 10950
rect 5554 10920 5782 10947
rect 5554 10914 5719 10920
rect 5554 10911 5651 10914
rect 5554 10877 5583 10911
rect 5617 10880 5651 10911
rect 5685 10886 5719 10914
rect 5753 10886 5782 10920
rect 5685 10880 5782 10886
rect 5617 10877 5782 10880
rect 5554 10850 5782 10877
rect 5554 10844 5719 10850
rect 5554 10841 5651 10844
rect 5554 10807 5583 10841
rect 5617 10810 5651 10841
rect 5685 10816 5719 10844
rect 5753 10816 5782 10850
rect 5685 10810 5782 10816
rect 5617 10807 5782 10810
rect 5554 10780 5782 10807
rect 5554 10774 5719 10780
rect 5554 10771 5651 10774
rect 5554 10737 5583 10771
rect 5617 10740 5651 10771
rect 5685 10746 5719 10774
rect 5753 10746 5782 10780
rect 5685 10740 5782 10746
rect 5617 10737 5782 10740
rect 5554 10710 5782 10737
rect 5554 10704 5719 10710
rect 5554 10701 5651 10704
rect 5554 10667 5583 10701
rect 5617 10670 5651 10701
rect 5685 10676 5719 10704
rect 5753 10676 5782 10710
rect 5685 10670 5782 10676
rect 5617 10667 5782 10670
rect 5554 10640 5782 10667
rect 5554 10634 5719 10640
rect 5554 10631 5651 10634
rect 5554 10597 5583 10631
rect 5617 10600 5651 10631
rect 5685 10606 5719 10634
rect 5753 10606 5782 10640
rect 5685 10600 5782 10606
rect 5617 10597 5782 10600
rect 5554 10570 5782 10597
rect 5554 10564 5719 10570
rect 5554 10561 5651 10564
rect 5554 10531 5583 10561
rect 5617 10531 5651 10561
rect 5685 10536 5719 10564
rect 5753 10536 5782 10570
rect 5685 10531 5782 10536
rect -76 10497 -48 10521
rect -14 10497 25 10531
rect 59 10497 98 10531
rect 132 10497 171 10531
rect 205 10497 244 10531
rect 278 10497 317 10531
rect 351 10497 390 10531
rect 424 10497 463 10531
rect 497 10497 536 10531
rect 570 10497 609 10531
rect 643 10497 682 10531
rect 716 10497 755 10531
rect 789 10497 828 10531
rect 862 10497 901 10531
rect 935 10497 974 10531
rect 1008 10497 1047 10531
rect 1081 10497 1120 10531
rect 1154 10497 1193 10531
rect 1227 10497 1266 10531
rect 1300 10497 1339 10531
rect 1373 10497 1412 10531
rect 1446 10497 1485 10531
rect 1519 10497 1558 10531
rect 1592 10497 1631 10531
rect 1665 10497 1704 10531
rect 1738 10497 1777 10531
rect 1811 10497 1850 10531
rect 1884 10497 1923 10531
rect -76 10492 1923 10497
rect -76 10322 -52 10492
rect 1546 10459 1581 10492
rect 1615 10459 1650 10492
rect 1684 10459 1719 10492
rect 1753 10459 1788 10492
rect 1822 10459 1857 10492
rect 1546 10425 1558 10459
rect 1615 10458 1631 10459
rect 1684 10458 1704 10459
rect 1753 10458 1777 10459
rect 1822 10458 1850 10459
rect 1891 10458 1923 10492
rect 1592 10425 1631 10458
rect 1665 10425 1704 10458
rect 1738 10425 1777 10458
rect 1811 10425 1850 10458
rect 1884 10425 1923 10458
rect 1546 10424 1923 10425
rect 1614 10390 1649 10424
rect 1683 10390 1718 10424
rect 1752 10390 1787 10424
rect 1821 10390 1856 10424
rect 1890 10390 1923 10424
rect 1614 10387 1923 10390
rect 1614 10353 1631 10387
rect 1665 10356 1704 10387
rect 1738 10356 1777 10387
rect 1811 10356 1850 10387
rect 1884 10356 1923 10387
rect 1682 10353 1704 10356
rect 1750 10353 1777 10356
rect 1818 10353 1850 10356
rect 1614 10322 1648 10353
rect 1682 10322 1716 10353
rect 1750 10322 1784 10353
rect 1818 10322 1852 10353
rect 1886 10322 1920 10356
rect 5773 10353 5782 10531
rect 1954 10322 1988 10353
rect 2022 10322 2057 10353
rect 2091 10322 2126 10353
rect 2160 10322 2195 10353
rect 2229 10322 2264 10353
rect 2298 10322 2333 10353
rect 2367 10322 2402 10353
rect 2436 10322 2471 10353
rect 2505 10322 2540 10353
rect 2574 10322 2609 10353
rect 2643 10322 2678 10353
rect 2712 10322 2747 10353
rect 2781 10322 2816 10353
rect 2850 10322 2885 10353
rect 2919 10322 2954 10353
rect 2988 10322 3023 10353
rect 3057 10322 3092 10353
rect 3126 10322 3161 10353
rect 3195 10322 3230 10353
rect 3264 10322 3299 10353
rect 3333 10322 3368 10353
rect 3402 10322 3437 10353
rect 3471 10322 3506 10353
rect 3540 10322 3575 10353
rect 3609 10322 3644 10353
rect 3678 10322 3713 10353
rect 3747 10322 3782 10353
rect 3816 10322 3851 10353
rect 3885 10322 3920 10353
rect 3954 10322 3989 10353
rect 4023 10322 4058 10353
rect 4092 10322 4127 10353
rect 4161 10322 4196 10353
rect 4230 10322 4265 10353
rect 4299 10322 4334 10353
rect 4368 10322 4403 10353
rect 4437 10322 4472 10353
rect 4506 10322 4541 10353
rect 4575 10322 4610 10353
rect 4644 10322 4679 10353
rect 4713 10322 4748 10353
rect 4782 10322 4817 10353
rect 4851 10322 4886 10353
rect 4920 10322 4955 10353
rect 4989 10322 5024 10353
rect 5058 10322 5093 10353
rect 5127 10322 5162 10353
rect 5196 10322 5231 10353
rect 5265 10322 5300 10353
rect 5334 10322 5369 10353
rect 5403 10322 5438 10353
rect 5472 10322 5507 10353
rect 5541 10322 5576 10353
rect 5610 10322 5645 10353
rect 5679 10322 5714 10353
rect 5748 10322 5782 10353
rect -76 10293 5782 10322
rect 14611 10247 15055 10252
rect 14611 10213 14623 10247
rect 14657 10213 14695 10247
rect 14729 10213 14949 10247
rect 14983 10213 15021 10247
rect 14611 10208 15055 10213
rect 17 10110 56 10144
rect 90 10110 129 10144
rect 163 10110 202 10144
rect 236 10110 275 10144
rect 309 10110 348 10144
rect 382 10110 421 10144
rect 455 10110 494 10144
rect 528 10110 567 10144
rect 601 10110 640 10144
rect 674 10110 713 10144
rect 747 10110 786 10144
rect 820 10110 859 10144
rect 893 10110 932 10144
rect 966 10110 1005 10144
rect 1039 10110 1078 10144
rect 1112 10110 1151 10144
rect 1185 10110 1224 10144
rect 1258 10110 1297 10144
rect 1331 10110 1370 10144
rect 1404 10110 1443 10144
rect 1477 10110 1516 10144
rect 1550 10110 1589 10144
rect 1623 10110 1662 10144
rect 1696 10110 1735 10144
rect 1769 10110 1808 10144
rect 1842 10110 1881 10144
rect 1915 10110 1954 10144
rect 1988 10110 2027 10144
rect 2061 10110 2100 10144
rect 2134 10110 2173 10144
rect 2207 10110 2246 10144
rect 2280 10110 2319 10144
rect 2353 10110 2392 10144
rect 2426 10110 2465 10144
rect 2499 10110 2538 10144
rect 2572 10110 2611 10144
rect 2645 10110 2684 10144
rect 2718 10110 2757 10144
rect 2791 10110 2830 10144
rect 2864 10110 2903 10144
rect 2937 10110 2976 10144
rect 3010 10110 3049 10144
rect 3083 10110 3122 10144
rect 3156 10110 3195 10144
rect 3229 10110 3268 10144
rect 3302 10110 3341 10144
rect 3375 10110 3414 10144
rect 3448 10110 3487 10144
rect 3521 10110 3560 10144
rect 3594 10110 3633 10144
rect 3667 10110 3706 10144
rect 3740 10110 3779 10144
rect 3813 10110 3852 10144
rect 3886 10110 3925 10144
rect 3959 10110 3998 10144
rect 4032 10110 4071 10144
rect 4105 10110 4144 10144
rect 4178 10110 4216 10144
rect 4250 10110 4288 10144
rect 4322 10110 4360 10144
rect 4394 10110 4432 10144
rect 4466 10110 4504 10144
rect 4538 10110 4576 10144
rect 4610 10110 4648 10144
rect 4682 10110 4720 10144
rect 4754 10110 4792 10144
rect 4826 10110 4864 10144
rect 4898 10110 4936 10144
rect 4970 10110 5008 10144
rect 5042 10110 5080 10144
rect 5114 10110 5152 10144
rect 5186 10110 5224 10144
rect 5258 10110 5296 10144
rect 5330 10110 5368 10144
rect 5402 10110 5440 10144
rect 5474 10110 5512 10144
rect 5546 10110 5584 10144
rect 5618 10110 5656 10144
rect 5690 10110 5728 10144
rect 5762 10110 5800 10144
rect 5834 10110 5872 10144
rect 5906 10110 5944 10144
rect 5978 10110 6016 10144
rect 6050 10110 6088 10144
rect 6122 10110 6160 10144
rect 6194 10110 6232 10144
rect 6266 10110 6304 10144
rect 6338 10110 6376 10144
rect 6410 10110 6448 10144
rect 6482 10110 6520 10144
rect 6554 10110 6592 10144
rect 6626 10110 6664 10144
rect 6698 10110 6736 10144
rect 6770 10110 6808 10144
rect 6842 10110 6880 10144
rect 6914 10110 6952 10144
rect 6986 10110 7024 10144
rect 7058 10110 7096 10144
rect 7130 10110 7168 10144
rect 7202 10110 7240 10144
rect 7274 10110 7312 10144
rect 7346 10110 7384 10144
rect 7418 10110 7456 10144
rect 7490 10110 7528 10144
rect 7562 10110 7600 10144
rect 7634 10110 7672 10144
rect 7706 10110 7744 10144
rect 7778 10110 7816 10144
rect 7850 10110 7888 10144
rect 7922 10110 7960 10144
rect 7994 10110 8032 10144
rect 8066 10110 8104 10144
rect 8138 10110 8176 10144
rect 8210 10110 8248 10144
rect 8282 10110 8320 10144
rect 8354 10110 8392 10144
rect 8426 10110 8464 10144
rect 8498 10110 8536 10144
rect 8570 10110 8608 10144
rect 8642 10110 8680 10144
rect 8714 10110 8752 10144
rect 8786 10110 8824 10144
rect 8858 10110 8896 10144
rect 8930 10110 8968 10144
rect 9002 10110 9040 10144
rect 9074 10110 9112 10144
rect 9146 10110 9184 10144
rect 9218 10110 9256 10144
rect 9290 10110 9328 10144
rect 9362 10110 9400 10144
rect 9434 10110 9472 10144
rect 9506 10110 9544 10144
rect 9578 10110 9616 10144
rect 9650 10110 9688 10144
rect 9722 10110 9760 10144
rect 9794 10110 9832 10144
rect 9866 10110 9904 10144
rect 9938 10110 9976 10144
rect 10010 10110 10048 10144
rect 10082 10110 10120 10144
rect 10154 10110 10192 10144
rect 10226 10110 10264 10144
rect 10298 10110 10336 10144
rect 10370 10110 10408 10144
rect 10442 10110 10480 10144
rect 10514 10110 10552 10144
rect 10586 10110 10624 10144
rect 10658 10110 10696 10144
rect 10730 10110 10768 10144
rect 10802 10110 10840 10144
rect 10874 10110 10912 10144
rect 10946 10110 10984 10144
rect 11018 10110 11056 10144
rect 11090 10110 11128 10144
rect 11162 10110 11200 10144
rect 11234 10110 11272 10144
rect 11306 10110 11344 10144
rect 11378 10110 11416 10144
rect 11450 10110 11488 10144
rect 11522 10110 11560 10144
rect 11594 10110 11632 10144
rect 11666 10110 11704 10144
rect 11738 10110 11776 10144
rect 11810 10110 11848 10144
rect 11882 10110 11920 10144
rect 11954 10110 11992 10144
rect 12026 10110 12064 10144
rect 12098 10110 12136 10144
rect 12170 10110 12208 10144
rect 12242 10141 12280 10144
rect 12314 10141 12352 10144
rect 12386 10141 12424 10144
rect 12458 10141 12496 10144
rect 12530 10141 12568 10144
rect 12602 10141 12640 10144
rect 12674 10141 12712 10144
rect 12980 10141 13020 10144
rect 13054 10141 13093 10144
rect 13127 10141 13166 10144
rect 13200 10141 13239 10144
rect 13273 10141 13312 10144
rect 13346 10141 13385 10144
rect 13419 10141 13458 10144
rect 13492 10141 13531 10144
rect 13565 10141 13604 10144
rect 13638 10141 13677 10144
rect 13711 10141 13750 10144
rect 13784 10141 13823 10144
rect 13857 10141 13896 10144
rect 13930 10141 13969 10144
rect 14003 10141 14042 10144
rect 14076 10141 14115 10144
rect 14149 10141 14188 10144
rect 14222 10141 14261 10144
rect 14295 10141 14334 10144
rect 14368 10141 14407 10144
rect 14441 10141 14480 10144
rect 14514 10141 14553 10144
rect 14990 10141 15042 10144
rect 15076 10141 15128 10144
rect 15162 10141 15214 10144
rect 12259 10110 12280 10141
rect 12329 10110 12352 10141
rect 12399 10110 12424 10141
rect 12469 10110 12496 10141
rect 12538 10110 12568 10141
rect 12607 10110 12640 10141
rect 12201 10107 12225 10110
rect 12259 10107 12295 10110
rect 12329 10107 12365 10110
rect 12399 10107 12435 10110
rect 12469 10107 12504 10110
rect 12538 10107 12573 10110
rect 12607 10107 12642 10110
rect 12676 10107 12711 10141
rect 12746 10110 12780 10141
rect 12745 10107 12780 10110
rect 12814 10107 12849 10141
rect 12883 10107 12918 10141
rect 12980 10110 12987 10141
rect 13054 10110 13056 10141
rect 12952 10107 12987 10110
rect 13021 10107 13056 10110
rect 13090 10110 13093 10141
rect 13159 10110 13166 10141
rect 13228 10110 13239 10141
rect 13297 10110 13312 10141
rect 13366 10110 13385 10141
rect 13435 10110 13458 10141
rect 13504 10110 13531 10141
rect 13573 10110 13604 10141
rect 13090 10107 13125 10110
rect 13159 10107 13194 10110
rect 13228 10107 13263 10110
rect 13297 10107 13332 10110
rect 13366 10107 13401 10110
rect 13435 10107 13470 10110
rect 13504 10107 13539 10110
rect 13573 10107 13608 10110
rect 13642 10107 13677 10141
rect 13711 10107 13746 10141
rect 13784 10110 13815 10141
rect 13857 10110 13884 10141
rect 13930 10110 13953 10141
rect 14003 10110 14022 10141
rect 14076 10110 14091 10141
rect 14149 10110 14160 10141
rect 14222 10110 14229 10141
rect 14295 10110 14298 10141
rect 13780 10107 13815 10110
rect 13849 10107 13884 10110
rect 13918 10107 13953 10110
rect 13987 10107 14022 10110
rect 14056 10107 14091 10110
rect 14125 10107 14160 10110
rect 14194 10107 14229 10110
rect 14263 10107 14298 10110
rect 14332 10110 14334 10141
rect 14401 10110 14407 10141
rect 14470 10110 14480 10141
rect 14539 10110 14553 10141
rect 14332 10107 14367 10110
rect 14401 10107 14436 10110
rect 14470 10107 14505 10110
rect 14539 10107 14574 10110
rect 14608 10107 14643 10141
rect 14677 10107 14712 10141
rect 14746 10107 14781 10141
rect 14815 10107 14850 10141
rect 14884 10107 14919 10141
rect 14953 10110 14956 10141
rect 15022 10110 15042 10141
rect 14953 10107 14988 10110
rect 15022 10107 15057 10110
rect 15091 10107 15126 10141
rect 15162 10110 15195 10141
rect 15248 10110 15299 10144
rect 15160 10107 15195 10110
rect 15229 10107 15333 10110
rect 15299 10072 15333 10073
rect -17 9993 17 10038
rect -17 9915 17 9959
rect 14658 9963 14692 10001
rect 14824 10006 14960 10024
rect 14858 9972 14926 10006
rect 14824 9954 14960 9972
rect 15299 9993 15333 10004
rect 15299 9915 15333 9935
rect 15299 9831 15333 9866
rect 4110 9749 4144 9787
rect 4422 9749 4456 9787
rect 4912 9749 4946 9787
rect 5264 9749 5298 9787
rect 6410 9749 6444 9787
rect 6762 9749 6796 9787
rect 7134 9749 7168 9787
rect 7486 9749 7520 9787
rect 15299 9762 15333 9797
rect 15299 9693 15333 9728
rect 15299 9624 15333 9659
rect 15299 9555 15333 9590
rect 15299 9486 15333 9521
rect 15299 9417 15333 9452
rect 15299 9348 15333 9383
rect 15299 9279 15333 9314
rect 15299 9210 15333 9245
rect 15299 9141 15333 9176
rect 11612 8281 11663 9102
rect 15299 9072 15333 9107
rect 15299 9003 15333 9038
rect 15299 8934 15333 8969
rect 15299 8865 15333 8900
rect 15299 8796 15333 8831
rect 15299 8727 15333 8762
rect 15299 8658 15333 8693
rect 15299 8589 15333 8624
rect 15299 8520 15333 8555
rect 15299 8452 15333 8486
rect 15299 8384 15333 8418
rect 15299 8316 15333 8350
rect 11612 8232 14634 8281
rect 15299 8248 15333 8282
rect 11612 7447 11684 8232
rect 15299 8180 15333 8214
rect 14868 7836 15006 8124
rect 14847 7812 15006 7836
rect 14881 7778 14915 7812
rect 14949 7778 15006 7812
rect 15299 8112 15333 8146
rect 15299 8044 15333 8078
rect 15299 7976 15333 8010
rect 15299 7908 15333 7942
rect 14847 7742 15006 7778
rect 15038 7772 15062 7806
rect 15096 7772 15163 7806
rect 15197 7772 15265 7806
rect 15299 7772 15333 7874
rect 15549 9754 15578 11181
rect 15549 9749 15714 9754
rect 15748 9749 15777 11823
rect 15549 9719 15777 9749
rect 15549 9685 15578 9719
rect 15612 9685 15646 9719
rect 15680 9715 15777 9719
rect 15680 9685 15714 9715
rect 15549 9681 15714 9685
rect 15748 9681 15777 9715
rect 15549 9650 15777 9681
rect 15549 9616 15578 9650
rect 15612 9616 15646 9650
rect 15680 9647 15777 9650
rect 15680 9616 15714 9647
rect 15549 9613 15714 9616
rect 15748 9613 15777 9647
rect 15549 9581 15777 9613
rect 15549 9547 15578 9581
rect 15612 9547 15646 9581
rect 15680 9579 15777 9581
rect 15680 9547 15714 9579
rect 15549 9545 15714 9547
rect 15748 9545 15777 9579
rect 15549 9512 15777 9545
rect 15549 9478 15578 9512
rect 15612 9478 15646 9512
rect 15680 9511 15777 9512
rect 15680 9478 15714 9511
rect 15549 9477 15714 9478
rect 15748 9477 15777 9511
rect 15549 9443 15777 9477
rect 15549 9409 15578 9443
rect 15612 9409 15646 9443
rect 15680 9409 15714 9443
rect 15748 9409 15777 9443
rect 15549 9374 15777 9409
rect 15549 9340 15578 9374
rect 15612 9340 15646 9374
rect 15680 9340 15714 9374
rect 15748 9340 15777 9374
rect 15549 9305 15777 9340
rect 15549 9271 15578 9305
rect 15612 9271 15646 9305
rect 15680 9271 15714 9305
rect 15748 9271 15777 9305
rect 15549 9236 15777 9271
rect 15549 9202 15578 9236
rect 15612 9202 15646 9236
rect 15680 9202 15714 9236
rect 15748 9202 15777 9236
rect 15549 9167 15777 9202
rect 15549 9133 15578 9167
rect 15612 9133 15646 9167
rect 15680 9133 15714 9167
rect 15748 9133 15777 9167
rect 15549 9098 15777 9133
rect 15549 9064 15578 9098
rect 15612 9064 15646 9098
rect 15680 9064 15714 9098
rect 15748 9064 15777 9098
rect 15549 9029 15777 9064
rect 15549 8995 15578 9029
rect 15612 8995 15646 9029
rect 15680 8995 15714 9029
rect 15748 8995 15777 9029
rect 15549 8960 15777 8995
rect 15549 8926 15578 8960
rect 15612 8926 15646 8960
rect 15680 8926 15714 8960
rect 15748 8926 15777 8960
rect 15549 8891 15777 8926
rect 15549 8857 15578 8891
rect 15612 8857 15646 8891
rect 15680 8857 15714 8891
rect 15748 8857 15777 8891
rect 15549 8822 15777 8857
rect 15549 8788 15578 8822
rect 15612 8788 15646 8822
rect 15680 8788 15714 8822
rect 15748 8788 15777 8822
rect 15549 8753 15777 8788
rect 15549 8719 15578 8753
rect 15612 8719 15646 8753
rect 15680 8719 15714 8753
rect 15748 8719 15777 8753
rect 15549 8684 15777 8719
rect 15549 8650 15578 8684
rect 15612 8650 15646 8684
rect 15680 8650 15714 8684
rect 15748 8650 15777 8684
rect 15549 8615 15777 8650
rect 15549 8581 15578 8615
rect 15612 8581 15646 8615
rect 15680 8581 15714 8615
rect 15748 8581 15777 8615
rect 15549 8546 15777 8581
rect 15549 8512 15578 8546
rect 15612 8512 15646 8546
rect 15680 8512 15714 8546
rect 15748 8512 15777 8546
rect 15549 8477 15777 8512
rect 15549 8443 15578 8477
rect 15612 8443 15646 8477
rect 15680 8443 15714 8477
rect 15748 8443 15777 8477
rect 15549 8408 15777 8443
rect 15549 8374 15578 8408
rect 15612 8374 15646 8408
rect 15680 8374 15714 8408
rect 15748 8374 15777 8408
rect 15549 8339 15777 8374
rect 15549 8305 15578 8339
rect 15612 8305 15646 8339
rect 15680 8305 15714 8339
rect 15748 8305 15777 8339
rect 15549 8270 15777 8305
rect 15549 8236 15578 8270
rect 15612 8236 15646 8270
rect 15680 8236 15714 8270
rect 15748 8236 15777 8270
rect 15549 8201 15777 8236
rect 15549 8167 15578 8201
rect 15612 8167 15646 8201
rect 15680 8167 15714 8201
rect 15748 8167 15777 8201
rect 15549 8132 15777 8167
rect 15549 8098 15578 8132
rect 15612 8098 15646 8132
rect 15680 8098 15714 8132
rect 15748 8098 15777 8132
rect 15549 8063 15777 8098
rect 15549 8029 15578 8063
rect 15612 8029 15646 8063
rect 15680 8029 15714 8063
rect 15748 8029 15777 8063
rect 15549 7994 15777 8029
rect 15549 7960 15578 7994
rect 15612 7960 15646 7994
rect 15680 7960 15714 7994
rect 15748 7960 15777 7994
rect 15549 7925 15777 7960
rect 15549 7891 15578 7925
rect 15612 7891 15646 7925
rect 15680 7891 15714 7925
rect 15748 7891 15777 7925
rect 15549 7856 15777 7891
rect 15549 7822 15578 7856
rect 15612 7822 15646 7856
rect 15680 7822 15714 7856
rect 15748 7822 15777 7856
rect 15549 7787 15777 7822
rect 14881 7708 14915 7742
rect 14949 7708 15006 7742
rect 14847 7672 15006 7708
rect 14881 7638 14915 7672
rect 14949 7638 15006 7672
rect 14847 7602 15006 7638
rect 14881 7568 14915 7602
rect 14949 7568 15006 7602
rect 14847 7532 15006 7568
rect 14881 7498 14915 7532
rect 14949 7498 15006 7532
rect 14847 7462 15006 7498
rect 14881 7428 14915 7462
rect 14949 7428 15006 7462
rect 14847 7391 15006 7428
rect 14881 7357 14915 7391
rect 14949 7357 15006 7391
rect 14847 7320 15006 7357
rect 14881 7286 14915 7320
rect 14949 7286 15006 7320
rect 14847 7249 15006 7286
rect 14881 7215 14915 7249
rect 14949 7215 15006 7249
rect 14847 7178 15006 7215
rect 14881 7144 14915 7178
rect 14949 7144 15006 7178
rect 14847 7107 15006 7144
rect 14881 7073 14915 7107
rect 14949 7073 15006 7107
rect 14847 7036 15006 7073
rect 14881 7002 14915 7036
rect 14949 7002 15006 7036
rect 14847 6965 15006 7002
rect 11514 6908 11548 6946
rect 14881 6931 14915 6965
rect 14949 6931 15006 6965
rect 14847 6894 15006 6931
rect 14881 6860 14915 6894
rect 14949 6860 15006 6894
rect 14847 6823 15006 6860
rect 14881 6789 14915 6823
rect 14949 6789 15006 6823
rect 14847 6752 15006 6789
rect 14881 6718 14915 6752
rect 14949 6718 15006 6752
rect 14847 6681 15006 6718
rect 14881 6647 14915 6681
rect 14949 6647 15006 6681
rect 14847 6610 15006 6647
rect 14881 6576 14915 6610
rect 14949 6576 15006 6610
rect 14847 6539 15006 6576
rect 14881 6505 14915 6539
rect 14949 6505 15006 6539
rect 14847 6468 15006 6505
rect 14881 6434 14915 6468
rect 14949 6434 15006 6468
rect 14847 6397 15006 6434
rect 14881 6363 14915 6397
rect 14949 6363 15006 6397
rect 14847 6326 15006 6363
rect 14881 6292 14915 6326
rect 14949 6292 15006 6326
rect 14847 6268 15006 6292
rect 14868 6030 15006 6268
rect 15549 7753 15578 7787
rect 15612 7753 15646 7787
rect 15680 7753 15714 7787
rect 15748 7753 15777 7787
rect 15549 7718 15777 7753
rect 15549 7684 15578 7718
rect 15612 7684 15646 7718
rect 15680 7684 15714 7718
rect 15748 7684 15777 7718
rect 15549 7649 15777 7684
rect 15549 7615 15578 7649
rect 15612 7615 15646 7649
rect 15680 7615 15714 7649
rect 15748 7615 15777 7649
rect 15549 7580 15777 7615
rect 15549 7546 15578 7580
rect 15612 7546 15646 7580
rect 15680 7546 15714 7580
rect 15748 7546 15777 7580
rect 15549 7511 15777 7546
rect 15549 7477 15578 7511
rect 15612 7477 15646 7511
rect 15680 7477 15714 7511
rect 15748 7477 15777 7511
rect 15549 7442 15777 7477
rect 15549 7408 15578 7442
rect 15612 7408 15646 7442
rect 15680 7408 15714 7442
rect 15748 7408 15777 7442
rect 15549 7373 15777 7408
rect 15549 7339 15578 7373
rect 15612 7339 15646 7373
rect 15680 7339 15714 7373
rect 15748 7339 15777 7373
rect 15549 7304 15777 7339
rect 15549 7270 15578 7304
rect 15612 7270 15646 7304
rect 15680 7270 15714 7304
rect 15748 7270 15777 7304
rect 15549 7235 15777 7270
rect 15549 7201 15578 7235
rect 15612 7201 15646 7235
rect 15680 7201 15714 7235
rect 15748 7201 15777 7235
rect 15549 7166 15777 7201
rect 15549 7132 15578 7166
rect 15612 7132 15646 7166
rect 15680 7132 15714 7166
rect 15748 7132 15777 7166
rect 15549 7097 15777 7132
rect 15549 7063 15578 7097
rect 15612 7063 15646 7097
rect 15680 7063 15714 7097
rect 15748 7063 15777 7097
rect 15549 7028 15777 7063
rect 15549 6994 15578 7028
rect 15612 6994 15646 7028
rect 15680 6994 15714 7028
rect 15748 6994 15777 7028
rect 15549 6959 15777 6994
rect 15549 6925 15578 6959
rect 15612 6925 15646 6959
rect 15680 6925 15714 6959
rect 15748 6925 15777 6959
rect 15549 6890 15777 6925
rect 15549 6856 15578 6890
rect 15612 6856 15646 6890
rect 15680 6856 15714 6890
rect 15748 6856 15777 6890
rect 15549 6821 15777 6856
rect 15549 6787 15578 6821
rect 15612 6787 15646 6821
rect 15680 6787 15714 6821
rect 15748 6787 15777 6821
rect 15549 6752 15777 6787
rect 15549 6718 15578 6752
rect 15612 6718 15646 6752
rect 15680 6718 15714 6752
rect 15748 6718 15777 6752
rect 15549 6683 15777 6718
rect 15549 6649 15578 6683
rect 15612 6649 15646 6683
rect 15680 6649 15714 6683
rect 15748 6649 15777 6683
rect 15549 6614 15777 6649
rect 15549 6580 15578 6614
rect 15612 6580 15646 6614
rect 15680 6580 15714 6614
rect 15748 6580 15777 6614
rect 15549 6545 15777 6580
rect 15549 6511 15578 6545
rect 15612 6511 15646 6545
rect 15680 6511 15714 6545
rect 15748 6511 15777 6545
rect 15549 6476 15777 6511
rect 15549 6442 15578 6476
rect 15612 6442 15646 6476
rect 15680 6442 15714 6476
rect 15748 6442 15777 6476
rect 15549 6407 15777 6442
rect 15549 6373 15578 6407
rect 15612 6373 15646 6407
rect 15680 6373 15714 6407
rect 15748 6373 15777 6407
rect 15549 6338 15777 6373
rect 15549 6304 15578 6338
rect 15612 6304 15646 6338
rect 15680 6304 15714 6338
rect 15748 6304 15777 6338
rect 15549 6269 15777 6304
rect 15549 6235 15578 6269
rect 15612 6235 15646 6269
rect 15680 6235 15714 6269
rect 15748 6235 15777 6269
rect 15549 6200 15777 6235
rect 15549 6166 15578 6200
rect 15612 6166 15646 6200
rect 15680 6166 15714 6200
rect 15748 6166 15777 6200
rect 15549 6131 15777 6166
rect 15549 6097 15578 6131
rect 15612 6097 15646 6131
rect 15680 6097 15714 6131
rect 15748 6097 15777 6131
rect 15549 6062 15777 6097
rect 15549 6028 15578 6062
rect 15612 6028 15646 6062
rect 15680 6028 15714 6062
rect 15748 6028 15777 6062
rect 11424 5878 11458 5916
rect 14553 5936 14587 5974
rect 15549 5993 15777 6028
rect 15549 5959 15578 5993
rect 15612 5959 15646 5993
rect 15680 5959 15714 5993
rect 15748 5959 15777 5993
rect 15549 5924 15777 5959
rect 15549 5890 15578 5924
rect 15612 5890 15646 5924
rect 15680 5890 15714 5924
rect 15748 5890 15777 5924
rect 15549 5855 15777 5890
rect 15549 5821 15578 5855
rect 15612 5821 15646 5855
rect 15680 5821 15714 5855
rect 15748 5821 15777 5855
rect 15549 5786 15777 5821
rect 15549 5752 15578 5786
rect 15612 5752 15646 5786
rect 15680 5752 15714 5786
rect 15748 5752 15777 5786
rect 15549 5717 15777 5752
rect 15549 5683 15578 5717
rect 15612 5683 15646 5717
rect 15680 5683 15714 5717
rect 15748 5683 15777 5717
rect 15549 5648 15777 5683
rect 15549 5614 15578 5648
rect 15612 5614 15646 5648
rect 15680 5614 15714 5648
rect 15748 5614 15777 5648
rect 15549 5579 15777 5614
rect 15549 5545 15578 5579
rect 15612 5545 15646 5579
rect 15680 5545 15714 5579
rect 15748 5545 15777 5579
rect 15549 5510 15777 5545
rect 15549 5476 15578 5510
rect 15612 5476 15646 5510
rect 15680 5476 15714 5510
rect 15748 5476 15777 5510
rect 15549 5441 15777 5476
rect 15549 5407 15578 5441
rect 15612 5407 15646 5441
rect 15680 5407 15714 5441
rect 15748 5407 15777 5441
rect 15549 5372 15777 5407
rect 15549 5338 15578 5372
rect 15612 5338 15646 5372
rect 15680 5338 15714 5372
rect 15748 5338 15777 5372
rect 15549 5303 15777 5338
rect 15549 5269 15578 5303
rect 15612 5269 15646 5303
rect 15680 5269 15714 5303
rect 15748 5269 15777 5303
rect 15549 5234 15777 5269
rect 15549 5200 15578 5234
rect 15612 5200 15646 5234
rect 15680 5200 15714 5234
rect 15748 5200 15777 5234
rect 15549 5181 15777 5200
rect 15170 5165 16042 5181
rect 15170 5164 15578 5165
rect 15612 5164 15646 5165
rect 15680 5164 15714 5165
rect 15748 5164 16042 5165
rect 15204 5130 15247 5164
rect 15281 5130 15324 5164
rect 15358 5130 15400 5164
rect 15434 5130 15476 5164
rect 15510 5130 15552 5164
rect 15612 5131 15628 5164
rect 15680 5131 15704 5164
rect 15748 5131 15780 5164
rect 15586 5130 15628 5131
rect 15662 5130 15704 5131
rect 15738 5130 15780 5131
rect 15814 5130 15856 5164
rect 15890 5130 15932 5164
rect 15966 5130 16008 5164
rect 15170 5123 16042 5130
rect 15170 5092 16045 5123
rect 15204 5058 15247 5092
rect 15281 5058 15324 5092
rect 15358 5058 15400 5092
rect 15434 5058 15476 5092
rect 15510 5058 15552 5092
rect 15586 5058 15628 5092
rect 15662 5058 15704 5092
rect 15738 5058 15780 5092
rect 15814 5058 15856 5092
rect 15890 5058 15932 5092
rect 15966 5058 16008 5092
rect 16042 5058 16045 5092
rect 15170 5020 16045 5058
rect 15204 4986 15247 5020
rect 15281 4986 15324 5020
rect 15358 4986 15400 5020
rect 15434 4986 15476 5020
rect 15510 4986 15552 5020
rect 15586 4986 15628 5020
rect 15662 4986 15704 5020
rect 15738 4986 15780 5020
rect 15814 4986 15856 5020
rect 15890 4986 15932 5020
rect 15966 4986 16008 5020
rect 16042 4986 16045 5020
rect 15170 4756 16045 4986
rect 425 4718 448 4734
rect 15829 4688 16045 4756
rect 11613 3617 11633 3651
rect 11667 3617 11687 3651
rect 11613 3579 11687 3617
rect 11613 3545 11633 3579
rect 11667 3545 11687 3579
rect 11613 2680 11687 3545
rect 11631 2419 11648 2429
rect 11952 2407 12058 2558
rect 12407 2457 12843 2528
rect 15139 2525 15183 2562
rect 12441 2423 12488 2457
rect 12522 2423 12569 2457
rect 12603 2423 12649 2457
rect 12683 2423 12729 2457
rect 12763 2423 12809 2457
rect 7418 2368 7552 2402
rect 7586 2368 7624 2402
rect 11986 2373 12024 2407
rect 11952 2370 12058 2373
<< viali >>
rect 1954 13572 1988 13606
rect 2032 13572 2066 13606
rect 2110 13572 2144 13606
rect 2188 13572 2222 13606
rect 2266 13572 2300 13606
rect 2344 13572 2378 13606
rect 2422 13572 2456 13606
rect 2500 13572 2534 13606
rect 2578 13572 2612 13606
rect 1954 13498 1988 13532
rect 2032 13498 2066 13532
rect 2110 13498 2144 13532
rect 2188 13498 2222 13532
rect 2266 13498 2300 13532
rect 2344 13498 2378 13532
rect 2422 13498 2456 13532
rect 2500 13498 2534 13532
rect 2578 13498 2612 13532
rect 1954 13424 1988 13458
rect 2032 13424 2066 13458
rect 2110 13424 2144 13458
rect 2188 13424 2222 13458
rect 2266 13424 2300 13458
rect 2344 13424 2378 13458
rect 2422 13424 2456 13458
rect 2500 13424 2534 13458
rect 2578 13424 2612 13458
rect 1954 13349 1988 13383
rect 2032 13349 2066 13383
rect 2110 13349 2144 13383
rect 2188 13349 2222 13383
rect 2266 13349 2300 13383
rect 2344 13349 2378 13383
rect 2422 13349 2456 13383
rect 2500 13349 2534 13383
rect 2578 13349 2612 13383
rect 1954 13274 1988 13308
rect 2032 13274 2066 13308
rect 2110 13274 2144 13308
rect 2188 13274 2222 13308
rect 2266 13274 2300 13308
rect 2344 13274 2378 13308
rect 2422 13274 2456 13308
rect 2500 13274 2534 13308
rect 2578 13274 2612 13308
rect 1954 13199 1988 13233
rect 2032 13199 2066 13233
rect 2110 13199 2144 13233
rect 2188 13199 2222 13233
rect 2266 13199 2300 13233
rect 2344 13199 2378 13233
rect 2422 13199 2456 13233
rect 2500 13199 2534 13233
rect 2578 13199 2612 13233
rect 1954 13124 1988 13158
rect 2032 13124 2066 13158
rect 2110 13124 2144 13158
rect 2188 13124 2222 13158
rect 2266 13124 2300 13158
rect 2344 13124 2378 13158
rect 2422 13124 2456 13158
rect 2500 13124 2534 13158
rect 2578 13124 2612 13158
rect 1954 13049 1988 13083
rect 2032 13049 2066 13083
rect 2110 13049 2144 13083
rect 2188 13049 2222 13083
rect 2266 13049 2300 13083
rect 2344 13049 2378 13083
rect 2422 13049 2456 13083
rect 2500 13049 2534 13083
rect 2578 13049 2612 13083
rect 1954 12974 1988 13008
rect 2032 12974 2066 13008
rect 2110 12974 2144 13008
rect 2188 12974 2222 13008
rect 2266 12974 2300 13008
rect 2344 12974 2378 13008
rect 2422 12974 2456 13008
rect 2500 12974 2534 13008
rect 2578 12974 2612 13008
rect 1954 12899 1988 12933
rect 2032 12899 2066 12933
rect 2110 12899 2144 12933
rect 2188 12899 2222 12933
rect 2266 12899 2300 12933
rect 2344 12899 2378 12933
rect 2422 12899 2456 12933
rect 2500 12899 2534 12933
rect 2578 12899 2612 12933
rect 1934 12330 1968 12364
rect 2008 12330 2042 12364
rect 2082 12330 2116 12364
rect 2156 12330 2190 12364
rect 2230 12330 2264 12364
rect 2304 12330 2338 12364
rect 2378 12330 2412 12364
rect 2452 12330 2486 12364
rect 2526 12330 2560 12364
rect 2600 12330 2634 12364
rect 2674 12330 2708 12364
rect 2748 12330 2782 12364
rect 2822 12330 2856 12364
rect 2896 12330 2930 12364
rect 2970 12330 3004 12364
rect 3044 12330 3078 12364
rect 3118 12330 3152 12364
rect 3192 12330 3226 12364
rect 3266 12330 3300 12364
rect 3340 12330 3374 12364
rect 3414 12330 3448 12364
rect 3488 12330 3522 12364
rect 3562 12330 3596 12364
rect 3636 12330 3670 12364
rect 3710 12330 3744 12364
rect 3784 12330 3818 12364
rect 3858 12330 3892 12364
rect 3931 12330 3965 12364
rect 4004 12330 4038 12364
rect 4077 12330 4111 12364
rect 4150 12330 4184 12364
rect 4223 12330 4257 12364
rect 1934 12248 1968 12282
rect 2008 12248 2042 12282
rect 2082 12248 2116 12282
rect 2156 12248 2190 12282
rect 2230 12248 2264 12282
rect 2304 12248 2338 12282
rect 2378 12248 2412 12282
rect 2452 12248 2486 12282
rect 2526 12248 2560 12282
rect 2600 12248 2634 12282
rect 2674 12248 2708 12282
rect 2748 12248 2782 12282
rect 2822 12248 2856 12282
rect 2896 12248 2930 12282
rect 2970 12248 3004 12282
rect 3044 12248 3078 12282
rect 3118 12248 3152 12282
rect 3192 12248 3226 12282
rect 3266 12248 3300 12282
rect 3340 12248 3374 12282
rect 3414 12248 3448 12282
rect 3488 12248 3522 12282
rect 3562 12248 3596 12282
rect 3636 12248 3670 12282
rect 3710 12248 3744 12282
rect 3784 12248 3818 12282
rect 3858 12248 3892 12282
rect 3931 12248 3965 12282
rect 4004 12248 4038 12282
rect 4077 12248 4111 12282
rect 4150 12248 4184 12282
rect 4223 12248 4257 12282
rect -2911 12203 -2877 12237
rect -2838 12203 -2804 12237
rect -2765 12203 -2731 12237
rect -2692 12203 -2658 12237
rect -2619 12203 -2585 12237
rect -2546 12203 -2512 12237
rect -2473 12203 -2439 12237
rect -2400 12203 -2366 12237
rect -2327 12203 -2293 12237
rect -2254 12203 -2220 12237
rect -2181 12203 -2147 12237
rect -2108 12203 -2074 12237
rect -2035 12203 -2001 12237
rect -1962 12203 -1928 12237
rect -1889 12203 -1855 12237
rect -1816 12203 -1782 12237
rect -2911 12131 -2877 12165
rect -2838 12131 -2804 12165
rect -2765 12131 -2731 12165
rect -2692 12131 -2658 12165
rect -2619 12131 -2585 12165
rect -2546 12131 -2512 12165
rect -2473 12131 -2439 12165
rect -2400 12131 -2366 12165
rect -2327 12131 -2293 12165
rect -2254 12131 -2220 12165
rect -2181 12131 -2147 12165
rect -2108 12131 -2074 12165
rect -2035 12131 -2001 12165
rect -1962 12131 -1928 12165
rect -1889 12131 -1855 12165
rect -1816 12131 -1782 12165
rect -2911 12059 -2877 12093
rect -2838 12059 -2804 12093
rect -2765 12059 -2731 12093
rect -2692 12059 -2658 12093
rect -2619 12059 -2585 12093
rect -2546 12059 -2512 12093
rect -2473 12059 -2439 12093
rect -2400 12059 -2366 12093
rect -2327 12059 -2293 12093
rect -2254 12059 -2220 12093
rect -2181 12059 -2147 12093
rect -2108 12059 -2074 12093
rect -2035 12059 -2001 12093
rect -1962 12059 -1928 12093
rect -1889 12059 -1855 12093
rect -1816 12059 -1782 12093
rect -2911 11987 -2877 12021
rect -2838 11987 -2804 12021
rect -2765 11987 -2731 12021
rect -2692 11987 -2658 12021
rect -2619 11987 -2585 12021
rect -2546 11987 -2512 12021
rect -2473 11987 -2439 12021
rect -2400 11987 -2366 12021
rect -2327 11987 -2293 12021
rect -2254 11987 -2220 12021
rect -2181 11987 -2147 12021
rect -2108 11987 -2074 12021
rect -2035 11987 -2001 12021
rect -1962 11987 -1928 12021
rect -1889 11987 -1855 12021
rect -1816 11987 -1782 12021
rect -2911 11915 -2877 11949
rect -2838 11915 -2804 11949
rect -2765 11915 -2731 11949
rect -2692 11915 -2658 11949
rect -2619 11915 -2585 11949
rect -2546 11915 -2512 11949
rect -2473 11915 -2439 11949
rect -2400 11915 -2366 11949
rect -2327 11915 -2293 11949
rect -2254 11915 -2220 11949
rect -2181 11915 -2147 11949
rect -2108 11915 -2074 11949
rect -2035 11915 -2001 11949
rect -1962 11915 -1928 11949
rect -1889 11915 -1855 11949
rect -1816 11915 -1782 11949
rect -2911 11843 -2877 11877
rect -2838 11843 -2804 11877
rect -2765 11843 -2731 11877
rect -2692 11843 -2658 11877
rect -2619 11843 -2585 11877
rect -2546 11843 -2512 11877
rect -2473 11843 -2439 11877
rect -2400 11843 -2366 11877
rect -2327 11843 -2293 11877
rect -2254 11843 -2220 11877
rect -2181 11843 -2147 11877
rect -2108 11843 -2074 11877
rect -2035 11843 -2001 11877
rect -1962 11843 -1928 11877
rect -1889 11843 -1855 11877
rect -1816 11843 -1782 11877
rect -2911 11771 -2877 11805
rect -2838 11771 -2804 11805
rect -2765 11771 -2731 11805
rect -2692 11771 -2658 11805
rect -2619 11771 -2585 11805
rect -2546 11771 -2512 11805
rect -2473 11771 -2439 11805
rect -2400 11771 -2366 11805
rect -2327 11771 -2293 11805
rect -2254 11771 -2220 11805
rect -2181 11771 -2147 11805
rect -2108 11771 -2074 11805
rect -2035 11771 -2001 11805
rect -1962 11771 -1928 11805
rect -1889 11771 -1855 11805
rect -1816 11771 -1782 11805
rect -1743 11771 307 12237
rect 1934 12166 1968 12200
rect 2008 12166 2042 12200
rect 2082 12166 2116 12200
rect 2156 12166 2190 12200
rect 2230 12166 2264 12200
rect 2304 12166 2338 12200
rect 2378 12166 2412 12200
rect 2452 12166 2486 12200
rect 2526 12166 2560 12200
rect 2600 12166 2634 12200
rect 2674 12166 2708 12200
rect 2748 12166 2782 12200
rect 2822 12166 2856 12200
rect 2896 12166 2930 12200
rect 2970 12166 3004 12200
rect 3044 12166 3078 12200
rect 3118 12166 3152 12200
rect 3192 12166 3226 12200
rect 3266 12166 3300 12200
rect 3340 12166 3374 12200
rect 3414 12166 3448 12200
rect 3488 12166 3522 12200
rect 3562 12166 3596 12200
rect 3636 12166 3670 12200
rect 3710 12166 3744 12200
rect 3784 12166 3818 12200
rect 3858 12166 3892 12200
rect 3931 12166 3965 12200
rect 4004 12166 4038 12200
rect 4077 12166 4111 12200
rect 4150 12166 4184 12200
rect 4223 12166 4257 12200
rect 1934 12084 1968 12118
rect 2008 12084 2042 12118
rect 2082 12084 2116 12118
rect 2156 12084 2190 12118
rect 2230 12084 2264 12118
rect 2304 12084 2338 12118
rect 2378 12084 2412 12118
rect 2452 12084 2486 12118
rect 2526 12084 2560 12118
rect 2600 12084 2634 12118
rect 2674 12084 2708 12118
rect 2748 12084 2782 12118
rect 2822 12084 2856 12118
rect 2896 12084 2930 12118
rect 2970 12084 3004 12118
rect 3044 12084 3078 12118
rect 3118 12084 3152 12118
rect 3192 12084 3226 12118
rect 3266 12084 3300 12118
rect 3340 12084 3374 12118
rect 3414 12084 3448 12118
rect 3488 12084 3522 12118
rect 3562 12084 3596 12118
rect 3636 12084 3670 12118
rect 3710 12084 3744 12118
rect 3784 12084 3818 12118
rect 3858 12084 3892 12118
rect 3931 12084 3965 12118
rect 4004 12084 4038 12118
rect 4077 12084 4111 12118
rect 4150 12084 4184 12118
rect 4223 12084 4257 12118
rect 1934 12002 1968 12036
rect 2008 12002 2042 12036
rect 2082 12002 2116 12036
rect 2156 12002 2190 12036
rect 2230 12002 2264 12036
rect 2304 12002 2338 12036
rect 2378 12002 2412 12036
rect 2452 12002 2486 12036
rect 2526 12002 2560 12036
rect 2600 12002 2634 12036
rect 2674 12002 2708 12036
rect 2748 12002 2782 12036
rect 2822 12002 2856 12036
rect 2896 12002 2930 12036
rect 2970 12002 3004 12036
rect 3044 12002 3078 12036
rect 3118 12002 3152 12036
rect 3192 12002 3226 12036
rect 3266 12002 3300 12036
rect 3340 12002 3374 12036
rect 3414 12002 3448 12036
rect 3488 12002 3522 12036
rect 3562 12002 3596 12036
rect 3636 12002 3670 12036
rect 3710 12002 3744 12036
rect 3784 12002 3818 12036
rect 3858 12002 3892 12036
rect 3931 12002 3965 12036
rect 4004 12002 4038 12036
rect 4077 12002 4111 12036
rect 4150 12002 4184 12036
rect 4223 12002 4257 12036
rect 367 11942 401 11976
rect 441 11942 475 11976
rect 515 11942 549 11976
rect 588 11942 622 11976
rect 661 11942 695 11976
rect 734 11942 768 11976
rect 807 11942 841 11976
rect 880 11942 914 11976
rect 953 11942 987 11976
rect 1026 11942 1060 11976
rect 1099 11942 1133 11976
rect 1172 11942 1206 11976
rect 1245 11942 1279 11976
rect 1318 11942 1352 11976
rect 1391 11942 1425 11976
rect 1464 11942 1498 11976
rect 1537 11942 1571 11976
rect 1610 11942 1644 11976
rect 1683 11942 1717 11976
rect 367 11854 401 11888
rect 441 11854 475 11888
rect 515 11854 549 11888
rect 588 11854 622 11888
rect 661 11854 695 11888
rect 734 11854 768 11888
rect 807 11854 841 11888
rect 880 11854 914 11888
rect 953 11854 987 11888
rect 1026 11854 1060 11888
rect 1099 11854 1133 11888
rect 1172 11854 1206 11888
rect 1245 11854 1279 11888
rect 1318 11854 1352 11888
rect 1391 11854 1425 11888
rect 1464 11854 1498 11888
rect 1537 11854 1571 11888
rect 1610 11854 1644 11888
rect 1683 11854 1717 11888
rect 367 11766 401 11800
rect 441 11766 475 11800
rect 515 11766 549 11800
rect 588 11766 622 11800
rect 661 11766 695 11800
rect 734 11766 768 11800
rect 807 11766 841 11800
rect 880 11766 914 11800
rect 953 11766 987 11800
rect 1026 11766 1060 11800
rect 1099 11766 1133 11800
rect 1172 11766 1206 11800
rect 1245 11766 1279 11800
rect 1318 11766 1352 11800
rect 1391 11766 1425 11800
rect 1464 11766 1498 11800
rect 1537 11766 1571 11800
rect 1610 11766 1644 11800
rect 1683 11766 1717 11800
rect -48 10497 -14 10531
rect 25 10497 59 10531
rect 98 10497 132 10531
rect 171 10497 205 10531
rect 244 10497 278 10531
rect 317 10497 351 10531
rect 390 10497 424 10531
rect 463 10497 497 10531
rect 536 10497 570 10531
rect 609 10497 643 10531
rect 682 10497 716 10531
rect 755 10497 789 10531
rect 828 10497 862 10531
rect 901 10497 935 10531
rect 974 10497 1008 10531
rect 1047 10497 1081 10531
rect 1120 10497 1154 10531
rect 1193 10497 1227 10531
rect 1266 10497 1300 10531
rect 1339 10497 1373 10531
rect 1412 10497 1446 10531
rect 1485 10497 1519 10531
rect 1558 10497 1592 10531
rect 1631 10497 1665 10531
rect 1704 10497 1738 10531
rect 1777 10497 1811 10531
rect 1850 10497 1884 10531
rect 1923 10527 5583 10531
rect 5583 10527 5617 10531
rect 5617 10530 5651 10531
rect 5651 10530 5685 10531
rect 5685 10530 5773 10531
rect 5617 10527 5773 10530
rect 1923 10500 5773 10527
rect 1923 10494 5719 10500
rect 1923 10492 5651 10494
rect -48 10425 -14 10459
rect 25 10425 59 10459
rect 98 10425 132 10459
rect 171 10425 205 10459
rect 244 10425 278 10459
rect 317 10425 351 10459
rect 390 10425 424 10459
rect 463 10425 497 10459
rect 536 10425 570 10459
rect 609 10425 643 10459
rect 682 10425 716 10459
rect 755 10425 789 10459
rect 828 10425 862 10459
rect 901 10425 935 10459
rect 974 10425 1008 10459
rect 1047 10425 1081 10459
rect 1120 10425 1154 10459
rect 1193 10425 1227 10459
rect 1266 10425 1300 10459
rect 1339 10425 1373 10459
rect 1412 10425 1446 10459
rect 1485 10425 1519 10459
rect 1558 10458 1581 10459
rect 1581 10458 1592 10459
rect 1631 10458 1650 10459
rect 1650 10458 1665 10459
rect 1704 10458 1719 10459
rect 1719 10458 1738 10459
rect 1777 10458 1788 10459
rect 1788 10458 1811 10459
rect 1850 10458 1857 10459
rect 1857 10458 1884 10459
rect 1923 10458 1926 10492
rect 1926 10458 1960 10492
rect 1960 10458 1995 10492
rect 1995 10458 2029 10492
rect 2029 10458 2064 10492
rect 2064 10458 2098 10492
rect 2098 10458 2133 10492
rect 2133 10458 2167 10492
rect 2167 10458 2202 10492
rect 2202 10458 2236 10492
rect 2236 10458 2271 10492
rect 2271 10458 2305 10492
rect 2305 10458 2340 10492
rect 2340 10458 2374 10492
rect 2374 10458 2409 10492
rect 2409 10458 2443 10492
rect 2443 10458 2478 10492
rect 2478 10458 2512 10492
rect 2512 10458 2547 10492
rect 2547 10458 2581 10492
rect 2581 10458 2616 10492
rect 2616 10458 2650 10492
rect 2650 10458 2685 10492
rect 2685 10458 2719 10492
rect 2719 10458 2754 10492
rect 2754 10458 2788 10492
rect 2788 10458 2823 10492
rect 2823 10458 2857 10492
rect 2857 10458 2892 10492
rect 2892 10458 2926 10492
rect 2926 10458 2961 10492
rect 2961 10458 2995 10492
rect 2995 10458 3030 10492
rect 3030 10458 3064 10492
rect 3064 10458 3099 10492
rect 3099 10458 3133 10492
rect 3133 10458 3168 10492
rect 3168 10458 3202 10492
rect 3202 10458 3237 10492
rect 3237 10458 3271 10492
rect 3271 10458 3306 10492
rect 3306 10458 3340 10492
rect 3340 10458 3375 10492
rect 3375 10458 3409 10492
rect 3409 10458 3444 10492
rect 3444 10458 3478 10492
rect 3478 10458 3513 10492
rect 3513 10458 3547 10492
rect 3547 10458 3582 10492
rect 3582 10458 3616 10492
rect 3616 10458 3651 10492
rect 3651 10458 3685 10492
rect 3685 10458 3720 10492
rect 3720 10458 3754 10492
rect 3754 10458 3789 10492
rect 3789 10458 3823 10492
rect 3823 10458 3858 10492
rect 3858 10458 3892 10492
rect 3892 10458 3927 10492
rect 3927 10458 3961 10492
rect 3961 10458 3996 10492
rect 3996 10458 4030 10492
rect 4030 10458 4065 10492
rect 4065 10458 4099 10492
rect 4099 10458 4134 10492
rect 4134 10458 4168 10492
rect 4168 10458 4203 10492
rect 4203 10458 4237 10492
rect 4237 10458 4272 10492
rect 4272 10458 4306 10492
rect 4306 10458 4341 10492
rect 4341 10458 4375 10492
rect 4375 10458 4410 10492
rect 4410 10458 4444 10492
rect 4444 10458 4479 10492
rect 4479 10458 4513 10492
rect 4513 10458 4548 10492
rect 4548 10458 4582 10492
rect 4582 10458 4617 10492
rect 4617 10458 4651 10492
rect 4651 10458 4686 10492
rect 4686 10458 4720 10492
rect 4720 10458 4755 10492
rect 4755 10458 4789 10492
rect 4789 10458 4824 10492
rect 4824 10458 4858 10492
rect 4858 10458 4893 10492
rect 4893 10458 4927 10492
rect 4927 10458 4962 10492
rect 4962 10458 4996 10492
rect 4996 10458 5031 10492
rect 5031 10458 5065 10492
rect 5065 10458 5100 10492
rect 5100 10458 5134 10492
rect 5134 10458 5169 10492
rect 5169 10458 5203 10492
rect 5203 10458 5238 10492
rect 5238 10458 5272 10492
rect 5272 10458 5307 10492
rect 5307 10458 5341 10492
rect 5341 10458 5376 10492
rect 5376 10458 5410 10492
rect 5410 10458 5445 10492
rect 5445 10458 5479 10492
rect 5479 10458 5514 10492
rect 5514 10458 5548 10492
rect 5548 10458 5583 10492
rect 5583 10458 5617 10492
rect 5617 10460 5651 10492
rect 5651 10460 5685 10494
rect 5685 10466 5719 10494
rect 5719 10466 5753 10500
rect 5753 10466 5773 10500
rect 5685 10460 5773 10466
rect 5617 10458 5773 10460
rect 1558 10425 1592 10458
rect 1631 10425 1665 10458
rect 1704 10425 1738 10458
rect 1777 10425 1811 10458
rect 1850 10425 1884 10458
rect 1923 10431 5773 10458
rect 1923 10424 5719 10431
rect 1923 10390 1925 10424
rect 1925 10390 1959 10424
rect 1959 10390 1994 10424
rect 1994 10390 2028 10424
rect 2028 10390 2063 10424
rect 2063 10390 2097 10424
rect 2097 10390 2132 10424
rect 2132 10390 2166 10424
rect 2166 10390 2201 10424
rect 2201 10390 2235 10424
rect 2235 10390 2270 10424
rect 2270 10390 2304 10424
rect 2304 10390 2339 10424
rect 2339 10390 2373 10424
rect 2373 10390 2408 10424
rect 2408 10390 2442 10424
rect 2442 10390 2477 10424
rect 2477 10390 2511 10424
rect 2511 10390 2546 10424
rect 2546 10390 2580 10424
rect 2580 10390 2615 10424
rect 2615 10390 2649 10424
rect 2649 10390 2684 10424
rect 2684 10390 2718 10424
rect 2718 10390 2753 10424
rect 2753 10390 2787 10424
rect 2787 10390 2822 10424
rect 2822 10390 2856 10424
rect 2856 10390 2891 10424
rect 2891 10390 2925 10424
rect 2925 10390 2960 10424
rect 2960 10390 2994 10424
rect 2994 10390 3029 10424
rect 3029 10390 3063 10424
rect 3063 10390 3098 10424
rect 3098 10390 3132 10424
rect 3132 10390 3167 10424
rect 3167 10390 3201 10424
rect 3201 10390 3236 10424
rect 3236 10390 3270 10424
rect 3270 10390 3305 10424
rect 3305 10390 3339 10424
rect 3339 10390 3374 10424
rect 3374 10390 3408 10424
rect 3408 10390 3443 10424
rect 3443 10390 3477 10424
rect 3477 10390 3512 10424
rect 3512 10390 3546 10424
rect 3546 10390 3581 10424
rect 3581 10390 3615 10424
rect 3615 10390 3650 10424
rect 3650 10390 3684 10424
rect 3684 10390 3719 10424
rect 3719 10390 3753 10424
rect 3753 10390 3788 10424
rect 3788 10390 3822 10424
rect 3822 10390 3857 10424
rect 3857 10390 3891 10424
rect 3891 10390 3926 10424
rect 3926 10390 3960 10424
rect 3960 10390 3995 10424
rect 3995 10390 4029 10424
rect 4029 10390 4064 10424
rect 4064 10390 4098 10424
rect 4098 10390 4133 10424
rect 4133 10390 4167 10424
rect 4167 10390 4202 10424
rect 4202 10390 4236 10424
rect 4236 10390 4271 10424
rect 4271 10390 4305 10424
rect 4305 10390 4340 10424
rect 4340 10390 4374 10424
rect 4374 10390 4409 10424
rect 4409 10390 4443 10424
rect 4443 10390 4478 10424
rect 4478 10390 4512 10424
rect 4512 10390 4547 10424
rect 4547 10390 4581 10424
rect 4581 10390 4616 10424
rect 4616 10390 4650 10424
rect 4650 10390 4685 10424
rect 4685 10390 4719 10424
rect 4719 10390 4754 10424
rect 4754 10390 4788 10424
rect 4788 10390 4823 10424
rect 4823 10390 4857 10424
rect 4857 10390 4892 10424
rect 4892 10390 4926 10424
rect 4926 10390 4961 10424
rect 4961 10390 4995 10424
rect 4995 10390 5030 10424
rect 5030 10390 5064 10424
rect 5064 10390 5099 10424
rect 5099 10390 5133 10424
rect 5133 10390 5168 10424
rect 5168 10390 5202 10424
rect 5202 10390 5237 10424
rect 5237 10390 5271 10424
rect 5271 10390 5306 10424
rect 5306 10390 5340 10424
rect 5340 10390 5375 10424
rect 5375 10390 5409 10424
rect 5409 10390 5444 10424
rect 5444 10390 5478 10424
rect 5478 10390 5513 10424
rect 5513 10390 5547 10424
rect 5547 10390 5582 10424
rect 5582 10390 5616 10424
rect 5616 10390 5651 10424
rect 5651 10390 5685 10424
rect 5685 10397 5719 10424
rect 5719 10397 5753 10431
rect 5753 10397 5773 10431
rect 5685 10390 5773 10397
rect -48 10353 -14 10387
rect 25 10353 59 10387
rect 98 10353 132 10387
rect 171 10353 205 10387
rect 244 10353 278 10387
rect 317 10353 351 10387
rect 390 10353 424 10387
rect 463 10353 497 10387
rect 536 10353 570 10387
rect 609 10353 643 10387
rect 682 10353 716 10387
rect 755 10353 789 10387
rect 828 10353 862 10387
rect 901 10353 935 10387
rect 974 10353 1008 10387
rect 1047 10353 1081 10387
rect 1120 10353 1154 10387
rect 1193 10353 1227 10387
rect 1266 10353 1300 10387
rect 1339 10353 1373 10387
rect 1412 10353 1446 10387
rect 1485 10353 1519 10387
rect 1558 10353 1592 10387
rect 1631 10356 1665 10387
rect 1704 10356 1738 10387
rect 1777 10356 1811 10387
rect 1850 10356 1884 10387
rect 1923 10356 5773 10390
rect 1631 10353 1648 10356
rect 1648 10353 1665 10356
rect 1704 10353 1716 10356
rect 1716 10353 1738 10356
rect 1777 10353 1784 10356
rect 1784 10353 1811 10356
rect 1850 10353 1852 10356
rect 1852 10353 1884 10356
rect 1923 10353 1954 10356
rect 1954 10353 1988 10356
rect 1988 10353 2022 10356
rect 2022 10353 2057 10356
rect 2057 10353 2091 10356
rect 2091 10353 2126 10356
rect 2126 10353 2160 10356
rect 2160 10353 2195 10356
rect 2195 10353 2229 10356
rect 2229 10353 2264 10356
rect 2264 10353 2298 10356
rect 2298 10353 2333 10356
rect 2333 10353 2367 10356
rect 2367 10353 2402 10356
rect 2402 10353 2436 10356
rect 2436 10353 2471 10356
rect 2471 10353 2505 10356
rect 2505 10353 2540 10356
rect 2540 10353 2574 10356
rect 2574 10353 2609 10356
rect 2609 10353 2643 10356
rect 2643 10353 2678 10356
rect 2678 10353 2712 10356
rect 2712 10353 2747 10356
rect 2747 10353 2781 10356
rect 2781 10353 2816 10356
rect 2816 10353 2850 10356
rect 2850 10353 2885 10356
rect 2885 10353 2919 10356
rect 2919 10353 2954 10356
rect 2954 10353 2988 10356
rect 2988 10353 3023 10356
rect 3023 10353 3057 10356
rect 3057 10353 3092 10356
rect 3092 10353 3126 10356
rect 3126 10353 3161 10356
rect 3161 10353 3195 10356
rect 3195 10353 3230 10356
rect 3230 10353 3264 10356
rect 3264 10353 3299 10356
rect 3299 10353 3333 10356
rect 3333 10353 3368 10356
rect 3368 10353 3402 10356
rect 3402 10353 3437 10356
rect 3437 10353 3471 10356
rect 3471 10353 3506 10356
rect 3506 10353 3540 10356
rect 3540 10353 3575 10356
rect 3575 10353 3609 10356
rect 3609 10353 3644 10356
rect 3644 10353 3678 10356
rect 3678 10353 3713 10356
rect 3713 10353 3747 10356
rect 3747 10353 3782 10356
rect 3782 10353 3816 10356
rect 3816 10353 3851 10356
rect 3851 10353 3885 10356
rect 3885 10353 3920 10356
rect 3920 10353 3954 10356
rect 3954 10353 3989 10356
rect 3989 10353 4023 10356
rect 4023 10353 4058 10356
rect 4058 10353 4092 10356
rect 4092 10353 4127 10356
rect 4127 10353 4161 10356
rect 4161 10353 4196 10356
rect 4196 10353 4230 10356
rect 4230 10353 4265 10356
rect 4265 10353 4299 10356
rect 4299 10353 4334 10356
rect 4334 10353 4368 10356
rect 4368 10353 4403 10356
rect 4403 10353 4437 10356
rect 4437 10353 4472 10356
rect 4472 10353 4506 10356
rect 4506 10353 4541 10356
rect 4541 10353 4575 10356
rect 4575 10353 4610 10356
rect 4610 10353 4644 10356
rect 4644 10353 4679 10356
rect 4679 10353 4713 10356
rect 4713 10353 4748 10356
rect 4748 10353 4782 10356
rect 4782 10353 4817 10356
rect 4817 10353 4851 10356
rect 4851 10353 4886 10356
rect 4886 10353 4920 10356
rect 4920 10353 4955 10356
rect 4955 10353 4989 10356
rect 4989 10353 5024 10356
rect 5024 10353 5058 10356
rect 5058 10353 5093 10356
rect 5093 10353 5127 10356
rect 5127 10353 5162 10356
rect 5162 10353 5196 10356
rect 5196 10353 5231 10356
rect 5231 10353 5265 10356
rect 5265 10353 5300 10356
rect 5300 10353 5334 10356
rect 5334 10353 5369 10356
rect 5369 10353 5403 10356
rect 5403 10353 5438 10356
rect 5438 10353 5472 10356
rect 5472 10353 5507 10356
rect 5507 10353 5541 10356
rect 5541 10353 5576 10356
rect 5576 10353 5610 10356
rect 5610 10353 5645 10356
rect 5645 10353 5679 10356
rect 5679 10353 5714 10356
rect 5714 10353 5748 10356
rect 5748 10353 5773 10356
rect 14623 10213 14657 10247
rect 14695 10213 14729 10247
rect 14949 10213 14983 10247
rect 15021 10213 15055 10247
rect -17 10110 17 10144
rect 56 10110 90 10144
rect 129 10110 163 10144
rect 202 10110 236 10144
rect 275 10110 309 10144
rect 348 10110 382 10144
rect 421 10110 455 10144
rect 494 10110 528 10144
rect 567 10110 601 10144
rect 640 10110 674 10144
rect 713 10110 747 10144
rect 786 10110 820 10144
rect 859 10110 893 10144
rect 932 10110 966 10144
rect 1005 10110 1039 10144
rect 1078 10110 1112 10144
rect 1151 10110 1185 10144
rect 1224 10110 1258 10144
rect 1297 10110 1331 10144
rect 1370 10110 1404 10144
rect 1443 10110 1477 10144
rect 1516 10110 1550 10144
rect 1589 10110 1623 10144
rect 1662 10110 1696 10144
rect 1735 10110 1769 10144
rect 1808 10110 1842 10144
rect 1881 10110 1915 10144
rect 1954 10110 1988 10144
rect 2027 10110 2061 10144
rect 2100 10110 2134 10144
rect 2173 10110 2207 10144
rect 2246 10110 2280 10144
rect 2319 10110 2353 10144
rect 2392 10110 2426 10144
rect 2465 10110 2499 10144
rect 2538 10110 2572 10144
rect 2611 10110 2645 10144
rect 2684 10110 2718 10144
rect 2757 10110 2791 10144
rect 2830 10110 2864 10144
rect 2903 10110 2937 10144
rect 2976 10110 3010 10144
rect 3049 10110 3083 10144
rect 3122 10110 3156 10144
rect 3195 10110 3229 10144
rect 3268 10110 3302 10144
rect 3341 10110 3375 10144
rect 3414 10110 3448 10144
rect 3487 10110 3521 10144
rect 3560 10110 3594 10144
rect 3633 10110 3667 10144
rect 3706 10110 3740 10144
rect 3779 10110 3813 10144
rect 3852 10110 3886 10144
rect 3925 10110 3959 10144
rect 3998 10110 4032 10144
rect 4071 10110 4105 10144
rect 4144 10110 4178 10144
rect 4216 10110 4250 10144
rect 4288 10110 4322 10144
rect 4360 10110 4394 10144
rect 4432 10110 4466 10144
rect 4504 10110 4538 10144
rect 4576 10110 4610 10144
rect 4648 10110 4682 10144
rect 4720 10110 4754 10144
rect 4792 10110 4826 10144
rect 4864 10110 4898 10144
rect 4936 10110 4970 10144
rect 5008 10110 5042 10144
rect 5080 10110 5114 10144
rect 5152 10110 5186 10144
rect 5224 10110 5258 10144
rect 5296 10110 5330 10144
rect 5368 10110 5402 10144
rect 5440 10110 5474 10144
rect 5512 10110 5546 10144
rect 5584 10110 5618 10144
rect 5656 10110 5690 10144
rect 5728 10110 5762 10144
rect 5800 10110 5834 10144
rect 5872 10110 5906 10144
rect 5944 10110 5978 10144
rect 6016 10110 6050 10144
rect 6088 10110 6122 10144
rect 6160 10110 6194 10144
rect 6232 10110 6266 10144
rect 6304 10110 6338 10144
rect 6376 10110 6410 10144
rect 6448 10110 6482 10144
rect 6520 10110 6554 10144
rect 6592 10110 6626 10144
rect 6664 10110 6698 10144
rect 6736 10110 6770 10144
rect 6808 10110 6842 10144
rect 6880 10110 6914 10144
rect 6952 10110 6986 10144
rect 7024 10110 7058 10144
rect 7096 10110 7130 10144
rect 7168 10110 7202 10144
rect 7240 10110 7274 10144
rect 7312 10110 7346 10144
rect 7384 10110 7418 10144
rect 7456 10110 7490 10144
rect 7528 10110 7562 10144
rect 7600 10110 7634 10144
rect 7672 10110 7706 10144
rect 7744 10110 7778 10144
rect 7816 10110 7850 10144
rect 7888 10110 7922 10144
rect 7960 10110 7994 10144
rect 8032 10110 8066 10144
rect 8104 10110 8138 10144
rect 8176 10110 8210 10144
rect 8248 10110 8282 10144
rect 8320 10110 8354 10144
rect 8392 10110 8426 10144
rect 8464 10110 8498 10144
rect 8536 10110 8570 10144
rect 8608 10110 8642 10144
rect 8680 10110 8714 10144
rect 8752 10110 8786 10144
rect 8824 10110 8858 10144
rect 8896 10110 8930 10144
rect 8968 10110 9002 10144
rect 9040 10110 9074 10144
rect 9112 10110 9146 10144
rect 9184 10110 9218 10144
rect 9256 10110 9290 10144
rect 9328 10110 9362 10144
rect 9400 10110 9434 10144
rect 9472 10110 9506 10144
rect 9544 10110 9578 10144
rect 9616 10110 9650 10144
rect 9688 10110 9722 10144
rect 9760 10110 9794 10144
rect 9832 10110 9866 10144
rect 9904 10110 9938 10144
rect 9976 10110 10010 10144
rect 10048 10110 10082 10144
rect 10120 10110 10154 10144
rect 10192 10110 10226 10144
rect 10264 10110 10298 10144
rect 10336 10110 10370 10144
rect 10408 10110 10442 10144
rect 10480 10110 10514 10144
rect 10552 10110 10586 10144
rect 10624 10110 10658 10144
rect 10696 10110 10730 10144
rect 10768 10110 10802 10144
rect 10840 10110 10874 10144
rect 10912 10110 10946 10144
rect 10984 10110 11018 10144
rect 11056 10110 11090 10144
rect 11128 10110 11162 10144
rect 11200 10110 11234 10144
rect 11272 10110 11306 10144
rect 11344 10110 11378 10144
rect 11416 10110 11450 10144
rect 11488 10110 11522 10144
rect 11560 10110 11594 10144
rect 11632 10110 11666 10144
rect 11704 10110 11738 10144
rect 11776 10110 11810 10144
rect 11848 10110 11882 10144
rect 11920 10110 11954 10144
rect 11992 10110 12026 10144
rect 12064 10110 12098 10144
rect 12136 10110 12170 10144
rect 12208 10141 12242 10144
rect 12280 10141 12314 10144
rect 12352 10141 12386 10144
rect 12424 10141 12458 10144
rect 12496 10141 12530 10144
rect 12568 10141 12602 10144
rect 12640 10141 12674 10144
rect 12712 10141 12746 10144
rect 12946 10141 12980 10144
rect 13020 10141 13054 10144
rect 13093 10141 13127 10144
rect 13166 10141 13200 10144
rect 13239 10141 13273 10144
rect 13312 10141 13346 10144
rect 13385 10141 13419 10144
rect 13458 10141 13492 10144
rect 13531 10141 13565 10144
rect 13604 10141 13638 10144
rect 13677 10141 13711 10144
rect 13750 10141 13784 10144
rect 13823 10141 13857 10144
rect 13896 10141 13930 10144
rect 13969 10141 14003 10144
rect 14042 10141 14076 10144
rect 14115 10141 14149 10144
rect 14188 10141 14222 10144
rect 14261 10141 14295 10144
rect 14334 10141 14368 10144
rect 14407 10141 14441 10144
rect 14480 10141 14514 10144
rect 14553 10141 14587 10144
rect 14956 10141 14990 10144
rect 15042 10141 15076 10144
rect 15128 10141 15162 10144
rect 15214 10141 15248 10144
rect 12208 10110 12225 10141
rect 12225 10110 12242 10141
rect 12280 10110 12295 10141
rect 12295 10110 12314 10141
rect 12352 10110 12365 10141
rect 12365 10110 12386 10141
rect 12424 10110 12435 10141
rect 12435 10110 12458 10141
rect 12496 10110 12504 10141
rect 12504 10110 12530 10141
rect 12568 10110 12573 10141
rect 12573 10110 12602 10141
rect 12640 10110 12642 10141
rect 12642 10110 12674 10141
rect 12712 10110 12745 10141
rect 12745 10110 12746 10141
rect 12946 10110 12952 10141
rect 12952 10110 12980 10141
rect 13020 10110 13021 10141
rect 13021 10110 13054 10141
rect 13093 10110 13125 10141
rect 13125 10110 13127 10141
rect 13166 10110 13194 10141
rect 13194 10110 13200 10141
rect 13239 10110 13263 10141
rect 13263 10110 13273 10141
rect 13312 10110 13332 10141
rect 13332 10110 13346 10141
rect 13385 10110 13401 10141
rect 13401 10110 13419 10141
rect 13458 10110 13470 10141
rect 13470 10110 13492 10141
rect 13531 10110 13539 10141
rect 13539 10110 13565 10141
rect 13604 10110 13608 10141
rect 13608 10110 13638 10141
rect 13677 10110 13711 10141
rect 13750 10110 13780 10141
rect 13780 10110 13784 10141
rect 13823 10110 13849 10141
rect 13849 10110 13857 10141
rect 13896 10110 13918 10141
rect 13918 10110 13930 10141
rect 13969 10110 13987 10141
rect 13987 10110 14003 10141
rect 14042 10110 14056 10141
rect 14056 10110 14076 10141
rect 14115 10110 14125 10141
rect 14125 10110 14149 10141
rect 14188 10110 14194 10141
rect 14194 10110 14222 10141
rect 14261 10110 14263 10141
rect 14263 10110 14295 10141
rect 14334 10110 14367 10141
rect 14367 10110 14368 10141
rect 14407 10110 14436 10141
rect 14436 10110 14441 10141
rect 14480 10110 14505 10141
rect 14505 10110 14514 10141
rect 14553 10110 14574 10141
rect 14574 10110 14587 10141
rect 14956 10110 14988 10141
rect 14988 10110 14990 10141
rect 15042 10110 15057 10141
rect 15057 10110 15076 10141
rect 15128 10110 15160 10141
rect 15160 10110 15162 10141
rect 15214 10110 15229 10141
rect 15229 10110 15248 10141
rect 15299 10110 15333 10144
rect -17 10038 17 10072
rect 15299 10038 15333 10072
rect -17 9959 17 9993
rect 14658 10001 14692 10035
rect 14658 9929 14692 9963
rect 14824 9972 14858 10006
rect 14926 9972 14960 10006
rect 15299 9969 15333 9993
rect 15299 9959 15333 9969
rect -17 9881 17 9915
rect 15299 9900 15333 9915
rect 15299 9881 15333 9900
rect 4110 9787 4144 9821
rect 4110 9715 4144 9749
rect 4422 9787 4456 9821
rect 4422 9715 4456 9749
rect 4912 9787 4946 9821
rect 4912 9715 4946 9749
rect 5264 9787 5298 9821
rect 5264 9715 5298 9749
rect 6410 9787 6444 9821
rect 6410 9715 6444 9749
rect 6762 9787 6796 9821
rect 6762 9715 6796 9749
rect 7134 9787 7168 9821
rect 7134 9715 7168 9749
rect 7486 9787 7520 9821
rect 7486 9715 7520 9749
rect 14553 5974 14587 6008
rect 11424 5916 11458 5950
rect 14553 5902 14587 5936
rect 11424 5844 11458 5878
rect 15170 5130 15204 5164
rect 15247 5130 15281 5164
rect 15324 5130 15358 5164
rect 15400 5130 15434 5164
rect 15476 5130 15510 5164
rect 15552 5131 15578 5164
rect 15578 5131 15586 5164
rect 15628 5131 15646 5164
rect 15646 5131 15662 5164
rect 15704 5131 15714 5164
rect 15714 5131 15738 5164
rect 15552 5130 15586 5131
rect 15628 5130 15662 5131
rect 15704 5130 15738 5131
rect 15780 5130 15814 5164
rect 15856 5130 15890 5164
rect 15932 5130 15966 5164
rect 16008 5130 16042 5164
rect 15170 5058 15204 5092
rect 15247 5058 15281 5092
rect 15324 5058 15358 5092
rect 15400 5058 15434 5092
rect 15476 5058 15510 5092
rect 15552 5058 15586 5092
rect 15628 5058 15662 5092
rect 15704 5058 15738 5092
rect 15780 5058 15814 5092
rect 15856 5058 15890 5092
rect 15932 5058 15966 5092
rect 16008 5058 16042 5092
rect 15170 4986 15204 5020
rect 15247 4986 15281 5020
rect 15324 4986 15358 5020
rect 15400 4986 15434 5020
rect 15476 4986 15510 5020
rect 15552 4986 15586 5020
rect 15628 4986 15662 5020
rect 15704 4986 15738 5020
rect 15780 4986 15814 5020
rect 15856 4986 15890 5020
rect 15932 4986 15966 5020
rect 16008 4986 16042 5020
rect 11633 3617 11667 3651
rect 11633 3545 11667 3579
rect 12407 2423 12441 2457
rect 12488 2423 12522 2457
rect 12569 2423 12603 2457
rect 12649 2423 12683 2457
rect 12729 2423 12763 2457
rect 12809 2423 12843 2457
rect 7552 2368 7586 2402
rect 7624 2368 7658 2402
rect 11952 2373 11986 2407
rect 12024 2373 12058 2407
<< metal1 >>
rect 1948 13606 2618 13618
rect 1948 13572 1954 13606
rect 1988 13572 2032 13606
rect 2066 13600 2110 13606
rect 2144 13600 2188 13606
rect 2222 13600 2266 13606
rect 2300 13600 2344 13606
rect 2378 13600 2422 13606
rect 2456 13600 2500 13606
rect 2534 13600 2578 13606
rect 2066 13572 2080 13600
rect 2144 13572 2146 13600
rect 2264 13572 2266 13600
rect 1948 13548 2080 13572
rect 2132 13548 2146 13572
rect 2198 13548 2212 13572
rect 2264 13548 2278 13572
rect 2330 13548 2344 13600
rect 2396 13548 2410 13600
rect 2462 13548 2476 13600
rect 2534 13572 2542 13600
rect 2612 13572 2618 13606
rect 2528 13548 2542 13572
rect 2594 13548 2618 13572
rect 1948 13536 2618 13548
rect 1948 13532 2080 13536
rect 2132 13532 2146 13536
rect 2198 13532 2212 13536
rect 2264 13532 2278 13536
rect 1948 13498 1954 13532
rect 1988 13498 2032 13532
rect 2066 13498 2080 13532
rect 2144 13498 2146 13532
rect 2264 13498 2266 13532
rect 1948 13484 2080 13498
rect 2132 13484 2146 13498
rect 2198 13484 2212 13498
rect 2264 13484 2278 13498
rect 2330 13484 2344 13536
rect 2396 13484 2410 13536
rect 2462 13484 2476 13536
rect 2528 13532 2542 13536
rect 2594 13532 2618 13536
rect 2534 13498 2542 13532
rect 2612 13498 2618 13532
rect 2528 13484 2542 13498
rect 2594 13484 2618 13498
rect 1948 13472 2618 13484
rect 1948 13458 2080 13472
rect 2132 13458 2146 13472
rect 2198 13458 2212 13472
rect 2264 13458 2278 13472
rect 1948 13424 1954 13458
rect 1988 13424 2032 13458
rect 2066 13424 2080 13458
rect 2144 13424 2146 13458
rect 2264 13424 2266 13458
rect 1948 13420 2080 13424
rect 2132 13420 2146 13424
rect 2198 13420 2212 13424
rect 2264 13420 2278 13424
rect 2330 13420 2344 13472
rect 2396 13420 2410 13472
rect 2462 13420 2476 13472
rect 2528 13458 2542 13472
rect 2594 13458 2618 13472
rect 2534 13424 2542 13458
rect 2612 13424 2618 13458
rect 2528 13420 2542 13424
rect 2594 13420 2618 13424
rect 1948 13408 2618 13420
rect 1948 13383 2080 13408
rect 2132 13383 2146 13408
rect 2198 13383 2212 13408
rect 2264 13383 2278 13408
rect 1948 13349 1954 13383
rect 1988 13349 2032 13383
rect 2066 13356 2080 13383
rect 2144 13356 2146 13383
rect 2264 13356 2266 13383
rect 2330 13356 2344 13408
rect 2396 13356 2410 13408
rect 2462 13356 2476 13408
rect 2528 13383 2542 13408
rect 2594 13383 2618 13408
rect 2534 13356 2542 13383
rect 2066 13349 2110 13356
rect 2144 13349 2188 13356
rect 2222 13349 2266 13356
rect 2300 13349 2344 13356
rect 2378 13349 2422 13356
rect 2456 13349 2500 13356
rect 2534 13349 2578 13356
rect 2612 13349 2618 13383
rect 1948 13344 2618 13349
rect 1948 13308 2080 13344
rect 2132 13308 2146 13344
rect 2198 13308 2212 13344
rect 2264 13308 2278 13344
rect 1948 13274 1954 13308
rect 1988 13274 2032 13308
rect 2066 13292 2080 13308
rect 2144 13292 2146 13308
rect 2264 13292 2266 13308
rect 2330 13292 2344 13344
rect 2396 13292 2410 13344
rect 2462 13292 2476 13344
rect 2528 13308 2542 13344
rect 2594 13308 2618 13344
rect 2534 13292 2542 13308
rect 2066 13280 2110 13292
rect 2144 13280 2188 13292
rect 2222 13280 2266 13292
rect 2300 13280 2344 13292
rect 2378 13280 2422 13292
rect 2456 13280 2500 13292
rect 2534 13280 2578 13292
rect 2066 13274 2080 13280
rect 2144 13274 2146 13280
rect 2264 13274 2266 13280
rect 1948 13233 2080 13274
rect 2132 13233 2146 13274
rect 2198 13233 2212 13274
rect 2264 13233 2278 13274
rect 1948 13199 1954 13233
rect 1988 13199 2032 13233
rect 2066 13228 2080 13233
rect 2144 13228 2146 13233
rect 2264 13228 2266 13233
rect 2330 13228 2344 13280
rect 2396 13228 2410 13280
rect 2462 13228 2476 13280
rect 2534 13274 2542 13280
rect 2612 13274 2618 13308
rect 2528 13233 2542 13274
rect 2594 13233 2618 13274
rect 2534 13228 2542 13233
rect 2066 13215 2110 13228
rect 2144 13215 2188 13228
rect 2222 13215 2266 13228
rect 2300 13215 2344 13228
rect 2378 13215 2422 13228
rect 2456 13215 2500 13228
rect 2534 13215 2578 13228
rect 2066 13199 2080 13215
rect 2144 13199 2146 13215
rect 2264 13199 2266 13215
rect 1948 13163 2080 13199
rect 2132 13163 2146 13199
rect 2198 13163 2212 13199
rect 2264 13163 2278 13199
rect 2330 13163 2344 13215
rect 2396 13163 2410 13215
rect 2462 13163 2476 13215
rect 2534 13199 2542 13215
rect 2612 13199 2618 13233
rect 2528 13163 2542 13199
rect 2594 13163 2618 13199
rect 1948 13158 2618 13163
rect 1948 13124 1954 13158
rect 1988 13124 2032 13158
rect 2066 13150 2110 13158
rect 2144 13150 2188 13158
rect 2222 13150 2266 13158
rect 2300 13150 2344 13158
rect 2378 13150 2422 13158
rect 2456 13150 2500 13158
rect 2534 13150 2578 13158
rect 2066 13124 2080 13150
rect 2144 13124 2146 13150
rect 2264 13124 2266 13150
rect 1948 13098 2080 13124
rect 2132 13098 2146 13124
rect 2198 13098 2212 13124
rect 2264 13098 2278 13124
rect 2330 13098 2344 13150
rect 2396 13098 2410 13150
rect 2462 13098 2476 13150
rect 2534 13124 2542 13150
rect 2612 13124 2618 13158
rect 2528 13098 2542 13124
rect 2594 13098 2618 13124
rect 1948 13085 2618 13098
rect 1948 13083 2080 13085
rect 2132 13083 2146 13085
rect 2198 13083 2212 13085
rect 2264 13083 2278 13085
rect 1948 13049 1954 13083
rect 1988 13049 2032 13083
rect 2066 13049 2080 13083
rect 2144 13049 2146 13083
rect 2264 13049 2266 13083
rect 1948 13033 2080 13049
rect 2132 13033 2146 13049
rect 2198 13033 2212 13049
rect 2264 13033 2278 13049
rect 2330 13033 2344 13085
rect 2396 13033 2410 13085
rect 2462 13033 2476 13085
rect 2528 13083 2542 13085
rect 2594 13083 2618 13085
rect 2534 13049 2542 13083
rect 2612 13049 2618 13083
rect 2528 13033 2542 13049
rect 2594 13033 2618 13049
rect 1948 13020 2618 13033
rect 1948 13008 2080 13020
rect 2132 13008 2146 13020
rect 2198 13008 2212 13020
rect 2264 13008 2278 13020
rect 1948 12974 1954 13008
rect 1988 12974 2032 13008
rect 2066 12974 2080 13008
rect 2144 12974 2146 13008
rect 2264 12974 2266 13008
rect 1948 12968 2080 12974
rect 2132 12968 2146 12974
rect 2198 12968 2212 12974
rect 2264 12968 2278 12974
rect 2330 12968 2344 13020
rect 2396 12968 2410 13020
rect 2462 12968 2476 13020
rect 2528 13008 2542 13020
rect 2594 13008 2618 13020
rect 2534 12974 2542 13008
rect 2612 12974 2618 13008
rect 2528 12968 2542 12974
rect 2594 12968 2618 12974
rect 1948 12955 2618 12968
rect 1948 12933 2080 12955
rect 2132 12933 2146 12955
rect 2198 12933 2212 12955
rect 2264 12933 2278 12955
rect 1948 12899 1954 12933
rect 1988 12899 2032 12933
rect 2066 12903 2080 12933
rect 2144 12903 2146 12933
rect 2264 12903 2266 12933
rect 2330 12903 2344 12955
rect 2396 12903 2410 12955
rect 2462 12903 2476 12955
rect 2528 12933 2542 12955
rect 2594 12933 2618 12955
rect 2534 12903 2542 12933
rect 2066 12899 2110 12903
rect 2144 12899 2188 12903
rect 2222 12899 2266 12903
rect 2300 12899 2344 12903
rect 2378 12899 2422 12903
rect 2456 12899 2500 12903
rect 2534 12899 2578 12903
rect 2612 12899 2618 12933
rect 1948 12887 2618 12899
rect 1922 12368 4269 12373
rect 1922 12364 2066 12368
rect 1922 12330 1934 12364
rect 1968 12330 2008 12364
rect 2042 12330 2066 12364
rect 1922 12316 2066 12330
rect 2118 12316 2131 12368
rect 2183 12364 2196 12368
rect 2248 12364 2261 12368
rect 2313 12364 2326 12368
rect 2378 12364 2390 12368
rect 2442 12364 2454 12368
rect 2190 12330 2196 12364
rect 2442 12330 2452 12364
rect 2183 12316 2196 12330
rect 2248 12316 2261 12330
rect 2313 12316 2326 12330
rect 2378 12316 2390 12330
rect 2442 12316 2454 12330
rect 2506 12316 2518 12368
rect 2570 12316 2582 12368
rect 2634 12364 4269 12368
rect 2634 12330 2674 12364
rect 2708 12330 2748 12364
rect 2782 12330 2822 12364
rect 2856 12330 2896 12364
rect 2930 12330 2970 12364
rect 3004 12330 3044 12364
rect 3078 12330 3118 12364
rect 3152 12330 3192 12364
rect 3226 12330 3266 12364
rect 3300 12330 3340 12364
rect 3374 12330 3414 12364
rect 3448 12330 3488 12364
rect 3522 12330 3562 12364
rect 3596 12330 3636 12364
rect 3670 12330 3710 12364
rect 3744 12330 3784 12364
rect 3818 12330 3858 12364
rect 3892 12330 3931 12364
rect 3965 12330 4004 12364
rect 4038 12363 4077 12364
rect 4111 12363 4150 12364
rect 4184 12363 4223 12364
rect 4257 12363 4269 12364
rect 4038 12330 4041 12363
rect 4111 12330 4127 12363
rect 4184 12330 4213 12363
rect 2634 12316 4041 12330
rect 1922 12311 4041 12316
rect 4093 12311 4127 12330
rect 4179 12311 4213 12330
rect 4265 12311 4269 12363
rect 1922 12282 4269 12311
tri 1895 12248 1922 12275 se
rect 1922 12248 1934 12282
rect 1968 12248 2008 12282
rect 2042 12254 2082 12282
rect 2116 12254 2156 12282
rect 2190 12254 2230 12282
rect 2264 12254 2304 12282
rect 2338 12254 2378 12282
rect 2412 12254 2452 12282
rect 2486 12254 2526 12282
rect 2560 12254 2600 12282
rect 2042 12248 2066 12254
rect -2923 12237 319 12248
tri 1894 12247 1895 12248 se
rect 1895 12247 2066 12248
rect -2923 12203 -2911 12237
rect -2877 12203 -2838 12237
rect -2804 12203 -2765 12237
rect -2731 12203 -2692 12237
rect -2658 12203 -2619 12237
rect -2585 12203 -2546 12237
rect -2512 12203 -2473 12237
rect -2439 12203 -2400 12237
rect -2366 12203 -2327 12237
rect -2293 12203 -2254 12237
rect -2220 12203 -2181 12237
rect -2147 12203 -2108 12237
rect -2074 12203 -2035 12237
rect -2001 12203 -1962 12237
rect -1928 12203 -1889 12237
rect -1855 12203 -1816 12237
rect -1782 12203 -1743 12237
rect -2923 12165 -1743 12203
rect -2923 12131 -2911 12165
rect -2877 12131 -2838 12165
rect -2804 12131 -2765 12165
rect -2731 12131 -2692 12165
rect -2658 12131 -2619 12165
rect -2585 12131 -2546 12165
rect -2512 12131 -2473 12165
rect -2439 12131 -2400 12165
rect -2366 12131 -2327 12165
rect -2293 12131 -2254 12165
rect -2220 12131 -2181 12165
rect -2147 12131 -2108 12165
rect -2074 12131 -2035 12165
rect -2001 12131 -1962 12165
rect -1928 12131 -1889 12165
rect -1855 12131 -1816 12165
rect -1782 12131 -1743 12165
rect -2923 12093 -1743 12131
rect -2923 12059 -2911 12093
rect -2877 12059 -2838 12093
rect -2804 12059 -2765 12093
rect -2731 12059 -2692 12093
rect -2658 12059 -2619 12093
rect -2585 12059 -2546 12093
rect -2512 12059 -2473 12093
rect -2439 12059 -2400 12093
rect -2366 12059 -2327 12093
rect -2293 12059 -2254 12093
rect -2220 12059 -2181 12093
rect -2147 12059 -2108 12093
rect -2074 12059 -2035 12093
rect -2001 12059 -1962 12093
rect -1928 12059 -1889 12093
rect -1855 12059 -1816 12093
rect -1782 12059 -1743 12093
rect -2923 12021 -1743 12059
rect -2923 11987 -2911 12021
rect -2877 11987 -2838 12021
rect -2804 11987 -2765 12021
rect -2731 11987 -2692 12021
rect -2658 11987 -2619 12021
rect -2585 11987 -2546 12021
rect -2512 11987 -2473 12021
rect -2439 11987 -2400 12021
rect -2366 11987 -2327 12021
rect -2293 11987 -2254 12021
rect -2220 11987 -2181 12021
rect -2147 11987 -2108 12021
rect -2074 11987 -2035 12021
rect -2001 11987 -1962 12021
rect -1928 11987 -1889 12021
rect -1855 11987 -1816 12021
rect -1782 11987 -1743 12021
rect -2923 11949 -1743 11987
rect -2923 11915 -2911 11949
rect -2877 11915 -2838 11949
rect -2804 11915 -2765 11949
rect -2731 11915 -2692 11949
rect -2658 11915 -2619 11949
rect -2585 11915 -2546 11949
rect -2512 11915 -2473 11949
rect -2439 11915 -2400 11949
rect -2366 11915 -2327 11949
rect -2293 11915 -2254 11949
rect -2220 11915 -2181 11949
rect -2147 11915 -2108 11949
rect -2074 11915 -2035 11949
rect -2001 11915 -1962 11949
rect -1928 11915 -1889 11949
rect -1855 11915 -1816 11949
rect -1782 11915 -1743 11949
rect -2923 11877 -1743 11915
rect -2923 11843 -2911 11877
rect -2877 11843 -2838 11877
rect -2804 11843 -2765 11877
rect -2731 11843 -2692 11877
rect -2658 11843 -2619 11877
rect -2585 11843 -2546 11877
rect -2512 11843 -2473 11877
rect -2439 11843 -2400 11877
rect -2366 11843 -2327 11877
rect -2293 11843 -2254 11877
rect -2220 11843 -2181 11877
rect -2147 11843 -2108 11877
rect -2074 11843 -2035 11877
rect -2001 11843 -1962 11877
rect -1928 11843 -1889 11877
rect -1855 11843 -1816 11877
rect -1782 11843 -1743 11877
rect -2923 11805 -1743 11843
rect -2923 11771 -2911 11805
rect -2877 11771 -2838 11805
rect -2804 11771 -2765 11805
rect -2731 11771 -2692 11805
rect -2658 11771 -2619 11805
rect -2585 11771 -2546 11805
rect -2512 11771 -2473 11805
rect -2439 11771 -2400 11805
rect -2366 11771 -2327 11805
rect -2293 11771 -2254 11805
rect -2220 11771 -2181 11805
rect -2147 11771 -2108 11805
rect -2074 11771 -2035 11805
rect -2001 11771 -1962 11805
rect -1928 11771 -1889 11805
rect -1855 11771 -1816 11805
rect -1782 11771 -1743 11805
rect 307 12202 319 12237
tri 319 12202 364 12247 sw
tri 1849 12202 1894 12247 se
rect 1894 12202 2066 12247
rect 2118 12202 2131 12254
rect 2190 12248 2196 12254
rect 2442 12248 2452 12254
rect 2183 12202 2196 12248
rect 2248 12202 2261 12248
rect 2313 12202 2326 12248
rect 2378 12202 2390 12248
rect 2442 12202 2454 12248
rect 2506 12202 2518 12254
rect 2570 12202 2582 12254
rect 2634 12248 2674 12282
rect 2708 12248 2748 12282
rect 2782 12248 2822 12282
rect 2856 12248 2896 12282
rect 2930 12248 2970 12282
rect 3004 12248 3044 12282
rect 3078 12248 3118 12282
rect 3152 12248 3192 12282
rect 3226 12248 3266 12282
rect 3300 12248 3340 12282
rect 3374 12248 3414 12282
rect 3448 12248 3488 12282
rect 3522 12248 3562 12282
rect 3596 12248 3636 12282
rect 3670 12248 3710 12282
rect 3744 12248 3784 12282
rect 3818 12248 3858 12282
rect 3892 12248 3931 12282
rect 3965 12248 4004 12282
rect 4038 12261 4077 12282
rect 4111 12261 4150 12282
rect 4184 12261 4223 12282
rect 4257 12261 4269 12282
rect 4038 12248 4041 12261
rect 4111 12248 4127 12261
rect 4184 12248 4213 12261
rect 2634 12209 4041 12248
rect 4093 12209 4127 12248
rect 4179 12209 4213 12248
rect 4265 12209 4269 12261
rect 2634 12202 4269 12209
rect 307 12200 364 12202
tri 364 12200 366 12202 sw
tri 1847 12200 1849 12202 se
rect 1849 12200 4269 12202
rect 307 12166 366 12200
tri 366 12166 400 12200 sw
tri 1813 12166 1847 12200 se
rect 1847 12166 1934 12200
rect 1968 12166 2008 12200
rect 2042 12166 2082 12200
rect 2116 12166 2156 12200
rect 2190 12166 2230 12200
rect 2264 12166 2304 12200
rect 2338 12166 2378 12200
rect 2412 12166 2452 12200
rect 2486 12166 2526 12200
rect 2560 12166 2600 12200
rect 2634 12166 2674 12200
rect 2708 12166 2748 12200
rect 2782 12166 2822 12200
rect 2856 12166 2896 12200
rect 2930 12166 2970 12200
rect 3004 12166 3044 12200
rect 3078 12166 3118 12200
rect 3152 12166 3192 12200
rect 3226 12166 3266 12200
rect 3300 12166 3340 12200
rect 3374 12166 3414 12200
rect 3448 12166 3488 12200
rect 3522 12166 3562 12200
rect 3596 12166 3636 12200
rect 3670 12166 3710 12200
rect 3744 12166 3784 12200
rect 3818 12166 3858 12200
rect 3892 12166 3931 12200
rect 3965 12166 4004 12200
rect 4038 12166 4077 12200
rect 4111 12166 4150 12200
rect 4184 12166 4223 12200
rect 4257 12166 4269 12200
rect 307 12118 400 12166
tri 400 12118 448 12166 sw
tri 1765 12118 1813 12166 se
rect 1813 12159 4269 12166
rect 1813 12118 4041 12159
rect 4093 12118 4127 12159
rect 4179 12118 4213 12159
rect 307 12084 448 12118
tri 448 12084 482 12118 sw
tri 1731 12084 1765 12118 se
rect 1765 12084 1934 12118
rect 1968 12084 2008 12118
rect 2042 12084 2082 12118
rect 2116 12084 2156 12118
rect 2190 12084 2230 12118
rect 2264 12084 2304 12118
rect 2338 12084 2378 12118
rect 2412 12084 2452 12118
rect 2486 12084 2526 12118
rect 2560 12084 2600 12118
rect 2634 12084 2674 12118
rect 2708 12084 2748 12118
rect 2782 12084 2822 12118
rect 2856 12084 2896 12118
rect 2930 12084 2970 12118
rect 3004 12084 3044 12118
rect 3078 12084 3118 12118
rect 3152 12084 3192 12118
rect 3226 12084 3266 12118
rect 3300 12084 3340 12118
rect 3374 12084 3414 12118
rect 3448 12084 3488 12118
rect 3522 12084 3562 12118
rect 3596 12084 3636 12118
rect 3670 12084 3710 12118
rect 3744 12084 3784 12118
rect 3818 12084 3858 12118
rect 3892 12084 3931 12118
rect 3965 12084 4004 12118
rect 4038 12107 4041 12118
rect 4111 12107 4127 12118
rect 4184 12107 4213 12118
rect 4265 12107 4269 12159
rect 4038 12084 4077 12107
rect 4111 12084 4150 12107
rect 4184 12084 4223 12107
rect 4257 12084 4269 12107
rect 307 12036 482 12084
tri 482 12036 530 12084 sw
tri 1683 12036 1731 12084 se
rect 1731 12056 4269 12084
rect 1731 12036 4041 12056
rect 4093 12036 4127 12056
rect 4179 12036 4213 12056
rect 307 12002 530 12036
tri 530 12002 564 12036 sw
tri 1649 12002 1683 12036 se
rect 1683 12002 1934 12036
rect 1968 12002 2008 12036
rect 2042 12002 2082 12036
rect 2116 12002 2156 12036
rect 2190 12002 2230 12036
rect 2264 12002 2304 12036
rect 2338 12002 2378 12036
rect 2412 12002 2452 12036
rect 2486 12002 2526 12036
rect 2560 12002 2600 12036
rect 2634 12002 2674 12036
rect 2708 12002 2748 12036
rect 2782 12002 2822 12036
rect 2856 12002 2896 12036
rect 2930 12002 2970 12036
rect 3004 12002 3044 12036
rect 3078 12002 3118 12036
rect 3152 12002 3192 12036
rect 3226 12002 3266 12036
rect 3300 12002 3340 12036
rect 3374 12002 3414 12036
rect 3448 12002 3488 12036
rect 3522 12002 3562 12036
rect 3596 12002 3636 12036
rect 3670 12002 3710 12036
rect 3744 12002 3784 12036
rect 3818 12002 3858 12036
rect 3892 12002 3931 12036
rect 3965 12002 4004 12036
rect 4038 12004 4041 12036
rect 4111 12004 4127 12036
rect 4184 12004 4213 12036
rect 4265 12004 4269 12056
rect 4038 12002 4077 12004
rect 4111 12002 4150 12004
rect 4184 12002 4223 12004
rect 4257 12002 4269 12004
rect 307 11998 564 12002
tri 564 11998 568 12002 sw
tri 1645 11998 1649 12002 se
rect 1649 11998 4269 12002
rect 307 11982 568 11998
tri 568 11982 584 11998 sw
tri 1629 11982 1645 11998 se
rect 1645 11993 4269 11998
rect 1645 11982 1932 11993
tri 1932 11982 1943 11993 nw
rect 307 11976 1729 11982
rect 307 11942 367 11976
rect 401 11942 441 11976
rect 475 11942 515 11976
rect 549 11942 588 11976
rect 622 11942 661 11976
rect 695 11942 734 11976
rect 768 11942 807 11976
rect 841 11942 880 11976
rect 914 11942 953 11976
rect 987 11942 1026 11976
rect 1060 11942 1099 11976
rect 1133 11942 1172 11976
rect 1206 11942 1245 11976
rect 1279 11942 1318 11976
rect 1352 11942 1391 11976
rect 1425 11942 1464 11976
rect 1498 11942 1537 11976
rect 1571 11942 1610 11976
rect 1644 11942 1683 11976
rect 1717 11942 1729 11976
rect 307 11888 1729 11942
rect 307 11854 367 11888
rect 401 11854 441 11888
rect 475 11854 515 11888
rect 549 11854 588 11888
rect 622 11854 661 11888
rect 695 11854 734 11888
rect 768 11854 807 11888
rect 841 11854 880 11888
rect 914 11854 953 11888
rect 987 11854 1026 11888
rect 1060 11854 1099 11888
rect 1133 11854 1172 11888
rect 1206 11854 1245 11888
rect 1279 11854 1318 11888
rect 1352 11854 1391 11888
rect 1425 11854 1464 11888
rect 1498 11854 1537 11888
rect 1571 11854 1610 11888
rect 1644 11854 1683 11888
rect 1717 11854 1729 11888
rect 307 11800 1729 11854
rect 307 11771 367 11800
rect -2923 11766 367 11771
rect 401 11766 441 11800
rect 475 11766 515 11800
rect 549 11766 588 11800
rect 622 11766 661 11800
rect 695 11766 734 11800
rect 768 11766 807 11800
rect 841 11766 880 11800
rect 914 11766 953 11800
rect 987 11766 1026 11800
rect 1060 11766 1099 11800
rect 1133 11766 1172 11800
rect 1206 11766 1245 11800
rect 1279 11766 1318 11800
rect 1352 11766 1391 11800
rect 1425 11766 1464 11800
rect 1498 11766 1537 11800
rect 1571 11766 1610 11800
rect 1644 11766 1683 11800
rect 1717 11766 1729 11800
tri 1729 11779 1932 11982 nw
rect -2923 11760 1729 11766
tri 13720 10870 13757 10907 se
tri 13894 10870 13925 10901 nw
tri 13805 10818 13806 10819 nw
rect 2913 10780 16806 10786
rect 2965 10734 16754 10780
rect 2965 10728 2978 10734
rect 2913 10722 2978 10728
tri 2978 10722 2990 10734 nw
tri 16729 10722 16741 10734 ne
rect 16741 10728 16754 10734
rect 16741 10722 16806 10728
rect 2913 10677 2965 10722
tri 2965 10709 2978 10722 nw
tri 16741 10709 16754 10722 ne
rect 16754 10716 16806 10722
tri 8129 10649 8153 10673 se
tri 8281 10658 8296 10673 sw
rect 16754 10658 16806 10664
rect 8281 10649 8296 10658
tri 8296 10649 8305 10658 sw
tri 8119 10639 8129 10649 se
rect 8129 10639 8153 10649
rect 14707 10621 14906 10649
tri 14906 10621 14934 10649 sw
tri 14888 10575 14934 10621 ne
tri 14934 10575 14980 10621 sw
tri 14934 10572 14937 10575 ne
tri 14508 10550 14510 10552 se
rect -60 10531 5785 10537
rect -60 10497 -48 10531
rect -14 10497 25 10531
rect 59 10497 98 10531
rect 132 10497 171 10531
rect 205 10497 244 10531
rect 278 10497 317 10531
rect 351 10497 390 10531
rect 424 10497 463 10531
rect 497 10497 536 10531
rect 570 10497 609 10531
rect 643 10497 682 10531
rect 716 10497 755 10531
rect 789 10497 828 10531
rect 862 10497 901 10531
rect 935 10497 974 10531
rect 1008 10497 1047 10531
rect 1081 10497 1120 10531
rect 1154 10497 1193 10531
rect 1227 10497 1266 10531
rect 1300 10497 1339 10531
rect 1373 10497 1412 10531
rect 1446 10497 1485 10531
rect 1519 10497 1558 10531
rect 1592 10497 1631 10531
rect 1665 10497 1704 10531
rect 1738 10497 1777 10531
rect 1811 10497 1850 10531
rect 1884 10497 1923 10531
rect -60 10459 1923 10497
rect -60 10425 -48 10459
rect -14 10425 25 10459
rect 59 10425 98 10459
rect 132 10425 171 10459
rect 205 10425 244 10459
rect 278 10425 317 10459
rect 351 10425 390 10459
rect 424 10425 463 10459
rect 497 10425 536 10459
rect 570 10425 609 10459
rect 643 10425 682 10459
rect 716 10425 755 10459
rect 789 10425 828 10459
rect 862 10425 901 10459
rect 935 10425 974 10459
rect 1008 10425 1047 10459
rect 1081 10425 1120 10459
rect 1154 10425 1193 10459
rect 1227 10425 1266 10459
rect 1300 10425 1339 10459
rect 1373 10425 1412 10459
rect 1446 10425 1485 10459
rect 1519 10425 1558 10459
rect 1592 10425 1631 10459
rect 1665 10425 1704 10459
rect 1738 10425 1777 10459
rect 1811 10425 1850 10459
rect 1884 10425 1923 10459
rect -60 10387 1923 10425
rect -60 10353 -48 10387
rect -14 10353 25 10387
rect 59 10353 98 10387
rect 132 10353 171 10387
rect 205 10353 244 10387
rect 278 10353 317 10387
rect 351 10353 390 10387
rect 424 10353 463 10387
rect 497 10353 536 10387
rect 570 10353 609 10387
rect 643 10353 682 10387
rect 716 10353 755 10387
rect 789 10353 828 10387
rect 862 10353 901 10387
rect 935 10353 974 10387
rect 1008 10353 1047 10387
rect 1081 10353 1120 10387
rect 1154 10353 1193 10387
rect 1227 10353 1266 10387
rect 1300 10353 1339 10387
rect 1373 10353 1412 10387
rect 1446 10353 1485 10387
rect 1519 10353 1558 10387
rect 1592 10353 1631 10387
rect 1665 10353 1704 10387
rect 1738 10353 1777 10387
rect 1811 10353 1850 10387
rect 1884 10353 1923 10387
rect 5773 10353 5785 10531
tri 14508 10502 14510 10504 ne
rect 6955 10418 6961 10470
rect 7013 10418 7025 10470
rect 7077 10418 9198 10470
rect 9356 10418 9386 10470
rect 9438 10418 9450 10470
rect 9502 10418 14884 10470
tri 14788 10394 14812 10418 ne
rect -60 10347 5785 10353
tri 4019 10338 4028 10347 ne
rect 4028 10338 4073 10347
tri 4028 10310 4056 10338 ne
rect 4056 10310 4073 10338
tri 4056 10293 4073 10310 ne
rect 4585 10338 4630 10347
tri 4630 10338 4639 10347 nw
rect 9983 10338 11947 10390
tri 14508 10352 14510 10354 se
rect 4585 10310 4602 10338
tri 4602 10310 4630 10338 nw
rect 7555 10310 7561 10338
tri 7561 10310 7589 10338 nw
tri 4585 10293 4602 10310 nw
rect 5583 10304 7426 10310
rect 7555 10306 7557 10310
tri 7557 10306 7561 10310 nw
tri 7555 10304 7557 10306 nw
rect 5635 10258 7426 10304
rect 9185 10258 11947 10310
tri 14508 10304 14510 10306 ne
rect 5635 10253 5655 10258
tri 5655 10253 5660 10258 nw
rect 5635 10252 5649 10253
rect 5583 10247 5649 10252
tri 5649 10247 5655 10253 nw
rect 14611 10247 14741 10253
rect 5583 10240 5635 10247
tri 5635 10233 5649 10247 nw
rect 5583 10182 5635 10188
rect 6073 10178 6079 10230
rect 6131 10178 6143 10230
rect 6195 10178 9135 10230
rect 9191 10183 9232 10235
rect 14611 10213 14623 10247
rect 14657 10213 14695 10247
rect 14729 10213 14741 10247
rect 14611 10207 14741 10213
tri 14611 10183 14635 10207 ne
rect 14635 10183 14698 10207
tri 14635 10178 14640 10183 ne
rect 14640 10178 14698 10183
tri 14640 10166 14652 10178 ne
rect -29 10144 87 10150
rect 139 10144 151 10150
rect 203 10144 215 10150
rect 267 10144 279 10150
rect -29 10122 -17 10144
rect 17 10122 56 10144
rect 23 10110 56 10122
rect 267 10110 275 10144
rect 23 10098 87 10110
rect 139 10098 151 10110
rect 203 10098 215 10110
rect 267 10098 279 10110
rect 331 10098 343 10150
rect 395 10098 407 10150
rect 459 10098 471 10150
rect 523 10144 1427 10150
rect 528 10110 567 10144
rect 601 10110 640 10144
rect 674 10110 713 10144
rect 747 10110 786 10144
rect 820 10110 859 10144
rect 893 10110 932 10144
rect 966 10110 1005 10144
rect 1039 10110 1078 10144
rect 1112 10110 1151 10144
rect 1185 10110 1224 10144
rect 1258 10110 1297 10144
rect 1331 10110 1370 10144
rect 1404 10110 1427 10144
rect 523 10098 1427 10110
rect 1479 10098 1491 10150
rect 1543 10144 1555 10150
rect 1607 10144 1619 10150
rect 1671 10144 1683 10150
rect 1735 10144 2247 10150
rect 1550 10110 1555 10144
rect 1769 10110 1808 10144
rect 1842 10110 1881 10144
rect 1915 10110 1954 10144
rect 1988 10110 2027 10144
rect 2061 10110 2100 10144
rect 2134 10110 2173 10144
rect 2207 10110 2246 10144
rect 1543 10098 1555 10110
rect 1607 10098 1619 10110
rect 1671 10098 1683 10110
rect 1735 10098 2247 10110
rect 2299 10098 2311 10150
rect 2363 10098 2375 10150
rect 2427 10098 2439 10150
rect 2491 10144 2503 10150
rect 2555 10144 2999 10150
rect 3051 10144 3063 10150
rect 3115 10144 3127 10150
rect 2499 10110 2503 10144
rect 2572 10110 2611 10144
rect 2645 10110 2684 10144
rect 2718 10110 2757 10144
rect 2791 10110 2830 10144
rect 2864 10110 2903 10144
rect 2937 10110 2976 10144
rect 3115 10110 3122 10144
rect 2491 10098 2503 10110
rect 2555 10098 2999 10110
rect 3051 10098 3063 10110
rect 3115 10098 3127 10110
rect 3179 10098 3191 10150
rect 3243 10098 3255 10150
rect 3307 10144 7645 10150
rect 7697 10144 7709 10150
rect 7761 10144 7773 10150
rect 7825 10144 7837 10150
rect 7889 10144 7901 10150
rect 7953 10144 7965 10150
rect 3307 10110 3341 10144
rect 3375 10110 3414 10144
rect 3448 10110 3487 10144
rect 3521 10110 3560 10144
rect 3594 10110 3633 10144
rect 3667 10110 3706 10144
rect 3740 10110 3779 10144
rect 3813 10110 3852 10144
rect 3886 10110 3925 10144
rect 3959 10110 3998 10144
rect 4032 10110 4071 10144
rect 4105 10110 4144 10144
rect 4178 10110 4216 10144
rect 4250 10110 4288 10144
rect 4322 10110 4360 10144
rect 4394 10110 4432 10144
rect 4466 10110 4504 10144
rect 4538 10110 4576 10144
rect 4610 10110 4648 10144
rect 4682 10110 4720 10144
rect 4754 10110 4792 10144
rect 4826 10110 4864 10144
rect 4898 10110 4936 10144
rect 4970 10110 5008 10144
rect 5042 10110 5080 10144
rect 5114 10110 5152 10144
rect 5186 10110 5224 10144
rect 5258 10110 5296 10144
rect 5330 10110 5368 10144
rect 5402 10110 5440 10144
rect 5474 10110 5512 10144
rect 5546 10110 5584 10144
rect 5618 10110 5656 10144
rect 5690 10110 5728 10144
rect 5762 10110 5800 10144
rect 5834 10110 5872 10144
rect 5906 10110 5944 10144
rect 5978 10110 6016 10144
rect 6050 10110 6088 10144
rect 6122 10110 6160 10144
rect 6194 10110 6232 10144
rect 6266 10110 6304 10144
rect 6338 10110 6376 10144
rect 6410 10110 6448 10144
rect 6482 10110 6520 10144
rect 6554 10110 6592 10144
rect 6626 10110 6664 10144
rect 6698 10110 6736 10144
rect 6770 10110 6808 10144
rect 6842 10110 6880 10144
rect 6914 10110 6952 10144
rect 6986 10110 7024 10144
rect 7058 10110 7096 10144
rect 7130 10110 7168 10144
rect 7202 10110 7240 10144
rect 7274 10110 7312 10144
rect 7346 10110 7384 10144
rect 7418 10110 7456 10144
rect 7490 10110 7528 10144
rect 7562 10110 7600 10144
rect 7634 10110 7645 10144
rect 7706 10110 7709 10144
rect 7953 10110 7960 10144
rect 3307 10098 7645 10110
rect 7697 10098 7709 10110
rect 7761 10098 7773 10110
rect 7825 10098 7837 10110
rect 7889 10098 7901 10110
rect 7953 10098 7965 10110
rect 8017 10098 8029 10150
rect 8081 10144 12758 10150
rect 8081 10110 8104 10144
rect 8138 10110 8176 10144
rect 8210 10110 8248 10144
rect 8282 10110 8320 10144
rect 8354 10110 8392 10144
rect 8426 10110 8464 10144
rect 8498 10110 8536 10144
rect 8570 10110 8608 10144
rect 8642 10110 8680 10144
rect 8714 10110 8752 10144
rect 8786 10110 8824 10144
rect 8858 10110 8896 10144
rect 8930 10110 8968 10144
rect 9002 10110 9040 10144
rect 9074 10110 9112 10144
rect 9146 10110 9184 10144
rect 9218 10110 9256 10144
rect 9290 10110 9328 10144
rect 9362 10110 9400 10144
rect 9434 10110 9472 10144
rect 9506 10110 9544 10144
rect 9578 10110 9616 10144
rect 9650 10110 9688 10144
rect 9722 10110 9760 10144
rect 9794 10110 9832 10144
rect 9866 10110 9904 10144
rect 9938 10110 9976 10144
rect 10010 10110 10048 10144
rect 10082 10110 10120 10144
rect 10154 10110 10192 10144
rect 10226 10110 10264 10144
rect 10298 10110 10336 10144
rect 10370 10110 10408 10144
rect 10442 10110 10480 10144
rect 10514 10110 10552 10144
rect 10586 10110 10624 10144
rect 10658 10110 10696 10144
rect 10730 10110 10768 10144
rect 10802 10110 10840 10144
rect 10874 10110 10912 10144
rect 10946 10110 10984 10144
rect 11018 10110 11056 10144
rect 11090 10110 11128 10144
rect 11162 10110 11200 10144
rect 11234 10110 11272 10144
rect 11306 10110 11344 10144
rect 11378 10110 11416 10144
rect 11450 10110 11488 10144
rect 11522 10110 11560 10144
rect 11594 10110 11632 10144
rect 11666 10110 11704 10144
rect 11738 10110 11776 10144
rect 11810 10110 11848 10144
rect 11882 10110 11920 10144
rect 11954 10110 11992 10144
rect 12026 10110 12064 10144
rect 12098 10110 12136 10144
rect 12170 10110 12208 10144
rect 12242 10110 12280 10144
rect 12314 10110 12352 10144
rect 12386 10110 12424 10144
rect 12458 10110 12496 10144
rect 12530 10110 12568 10144
rect 12602 10110 12640 10144
rect 12674 10110 12712 10144
rect 12746 10110 12758 10144
rect 8081 10098 12758 10110
rect 12934 10144 14599 10150
rect 12934 10110 12946 10144
rect 12980 10110 13020 10144
rect 13054 10110 13093 10144
rect 13127 10110 13166 10144
rect 13200 10110 13239 10144
rect 13273 10110 13312 10144
rect 13346 10110 13385 10144
rect 13419 10110 13458 10144
rect 13492 10110 13531 10144
rect 13565 10110 13604 10144
rect 13638 10110 13677 10144
rect 13711 10110 13750 10144
rect 13784 10110 13823 10144
rect 13857 10110 13896 10144
rect 13930 10110 13969 10144
rect 14003 10110 14042 10144
rect 14076 10110 14115 10144
rect 14149 10110 14188 10144
rect 14222 10110 14261 10144
rect 14295 10110 14334 10144
rect 14368 10110 14407 10144
rect 14441 10110 14480 10144
rect 14514 10110 14553 10144
rect 14587 10110 14599 10144
rect 12934 10098 14599 10110
tri 23 10073 48 10098 nw
rect -29 10058 -17 10070
rect 17 10058 23 10070
tri 14104 10064 14110 10070 se
rect -29 9994 23 10006
rect -29 9930 23 9942
rect 14652 10035 14698 10178
tri 14698 10166 14739 10207 nw
rect 14652 10001 14658 10035
rect 14692 10001 14698 10035
rect 14652 9963 14698 10001
rect 14652 9929 14658 9963
rect 14692 9929 14698 9963
rect 14812 10038 14884 10418
rect 14937 10253 14980 10575
tri 14980 10253 15018 10291 sw
rect 14937 10247 15067 10253
rect 14937 10213 14949 10247
rect 14983 10213 15021 10247
rect 15055 10213 15067 10247
rect 14937 10207 15067 10213
rect 14944 10144 15345 10150
rect 14944 10110 14956 10144
rect 14990 10110 15042 10144
rect 15076 10110 15128 10144
rect 15162 10110 15214 10144
rect 15248 10110 15299 10144
rect 15333 10110 15345 10144
rect 14944 10098 15345 10110
tri 15268 10084 15282 10098 ne
rect 15282 10084 15345 10098
tri 15282 10073 15293 10084 ne
rect 15293 10072 15345 10084
tri 14884 10038 14905 10059 sw
rect 15293 10038 15299 10072
rect 15333 10038 15345 10072
rect 14812 10030 14905 10038
tri 14905 10030 14913 10038 sw
rect 14812 10006 14972 10030
rect 14812 9972 14824 10006
rect 14858 9972 14926 10006
rect 14960 9972 14972 10006
rect 14812 9948 14972 9972
rect 15293 9993 15345 10038
rect 15293 9959 15299 9993
rect 15333 9959 15345 9993
rect 14652 9917 14698 9929
rect -29 9872 23 9878
rect 15293 9915 15345 9959
rect 15293 9881 15299 9915
rect 15333 9881 15345 9915
tri 23 9872 25 9874 sw
tri 15291 9872 15293 9874 se
rect 15293 9872 15345 9881
rect -29 9849 25 9872
tri 25 9849 48 9872 sw
tri 15288 9869 15291 9872 se
rect 15291 9869 15345 9872
tri 15268 9849 15288 9869 se
rect 15288 9849 15345 9869
rect -29 9703 23 9849
rect 1881 9827 1997 9833
rect 1881 9705 1997 9711
rect 4104 9821 4150 9833
rect 4104 9787 4110 9821
rect 4144 9787 4150 9821
rect 4104 9749 4150 9787
rect 4104 9715 4110 9749
rect 4144 9715 4150 9749
rect 4104 9703 4150 9715
rect 4416 9821 4462 9833
rect 4416 9787 4422 9821
rect 4456 9787 4462 9821
rect 4416 9749 4462 9787
rect 4416 9715 4422 9749
rect 4456 9715 4462 9749
rect 4416 9703 4462 9715
rect 4906 9821 4952 9833
rect 4906 9787 4912 9821
rect 4946 9787 4952 9821
rect 4906 9749 4952 9787
rect 4906 9715 4912 9749
rect 4946 9715 4952 9749
rect 4906 9703 4952 9715
rect 5258 9821 5304 9833
rect 5258 9787 5264 9821
rect 5298 9787 5304 9821
rect 5258 9749 5304 9787
rect 5258 9715 5264 9749
rect 5298 9715 5304 9749
rect 5258 9703 5304 9715
rect 6404 9821 6450 9833
rect 6404 9787 6410 9821
rect 6444 9787 6450 9821
rect 6404 9749 6450 9787
rect 6404 9715 6410 9749
rect 6444 9715 6450 9749
rect 6404 9703 6450 9715
rect 6756 9821 6802 9833
rect 6756 9787 6762 9821
rect 6796 9787 6802 9821
rect 6756 9749 6802 9787
rect 6756 9715 6762 9749
rect 6796 9715 6802 9749
rect 6756 9703 6802 9715
rect 7128 9821 7174 9833
rect 7128 9787 7134 9821
rect 7168 9787 7174 9821
rect 7128 9749 7174 9787
rect 7128 9715 7134 9749
rect 7168 9715 7174 9749
rect 7128 9703 7174 9715
rect 7480 9821 7526 9833
rect 7480 9787 7486 9821
rect 7520 9787 7526 9821
rect 7480 9749 7526 9787
rect 7480 9715 7486 9749
rect 7520 9715 7526 9749
rect 7480 9703 7526 9715
rect 12576 9831 15345 9849
rect 12576 9715 14841 9831
rect 15021 9715 15345 9831
rect 12576 9703 15345 9715
tri 15252 9697 15258 9703 ne
rect 15258 9697 15293 9703
tri 15339 9697 15345 9703 nw
tri 15258 9662 15293 9697 ne
tri 8205 9589 8239 9623 nw
tri 8363 9589 8397 9623 ne
rect 13960 9516 13980 9536
rect 7860 9411 8247 9463
rect 8299 9411 8311 9463
rect 8363 9411 8369 9463
rect 9018 9411 9306 9463
rect 9358 9411 9370 9463
rect 9422 9411 9428 9463
rect 9456 9375 9989 9427
rect 10041 9375 10053 9427
rect 10105 9375 10138 9427
rect 6955 9299 6961 9351
rect 7013 9299 7025 9351
rect 7077 9299 7708 9351
rect 1881 9181 1997 9187
rect 13458 9114 13510 9120
tri 13433 9044 13458 9069 se
rect 13458 9050 13510 9062
rect 1881 8995 1997 9001
tri 11869 8995 11918 9044 se
rect 11918 8998 13458 9044
rect 11918 8995 13510 8998
tri 11866 8992 11869 8995 se
rect 11869 8992 13510 8995
tri 11835 8961 11866 8992 se
rect 11866 8961 11928 8992
tri 11928 8961 11959 8992 nw
rect 11508 8909 11876 8961
tri 11876 8909 11928 8961 nw
rect 16494 8726 17092 8732
rect 16546 8680 17092 8726
rect 12484 8463 12614 8665
rect 16494 8662 16546 8674
tri 16546 8644 16582 8680 nw
rect 16494 8604 16546 8610
rect 16586 8612 17092 8618
rect 16638 8566 17092 8612
rect 16586 8548 16638 8560
tri 16638 8530 16674 8566 nw
rect 16586 8490 16638 8496
rect 16678 8441 16684 8493
rect 16736 8441 16748 8493
rect 16800 8441 17000 8493
rect 6999 8365 7005 8417
rect 7057 8412 8601 8417
tri 8601 8412 8606 8417 sw
rect 7057 8365 8606 8412
rect 6999 8353 7063 8365
rect 6999 8301 7005 8353
rect 7057 8301 7063 8353
tri 7063 8340 7088 8365 nw
tri 8579 8340 8604 8365 ne
rect 8604 8340 8606 8365
tri 8604 8338 8606 8340 ne
tri 8606 8338 8680 8412 sw
tri 8606 8301 8643 8338 ne
rect 8643 8301 9890 8338
tri 8643 8286 8658 8301 ne
rect 8658 8286 9890 8301
rect 9942 8286 9954 8338
rect 10006 8286 10012 8338
rect 13845 8196 14462 8203
rect 13845 8144 13851 8196
rect 13903 8144 13921 8196
rect 13973 8144 13990 8196
rect 14042 8144 14059 8196
rect 14111 8144 14128 8196
rect 14180 8144 14197 8196
rect 14249 8144 14266 8196
rect 14318 8144 14335 8196
rect 14387 8144 14404 8196
rect 14456 8144 14462 8196
rect 13845 8132 14462 8144
rect 13845 8080 13851 8132
rect 13903 8080 13921 8132
rect 13973 8080 13990 8132
rect 14042 8080 14059 8132
rect 14111 8080 14128 8132
rect 14180 8080 14197 8132
rect 14249 8080 14266 8132
rect 14318 8080 14335 8132
rect 14387 8080 14404 8132
rect 14456 8080 14462 8132
rect 13845 8073 14462 8080
tri 11991 7893 12043 7945 se
rect 12043 7893 13305 7945
rect 13357 7893 13369 7945
rect 13421 7893 13427 7945
tri 11969 7871 11991 7893 se
rect 11991 7871 12043 7893
tri 12043 7871 12065 7893 nw
tri 11955 7857 11969 7871 se
rect 11969 7857 12029 7871
tri 12029 7857 12043 7871 nw
rect 10569 7805 10575 7857
rect 10627 7805 10639 7857
rect 10691 7805 11977 7857
tri 11977 7805 12029 7857 nw
rect 6233 7748 6239 7800
rect 6291 7748 7005 7800
rect 7057 7748 7063 7800
rect 6233 7736 7063 7748
rect 2913 7719 2965 7725
rect 6233 7684 6239 7736
rect 6291 7684 7005 7736
rect 7057 7684 7063 7736
rect 12015 7715 16459 7721
rect 2913 7655 2965 7667
tri 2965 7649 2990 7674 sw
rect 12067 7663 16407 7715
rect 12015 7651 16459 7663
rect 2965 7603 4806 7649
rect 2913 7597 4806 7603
rect 4858 7597 4870 7649
rect 4922 7597 4928 7649
rect 12067 7599 16407 7651
rect 12015 7593 16459 7599
rect 13845 7558 14462 7565
rect 13845 7506 13851 7558
rect 13903 7506 13921 7558
rect 13973 7506 13990 7558
rect 14042 7506 14059 7558
rect 14111 7506 14128 7558
rect 14180 7506 14197 7558
rect 14249 7506 14266 7558
rect 14318 7506 14335 7558
rect 14387 7506 14404 7558
rect 14456 7506 14462 7558
rect 13845 7494 14462 7506
rect 13845 7442 13851 7494
rect 13903 7442 13921 7494
rect 13973 7442 13990 7494
rect 14042 7442 14059 7494
rect 14111 7442 14128 7494
rect 14180 7442 14197 7494
rect 14249 7442 14266 7494
rect 14318 7442 14335 7494
rect 14387 7442 14404 7494
rect 14456 7442 14462 7494
rect 13845 7435 14462 7442
tri 15424 7435 15490 7501 se
rect 15490 7449 17092 7501
tri 15490 7435 15504 7449 nw
tri 15398 7409 15424 7435 se
rect 15424 7409 15464 7435
tri 15464 7409 15490 7435 nw
tri 15396 7407 15398 7409 se
rect 15398 7407 15462 7409
tri 15462 7407 15464 7409 nw
rect 9884 7355 9890 7407
rect 9942 7355 9954 7407
rect 10006 7361 13423 7407
rect 13507 7367 13541 7401
rect 13625 7361 15416 7407
tri 15416 7361 15462 7407 nw
rect 16225 7403 17092 7409
rect 10006 7355 10012 7361
tri 10012 7355 10018 7361 nw
rect 16277 7357 17092 7403
rect 16225 7339 16277 7351
rect 12251 7281 12257 7327
tri 12245 7280 12246 7281 ne
rect 12246 7280 12257 7281
rect 677 7274 6175 7280
rect 729 7228 6175 7274
rect 6227 7228 6239 7280
rect 6291 7228 6297 7280
tri 12246 7278 12248 7280 ne
rect 12248 7278 12257 7280
rect 729 7226 752 7228
tri 752 7226 754 7228 nw
rect 10493 7226 10499 7278
rect 10551 7226 10563 7278
rect 10615 7226 10621 7278
tri 12248 7275 12251 7278 ne
rect 12251 7275 12257 7278
rect 12309 7275 12321 7327
rect 12373 7275 12379 7327
rect 14245 7281 14533 7327
tri 16277 7332 16302 7357 nw
rect 16225 7281 16277 7287
rect 16407 7323 16459 7329
tri 12379 7275 12385 7281 nw
rect 16407 7269 16459 7271
tri 16459 7269 16468 7278 sw
rect 16407 7259 16468 7269
rect 677 7210 729 7222
tri 729 7203 752 7226 nw
rect 16459 7253 16468 7259
tri 16468 7253 16484 7269 sw
tri 16572 7253 16588 7269 se
rect 16588 7253 17092 7269
rect 16459 7217 17092 7253
rect 16459 7207 16594 7217
rect 16407 7201 16594 7207
tri 16594 7201 16610 7217 nw
tri 16618 7161 16646 7189 se
rect 16646 7161 17092 7189
rect 677 7152 729 7158
rect 16407 7155 17092 7161
rect 16459 7137 17092 7155
rect 16459 7109 16640 7137
tri 16640 7109 16668 7137 nw
rect 16407 7091 16459 7103
tri 16459 7084 16484 7109 nw
rect 16407 7033 16459 7039
rect 10460 6839 10466 7019
rect 10582 6839 10588 7019
rect 11858 6838 11972 6952
rect 14826 6878 14832 6994
rect 15012 6878 15018 6994
rect 23171 6966 23223 6972
tri 23125 6890 23171 6936 se
rect 23171 6902 23223 6914
tri 17716 6878 17728 6890 se
rect 17728 6878 23171 6890
tri 17677 6839 17716 6878 se
rect 17716 6850 23171 6878
rect 17716 6844 23223 6850
rect 17716 6839 17736 6844
tri 17676 6838 17677 6839 se
rect 17677 6838 17736 6839
tri 17670 6832 17676 6838 se
rect 17676 6832 17736 6838
tri 17736 6832 17748 6844 nw
tri 16234 6785 16281 6832 se
rect 16281 6786 17690 6832
tri 17690 6786 17736 6832 nw
rect 16035 6779 16087 6785
tri 5790 6736 5808 6754 se
rect 5808 6736 5814 6754
rect 1820 6684 1826 6736
rect 1878 6684 1890 6736
rect 1942 6702 5814 6736
rect 5866 6702 5878 6754
rect 5930 6702 5936 6754
tri 15984 6703 16035 6754 se
tri 16215 6766 16234 6785 se
rect 16234 6766 16281 6785
tri 16281 6766 16301 6786 nw
rect 16035 6715 16087 6727
tri 13453 6702 13454 6703 se
rect 13454 6702 16035 6703
rect 1942 6684 1948 6702
tri 1948 6684 1966 6702 nw
tri 13435 6684 13453 6702 se
rect 13453 6684 16035 6702
tri 13408 6657 13435 6684 se
rect 13435 6663 16035 6684
rect 13435 6657 16087 6663
tri 16179 6730 16215 6766 se
rect 16215 6730 16245 6766
tri 16245 6730 16281 6766 nw
tri 13388 6637 13408 6657 se
rect 13408 6637 13454 6657
tri 13454 6637 13474 6657 nw
tri 13365 6614 13388 6637 se
rect 13388 6614 13431 6637
tri 13431 6614 13454 6637 nw
tri 13339 6588 13365 6614 se
rect 13365 6588 13405 6614
tri 13405 6588 13431 6614 nw
tri 15202 6588 15228 6614 se
rect 15228 6608 16001 6614
rect 15228 6588 15949 6608
rect 12402 6548 12436 6582
rect 13188 6542 13359 6588
tri 13359 6542 13405 6588 nw
rect 13866 6548 13900 6582
rect 14299 6568 15949 6588
rect 14299 6542 15222 6568
tri 15222 6542 15248 6568 nw
tri 15924 6543 15949 6568 ne
rect 15949 6544 16001 6556
rect 5675 6451 5681 6503
rect 5733 6451 5739 6503
rect 5675 6439 5739 6451
rect 5675 6387 5681 6439
rect 5733 6387 5739 6439
rect 5675 6375 5739 6387
rect 5675 6323 5681 6375
rect 5733 6323 5739 6375
rect 5969 6451 5975 6503
rect 6027 6451 6033 6503
rect 15949 6486 16001 6492
rect 5969 6439 6033 6451
rect 5969 6387 5975 6439
rect 6027 6387 6033 6439
rect 5969 6375 6033 6387
rect 5969 6323 5975 6375
rect 6027 6323 6033 6375
rect 1284 6186 1336 6192
tri 16150 6135 16179 6164 se
rect 16179 6144 16225 6730
tri 16225 6710 16245 6730 nw
rect 1284 6122 1336 6134
tri 1336 6110 1361 6135 sw
tri 16125 6110 16150 6135 se
rect 16150 6110 16179 6135
rect 1336 6070 2355 6110
tri 16115 6100 16125 6110 se
rect 16125 6100 16179 6110
rect 1284 6064 2355 6070
rect 7619 6056 8292 6100
rect 7619 6036 7682 6056
tri 7682 6036 7702 6056 nw
tri 8261 6036 8281 6056 ne
rect 8281 6048 8292 6056
rect 8344 6048 8350 6100
tri 16113 6098 16115 6100 se
rect 16115 6098 16179 6100
tri 16179 6098 16225 6144 nw
tri 16073 6058 16113 6098 se
rect 8281 6036 8350 6048
tri 2234 6030 2240 6036 se
rect 2240 5984 2246 6036
rect 2298 5984 2310 6036
rect 2362 5984 2368 6036
tri 2368 6030 2374 6036 sw
rect 7619 6028 7677 6036
tri 7677 6031 7682 6036 nw
tri 8281 6031 8286 6036 ne
rect 8286 5984 8292 6036
rect 8344 5984 8350 6036
rect 9496 6032 9504 6058
tri 9504 6032 9530 6058 nw
tri 16047 6032 16073 6058 se
rect 16073 6032 16113 6058
tri 16113 6032 16179 6098 nw
rect 9496 6030 9502 6032
tri 9502 6030 9504 6032 nw
tri 16045 6030 16047 6032 se
rect 16047 6030 16095 6032
tri 9496 6024 9502 6030 nw
rect 12171 6024 14234 6030
rect 12223 6014 14234 6024
tri 14234 6014 14250 6030 sw
tri 16029 6014 16045 6030 se
rect 16045 6014 16095 6030
tri 16095 6014 16113 6032 nw
rect 12223 6008 14250 6014
tri 14250 6008 14256 6014 sw
rect 14541 6008 16049 6014
rect 12223 6006 14256 6008
tri 14256 6006 14258 6008 sw
rect 12223 5978 14258 6006
rect 12223 5974 12244 5978
tri 12244 5974 12248 5978 nw
tri 14212 5974 14216 5978 ne
rect 14216 5974 14258 5978
tri 14258 5974 14290 6006 sw
rect 14541 5974 14553 6008
rect 14587 5974 16049 6008
rect 12015 5960 12067 5966
rect 11412 5950 11470 5956
rect 11412 5916 11424 5950
rect 11458 5916 11470 5950
rect 2788 5876 2915 5882
rect 2840 5824 2915 5876
rect 11412 5878 11470 5916
rect 11412 5844 11424 5878
rect 11458 5872 11470 5878
tri 11470 5872 11495 5897 sw
tri 11990 5872 12015 5897 se
rect 12015 5896 12067 5908
rect 12171 5960 12223 5972
tri 12223 5953 12244 5974 nw
tri 14216 5953 14237 5974 ne
rect 14237 5953 14290 5974
tri 14237 5936 14254 5953 ne
rect 14254 5936 14290 5953
tri 14290 5936 14328 5974 sw
rect 14541 5968 16049 5974
tri 16049 5968 16095 6014 nw
rect 14541 5936 14599 5968
tri 14599 5943 14624 5968 nw
tri 14254 5932 14258 5936 ne
rect 14258 5932 14328 5936
tri 14328 5932 14332 5936 sw
rect 12171 5902 12223 5908
tri 14258 5902 14288 5932 ne
rect 14288 5902 14332 5932
tri 14332 5902 14362 5932 sw
rect 14541 5902 14553 5936
rect 14587 5902 14599 5936
rect 11458 5844 12015 5872
tri 14288 5858 14332 5902 ne
rect 14332 5896 14362 5902
tri 14362 5896 14368 5902 sw
rect 14541 5896 14599 5902
rect 16225 5906 16277 5912
rect 14332 5858 14368 5896
tri 14368 5858 14406 5896 sw
rect 11412 5838 12067 5844
tri 14332 5838 14352 5858 ne
rect 14352 5838 14406 5858
tri 14406 5838 14426 5858 sw
rect 16225 5842 16277 5854
rect 2788 5812 2915 5824
rect 926 5800 1049 5806
tri 901 5736 926 5761 se
rect 978 5753 1049 5800
rect 2840 5760 2915 5812
tri 14352 5808 14382 5838 ne
rect 14382 5809 14426 5838
tri 14426 5809 14455 5838 sw
rect 14382 5808 14455 5809
tri 8722 5784 8746 5808 se
tri 14382 5784 14406 5808 ne
rect 14406 5784 14455 5808
tri 14455 5784 14480 5809 sw
tri 16200 5784 16225 5809 se
rect 16225 5784 16277 5790
tri 8712 5774 8722 5784 se
rect 8722 5774 8746 5784
tri 14406 5774 14416 5784 ne
rect 14416 5774 16277 5784
rect 2788 5754 2915 5760
tri 14416 5754 14436 5774 ne
rect 14436 5754 16277 5774
tri 14436 5753 14437 5754 ne
rect 14437 5753 16277 5754
rect 978 5748 992 5753
tri 14437 5752 14438 5753 ne
rect 14438 5752 16277 5753
rect 926 5736 992 5748
rect 978 5684 992 5736
tri 8712 5732 8732 5752 ne
rect 8732 5732 8746 5752
tri 14438 5732 14458 5752 ne
rect 14458 5732 16277 5752
tri 8732 5718 8746 5732 ne
rect 926 5678 992 5684
tri 16355 5678 16377 5700 se
tri 16277 5600 16355 5678 se
rect 16355 5600 16377 5678
tri 16254 5236 16354 5336 ne
tri 4067 5198 4073 5204 se
tri 4585 5198 4591 5204 sw
tri 12666 5198 12672 5204 se
rect 12672 5152 12678 5204
rect 12730 5152 12742 5204
rect 12794 5152 12806 5204
rect 12858 5152 12864 5204
tri 12864 5198 12870 5204 sw
rect 15158 5180 16054 5187
rect 15158 5164 15714 5180
rect 15766 5164 15786 5180
rect 15838 5164 15858 5180
rect 15158 5130 15170 5164
rect 15204 5130 15247 5164
rect 15281 5130 15324 5164
rect 15358 5130 15400 5164
rect 15434 5130 15476 5164
rect 15510 5130 15552 5164
rect 15586 5130 15628 5164
rect 15662 5130 15704 5164
rect 15766 5130 15780 5164
rect 15838 5130 15856 5164
rect 15158 5128 15714 5130
rect 15766 5128 15786 5130
rect 15838 5128 15858 5130
rect 15910 5128 15930 5180
rect 15982 5128 16002 5180
rect 15158 5101 16054 5128
rect 15158 5092 15714 5101
rect 15766 5092 15786 5101
rect 15838 5092 15858 5101
rect 15158 5058 15170 5092
rect 15204 5058 15247 5092
rect 15281 5058 15324 5092
rect 15358 5058 15400 5092
rect 15434 5058 15476 5092
rect 15510 5058 15552 5092
rect 15586 5058 15628 5092
rect 15662 5058 15704 5092
rect 15766 5058 15780 5092
rect 15838 5058 15856 5092
rect 15158 5049 15714 5058
rect 15766 5049 15786 5058
rect 15838 5049 15858 5058
rect 15910 5049 15930 5101
rect 15982 5049 16002 5101
rect 15158 5021 16054 5049
rect 15158 5020 15714 5021
rect 15766 5020 15786 5021
rect 15838 5020 15858 5021
rect 15158 4986 15170 5020
rect 15204 4986 15247 5020
rect 15281 4986 15324 5020
rect 15358 4986 15400 5020
rect 15434 4986 15476 5020
rect 15510 4986 15552 5020
rect 15586 4986 15628 5020
rect 15662 4986 15704 5020
rect 15766 4986 15780 5020
rect 15838 4986 15856 5020
rect 15158 4969 15714 4986
rect 15766 4969 15786 4986
rect 15838 4969 15858 4986
rect 15910 4969 15930 5021
rect 15982 4969 16002 5021
rect 15158 4963 16054 4969
rect 1458 4838 1890 4884
tri 1859 4813 1884 4838 ne
rect 1884 4832 1890 4838
rect 1942 4832 1948 4884
tri 3536 4864 3542 4870 se
rect 1884 4820 1948 4832
rect 1884 4768 1890 4820
rect 1942 4768 1948 4820
rect 3542 4818 3548 4870
rect 3600 4818 3612 4870
rect 3664 4818 3670 4870
tri 3670 4864 3676 4870 sw
rect 12015 4810 12067 4816
rect 12015 4746 12067 4758
tri 13212 4750 13215 4753 se
tri 12067 4740 12077 4750 sw
tri 13202 4740 13212 4750 se
rect 13212 4740 13215 4750
rect 12067 4737 12077 4740
tri 12077 4737 12080 4740 sw
tri 13199 4737 13202 4740 se
rect 13202 4737 13215 4740
tri 13713 4737 13716 4740 se
rect 13716 4737 16183 4740
tri 16183 4737 16186 4740 sw
rect 12067 4725 12080 4737
tri 12080 4725 12092 4737 sw
tri 13187 4725 13199 4737 se
rect 13199 4725 13215 4737
tri 13701 4725 13713 4737 se
rect 13713 4725 16186 4737
rect 12067 4694 16186 4725
rect 12015 4688 16186 4694
tri 16186 4688 16235 4737 sw
tri 16161 4663 16186 4688 ne
rect 16186 4663 16235 4688
tri 16235 4663 16260 4688 sw
tri 16186 4660 16189 4663 ne
rect 16189 4660 16260 4663
rect 117 4480 123 4660
rect 239 4480 245 4660
tri 16189 4653 16196 4660 ne
rect 16196 4653 16260 4660
rect 10460 4473 10466 4653
rect 10582 4473 10588 4653
tri 16196 4641 16208 4653 ne
rect 50 4468 60 4472
rect 2236 4266 2288 4272
tri 2211 4195 2236 4220 ne
rect 2236 4202 2288 4214
tri 2288 4195 2313 4220 nw
rect 2236 4144 2288 4150
rect 12251 4140 12257 4192
rect 12309 4140 12321 4192
rect 12373 4140 12379 4192
rect 401 4085 658 4091
rect 401 3969 410 4085
rect 526 3969 658 4085
rect 12390 4048 12434 4100
rect 401 3963 658 3969
rect 4242 3809 4248 3861
rect 4300 3809 4312 3861
rect 4364 3809 4370 3861
rect 54 3766 175 3772
rect 106 3714 175 3766
rect 16208 3729 16260 4653
tri 16675 3840 16723 3888 ne
tri 16775 3840 16823 3888 nw
tri 16208 3728 16209 3729 ne
rect 16209 3728 16260 3729
tri 16260 3728 16283 3751 sw
rect 54 3702 175 3714
rect 106 3650 175 3702
tri 16209 3701 16236 3728 ne
rect 16236 3701 16283 3728
rect 4071 3667 4105 3701
tri 16236 3677 16260 3701 ne
rect 16260 3677 16283 3701
tri 16260 3671 16266 3677 ne
rect 16266 3671 16283 3677
tri 16283 3671 16340 3728 sw
rect 54 3644 175 3650
rect 7335 3619 7341 3671
rect 7393 3619 7405 3671
rect 7457 3665 9442 3671
tri 9442 3665 9448 3671 sw
tri 16266 3665 16272 3671 ne
rect 16272 3665 16340 3671
rect 7457 3657 9448 3665
tri 9448 3657 9456 3665 sw
tri 16272 3657 16280 3665 ne
rect 16280 3657 16340 3665
tri 16340 3657 16354 3671 sw
rect 7457 3651 9456 3657
tri 9456 3651 9462 3657 sw
rect 11621 3651 11679 3657
tri 16280 3654 16283 3657 ne
rect 16283 3654 16354 3657
tri 16354 3654 16357 3657 sw
rect 7457 3619 9462 3651
tri 9462 3619 9494 3651 sw
tri 9420 3617 9422 3619 ne
rect 9422 3617 9494 3619
tri 9494 3617 9496 3619 sw
rect 11621 3617 11633 3651
rect 11667 3617 11679 3651
tri 9422 3591 9448 3617 ne
rect 9448 3616 9496 3617
tri 9496 3616 9497 3617 sw
rect 9448 3591 9497 3616
tri 9497 3591 9522 3616 sw
tri 11596 3591 11621 3616 se
rect 11621 3591 11679 3617
tri 16283 3602 16335 3654 ne
rect 16335 3602 17240 3654
rect 17292 3602 17304 3654
rect 17356 3602 17362 3654
rect 4242 3539 4248 3591
rect 4300 3539 4312 3591
rect 4364 3539 4376 3591
rect 4428 3539 4440 3591
rect 4492 3579 4498 3591
tri 4498 3579 4510 3591 sw
tri 9448 3579 9460 3591 ne
rect 9460 3579 11247 3591
rect 4492 3545 4510 3579
tri 4510 3545 4544 3579 sw
tri 9460 3545 9494 3579 ne
rect 9494 3545 11247 3579
rect 4492 3539 4544 3545
tri 4544 3539 4550 3545 sw
tri 9494 3539 9500 3545 ne
rect 9500 3539 11247 3545
rect 11299 3539 11311 3591
rect 11363 3579 11679 3591
rect 11363 3545 11633 3579
rect 11667 3545 11679 3579
rect 11363 3539 11679 3545
rect 410 3501 526 3507
rect 410 3315 526 3321
rect 7178 3500 7294 3506
rect 19766 3499 20585 3507
rect 19766 3447 19772 3499
rect 19824 3447 19841 3499
rect 19893 3447 19910 3499
rect 19962 3447 19979 3499
rect 20031 3447 20048 3499
rect 20100 3447 20117 3499
rect 20169 3447 20186 3499
rect 20238 3447 20255 3499
rect 20307 3447 20323 3499
rect 20375 3447 20391 3499
rect 20443 3447 20459 3499
rect 20511 3447 20527 3499
rect 20579 3447 20585 3499
rect 7178 3314 7294 3320
rect 12185 3431 12237 3437
rect 12185 3367 12237 3379
rect 12185 3309 12237 3315
rect 19766 3435 20585 3447
rect 19766 3383 19772 3435
rect 19824 3383 19841 3435
rect 19893 3383 19910 3435
rect 19962 3383 19979 3435
rect 20031 3383 20048 3435
rect 20100 3383 20117 3435
rect 20169 3383 20186 3435
rect 20238 3383 20255 3435
rect 20307 3383 20323 3435
rect 20375 3383 20391 3435
rect 20443 3383 20459 3435
rect 20511 3383 20527 3435
rect 20579 3383 20585 3435
rect 21156 3505 21348 3507
rect 21156 3389 21162 3505
rect 21342 3389 21348 3505
rect 21156 3387 21348 3389
rect 19766 3371 20585 3383
rect 19766 3319 19772 3371
rect 19824 3319 19841 3371
rect 19893 3319 19910 3371
rect 19962 3319 19979 3371
rect 20031 3319 20048 3371
rect 20100 3319 20117 3371
rect 20169 3319 20186 3371
rect 20238 3319 20255 3371
rect 20307 3319 20323 3371
rect 20375 3319 20391 3371
rect 20443 3319 20459 3371
rect 20511 3319 20527 3371
rect 20579 3319 20585 3371
rect 19766 3311 20585 3319
tri 6629 3281 6657 3309 ne
rect 6657 3281 6663 3309
rect 2003 3275 2055 3281
tri 6657 3275 6663 3281 ne
tri 1978 3210 2003 3235 ne
rect 2003 3211 2055 3223
tri 2055 3210 2080 3235 nw
tri 6662 3210 6663 3211 se
tri 6629 3177 6662 3210 se
rect 6662 3177 6663 3210
rect 2003 3153 2055 3159
rect 54 3096 106 3102
rect 1364 3096 1416 3102
rect 54 3032 106 3044
tri 106 3026 131 3051 sw
tri 1339 3026 1364 3051 se
rect 1364 3032 1416 3044
rect 106 2980 1364 3026
rect 12185 3027 12237 3033
rect 54 2974 1416 2980
tri 12173 2974 12185 2986 se
rect 12185 2974 12237 2975
tri 12160 2961 12173 2974 se
rect 12173 2963 12237 2974
rect 12173 2961 12185 2963
rect 7014 2906 7020 2958
rect 7072 2906 7084 2958
rect 7136 2906 7142 2958
rect 12185 2905 12237 2911
rect 247 2714 285 2758
tri 20663 2706 20669 2712 se
rect 20669 2706 20675 2712
rect 20663 2660 20675 2706
rect 20727 2660 20739 2712
rect 20791 2660 20803 2712
rect 20855 2660 20867 2712
rect 20919 2706 20925 2712
tri 20925 2706 20931 2712 sw
rect 20919 2660 20931 2706
rect 48 2606 56 2617
rect 126 2519 132 2635
rect 312 2519 318 2635
rect 1006 2584 1012 2636
rect 1064 2584 1101 2636
rect 1153 2584 1190 2636
rect 1242 2584 1278 2636
rect 1330 2584 1336 2636
rect 1006 2570 1336 2584
rect 1006 2518 1012 2570
rect 1064 2518 1101 2570
rect 1153 2518 1190 2570
rect 1242 2518 1278 2570
rect 1330 2518 1336 2570
rect 2396 2519 2402 2635
rect 2518 2519 2524 2635
rect 3622 2438 3628 2490
rect 3680 2438 3692 2490
rect 3744 2438 5578 2490
rect 5630 2438 5642 2490
rect 5694 2438 5700 2490
rect 8956 2450 8989 2483
rect 10128 2450 10162 2484
rect 12395 2457 12855 2463
tri 12392 2438 12395 2441 se
rect 12395 2438 12407 2457
tri 12377 2423 12392 2438 se
rect 12392 2423 12407 2438
rect 12441 2423 12488 2457
rect 12522 2423 12569 2457
rect 12603 2423 12649 2457
rect 12683 2423 12729 2457
rect 12763 2423 12809 2457
rect 12843 2423 12855 2457
tri 12371 2417 12377 2423 se
rect 12377 2417 12855 2423
tri 12370 2416 12371 2417 se
rect 12371 2416 12855 2417
tri 7409 2407 7418 2416 se
rect 7418 2407 7546 2416
tri 7404 2402 7409 2407 se
rect 7409 2402 7546 2407
rect 7418 2364 7546 2402
rect 7598 2364 7610 2416
rect 7662 2408 7668 2416
tri 7668 2408 7670 2410 sw
rect 7662 2364 7670 2408
rect 11940 2407 12413 2416
rect 11940 2373 11952 2407
rect 11986 2373 12024 2407
rect 12058 2373 12413 2407
rect 11940 2364 12413 2373
rect 12465 2364 12477 2416
rect 12529 2364 12541 2416
rect 12593 2364 12605 2416
rect 12657 2364 12669 2416
rect 12721 2364 12733 2416
rect 12785 2364 12797 2416
rect 12849 2364 12855 2416
rect 7418 2362 7670 2364
rect 16407 2320 16459 2326
rect 4972 2286 5009 2320
tri 16391 2286 16407 2302 se
tri 16355 2250 16391 2286 se
rect 16391 2268 16407 2286
rect 16391 2256 16459 2268
rect 16391 2250 16407 2256
tri 16459 2250 16511 2302 sw
rect 16407 2198 16459 2204
tri 14745 2101 14808 2164 sw
tri 14753 1902 14760 1909 nw
rect 16145 1842 16185 2044
rect 20651 2032 20933 2035
rect 20651 1980 20657 2032
rect 20709 1980 20730 2032
rect 20782 1980 20803 2032
rect 20855 1980 20875 2032
rect 20927 1980 20933 2032
rect 20651 1968 20933 1980
rect 20651 1916 20657 1968
rect 20709 1916 20730 1968
rect 20782 1916 20803 1968
rect 20855 1916 20875 1968
rect 20927 1916 20933 1968
rect 20651 1904 20933 1916
rect 20651 1852 20657 1904
rect 20709 1852 20730 1904
rect 20782 1852 20803 1904
rect 20855 1852 20875 1904
rect 20927 1852 20933 1904
rect 20651 1849 20933 1852
<< via1 >>
rect 2080 13572 2110 13600
rect 2110 13572 2132 13600
rect 2146 13572 2188 13600
rect 2188 13572 2198 13600
rect 2212 13572 2222 13600
rect 2222 13572 2264 13600
rect 2278 13572 2300 13600
rect 2300 13572 2330 13600
rect 2080 13548 2132 13572
rect 2146 13548 2198 13572
rect 2212 13548 2264 13572
rect 2278 13548 2330 13572
rect 2344 13572 2378 13600
rect 2378 13572 2396 13600
rect 2344 13548 2396 13572
rect 2410 13572 2422 13600
rect 2422 13572 2456 13600
rect 2456 13572 2462 13600
rect 2410 13548 2462 13572
rect 2476 13572 2500 13600
rect 2500 13572 2528 13600
rect 2542 13572 2578 13600
rect 2578 13572 2594 13600
rect 2476 13548 2528 13572
rect 2542 13548 2594 13572
rect 2080 13532 2132 13536
rect 2146 13532 2198 13536
rect 2212 13532 2264 13536
rect 2278 13532 2330 13536
rect 2080 13498 2110 13532
rect 2110 13498 2132 13532
rect 2146 13498 2188 13532
rect 2188 13498 2198 13532
rect 2212 13498 2222 13532
rect 2222 13498 2264 13532
rect 2278 13498 2300 13532
rect 2300 13498 2330 13532
rect 2080 13484 2132 13498
rect 2146 13484 2198 13498
rect 2212 13484 2264 13498
rect 2278 13484 2330 13498
rect 2344 13532 2396 13536
rect 2344 13498 2378 13532
rect 2378 13498 2396 13532
rect 2344 13484 2396 13498
rect 2410 13532 2462 13536
rect 2410 13498 2422 13532
rect 2422 13498 2456 13532
rect 2456 13498 2462 13532
rect 2410 13484 2462 13498
rect 2476 13532 2528 13536
rect 2542 13532 2594 13536
rect 2476 13498 2500 13532
rect 2500 13498 2528 13532
rect 2542 13498 2578 13532
rect 2578 13498 2594 13532
rect 2476 13484 2528 13498
rect 2542 13484 2594 13498
rect 2080 13458 2132 13472
rect 2146 13458 2198 13472
rect 2212 13458 2264 13472
rect 2278 13458 2330 13472
rect 2080 13424 2110 13458
rect 2110 13424 2132 13458
rect 2146 13424 2188 13458
rect 2188 13424 2198 13458
rect 2212 13424 2222 13458
rect 2222 13424 2264 13458
rect 2278 13424 2300 13458
rect 2300 13424 2330 13458
rect 2080 13420 2132 13424
rect 2146 13420 2198 13424
rect 2212 13420 2264 13424
rect 2278 13420 2330 13424
rect 2344 13458 2396 13472
rect 2344 13424 2378 13458
rect 2378 13424 2396 13458
rect 2344 13420 2396 13424
rect 2410 13458 2462 13472
rect 2410 13424 2422 13458
rect 2422 13424 2456 13458
rect 2456 13424 2462 13458
rect 2410 13420 2462 13424
rect 2476 13458 2528 13472
rect 2542 13458 2594 13472
rect 2476 13424 2500 13458
rect 2500 13424 2528 13458
rect 2542 13424 2578 13458
rect 2578 13424 2594 13458
rect 2476 13420 2528 13424
rect 2542 13420 2594 13424
rect 2080 13383 2132 13408
rect 2146 13383 2198 13408
rect 2212 13383 2264 13408
rect 2278 13383 2330 13408
rect 2080 13356 2110 13383
rect 2110 13356 2132 13383
rect 2146 13356 2188 13383
rect 2188 13356 2198 13383
rect 2212 13356 2222 13383
rect 2222 13356 2264 13383
rect 2278 13356 2300 13383
rect 2300 13356 2330 13383
rect 2344 13383 2396 13408
rect 2344 13356 2378 13383
rect 2378 13356 2396 13383
rect 2410 13383 2462 13408
rect 2410 13356 2422 13383
rect 2422 13356 2456 13383
rect 2456 13356 2462 13383
rect 2476 13383 2528 13408
rect 2542 13383 2594 13408
rect 2476 13356 2500 13383
rect 2500 13356 2528 13383
rect 2542 13356 2578 13383
rect 2578 13356 2594 13383
rect 2080 13308 2132 13344
rect 2146 13308 2198 13344
rect 2212 13308 2264 13344
rect 2278 13308 2330 13344
rect 2080 13292 2110 13308
rect 2110 13292 2132 13308
rect 2146 13292 2188 13308
rect 2188 13292 2198 13308
rect 2212 13292 2222 13308
rect 2222 13292 2264 13308
rect 2278 13292 2300 13308
rect 2300 13292 2330 13308
rect 2344 13308 2396 13344
rect 2344 13292 2378 13308
rect 2378 13292 2396 13308
rect 2410 13308 2462 13344
rect 2410 13292 2422 13308
rect 2422 13292 2456 13308
rect 2456 13292 2462 13308
rect 2476 13308 2528 13344
rect 2542 13308 2594 13344
rect 2476 13292 2500 13308
rect 2500 13292 2528 13308
rect 2542 13292 2578 13308
rect 2578 13292 2594 13308
rect 2080 13274 2110 13280
rect 2110 13274 2132 13280
rect 2146 13274 2188 13280
rect 2188 13274 2198 13280
rect 2212 13274 2222 13280
rect 2222 13274 2264 13280
rect 2278 13274 2300 13280
rect 2300 13274 2330 13280
rect 2080 13233 2132 13274
rect 2146 13233 2198 13274
rect 2212 13233 2264 13274
rect 2278 13233 2330 13274
rect 2080 13228 2110 13233
rect 2110 13228 2132 13233
rect 2146 13228 2188 13233
rect 2188 13228 2198 13233
rect 2212 13228 2222 13233
rect 2222 13228 2264 13233
rect 2278 13228 2300 13233
rect 2300 13228 2330 13233
rect 2344 13274 2378 13280
rect 2378 13274 2396 13280
rect 2344 13233 2396 13274
rect 2344 13228 2378 13233
rect 2378 13228 2396 13233
rect 2410 13274 2422 13280
rect 2422 13274 2456 13280
rect 2456 13274 2462 13280
rect 2410 13233 2462 13274
rect 2410 13228 2422 13233
rect 2422 13228 2456 13233
rect 2456 13228 2462 13233
rect 2476 13274 2500 13280
rect 2500 13274 2528 13280
rect 2542 13274 2578 13280
rect 2578 13274 2594 13280
rect 2476 13233 2528 13274
rect 2542 13233 2594 13274
rect 2476 13228 2500 13233
rect 2500 13228 2528 13233
rect 2542 13228 2578 13233
rect 2578 13228 2594 13233
rect 2080 13199 2110 13215
rect 2110 13199 2132 13215
rect 2146 13199 2188 13215
rect 2188 13199 2198 13215
rect 2212 13199 2222 13215
rect 2222 13199 2264 13215
rect 2278 13199 2300 13215
rect 2300 13199 2330 13215
rect 2080 13163 2132 13199
rect 2146 13163 2198 13199
rect 2212 13163 2264 13199
rect 2278 13163 2330 13199
rect 2344 13199 2378 13215
rect 2378 13199 2396 13215
rect 2344 13163 2396 13199
rect 2410 13199 2422 13215
rect 2422 13199 2456 13215
rect 2456 13199 2462 13215
rect 2410 13163 2462 13199
rect 2476 13199 2500 13215
rect 2500 13199 2528 13215
rect 2542 13199 2578 13215
rect 2578 13199 2594 13215
rect 2476 13163 2528 13199
rect 2542 13163 2594 13199
rect 2080 13124 2110 13150
rect 2110 13124 2132 13150
rect 2146 13124 2188 13150
rect 2188 13124 2198 13150
rect 2212 13124 2222 13150
rect 2222 13124 2264 13150
rect 2278 13124 2300 13150
rect 2300 13124 2330 13150
rect 2080 13098 2132 13124
rect 2146 13098 2198 13124
rect 2212 13098 2264 13124
rect 2278 13098 2330 13124
rect 2344 13124 2378 13150
rect 2378 13124 2396 13150
rect 2344 13098 2396 13124
rect 2410 13124 2422 13150
rect 2422 13124 2456 13150
rect 2456 13124 2462 13150
rect 2410 13098 2462 13124
rect 2476 13124 2500 13150
rect 2500 13124 2528 13150
rect 2542 13124 2578 13150
rect 2578 13124 2594 13150
rect 2476 13098 2528 13124
rect 2542 13098 2594 13124
rect 2080 13083 2132 13085
rect 2146 13083 2198 13085
rect 2212 13083 2264 13085
rect 2278 13083 2330 13085
rect 2080 13049 2110 13083
rect 2110 13049 2132 13083
rect 2146 13049 2188 13083
rect 2188 13049 2198 13083
rect 2212 13049 2222 13083
rect 2222 13049 2264 13083
rect 2278 13049 2300 13083
rect 2300 13049 2330 13083
rect 2080 13033 2132 13049
rect 2146 13033 2198 13049
rect 2212 13033 2264 13049
rect 2278 13033 2330 13049
rect 2344 13083 2396 13085
rect 2344 13049 2378 13083
rect 2378 13049 2396 13083
rect 2344 13033 2396 13049
rect 2410 13083 2462 13085
rect 2410 13049 2422 13083
rect 2422 13049 2456 13083
rect 2456 13049 2462 13083
rect 2410 13033 2462 13049
rect 2476 13083 2528 13085
rect 2542 13083 2594 13085
rect 2476 13049 2500 13083
rect 2500 13049 2528 13083
rect 2542 13049 2578 13083
rect 2578 13049 2594 13083
rect 2476 13033 2528 13049
rect 2542 13033 2594 13049
rect 2080 13008 2132 13020
rect 2146 13008 2198 13020
rect 2212 13008 2264 13020
rect 2278 13008 2330 13020
rect 2080 12974 2110 13008
rect 2110 12974 2132 13008
rect 2146 12974 2188 13008
rect 2188 12974 2198 13008
rect 2212 12974 2222 13008
rect 2222 12974 2264 13008
rect 2278 12974 2300 13008
rect 2300 12974 2330 13008
rect 2080 12968 2132 12974
rect 2146 12968 2198 12974
rect 2212 12968 2264 12974
rect 2278 12968 2330 12974
rect 2344 13008 2396 13020
rect 2344 12974 2378 13008
rect 2378 12974 2396 13008
rect 2344 12968 2396 12974
rect 2410 13008 2462 13020
rect 2410 12974 2422 13008
rect 2422 12974 2456 13008
rect 2456 12974 2462 13008
rect 2410 12968 2462 12974
rect 2476 13008 2528 13020
rect 2542 13008 2594 13020
rect 2476 12974 2500 13008
rect 2500 12974 2528 13008
rect 2542 12974 2578 13008
rect 2578 12974 2594 13008
rect 2476 12968 2528 12974
rect 2542 12968 2594 12974
rect 2080 12933 2132 12955
rect 2146 12933 2198 12955
rect 2212 12933 2264 12955
rect 2278 12933 2330 12955
rect 2080 12903 2110 12933
rect 2110 12903 2132 12933
rect 2146 12903 2188 12933
rect 2188 12903 2198 12933
rect 2212 12903 2222 12933
rect 2222 12903 2264 12933
rect 2278 12903 2300 12933
rect 2300 12903 2330 12933
rect 2344 12933 2396 12955
rect 2344 12903 2378 12933
rect 2378 12903 2396 12933
rect 2410 12933 2462 12955
rect 2410 12903 2422 12933
rect 2422 12903 2456 12933
rect 2456 12903 2462 12933
rect 2476 12933 2528 12955
rect 2542 12933 2594 12955
rect 2476 12903 2500 12933
rect 2500 12903 2528 12933
rect 2542 12903 2578 12933
rect 2578 12903 2594 12933
rect 2066 12364 2118 12368
rect 2066 12330 2082 12364
rect 2082 12330 2116 12364
rect 2116 12330 2118 12364
rect 2066 12316 2118 12330
rect 2131 12364 2183 12368
rect 2196 12364 2248 12368
rect 2261 12364 2313 12368
rect 2326 12364 2378 12368
rect 2390 12364 2442 12368
rect 2454 12364 2506 12368
rect 2131 12330 2156 12364
rect 2156 12330 2183 12364
rect 2196 12330 2230 12364
rect 2230 12330 2248 12364
rect 2261 12330 2264 12364
rect 2264 12330 2304 12364
rect 2304 12330 2313 12364
rect 2326 12330 2338 12364
rect 2338 12330 2378 12364
rect 2390 12330 2412 12364
rect 2412 12330 2442 12364
rect 2454 12330 2486 12364
rect 2486 12330 2506 12364
rect 2131 12316 2183 12330
rect 2196 12316 2248 12330
rect 2261 12316 2313 12330
rect 2326 12316 2378 12330
rect 2390 12316 2442 12330
rect 2454 12316 2506 12330
rect 2518 12364 2570 12368
rect 2518 12330 2526 12364
rect 2526 12330 2560 12364
rect 2560 12330 2570 12364
rect 2518 12316 2570 12330
rect 2582 12364 2634 12368
rect 2582 12330 2600 12364
rect 2600 12330 2634 12364
rect 4041 12330 4077 12363
rect 4077 12330 4093 12363
rect 4127 12330 4150 12363
rect 4150 12330 4179 12363
rect 4213 12330 4223 12363
rect 4223 12330 4257 12363
rect 4257 12330 4265 12363
rect 2582 12316 2634 12330
rect 4041 12311 4093 12330
rect 4127 12311 4179 12330
rect 4213 12311 4265 12330
rect 2066 12248 2082 12254
rect 2082 12248 2116 12254
rect 2116 12248 2118 12254
rect 2066 12202 2118 12248
rect 2131 12248 2156 12254
rect 2156 12248 2183 12254
rect 2196 12248 2230 12254
rect 2230 12248 2248 12254
rect 2261 12248 2264 12254
rect 2264 12248 2304 12254
rect 2304 12248 2313 12254
rect 2326 12248 2338 12254
rect 2338 12248 2378 12254
rect 2390 12248 2412 12254
rect 2412 12248 2442 12254
rect 2454 12248 2486 12254
rect 2486 12248 2506 12254
rect 2131 12202 2183 12248
rect 2196 12202 2248 12248
rect 2261 12202 2313 12248
rect 2326 12202 2378 12248
rect 2390 12202 2442 12248
rect 2454 12202 2506 12248
rect 2518 12248 2526 12254
rect 2526 12248 2560 12254
rect 2560 12248 2570 12254
rect 2518 12202 2570 12248
rect 2582 12248 2600 12254
rect 2600 12248 2634 12254
rect 4041 12248 4077 12261
rect 4077 12248 4093 12261
rect 4127 12248 4150 12261
rect 4150 12248 4179 12261
rect 4213 12248 4223 12261
rect 4223 12248 4257 12261
rect 4257 12248 4265 12261
rect 2582 12202 2634 12248
rect 4041 12209 4093 12248
rect 4127 12209 4179 12248
rect 4213 12209 4265 12248
rect 4041 12118 4093 12159
rect 4127 12118 4179 12159
rect 4213 12118 4265 12159
rect 4041 12107 4077 12118
rect 4077 12107 4093 12118
rect 4127 12107 4150 12118
rect 4150 12107 4179 12118
rect 4213 12107 4223 12118
rect 4223 12107 4257 12118
rect 4257 12107 4265 12118
rect 4041 12036 4093 12056
rect 4127 12036 4179 12056
rect 4213 12036 4265 12056
rect 4041 12004 4077 12036
rect 4077 12004 4093 12036
rect 4127 12004 4150 12036
rect 4150 12004 4179 12036
rect 4213 12004 4223 12036
rect 4223 12004 4257 12036
rect 4257 12004 4265 12036
rect 2913 10728 2965 10780
rect 16754 10728 16806 10780
rect 16754 10664 16806 10716
rect 6961 10418 7013 10470
rect 7025 10418 7077 10470
rect 9386 10418 9438 10470
rect 9450 10418 9502 10470
rect 5583 10252 5635 10304
rect 5583 10188 5635 10240
rect 6079 10178 6131 10230
rect 6143 10178 6195 10230
rect 87 10144 139 10150
rect 151 10144 203 10150
rect 215 10144 267 10150
rect 279 10144 331 10150
rect -29 10110 -17 10122
rect -17 10110 17 10122
rect 17 10110 23 10122
rect 87 10110 90 10144
rect 90 10110 129 10144
rect 129 10110 139 10144
rect 151 10110 163 10144
rect 163 10110 202 10144
rect 202 10110 203 10144
rect 215 10110 236 10144
rect 236 10110 267 10144
rect 279 10110 309 10144
rect 309 10110 331 10144
rect -29 10072 23 10110
rect 87 10098 139 10110
rect 151 10098 203 10110
rect 215 10098 267 10110
rect 279 10098 331 10110
rect 343 10144 395 10150
rect 343 10110 348 10144
rect 348 10110 382 10144
rect 382 10110 395 10144
rect 343 10098 395 10110
rect 407 10144 459 10150
rect 407 10110 421 10144
rect 421 10110 455 10144
rect 455 10110 459 10144
rect 407 10098 459 10110
rect 471 10144 523 10150
rect 1427 10144 1479 10150
rect 471 10110 494 10144
rect 494 10110 523 10144
rect 1427 10110 1443 10144
rect 1443 10110 1477 10144
rect 1477 10110 1479 10144
rect 471 10098 523 10110
rect 1427 10098 1479 10110
rect 1491 10144 1543 10150
rect 1555 10144 1607 10150
rect 1619 10144 1671 10150
rect 1683 10144 1735 10150
rect 2247 10144 2299 10150
rect 1491 10110 1516 10144
rect 1516 10110 1543 10144
rect 1555 10110 1589 10144
rect 1589 10110 1607 10144
rect 1619 10110 1623 10144
rect 1623 10110 1662 10144
rect 1662 10110 1671 10144
rect 1683 10110 1696 10144
rect 1696 10110 1735 10144
rect 2247 10110 2280 10144
rect 2280 10110 2299 10144
rect 1491 10098 1543 10110
rect 1555 10098 1607 10110
rect 1619 10098 1671 10110
rect 1683 10098 1735 10110
rect 2247 10098 2299 10110
rect 2311 10144 2363 10150
rect 2311 10110 2319 10144
rect 2319 10110 2353 10144
rect 2353 10110 2363 10144
rect 2311 10098 2363 10110
rect 2375 10144 2427 10150
rect 2375 10110 2392 10144
rect 2392 10110 2426 10144
rect 2426 10110 2427 10144
rect 2375 10098 2427 10110
rect 2439 10144 2491 10150
rect 2503 10144 2555 10150
rect 2999 10144 3051 10150
rect 3063 10144 3115 10150
rect 3127 10144 3179 10150
rect 2439 10110 2465 10144
rect 2465 10110 2491 10144
rect 2503 10110 2538 10144
rect 2538 10110 2555 10144
rect 2999 10110 3010 10144
rect 3010 10110 3049 10144
rect 3049 10110 3051 10144
rect 3063 10110 3083 10144
rect 3083 10110 3115 10144
rect 3127 10110 3156 10144
rect 3156 10110 3179 10144
rect 2439 10098 2491 10110
rect 2503 10098 2555 10110
rect 2999 10098 3051 10110
rect 3063 10098 3115 10110
rect 3127 10098 3179 10110
rect 3191 10144 3243 10150
rect 3191 10110 3195 10144
rect 3195 10110 3229 10144
rect 3229 10110 3243 10144
rect 3191 10098 3243 10110
rect 3255 10144 3307 10150
rect 7645 10144 7697 10150
rect 7709 10144 7761 10150
rect 7773 10144 7825 10150
rect 7837 10144 7889 10150
rect 7901 10144 7953 10150
rect 7965 10144 8017 10150
rect 3255 10110 3268 10144
rect 3268 10110 3302 10144
rect 3302 10110 3307 10144
rect 7645 10110 7672 10144
rect 7672 10110 7697 10144
rect 7709 10110 7744 10144
rect 7744 10110 7761 10144
rect 7773 10110 7778 10144
rect 7778 10110 7816 10144
rect 7816 10110 7825 10144
rect 7837 10110 7850 10144
rect 7850 10110 7888 10144
rect 7888 10110 7889 10144
rect 7901 10110 7922 10144
rect 7922 10110 7953 10144
rect 7965 10110 7994 10144
rect 7994 10110 8017 10144
rect 3255 10098 3307 10110
rect 7645 10098 7697 10110
rect 7709 10098 7761 10110
rect 7773 10098 7825 10110
rect 7837 10098 7889 10110
rect 7901 10098 7953 10110
rect 7965 10098 8017 10110
rect 8029 10144 8081 10150
rect 8029 10110 8032 10144
rect 8032 10110 8066 10144
rect 8066 10110 8081 10144
rect 8029 10098 8081 10110
rect -29 10070 -17 10072
rect -17 10070 17 10072
rect 17 10070 23 10072
rect -29 10038 -17 10058
rect -17 10038 17 10058
rect 17 10038 23 10058
rect -29 10006 23 10038
rect -29 9993 23 9994
rect -29 9959 -17 9993
rect -17 9959 17 9993
rect 17 9959 23 9993
rect -29 9942 23 9959
rect -29 9915 23 9930
rect -29 9881 -17 9915
rect -17 9881 17 9915
rect 17 9881 23 9915
rect -29 9878 23 9881
rect 1881 9711 1997 9827
rect 14841 9715 15021 9831
rect 8247 9411 8299 9463
rect 8311 9411 8363 9463
rect 9306 9411 9358 9463
rect 9370 9411 9422 9463
rect 9989 9375 10041 9427
rect 10053 9375 10105 9427
rect 6961 9299 7013 9351
rect 7025 9299 7077 9351
rect 1881 9001 1997 9181
rect 13458 9062 13510 9114
rect 13458 8998 13510 9050
rect 16494 8674 16546 8726
rect 16494 8610 16546 8662
rect 16586 8560 16638 8612
rect 16586 8496 16638 8548
rect 16684 8441 16736 8493
rect 16748 8441 16800 8493
rect 7005 8365 7057 8417
rect 7005 8301 7057 8353
rect 9890 8286 9942 8338
rect 9954 8286 10006 8338
rect 13851 8144 13903 8196
rect 13921 8144 13973 8196
rect 13990 8144 14042 8196
rect 14059 8144 14111 8196
rect 14128 8144 14180 8196
rect 14197 8144 14249 8196
rect 14266 8144 14318 8196
rect 14335 8144 14387 8196
rect 14404 8144 14456 8196
rect 13851 8080 13903 8132
rect 13921 8080 13973 8132
rect 13990 8080 14042 8132
rect 14059 8080 14111 8132
rect 14128 8080 14180 8132
rect 14197 8080 14249 8132
rect 14266 8080 14318 8132
rect 14335 8080 14387 8132
rect 14404 8080 14456 8132
rect 13305 7893 13357 7945
rect 13369 7893 13421 7945
rect 10575 7805 10627 7857
rect 10639 7805 10691 7857
rect 6239 7748 6291 7800
rect 7005 7748 7057 7800
rect 2913 7667 2965 7719
rect 6239 7684 6291 7736
rect 7005 7684 7057 7736
rect 2913 7603 2965 7655
rect 12015 7663 12067 7715
rect 16407 7663 16459 7715
rect 4806 7597 4858 7649
rect 4870 7597 4922 7649
rect 12015 7599 12067 7651
rect 16407 7599 16459 7651
rect 13851 7506 13903 7558
rect 13921 7506 13973 7558
rect 13990 7506 14042 7558
rect 14059 7506 14111 7558
rect 14128 7506 14180 7558
rect 14197 7506 14249 7558
rect 14266 7506 14318 7558
rect 14335 7506 14387 7558
rect 14404 7506 14456 7558
rect 13851 7442 13903 7494
rect 13921 7442 13973 7494
rect 13990 7442 14042 7494
rect 14059 7442 14111 7494
rect 14128 7442 14180 7494
rect 14197 7442 14249 7494
rect 14266 7442 14318 7494
rect 14335 7442 14387 7494
rect 14404 7442 14456 7494
rect 9890 7355 9942 7407
rect 9954 7355 10006 7407
rect 16225 7351 16277 7403
rect 677 7222 729 7274
rect 6175 7228 6227 7280
rect 6239 7228 6291 7280
rect 10499 7226 10551 7278
rect 10563 7226 10615 7278
rect 12257 7275 12309 7327
rect 12321 7275 12373 7327
rect 16225 7287 16277 7339
rect 16407 7271 16459 7323
rect 677 7158 729 7210
rect 16407 7207 16459 7259
rect 16407 7103 16459 7155
rect 16407 7039 16459 7091
rect 10466 6839 10582 7019
rect 14832 6878 15012 6994
rect 23171 6914 23223 6966
rect 23171 6850 23223 6902
rect 1826 6684 1878 6736
rect 1890 6684 1942 6736
rect 5814 6702 5866 6754
rect 5878 6702 5930 6754
rect 16035 6727 16087 6779
rect 16035 6663 16087 6715
rect 15949 6556 16001 6608
rect 5681 6451 5733 6503
rect 5681 6387 5733 6439
rect 5681 6323 5733 6375
rect 5975 6451 6027 6503
rect 15949 6492 16001 6544
rect 5975 6387 6027 6439
rect 5975 6323 6027 6375
rect 1284 6134 1336 6186
rect 1284 6070 1336 6122
rect 8292 6048 8344 6100
rect 2246 5984 2298 6036
rect 2310 5984 2362 6036
rect 8292 5984 8344 6036
rect 12171 5972 12223 6024
rect 2788 5824 2840 5876
rect 12015 5908 12067 5960
rect 12171 5908 12223 5960
rect 12015 5844 12067 5896
rect 16225 5854 16277 5906
rect 926 5748 978 5800
rect 2788 5760 2840 5812
rect 16225 5790 16277 5842
rect 926 5684 978 5736
rect 12678 5152 12730 5204
rect 12742 5152 12794 5204
rect 12806 5152 12858 5204
rect 15714 5164 15766 5180
rect 15786 5164 15838 5180
rect 15858 5164 15910 5180
rect 15714 5130 15738 5164
rect 15738 5130 15766 5164
rect 15786 5130 15814 5164
rect 15814 5130 15838 5164
rect 15858 5130 15890 5164
rect 15890 5130 15910 5164
rect 15714 5128 15766 5130
rect 15786 5128 15838 5130
rect 15858 5128 15910 5130
rect 15930 5164 15982 5180
rect 15930 5130 15932 5164
rect 15932 5130 15966 5164
rect 15966 5130 15982 5164
rect 15930 5128 15982 5130
rect 16002 5164 16054 5180
rect 16002 5130 16008 5164
rect 16008 5130 16042 5164
rect 16042 5130 16054 5164
rect 16002 5128 16054 5130
rect 15714 5092 15766 5101
rect 15786 5092 15838 5101
rect 15858 5092 15910 5101
rect 15714 5058 15738 5092
rect 15738 5058 15766 5092
rect 15786 5058 15814 5092
rect 15814 5058 15838 5092
rect 15858 5058 15890 5092
rect 15890 5058 15910 5092
rect 15714 5049 15766 5058
rect 15786 5049 15838 5058
rect 15858 5049 15910 5058
rect 15930 5092 15982 5101
rect 15930 5058 15932 5092
rect 15932 5058 15966 5092
rect 15966 5058 15982 5092
rect 15930 5049 15982 5058
rect 16002 5092 16054 5101
rect 16002 5058 16008 5092
rect 16008 5058 16042 5092
rect 16042 5058 16054 5092
rect 16002 5049 16054 5058
rect 15714 5020 15766 5021
rect 15786 5020 15838 5021
rect 15858 5020 15910 5021
rect 15714 4986 15738 5020
rect 15738 4986 15766 5020
rect 15786 4986 15814 5020
rect 15814 4986 15838 5020
rect 15858 4986 15890 5020
rect 15890 4986 15910 5020
rect 15714 4969 15766 4986
rect 15786 4969 15838 4986
rect 15858 4969 15910 4986
rect 15930 5020 15982 5021
rect 15930 4986 15932 5020
rect 15932 4986 15966 5020
rect 15966 4986 15982 5020
rect 15930 4969 15982 4986
rect 16002 5020 16054 5021
rect 16002 4986 16008 5020
rect 16008 4986 16042 5020
rect 16042 4986 16054 5020
rect 16002 4969 16054 4986
rect 1890 4832 1942 4884
rect 1890 4768 1942 4820
rect 3548 4818 3600 4870
rect 3612 4818 3664 4870
rect 12015 4758 12067 4810
rect 12015 4694 12067 4746
rect 123 4480 239 4660
rect 10466 4473 10582 4653
rect 2236 4214 2288 4266
rect 2236 4150 2288 4202
rect 12257 4140 12309 4192
rect 12321 4140 12373 4192
rect 410 3969 526 4085
rect 4248 3809 4300 3861
rect 4312 3809 4364 3861
rect 54 3714 106 3766
rect 54 3650 106 3702
rect 7341 3619 7393 3671
rect 7405 3619 7457 3671
rect 17240 3602 17292 3654
rect 17304 3602 17356 3654
rect 4248 3539 4300 3591
rect 4312 3539 4364 3591
rect 4376 3539 4428 3591
rect 4440 3539 4492 3591
rect 11247 3539 11299 3591
rect 11311 3539 11363 3591
rect 410 3321 526 3501
rect 7178 3320 7294 3500
rect 19772 3447 19824 3499
rect 19841 3447 19893 3499
rect 19910 3447 19962 3499
rect 19979 3447 20031 3499
rect 20048 3447 20100 3499
rect 20117 3447 20169 3499
rect 20186 3447 20238 3499
rect 20255 3447 20307 3499
rect 20323 3447 20375 3499
rect 20391 3447 20443 3499
rect 20459 3447 20511 3499
rect 20527 3447 20579 3499
rect 12185 3379 12237 3431
rect 12185 3315 12237 3367
rect 19772 3383 19824 3435
rect 19841 3383 19893 3435
rect 19910 3383 19962 3435
rect 19979 3383 20031 3435
rect 20048 3383 20100 3435
rect 20117 3383 20169 3435
rect 20186 3383 20238 3435
rect 20255 3383 20307 3435
rect 20323 3383 20375 3435
rect 20391 3383 20443 3435
rect 20459 3383 20511 3435
rect 20527 3383 20579 3435
rect 21162 3389 21342 3505
rect 19772 3319 19824 3371
rect 19841 3319 19893 3371
rect 19910 3319 19962 3371
rect 19979 3319 20031 3371
rect 20048 3319 20100 3371
rect 20117 3319 20169 3371
rect 20186 3319 20238 3371
rect 20255 3319 20307 3371
rect 20323 3319 20375 3371
rect 20391 3319 20443 3371
rect 20459 3319 20511 3371
rect 20527 3319 20579 3371
rect 2003 3223 2055 3275
rect 2003 3159 2055 3211
rect 54 3044 106 3096
rect 54 2980 106 3032
rect 1364 3044 1416 3096
rect 1364 2980 1416 3032
rect 12185 2975 12237 3027
rect 7020 2906 7072 2958
rect 7084 2906 7136 2958
rect 12185 2911 12237 2963
rect 20675 2660 20727 2712
rect 20739 2660 20791 2712
rect 20803 2660 20855 2712
rect 20867 2660 20919 2712
rect 132 2519 312 2635
rect 1012 2584 1064 2636
rect 1101 2584 1153 2636
rect 1190 2584 1242 2636
rect 1278 2584 1330 2636
rect 1012 2518 1064 2570
rect 1101 2518 1153 2570
rect 1190 2518 1242 2570
rect 1278 2518 1330 2570
rect 2402 2519 2518 2635
rect 3628 2438 3680 2490
rect 3692 2438 3744 2490
rect 5578 2438 5630 2490
rect 5642 2438 5694 2490
rect 7546 2402 7598 2416
rect 7546 2368 7552 2402
rect 7552 2368 7586 2402
rect 7586 2368 7598 2402
rect 7546 2364 7598 2368
rect 7610 2402 7662 2416
rect 7610 2368 7624 2402
rect 7624 2368 7658 2402
rect 7658 2368 7662 2402
rect 7610 2364 7662 2368
rect 12413 2364 12465 2416
rect 12477 2364 12529 2416
rect 12541 2364 12593 2416
rect 12605 2364 12657 2416
rect 12669 2364 12721 2416
rect 12733 2364 12785 2416
rect 12797 2364 12849 2416
rect 16407 2268 16459 2320
rect 16407 2204 16459 2256
rect 20657 1980 20709 2032
rect 20730 1980 20782 2032
rect 20803 1980 20855 2032
rect 20875 1980 20927 2032
rect 20657 1916 20709 1968
rect 20730 1916 20782 1968
rect 20803 1916 20855 1968
rect 20875 1916 20927 1968
rect 20657 1852 20709 1904
rect 20730 1852 20782 1904
rect 20803 1852 20855 1904
rect 20875 1852 20927 1904
<< metal2 >>
rect 2077 13600 2597 13606
rect 2077 13548 2080 13600
rect 2132 13548 2146 13600
rect 2198 13548 2212 13600
rect 2264 13548 2278 13600
rect 2330 13548 2344 13600
rect 2396 13548 2410 13600
rect 2462 13548 2476 13600
rect 2528 13548 2542 13600
rect 2594 13548 2597 13600
rect 2077 13536 2597 13548
rect 2077 13484 2080 13536
rect 2132 13484 2146 13536
rect 2198 13484 2212 13536
rect 2264 13484 2278 13536
rect 2330 13484 2344 13536
rect 2396 13484 2410 13536
rect 2462 13484 2476 13536
rect 2528 13484 2542 13536
rect 2594 13484 2597 13536
rect 2077 13472 2597 13484
rect 2077 13420 2080 13472
rect 2132 13420 2146 13472
rect 2198 13420 2212 13472
rect 2264 13420 2278 13472
rect 2330 13420 2344 13472
rect 2396 13420 2410 13472
rect 2462 13420 2476 13472
rect 2528 13420 2542 13472
rect 2594 13420 2597 13472
rect 2077 13408 2597 13420
rect 2077 13356 2080 13408
rect 2132 13356 2146 13408
rect 2198 13356 2212 13408
rect 2264 13356 2278 13408
rect 2330 13356 2344 13408
rect 2396 13356 2410 13408
rect 2462 13356 2476 13408
rect 2528 13356 2542 13408
rect 2594 13356 2597 13408
rect 2077 13344 2597 13356
rect 2077 13292 2080 13344
rect 2132 13292 2146 13344
rect 2198 13292 2212 13344
rect 2264 13292 2278 13344
rect 2330 13292 2344 13344
rect 2396 13292 2410 13344
rect 2462 13292 2476 13344
rect 2528 13292 2542 13344
rect 2594 13292 2597 13344
rect 2077 13280 2597 13292
rect 2077 13228 2080 13280
rect 2132 13228 2146 13280
rect 2198 13228 2212 13280
rect 2264 13228 2278 13280
rect 2330 13228 2344 13280
rect 2396 13228 2410 13280
rect 2462 13228 2476 13280
rect 2528 13228 2542 13280
rect 2594 13228 2597 13280
rect 2077 13215 2597 13228
rect 2077 13163 2080 13215
rect 2132 13163 2146 13215
rect 2198 13163 2212 13215
rect 2264 13163 2278 13215
rect 2330 13163 2344 13215
rect 2396 13163 2410 13215
rect 2462 13163 2476 13215
rect 2528 13163 2542 13215
rect 2594 13163 2597 13215
rect 2077 13150 2597 13163
rect 2077 13098 2080 13150
rect 2132 13098 2146 13150
rect 2198 13098 2212 13150
rect 2264 13098 2278 13150
rect 2330 13098 2344 13150
rect 2396 13098 2410 13150
rect 2462 13098 2476 13150
rect 2528 13098 2542 13150
rect 2594 13098 2597 13150
rect 2077 13085 2597 13098
rect 2077 13033 2080 13085
rect 2132 13033 2146 13085
rect 2198 13033 2212 13085
rect 2264 13033 2278 13085
rect 2330 13033 2344 13085
rect 2396 13033 2410 13085
rect 2462 13033 2476 13085
rect 2528 13033 2542 13085
rect 2594 13033 2597 13085
rect 2077 13020 2597 13033
rect 2077 12968 2080 13020
rect 2132 12968 2146 13020
rect 2198 12968 2212 13020
rect 2264 12968 2278 13020
rect 2330 12968 2344 13020
rect 2396 12968 2410 13020
rect 2462 12968 2476 13020
rect 2528 12968 2542 13020
rect 2594 12968 2597 13020
rect 2077 12955 2597 12968
rect 2077 12903 2080 12955
rect 2132 12903 2146 12955
rect 2198 12903 2212 12955
rect 2264 12903 2278 12955
rect 2330 12903 2344 12955
rect 2396 12903 2410 12955
rect 2462 12903 2476 12955
rect 2528 12903 2542 12955
rect 2594 12903 2597 12955
rect 2077 12897 2597 12903
rect 2060 12316 2066 12368
rect 2118 12316 2131 12368
rect 2183 12316 2196 12368
rect 2248 12316 2261 12368
rect 2313 12316 2326 12368
rect 2378 12316 2390 12368
rect 2442 12316 2454 12368
rect 2506 12316 2518 12368
rect 2570 12316 2582 12368
rect 2634 12316 2640 12368
rect 2060 12254 2640 12316
rect 2060 12202 2066 12254
rect 2118 12202 2131 12254
rect 2183 12202 2196 12254
rect 2248 12202 2261 12254
rect 2313 12202 2326 12254
rect 2378 12202 2390 12254
rect 2442 12202 2454 12254
rect 2506 12202 2518 12254
rect 2570 12202 2582 12254
rect 2634 12202 2640 12254
rect 4041 12363 4265 12369
rect 4093 12311 4127 12363
rect 4179 12311 4213 12363
rect 4041 12261 4265 12311
rect 4093 12209 4127 12261
rect 4179 12209 4213 12261
rect 4041 12159 4265 12209
rect 4093 12107 4127 12159
rect 4179 12107 4213 12159
rect 4041 12056 4265 12107
rect 4093 12004 4127 12056
rect 4179 12004 4213 12056
rect 4041 11998 4265 12004
rect 1837 11671 2145 11836
tri 1837 11483 2025 11671 ne
rect 1881 11404 1997 11421
rect 1881 11348 1911 11404
rect 1967 11348 1997 11404
rect 1881 11324 1997 11348
rect 1881 11268 1911 11324
rect 1967 11268 1997 11324
rect 1881 11244 1997 11268
rect 1881 11188 1911 11244
rect 1967 11188 1997 11244
rect 1881 11163 1997 11188
rect -71 10150 529 10818
rect -71 10122 87 10150
rect -71 10070 -29 10122
rect 23 10098 87 10122
rect 139 10098 151 10150
rect 203 10098 215 10150
rect 267 10098 279 10150
rect 331 10098 343 10150
rect 395 10098 407 10150
rect 459 10098 471 10150
rect 523 10098 529 10150
rect 23 10070 529 10098
rect -71 10058 529 10070
rect -71 10006 -29 10058
rect 23 10006 529 10058
rect -71 9994 529 10006
rect -71 9942 -29 9994
rect 23 9942 529 9994
rect -71 9930 529 9942
rect -71 9878 -29 9930
rect 23 9878 529 9930
rect -71 5374 529 9878
rect 799 10562 1365 10818
rect 799 10506 861 10562
rect 917 10506 941 10562
rect 997 10506 1365 10562
rect 799 10481 1365 10506
rect 799 10425 861 10481
rect 917 10425 941 10481
rect 997 10425 1365 10481
rect 799 10400 1365 10425
rect 799 10344 861 10400
rect 917 10344 941 10400
rect 997 10344 1365 10400
rect 799 10319 1365 10344
rect 799 10263 861 10319
rect 917 10263 941 10319
rect 997 10263 1365 10319
rect 799 10238 1365 10263
rect 799 10182 861 10238
rect 917 10182 941 10238
rect 997 10182 1365 10238
rect 799 10157 1365 10182
rect 799 10101 861 10157
rect 917 10101 941 10157
rect 997 10101 1365 10157
rect 799 10076 1365 10101
rect 799 10020 861 10076
rect 917 10020 941 10076
rect 997 10020 1365 10076
rect 799 9995 1365 10020
rect 799 9939 861 9995
rect 917 9939 941 9995
rect 997 9939 1365 9995
rect 799 9914 1365 9939
rect 799 9858 861 9914
rect 917 9858 941 9914
rect 997 9858 1365 9914
rect 799 9832 1365 9858
rect 799 9776 861 9832
rect 917 9776 941 9832
rect 997 9776 1365 9832
rect 799 9750 1365 9776
rect 799 9694 861 9750
rect 917 9694 941 9750
rect 997 9694 1365 9750
rect 1421 10150 1741 11132
rect 1421 10098 1427 10150
rect 1479 10098 1491 10150
rect 1543 10098 1555 10150
rect 1607 10098 1619 10150
rect 1671 10098 1683 10150
rect 1735 10098 1741 10150
rect 1421 9709 1741 10098
rect 1881 11107 1911 11163
rect 1967 11107 1997 11163
rect 1881 9827 1997 11107
rect 1881 9705 1997 9711
tri 1881 9704 1882 9705 ne
rect 799 9668 1365 9694
rect 799 9612 861 9668
rect 917 9612 941 9668
rect 997 9612 1365 9668
rect 799 9586 1365 9612
rect 799 9535 861 9586
tri 799 9497 837 9535 ne
rect 837 9530 861 9535
rect 917 9530 941 9586
rect 997 9530 1365 9586
rect 837 9504 1365 9530
rect 837 9448 861 9504
rect 917 9448 941 9504
rect 997 9448 1365 9504
rect 837 9422 1365 9448
rect 837 9366 861 9422
rect 917 9366 941 9422
rect 997 9366 1365 9422
rect 837 9340 1365 9366
rect 837 9284 861 9340
rect 917 9284 941 9340
rect 997 9284 1365 9340
rect 837 9258 1365 9284
rect 837 9202 861 9258
rect 917 9202 941 9258
rect 997 9202 1365 9258
rect 837 9176 1365 9202
rect 837 9120 861 9176
rect 917 9120 941 9176
rect 997 9120 1365 9176
rect 837 9094 1365 9120
rect 837 9038 861 9094
rect 917 9038 941 9094
rect 997 9038 1365 9094
rect 837 9012 1365 9038
rect 837 8956 861 9012
rect 917 8956 941 9012
rect 997 8956 1365 9012
tri 1881 9187 1882 9188 se
rect 1882 9187 1997 9705
rect 1881 9181 1997 9187
rect 1881 8995 1997 9001
rect 837 8930 1365 8956
rect 837 8874 861 8930
rect 917 8874 941 8930
rect 997 8874 1365 8930
rect 837 8848 1365 8874
rect 837 8792 861 8848
rect 917 8792 941 8848
rect 997 8792 1365 8848
rect 837 8766 1365 8792
rect 837 8710 861 8766
rect 917 8710 941 8766
rect 997 8710 1365 8766
rect 837 8684 1365 8710
rect 837 8628 861 8684
rect 917 8628 941 8684
rect 997 8628 1365 8684
rect 837 8602 1365 8628
rect 837 8546 861 8602
rect 917 8546 941 8602
rect 997 8546 1365 8602
rect 837 8520 1365 8546
rect 837 8464 861 8520
rect 917 8464 941 8520
rect 997 8464 1365 8520
rect 837 8438 1365 8464
rect 837 8382 861 8438
rect 917 8382 941 8438
rect 997 8382 1365 8438
rect 837 8356 1365 8382
rect 837 8300 861 8356
rect 917 8300 941 8356
rect 997 8300 1365 8356
rect 837 8274 1365 8300
rect 837 8218 861 8274
rect 917 8218 941 8274
rect 997 8218 1365 8274
rect 837 8192 1365 8218
rect 837 8136 861 8192
rect 917 8136 941 8192
rect 997 8136 1365 8192
rect 837 8110 1365 8136
rect 837 8054 861 8110
rect 917 8054 941 8110
rect 997 8054 1365 8110
rect 837 8028 1365 8054
rect 837 7972 861 8028
rect 917 7972 941 8028
rect 997 7972 1365 8028
rect 837 7946 1365 7972
rect 837 7890 861 7946
rect 917 7890 941 7946
rect 997 7890 1365 7946
rect 837 7864 1365 7890
rect 837 7808 861 7864
rect 917 7808 941 7864
rect 997 7808 1365 7864
rect 677 7274 729 7280
rect 677 7210 729 7222
rect 677 7152 729 7158
rect 837 6319 1365 7808
rect 1789 6839 1836 6860
tri 1836 6839 1857 6860 nw
tri 1789 6792 1836 6839 nw
rect 1820 6684 1826 6736
rect 1878 6684 1890 6736
rect 1942 6684 1948 6736
tri 1859 6663 1880 6684 ne
rect 1880 6663 1948 6684
tri 1880 6659 1884 6663 ne
rect 1745 6556 1789 6592
tri 1789 6556 1825 6592 sw
rect 1745 6544 1825 6556
tri 1825 6544 1837 6556 sw
rect 1745 6525 1837 6544
tri 1837 6525 1856 6544 sw
rect 1284 6186 1336 6192
rect 1284 6122 1336 6134
rect -71 5268 423 5374
tri 423 5268 529 5374 nw
rect 926 5800 978 5806
rect 926 5736 978 5748
rect -71 5204 359 5268
tri 359 5204 423 5268 nw
rect -71 5152 307 5204
tri 307 5152 359 5204 nw
rect -71 5128 283 5152
tri 283 5128 307 5152 nw
rect -71 4660 267 5128
tri 267 5112 283 5128 nw
rect -71 4480 123 4660
rect 239 4480 267 4660
tri 513 4150 530 4167 se
tri 507 4144 513 4150 se
rect 513 4144 530 4150
tri 503 4140 507 4144 se
rect 507 4140 530 4144
tri 454 4091 503 4140 se
rect 503 4091 530 4140
rect 346 4085 658 4091
rect 346 3969 410 4085
rect 526 3969 658 4085
rect 54 3766 106 3772
rect 54 3702 106 3714
rect 54 3096 106 3650
rect 54 3032 106 3044
rect 54 2974 106 2980
rect 346 3501 658 3969
rect 346 3321 410 3501
rect 526 3321 658 3501
rect 346 3315 658 3321
rect 346 3314 657 3315
tri 657 3314 658 3315 nw
rect 346 3281 624 3314
tri 624 3281 657 3314 nw
rect 346 3275 618 3281
tri 618 3275 624 3281 nw
rect 126 2519 132 2635
rect 312 2519 318 2635
rect 126 2137 318 2519
rect 346 2321 582 3275
tri 582 3239 618 3275 nw
rect 926 2321 978 5684
rect 1284 4257 1336 6070
rect 1745 6058 1856 6525
rect 1473 5409 1856 6058
tri 1473 5282 1600 5409 ne
rect 1600 5282 1856 5409
rect 1444 5259 1572 5268
rect 1444 5203 1480 5259
rect 1536 5203 1572 5259
rect 1444 5173 1572 5203
rect 1444 5117 1480 5173
rect 1536 5117 1572 5173
rect 1444 5087 1572 5117
rect 1444 5031 1480 5087
rect 1536 5031 1572 5087
rect 1444 5001 1572 5031
rect 1444 4945 1480 5001
rect 1536 4945 1572 5001
rect 1444 4915 1572 4945
rect 1444 4859 1480 4915
rect 1536 4859 1572 4915
rect 1444 4828 1572 4859
rect 1444 4772 1480 4828
rect 1536 4772 1572 4828
rect 1444 4741 1572 4772
rect 1884 4884 1948 6663
rect 2025 6048 2145 11671
rect 2241 10150 2561 11132
rect 2241 10098 2247 10150
rect 2299 10098 2311 10150
rect 2363 10098 2375 10150
rect 2427 10098 2439 10150
rect 2491 10098 2503 10150
rect 2555 10098 2561 10150
rect 2241 6854 2561 10098
rect 2913 10780 2965 10786
rect 2913 7719 2965 10728
rect 2913 7655 2965 7667
rect 2913 7597 2965 7603
rect 2993 10150 3313 11132
rect 3537 10801 3937 11132
tri 5947 10847 6055 10955 se
rect 6055 10847 6455 11350
tri 3537 10780 3558 10801 ne
rect 3558 10786 3937 10801
tri 3937 10786 3998 10847 sw
tri 5886 10786 5947 10847 se
rect 5947 10786 6455 10847
tri 8470 11051 8551 11132 se
rect 8551 11051 8951 11132
rect 3558 10780 3998 10786
tri 3998 10780 4004 10786 sw
tri 5881 10781 5886 10786 se
rect 5886 10781 6455 10786
tri 5880 10780 5881 10781 se
rect 5881 10780 6455 10781
tri 6455 10780 6456 10781 sw
tri 3558 10759 3579 10780 ne
rect 3579 10759 4004 10780
tri 4004 10759 4025 10780 sw
tri 5866 10766 5880 10780 se
rect 5880 10766 6456 10780
tri 3579 10728 3610 10759 ne
rect 3610 10728 4025 10759
tri 5309 10728 5347 10766 se
rect 5347 10728 6456 10766
tri 6456 10728 6508 10780 sw
tri 3610 10716 3622 10728 ne
rect 3622 10716 4025 10728
tri 5297 10716 5309 10728 se
rect 5309 10716 6508 10728
tri 6508 10716 6520 10728 sw
tri 3622 10664 3674 10716 ne
rect 3674 10664 4025 10716
tri 5245 10664 5297 10716 se
rect 5297 10664 6520 10716
tri 6520 10664 6572 10716 sw
tri 3674 10658 3680 10664 ne
rect 3680 10658 4025 10664
tri 3680 10633 3705 10658 ne
rect 2993 10098 2999 10150
rect 3051 10098 3063 10150
rect 3115 10098 3127 10150
rect 3179 10098 3191 10150
rect 3243 10098 3255 10150
rect 3307 10098 3313 10150
tri 2561 6854 2716 7009 sw
rect 2241 6203 2716 6854
rect 2993 6864 3313 10098
tri 3313 6864 3346 6897 sw
rect 2993 6679 3346 6864
tri 2993 6663 3009 6679 ne
rect 3009 6663 3346 6679
tri 3009 6646 3026 6663 ne
tri 2241 6181 2263 6203 ne
rect 2263 6181 2716 6203
tri 2263 6107 2337 6181 ne
rect 2337 6107 2716 6181
tri 2337 6100 2344 6107 ne
rect 2344 6100 2716 6107
tri 2344 6093 2351 6100 ne
rect 2351 6093 2716 6100
tri 2145 6048 2190 6093 sw
tri 2351 6048 2396 6093 ne
rect 2025 6043 2190 6048
tri 2025 6036 2032 6043 ne
rect 2032 6036 2190 6043
tri 2190 6036 2202 6048 sw
tri 2032 6030 2038 6036 ne
rect 2038 6030 2202 6036
tri 2202 6030 2208 6036 sw
tri 2038 5984 2084 6030 ne
rect 2084 5984 2208 6030
rect 2240 5984 2246 6036
rect 2298 5984 2310 6036
rect 2362 5984 2368 6036
tri 2084 5980 2088 5984 ne
rect 1884 4832 1890 4884
rect 1942 4832 1948 4884
rect 1884 4820 1948 4832
rect 1884 4768 1890 4820
rect 1942 4768 1948 4820
rect 1444 4685 1480 4741
rect 1536 4685 1572 4741
rect 1444 4676 1572 4685
tri 1572 4430 1597 4455 sw
rect 1444 4310 1652 4430
tri 1575 4292 1593 4310 ne
rect 1593 4292 1600 4310
tri 1593 4285 1600 4292 ne
tri 1336 4257 1342 4263 sw
rect 1284 4241 1342 4257
tri 1284 4214 1311 4241 ne
rect 1311 4214 1342 4241
tri 1342 4214 1385 4257 sw
tri 1311 4202 1323 4214 ne
rect 1323 4202 1385 4214
tri 1385 4202 1397 4214 sw
tri 1323 4183 1342 4202 ne
rect 1342 4183 1397 4202
tri 1397 4183 1416 4202 sw
tri 1342 4167 1358 4183 ne
rect 1358 4167 1416 4183
tri 1358 4161 1364 4167 ne
rect 1006 4150 1322 4152
tri 1322 4150 1324 4152 sw
rect 1006 4144 1324 4150
tri 1324 4144 1330 4150 sw
rect 1006 4140 1330 4144
tri 1330 4140 1334 4144 sw
rect 1006 4138 1334 4140
tri 1334 4138 1336 4140 sw
rect 1006 2636 1336 4138
rect 1364 3636 1416 4167
tri 1416 3636 1422 3642 sw
rect 1364 3620 1422 3636
tri 1364 3619 1365 3620 ne
rect 1365 3619 1422 3620
tri 1422 3619 1439 3636 sw
tri 1365 3602 1382 3619 ne
rect 1382 3602 1439 3619
tri 1439 3602 1456 3619 sw
tri 1382 3591 1393 3602 ne
rect 1393 3591 1456 3602
tri 1456 3591 1467 3602 sw
tri 1393 3562 1422 3591 ne
rect 1422 3562 1467 3591
tri 1467 3562 1496 3591 sw
tri 1422 3540 1444 3562 ne
rect 1006 2584 1012 2636
rect 1064 2584 1101 2636
rect 1153 2584 1190 2636
rect 1242 2584 1278 2636
rect 1330 2584 1336 2636
rect 1006 2570 1336 2584
rect 1006 2518 1012 2570
rect 1064 2518 1101 2570
rect 1153 2518 1190 2570
rect 1242 2518 1278 2570
rect 1330 2518 1336 2570
rect 1006 2321 1336 2518
rect 1364 3096 1416 3102
rect 1364 3032 1416 3044
rect 1364 2321 1416 2980
rect 1444 2321 1496 3562
rect 2003 3275 2055 3281
rect 2003 3211 2055 3223
rect 2003 2336 2055 3159
rect 2088 2321 2208 5984
tri 2291 5972 2303 5984 ne
rect 2303 5972 2368 5984
tri 2303 5960 2315 5972 ne
rect 2315 5960 2368 5972
tri 2315 5959 2316 5960 ne
rect 2236 4266 2288 4272
rect 2236 4202 2288 4214
rect 2236 2321 2288 4150
rect 2316 2321 2368 5960
rect 2396 4464 2716 6093
rect 2788 5876 2840 5882
rect 2788 5812 2840 5824
tri 2755 2975 2788 3008 se
rect 2788 2986 2840 5760
rect 3026 4464 3346 6663
rect 3705 6314 4025 10658
tri 5158 10577 5245 10664 se
rect 5245 10658 6572 10664
tri 6572 10658 6578 10664 sw
rect 5245 10621 6578 10658
tri 6578 10621 6615 10658 sw
rect 5245 10587 6615 10621
tri 6615 10587 6649 10621 sw
rect 5245 10577 6649 10587
tri 4989 10549 5017 10577 se
rect 5017 10549 6649 10577
rect 4989 10545 6649 10549
tri 6649 10545 6691 10587 sw
rect 4989 10366 6691 10545
rect 4989 10310 5445 10366
tri 5445 10310 5501 10366 nw
tri 6207 10310 6263 10366 ne
rect 6263 10310 6691 10366
rect 4989 10304 5439 10310
tri 5439 10304 5445 10310 nw
rect 5583 10304 5635 10310
rect 4989 10252 5387 10304
tri 5387 10252 5439 10304 nw
rect 4989 10240 5375 10252
tri 5375 10240 5387 10252 nw
rect 5583 10240 5635 10252
rect 4073 5151 4593 10041
rect 4800 7597 4806 7649
rect 4858 7597 4870 7649
rect 4922 7597 4928 7649
tri 4851 7593 4855 7597 ne
rect 4855 7593 4928 7597
tri 4855 7572 4876 7593 ne
rect 4876 6279 4928 7593
rect 4989 6315 5359 10240
tri 5359 10224 5375 10240 nw
tri 6263 10230 6343 10310 ne
rect 6343 10230 6691 10310
rect 5583 9347 5635 10188
rect 6073 10178 6079 10230
rect 6131 10178 6143 10230
rect 6195 10178 6201 10230
tri 6343 10224 6349 10230 ne
rect 6073 9347 6125 10178
tri 6125 10153 6150 10178 nw
rect 6233 7748 6239 7800
rect 6291 7748 6297 7800
rect 6233 7736 6297 7748
rect 6233 7684 6239 7736
rect 6291 7684 6297 7736
rect 5675 6503 5739 7443
rect 5808 6702 5814 6754
rect 5866 6702 5878 6754
rect 5930 6702 5936 6754
tri 5859 6677 5884 6702 ne
rect 5675 6451 5681 6503
rect 5733 6451 5739 6503
rect 5675 6439 5739 6451
rect 5675 6387 5681 6439
rect 5733 6387 5739 6439
rect 5675 6375 5739 6387
rect 5675 6323 5681 6375
rect 5733 6323 5739 6375
tri 4876 6255 4900 6279 ne
rect 4900 6259 4928 6279
tri 4928 6259 4970 6301 sw
rect 4900 6255 4970 6259
tri 4970 6255 4974 6259 sw
tri 4900 6227 4928 6255 ne
rect 4928 6231 4974 6255
tri 4974 6231 4998 6255 sw
rect 4928 6227 4998 6231
tri 4928 6181 4974 6227 ne
rect 4974 6197 4998 6227
tri 4998 6197 5032 6231 sw
rect 4974 6181 5032 6197
tri 5032 6181 5048 6197 sw
tri 4974 6107 5048 6181 ne
tri 5048 6107 5122 6181 sw
tri 5048 6100 5055 6107 ne
rect 5055 6100 5122 6107
tri 5122 6100 5129 6107 sw
tri 5055 6048 5107 6100 ne
rect 5107 6048 5129 6100
tri 5129 6048 5181 6100 sw
tri 5107 6036 5119 6048 ne
rect 5119 6036 5181 6048
tri 5181 6036 5193 6048 sw
tri 5119 6033 5122 6036 ne
rect 5122 6033 5193 6036
tri 5193 6033 5196 6036 sw
tri 5122 5984 5171 6033 ne
rect 5171 5984 5196 6033
tri 5196 5984 5245 6033 sw
tri 5171 5972 5183 5984 ne
rect 5183 5972 5245 5984
tri 5245 5972 5257 5984 sw
tri 5183 5960 5195 5972 ne
rect 5195 5960 5257 5972
tri 5257 5960 5269 5972 sw
tri 5195 5959 5196 5960 ne
rect 5196 5959 5269 5960
tri 5269 5959 5270 5960 sw
tri 5196 5908 5247 5959 ne
rect 5247 5908 5270 5959
tri 5270 5908 5321 5959 sw
tri 5247 5906 5249 5908 ne
rect 5249 5906 5321 5908
tri 5321 5906 5323 5908 sw
tri 5249 5896 5259 5906 ne
rect 5259 5896 5323 5906
tri 5323 5896 5333 5906 sw
tri 5259 5885 5270 5896 ne
rect 5270 5885 5333 5896
tri 5333 5885 5344 5896 sw
tri 5270 5882 5273 5885 ne
rect 5273 5882 5344 5885
tri 5344 5882 5347 5885 sw
tri 5273 5844 5311 5882 ne
rect 5311 5844 5347 5882
tri 5347 5844 5385 5882 sw
tri 5311 5842 5313 5844 ne
rect 5313 5842 5385 5844
tri 5385 5842 5387 5844 sw
tri 5313 5811 5344 5842 ne
rect 5344 5811 5387 5842
tri 5387 5811 5418 5842 sw
tri 5344 5790 5365 5811 ne
rect 5365 5790 5418 5811
tri 5365 5789 5366 5790 ne
rect 4073 5128 4570 5151
tri 4570 5128 4593 5151 nw
rect 3542 4818 3548 4870
rect 3600 4818 3612 4870
rect 3664 4818 3670 4870
tri 3597 4810 3605 4818 ne
rect 3605 4810 3670 4818
tri 3605 4793 3622 4810 ne
rect 2788 2975 2829 2986
tri 2829 2975 2840 2986 nw
tri 2743 2963 2755 2975 se
rect 2755 2963 2817 2975
tri 2817 2963 2829 2975 nw
tri 2738 2958 2743 2963 se
rect 2743 2958 2812 2963
tri 2812 2958 2817 2963 nw
tri 2714 2934 2738 2958 se
rect 2738 2934 2788 2958
tri 2788 2934 2812 2958 nw
tri 2686 2906 2714 2934 se
rect 2714 2906 2760 2934
tri 2760 2906 2788 2934 nw
tri 2640 2860 2686 2906 se
rect 2686 2860 2714 2906
tri 2714 2860 2760 2906 nw
tri 2566 2786 2640 2860 se
tri 2640 2786 2714 2860 nw
tri 2552 2772 2566 2786 se
rect 2566 2772 2626 2786
tri 2626 2772 2640 2786 nw
rect 2396 2519 2402 2635
rect 2518 2519 2524 2635
rect 2396 2321 2524 2519
rect 2552 2321 2604 2772
tri 2604 2750 2626 2772 nw
rect 2872 2321 3192 4152
rect 3622 2497 3670 4810
rect 3698 4230 3814 4688
rect 4073 4385 4568 5128
tri 4568 5126 4570 5128 nw
tri 4073 4284 4174 4385 ne
tri 3698 4218 3710 4230 ne
rect 3710 4218 3814 4230
tri 3710 4192 3736 4218 ne
rect 3736 4192 3814 4218
tri 3736 4188 3740 4192 ne
rect 3740 4188 3814 4192
tri 3740 4144 3784 4188 ne
rect 3784 4144 3814 4188
tri 3814 4144 3858 4188 sw
tri 3784 4140 3788 4144 ne
rect 3788 4140 3858 4144
tri 3788 4122 3806 4140 ne
rect 3806 4091 3858 4140
rect 4174 4149 4568 4385
rect 4174 4140 4559 4149
tri 4559 4140 4568 4149 nw
rect 4174 4137 4556 4140
tri 4556 4137 4559 4140 nw
rect 4174 4109 4528 4137
tri 4528 4109 4556 4137 nw
tri 4568 4109 4596 4137 se
rect 4596 4123 4712 4688
rect 5366 4330 5418 5790
tri 5366 4292 5404 4330 ne
rect 5404 4292 5418 4330
tri 5418 4292 5478 4352 sw
tri 5404 4278 5418 4292 ne
rect 5418 4278 5478 4292
tri 5418 4272 5424 4278 ne
rect 5424 4272 5478 4278
tri 5478 4272 5498 4292 sw
tri 5424 4218 5478 4272 ne
rect 5478 4218 5498 4272
tri 5498 4218 5552 4272 sw
tri 5478 4192 5504 4218 ne
rect 5504 4192 5552 4218
tri 5552 4192 5578 4218 sw
tri 5504 4144 5552 4192 ne
rect 5552 4157 5578 4192
tri 5578 4157 5613 4192 sw
rect 5552 4144 5613 4157
tri 5613 4144 5626 4157 sw
tri 5552 4140 5556 4144 ne
rect 5556 4140 5626 4144
tri 5626 4140 5630 4144 sw
rect 4596 4109 4680 4123
rect 4174 3861 4522 4109
tri 4522 4103 4528 4109 nw
tri 4562 4103 4568 4109 se
rect 4568 4103 4680 4109
tri 4550 4091 4562 4103 se
rect 4562 4091 4680 4103
tri 4680 4091 4712 4123 nw
tri 5556 4091 5605 4140 ne
rect 5605 4113 5630 4140
tri 5630 4113 5657 4140 sw
rect 5605 4091 5657 4113
tri 5657 4091 5679 4113 sw
rect 4550 4070 4659 4091
tri 4659 4070 4680 4091 nw
tri 5605 4070 5626 4091 ne
rect 5626 4079 5679 4091
tri 5679 4079 5691 4091 sw
rect 5626 4070 5691 4079
tri 5691 4070 5700 4079 sw
rect 4550 4048 4637 4070
tri 4637 4048 4659 4070 nw
tri 5626 4048 5648 4070 ne
rect 4550 3963 4602 4048
tri 4602 4013 4637 4048 nw
rect 4174 3809 4248 3861
rect 4300 3809 4312 3861
rect 4364 3809 4522 3861
rect 4174 3591 4522 3809
rect 5648 3707 5700 4070
tri 5700 3707 5734 3741 sw
rect 5648 3655 5776 3707
rect 4174 3539 4248 3591
rect 4300 3539 4312 3591
rect 4364 3539 4376 3591
rect 4428 3539 4440 3591
rect 4492 3539 4522 3591
tri 3670 2497 3688 2515 sw
rect 3622 2490 3688 2497
tri 3688 2490 3695 2497 sw
rect 3622 2438 3628 2490
rect 3680 2438 3692 2490
rect 3744 2438 3750 2490
tri 3794 2438 3806 2450 se
rect 3806 2438 3858 3315
tri 4172 3165 4174 3167 se
rect 4174 3165 4522 3539
tri 4154 2906 4172 2924 se
rect 4172 2906 4522 3165
tri 3772 2416 3794 2438 se
rect 3794 2428 3858 2438
rect 3794 2416 3846 2428
tri 3846 2416 3858 2428 nw
tri 3981 2733 4154 2906 se
rect 4154 2733 4522 2906
rect 3981 2670 4522 2733
rect 3981 2660 4512 2670
tri 4512 2660 4522 2670 nw
rect 3981 2490 4342 2660
tri 4342 2490 4512 2660 nw
tri 3745 2389 3772 2416 se
rect 3772 2389 3819 2416
tri 3819 2389 3846 2416 nw
rect 3745 2382 3812 2389
tri 3812 2382 3819 2389 nw
rect 3745 2302 3797 2382
tri 3797 2367 3812 2382 nw
rect 3981 2302 4301 2490
tri 4301 2449 4342 2490 nw
rect 5572 2438 5578 2490
rect 5630 2438 5642 2490
rect 5694 2438 5700 2490
tri 5623 2416 5645 2438 ne
rect 5645 2416 5700 2438
tri 5645 2413 5648 2416 ne
rect 5648 2321 5700 2416
rect 5884 2321 5936 6702
rect 5969 6503 6033 7443
tri 6208 7280 6233 7305 se
rect 6233 7280 6297 7684
rect 6169 7228 6175 7280
rect 6227 7228 6239 7280
rect 6291 7228 6297 7280
rect 5969 6451 5975 6503
rect 6027 6451 6033 6503
rect 5969 6439 6033 6451
rect 5969 6387 5975 6439
rect 6027 6387 6033 6439
rect 5969 6375 6033 6387
rect 5969 6323 5975 6375
rect 6027 6323 6033 6375
rect 6349 6315 6691 10230
rect 6955 10418 6961 10470
rect 7013 10418 7025 10470
rect 7077 10418 7083 10470
rect 6955 9375 7007 10418
tri 7007 10393 7032 10418 nw
rect 7620 10150 8100 10815
tri 8205 10587 8239 10621 nw
rect 7620 10098 7645 10150
rect 7697 10098 7709 10150
rect 7761 10098 7773 10150
rect 7825 10098 7837 10150
rect 7889 10098 7901 10150
rect 7953 10098 7965 10150
rect 8017 10098 8029 10150
rect 8081 10098 8100 10150
tri 7007 9375 7008 9376 sw
rect 6955 9360 7008 9375
tri 7008 9360 7023 9375 sw
rect 6955 9351 7023 9360
tri 7023 9351 7032 9360 sw
rect 6955 9299 6961 9351
rect 7013 9299 7025 9351
rect 7077 9299 7083 9351
rect 6875 8821 6927 8873
rect 6999 8365 7005 8417
rect 7057 8365 7063 8417
rect 6999 8353 7063 8365
rect 6999 8301 7005 8353
rect 7057 8301 7063 8353
rect 6999 7800 7063 8301
rect 6999 7748 7005 7800
rect 7057 7748 7063 7800
rect 6999 7736 7063 7748
rect 6999 7684 7005 7736
rect 7057 7684 7063 7736
tri 7502 5616 7620 5734 se
rect 7620 5616 8100 10098
tri 8292 9463 8317 9488 se
rect 8317 9463 8369 10041
rect 8470 9760 8951 11051
rect 16754 10780 16806 10786
rect 16754 10716 16806 10728
rect 9380 10418 9386 10470
rect 9438 10418 9450 10470
rect 9502 10418 9508 10470
tri 9424 10386 9456 10418 ne
tri 9446 10041 9456 10051 se
rect 9456 10041 9508 10418
tri 8470 9715 8515 9760 ne
rect 8515 9715 8951 9760
tri 8515 9705 8525 9715 ne
rect 8525 9705 8951 9715
tri 8525 9676 8554 9705 ne
tri 8415 9513 8449 9547 nw
rect 8241 9411 8247 9463
rect 8299 9411 8311 9463
rect 8363 9411 8369 9463
tri 8545 9351 8554 9360 se
rect 8554 9351 8951 9705
rect 9300 9463 9352 10041
tri 9419 10014 9446 10041 se
rect 9446 10014 9508 10041
tri 9352 9463 9377 9488 sw
rect 9300 9411 9306 9463
rect 9358 9411 9370 9463
rect 9422 9411 9428 9463
rect 9983 9427 10111 10338
rect 9983 9375 9989 9427
rect 10041 9375 10053 9427
rect 10105 9375 10111 9427
tri 8493 9299 8545 9351 se
rect 8545 9299 8951 9351
tri 8470 9276 8493 9299 se
rect 8493 9276 8951 9299
rect 8470 7404 8951 9276
rect 9884 8286 9890 8338
rect 9942 8286 9954 8338
rect 10006 8286 10012 8338
tri 9340 7893 9362 7915 sw
rect 9340 7867 9362 7893
tri 9362 7867 9388 7893 sw
tri 8470 7355 8519 7404 ne
rect 8519 7355 8951 7404
rect 9884 7407 10012 8286
rect 9884 7355 9890 7407
rect 9942 7355 9954 7407
rect 10006 7355 10012 7407
rect 10569 7805 10575 7857
rect 10627 7805 10639 7857
rect 10691 7805 10697 7857
rect 10569 7800 10650 7805
tri 10650 7800 10655 7805 nw
tri 8519 7351 8523 7355 ne
rect 8523 7351 8951 7355
tri 8523 7348 8526 7351 ne
rect 8526 6314 8951 7351
tri 10544 7278 10569 7303 se
rect 10569 7278 10621 7800
tri 10621 7771 10650 7800 nw
rect 10493 7226 10499 7278
rect 10551 7226 10563 7278
rect 10615 7226 10621 7278
rect 10457 7019 10594 7040
rect 10457 6839 10466 7019
rect 10582 6839 10594 7019
rect 8830 6231 8882 6259
tri 8796 6201 8826 6231 ne
rect 8826 6201 8882 6231
rect 8286 6137 8564 6201
tri 8826 6197 8830 6201 ne
rect 8286 6100 8350 6137
tri 8350 6112 8375 6137 nw
tri 8475 6112 8500 6137 ne
rect 8286 6048 8292 6100
rect 8344 6048 8350 6100
rect 8286 6036 8350 6048
rect 8286 5984 8292 6036
rect 8344 5984 8350 6036
rect 7502 5296 8100 5616
rect 7502 5204 8008 5296
tri 8008 5204 8100 5296 nw
rect 6980 4113 7307 5122
rect 7502 4480 7982 5204
tri 7982 5178 8008 5204 nw
tri 7119 4091 7141 4113 ne
rect 7141 4091 7307 4113
tri 7141 4079 7153 4091 ne
rect 7153 3500 7307 4091
rect 7153 3320 7178 3500
rect 7294 3320 7307 3500
tri 7119 3110 7153 3144 se
rect 7153 3110 7307 3320
rect 6980 2958 7307 3110
rect 6980 2906 7020 2958
rect 7072 2906 7084 2958
rect 7136 2906 7307 2958
rect 6980 2302 7307 2906
rect 7335 3619 7341 3671
rect 7393 3619 7405 3671
rect 7457 3619 7463 3671
rect 7335 2519 7463 3619
tri 7463 2519 7475 2531 sw
rect 7335 2497 7475 2519
tri 7475 2497 7497 2519 sw
rect 7335 2416 7668 2497
tri 7506 2382 7540 2416 ne
rect 7540 2364 7546 2416
rect 7598 2364 7610 2416
rect 7662 2364 7668 2416
rect 8010 2302 8382 5122
tri 8427 2549 8500 2622 se
rect 8500 2553 8564 6137
rect 8830 5756 8882 6201
tri 9398 5327 9432 5361 se
tri 9040 5241 9074 5275 nw
rect 10457 4653 10594 6839
rect 10457 4473 10466 4653
rect 10582 4473 10594 4653
rect 10457 4458 10594 4473
rect 10805 4301 11907 10041
tri 12552 8369 12563 8380 se
rect 12563 8369 13107 10041
tri 12521 8338 12552 8369 se
rect 12552 8338 13107 8369
tri 12478 8295 12521 8338 se
rect 12521 8295 13107 8338
tri 12469 8286 12478 8295 se
rect 12478 8286 13107 8295
tri 12407 8224 12469 8286 se
rect 12469 8224 13107 8286
rect 12407 8207 13107 8224
rect 12407 8203 13103 8207
tri 13103 8203 13107 8207 nw
rect 12407 8196 13096 8203
tri 13096 8196 13103 8203 nw
rect 12407 8144 13044 8196
tri 13044 8144 13096 8196 nw
rect 12407 8132 13032 8144
tri 13032 8132 13044 8144 nw
rect 12015 7715 12067 7721
rect 12015 7651 12067 7663
rect 12015 5960 12067 7599
rect 12251 7275 12257 7327
rect 12309 7275 12321 7327
rect 12373 7275 12379 7327
rect 12015 5896 12067 5908
rect 12015 5838 12067 5844
rect 12171 6024 12223 6030
rect 12171 5960 12223 5972
tri 12146 4820 12171 4845 se
rect 12171 4820 12223 5908
rect 12015 4810 12067 4816
rect 12015 4746 12067 4758
tri 11975 4245 12015 4285 se
rect 12015 4255 12067 4694
rect 12015 4245 12057 4255
tri 12057 4245 12067 4255 nw
tri 11530 4199 11576 4245 se
rect 11576 4199 12011 4245
tri 12011 4199 12057 4245 nw
rect 11530 4193 12005 4199
tri 12005 4193 12011 4199 nw
rect 11530 4192 11610 4193
tri 11610 4192 11611 4193 nw
rect 12251 4192 12379 7275
rect 11530 4170 11588 4192
tri 11588 4170 11610 4192 nw
rect 8500 2549 8560 2553
tri 8560 2549 8564 2553 nw
rect 9642 4148 9886 4170
rect 9642 4092 9653 4148
rect 9709 4092 9735 4148
rect 9791 4092 9817 4148
rect 9873 4092 9886 4148
rect 9642 4065 9886 4092
rect 9642 4009 9653 4065
rect 9709 4009 9735 4065
rect 9791 4009 9817 4065
rect 9873 4009 9886 4065
rect 9642 3982 9886 4009
rect 9642 3926 9653 3982
rect 9709 3926 9735 3982
rect 9791 3926 9817 3982
rect 9873 3926 9886 3982
rect 9642 3899 9886 3926
rect 9642 3843 9653 3899
rect 9709 3843 9735 3899
rect 9791 3843 9817 3899
rect 9873 3843 9886 3899
rect 9642 3816 9886 3843
rect 9642 3760 9653 3816
rect 9709 3760 9735 3816
rect 9791 3760 9817 3816
rect 9873 3760 9886 3816
rect 9642 3733 9886 3760
rect 9642 3677 9653 3733
rect 9709 3677 9735 3733
rect 9791 3677 9817 3733
rect 9873 3677 9886 3733
rect 9642 3650 9886 3677
rect 9642 3594 9653 3650
rect 9709 3594 9735 3650
rect 9791 3594 9817 3650
rect 9873 3594 9886 3650
rect 9642 3567 9886 3594
rect 9642 3511 9653 3567
rect 9709 3511 9735 3567
rect 9791 3511 9817 3567
rect 9873 3511 9886 3567
rect 11241 3539 11247 3591
rect 11299 3539 11311 3591
rect 11363 3539 11369 3591
tri 11292 3514 11317 3539 ne
rect 9642 3483 9886 3511
rect 9642 3427 9653 3483
rect 9709 3427 9735 3483
rect 9791 3427 9817 3483
rect 9873 3427 9886 3483
rect 9642 3399 9886 3427
rect 9642 3343 9653 3399
rect 9709 3343 9735 3399
rect 9791 3343 9817 3399
rect 9873 3343 9886 3399
rect 8427 2531 8542 2549
tri 8542 2531 8560 2549 nw
rect 8427 2519 8530 2531
tri 8530 2519 8542 2531 nw
rect 8427 2497 8508 2519
tri 8508 2497 8530 2519 nw
rect 8427 2490 8501 2497
tri 8501 2490 8508 2497 nw
rect 8427 2302 8491 2490
tri 8491 2480 8501 2490 nw
rect 8547 2370 8651 2410
rect 9642 2302 9886 3343
rect 11317 2448 11369 3539
rect 11530 2451 11582 4170
tri 11582 4164 11588 4170 nw
tri 11530 2448 11533 2451 ne
rect 11533 2448 11582 2451
tri 11533 2428 11553 2448 ne
rect 11553 2365 11582 2448
rect 11610 4143 11930 4152
rect 11610 4087 11618 4143
rect 11674 4087 11698 4143
rect 11754 4087 11778 4143
rect 11834 4087 11858 4143
rect 11914 4087 11930 4143
rect 12251 4140 12257 4192
rect 12309 4140 12321 4192
rect 12373 4140 12379 4192
rect 12407 5464 13005 8132
tri 13005 8105 13032 8132 nw
tri 13341 7945 13375 7979 se
rect 13375 7945 13427 10041
rect 13458 9114 13510 10041
rect 13458 9050 13510 9062
rect 13458 8992 13510 8998
rect 14824 9831 15034 9849
rect 14824 9715 14841 9831
rect 15021 9715 15034 9831
rect 13299 7893 13305 7945
rect 13357 7893 13369 7945
rect 13421 7893 13427 7945
rect 13845 8196 14462 8203
rect 13845 8144 13851 8196
rect 13903 8144 13921 8196
rect 13973 8144 13990 8196
rect 14042 8144 14059 8196
rect 14111 8144 14128 8196
rect 14180 8144 14197 8196
rect 14249 8144 14266 8196
rect 14318 8144 14335 8196
rect 14387 8144 14404 8196
rect 14456 8144 14462 8196
rect 13845 8132 14462 8144
rect 13845 8080 13851 8132
rect 13903 8080 13921 8132
rect 13973 8080 13990 8132
rect 14042 8080 14059 8132
rect 14111 8080 14128 8132
rect 14180 8080 14197 8132
rect 14249 8080 14266 8132
rect 14318 8080 14335 8132
rect 14387 8080 14404 8132
rect 14456 8080 14462 8132
rect 13845 7558 14462 8080
rect 13845 7506 13851 7558
rect 13903 7506 13921 7558
rect 13973 7506 13990 7558
rect 14042 7506 14059 7558
rect 14111 7506 14128 7558
rect 14180 7506 14197 7558
rect 14249 7506 14266 7558
rect 14318 7506 14335 7558
rect 14387 7506 14404 7558
rect 14456 7506 14462 7558
rect 13845 7494 14462 7506
rect 13845 7442 13851 7494
rect 13903 7442 13921 7494
rect 13973 7442 13990 7494
rect 14042 7442 14059 7494
rect 14111 7442 14128 7494
rect 14180 7442 14197 7494
rect 14249 7442 14266 7494
rect 14318 7442 14335 7494
rect 14387 7442 14404 7494
rect 14456 7442 14462 7494
rect 13845 7435 14462 7442
rect 14824 6994 15034 9715
rect 16494 8726 16546 8732
rect 16494 8662 16546 8674
tri 16463 8338 16494 8369 se
rect 16494 8347 16546 8610
tri 16420 8295 16463 8338 se
rect 16463 8295 16494 8338
tri 16494 8295 16546 8347 nw
rect 16586 8612 16638 8618
rect 16586 8548 16638 8560
tri 16411 8286 16420 8295 se
tri 16346 8221 16411 8286 se
rect 16411 8221 16420 8286
tri 16420 8221 16494 8295 nw
tri 16523 8221 16586 8284 se
rect 16586 8262 16638 8496
tri 16729 8493 16754 8518 se
rect 16754 8493 16806 10664
rect 16678 8441 16684 8493
rect 16736 8441 16748 8493
rect 16800 8441 16806 8493
tri 16328 8203 16346 8221 se
tri 16272 8147 16328 8203 se
rect 16328 8147 16346 8203
tri 16346 8147 16420 8221 nw
tri 16512 8210 16523 8221 se
rect 16523 8210 16586 8221
tri 16586 8210 16638 8262 nw
tri 16449 8147 16512 8210 se
tri 16198 8073 16272 8147 se
tri 16272 8073 16346 8147 nw
tri 16438 8136 16449 8147 se
rect 16449 8136 16512 8147
tri 16512 8136 16586 8210 nw
tri 16375 8073 16438 8136 se
tri 16124 7999 16198 8073 se
tri 16198 7999 16272 8073 nw
tri 16364 8062 16375 8073 se
rect 16375 8062 16438 8073
tri 16438 8062 16512 8136 nw
tri 16301 7999 16364 8062 se
tri 16104 7979 16124 7999 se
tri 16070 7945 16104 7979 se
rect 16104 7945 16124 7979
tri 16050 7925 16070 7945 se
rect 16070 7925 16124 7945
tri 16124 7925 16198 7999 nw
tri 16290 7988 16301 7999 se
rect 16301 7988 16364 7999
tri 16364 7988 16438 8062 nw
tri 16227 7925 16290 7988 se
tri 16018 7893 16050 7925 se
tri 15992 7867 16018 7893 se
rect 16018 7867 16050 7893
tri 15982 7857 15992 7867 se
rect 15992 7857 16050 7867
tri 15976 7851 15982 7857 se
rect 15982 7851 16050 7857
tri 16050 7851 16124 7925 nw
tri 16216 7914 16227 7925 se
rect 16227 7914 16290 7925
tri 16290 7914 16364 7988 nw
tri 16153 7851 16216 7914 se
rect 14824 6878 14832 6994
rect 15012 6878 15034 6994
rect 14824 6032 15034 6878
tri 15949 7824 15976 7851 se
rect 15976 7824 16023 7851
tri 16023 7824 16050 7851 nw
tri 16142 7840 16153 7851 se
rect 16153 7840 16216 7851
tri 16216 7840 16290 7914 nw
tri 16126 7824 16142 7840 se
rect 15949 7805 16004 7824
tri 16004 7805 16023 7824 nw
tri 16107 7805 16126 7824 se
rect 16126 7805 16142 7824
rect 15949 6608 16001 7805
tri 16001 7802 16004 7805 nw
tri 16104 7802 16107 7805 se
rect 16107 7802 16142 7805
tri 16068 7766 16104 7802 se
rect 16104 7766 16142 7802
tri 16142 7766 16216 7840 nw
tri 16041 7739 16068 7766 se
rect 16068 7739 16115 7766
tri 16115 7739 16142 7766 nw
rect 16041 7721 16097 7739
tri 16097 7721 16115 7739 nw
tri 16035 6785 16041 6791 se
rect 16041 6785 16093 7721
tri 16093 7717 16097 7721 nw
rect 16407 7715 16459 7721
rect 16407 7651 16459 7663
rect 16035 6779 16093 6785
rect 16087 6727 16093 6779
rect 16035 6715 16093 6727
rect 16087 6663 16093 6715
rect 16035 6657 16093 6663
rect 16225 7403 16277 7409
rect 16225 7339 16277 7351
rect 15949 6544 16001 6556
rect 15949 6486 16001 6492
rect 16225 5906 16277 7287
rect 16407 7323 16459 7599
rect 16407 7259 16459 7271
rect 16407 7201 16459 7207
rect 16225 5842 16277 5854
rect 16225 5784 16277 5790
rect 16407 7155 16459 7161
rect 16407 7091 16459 7103
rect 12407 5204 12864 5464
tri 12864 5323 13005 5464 nw
rect 12407 5152 12678 5204
rect 12730 5152 12742 5204
rect 12794 5152 12806 5204
rect 12858 5152 12864 5204
rect 11610 4060 11930 4087
rect 11610 4004 11618 4060
rect 11674 4004 11698 4060
rect 11754 4004 11778 4060
rect 11834 4004 11858 4060
rect 11914 4004 11930 4060
rect 11610 3977 11930 4004
rect 11610 3921 11618 3977
rect 11674 3921 11698 3977
rect 11754 3921 11778 3977
rect 11834 3921 11858 3977
rect 11914 3921 11930 3977
rect 11610 3894 11930 3921
rect 11610 3838 11618 3894
rect 11674 3838 11698 3894
rect 11754 3838 11778 3894
rect 11834 3838 11858 3894
rect 11914 3838 11930 3894
rect 11610 3811 11930 3838
rect 11610 3755 11618 3811
rect 11674 3755 11698 3811
rect 11754 3755 11778 3811
rect 11834 3755 11858 3811
rect 11914 3755 11930 3811
rect 11610 3728 11930 3755
rect 11610 3672 11618 3728
rect 11674 3672 11698 3728
rect 11754 3672 11778 3728
rect 11834 3672 11858 3728
rect 11914 3672 11930 3728
rect 11610 3645 11930 3672
rect 11610 3589 11618 3645
rect 11674 3589 11698 3645
rect 11754 3589 11778 3645
rect 11834 3589 11858 3645
rect 11914 3589 11930 3645
rect 11610 3562 11930 3589
rect 11610 3506 11618 3562
rect 11674 3506 11698 3562
rect 11754 3506 11778 3562
rect 11834 3506 11858 3562
rect 11914 3506 11930 3562
rect 11610 3478 11930 3506
rect 11610 3422 11618 3478
rect 11674 3422 11698 3478
rect 11754 3422 11778 3478
rect 11834 3422 11858 3478
rect 11914 3422 11930 3478
rect 11610 3394 11930 3422
rect 11610 3338 11618 3394
rect 11674 3338 11698 3394
rect 11754 3338 11778 3394
rect 11834 3338 11858 3394
rect 11914 3338 11930 3394
tri 9932 2336 9957 2361 ne
rect 9957 2336 9960 2361
tri 9957 2333 9960 2336 ne
rect 10012 2336 10048 2361
tri 10048 2336 10073 2361 nw
rect 10012 2330 10042 2336
tri 10042 2330 10048 2336 nw
rect 10012 2320 10032 2330
tri 10032 2320 10042 2330 nw
rect 10012 2302 10014 2320
tri 10014 2302 10032 2320 nw
rect 11610 2302 11930 3338
rect 12185 3431 12237 3437
rect 12185 3367 12237 3379
rect 12185 3027 12237 3315
rect 12185 2963 12237 2975
rect 12185 2905 12237 2911
rect 12407 2416 12864 5152
rect 15714 5180 16351 5189
rect 15766 5128 15786 5180
rect 15838 5128 15858 5180
rect 15910 5128 15930 5180
rect 15982 5128 16002 5180
rect 16054 5128 16351 5180
rect 13679 4192 14074 5122
rect 15714 5101 16351 5128
rect 15766 5049 15786 5101
rect 15838 5049 15858 5101
rect 15910 5049 15930 5101
rect 15982 5049 16002 5101
rect 16054 5049 16351 5101
rect 15714 5021 16351 5049
rect 15766 4969 15786 5021
rect 15838 4969 15858 5021
rect 15910 4969 15930 5021
rect 15982 4969 16002 5021
rect 16054 4969 16351 5021
rect 15714 4945 16351 4969
tri 15714 4884 15775 4945 ne
rect 15775 4884 16351 4945
tri 15775 4870 15789 4884 ne
rect 15789 4870 16351 4884
tri 15789 4818 15841 4870 ne
rect 15841 4818 16351 4870
tri 15841 4816 15843 4818 ne
rect 15843 4816 16351 4818
tri 15843 4715 15944 4816 ne
rect 15944 4423 16351 4816
tri 13679 4140 13731 4192 ne
rect 13731 4140 14074 4192
tri 13731 4091 13780 4140 ne
rect 13780 4091 14074 4140
tri 13780 4042 13829 4091 ne
tri 13798 3505 13829 3536 se
rect 13829 3505 14074 4091
rect 15111 4076 15387 4230
tri 13795 3502 13798 3505 se
rect 13798 3502 14074 3505
rect 13829 3322 14074 3502
tri 13795 3319 13798 3322 ne
rect 13798 3319 14074 3322
tri 13798 3309 13808 3319 ne
rect 13808 3309 14074 3319
tri 13808 3288 13829 3309 ne
rect 12407 2364 12413 2416
rect 12465 2364 12477 2416
rect 12529 2364 12541 2416
rect 12593 2364 12605 2416
rect 12657 2364 12669 2416
rect 12721 2364 12733 2416
rect 12785 2364 12797 2416
rect 12849 2364 12864 2416
rect 12407 2302 12864 2364
tri 13766 2793 13829 2856 se
rect 13829 2793 14074 3309
rect 13766 2733 14074 2793
rect 13766 2712 14053 2733
tri 14053 2712 14074 2733 nw
tri 10012 2300 10014 2302 nw
rect 13766 2301 14011 2712
tri 14011 2670 14053 2712 nw
tri 14787 2326 14791 2330 sw
rect 14787 2320 14791 2326
tri 14791 2320 14797 2326 sw
rect 14787 2302 14797 2320
tri 14797 2302 14815 2320 sw
tri 14471 1980 14475 1984 ne
rect 14475 1980 14495 1984
tri 14475 1968 14487 1980 ne
rect 14487 1968 14495 1980
tri 14487 1960 14495 1968 ne
rect 16031 1881 16351 4423
rect 16407 2320 16459 7039
rect 23171 6966 23223 6972
rect 23171 6902 23223 6914
rect 23171 6844 23223 6850
rect 17234 3602 17240 3654
rect 17292 3602 17304 3654
rect 17356 3602 17362 3654
rect 19766 3499 20585 3507
rect 19766 3447 19772 3499
rect 19824 3447 19841 3499
rect 19893 3447 19910 3499
rect 19962 3447 19979 3499
rect 20031 3447 20048 3499
rect 20100 3447 20117 3499
rect 20169 3447 20186 3499
rect 20238 3447 20255 3499
rect 20307 3447 20323 3499
rect 20375 3447 20391 3499
rect 20443 3447 20459 3499
rect 20511 3447 20527 3499
rect 20579 3447 20585 3499
rect 19766 3435 20585 3447
rect 19766 3383 19772 3435
rect 19824 3383 19841 3435
rect 19893 3383 19910 3435
rect 19962 3383 19979 3435
rect 20031 3383 20048 3435
rect 20100 3383 20117 3435
rect 20169 3383 20186 3435
rect 20238 3383 20255 3435
rect 20307 3383 20323 3435
rect 20375 3383 20391 3435
rect 20443 3383 20459 3435
rect 20511 3383 20527 3435
rect 20579 3383 20585 3435
rect 21156 3505 21348 3507
rect 21156 3389 21162 3505
rect 21342 3389 21348 3505
rect 21156 3387 21348 3389
rect 19766 3371 20585 3383
rect 19766 3319 19772 3371
rect 19824 3319 19841 3371
rect 19893 3319 19910 3371
rect 19962 3319 19979 3371
rect 20031 3319 20048 3371
rect 20100 3319 20117 3371
rect 20169 3319 20186 3371
rect 20238 3319 20255 3371
rect 20307 3319 20323 3371
rect 20375 3319 20391 3371
rect 20443 3319 20459 3371
rect 20511 3319 20527 3371
rect 20579 3319 20585 3371
rect 19766 3311 20585 3319
rect 20669 2660 20675 2712
rect 20727 2660 20739 2712
rect 20791 2660 20803 2712
rect 20855 2660 20867 2712
rect 20919 2660 20925 2712
rect 16407 2256 16459 2268
rect 16407 2198 16459 2204
rect 20651 2032 20933 2035
rect 20651 1980 20657 2032
rect 20709 1980 20730 2032
rect 20782 1980 20803 2032
rect 20855 1980 20875 2032
rect 20927 1980 20933 2032
rect 20651 1968 20933 1980
rect 20651 1916 20657 1968
rect 20709 1916 20730 1968
rect 20782 1916 20803 1968
rect 20855 1916 20875 1968
rect 20927 1916 20933 1968
rect 20651 1904 20933 1916
rect 20651 1852 20657 1904
rect 20709 1852 20730 1904
rect 20782 1852 20803 1904
rect 20855 1852 20875 1904
rect 20927 1852 20933 1904
rect 20651 1849 20933 1852
<< via2 >>
rect 1911 11348 1967 11404
rect 1911 11268 1967 11324
rect 1911 11188 1967 11244
rect 861 10506 917 10562
rect 941 10506 997 10562
rect 861 10425 917 10481
rect 941 10425 997 10481
rect 861 10344 917 10400
rect 941 10344 997 10400
rect 861 10263 917 10319
rect 941 10263 997 10319
rect 861 10182 917 10238
rect 941 10182 997 10238
rect 861 10101 917 10157
rect 941 10101 997 10157
rect 861 10020 917 10076
rect 941 10020 997 10076
rect 861 9939 917 9995
rect 941 9939 997 9995
rect 861 9858 917 9914
rect 941 9858 997 9914
rect 861 9776 917 9832
rect 941 9776 997 9832
rect 861 9694 917 9750
rect 941 9694 997 9750
rect 1911 11107 1967 11163
rect 861 9612 917 9668
rect 941 9612 997 9668
rect 861 9530 917 9586
rect 941 9530 997 9586
rect 861 9448 917 9504
rect 941 9448 997 9504
rect 861 9366 917 9422
rect 941 9366 997 9422
rect 861 9284 917 9340
rect 941 9284 997 9340
rect 861 9202 917 9258
rect 941 9202 997 9258
rect 861 9120 917 9176
rect 941 9120 997 9176
rect 861 9038 917 9094
rect 941 9038 997 9094
rect 861 8956 917 9012
rect 941 8956 997 9012
rect 861 8874 917 8930
rect 941 8874 997 8930
rect 861 8792 917 8848
rect 941 8792 997 8848
rect 861 8710 917 8766
rect 941 8710 997 8766
rect 861 8628 917 8684
rect 941 8628 997 8684
rect 861 8546 917 8602
rect 941 8546 997 8602
rect 861 8464 917 8520
rect 941 8464 997 8520
rect 861 8382 917 8438
rect 941 8382 997 8438
rect 861 8300 917 8356
rect 941 8300 997 8356
rect 861 8218 917 8274
rect 941 8218 997 8274
rect 861 8136 917 8192
rect 941 8136 997 8192
rect 861 8054 917 8110
rect 941 8054 997 8110
rect 861 7972 917 8028
rect 941 7972 997 8028
rect 861 7890 917 7946
rect 941 7890 997 7946
rect 861 7808 917 7864
rect 941 7808 997 7864
rect 1480 5203 1536 5259
rect 1480 5117 1536 5173
rect 1480 5031 1536 5087
rect 1480 4945 1536 5001
rect 1480 4859 1536 4915
rect 1480 4772 1536 4828
rect 1480 4685 1536 4741
rect 9653 4092 9709 4148
rect 9735 4092 9791 4148
rect 9817 4092 9873 4148
rect 9653 4009 9709 4065
rect 9735 4009 9791 4065
rect 9817 4009 9873 4065
rect 9653 3926 9709 3982
rect 9735 3926 9791 3982
rect 9817 3926 9873 3982
rect 9653 3843 9709 3899
rect 9735 3843 9791 3899
rect 9817 3843 9873 3899
rect 9653 3760 9709 3816
rect 9735 3760 9791 3816
rect 9817 3760 9873 3816
rect 9653 3677 9709 3733
rect 9735 3677 9791 3733
rect 9817 3677 9873 3733
rect 9653 3594 9709 3650
rect 9735 3594 9791 3650
rect 9817 3594 9873 3650
rect 9653 3511 9709 3567
rect 9735 3511 9791 3567
rect 9817 3511 9873 3567
rect 9653 3427 9709 3483
rect 9735 3427 9791 3483
rect 9817 3427 9873 3483
rect 9653 3343 9709 3399
rect 9735 3343 9791 3399
rect 9817 3343 9873 3399
rect 11618 4087 11674 4143
rect 11698 4087 11754 4143
rect 11778 4087 11834 4143
rect 11858 4087 11914 4143
rect 11618 4004 11674 4060
rect 11698 4004 11754 4060
rect 11778 4004 11834 4060
rect 11858 4004 11914 4060
rect 11618 3921 11674 3977
rect 11698 3921 11754 3977
rect 11778 3921 11834 3977
rect 11858 3921 11914 3977
rect 11618 3838 11674 3894
rect 11698 3838 11754 3894
rect 11778 3838 11834 3894
rect 11858 3838 11914 3894
rect 11618 3755 11674 3811
rect 11698 3755 11754 3811
rect 11778 3755 11834 3811
rect 11858 3755 11914 3811
rect 11618 3672 11674 3728
rect 11698 3672 11754 3728
rect 11778 3672 11834 3728
rect 11858 3672 11914 3728
rect 11618 3589 11674 3645
rect 11698 3589 11754 3645
rect 11778 3589 11834 3645
rect 11858 3589 11914 3645
rect 11618 3506 11674 3562
rect 11698 3506 11754 3562
rect 11778 3506 11834 3562
rect 11858 3506 11914 3562
rect 11618 3422 11674 3478
rect 11698 3422 11754 3478
rect 11778 3422 11834 3478
rect 11858 3422 11914 3478
rect 11618 3338 11674 3394
rect 11698 3338 11754 3394
rect 11778 3338 11834 3394
rect 11858 3338 11914 3394
<< metal3 >>
rect 1882 11404 1996 11409
rect 1882 11348 1911 11404
rect 1967 11348 1996 11404
rect 1882 11324 1996 11348
rect 1882 11268 1911 11324
rect 1967 11268 1996 11324
rect 1882 11244 1996 11268
rect 1882 11188 1911 11244
rect 1967 11188 1996 11244
rect 1882 11163 1996 11188
rect 1882 11107 1911 11163
rect 1967 11107 1996 11163
rect 1882 11102 1996 11107
rect 181 10562 8894 10594
rect 181 10506 861 10562
rect 917 10506 941 10562
rect 997 10506 8894 10562
rect 181 10481 8894 10506
rect 181 10425 861 10481
rect 917 10425 941 10481
rect 997 10425 8894 10481
rect 181 10400 8894 10425
rect 181 10344 861 10400
rect 917 10344 941 10400
rect 997 10344 8894 10400
rect 181 10319 8894 10344
rect 181 10263 861 10319
rect 917 10263 941 10319
rect 997 10263 8894 10319
rect 181 10238 8894 10263
rect 181 10182 861 10238
rect 917 10182 941 10238
rect 997 10182 8894 10238
rect 181 10157 8894 10182
rect 181 10101 861 10157
rect 917 10101 941 10157
rect 997 10101 8894 10157
rect 181 10076 8894 10101
rect 181 10020 861 10076
rect 917 10020 941 10076
rect 997 10020 8894 10076
rect 181 9995 8894 10020
rect 181 9939 861 9995
rect 917 9939 941 9995
rect 997 9939 8894 9995
rect 181 9914 8894 9939
rect 181 9858 861 9914
rect 917 9858 941 9914
rect 997 9858 8894 9914
rect 181 9832 8894 9858
rect 181 9776 861 9832
rect 917 9776 941 9832
rect 997 9776 8894 9832
rect 181 9750 8894 9776
rect 181 9694 861 9750
rect 917 9694 941 9750
rect 997 9694 8894 9750
rect 181 9668 8894 9694
rect 181 9612 861 9668
rect 917 9612 941 9668
rect 997 9612 8894 9668
rect 181 9586 8894 9612
rect 181 9530 861 9586
rect 917 9530 941 9586
rect 997 9530 8894 9586
rect 181 9504 8894 9530
rect 181 9448 861 9504
rect 917 9448 941 9504
rect 997 9448 8894 9504
rect 181 9422 8894 9448
rect 181 9366 861 9422
rect 917 9366 941 9422
rect 997 9366 8894 9422
rect 181 9340 8894 9366
rect 181 9284 861 9340
rect 917 9284 941 9340
rect 997 9284 8894 9340
rect 181 9258 8894 9284
rect 181 9202 861 9258
rect 917 9202 941 9258
rect 997 9202 8894 9258
rect 181 9176 8894 9202
rect 181 9120 861 9176
rect 917 9120 941 9176
rect 997 9120 8894 9176
rect 181 9094 8894 9120
rect 181 9038 861 9094
rect 917 9038 941 9094
rect 997 9038 8894 9094
rect 181 9012 8894 9038
rect 181 8956 861 9012
rect 917 8956 941 9012
rect 997 8956 8894 9012
rect 181 8930 8894 8956
rect 181 8874 861 8930
rect 917 8874 941 8930
rect 997 8874 8894 8930
rect 181 8848 8894 8874
rect 181 8792 861 8848
rect 917 8792 941 8848
rect 997 8792 8894 8848
rect 181 8766 8894 8792
rect 181 8710 861 8766
rect 917 8710 941 8766
rect 997 8710 8894 8766
rect 181 8684 8894 8710
rect 181 8628 861 8684
rect 917 8628 941 8684
rect 997 8628 8894 8684
rect 181 8602 8894 8628
rect 181 8546 861 8602
rect 917 8546 941 8602
rect 997 8546 8894 8602
rect 181 8520 8894 8546
rect 181 8464 861 8520
rect 917 8464 941 8520
rect 997 8464 8894 8520
rect 181 8438 8894 8464
rect 181 8382 861 8438
rect 917 8382 941 8438
rect 997 8382 8894 8438
rect 181 8356 8894 8382
rect 181 8300 861 8356
rect 917 8300 941 8356
rect 997 8300 8894 8356
rect 181 8274 8894 8300
rect 181 8218 861 8274
rect 917 8218 941 8274
rect 997 8218 8894 8274
rect 181 8192 8894 8218
rect 181 8136 861 8192
rect 917 8136 941 8192
rect 997 8136 8894 8192
rect 181 8110 8894 8136
rect 181 8054 861 8110
rect 917 8054 941 8110
rect 997 8054 8894 8110
rect 181 8028 8894 8054
rect 181 7972 861 8028
rect 917 7972 941 8028
rect 997 7972 8894 8028
rect 181 7946 8894 7972
rect 181 7890 861 7946
rect 917 7890 941 7946
rect 997 7890 8894 7946
rect 181 7864 8894 7890
rect 181 7808 861 7864
rect 917 7808 941 7864
rect 997 7808 8894 7864
rect 181 7760 8894 7808
rect 189 6034 8951 6892
rect 566 5259 12886 5535
rect 566 5203 1480 5259
rect 1536 5203 12886 5259
rect 566 5173 12886 5203
rect 566 5117 1480 5173
rect 1536 5117 12886 5173
rect 566 5087 12886 5117
rect 566 5031 1480 5087
rect 1536 5031 12886 5087
rect 566 5001 12886 5031
rect 566 4945 1480 5001
rect 1536 4945 12886 5001
rect 566 4915 12886 4945
rect 566 4859 1480 4915
rect 1536 4859 12886 4915
rect 566 4828 12886 4859
rect 566 4772 1480 4828
rect 1536 4772 12886 4828
rect 566 4741 12886 4772
rect 566 4685 1480 4741
rect 1536 4685 12886 4741
rect 566 4632 12886 4685
rect 974 4148 11977 4176
rect 974 4092 9653 4148
rect 9709 4092 9735 4148
rect 9791 4092 9817 4148
rect 9873 4143 11977 4148
rect 9873 4092 11618 4143
rect 974 4087 11618 4092
rect 11674 4087 11698 4143
rect 11754 4087 11778 4143
rect 11834 4087 11858 4143
rect 11914 4087 11977 4143
rect 974 4065 11977 4087
rect 974 4009 9653 4065
rect 9709 4009 9735 4065
rect 9791 4009 9817 4065
rect 9873 4060 11977 4065
rect 9873 4009 11618 4060
rect 974 4004 11618 4009
rect 11674 4004 11698 4060
rect 11754 4004 11778 4060
rect 11834 4004 11858 4060
rect 11914 4004 11977 4060
rect 974 3982 11977 4004
rect 974 3926 9653 3982
rect 9709 3926 9735 3982
rect 9791 3926 9817 3982
rect 9873 3977 11977 3982
rect 9873 3926 11618 3977
rect 974 3921 11618 3926
rect 11674 3921 11698 3977
rect 11754 3921 11778 3977
rect 11834 3921 11858 3977
rect 11914 3921 11977 3977
rect 974 3899 11977 3921
rect 974 3843 9653 3899
rect 9709 3843 9735 3899
rect 9791 3843 9817 3899
rect 9873 3894 11977 3899
rect 9873 3843 11618 3894
rect 974 3838 11618 3843
rect 11674 3838 11698 3894
rect 11754 3838 11778 3894
rect 11834 3838 11858 3894
rect 11914 3838 11977 3894
rect 974 3816 11977 3838
rect 974 3760 9653 3816
rect 9709 3760 9735 3816
rect 9791 3760 9817 3816
rect 9873 3811 11977 3816
rect 9873 3760 11618 3811
rect 974 3755 11618 3760
rect 11674 3755 11698 3811
rect 11754 3755 11778 3811
rect 11834 3755 11858 3811
rect 11914 3755 11977 3811
rect 974 3733 11977 3755
rect 974 3677 9653 3733
rect 9709 3677 9735 3733
rect 9791 3677 9817 3733
rect 9873 3728 11977 3733
rect 9873 3677 11618 3728
rect 974 3672 11618 3677
rect 11674 3672 11698 3728
rect 11754 3672 11778 3728
rect 11834 3672 11858 3728
rect 11914 3672 11977 3728
rect 974 3650 11977 3672
rect 974 3594 9653 3650
rect 9709 3594 9735 3650
rect 9791 3594 9817 3650
rect 9873 3645 11977 3650
rect 9873 3594 11618 3645
rect 974 3589 11618 3594
rect 11674 3589 11698 3645
rect 11754 3589 11778 3645
rect 11834 3589 11858 3645
rect 11914 3589 11977 3645
rect 974 3567 11977 3589
rect 974 3511 9653 3567
rect 9709 3511 9735 3567
rect 9791 3511 9817 3567
rect 9873 3562 11977 3567
rect 9873 3511 11618 3562
rect 974 3506 11618 3511
rect 11674 3506 11698 3562
rect 11754 3506 11778 3562
rect 11834 3506 11858 3562
rect 11914 3506 11977 3562
rect 974 3483 11977 3506
rect 974 3427 9653 3483
rect 9709 3427 9735 3483
rect 9791 3427 9817 3483
rect 9873 3478 11977 3483
rect 9873 3427 11618 3478
rect 974 3422 11618 3427
rect 11674 3422 11698 3478
rect 11754 3422 11778 3478
rect 11834 3422 11858 3478
rect 11914 3422 11977 3478
rect 974 3399 11977 3422
rect 974 3343 9653 3399
rect 9709 3343 9735 3399
rect 9791 3343 9817 3399
rect 9873 3394 11977 3399
rect 9873 3343 11618 3394
rect 974 3338 11618 3343
rect 11674 3338 11698 3394
rect 11754 3338 11778 3394
rect 11834 3338 11858 3394
rect 11914 3338 11977 3394
rect 974 3318 11977 3338
<< comment >>
rect 7416 2349 7678 2416
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_0
timestamp 1701704242
transform 1 0 11424 0 -1 5950
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_1
timestamp 1701704242
transform 1 0 11633 0 1 3545
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_2
timestamp 1701704242
transform 1 0 14553 0 1 5902
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1701704242
transform 0 -1 4144 1 0 9715
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1701704242
transform 0 -1 4456 1 0 9715
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1701704242
transform 0 -1 4946 1 0 9715
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_3
timestamp 1701704242
transform 0 -1 5298 1 0 9715
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_4
timestamp 1701704242
transform 0 -1 6444 1 0 9715
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_5
timestamp 1701704242
transform 0 -1 6796 1 0 9715
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_6
timestamp 1701704242
transform 0 -1 7168 1 0 9715
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_7
timestamp 1701704242
transform 0 -1 7520 1 0 9715
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_8
timestamp 1701704242
transform 1 0 7552 0 1 2368
box 0 0 1 1
use L1M1_CDNS_52468879185336  L1M1_CDNS_52468879185336_0
timestamp 1701704242
transform 0 -1 15333 1 0 8293
box -12 -6 1558 40
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_0
timestamp 1701704242
transform 0 -1 16546 -1 0 8732
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_1
timestamp 1701704242
transform 0 -1 729 -1 0 7280
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_2
timestamp 1701704242
transform 0 -1 2288 -1 0 4272
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_3
timestamp 1701704242
transform 0 -1 2055 -1 0 3281
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_4
timestamp 1701704242
transform 0 -1 2840 -1 0 5882
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_5
timestamp 1701704242
transform 0 -1 16638 -1 0 8618
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_6
timestamp 1701704242
transform 0 -1 16806 -1 0 10786
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_7
timestamp 1701704242
transform 0 1 5583 -1 0 10310
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_8
timestamp 1701704242
transform 0 1 16407 -1 0 2326
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_9
timestamp 1701704242
transform -1 0 10012 0 1 7355
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_10
timestamp 1701704242
transform -1 0 10012 0 1 8286
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_11
timestamp 1701704242
transform -1 0 2368 0 1 5984
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_12
timestamp 1701704242
transform -1 0 5936 0 1 6702
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_13
timestamp 1701704242
transform -1 0 3670 0 1 4818
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_14
timestamp 1701704242
transform -1 0 8369 0 1 9411
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_15
timestamp 1701704242
transform -1 0 10621 0 1 7226
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_16
timestamp 1701704242
transform -1 0 13427 0 1 7893
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_17
timestamp 1701704242
transform -1 0 4928 0 1 7597
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_18
timestamp 1701704242
transform -1 0 17362 0 1 3602
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_19
timestamp 1701704242
transform -1 0 11369 0 -1 3591
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_20
timestamp 1701704242
transform -1 0 6201 0 -1 10230
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_21
timestamp 1701704242
transform -1 0 1948 0 -1 6736
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_22
timestamp 1701704242
transform 0 1 13458 1 0 8992
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_23
timestamp 1701704242
transform 0 1 2913 1 0 7597
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_24
timestamp 1701704242
transform 0 1 15949 1 0 6486
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_25
timestamp 1701704242
transform 0 1 16035 1 0 6657
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_26
timestamp 1701704242
transform 0 -1 12067 1 0 7593
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_27
timestamp 1701704242
transform 0 -1 12067 1 0 5838
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_28
timestamp 1701704242
transform 0 -1 978 1 0 5678
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_29
timestamp 1701704242
transform 0 -1 106 1 0 3644
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_30
timestamp 1701704242
transform 0 -1 1416 1 0 2974
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_31
timestamp 1701704242
transform 0 -1 106 1 0 2974
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_32
timestamp 1701704242
transform 0 -1 1336 1 0 6064
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_33
timestamp 1701704242
transform 0 -1 16459 1 0 7201
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_34
timestamp 1701704242
transform 0 -1 16277 1 0 5784
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_35
timestamp 1701704242
transform 0 -1 12223 1 0 5902
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_36
timestamp 1701704242
transform 0 -1 16459 1 0 7033
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_37
timestamp 1701704242
transform 0 -1 16459 1 0 7593
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_38
timestamp 1701704242
transform 0 -1 16277 1 0 7281
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_39
timestamp 1701704242
transform 0 -1 12237 1 0 2905
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_40
timestamp 1701704242
transform 0 -1 12237 1 0 3309
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_41
timestamp 1701704242
transform 0 -1 12067 1 0 4688
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_42
timestamp 1701704242
transform 1 0 5572 0 -1 2490
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_43
timestamp 1701704242
transform 1 0 10569 0 -1 7857
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_44
timestamp 1701704242
transform 1 0 16678 0 -1 8493
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_45
timestamp 1701704242
transform 1 0 12251 0 1 4140
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_46
timestamp 1701704242
transform 1 0 6169 0 1 7228
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_47
timestamp 1701704242
transform 1 0 3622 0 1 2438
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_48
timestamp 1701704242
transform 1 0 7335 0 1 3619
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_49
timestamp 1701704242
transform 1 0 7540 0 1 2364
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_50
timestamp 1701704242
transform 1 0 4242 0 1 3809
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_51
timestamp 1701704242
transform 1 0 9300 0 1 9411
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_52
timestamp 1701704242
transform 1 0 6955 0 1 9299
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_53
timestamp 1701704242
transform 1 0 6955 0 1 10418
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_54
timestamp 1701704242
transform 1 0 9983 0 1 9375
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_55
timestamp 1701704242
transform 1 0 12251 0 1 7275
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_56
timestamp 1701704242
transform 1 0 7014 0 1 2906
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_0
timestamp 1701704242
transform 0 -1 7294 -1 0 3506
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_1
timestamp 1701704242
transform 0 1 410 -1 0 3507
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_2
timestamp 1701704242
transform 0 1 1881 -1 0 9187
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_3
timestamp 1701704242
transform 1 0 126 0 -1 2635
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_4
timestamp 1701704242
transform 1 0 14835 0 1 9715
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_5
timestamp 1701704242
transform 1 0 14826 0 1 6878
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_0
timestamp 1701704242
transform 0 1 410 -1 0 4091
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_1
timestamp 1701704242
transform 0 1 1881 -1 0 9833
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_2
timestamp 1701704242
transform 1 0 2396 0 -1 2635
box 0 0 1 1
use M1M2_CDNS_52468879185200  M1M2_CDNS_52468879185200_0
timestamp 1701704242
transform 1 0 117 0 -1 4660
box 0 0 1 1
use M1M2_CDNS_52468879185200  M1M2_CDNS_52468879185200_1
timestamp 1701704242
transform 1 0 10460 0 1 6839
box 0 0 1 1
use M1M2_CDNS_52468879185200  M1M2_CDNS_52468879185200_2
timestamp 1701704242
transform 1 0 10460 0 1 4473
box 0 0 1 1
use M1M2_CDNS_52468879185201  M1M2_CDNS_52468879185201_0
timestamp 1701704242
transform 0 1 12422 -1 0 3234
box 0 0 320 116
use M1M2_CDNS_52468879185201  M1M2_CDNS_52468879185201_1
timestamp 1701704242
transform 1 0 5010 0 -1 7559
box 0 0 320 116
use M1M2_CDNS_52468879185201  M1M2_CDNS_52468879185201_2
timestamp 1701704242
transform 1 0 5010 0 -1 8172
box 0 0 320 116
use M1M2_CDNS_52468879185201  M1M2_CDNS_52468879185201_3
timestamp 1701704242
transform 1 0 6357 0 -1 7559
box 0 0 320 116
use M1M2_CDNS_52468879185201  M1M2_CDNS_52468879185201_4
timestamp 1701704242
transform 1 0 6357 0 -1 8172
box 0 0 320 116
use M1M2_CDNS_52468879185201  M1M2_CDNS_52468879185201_5
timestamp 1701704242
transform 1 0 3705 0 -1 7559
box 0 0 320 116
use M1M2_CDNS_52468879185201  M1M2_CDNS_52468879185201_6
timestamp 1701704242
transform 1 0 3705 0 -1 8172
box 0 0 320 116
use M1M2_CDNS_52468879185201  M1M2_CDNS_52468879185201_7
timestamp 1701704242
transform 1 0 2241 0 -1 9834
box 0 0 320 116
use M1M2_CDNS_52468879185201  M1M2_CDNS_52468879185201_8
timestamp 1701704242
transform 1 0 1421 0 -1 9834
box 0 0 320 116
use M1M2_CDNS_52468879185201  M1M2_CDNS_52468879185201_9
timestamp 1701704242
transform 1 0 2993 0 -1 9834
box 0 0 320 116
use M1M2_CDNS_52468879185202  M1M2_CDNS_52468879185202_0
timestamp 1701704242
transform 1 0 2241 0 -1 10150
box 0 0 1 1
use M1M2_CDNS_52468879185202  M1M2_CDNS_52468879185202_1
timestamp 1701704242
transform 1 0 1421 0 -1 10150
box 0 0 1 1
use M1M2_CDNS_52468879185202  M1M2_CDNS_52468879185202_2
timestamp 1701704242
transform 1 0 2993 0 -1 10150
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_0
timestamp 1701704242
transform 1 0 12672 0 1 5152
box 0 0 1 1
use M1M2_CDNS_52468879185209  M1M2_CDNS_52468879185209_0
timestamp 1701704242
transform 0 -1 4498 -1 0 4428
box 0 0 128 244
use M1M2_CDNS_52468879185209  M1M2_CDNS_52468879185209_1
timestamp 1701704242
transform 1 0 10460 0 1 5380
box 0 0 128 244
use M1M2_CDNS_52468879185297  M1M2_CDNS_52468879185297_0
timestamp 1701704242
transform -1 0 4498 0 1 3539
box 0 0 1 1
use M1M2_CDNS_52468879185297  M1M2_CDNS_52468879185297_1
timestamp 1701704242
transform 0 -1 23 1 0 9872
box 0 0 1 1
use M1M2_CDNS_52468879185297  M1M2_CDNS_52468879185297_2
timestamp 1701704242
transform 1 0 20669 0 1 2660
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_0
timestamp 1701704242
transform -1 0 8350 0 -1 6100
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_1
timestamp 1701704242
transform 1 0 1884 0 -1 4884
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_2
timestamp 1701704242
transform 1 0 6233 0 1 7684
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_3
timestamp 1701704242
transform 1 0 6999 0 1 7684
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_4
timestamp 1701704242
transform 1 0 6999 0 1 8301
box 0 0 1 1
use M1M2_CDNS_52468879185371  M1M2_CDNS_52468879185371_0
timestamp 1701704242
transform 1 0 5969 0 1 6323
box 0 0 1 1
use M1M2_CDNS_52468879185371  M1M2_CDNS_52468879185371_1
timestamp 1701704242
transform 1 0 5675 0 1 6323
box 0 0 1 1
use M1M2_CDNS_52468879185967  M1M2_CDNS_52468879185967_0
timestamp 1701704242
transform 1 0 1525 0 -1 2635
box 0 0 448 116
use M1M2_CDNS_52468879185967  M1M2_CDNS_52468879185967_1
timestamp 1701704242
transform 1 0 8489 0 -1 7557
box 0 0 448 116
use M1M2_CDNS_52468879185967  M1M2_CDNS_52468879185967_2
timestamp 1701704242
transform 1 0 8489 0 -1 8175
box 0 0 448 116
use M1M2_CDNS_52468879185967  M1M2_CDNS_52468879185967_3
timestamp 1701704242
transform 1 0 7639 0 -1 9832
box 0 0 448 116
use M1M2_CDNS_52468879185970  M1M2_CDNS_52468879185970_0
timestamp 1701704242
transform 0 -1 2965 -1 0 10786
box 0 0 1 1
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_0
timestamp 1701704242
transform 1 0 13877 0 1 3322
box 0 0 192 180
use M1M2_CDNS_524688791851032  M1M2_CDNS_524688791851032_0
timestamp 1701704242
transform 0 1 8010 -1 0 5120
box 0 0 192 372
use M1M2_CDNS_524688791851032  M1M2_CDNS_524688791851032_1
timestamp 1701704242
transform 0 1 8010 -1 0 3506
box 0 0 192 372
use M1M2_CDNS_524688791851077  M1M2_CDNS_524688791851077_0
timestamp 1701704242
transform -1 0 3192 0 -1 2852
box 0 0 320 180
use M1M2_CDNS_524688791851077  M1M2_CDNS_524688791851077_1
timestamp 1701704242
transform 1 0 5010 0 -1 8652
box 0 0 320 180
use M1M2_CDNS_524688791851077  M1M2_CDNS_524688791851077_2
timestamp 1701704242
transform 1 0 6357 0 -1 8652
box 0 0 320 180
use M1M2_CDNS_524688791851077  M1M2_CDNS_524688791851077_3
timestamp 1701704242
transform 1 0 3705 0 -1 8652
box 0 0 320 180
use M1M2_CDNS_524688791851077  M1M2_CDNS_524688791851077_4
timestamp 1701704242
transform 1 0 2396 0 -1 4660
box 0 0 320 180
use M1M2_CDNS_524688791851077  M1M2_CDNS_524688791851077_5
timestamp 1701704242
transform 1 0 2241 0 -1 7032
box 0 0 320 180
use M1M2_CDNS_524688791851077  M1M2_CDNS_524688791851077_6
timestamp 1701704242
transform 1 0 2241 0 -1 9191
box 0 0 320 180
use M1M2_CDNS_524688791851077  M1M2_CDNS_524688791851077_7
timestamp 1701704242
transform 1 0 3026 0 -1 4660
box 0 0 320 180
use M1M2_CDNS_524688791851077  M1M2_CDNS_524688791851077_8
timestamp 1701704242
transform 1 0 2993 0 -1 7040
box 0 0 320 180
use M1M2_CDNS_524688791851077  M1M2_CDNS_524688791851077_9
timestamp 1701704242
transform 1 0 2993 0 -1 9191
box 0 0 320 180
use M1M2_CDNS_524688791851077  M1M2_CDNS_524688791851077_10
timestamp 1701704242
transform 1 0 5010 0 1 6323
box 0 0 320 180
use M1M2_CDNS_524688791851077  M1M2_CDNS_524688791851077_11
timestamp 1701704242
transform 1 0 6357 0 1 6323
box 0 0 320 180
use M1M2_CDNS_524688791851077  M1M2_CDNS_524688791851077_12
timestamp 1701704242
transform 1 0 3705 0 1 6323
box 0 0 320 180
use M1M2_CDNS_524688791851084  M1M2_CDNS_524688791851084_0
timestamp 1701704242
transform 1 0 4073 0 1 5152
box 0 0 512 52
use M1M2_CDNS_524688791851113  M1M2_CDNS_524688791851113_0
timestamp 1701704242
transform -1 0 529 0 -1 10150
box 0 0 1 1
use M1M2_CDNS_524688791851113  M1M2_CDNS_524688791851113_1
timestamp 1701704242
transform 1 0 7639 0 -1 10150
box 0 0 1 1
use M1M2_CDNS_524688791851113  M1M2_CDNS_524688791851113_2
timestamp 1701704242
transform 1 0 12407 0 1 2364
box 0 0 1 1
use M1M2_CDNS_524688791851144  M1M2_CDNS_524688791851144_0
timestamp 1701704242
transform 1 0 117 0 -1 7040
box 0 0 384 180
use M1M2_CDNS_524688791851144  M1M2_CDNS_524688791851144_1
timestamp 1701704242
transform 1 0 13685 0 -1 5111
box 0 0 384 180
use M1M2_CDNS_524688791851144  M1M2_CDNS_524688791851144_2
timestamp 1701704242
transform 1 0 117 0 -1 9191
box 0 0 384 180
use M1M2_CDNS_524688791851144  M1M2_CDNS_524688791851144_3
timestamp 1701704242
transform 1 0 1473 0 -1 7040
box 0 0 384 180
use M1M2_CDNS_524688791851144  M1M2_CDNS_524688791851144_4
timestamp 1701704242
transform 1 0 8546 0 1 6323
box 0 0 384 180
use M1M2_CDNS_524688791851151  M1M2_CDNS_524688791851151_0
timestamp 1701704242
transform 1 0 841 0 -1 8652
box 0 0 512 180
use M1M2_CDNS_524688791851151  M1M2_CDNS_524688791851151_1
timestamp 1701704242
transform 1 0 841 0 1 6323
box 0 0 512 180
use M1M2_CDNS_524688791851177  M1M2_CDNS_524688791851177_0
timestamp 1701704242
transform 1 0 117 0 -1 9849
box 0 0 384 116
use M1M2_CDNS_524688791851185  M1M2_CDNS_524688791851185_0
timestamp 1701704242
transform 1 0 2396 0 -1 5647
box 0 0 320 244
use M1M2_CDNS_524688791851185  M1M2_CDNS_524688791851185_1
timestamp 1701704242
transform 1 0 3026 0 -1 5647
box 0 0 320 244
use M1M2_CDNS_524688791851186  M1M2_CDNS_524688791851186_0
timestamp 1701704242
transform 0 -1 7294 -1 0 5118
box 0 0 192 308
use M1M2_CDNS_524688791851186  M1M2_CDNS_524688791851186_1
timestamp 1701704242
transform 0 1 1016 -1 0 2861
box 0 0 192 308
use M1M2_CDNS_524688791851188  M1M2_CDNS_524688791851188_0
timestamp 1701704242
transform 1 0 841 0 -1 8172
box 0 0 512 116
use M1M2_CDNS_524688791851188  M1M2_CDNS_524688791851188_1
timestamp 1701704242
transform 1 0 841 0 -1 7559
box 0 0 512 116
use M1M2_CDNS_524688791851249  M1M2_CDNS_524688791851249_0
timestamp 1701704242
transform 0 1 12416 -1 0 4429
box 0 0 128 436
use M1M2_CDNS_524688791851250  M1M2_CDNS_524688791851250_0
timestamp 1701704242
transform 1 0 8489 0 -1 8653
box 0 0 448 180
use M1M2_CDNS_524688791851250  M1M2_CDNS_524688791851250_1
timestamp 1701704242
transform 1 0 7519 0 -1 4660
box 0 0 448 180
use M1M2_CDNS_524688791851250  M1M2_CDNS_524688791851250_2
timestamp 1701704242
transform 1 0 7639 0 -1 7030
box 0 0 448 180
use M1M2_CDNS_524688791851250  M1M2_CDNS_524688791851250_3
timestamp 1701704242
transform 1 0 7639 0 -1 9181
box 0 0 448 180
use M1M2_CDNS_524688791851390  M1M2_CDNS_524688791851390_0
timestamp 1701704242
transform 1 0 117 0 -1 5650
box 0 0 384 244
use M1M2_CDNS_524688791851391  M1M2_CDNS_524688791851391_0
timestamp 1701704242
transform 1 0 7519 0 1 5379
box 0 0 576 244
use M1M2_CDNS_524688791851392  M1M2_CDNS_524688791851392_0
timestamp 1701704242
transform 0 -1 11893 -1 0 4429
box 0 0 128 1076
use M1M2_CDNS_524688791851393  M1M2_CDNS_524688791851393_0
timestamp 1701704242
transform 1 0 16095 0 -1 3266
box 0 0 256 372
use M1M2_CDNS_524688791851394  M1M2_CDNS_524688791851394_0
timestamp 1701704242
transform 1 0 4073 0 1 10293
box 0 0 512 244
use sky130_fd_io__sio_com_m2m3_strap  sky130_fd_io__sio_com_m2m3_strap_0
timestamp 1701704242
transform 1 0 982 0 1 3318
box 0 0 364 858
use sky130_fd_io__sio_com_m2m3_strap  sky130_fd_io__sio_com_m2m3_strap_1
timestamp 1701704242
transform 1 0 1025 0 1 9736
box 0 0 364 858
use sky130_fd_io__sio_com_m2m3_strap  sky130_fd_io__sio_com_m2m3_strap_2
timestamp 1701704242
transform 1 0 2850 0 1 3318
box 0 0 364 858
use sky130_fd_io__sio_com_m2m3_strap  sky130_fd_io__sio_com_m2m3_strap_3
timestamp 1701704242
transform 1 0 12522 0 1 4676
box 0 0 364 858
use sky130_fd_io__sio_com_m2m3_strap  sky130_fd_io__sio_com_m2m3_strap_4
timestamp 1701704242
transform 1 0 4156 0 1 4676
box 0 0 364 858
use sky130_fd_io__sio_com_m2m3_strap  sky130_fd_io__sio_com_m2m3_strap_5
timestamp 1701704242
transform 1 0 1025 0 1 8748
box 0 0 364 858
use sky130_fd_io__sio_com_m2m3_strap  sky130_fd_io__sio_com_m2m3_strap_6
timestamp 1701704242
transform 1 0 1025 0 1 7760
box 0 0 364 858
use sky130_fd_io__sio_com_m2m3_strap  sky130_fd_io__sio_com_m2m3_strap_7
timestamp 1701704242
transform 1 0 11567 0 1 4676
box 0 0 364 858
use sky130_fd_io__sio_com_m2m3_strap  sky130_fd_io__sio_com_m2m3_strap_8
timestamp 1701704242
transform 1 0 10781 0 1 4676
box 0 0 364 858
use sky130_fd_io__sio_com_m2m3_strap  sky130_fd_io__sio_com_m2m3_strap_9
timestamp 1701704242
transform 1 0 189 0 1 6034
box 0 0 364 858
use sky130_fd_io__sio_com_m2m3_strap  sky130_fd_io__sio_com_m2m3_strap_10
timestamp 1701704242
transform 1 0 1449 0 1 6034
box 0 0 364 858
use sky130_fd_io__sio_com_m2m3_strap  sky130_fd_io__sio_com_m2m3_strap_11
timestamp 1701704242
transform 1 0 4991 0 1 9736
box 0 0 364 858
use sky130_fd_io__sio_com_m2m3_strap  sky130_fd_io__sio_com_m2m3_strap_12
timestamp 1701704242
transform 1 0 4991 0 1 8748
box 0 0 364 858
use sky130_fd_io__sio_com_m2m3_strap  sky130_fd_io__sio_com_m2m3_strap_13
timestamp 1701704242
transform 1 0 4991 0 1 7760
box 0 0 364 858
use sky130_fd_io__sio_com_m2m3_strap  sky130_fd_io__sio_com_m2m3_strap_14
timestamp 1701704242
transform 1 0 6325 0 1 9736
box 0 0 364 858
use sky130_fd_io__sio_com_m2m3_strap  sky130_fd_io__sio_com_m2m3_strap_15
timestamp 1701704242
transform 1 0 6325 0 1 8748
box 0 0 364 858
use sky130_fd_io__sio_com_m2m3_strap  sky130_fd_io__sio_com_m2m3_strap_16
timestamp 1701704242
transform 1 0 6325 0 1 7760
box 0 0 364 858
use sky130_fd_io__sio_com_m2m3_strap  sky130_fd_io__sio_com_m2m3_strap_17
timestamp 1701704242
transform 1 0 3681 0 1 8748
box 0 0 364 858
use sky130_fd_io__sio_com_m2m3_strap  sky130_fd_io__sio_com_m2m3_strap_18
timestamp 1701704242
transform 1 0 3681 0 1 9736
box 0 0 364 858
use sky130_fd_io__sio_com_m2m3_strap  sky130_fd_io__sio_com_m2m3_strap_19
timestamp 1701704242
transform 1 0 3681 0 1 7760
box 0 0 364 858
use sky130_fd_io__sio_com_m2m3_strap  sky130_fd_io__sio_com_m2m3_strap_20
timestamp 1701704242
transform 1 0 8530 0 1 9736
box 0 0 364 858
use sky130_fd_io__sio_com_m2m3_strap  sky130_fd_io__sio_com_m2m3_strap_21
timestamp 1701704242
transform 1 0 8530 0 1 8748
box 0 0 364 858
use sky130_fd_io__sio_com_m2m3_strap  sky130_fd_io__sio_com_m2m3_strap_22
timestamp 1701704242
transform 1 0 8530 0 1 7760
box 0 0 364 858
use sky130_fd_io__sio_com_m2m3_strap  sky130_fd_io__sio_com_m2m3_strap_23
timestamp 1701704242
transform 1 0 7682 0 1 6034
box 0 0 364 858
use sky130_fd_io__sio_com_m2m3_strap  sky130_fd_io__sio_com_m2m3_strap_24
timestamp 1701704242
transform 1 0 2362 0 1 6034
box 0 0 364 858
use sky130_fd_io__sio_com_m2m3_strap  sky130_fd_io__sio_com_m2m3_strap_25
timestamp 1701704242
transform 1 0 3002 0 1 6034
box 0 0 364 858
use sky130_fd_io__sio_obpredrvr_reg  sky130_fd_io__sio_obpredrvr_reg_0
timestamp 1701704242
transform 1 0 11766 0 -1 8268
box -108 10 2896 2150
use sky130_fd_io__sio_octl_dat  sky130_fd_io__sio_octl_dat_0
timestamp 1701704242
transform 1 0 0 0 1 0
box -185 1361 22297 10673
<< labels >>
flabel metal1 s 16145 1842 16185 2044 3 FreeSans 300 0 0 0 vcc_io
port 13 nsew
flabel metal1 s 12402 6548 12436 6582 7 FreeSans 200 0 0 0 pu_h_n<5>
port 3 nsew
flabel metal1 s 13866 6548 13900 6582 7 FreeSans 200 0 0 0 pu_h_n<4>
port 4 nsew
flabel metal1 s 9206 10236 9206 10236 0 FreeSans 200 270 0 0 pu_h_n<3>
flabel metal1 s 7384 10258 7424 10310 3 FreeSans 300 180 0 0 pu_h_n<2>
port 5 nsew
flabel metal1 s 10024 9375 10064 9427 3 FreeSans 300 180 0 0 pu_h_n<1>
port 6 nsew
flabel metal1 s 7029 10418 7068 10470 3 FreeSans 300 180 0 0 pu_h_n<0>
port 7 nsew
flabel metal1 s 8956 2450 8989 2483 0 FreeSans 200 0 0 0 oe_n
port 8 nsew
flabel metal1 s 10128 2450 10162 2484 0 FreeSans 400 0 0 0 din
port 9 nsew
flabel metal1 s 13507 7367 13541 7401 0 FreeSans 200 0 0 0 slow_h_n
port 10 nsew
flabel metal1 s 12390 4048 12434 4100 7 FreeSans 400 0 0 0 vreg_en_h
port 11 nsew
flabel metal1 s 4972 2286 5009 2320 0 FreeSans 200 0 0 0 hld_i_h_n
port 12 nsew
flabel metal1 s 4071 3667 4105 3701 0 FreeSans 200 0 0 0 vreg_en
port 14 nsew
flabel metal1 s 13960 9516 13980 9536 0 FreeSans 200 0 0 0 pd_h<4>
port 2 nsew
flabel metal3 s 636 4670 888 5487 3 FreeSans 200 0 0 0 vgnd
port 15 nsew
flabel metal3 s 1036 3356 1393 4153 3 FreeSans 200 0 0 0 vpwr
port 16 nsew
flabel metal3 s 273 7783 543 10498 3 FreeSans 200 0 0 0 vgnd_io
port 17 nsew
flabel metal3 s 332 6061 612 6854 0 FreeSans 200 0 0 0 vcc_io
port 13 nsew
flabel locali s 14553 5946 14587 5989 0 FreeSans 200 0 0 0 oe_hs_h
port 18 nsew
flabel metal2 s 15111 4076 15387 4230 7 FreeSans 200 90 0 0 vpwr_ka
port 19 nsew
flabel metal2 s 6875 8821 6927 8873 3 FreeSans 200 0 0 0 drvhi_h
port 20 nsew
flabel metal2 s 13458 9983 13510 10041 3 FreeSans 200 270 0 0 pd_h<3>
port 21 nsew
flabel metal2 s 12015 7235 12067 7281 7 FreeSans 200 90 0 0 puen_reg_h
port 22 nsew
flabel metal2 s 2003 2336 2055 2377 3 FreeSans 200 90 0 0 hld_i_vpwr
port 23 nsew
flabel metal2 s 13375 9984 13427 10041 0 FreeSans 200 90 0 0 pd_h<2>
port 24 nsew
flabel metal2 s 8547 2370 8651 2410 0 FreeSans 100 0 0 0 hld_i_ovr_h
port 25 nsew
flabel metal2 s 1444 2321 1496 2370 3 FreeSans 200 90 0 0 dm_h<0>
port 26 nsew
flabel metal2 s 7335 2432 7463 2464 3 FreeSans 200 90 0 0 od_h
port 27 nsew
flabel metal2 s 2236 2321 2288 2364 3 FreeSans 200 90 0 0 od_h
port 27 nsew
flabel metal2 s 9300 9994 9352 10041 7 FreeSans 200 90 0 0 pd_h<1>
port 28 nsew
flabel metal2 s 8317 9997 8369 10041 7 FreeSans 200 90 0 0 pd_h<0>
port 29 nsew
flabel metal2 s 5884 2321 5936 2364 3 FreeSans 200 90 0 0 dm_h_n<2>
port 30 nsew
flabel metal2 s 2316 2321 2368 2364 3 FreeSans 200 90 0 0 dm_h_n<1>
port 31 nsew
flabel metal2 s 926 2321 978 2370 3 FreeSans 200 90 0 0 dm_h_n<0>
port 32 nsew
flabel metal2 s 5648 2321 5700 2364 3 FreeSans 200 90 0 0 dm_h<2>
port 33 nsew
flabel metal2 s 2552 2321 2604 2364 3 FreeSans 200 90 0 0 dm_h<1>
port 34 nsew
flabel metal2 s 1364 2321 1416 2370 3 FreeSans 200 90 0 0 slow
port 35 nsew
<< properties >>
string GDS_END 88430812
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 88155398
string path 37.700 117.000 37.700 131.600 
<< end >>
