magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< metal3 >>
rect 0 1190 544 1196
rect 0 0 544 6
<< via3 >>
rect 0 6 544 1190
<< metal4 >>
rect -1 1190 545 1191
rect -1 6 0 1190
rect 544 6 545 1190
rect -1 5 545 6
<< properties >>
string GDS_END 93362692
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 93355840
<< end >>
