magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -38 261 1234 582
<< pwell >>
rect 1 21 1169 203
rect 29 -17 63 21
<< scnmos >>
rect 82 47 112 177
rect 166 47 196 177
rect 250 47 280 177
rect 334 47 364 177
rect 530 47 560 177
rect 614 47 644 177
rect 698 47 728 177
rect 789 47 819 177
rect 977 47 1007 177
rect 1061 47 1091 177
<< scpmoshvt >>
rect 82 297 112 497
rect 166 297 196 497
rect 250 297 280 497
rect 334 297 364 497
rect 530 297 560 497
rect 614 297 644 497
rect 698 297 728 497
rect 789 297 819 497
rect 977 297 1007 497
rect 1061 297 1091 497
<< ndiff >>
rect 27 95 82 177
rect 27 61 38 95
rect 72 61 82 95
rect 27 47 82 61
rect 112 163 166 177
rect 112 129 122 163
rect 156 129 166 163
rect 112 47 166 129
rect 196 163 250 177
rect 196 129 206 163
rect 240 129 250 163
rect 196 95 250 129
rect 196 61 206 95
rect 240 61 250 95
rect 196 47 250 61
rect 280 95 334 177
rect 280 61 290 95
rect 324 61 334 95
rect 280 47 334 61
rect 364 163 420 177
rect 364 129 374 163
rect 408 129 420 163
rect 364 95 420 129
rect 364 61 374 95
rect 408 61 420 95
rect 364 47 420 61
rect 474 163 530 177
rect 474 129 486 163
rect 520 129 530 163
rect 474 95 530 129
rect 474 61 486 95
rect 520 61 530 95
rect 474 47 530 61
rect 560 163 614 177
rect 560 129 570 163
rect 604 129 614 163
rect 560 95 614 129
rect 560 61 570 95
rect 604 61 614 95
rect 560 47 614 61
rect 644 95 698 177
rect 644 61 654 95
rect 688 61 698 95
rect 644 47 698 61
rect 728 163 789 177
rect 728 129 745 163
rect 779 129 789 163
rect 728 95 789 129
rect 728 61 745 95
rect 779 61 789 95
rect 728 47 789 61
rect 819 95 871 177
rect 819 61 829 95
rect 863 61 871 95
rect 819 47 871 61
rect 925 95 977 177
rect 925 61 933 95
rect 967 61 977 95
rect 925 47 977 61
rect 1007 163 1061 177
rect 1007 129 1017 163
rect 1051 129 1061 163
rect 1007 47 1061 129
rect 1091 163 1143 177
rect 1091 129 1101 163
rect 1135 129 1143 163
rect 1091 95 1143 129
rect 1091 61 1101 95
rect 1135 61 1143 95
rect 1091 47 1143 61
<< pdiff >>
rect 27 477 82 497
rect 27 443 38 477
rect 72 443 82 477
rect 27 409 82 443
rect 27 375 38 409
rect 72 375 82 409
rect 27 297 82 375
rect 112 477 166 497
rect 112 443 122 477
rect 156 443 166 477
rect 112 297 166 443
rect 196 477 250 497
rect 196 443 206 477
rect 240 443 250 477
rect 196 409 250 443
rect 196 375 206 409
rect 240 375 250 409
rect 196 297 250 375
rect 280 477 334 497
rect 280 443 290 477
rect 324 443 334 477
rect 280 297 334 443
rect 364 477 420 497
rect 364 443 374 477
rect 408 443 420 477
rect 364 409 420 443
rect 364 375 374 409
rect 408 375 420 409
rect 364 297 420 375
rect 474 477 530 497
rect 474 443 486 477
rect 520 443 530 477
rect 474 297 530 443
rect 560 477 614 497
rect 560 443 570 477
rect 604 443 614 477
rect 560 297 614 443
rect 644 477 698 497
rect 644 443 654 477
rect 688 443 698 477
rect 644 297 698 443
rect 728 409 789 497
rect 728 375 745 409
rect 779 375 789 409
rect 728 297 789 375
rect 819 477 871 497
rect 819 443 829 477
rect 863 443 871 477
rect 819 297 871 443
rect 925 477 977 497
rect 925 443 933 477
rect 967 443 977 477
rect 925 297 977 443
rect 1007 409 1061 497
rect 1007 375 1017 409
rect 1051 375 1061 409
rect 1007 341 1061 375
rect 1007 307 1017 341
rect 1051 307 1061 341
rect 1007 297 1061 307
rect 1091 477 1147 497
rect 1091 443 1101 477
rect 1135 443 1147 477
rect 1091 409 1147 443
rect 1091 375 1101 409
rect 1135 375 1147 409
rect 1091 297 1147 375
<< ndiffc >>
rect 38 61 72 95
rect 122 129 156 163
rect 206 129 240 163
rect 206 61 240 95
rect 290 61 324 95
rect 374 129 408 163
rect 374 61 408 95
rect 486 129 520 163
rect 486 61 520 95
rect 570 129 604 163
rect 570 61 604 95
rect 654 61 688 95
rect 745 129 779 163
rect 745 61 779 95
rect 829 61 863 95
rect 933 61 967 95
rect 1017 129 1051 163
rect 1101 129 1135 163
rect 1101 61 1135 95
<< pdiffc >>
rect 38 443 72 477
rect 38 375 72 409
rect 122 443 156 477
rect 206 443 240 477
rect 206 375 240 409
rect 290 443 324 477
rect 374 443 408 477
rect 374 375 408 409
rect 486 443 520 477
rect 570 443 604 477
rect 654 443 688 477
rect 745 375 779 409
rect 829 443 863 477
rect 933 443 967 477
rect 1017 375 1051 409
rect 1017 307 1051 341
rect 1101 443 1135 477
rect 1101 375 1135 409
<< poly >>
rect 82 497 112 523
rect 166 497 196 523
rect 250 497 280 523
rect 334 497 364 523
rect 530 497 560 523
rect 614 497 644 523
rect 698 497 728 523
rect 789 497 819 523
rect 977 497 1007 523
rect 1061 497 1091 523
rect 82 265 112 297
rect 166 265 196 297
rect 82 249 196 265
rect 82 215 113 249
rect 147 215 196 249
rect 82 199 196 215
rect 82 177 112 199
rect 166 177 196 199
rect 250 265 280 297
rect 334 265 364 297
rect 530 265 560 297
rect 614 265 644 297
rect 250 249 644 265
rect 250 215 267 249
rect 301 215 335 249
rect 369 215 403 249
rect 437 215 475 249
rect 509 215 644 249
rect 250 199 644 215
rect 250 177 280 199
rect 334 177 364 199
rect 530 177 560 199
rect 614 177 644 199
rect 698 265 728 297
rect 789 265 819 297
rect 698 249 819 265
rect 698 215 734 249
rect 768 215 819 249
rect 698 199 819 215
rect 698 177 728 199
rect 789 177 819 199
rect 977 265 1007 297
rect 1061 265 1091 297
rect 977 249 1091 265
rect 977 215 1009 249
rect 1043 215 1091 249
rect 977 199 1091 215
rect 977 177 1007 199
rect 1061 177 1091 199
rect 82 21 112 47
rect 166 21 196 47
rect 250 21 280 47
rect 334 21 364 47
rect 530 21 560 47
rect 614 21 644 47
rect 698 21 728 47
rect 789 21 819 47
rect 977 21 1007 47
rect 1061 21 1091 47
<< polycont >>
rect 113 215 147 249
rect 267 215 301 249
rect 335 215 369 249
rect 403 215 437 249
rect 475 215 509 249
rect 734 215 768 249
rect 1009 215 1043 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 17 477 80 493
rect 17 443 38 477
rect 72 443 80 477
rect 17 409 80 443
rect 114 477 164 527
rect 114 443 122 477
rect 156 443 164 477
rect 114 427 164 443
rect 198 477 248 493
rect 198 443 206 477
rect 240 443 248 477
rect 17 375 38 409
rect 72 393 80 409
rect 198 409 248 443
rect 282 477 332 527
rect 282 443 290 477
rect 324 443 332 477
rect 282 427 332 443
rect 366 477 416 493
rect 366 443 374 477
rect 408 443 416 477
rect 198 393 206 409
rect 72 375 206 393
rect 240 393 248 409
rect 366 409 416 443
rect 478 477 528 493
rect 478 443 486 477
rect 520 459 528 477
rect 478 425 493 443
rect 527 425 528 459
rect 562 477 612 527
rect 562 443 570 477
rect 604 443 612 477
rect 562 427 612 443
rect 646 477 871 493
rect 646 443 654 477
rect 688 459 829 477
rect 646 425 677 443
rect 821 443 829 459
rect 863 443 871 477
rect 821 427 871 443
rect 925 477 975 527
rect 925 443 933 477
rect 967 443 975 477
rect 925 427 975 443
rect 1093 477 1179 527
rect 1093 443 1101 477
rect 1135 443 1179 477
rect 366 393 374 409
rect 240 375 374 393
rect 408 391 416 409
rect 745 409 787 425
rect 408 375 696 391
rect 17 357 696 375
rect 779 393 787 409
rect 1009 409 1059 425
rect 1009 393 1017 409
rect 779 375 1017 393
rect 1051 375 1059 409
rect 745 359 1059 375
rect 1093 409 1179 443
rect 1093 375 1101 409
rect 1135 375 1179 409
rect 1093 359 1179 375
rect 17 179 63 357
rect 662 325 696 357
rect 1009 341 1059 359
rect 158 289 620 323
rect 662 291 961 325
rect 158 257 192 289
rect 97 249 192 257
rect 586 257 620 289
rect 97 215 113 249
rect 147 215 192 249
rect 251 249 541 255
rect 251 215 267 249
rect 301 215 335 249
rect 369 215 403 249
rect 437 215 475 249
rect 509 215 541 249
rect 586 249 791 257
rect 586 215 734 249
rect 768 215 791 249
rect 927 249 961 291
rect 1009 307 1017 341
rect 1051 325 1059 341
rect 1051 307 1179 325
rect 1009 283 1179 307
rect 927 215 1009 249
rect 1043 215 1059 249
rect 17 163 172 179
rect 17 129 122 163
rect 156 129 172 163
rect 206 163 424 181
rect 240 145 374 163
rect 240 129 256 145
rect 206 95 256 129
rect 358 129 374 145
rect 408 129 424 163
rect 21 61 38 95
rect 72 61 206 95
rect 240 61 256 95
rect 21 51 256 61
rect 290 95 324 111
rect 290 17 324 61
rect 358 95 424 129
rect 358 61 374 95
rect 408 61 424 95
rect 358 51 424 61
rect 486 163 520 181
rect 486 95 520 129
rect 486 17 520 61
rect 554 163 1067 181
rect 554 129 570 163
rect 604 145 745 163
rect 604 129 620 145
rect 554 95 620 129
rect 722 129 745 145
rect 779 145 1017 163
rect 779 129 795 145
rect 1001 129 1017 145
rect 1051 129 1067 163
rect 1101 163 1179 283
rect 1135 129 1179 163
rect 554 61 570 95
rect 604 61 620 95
rect 554 51 620 61
rect 654 95 688 111
rect 654 17 688 61
rect 722 95 795 129
rect 722 61 745 95
rect 779 61 795 95
rect 722 51 795 61
rect 829 95 863 111
rect 1101 95 1179 129
rect 917 61 933 95
rect 967 61 1101 95
rect 1135 61 1179 95
rect 829 17 863 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 493 443 520 459
rect 520 443 527 459
rect 493 425 527 443
rect 677 443 688 459
rect 688 443 711 459
rect 677 425 711 443
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 481 459 539 465
rect 481 425 493 459
rect 527 456 539 459
rect 665 459 723 465
rect 665 456 677 459
rect 527 428 677 456
rect 527 425 539 428
rect 481 419 539 425
rect 665 425 677 428
rect 711 425 723 459
rect 665 419 723 425
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< labels >>
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel locali s 1141 289 1175 323 0 FreeSans 400 0 0 0 Y
port 7 nsew signal output
flabel locali s 397 221 431 255 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 213 289 247 323 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 xnor2_2
rlabel metal1 s 0 -48 1196 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1196 592 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1196 544
string GDS_END 626992
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 618312
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 2.720 5.980 2.720 
<< end >>
