magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< nwell >>
rect 6630 124 6846 534
rect 6952 124 7168 534
rect 6630 96 7168 124
rect 6654 -370 7086 96
<< pwell >>
rect 18 1429 714 1681
rect 72 1328 714 1429
rect 72 10 724 1328
<< mvnmos >>
rect 97 1455 197 1655
rect 379 1455 479 1655
rect 535 1455 635 1655
rect 98 1149 698 1249
rect 98 993 698 1093
rect 98 837 698 937
rect 98 681 698 781
rect 98 525 698 625
rect 98 369 698 469
rect 98 89 698 189
<< mvpmos >>
rect 6696 215 6780 415
rect 7018 215 7102 415
rect 6720 -95 7020 5
rect 6720 -251 7020 -151
<< mvndiff >>
rect 44 1643 97 1655
rect 44 1609 52 1643
rect 86 1609 97 1643
rect 44 1575 97 1609
rect 44 1541 52 1575
rect 86 1541 97 1575
rect 44 1507 97 1541
rect 44 1473 52 1507
rect 86 1473 97 1507
rect 44 1455 97 1473
rect 197 1643 250 1655
rect 197 1609 208 1643
rect 242 1609 250 1643
rect 197 1575 250 1609
rect 197 1541 208 1575
rect 242 1541 250 1575
rect 197 1507 250 1541
rect 197 1473 208 1507
rect 242 1473 250 1507
rect 197 1455 250 1473
rect 326 1643 379 1655
rect 326 1609 334 1643
rect 368 1609 379 1643
rect 326 1575 379 1609
rect 326 1541 334 1575
rect 368 1541 379 1575
rect 326 1507 379 1541
rect 326 1473 334 1507
rect 368 1473 379 1507
rect 326 1455 379 1473
rect 479 1643 535 1655
rect 479 1609 490 1643
rect 524 1609 535 1643
rect 479 1575 535 1609
rect 479 1541 490 1575
rect 524 1541 535 1575
rect 479 1507 535 1541
rect 479 1473 490 1507
rect 524 1473 535 1507
rect 479 1455 535 1473
rect 635 1643 688 1655
rect 635 1609 646 1643
rect 680 1609 688 1643
rect 635 1575 688 1609
rect 635 1541 646 1575
rect 680 1541 688 1575
rect 635 1507 688 1541
rect 635 1473 646 1507
rect 680 1473 688 1507
rect 635 1455 688 1473
rect 98 1294 698 1302
rect 98 1260 176 1294
rect 210 1260 244 1294
rect 278 1260 312 1294
rect 346 1260 380 1294
rect 414 1260 448 1294
rect 482 1260 516 1294
rect 550 1260 584 1294
rect 618 1260 652 1294
rect 686 1260 698 1294
rect 98 1249 698 1260
rect 98 1138 698 1149
rect 98 1104 176 1138
rect 210 1104 244 1138
rect 278 1104 312 1138
rect 346 1104 380 1138
rect 414 1104 448 1138
rect 482 1104 516 1138
rect 550 1104 584 1138
rect 618 1104 652 1138
rect 686 1104 698 1138
rect 98 1093 698 1104
rect 98 982 698 993
rect 98 948 176 982
rect 210 948 244 982
rect 278 948 312 982
rect 346 948 380 982
rect 414 948 448 982
rect 482 948 516 982
rect 550 948 584 982
rect 618 948 652 982
rect 686 948 698 982
rect 98 937 698 948
rect 98 826 698 837
rect 98 792 176 826
rect 210 792 244 826
rect 278 792 312 826
rect 346 792 380 826
rect 414 792 448 826
rect 482 792 516 826
rect 550 792 584 826
rect 618 792 652 826
rect 686 792 698 826
rect 98 781 698 792
rect 98 670 698 681
rect 98 636 176 670
rect 210 636 244 670
rect 278 636 312 670
rect 346 636 380 670
rect 414 636 448 670
rect 482 636 516 670
rect 550 636 584 670
rect 618 636 652 670
rect 686 636 698 670
rect 98 625 698 636
rect 98 514 698 525
rect 98 480 176 514
rect 210 480 244 514
rect 278 480 312 514
rect 346 480 380 514
rect 414 480 448 514
rect 482 480 516 514
rect 550 480 584 514
rect 618 480 652 514
rect 686 480 698 514
rect 98 469 698 480
rect 98 358 698 369
rect 98 324 176 358
rect 210 324 244 358
rect 278 324 312 358
rect 346 324 380 358
rect 414 324 448 358
rect 482 324 516 358
rect 550 324 584 358
rect 618 324 652 358
rect 686 324 698 358
rect 98 316 698 324
rect 98 234 698 242
rect 98 200 176 234
rect 210 200 244 234
rect 278 200 312 234
rect 346 200 380 234
rect 414 200 448 234
rect 482 200 516 234
rect 550 200 584 234
rect 618 200 652 234
rect 686 200 698 234
rect 98 189 698 200
rect 98 78 698 89
rect 98 44 176 78
rect 210 44 244 78
rect 278 44 312 78
rect 346 44 380 78
rect 414 44 448 78
rect 482 44 516 78
rect 550 44 584 78
rect 618 44 652 78
rect 686 44 698 78
rect 98 36 698 44
<< mvpdiff >>
rect 6696 460 6780 468
rect 6696 426 6708 460
rect 6742 426 6780 460
rect 6696 415 6780 426
rect 7018 460 7102 468
rect 7018 426 7030 460
rect 7064 426 7102 460
rect 7018 415 7102 426
rect 6696 204 6780 215
rect 6696 170 6708 204
rect 6742 170 6780 204
rect 6696 162 6780 170
rect 7018 204 7102 215
rect 7018 170 7030 204
rect 7064 170 7102 204
rect 7018 162 7102 170
rect 6720 50 7020 58
rect 6720 16 6732 50
rect 6766 16 6800 50
rect 6834 16 6868 50
rect 6902 16 6936 50
rect 6970 16 7020 50
rect 6720 5 7020 16
rect 6720 -106 7020 -95
rect 6720 -140 6732 -106
rect 6766 -140 6800 -106
rect 6834 -140 6868 -106
rect 6902 -140 6936 -106
rect 6970 -140 7020 -106
rect 6720 -151 7020 -140
rect 6720 -262 7020 -251
rect 6720 -296 6732 -262
rect 6766 -296 6800 -262
rect 6834 -296 6868 -262
rect 6902 -296 6936 -262
rect 6970 -296 7020 -262
rect 6720 -304 7020 -296
<< mvndiffc >>
rect 52 1609 86 1643
rect 52 1541 86 1575
rect 52 1473 86 1507
rect 208 1609 242 1643
rect 208 1541 242 1575
rect 208 1473 242 1507
rect 334 1609 368 1643
rect 334 1541 368 1575
rect 334 1473 368 1507
rect 490 1609 524 1643
rect 490 1541 524 1575
rect 490 1473 524 1507
rect 646 1609 680 1643
rect 646 1541 680 1575
rect 646 1473 680 1507
rect 176 1260 210 1294
rect 244 1260 278 1294
rect 312 1260 346 1294
rect 380 1260 414 1294
rect 448 1260 482 1294
rect 516 1260 550 1294
rect 584 1260 618 1294
rect 652 1260 686 1294
rect 176 1104 210 1138
rect 244 1104 278 1138
rect 312 1104 346 1138
rect 380 1104 414 1138
rect 448 1104 482 1138
rect 516 1104 550 1138
rect 584 1104 618 1138
rect 652 1104 686 1138
rect 176 948 210 982
rect 244 948 278 982
rect 312 948 346 982
rect 380 948 414 982
rect 448 948 482 982
rect 516 948 550 982
rect 584 948 618 982
rect 652 948 686 982
rect 176 792 210 826
rect 244 792 278 826
rect 312 792 346 826
rect 380 792 414 826
rect 448 792 482 826
rect 516 792 550 826
rect 584 792 618 826
rect 652 792 686 826
rect 176 636 210 670
rect 244 636 278 670
rect 312 636 346 670
rect 380 636 414 670
rect 448 636 482 670
rect 516 636 550 670
rect 584 636 618 670
rect 652 636 686 670
rect 176 480 210 514
rect 244 480 278 514
rect 312 480 346 514
rect 380 480 414 514
rect 448 480 482 514
rect 516 480 550 514
rect 584 480 618 514
rect 652 480 686 514
rect 176 324 210 358
rect 244 324 278 358
rect 312 324 346 358
rect 380 324 414 358
rect 448 324 482 358
rect 516 324 550 358
rect 584 324 618 358
rect 652 324 686 358
rect 176 200 210 234
rect 244 200 278 234
rect 312 200 346 234
rect 380 200 414 234
rect 448 200 482 234
rect 516 200 550 234
rect 584 200 618 234
rect 652 200 686 234
rect 176 44 210 78
rect 244 44 278 78
rect 312 44 346 78
rect 380 44 414 78
rect 448 44 482 78
rect 516 44 550 78
rect 584 44 618 78
rect 652 44 686 78
<< mvpdiffc >>
rect 6708 426 6742 460
rect 7030 426 7064 460
rect 6708 170 6742 204
rect 7030 170 7064 204
rect 6732 16 6766 50
rect 6800 16 6834 50
rect 6868 16 6902 50
rect 6936 16 6970 50
rect 6732 -140 6766 -106
rect 6800 -140 6834 -106
rect 6868 -140 6902 -106
rect 6936 -140 6970 -106
rect 6732 -296 6766 -262
rect 6800 -296 6834 -262
rect 6868 -296 6902 -262
rect 6936 -296 6970 -262
<< poly >>
rect 97 1655 197 1687
rect 379 1655 479 1687
rect 535 1655 635 1687
rect 97 1423 197 1455
rect 379 1423 479 1455
rect 50 1407 197 1423
rect 50 1373 66 1407
rect 100 1373 147 1407
rect 181 1373 197 1407
rect 50 1357 197 1373
rect 345 1407 479 1423
rect 345 1373 361 1407
rect 395 1373 429 1407
rect 463 1373 479 1407
rect 345 1357 479 1373
rect 535 1423 635 1455
rect 535 1407 669 1423
rect 535 1373 551 1407
rect 585 1373 619 1407
rect 653 1373 669 1407
rect 535 1357 669 1373
rect 0 1233 98 1249
rect 0 1199 16 1233
rect 50 1199 98 1233
rect 0 1164 98 1199
rect 0 1130 16 1164
rect 50 1149 98 1164
rect 698 1149 730 1249
rect 50 1130 66 1149
rect 0 1095 66 1130
rect 0 1061 16 1095
rect 50 1093 66 1095
rect 50 1061 98 1093
rect 0 1026 98 1061
rect 0 992 16 1026
rect 50 993 98 1026
rect 698 993 730 1093
rect 50 992 66 993
rect 0 957 66 992
rect 0 923 16 957
rect 50 937 66 957
rect 50 923 98 937
rect 0 887 98 923
rect 0 853 16 887
rect 50 853 98 887
rect 0 837 98 853
rect 698 837 730 937
rect 0 765 98 781
rect 0 731 16 765
rect 50 731 98 765
rect 0 696 98 731
rect 0 662 16 696
rect 50 681 98 696
rect 698 681 730 781
rect 50 662 66 681
rect 0 627 66 662
rect 0 593 16 627
rect 50 625 66 627
rect 50 593 98 625
rect 0 558 98 593
rect 0 524 16 558
rect 50 525 98 558
rect 698 525 730 625
rect 50 524 66 525
rect 0 489 66 524
rect 0 455 16 489
rect 50 469 66 489
rect 50 455 98 469
rect 0 419 98 455
rect 0 385 16 419
rect 50 385 98 419
rect 0 369 98 385
rect 698 369 730 469
rect 0 190 66 206
rect 0 156 16 190
rect 50 189 66 190
rect 6664 215 6696 415
rect 6780 399 6878 415
rect 6780 365 6828 399
rect 6862 365 6878 399
rect 6780 265 6878 365
rect 6780 231 6828 265
rect 6862 231 6878 265
rect 6780 215 6878 231
rect 6920 399 7018 415
rect 6920 365 6936 399
rect 6970 365 7018 399
rect 6920 265 7018 365
rect 6920 231 6936 265
rect 6970 231 7018 265
rect 6920 215 7018 231
rect 7102 215 7134 415
rect 50 156 98 189
rect 0 122 98 156
rect 0 88 16 122
rect 50 89 98 122
rect 698 89 730 189
rect 50 88 66 89
rect 0 72 66 88
rect 7052 23 7118 39
rect 7052 5 7068 23
rect 6688 -95 6720 5
rect 7020 -11 7068 5
rect 7102 -11 7118 23
rect 7020 -45 7118 -11
rect 7020 -79 7068 -45
rect 7102 -79 7118 -45
rect 7020 -95 7118 -79
rect 6688 -251 6720 -151
rect 7020 -167 7118 -151
rect 7020 -201 7068 -167
rect 7102 -201 7118 -167
rect 7020 -235 7118 -201
rect 7020 -251 7068 -235
rect 7052 -269 7068 -251
rect 7102 -269 7118 -235
rect 7052 -285 7118 -269
<< polycont >>
rect 66 1373 100 1407
rect 147 1373 181 1407
rect 361 1373 395 1407
rect 429 1373 463 1407
rect 551 1373 585 1407
rect 619 1373 653 1407
rect 16 1199 50 1233
rect 16 1130 50 1164
rect 16 1061 50 1095
rect 16 992 50 1026
rect 16 923 50 957
rect 16 853 50 887
rect 16 731 50 765
rect 16 662 50 696
rect 16 593 50 627
rect 16 524 50 558
rect 16 455 50 489
rect 16 385 50 419
rect 16 156 50 190
rect 6828 365 6862 399
rect 6828 231 6862 265
rect 6936 365 6970 399
rect 6936 231 6970 265
rect 16 88 50 122
rect 7068 -11 7102 23
rect 7068 -79 7102 -45
rect 7068 -201 7102 -167
rect 7068 -269 7102 -235
<< locali >>
rect -126 1703 567 1761
rect 52 1643 86 1659
rect 52 1575 86 1609
rect 52 1507 86 1541
rect 52 1457 86 1469
rect 208 1643 292 1659
rect 242 1609 292 1643
rect 208 1575 292 1609
rect 242 1541 292 1575
rect 208 1507 292 1541
rect 242 1473 292 1507
rect 208 1457 292 1473
rect 334 1647 368 1659
rect 334 1575 368 1609
rect 334 1507 368 1541
rect 334 1457 368 1469
rect 460 1643 567 1703
rect 460 1609 490 1643
rect 524 1609 567 1643
rect 460 1575 567 1609
rect 460 1541 490 1575
rect 524 1541 567 1575
rect 460 1507 567 1541
rect 460 1473 490 1507
rect 524 1473 567 1507
rect 460 1457 567 1473
rect 646 1647 680 1659
rect 646 1575 680 1609
rect 646 1507 680 1541
rect 646 1457 680 1469
rect 252 1413 292 1457
rect 252 1407 479 1413
rect 50 1373 66 1407
rect 108 1373 147 1407
rect 252 1373 357 1407
rect 395 1373 429 1407
rect 467 1373 479 1407
rect 535 1373 547 1407
rect 585 1373 619 1407
rect 657 1373 669 1407
rect 160 1260 176 1294
rect 210 1260 244 1294
rect 278 1260 312 1294
rect 346 1260 380 1294
rect 414 1260 448 1294
rect 482 1260 516 1294
rect 550 1260 584 1294
rect 630 1260 652 1294
rect 16 1233 50 1249
rect 16 1164 50 1199
rect 16 1095 50 1130
rect 160 1104 176 1138
rect 238 1104 244 1138
rect 310 1104 312 1138
rect 346 1104 380 1138
rect 414 1104 448 1138
rect 482 1104 516 1138
rect 550 1104 584 1138
rect 618 1104 652 1138
rect 686 1104 702 1138
rect 16 1026 50 1061
rect 16 957 50 992
rect 160 948 176 982
rect 210 948 244 982
rect 278 948 312 982
rect 346 948 380 982
rect 414 948 448 982
rect 482 948 516 982
rect 550 948 584 982
rect 630 948 652 982
rect 16 887 50 923
rect 16 837 50 853
rect 160 792 176 826
rect 238 792 244 826
rect 310 792 312 826
rect 346 792 380 826
rect 414 792 448 826
rect 482 792 516 826
rect 550 792 584 826
rect 618 792 652 826
rect 686 792 702 826
rect 16 765 50 781
rect 16 696 50 731
rect 16 627 50 662
rect 160 636 176 670
rect 210 636 244 670
rect 278 636 312 670
rect 346 636 380 670
rect 414 636 448 670
rect 550 636 554 670
rect 618 636 652 670
rect 686 636 702 670
rect 16 558 50 593
rect 16 489 50 524
rect 160 480 176 514
rect 238 480 244 514
rect 310 480 312 514
rect 346 480 380 514
rect 414 480 448 514
rect 482 480 516 514
rect 550 480 584 514
rect 618 480 652 514
rect 686 480 702 514
rect 16 419 50 455
rect 6692 426 6708 460
rect 6742 426 6758 460
rect 7014 426 7030 460
rect 7064 426 7080 460
rect 16 369 50 385
rect 6828 399 6862 415
rect 160 324 176 358
rect 210 324 244 358
rect 278 324 312 358
rect 346 324 380 358
rect 414 324 448 358
rect 550 324 554 358
rect 618 324 652 358
rect 686 324 702 358
rect 6828 334 6862 365
rect 6928 399 6978 415
rect 6928 365 6936 399
rect 6970 365 6978 399
rect 6828 300 6834 334
rect 16 190 50 206
rect 160 200 176 234
rect 238 200 244 234
rect 310 200 312 234
rect 346 200 380 234
rect 414 200 448 234
rect 482 200 516 234
rect 550 200 584 234
rect 618 200 652 234
rect 686 200 702 234
rect 6747 204 6781 242
rect 6828 265 6868 300
rect 6862 262 6868 265
rect 6828 228 6834 231
rect 6928 265 6978 365
rect 6928 231 6936 265
rect 6970 231 6978 265
rect 6828 215 6862 228
rect 6692 170 6708 204
rect 6742 170 6747 204
rect 6928 179 6978 231
rect 7037 204 7071 242
rect 6781 170 6978 179
rect 7014 170 7030 204
rect 7071 170 7080 204
rect 16 122 74 156
rect 50 118 74 122
rect 6699 121 6978 170
rect 16 84 40 88
rect 16 72 50 84
rect 159 44 176 78
rect 210 44 244 78
rect 278 44 312 78
rect 346 44 380 78
rect 414 44 448 78
rect 482 44 516 78
rect 550 44 584 78
rect 618 44 652 78
rect 686 44 702 78
rect 159 30 702 44
rect -126 -31 702 30
rect 6716 16 6732 50
rect 6766 16 6800 50
rect 6834 16 6836 50
rect 6902 16 6908 50
rect 6970 16 6986 50
rect 7068 23 7102 39
rect 7068 -45 7102 -11
rect 7068 -95 7102 -83
rect 6716 -140 6732 -106
rect 6766 -140 6800 -106
rect 6834 -140 6868 -106
rect 6902 -140 6936 -106
rect 6970 -140 6986 -106
rect 7068 -167 7102 -151
rect 7068 -235 7102 -201
rect 6716 -296 6732 -262
rect 6766 -296 6778 -262
rect 6834 -296 6850 -262
rect 6902 -296 6936 -262
rect 6970 -296 6986 -262
rect 7102 -269 7126 -251
rect 7088 -285 7126 -269
<< viali >>
rect 52 1541 86 1575
rect 52 1473 86 1503
rect 52 1469 86 1473
rect 334 1643 368 1647
rect 334 1613 368 1643
rect 334 1541 368 1575
rect 334 1473 368 1503
rect 334 1469 368 1473
rect 646 1643 680 1647
rect 646 1613 680 1643
rect 646 1541 680 1575
rect 646 1473 680 1503
rect 646 1469 680 1473
rect 74 1373 100 1407
rect 100 1373 108 1407
rect 163 1373 181 1407
rect 181 1373 197 1407
rect 357 1373 361 1407
rect 361 1373 391 1407
rect 433 1373 463 1407
rect 463 1373 467 1407
rect 547 1373 551 1407
rect 551 1373 581 1407
rect 623 1373 653 1407
rect 653 1373 657 1407
rect 596 1260 618 1294
rect 618 1260 630 1294
rect 668 1260 686 1294
rect 686 1260 702 1294
rect 204 1104 210 1138
rect 210 1104 238 1138
rect 276 1104 278 1138
rect 278 1104 310 1138
rect 596 948 618 982
rect 618 948 630 982
rect 668 948 686 982
rect 686 948 702 982
rect 204 792 210 826
rect 210 792 238 826
rect 276 792 278 826
rect 278 792 310 826
rect 482 636 516 670
rect 554 636 584 670
rect 584 636 588 670
rect 204 480 210 514
rect 210 480 238 514
rect 276 480 278 514
rect 278 480 310 514
rect 482 324 516 358
rect 554 324 584 358
rect 584 324 588 358
rect 6834 300 6868 334
rect 6747 242 6781 276
rect 204 200 210 234
rect 210 200 238 234
rect 276 200 278 234
rect 278 200 310 234
rect 6834 231 6862 262
rect 6862 231 6868 262
rect 6834 228 6868 231
rect 40 156 50 190
rect 50 156 74 190
rect 6747 170 6781 204
rect 7037 242 7071 276
rect 7037 170 7064 204
rect 7064 170 7071 204
rect 40 88 50 118
rect 50 88 74 118
rect 40 84 74 88
rect 6836 16 6868 50
rect 6868 16 6870 50
rect 6908 16 6936 50
rect 6936 16 6942 50
rect 7068 -11 7102 23
rect 7068 -79 7102 -49
rect 7068 -83 7102 -79
rect 6778 -296 6800 -262
rect 6800 -296 6812 -262
rect 6850 -296 6868 -262
rect 6868 -296 6884 -262
rect 7054 -269 7068 -251
rect 7068 -269 7088 -251
rect 7054 -285 7088 -269
rect 7126 -285 7160 -251
<< metal1 >>
rect 267 1647 374 1659
rect 267 1613 334 1647
rect 368 1613 374 1647
rect -95 1575 92 1587
rect -95 1541 52 1575
rect 86 1541 92 1575
rect -95 1503 92 1541
rect -95 1469 52 1503
rect 86 1469 92 1503
rect -95 1457 92 1469
rect 267 1575 374 1613
rect 267 1541 334 1575
rect 368 1541 374 1575
rect 267 1503 374 1541
rect 267 1469 334 1503
rect 368 1469 374 1503
rect 267 1457 374 1469
rect 640 1647 780 1659
rect 640 1613 646 1647
rect 680 1613 780 1647
rect 640 1575 780 1613
rect 640 1541 646 1575
rect 680 1541 780 1575
rect 640 1503 780 1541
rect 640 1469 646 1503
rect 680 1469 780 1503
rect 640 1457 780 1469
tri 1 1407 7 1413 se
rect 7 1407 209 1413
tri -33 1373 1 1407 se
rect 1 1373 74 1407
rect 108 1373 163 1407
rect 197 1373 209 1407
tri -39 1367 -33 1373 se
rect -33 1367 209 1373
tri -54 1352 -39 1367 se
rect -39 1352 7 1367
tri 7 1352 22 1367 nw
tri -58 1348 -54 1352 se
rect -54 1348 3 1352
tri 3 1348 7 1352 nw
rect -58 1256 -20 1348
tri -20 1325 3 1348 nw
tri -58 1255 -57 1256 ne
rect -57 1255 -20 1256
rect 267 1263 315 1457
tri 315 1431 341 1457 nw
tri 709 1431 735 1457 ne
rect 735 1431 780 1457
tri 735 1424 742 1431 ne
rect 345 1407 495 1413
rect 345 1373 357 1407
rect 391 1373 433 1407
rect 467 1373 495 1407
rect 345 1367 495 1373
rect 535 1407 669 1413
rect 535 1373 547 1407
rect 581 1373 623 1407
rect 657 1406 669 1407
rect 657 1373 714 1406
rect 535 1367 714 1373
tri 378 1330 415 1367 ne
tri 315 1263 340 1288 sw
rect 267 1260 340 1263
tri 340 1260 343 1263 sw
rect 415 1260 495 1367
tri 547 1330 584 1367 ne
rect 584 1294 714 1367
tri 495 1260 521 1286 sw
rect 584 1260 596 1294
rect 630 1260 668 1294
rect 702 1260 714 1294
rect 267 1255 343 1260
tri 343 1255 348 1260 sw
rect 415 1255 521 1260
tri -57 1249 -51 1255 ne
tri -58 1063 -51 1070 se
rect -51 1063 -20 1255
tri 270 1185 340 1255 ne
rect 340 1252 348 1255
tri 348 1252 351 1255 sw
tri 415 1252 418 1255 ne
rect 418 1252 521 1255
rect 340 1231 351 1252
tri 351 1231 372 1252 sw
tri 418 1231 439 1252 ne
rect 439 1231 521 1252
tri 521 1231 550 1260 sw
rect 340 1200 372 1231
tri 372 1200 403 1231 sw
tri 439 1200 470 1231 ne
rect 340 1185 403 1200
tri 403 1185 418 1200 sw
tri 340 1155 370 1185 ne
rect -58 -47 -20 1063
rect 192 1138 322 1144
rect 192 1104 204 1138
rect 238 1104 276 1138
rect 310 1104 322 1138
rect 192 826 322 1104
rect 192 792 204 826
rect 238 792 276 826
rect 310 792 322 826
rect 192 514 322 792
rect 192 480 204 514
rect 238 480 276 514
rect 310 480 322 514
rect 192 234 322 480
rect 34 190 80 202
rect 192 200 204 234
rect 238 200 276 234
rect 310 200 322 234
rect 192 194 322 200
rect 34 156 40 190
rect 74 156 80 190
rect 34 118 80 156
rect 34 84 40 118
rect 74 84 80 118
rect 34 -129 80 84
rect 370 14 418 1185
rect 470 679 550 1231
rect 584 982 714 1260
rect 584 948 596 982
rect 630 948 668 982
rect 702 948 714 982
rect 584 942 714 948
tri 627 907 662 942 ne
tri 550 679 600 729 sw
rect 470 670 600 679
rect 470 636 482 670
rect 516 636 554 670
rect 588 636 600 670
rect 470 358 600 636
rect 470 324 482 358
rect 516 324 554 358
rect 588 324 600 358
rect 470 318 600 324
tri 507 300 525 318 ne
rect 525 300 600 318
tri 525 277 548 300 ne
rect 370 8 422 14
rect 370 -64 422 -44
rect 370 -122 422 -116
rect 548 8 600 300
rect 548 -64 600 -44
rect 548 -122 600 -116
rect 662 8 714 942
rect 662 -64 714 -44
rect 662 -122 714 -116
rect 742 14 780 1431
rect 6828 334 6874 346
rect 6828 300 6834 334
rect 6868 300 6874 334
rect 6828 288 6874 300
rect 6741 276 6787 288
rect 6741 242 6747 276
rect 6781 242 6787 276
rect 6741 204 6787 242
rect 6828 276 7085 288
rect 6828 262 7037 276
rect 6828 228 6834 262
rect 6868 242 7037 262
rect 7071 242 7085 276
rect 6868 228 7085 242
rect 6828 216 7085 228
rect 6741 170 6747 204
rect 6781 170 6787 204
rect 742 8 794 14
rect 742 -64 794 -44
rect 742 -122 794 -116
rect 6741 -154 6787 170
rect 6985 204 7085 216
rect 6985 170 7037 204
rect 7071 170 7085 204
rect 6985 158 7085 170
rect 6824 50 6954 56
rect 6824 16 6836 50
rect 6870 16 6908 50
rect 6942 16 6954 50
rect 6824 -70 6954 16
rect 6824 -122 6830 -70
rect 6882 -122 6894 -70
rect 6946 -122 6952 -70
tri 6787 -154 6815 -126 sw
rect 6741 -206 6747 -154
rect 6799 -206 6811 -154
rect 6863 -206 6869 -154
rect 6985 -242 7031 158
tri 7031 110 7079 158 nw
rect 7061 23 7113 35
rect 7061 -11 7068 23
rect 7102 -11 7113 23
rect 7061 -49 7113 -11
rect 7061 -83 7068 -49
rect 7102 -83 7113 -49
rect 7061 -84 7113 -83
rect 7061 -148 7113 -136
rect 7061 -206 7113 -200
tri 7031 -242 7042 -231 sw
rect 6766 -262 6896 -256
rect 6766 -296 6778 -262
rect 6812 -296 6850 -262
rect 6884 -296 6896 -262
rect 6985 -294 7048 -242
rect 7100 -294 7114 -242
rect 7166 -294 7172 -242
rect 6766 -324 6896 -296
rect 6766 -376 6774 -324
rect 6826 -376 6838 -324
rect 6890 -376 6896 -324
<< via1 >>
rect 370 -44 422 8
rect 370 -116 422 -64
rect 548 -44 600 8
rect 548 -116 600 -64
rect 662 -44 714 8
rect 662 -116 714 -64
rect 742 -44 794 8
rect 742 -116 794 -64
rect 6830 -122 6882 -70
rect 6894 -122 6946 -70
rect 6747 -206 6799 -154
rect 6811 -206 6863 -154
rect 7061 -136 7113 -84
rect 7061 -200 7113 -148
rect 7048 -251 7100 -242
rect 7048 -285 7054 -251
rect 7054 -285 7088 -251
rect 7088 -285 7100 -251
rect 7048 -294 7100 -285
rect 7114 -251 7166 -242
rect 7114 -285 7126 -251
rect 7126 -285 7160 -251
rect 7160 -285 7166 -251
rect 7114 -294 7166 -285
rect 6774 -376 6826 -324
rect 6838 -376 6890 -324
<< metal2 >>
rect 370 8 422 14
rect 370 -64 422 -44
rect 370 -294 422 -116
rect 548 8 600 14
rect 548 -64 600 -44
rect 548 -242 600 -116
rect 662 8 714 14
rect 662 -64 714 -44
rect 662 -148 714 -116
rect 742 8 794 14
rect 742 -64 794 -44
tri 794 -70 833 -31 sw
rect 794 -116 6830 -70
rect 742 -122 6830 -116
rect 6882 -122 6894 -70
rect 6946 -122 6952 -70
rect 7061 -84 7113 -78
tri 714 -148 726 -136 sw
rect 7061 -148 7113 -136
rect 662 -154 726 -148
tri 726 -154 732 -148 sw
rect 662 -185 6747 -154
tri 662 -206 683 -185 ne
rect 683 -206 6747 -185
rect 6799 -206 6811 -154
rect 6863 -200 7061 -154
rect 6863 -206 7113 -200
tri 600 -242 634 -208 sw
rect 548 -271 7048 -242
tri 548 -275 552 -271 ne
rect 552 -275 7048 -271
tri 422 -294 441 -275 sw
tri 552 -294 571 -275 ne
rect 571 -294 7048 -275
rect 7100 -294 7114 -242
rect 7166 -294 7172 -242
rect 370 -324 441 -294
tri 441 -324 471 -294 sw
rect 370 -344 6774 -324
tri 370 -376 402 -344 ne
rect 402 -376 6774 -344
rect 6826 -376 6838 -324
rect 6890 -376 6896 -324
use sky130_fd_pr__nfet_01v8__example_55959141808474  sky130_fd_pr__nfet_01v8__example_55959141808474_0
timestamp 1701704242
transform 1 0 97 0 -1 1655
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808483  sky130_fd_pr__nfet_01v8__example_55959141808483_0
timestamp 1701704242
transform 0 -1 698 1 0 369
box -1 0 881 1
use sky130_fd_pr__nfet_01v8__example_55959141808484  sky130_fd_pr__nfet_01v8__example_55959141808484_0
timestamp 1701704242
transform 0 -1 698 1 0 89
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808485  sky130_fd_pr__nfet_01v8__example_55959141808485_0
timestamp 1701704242
transform 1 0 379 0 -1 1655
box -1 0 257 1
use sky130_fd_pr__pfet_01v8__example_55959141808481  sky130_fd_pr__pfet_01v8__example_55959141808481_0
timestamp 1701704242
transform 0 1 6720 -1 0 -151
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808481  sky130_fd_pr__pfet_01v8__example_55959141808481_1
timestamp 1701704242
transform 0 1 6720 1 0 -95
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808482  sky130_fd_pr__pfet_01v8__example_55959141808482_0
timestamp 1701704242
transform 0 1 7018 -1 0 415
box -1 0 201 1
use sky130_fd_pr__pfet_01v8__example_55959141808482  sky130_fd_pr__pfet_01v8__example_55959141808482_1
timestamp 1701704242
transform 0 1 6696 -1 0 415
box -1 0 201 1
<< labels >>
flabel comment s 571 -38 571 -38 0 FreeSans 400 90 0 0 FBK
flabel comment s 391 -54 391 -54 0 FreeSans 400 90 0 0 OUT_H_N
<< properties >>
string GDS_END 64790902
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 64775598
<< end >>
