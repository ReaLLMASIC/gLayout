magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< pwell >>
rect -76 -26 1388 2026
<< mvnnmos >>
rect 0 0 400 2000
rect 456 0 856 2000
rect 912 0 1312 2000
<< mvndiff >>
rect -50 0 0 2000
rect 1312 0 1362 2000
<< poly >>
rect 0 2000 400 2026
rect 0 -26 400 0
rect 456 2000 856 2026
rect 456 -26 856 0
rect 912 2000 1312 2026
rect 912 -26 1312 0
<< metal1 >>
rect -51 -16 -5 1986
rect 405 -16 451 1986
rect 861 -16 907 1986
rect 1317 -16 1363 1986
use DFM1sd_CDNS_524688791851117  DFM1sd_CDNS_524688791851117_0
timestamp 1701704242
transform -1 0 0 0 1 0
box -26 -26 79 2026
use DFM1sd_CDNS_524688791851117  DFM1sd_CDNS_524688791851117_1
timestamp 1701704242
transform 1 0 1312 0 1 0
box -26 -26 79 2026
use hvDFM1sd2_CDNS_5246887918552  hvDFM1sd2_CDNS_5246887918552_0
timestamp 1701704242
transform 1 0 856 0 1 0
box -26 -26 82 2026
use hvDFM1sd2_CDNS_5246887918552  hvDFM1sd2_CDNS_5246887918552_1
timestamp 1701704242
transform 1 0 400 0 1 0
box -26 -26 82 2026
<< labels >>
flabel comment s -28 985 -28 985 0 FreeSans 300 0 0 0 S
flabel comment s 428 985 428 985 0 FreeSans 300 0 0 0 D
flabel comment s 884 985 884 985 0 FreeSans 300 0 0 0 S
flabel comment s 1340 985 1340 985 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 78947006
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 78945056
<< end >>
