magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< nwell >>
rect 21 1714 965 1822
rect -44 1498 1013 1714
rect -44 1382 839 1498
<< pwell >>
rect 207 1128 933 1254
rect 33 992 933 1128
rect 207 720 933 992
rect 33 536 933 720
rect -17 202 933 536
<< mvnmos >>
rect 112 1018 212 1102
rect 112 610 212 694
rect 286 228 386 1228
rect 442 228 542 1228
rect 598 228 698 1228
rect 754 228 854 1228
<< mvpmos >>
rect 72 1448 192 1648
rect 248 1448 368 1648
rect 424 1448 544 1648
rect 600 1448 720 1648
rect 794 1564 894 1648
<< mvndiff >>
rect 233 1158 286 1228
rect 233 1124 241 1158
rect 275 1124 286 1158
rect 233 1102 286 1124
rect 59 1090 112 1102
rect 59 1056 67 1090
rect 101 1056 112 1090
rect 59 1018 112 1056
rect 212 1090 286 1102
rect 212 1056 241 1090
rect 275 1056 286 1090
rect 212 1022 286 1056
rect 212 1018 241 1022
rect 233 988 241 1018
rect 275 988 286 1022
rect 233 954 286 988
rect 233 920 241 954
rect 275 920 286 954
rect 233 886 286 920
rect 233 852 241 886
rect 275 852 286 886
rect 233 818 286 852
rect 233 784 241 818
rect 275 784 286 818
rect 233 750 286 784
rect 233 716 241 750
rect 275 716 286 750
rect 233 694 286 716
rect 59 682 112 694
rect 59 648 67 682
rect 101 648 112 682
rect 59 610 112 648
rect 212 682 286 694
rect 212 648 241 682
rect 275 648 286 682
rect 212 614 286 648
rect 212 610 241 614
rect 233 580 241 610
rect 275 580 286 614
rect 233 546 286 580
rect 233 512 241 546
rect 275 512 286 546
rect 233 478 286 512
rect 233 444 241 478
rect 275 444 286 478
rect 233 410 286 444
rect 233 376 241 410
rect 275 376 286 410
rect 233 342 286 376
rect 233 308 241 342
rect 275 308 286 342
rect 233 274 286 308
rect 233 240 241 274
rect 275 240 286 274
rect 233 228 286 240
rect 386 1158 442 1228
rect 386 1124 397 1158
rect 431 1124 442 1158
rect 386 1090 442 1124
rect 386 1056 397 1090
rect 431 1056 442 1090
rect 386 1022 442 1056
rect 386 988 397 1022
rect 431 988 442 1022
rect 386 954 442 988
rect 386 920 397 954
rect 431 920 442 954
rect 386 886 442 920
rect 386 852 397 886
rect 431 852 442 886
rect 386 818 442 852
rect 386 784 397 818
rect 431 784 442 818
rect 386 750 442 784
rect 386 716 397 750
rect 431 716 442 750
rect 386 682 442 716
rect 386 648 397 682
rect 431 648 442 682
rect 386 614 442 648
rect 386 580 397 614
rect 431 580 442 614
rect 386 546 442 580
rect 386 512 397 546
rect 431 512 442 546
rect 386 478 442 512
rect 386 444 397 478
rect 431 444 442 478
rect 386 410 442 444
rect 386 376 397 410
rect 431 376 442 410
rect 386 342 442 376
rect 386 308 397 342
rect 431 308 442 342
rect 386 274 442 308
rect 386 240 397 274
rect 431 240 442 274
rect 386 228 442 240
rect 542 1158 598 1228
rect 542 1124 553 1158
rect 587 1124 598 1158
rect 542 1090 598 1124
rect 542 1056 553 1090
rect 587 1056 598 1090
rect 542 1022 598 1056
rect 542 988 553 1022
rect 587 988 598 1022
rect 542 954 598 988
rect 542 920 553 954
rect 587 920 598 954
rect 542 886 598 920
rect 542 852 553 886
rect 587 852 598 886
rect 542 818 598 852
rect 542 784 553 818
rect 587 784 598 818
rect 542 750 598 784
rect 542 716 553 750
rect 587 716 598 750
rect 542 682 598 716
rect 542 648 553 682
rect 587 648 598 682
rect 542 614 598 648
rect 542 580 553 614
rect 587 580 598 614
rect 542 546 598 580
rect 542 512 553 546
rect 587 512 598 546
rect 542 478 598 512
rect 542 444 553 478
rect 587 444 598 478
rect 542 410 598 444
rect 542 376 553 410
rect 587 376 598 410
rect 542 342 598 376
rect 542 308 553 342
rect 587 308 598 342
rect 542 274 598 308
rect 542 240 553 274
rect 587 240 598 274
rect 542 228 598 240
rect 698 1158 754 1228
rect 698 1124 709 1158
rect 743 1124 754 1158
rect 698 1090 754 1124
rect 698 1056 709 1090
rect 743 1056 754 1090
rect 698 1022 754 1056
rect 698 988 709 1022
rect 743 988 754 1022
rect 698 954 754 988
rect 698 920 709 954
rect 743 920 754 954
rect 698 886 754 920
rect 698 852 709 886
rect 743 852 754 886
rect 698 818 754 852
rect 698 784 709 818
rect 743 784 754 818
rect 698 750 754 784
rect 698 716 709 750
rect 743 716 754 750
rect 698 682 754 716
rect 698 648 709 682
rect 743 648 754 682
rect 698 614 754 648
rect 698 580 709 614
rect 743 580 754 614
rect 698 546 754 580
rect 698 512 709 546
rect 743 512 754 546
rect 698 478 754 512
rect 698 444 709 478
rect 743 444 754 478
rect 698 410 754 444
rect 698 376 709 410
rect 743 376 754 410
rect 698 342 754 376
rect 698 308 709 342
rect 743 308 754 342
rect 698 274 754 308
rect 698 240 709 274
rect 743 240 754 274
rect 698 228 754 240
rect 854 1158 907 1228
rect 854 1124 865 1158
rect 899 1124 907 1158
rect 854 1090 907 1124
rect 854 1056 865 1090
rect 899 1056 907 1090
rect 854 1022 907 1056
rect 854 988 865 1022
rect 899 988 907 1022
rect 854 954 907 988
rect 854 920 865 954
rect 899 920 907 954
rect 854 886 907 920
rect 854 852 865 886
rect 899 852 907 886
rect 854 818 907 852
rect 854 784 865 818
rect 899 784 907 818
rect 854 750 907 784
rect 854 716 865 750
rect 899 716 907 750
rect 854 682 907 716
rect 854 648 865 682
rect 899 648 907 682
rect 854 614 907 648
rect 854 580 865 614
rect 899 580 907 614
rect 854 546 907 580
rect 854 512 865 546
rect 899 512 907 546
rect 854 478 907 512
rect 854 444 865 478
rect 899 444 907 478
rect 854 410 907 444
rect 854 376 865 410
rect 899 376 907 410
rect 854 342 907 376
rect 854 308 865 342
rect 899 308 907 342
rect 854 274 907 308
rect 854 240 865 274
rect 899 240 907 274
rect 854 228 907 240
<< mvpdiff >>
rect 1 1636 72 1648
rect 1 1602 9 1636
rect 43 1602 72 1636
rect 1 1568 72 1602
rect 1 1534 9 1568
rect 43 1534 72 1568
rect 1 1500 72 1534
rect 1 1466 9 1500
rect 43 1466 72 1500
rect 1 1454 72 1466
rect 22 1448 72 1454
rect 192 1636 248 1648
rect 192 1602 203 1636
rect 237 1602 248 1636
rect 192 1568 248 1602
rect 192 1534 203 1568
rect 237 1534 248 1568
rect 192 1500 248 1534
rect 192 1466 203 1500
rect 237 1466 248 1500
rect 192 1448 248 1466
rect 368 1636 424 1648
rect 368 1602 379 1636
rect 413 1602 424 1636
rect 368 1568 424 1602
rect 368 1534 379 1568
rect 413 1534 424 1568
rect 368 1500 424 1534
rect 368 1466 379 1500
rect 413 1466 424 1500
rect 368 1448 424 1466
rect 544 1636 600 1648
rect 544 1602 555 1636
rect 589 1602 600 1636
rect 544 1568 600 1602
rect 544 1534 555 1568
rect 589 1534 600 1568
rect 544 1500 600 1534
rect 544 1466 555 1500
rect 589 1466 600 1500
rect 544 1448 600 1466
rect 720 1636 794 1648
rect 720 1602 731 1636
rect 765 1602 794 1636
rect 720 1568 794 1602
rect 720 1534 731 1568
rect 765 1564 794 1568
rect 894 1636 947 1648
rect 894 1602 905 1636
rect 939 1602 947 1636
rect 894 1564 947 1602
rect 765 1534 773 1564
rect 720 1500 773 1534
rect 720 1466 731 1500
rect 765 1466 773 1500
rect 720 1448 773 1466
<< mvndiffc >>
rect 241 1124 275 1158
rect 67 1056 101 1090
rect 241 1056 275 1090
rect 241 988 275 1022
rect 241 920 275 954
rect 241 852 275 886
rect 241 784 275 818
rect 241 716 275 750
rect 67 648 101 682
rect 241 648 275 682
rect 241 580 275 614
rect 241 512 275 546
rect 241 444 275 478
rect 241 376 275 410
rect 241 308 275 342
rect 241 240 275 274
rect 397 1124 431 1158
rect 397 1056 431 1090
rect 397 988 431 1022
rect 397 920 431 954
rect 397 852 431 886
rect 397 784 431 818
rect 397 716 431 750
rect 397 648 431 682
rect 397 580 431 614
rect 397 512 431 546
rect 397 444 431 478
rect 397 376 431 410
rect 397 308 431 342
rect 397 240 431 274
rect 553 1124 587 1158
rect 553 1056 587 1090
rect 553 988 587 1022
rect 553 920 587 954
rect 553 852 587 886
rect 553 784 587 818
rect 553 716 587 750
rect 553 648 587 682
rect 553 580 587 614
rect 553 512 587 546
rect 553 444 587 478
rect 553 376 587 410
rect 553 308 587 342
rect 553 240 587 274
rect 709 1124 743 1158
rect 709 1056 743 1090
rect 709 988 743 1022
rect 709 920 743 954
rect 709 852 743 886
rect 709 784 743 818
rect 709 716 743 750
rect 709 648 743 682
rect 709 580 743 614
rect 709 512 743 546
rect 709 444 743 478
rect 709 376 743 410
rect 709 308 743 342
rect 709 240 743 274
rect 865 1124 899 1158
rect 865 1056 899 1090
rect 865 988 899 1022
rect 865 920 899 954
rect 865 852 899 886
rect 865 784 899 818
rect 865 716 899 750
rect 865 648 899 682
rect 865 580 899 614
rect 865 512 899 546
rect 865 444 899 478
rect 865 376 899 410
rect 865 308 899 342
rect 865 240 899 274
<< mvpdiffc >>
rect 9 1602 43 1636
rect 9 1534 43 1568
rect 9 1466 43 1500
rect 203 1602 237 1636
rect 203 1534 237 1568
rect 203 1466 237 1500
rect 379 1602 413 1636
rect 379 1534 413 1568
rect 379 1466 413 1500
rect 555 1602 589 1636
rect 555 1534 589 1568
rect 555 1466 589 1500
rect 731 1602 765 1636
rect 731 1534 765 1568
rect 905 1602 939 1636
rect 731 1466 765 1500
<< psubdiff >>
rect 9 486 149 510
rect 43 452 115 486
rect 9 386 149 452
rect 43 352 115 386
rect 9 286 149 352
rect 43 252 115 286
rect 9 228 149 252
<< mvnsubdiff >>
rect 87 1722 111 1756
rect 145 1722 184 1756
rect 218 1722 257 1756
rect 291 1722 330 1756
rect 364 1722 403 1756
rect 437 1722 476 1756
rect 510 1722 549 1756
rect 583 1722 622 1756
rect 656 1722 695 1756
rect 729 1722 768 1756
rect 802 1722 841 1756
rect 875 1722 899 1756
<< psubdiffcont >>
rect 9 452 43 486
rect 115 452 149 486
rect 9 352 43 386
rect 115 352 149 386
rect 9 252 43 286
rect 115 252 149 286
<< mvnsubdiffcont >>
rect 111 1722 145 1756
rect 184 1722 218 1756
rect 257 1722 291 1756
rect 330 1722 364 1756
rect 403 1722 437 1756
rect 476 1722 510 1756
rect 549 1722 583 1756
rect 622 1722 656 1756
rect 695 1722 729 1756
rect 768 1722 802 1756
rect 841 1722 875 1756
<< poly >>
rect 72 1648 192 1680
rect 248 1648 368 1680
rect 424 1648 544 1680
rect 600 1648 720 1680
rect 794 1648 894 1680
rect 794 1515 894 1564
rect 794 1481 836 1515
rect 870 1481 894 1515
rect 72 1416 192 1448
rect 248 1416 368 1448
rect 72 1400 368 1416
rect 72 1366 88 1400
rect 122 1366 165 1400
rect 199 1366 242 1400
rect 276 1366 318 1400
rect 352 1366 368 1400
rect 72 1350 368 1366
rect 424 1416 544 1448
rect 600 1416 720 1448
rect 424 1400 720 1416
rect 424 1366 440 1400
rect 474 1366 516 1400
rect 550 1366 593 1400
rect 627 1366 670 1400
rect 704 1366 720 1400
rect 794 1447 894 1481
rect 794 1413 836 1447
rect 870 1413 894 1447
rect 794 1397 894 1413
rect 424 1350 720 1366
rect 112 1271 212 1288
rect 112 1237 145 1271
rect 179 1237 212 1271
rect 112 1203 212 1237
rect 286 1228 386 1260
rect 442 1228 542 1260
rect 598 1228 698 1260
rect 754 1228 854 1260
rect 112 1169 145 1203
rect 179 1169 212 1203
rect 112 1102 212 1169
rect 112 986 212 1018
rect 112 863 212 880
rect 112 829 145 863
rect 179 829 212 863
rect 112 795 212 829
rect 112 761 145 795
rect 179 761 212 795
rect 112 694 212 761
rect 112 578 212 610
rect 286 158 386 228
rect 286 124 319 158
rect 353 124 386 158
rect 286 90 386 124
rect 286 56 319 90
rect 353 56 386 90
rect 286 40 386 56
rect 442 158 542 228
rect 442 124 479 158
rect 513 124 542 158
rect 442 90 542 124
rect 442 56 479 90
rect 513 56 542 90
rect 442 40 542 56
rect 598 158 698 228
rect 598 124 629 158
rect 663 124 698 158
rect 598 90 698 124
rect 598 56 629 90
rect 663 56 698 90
rect 598 40 698 56
rect 754 156 854 228
rect 754 122 784 156
rect 818 122 854 156
rect 754 88 854 122
rect 754 54 784 88
rect 818 54 854 88
rect 754 38 854 54
<< polycont >>
rect 836 1481 870 1515
rect 88 1366 122 1400
rect 165 1366 199 1400
rect 242 1366 276 1400
rect 318 1366 352 1400
rect 440 1366 474 1400
rect 516 1366 550 1400
rect 593 1366 627 1400
rect 670 1366 704 1400
rect 836 1413 870 1447
rect 145 1237 179 1271
rect 145 1169 179 1203
rect 145 829 179 863
rect 145 761 179 795
rect 319 124 353 158
rect 319 56 353 90
rect 479 124 513 158
rect 479 56 513 90
rect 629 124 663 158
rect 629 56 663 90
rect 784 122 818 156
rect 784 54 818 88
<< locali >>
rect 87 1722 111 1756
rect 145 1724 146 1756
rect 180 1756 222 1758
rect 180 1724 184 1756
rect 145 1722 184 1724
rect 218 1724 222 1756
rect 256 1756 298 1758
rect 332 1756 374 1758
rect 408 1756 450 1758
rect 484 1756 526 1758
rect 560 1756 602 1758
rect 636 1756 678 1758
rect 712 1756 754 1758
rect 788 1756 831 1758
rect 256 1724 257 1756
rect 218 1722 257 1724
rect 291 1724 298 1756
rect 364 1724 374 1756
rect 437 1724 450 1756
rect 510 1724 526 1756
rect 583 1724 602 1756
rect 656 1724 678 1756
rect 729 1724 754 1756
rect 802 1724 831 1756
rect 291 1722 330 1724
rect 364 1722 403 1724
rect 437 1722 476 1724
rect 510 1722 549 1724
rect 583 1722 622 1724
rect 656 1722 695 1724
rect 729 1722 768 1724
rect 802 1722 841 1724
rect 875 1722 899 1756
rect 9 1638 43 1652
rect 9 1568 43 1602
rect 9 1500 43 1534
rect 9 1450 43 1462
rect 203 1580 237 1602
rect 203 1508 237 1534
rect 203 1450 237 1466
rect 379 1580 413 1602
rect 379 1508 413 1534
rect 379 1450 413 1466
rect 555 1580 589 1602
rect 555 1508 589 1534
rect 555 1450 589 1466
rect 867 1618 905 1652
rect 731 1580 765 1602
rect 905 1586 939 1602
rect 731 1508 765 1534
rect 731 1450 765 1466
rect 816 1522 831 1549
rect 865 1522 939 1549
rect 816 1515 939 1522
rect 816 1484 836 1515
rect 816 1450 831 1484
rect 870 1481 939 1515
rect 865 1450 939 1481
rect 816 1447 939 1450
rect 816 1413 836 1447
rect 870 1413 939 1447
rect 72 1366 88 1400
rect 122 1366 165 1400
rect 199 1366 242 1400
rect 276 1366 318 1400
rect 352 1366 368 1400
rect 424 1366 440 1400
rect 474 1366 516 1400
rect 550 1366 593 1400
rect 627 1366 670 1400
rect 704 1366 722 1400
rect 816 1397 939 1413
rect 127 1285 165 1319
rect 199 1285 225 1319
rect 93 1271 225 1285
rect 93 1237 145 1271
rect 179 1237 225 1271
rect 93 1205 225 1237
rect 93 1203 203 1205
rect 93 1169 145 1203
rect 179 1169 203 1203
rect 309 1181 363 1366
rect 424 1356 722 1366
rect 424 1322 436 1356
rect 470 1322 526 1356
rect 560 1322 616 1356
rect 650 1325 722 1356
rect 650 1322 678 1325
rect 424 1316 678 1322
rect 732 1248 770 1282
rect 93 1153 203 1169
rect 67 1034 101 1056
rect 139 1038 203 1153
rect 139 1004 163 1038
rect 197 1004 203 1038
rect 139 966 203 1004
rect 139 932 163 966
rect 197 932 203 966
rect 241 1158 275 1174
rect 241 1092 275 1124
rect 309 1147 320 1181
rect 354 1147 363 1181
rect 309 1109 363 1147
rect 309 1075 320 1109
rect 354 1075 363 1109
rect 309 1074 363 1075
rect 397 1158 431 1160
rect 397 1122 431 1124
rect 241 1022 275 1056
rect 241 954 275 984
rect 241 886 275 910
rect 66 845 67 879
rect 101 863 203 879
rect 101 845 145 863
rect 66 829 145 845
rect 179 829 203 863
rect 66 807 203 829
rect 66 773 67 807
rect 101 795 203 807
rect 101 773 145 795
rect 66 761 145 773
rect 179 761 203 795
rect 66 745 203 761
rect 241 818 275 836
rect 241 750 275 761
rect 67 626 101 648
rect 241 682 275 686
rect 241 645 275 648
rect 241 570 275 580
rect 43 486 129 510
rect 43 452 115 486
rect 149 452 163 476
rect 9 426 163 452
rect 43 392 129 426
rect 9 386 163 392
rect 43 352 115 386
rect 149 352 163 386
rect 9 342 163 352
rect 43 308 129 342
rect 9 286 163 308
rect 43 252 115 286
rect 149 258 163 286
rect 43 224 129 252
rect 241 495 275 512
rect 241 420 275 444
rect 241 345 275 376
rect 241 274 275 308
rect 241 224 275 236
rect 397 1050 431 1056
rect 397 978 431 988
rect 397 906 431 920
rect 397 834 431 852
rect 397 762 431 784
rect 397 690 431 716
rect 397 618 431 648
rect 397 546 431 580
rect 397 478 431 512
rect 397 410 431 440
rect 397 342 431 368
rect 397 274 431 296
rect 553 1158 587 1160
rect 553 1122 587 1124
rect 553 1050 587 1056
rect 553 978 587 988
rect 553 906 587 920
rect 553 834 587 852
rect 553 762 587 784
rect 553 690 587 716
rect 553 618 587 648
rect 553 546 587 580
rect 553 478 587 512
rect 553 410 587 440
rect 553 342 587 368
rect 553 274 587 296
rect 709 1158 743 1160
rect 709 1122 743 1124
rect 709 1050 743 1056
rect 709 978 743 988
rect 709 906 743 920
rect 709 834 743 852
rect 709 762 743 784
rect 709 690 743 716
rect 709 618 743 648
rect 709 546 743 580
rect 709 478 743 512
rect 709 410 743 440
rect 709 342 743 368
rect 709 274 743 296
rect 865 1158 899 1160
rect 865 1122 899 1124
rect 865 1050 899 1056
rect 865 978 899 988
rect 865 906 899 920
rect 865 834 899 852
rect 865 762 899 784
rect 865 690 899 716
rect 865 618 899 648
rect 865 546 899 580
rect 865 478 899 512
rect 865 410 899 440
rect 865 342 899 368
rect 865 274 899 296
rect 319 158 320 174
rect 353 124 354 147
rect 319 109 354 124
rect 319 90 320 109
rect 479 158 513 174
rect 479 90 513 124
rect 319 40 353 56
rect 479 40 513 56
rect 629 158 663 174
rect 629 90 663 124
rect 629 40 663 56
rect 784 156 818 172
rect 784 88 818 122
rect 784 38 818 54
<< viali >>
rect 146 1724 180 1758
rect 222 1724 256 1758
rect 298 1756 332 1758
rect 374 1756 408 1758
rect 450 1756 484 1758
rect 526 1756 560 1758
rect 602 1756 636 1758
rect 678 1756 712 1758
rect 754 1756 788 1758
rect 831 1756 865 1758
rect 298 1724 330 1756
rect 330 1724 332 1756
rect 374 1724 403 1756
rect 403 1724 408 1756
rect 450 1724 476 1756
rect 476 1724 484 1756
rect 526 1724 549 1756
rect 549 1724 560 1756
rect 602 1724 622 1756
rect 622 1724 636 1756
rect 678 1724 695 1756
rect 695 1724 712 1756
rect 754 1724 768 1756
rect 768 1724 788 1756
rect 831 1724 841 1756
rect 841 1724 865 1756
rect 9 1636 43 1638
rect 9 1604 43 1636
rect 9 1466 43 1496
rect 9 1462 43 1466
rect 203 1636 237 1652
rect 203 1618 237 1636
rect 203 1568 237 1580
rect 203 1546 237 1568
rect 203 1500 237 1508
rect 203 1474 237 1500
rect 379 1636 413 1652
rect 379 1618 413 1636
rect 379 1568 413 1580
rect 379 1546 413 1568
rect 379 1500 413 1508
rect 379 1474 413 1500
rect 555 1636 589 1652
rect 555 1618 589 1636
rect 555 1568 589 1580
rect 555 1546 589 1568
rect 555 1500 589 1508
rect 555 1474 589 1500
rect 731 1636 765 1652
rect 731 1618 765 1636
rect 833 1618 867 1652
rect 905 1636 939 1652
rect 905 1618 939 1636
rect 731 1568 765 1580
rect 731 1546 765 1568
rect 731 1500 765 1508
rect 731 1474 765 1500
rect 831 1522 865 1556
rect 831 1481 836 1484
rect 836 1481 865 1484
rect 831 1450 865 1481
rect 93 1285 127 1319
rect 165 1285 199 1319
rect 436 1322 470 1356
rect 526 1322 560 1356
rect 616 1322 650 1356
rect 698 1248 732 1282
rect 770 1248 804 1282
rect 67 1090 101 1106
rect 67 1072 101 1090
rect 67 1000 101 1034
rect 163 1004 197 1038
rect 163 932 197 966
rect 241 1090 275 1092
rect 241 1058 275 1090
rect 320 1147 354 1181
rect 320 1075 354 1109
rect 397 1160 431 1194
rect 397 1090 431 1122
rect 397 1088 431 1090
rect 241 988 275 1018
rect 241 984 275 988
rect 241 920 275 944
rect 241 910 275 920
rect 67 845 101 879
rect 67 773 101 807
rect 241 852 275 870
rect 241 836 275 852
rect 241 784 275 795
rect 241 761 275 784
rect 241 716 275 720
rect 67 682 101 698
rect 67 664 101 682
rect 67 592 101 626
rect 241 686 275 716
rect 241 614 275 645
rect 241 611 275 614
rect 241 546 275 570
rect 241 536 275 546
rect 9 486 43 510
rect 129 486 163 510
rect 9 476 43 486
rect 129 476 149 486
rect 149 476 163 486
rect 9 392 43 426
rect 129 392 163 426
rect 9 308 43 342
rect 129 308 163 342
rect 9 252 43 258
rect 129 252 149 258
rect 149 252 163 258
rect 9 224 43 252
rect 129 224 163 252
rect 241 478 275 495
rect 241 461 275 478
rect 241 410 275 420
rect 241 386 275 410
rect 241 342 275 345
rect 241 311 275 342
rect 241 240 275 270
rect 241 236 275 240
rect 397 1022 431 1050
rect 397 1016 431 1022
rect 397 954 431 978
rect 397 944 431 954
rect 397 886 431 906
rect 397 872 431 886
rect 397 818 431 834
rect 397 800 431 818
rect 397 750 431 762
rect 397 728 431 750
rect 397 682 431 690
rect 397 656 431 682
rect 397 614 431 618
rect 397 584 431 614
rect 397 512 431 546
rect 397 444 431 474
rect 397 440 431 444
rect 397 376 431 402
rect 397 368 431 376
rect 397 308 431 330
rect 397 296 431 308
rect 397 240 431 258
rect 397 224 431 240
rect 553 1160 587 1194
rect 553 1090 587 1122
rect 553 1088 587 1090
rect 553 1022 587 1050
rect 553 1016 587 1022
rect 553 954 587 978
rect 553 944 587 954
rect 553 886 587 906
rect 553 872 587 886
rect 553 818 587 834
rect 553 800 587 818
rect 553 750 587 762
rect 553 728 587 750
rect 553 682 587 690
rect 553 656 587 682
rect 553 614 587 618
rect 553 584 587 614
rect 553 512 587 546
rect 553 444 587 474
rect 553 440 587 444
rect 553 376 587 402
rect 553 368 587 376
rect 553 308 587 330
rect 553 296 587 308
rect 553 240 587 258
rect 553 224 587 240
rect 709 1160 743 1194
rect 709 1090 743 1122
rect 709 1088 743 1090
rect 709 1022 743 1050
rect 709 1016 743 1022
rect 709 954 743 978
rect 709 944 743 954
rect 709 886 743 906
rect 709 872 743 886
rect 709 818 743 834
rect 709 800 743 818
rect 709 750 743 762
rect 709 728 743 750
rect 709 682 743 690
rect 709 656 743 682
rect 709 614 743 618
rect 709 584 743 614
rect 709 512 743 546
rect 709 444 743 474
rect 709 440 743 444
rect 709 376 743 402
rect 709 368 743 376
rect 709 308 743 330
rect 709 296 743 308
rect 709 240 743 258
rect 709 224 743 240
rect 865 1160 899 1194
rect 865 1090 899 1122
rect 865 1088 899 1090
rect 865 1022 899 1050
rect 865 1016 899 1022
rect 865 954 899 978
rect 865 944 899 954
rect 865 886 899 906
rect 865 872 899 886
rect 865 818 899 834
rect 865 800 899 818
rect 865 750 899 762
rect 865 728 899 750
rect 865 682 899 690
rect 865 656 899 682
rect 865 614 899 618
rect 865 584 899 614
rect 865 512 899 546
rect 865 444 899 474
rect 865 440 899 444
rect 865 376 899 402
rect 865 368 899 376
rect 865 308 899 330
rect 865 296 899 308
rect 865 240 899 258
rect 865 224 899 240
rect 320 158 354 181
rect 320 147 353 158
rect 353 147 354 158
rect 320 90 354 109
rect 320 75 353 90
rect 353 75 354 90
<< metal1 >>
rect 21 1758 1000 1803
rect 21 1724 146 1758
rect 180 1724 222 1758
rect 256 1724 298 1758
rect 332 1724 374 1758
rect 408 1724 450 1758
rect 484 1724 526 1758
rect 560 1724 602 1758
rect 636 1724 678 1758
rect 712 1724 754 1758
rect 788 1724 831 1758
rect 865 1724 1000 1758
rect 21 1714 1000 1724
rect 21 1650 67 1714
rect 3 1638 67 1650
rect 3 1604 9 1638
rect 43 1604 67 1638
rect 3 1496 67 1604
rect 3 1462 9 1496
rect 43 1462 67 1496
rect 3 1450 67 1462
rect 197 1652 243 1664
rect 197 1618 203 1652
rect 237 1618 243 1652
rect 197 1580 243 1618
rect 197 1546 203 1580
rect 237 1546 243 1580
rect 197 1508 243 1546
rect 197 1474 203 1508
rect 237 1474 243 1508
tri 151 1362 197 1408 se
rect 197 1391 243 1474
rect 373 1652 419 1714
rect 373 1618 379 1652
rect 413 1618 419 1652
rect 373 1580 419 1618
rect 373 1546 379 1580
rect 413 1546 419 1580
rect 373 1508 419 1546
rect 549 1652 595 1664
rect 549 1618 555 1652
rect 589 1618 595 1652
rect 549 1580 595 1618
rect 549 1546 555 1580
rect 589 1546 595 1580
rect 549 1519 595 1546
rect 373 1474 379 1508
rect 413 1474 419 1508
rect 373 1462 419 1474
rect 543 1513 595 1519
rect 725 1652 771 1714
rect 899 1658 945 1664
rect 725 1618 731 1652
rect 765 1618 771 1652
rect 725 1580 771 1618
rect 821 1652 951 1658
rect 821 1618 833 1652
rect 867 1618 905 1652
rect 939 1618 951 1652
rect 821 1612 951 1618
rect 725 1546 731 1580
rect 765 1546 771 1580
rect 725 1508 771 1546
rect 725 1474 731 1508
rect 765 1474 771 1508
rect 725 1462 771 1474
rect 825 1556 871 1568
rect 825 1522 831 1556
rect 865 1522 871 1556
rect 825 1484 871 1522
rect 543 1449 595 1461
tri 817 1450 825 1458 se
rect 825 1450 831 1484
rect 865 1450 871 1484
tri 243 1391 267 1415 sw
tri 812 1445 817 1450 se
rect 817 1445 871 1450
tri 595 1438 602 1445 sw
tri 805 1438 812 1445 se
rect 812 1438 871 1445
rect 595 1432 602 1438
tri 602 1432 608 1438 sw
tri 799 1432 805 1438 se
rect 805 1432 824 1438
rect 595 1397 824 1432
rect 543 1391 824 1397
tri 824 1391 871 1438 nw
tri 890 1391 899 1400 se
rect 899 1391 945 1612
rect 197 1382 267 1391
tri 267 1382 276 1391 sw
tri 881 1382 890 1391 se
rect 890 1382 945 1391
rect 197 1362 276 1382
tri 276 1362 296 1382 sw
tri 860 1362 880 1382 se
rect 880 1380 945 1382
rect 880 1362 927 1380
tri 927 1362 945 1380 nw
rect 107 1356 905 1362
rect 107 1325 436 1356
rect 81 1322 436 1325
rect 470 1322 526 1356
rect 560 1322 616 1356
rect 650 1322 905 1356
tri 905 1340 927 1362 nw
rect 81 1319 905 1322
rect 81 1285 93 1319
rect 127 1285 165 1319
rect 199 1316 905 1319
rect 199 1288 220 1316
tri 220 1288 248 1316 nw
tri 834 1291 859 1316 ne
rect 199 1286 218 1288
tri 218 1286 220 1288 nw
tri 276 1286 278 1288 se
rect 278 1286 514 1288
rect 199 1285 214 1286
rect 81 1282 214 1285
tri 214 1282 218 1286 nw
tri 272 1282 276 1286 se
rect 276 1282 514 1286
rect 81 1279 211 1282
tri 211 1279 214 1282 nw
tri 269 1279 272 1282 se
rect 272 1279 514 1282
tri 238 1248 269 1279 se
rect 269 1248 514 1279
tri 232 1242 238 1248 se
rect 238 1247 514 1248
rect 238 1242 292 1247
tri 292 1242 297 1247 nw
tri 503 1242 508 1247 ne
tri 226 1236 232 1242 se
rect 232 1236 286 1242
tri 286 1236 292 1242 nw
rect 508 1236 514 1247
rect 566 1236 578 1288
rect 630 1282 816 1288
rect 630 1248 698 1282
rect 732 1248 770 1282
rect 804 1248 816 1282
rect 630 1242 816 1248
rect 630 1236 636 1242
tri 218 1228 226 1236 se
rect 226 1228 278 1236
tri 278 1228 286 1236 nw
tri 184 1194 218 1228 se
rect 218 1194 244 1228
tri 244 1194 278 1228 nw
rect 391 1194 437 1206
tri 183 1193 184 1194 se
rect 184 1193 243 1194
tri 243 1193 244 1194 nw
tri 171 1181 183 1193 se
rect 183 1181 231 1193
tri 231 1181 243 1193 nw
rect 309 1181 363 1193
tri 158 1168 171 1181 se
rect 171 1168 218 1181
tri 218 1168 231 1181 nw
tri 137 1147 158 1168 se
rect 158 1147 197 1168
tri 197 1147 218 1168 nw
rect 309 1147 320 1181
rect 354 1147 363 1181
tri 112 1122 137 1147 se
rect 137 1122 172 1147
tri 172 1122 197 1147 nw
tri 108 1118 112 1122 se
rect 112 1118 168 1122
tri 168 1118 172 1122 nw
rect 61 1109 159 1118
tri 159 1109 168 1118 nw
rect 309 1109 363 1147
rect 61 1106 154 1109
rect 61 1072 67 1106
rect 101 1104 154 1106
tri 154 1104 159 1109 nw
rect 101 1092 142 1104
tri 142 1092 154 1104 nw
rect 235 1092 281 1104
rect 101 1072 108 1092
rect 61 1058 108 1072
tri 108 1058 142 1092 nw
rect 235 1058 241 1092
rect 275 1058 281 1092
rect 61 1034 107 1058
tri 107 1057 108 1058 nw
rect 61 1000 67 1034
rect 101 1000 107 1034
rect 61 879 107 1000
rect 157 1038 203 1050
rect 157 1004 163 1038
rect 197 1004 203 1038
rect 157 966 203 1004
rect 157 932 163 966
rect 197 932 203 966
rect 157 920 203 932
rect 235 1018 281 1058
rect 235 984 241 1018
rect 275 984 281 1018
rect 235 944 281 984
rect 61 845 67 879
rect 101 845 107 879
rect 61 807 107 845
rect 61 773 67 807
rect 101 773 107 807
rect 61 761 107 773
rect 235 910 241 944
rect 275 910 281 944
rect 235 870 281 910
rect 235 836 241 870
rect 275 836 281 870
rect 235 795 281 836
rect 235 761 241 795
rect 275 761 281 795
rect 235 720 281 761
rect 235 710 241 720
rect 61 698 241 710
rect 61 664 67 698
rect 101 686 241 698
rect 275 686 281 720
rect 101 664 281 686
rect 61 645 281 664
rect 61 626 241 645
rect 61 592 67 626
rect 101 611 241 626
rect 275 611 281 645
rect 101 592 281 611
rect 61 580 281 592
rect 235 570 281 580
rect 235 536 241 570
rect 275 536 281 570
rect 235 522 281 536
rect 3 510 281 522
rect 3 476 9 510
rect 43 476 129 510
rect 163 495 281 510
rect 163 476 241 495
rect 3 461 241 476
rect 275 461 281 495
rect 3 426 281 461
rect 3 392 9 426
rect 43 392 129 426
rect 163 420 281 426
rect 163 392 241 420
rect 3 386 241 392
rect 275 386 281 420
rect 3 345 281 386
rect 3 342 241 345
rect 3 308 9 342
rect 43 308 129 342
rect 163 311 241 342
rect 275 311 281 345
rect 163 308 281 311
rect 3 270 281 308
rect 3 258 241 270
rect 3 224 9 258
rect 43 224 129 258
rect 163 236 241 258
rect 275 236 281 270
rect 163 224 281 236
rect 3 212 281 224
rect 309 1075 320 1109
rect 354 1075 363 1109
rect 309 181 363 1075
rect 391 1160 397 1194
rect 431 1160 437 1194
rect 391 1122 437 1160
rect 391 1088 397 1122
rect 431 1088 437 1122
rect 391 1050 437 1088
rect 391 1016 397 1050
rect 431 1016 437 1050
rect 391 978 437 1016
rect 391 944 397 978
rect 431 944 437 978
rect 391 906 437 944
rect 391 872 397 906
rect 431 872 437 906
rect 391 834 437 872
rect 391 800 397 834
rect 431 800 437 834
rect 391 762 437 800
rect 391 728 397 762
rect 431 728 437 762
rect 391 690 437 728
rect 391 656 397 690
rect 431 656 437 690
rect 391 618 437 656
rect 391 584 397 618
rect 431 584 437 618
rect 391 546 437 584
rect 391 512 397 546
rect 431 512 437 546
rect 391 474 437 512
rect 391 440 397 474
rect 431 440 437 474
rect 391 402 437 440
rect 391 368 397 402
rect 431 368 437 402
rect 391 330 437 368
rect 391 296 397 330
rect 431 296 437 330
rect 391 258 437 296
rect 391 224 397 258
rect 431 224 437 258
rect 391 212 437 224
rect 547 1194 593 1206
rect 547 1160 553 1194
rect 587 1160 593 1194
rect 547 1122 593 1160
rect 547 1088 553 1122
rect 587 1088 593 1122
rect 547 1050 593 1088
rect 547 1016 553 1050
rect 587 1016 593 1050
rect 547 978 593 1016
rect 547 944 553 978
rect 587 944 593 978
rect 547 906 593 944
rect 547 872 553 906
rect 587 872 593 906
rect 547 834 593 872
rect 547 800 553 834
rect 587 800 593 834
rect 547 762 593 800
rect 547 728 553 762
rect 587 728 593 762
rect 547 690 593 728
rect 547 656 553 690
rect 587 656 593 690
rect 547 618 593 656
rect 547 584 553 618
rect 587 584 593 618
rect 547 546 593 584
rect 547 512 553 546
rect 587 512 593 546
rect 547 474 593 512
rect 547 440 553 474
rect 587 440 593 474
rect 547 402 593 440
rect 547 368 553 402
rect 587 368 593 402
rect 547 330 593 368
rect 547 296 553 330
rect 587 296 593 330
rect 547 258 593 296
rect 547 224 553 258
rect 587 224 593 258
rect 547 212 593 224
rect 703 1194 749 1206
rect 703 1160 709 1194
rect 743 1160 749 1194
rect 703 1122 749 1160
rect 703 1088 709 1122
rect 743 1088 749 1122
rect 703 1050 749 1088
rect 703 1016 709 1050
rect 743 1016 749 1050
rect 703 978 749 1016
rect 703 944 709 978
rect 743 944 749 978
rect 703 906 749 944
rect 703 872 709 906
rect 743 872 749 906
rect 703 834 749 872
rect 703 800 709 834
rect 743 800 749 834
rect 703 762 749 800
rect 703 728 709 762
rect 743 728 749 762
rect 703 690 749 728
rect 703 656 709 690
rect 743 656 749 690
rect 703 618 749 656
rect 703 584 709 618
rect 743 584 749 618
rect 703 546 749 584
rect 703 512 709 546
rect 743 512 749 546
rect 703 474 749 512
rect 703 440 709 474
rect 743 440 749 474
rect 703 402 749 440
rect 703 368 709 402
rect 743 368 749 402
rect 703 330 749 368
rect 703 296 709 330
rect 743 296 749 330
rect 703 258 749 296
rect 703 224 709 258
rect 743 224 749 258
rect 703 212 749 224
rect 859 1194 905 1316
rect 859 1160 865 1194
rect 899 1160 905 1194
rect 859 1122 905 1160
rect 859 1088 865 1122
rect 899 1088 905 1122
rect 859 1050 905 1088
rect 859 1016 865 1050
rect 899 1016 905 1050
rect 859 978 905 1016
rect 859 944 865 978
rect 899 944 905 978
rect 859 906 905 944
rect 859 872 865 906
rect 899 872 905 906
rect 859 834 905 872
rect 859 800 865 834
rect 899 800 905 834
rect 859 762 905 800
rect 859 728 865 762
rect 899 728 905 762
rect 859 690 905 728
rect 859 656 865 690
rect 899 656 905 690
rect 859 618 905 656
rect 859 584 865 618
rect 899 584 905 618
rect 859 546 905 584
rect 859 512 865 546
rect 899 512 905 546
rect 859 474 905 512
rect 859 440 865 474
rect 899 440 905 474
rect 859 402 905 440
rect 859 368 865 402
rect 899 368 905 402
rect 859 330 905 368
rect 859 296 865 330
rect 899 296 905 330
rect 859 258 905 296
rect 859 224 865 258
rect 899 224 905 258
rect 859 212 905 224
rect 309 147 320 181
rect 354 147 363 181
rect 309 109 363 147
rect 309 75 320 109
rect 354 75 363 109
rect 309 33 363 75
<< via1 >>
rect 543 1508 595 1513
rect 543 1474 555 1508
rect 555 1474 589 1508
rect 589 1474 595 1508
rect 543 1461 595 1474
rect 543 1397 595 1449
rect 514 1236 566 1288
rect 578 1236 630 1288
<< metal2 >>
rect 543 1513 595 1519
rect 543 1449 595 1461
rect 543 1288 595 1397
rect 508 1236 514 1288
rect 566 1236 578 1288
rect 630 1236 636 1288
use sky130_fd_pr__dfl1__example_55959141808444  sky130_fd_pr__dfl1__example_55959141808444_0
timestamp 1701704242
transform 1 0 1 0 1 1454
box 0 0 1 1
use sky130_fd_pr__nfet_01v8__example_55959141808248  sky130_fd_pr__nfet_01v8__example_55959141808248_0
timestamp 1701704242
transform 1 0 754 0 1 228
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808445  sky130_fd_pr__nfet_01v8__example_55959141808445_0
timestamp 1701704242
transform 1 0 286 0 1 228
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808446  sky130_fd_pr__nfet_01v8__example_55959141808446_0
timestamp 1701704242
transform -1 0 212 0 -1 694
box -19 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808446  sky130_fd_pr__nfet_01v8__example_55959141808446_1
timestamp 1701704242
transform -1 0 212 0 -1 1102
box -19 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808447  sky130_fd_pr__nfet_01v8__example_55959141808447_0
timestamp 1701704242
transform 1 0 442 0 1 228
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808447  sky130_fd_pr__nfet_01v8__example_55959141808447_1
timestamp 1701704242
transform 1 0 598 0 1 228
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808448  sky130_fd_pr__pfet_01v8__example_55959141808448_0
timestamp 1701704242
transform 1 0 72 0 -1 1648
box 120 0 297 1
use sky130_fd_pr__pfet_01v8__example_55959141808450  sky130_fd_pr__pfet_01v8__example_55959141808450_0
timestamp 1701704242
transform -1 0 720 0 -1 1648
box -1 0 297 1
use sky130_fd_pr__pfet_01v8__example_55959141808451  sky130_fd_pr__pfet_01v8__example_55959141808451_0
timestamp 1701704242
transform 1 0 794 0 -1 1648
box -19 0 101 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1701704242
transform 1 0 833 0 1 1618
box 0 0 1 1
<< labels >>
flabel comment s 601 1277 601 1277 0 FreeSans 280 0 0 0 OUT_N
flabel metal1 s 871 1285 899 1313 3 FreeSans 280 180 0 0 OUT
port 1 nsew
flabel metal1 s 227 1732 321 1803 3 FreeSans 520 0 0 0 VPWR
port 2 nsew
flabel metal1 s 55 313 142 434 3 FreeSans 520 0 0 0 VGND
port 3 nsew
flabel locali s 790 109 818 137 3 FreeSans 280 270 0 0 IN1
port 4 nsew
flabel locali s 322 109 350 137 3 FreeSans 280 270 0 0 IN0
port 5 nsew
flabel locali s 482 109 510 137 3 FreeSans 280 270 0 0 IN3
port 6 nsew
flabel locali s 634 109 662 137 3 FreeSans 280 270 0 0 IN2
port 7 nsew
<< properties >>
string GDS_END 64877634
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 64863184
<< end >>
