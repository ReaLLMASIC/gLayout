magic
tech sky130A
magscale 1 2
timestamp 1701704242
use sky130_fd_pr__gendlring__example_559591418081  sky130_fd_pr__gendlring__example_559591418081_0
timestamp 1701704242
transform 1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__genrivetdlring__example_559591418082  sky130_fd_pr__genrivetdlring__example_559591418082_0
timestamp 1701704242
transform 1 0 -478 0 1 -478
box 0 0 1 1
<< properties >>
string GDS_END 9677918
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 9677050
<< end >>
