magic
tech sky130A
magscale 1 2
timestamp 1701704242
use sky130_fd_pr__dfl1__example_55959141808187  sky130_fd_pr__dfl1__example_55959141808187_0
timestamp 1701704242
transform -1 0 8 0 1 21
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808187  sky130_fd_pr__dfl1__example_55959141808187_1
timestamp 1701704242
transform 1 0 9392 0 1 21
box 0 0 1 1
<< properties >>
string GDS_END 58055272
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 58054734
<< end >>
