magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -107 515 811 1337
<< pwell >>
rect -67 367 67 455
rect 285 367 419 455
rect 637 367 771 455
<< mvpsubdiff >>
rect -41 427 41 429
rect -41 393 -17 427
rect 17 393 41 427
rect 311 427 393 429
rect 311 393 335 427
rect 369 393 393 427
rect 663 427 745 429
rect 663 393 687 427
rect 721 393 745 427
<< mvnsubdiff >>
rect -41 583 -17 617
rect 17 583 41 617
rect -41 581 41 583
rect 311 583 335 617
rect 369 583 393 617
rect 311 581 393 583
rect 663 583 687 617
rect 721 583 745 617
rect 663 581 745 583
<< mvpsubdiffcont >>
rect -17 393 17 427
rect 335 393 369 427
rect 687 393 721 427
<< mvnsubdiffcont >>
rect -17 583 17 617
rect 335 583 369 617
rect 687 583 721 617
<< poly >>
rect 21 1353 683 1369
rect 21 1319 37 1353
rect 71 1319 105 1353
rect 139 1319 213 1353
rect 247 1319 281 1353
rect 315 1319 389 1353
rect 423 1319 457 1353
rect 491 1319 565 1353
rect 599 1319 633 1353
rect 667 1319 683 1353
rect 21 1303 683 1319
rect 28 1297 676 1303
rect 52 345 148 645
rect 204 345 300 645
rect 404 345 500 645
rect 556 345 652 645
rect 21 71 683 93
rect 21 37 37 71
rect 71 37 105 71
rect 139 37 213 71
rect 247 37 281 71
rect 315 37 389 71
rect 423 37 457 71
rect 491 37 565 71
rect 599 37 633 71
rect 667 37 683 71
rect 21 21 683 37
<< polycont >>
rect 37 1319 71 1353
rect 105 1319 139 1353
rect 213 1319 247 1353
rect 281 1319 315 1353
rect 389 1319 423 1353
rect 457 1319 491 1353
rect 565 1319 599 1353
rect 633 1319 667 1353
rect 37 37 71 71
rect 105 37 139 71
rect 213 37 247 71
rect 281 37 315 71
rect 389 37 423 71
rect 457 37 491 71
rect 565 37 599 71
rect 633 37 667 71
<< locali >>
rect 37 1353 139 1369
rect 71 1319 105 1353
rect 37 1303 139 1319
rect 213 1353 491 1369
rect 247 1319 281 1353
rect 315 1319 389 1353
rect 423 1319 457 1353
rect 213 1303 491 1319
rect 565 1353 667 1369
rect 599 1319 633 1353
rect 565 1303 667 1319
rect -17 857 17 1209
rect -17 785 17 823
rect -17 713 17 751
rect -17 667 17 679
rect -17 567 17 583
rect -17 427 17 443
rect -17 259 17 297
rect -17 187 17 225
rect -17 121 17 153
rect 51 87 125 1303
rect 159 485 193 1270
rect 159 121 193 451
rect 227 87 301 1303
rect 335 857 369 1209
rect 335 785 369 823
rect 335 713 369 751
rect 335 667 369 679
rect 335 567 369 583
rect 335 427 369 443
rect 335 259 369 297
rect 335 187 369 225
rect 403 87 477 1303
rect 511 485 545 1270
rect 511 121 545 451
rect 579 87 653 1303
rect 687 857 721 1209
rect 687 785 721 823
rect 687 713 721 751
rect 687 667 721 679
rect 687 567 721 583
rect 687 427 721 443
rect 687 259 721 297
rect 687 187 721 225
rect 37 71 139 87
rect 71 37 105 71
rect 37 21 139 37
rect 213 71 491 87
rect 247 37 281 71
rect 315 37 389 71
rect 423 37 457 71
rect 213 21 491 37
rect 565 71 667 87
rect 599 37 633 71
rect 565 21 667 37
<< viali >>
rect -17 823 17 857
rect -17 751 17 785
rect -17 679 17 713
rect -17 617 17 633
rect -17 599 17 617
rect -17 393 17 411
rect -17 377 17 393
rect -17 297 17 331
rect -17 225 17 259
rect -17 153 17 187
rect 159 451 193 485
rect 335 823 369 857
rect 335 751 369 785
rect 335 679 369 713
rect 335 617 369 633
rect 335 599 369 617
rect 335 393 369 411
rect 335 377 369 393
rect 335 297 369 331
rect 335 225 369 259
rect 335 153 369 187
rect 511 451 545 485
rect 687 823 721 857
rect 687 751 721 785
rect 687 679 721 713
rect 687 617 721 633
rect 687 599 721 617
rect 687 393 721 411
rect 687 377 721 393
rect 687 297 721 331
rect 687 225 721 259
rect 687 153 721 187
<< metal1 >>
rect -29 857 733 869
rect -29 823 -17 857
rect 17 823 335 857
rect 369 823 687 857
rect 721 823 733 857
rect -29 785 733 823
rect -29 751 -17 785
rect 17 751 335 785
rect 369 751 687 785
rect 721 751 733 785
rect -29 713 733 751
rect -29 679 -17 713
rect 17 679 335 713
rect 369 679 687 713
rect 721 679 733 713
rect -29 667 733 679
rect -29 633 733 639
rect -29 599 -17 633
rect 17 599 335 633
rect 369 599 687 633
rect 721 599 733 633
rect -29 593 733 599
rect 147 485 557 491
rect 147 451 159 485
rect 193 451 511 485
rect 545 451 557 485
rect 147 445 557 451
rect -29 411 733 417
rect -29 377 -17 411
rect 17 377 335 411
rect 369 377 687 411
rect 721 377 733 411
rect -29 371 733 377
rect -29 331 733 343
rect -29 297 -17 331
rect 17 297 335 331
rect 369 297 687 331
rect 721 297 733 331
rect -29 259 733 297
rect -29 225 -17 259
rect 17 225 335 259
rect 369 225 687 259
rect 721 225 733 259
rect -29 187 733 225
rect -29 153 -17 187
rect 17 153 335 187
rect 369 153 687 187
rect 721 153 733 187
rect -29 141 733 153
use hvnTran_CDNS_52468879185529  hvnTran_CDNS_52468879185529_0
timestamp 1701704242
transform 1 0 28 0 -1 319
box -79 -26 727 226
use hvpTran_CDNS_52468879185530  hvpTran_CDNS_52468879185530_0
timestamp 1701704242
transform 1 0 28 0 1 671
box -119 -66 767 666
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_0
timestamp 1701704242
transform 0 -1 17 -1 0 331
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_1
timestamp 1701704242
transform 0 -1 369 -1 0 331
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_2
timestamp 1701704242
transform 0 -1 721 -1 0 331
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_3
timestamp 1701704242
transform 0 -1 17 1 0 679
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_4
timestamp 1701704242
transform 0 -1 721 1 0 679
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_5
timestamp 1701704242
transform 0 -1 369 1 0 679
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_0
timestamp 1701704242
transform 1 0 687 0 -1 411
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_1
timestamp 1701704242
transform 1 0 -17 0 -1 411
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_2
timestamp 1701704242
transform 1 0 335 0 -1 411
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_3
timestamp 1701704242
transform 1 0 687 0 -1 633
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_4
timestamp 1701704242
transform 1 0 335 0 -1 633
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_5
timestamp 1701704242
transform 1 0 -17 0 -1 633
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_6
timestamp 1701704242
transform 1 0 159 0 1 451
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_7
timestamp 1701704242
transform 1 0 511 0 1 451
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_0
timestamp 1701704242
transform -1 0 155 0 1 21
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_1
timestamp 1701704242
transform -1 0 331 0 1 21
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_2
timestamp 1701704242
transform -1 0 507 0 1 21
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_3
timestamp 1701704242
transform -1 0 683 0 1 21
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_4
timestamp 1701704242
transform -1 0 155 0 1 1303
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_5
timestamp 1701704242
transform -1 0 331 0 1 1303
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_6
timestamp 1701704242
transform -1 0 507 0 1 1303
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_7
timestamp 1701704242
transform -1 0 683 0 1 1303
box 0 0 1 1
<< labels >>
flabel comment s 366 61 366 61 0 FreeSans 100 0 0 0 no_jumper_check
flabel comment s 203 61 203 61 0 FreeSans 100 0 0 0 no_jumper_check
flabel comment s 541 61 541 61 0 FreeSans 100 0 0 0 no_jumper_check
flabel metal1 s 692 667 704 869 3 FreeSans 200 180 0 0 vpwr
port 1 nsew
flabel metal1 s 692 593 704 639 3 FreeSans 200 180 0 0 vpb
port 2 nsew
flabel metal1 s 692 371 704 417 3 FreeSans 200 180 0 0 vnb
port 3 nsew
flabel metal1 s 692 141 704 343 3 FreeSans 200 180 0 0 vgnd
port 4 nsew
flabel metal1 s 0 141 12 343 3 FreeSans 200 0 0 0 vgnd
port 4 nsew
flabel metal1 s 0 371 12 417 3 FreeSans 200 0 0 0 vnb
port 3 nsew
flabel metal1 s 0 593 12 639 3 FreeSans 200 0 0 0 vpb
port 2 nsew
flabel metal1 s 0 667 12 869 3 FreeSans 200 0 0 0 vpwr
port 1 nsew
flabel locali s 71 21 105 71 0 FreeSans 200 0 0 0 in
port 6 nsew
flabel locali s 511 1221 545 1270 0 FreeSans 200 0 0 0 out
port 7 nsew
flabel locali s 159 1221 193 1270 0 FreeSans 200 0 0 0 out
port 7 nsew
flabel locali s 159 121 193 171 0 FreeSans 200 0 0 0 out
port 7 nsew
flabel locali s 511 121 545 171 0 FreeSans 200 0 0 0 out
port 7 nsew
flabel locali s 599 21 633 71 0 FreeSans 200 0 0 0 in
port 6 nsew
flabel locali s 423 21 457 71 0 FreeSans 200 0 0 0 in
port 6 nsew
flabel locali s 246 21 280 71 0 FreeSans 200 0 0 0 in
port 6 nsew
flabel locali s 247 1319 281 1369 0 FreeSans 200 0 0 0 in
port 6 nsew
flabel locali s 71 1319 105 1369 0 FreeSans 200 0 0 0 in
port 6 nsew
flabel locali s 599 1319 633 1369 0 FreeSans 200 0 0 0 in
port 6 nsew
flabel locali s 423 1319 457 1369 0 FreeSans 200 0 0 0 in
port 6 nsew
<< properties >>
string GDS_END 79692690
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 79684828
<< end >>
