magic
tech sky130A
timestamp 1701704242
<< metal1 >>
rect 0 0 3 250
rect 893 0 896 250
<< via1 >>
rect 3 0 893 250
<< metal2 >>
rect 0 0 3 250
rect 893 0 896 250
<< properties >>
string GDS_END 93851234
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 93836766
<< end >>
