magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -38 261 2246 582
<< pwell >>
rect 1220 157 1404 201
rect 1989 157 2179 203
rect 1 145 909 157
rect 1101 145 2179 157
rect 1 21 2179 145
rect 29 -17 63 21
<< locali >>
rect 19 195 89 325
rect 339 153 383 344
rect 422 237 465 274
rect 422 153 513 237
rect 2093 61 2159 484
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2208 561
rect 35 393 69 493
rect 103 427 169 527
rect 35 359 169 393
rect 123 161 169 359
rect 35 127 169 161
rect 35 69 69 127
rect 103 17 169 93
rect 203 69 237 493
rect 271 378 357 493
rect 447 378 513 527
rect 271 103 305 378
rect 551 344 617 485
rect 653 365 692 527
rect 825 404 891 493
rect 983 435 1191 475
rect 825 364 903 404
rect 499 271 617 344
rect 556 235 617 271
rect 761 264 835 330
rect 556 169 727 235
rect 271 51 357 103
rect 447 17 513 103
rect 556 51 601 169
rect 761 137 795 264
rect 869 230 903 364
rect 829 196 903 230
rect 959 225 996 344
rect 1030 331 1123 401
rect 637 17 703 122
rect 829 51 883 196
rect 1030 191 1064 331
rect 1157 315 1191 435
rect 1225 367 1272 527
rect 1157 297 1272 315
rect 963 147 1064 191
rect 1102 263 1272 297
rect 1102 113 1136 263
rect 1238 249 1272 263
rect 1306 275 1372 493
rect 1414 421 1472 527
rect 1585 433 1762 471
rect 1174 213 1214 219
rect 1306 213 1489 275
rect 1558 249 1596 393
rect 1174 209 1489 213
rect 1174 153 1387 209
rect 1630 207 1694 399
rect 1001 51 1136 113
rect 1189 17 1268 112
rect 1306 51 1387 153
rect 1601 141 1694 207
rect 1728 265 1762 433
rect 1796 427 1848 527
rect 1908 381 1976 493
rect 1796 306 1976 381
rect 1728 199 1902 265
rect 1433 17 1488 123
rect 1728 107 1762 199
rect 1938 165 1976 306
rect 2010 293 2059 527
rect 1605 66 1762 107
rect 1810 17 1873 123
rect 1910 60 1976 165
rect 2010 17 2059 180
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2208 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
<< metal1 >>
rect 0 561 2208 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2208 561
rect 0 496 2208 527
rect 0 17 2208 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2208 17
rect 0 -48 2208 -17
<< obsm1 >>
rect 115 388 173 397
rect 1030 388 1088 397
rect 1548 388 1606 397
rect 115 360 1606 388
rect 115 351 173 360
rect 1030 351 1088 360
rect 1548 351 1606 360
rect 191 320 249 329
rect 948 320 1006 329
rect 1632 320 1690 329
rect 191 292 1690 320
rect 191 283 249 292
rect 948 283 1006 292
rect 1632 283 1690 292
rect 749 184 807 193
rect 1928 184 1986 193
rect 749 156 1986 184
rect 749 147 807 156
rect 1928 147 1986 156
rect 259 116 317 125
rect 825 116 883 125
rect 259 79 883 116
<< labels >>
rlabel locali s 19 195 89 325 6 CLK
port 1 nsew clock input
rlabel locali s 339 153 383 344 6 D
port 2 nsew signal input
rlabel locali s 422 153 513 237 6 DE
port 3 nsew signal input
rlabel locali s 422 237 465 274 6 DE
port 3 nsew signal input
rlabel metal1 s 0 -48 2208 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 21 2179 145 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1101 145 2179 157 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 145 909 157 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1989 157 2179 203 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1220 157 1404 201 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 2246 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 2208 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 2093 61 2159 484 6 Q
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 2208 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 3015124
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2997690
<< end >>
