magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -1188 -544 14070 3644
<< pwell >>
rect -1484 3718 14366 3940
rect -1484 -618 -1262 3718
rect 14144 -618 14366 3718
rect -1484 -840 14366 -618
<< mvpmosesd >>
tri -20 3080 0 3100 ne
tri -20 0 0 20 se
rect 0 0 110 3100
tri 110 3080 130 3100 nw
tri 392 3080 412 3100 ne
tri 110 0 130 20 sw
tri 392 0 412 20 se
rect 412 0 522 3100
tri 522 3080 542 3100 nw
tri 804 3080 824 3100 ne
tri 522 0 542 20 sw
tri 804 0 824 20 se
rect 824 0 934 3100
tri 934 3080 954 3100 nw
tri 1216 3080 1236 3100 ne
tri 934 0 954 20 sw
tri 1216 0 1236 20 se
rect 1236 0 1346 3100
tri 1346 3080 1366 3100 nw
tri 1628 3080 1648 3100 ne
tri 1346 0 1366 20 sw
tri 1628 0 1648 20 se
rect 1648 0 1758 3100
tri 1758 3080 1778 3100 nw
tri 2040 3080 2060 3100 ne
tri 1758 0 1778 20 sw
tri 2040 0 2060 20 se
rect 2060 0 2170 3100
tri 2170 3080 2190 3100 nw
tri 2452 3080 2472 3100 ne
tri 2170 0 2190 20 sw
tri 2452 0 2472 20 se
rect 2472 0 2582 3100
tri 2582 3080 2602 3100 nw
tri 2864 3080 2884 3100 ne
tri 2582 0 2602 20 sw
tri 2864 0 2884 20 se
rect 2884 0 2994 3100
tri 2994 3080 3014 3100 nw
tri 3276 3080 3296 3100 ne
tri 2994 0 3014 20 sw
tri 3276 0 3296 20 se
rect 3296 0 3406 3100
tri 3406 3080 3426 3100 nw
tri 3688 3080 3708 3100 ne
tri 3406 0 3426 20 sw
tri 3688 0 3708 20 se
rect 3708 0 3818 3100
tri 3818 3080 3838 3100 nw
tri 4100 3080 4120 3100 ne
tri 3818 0 3838 20 sw
tri 4100 0 4120 20 se
rect 4120 0 4230 3100
tri 4230 3080 4250 3100 nw
tri 4512 3080 4532 3100 ne
tri 4230 0 4250 20 sw
tri 4512 0 4532 20 se
rect 4532 0 4642 3100
tri 4642 3080 4662 3100 nw
tri 4924 3080 4944 3100 ne
tri 4642 0 4662 20 sw
tri 4924 0 4944 20 se
rect 4944 0 5054 3100
tri 5054 3080 5074 3100 nw
tri 5336 3080 5356 3100 ne
tri 5054 0 5074 20 sw
tri 5336 0 5356 20 se
rect 5356 0 5466 3100
tri 5466 3080 5486 3100 nw
tri 5748 3080 5768 3100 ne
tri 5466 0 5486 20 sw
tri 5748 0 5768 20 se
rect 5768 0 5878 3100
tri 5878 3080 5898 3100 nw
tri 6160 3080 6180 3100 ne
tri 5878 0 5898 20 sw
tri 6160 0 6180 20 se
rect 6180 0 6290 3100
tri 6290 3080 6310 3100 nw
tri 6572 3080 6592 3100 ne
tri 6290 0 6310 20 sw
tri 6572 0 6592 20 se
rect 6592 0 6702 3100
tri 6702 3080 6722 3100 nw
tri 6984 3080 7004 3100 ne
tri 6702 0 6722 20 sw
tri 6984 0 7004 20 se
rect 7004 0 7114 3100
tri 7114 3080 7134 3100 nw
tri 7396 3080 7416 3100 ne
tri 7114 0 7134 20 sw
tri 7396 0 7416 20 se
rect 7416 0 7526 3100
tri 7526 3080 7546 3100 nw
tri 7808 3080 7828 3100 ne
tri 7526 0 7546 20 sw
tri 7808 0 7828 20 se
rect 7828 0 7938 3100
tri 7938 3080 7958 3100 nw
tri 8220 3080 8240 3100 ne
tri 7938 0 7958 20 sw
tri 8220 0 8240 20 se
rect 8240 0 8350 3100
tri 8350 3080 8370 3100 nw
tri 8632 3080 8652 3100 ne
tri 8350 0 8370 20 sw
tri 8632 0 8652 20 se
rect 8652 0 8762 3100
tri 8762 3080 8782 3100 nw
tri 9044 3080 9064 3100 ne
tri 8762 0 8782 20 sw
tri 9044 0 9064 20 se
rect 9064 0 9174 3100
tri 9174 3080 9194 3100 nw
tri 9456 3080 9476 3100 ne
tri 9174 0 9194 20 sw
tri 9456 0 9476 20 se
rect 9476 0 9586 3100
tri 9586 3080 9606 3100 nw
tri 9868 3080 9888 3100 ne
tri 9586 0 9606 20 sw
tri 9868 0 9888 20 se
rect 9888 0 9998 3100
tri 9998 3080 10018 3100 nw
tri 10280 3080 10300 3100 ne
tri 9998 0 10018 20 sw
tri 10280 0 10300 20 se
rect 10300 0 10410 3100
tri 10410 3080 10430 3100 nw
tri 10692 3080 10712 3100 ne
tri 10410 0 10430 20 sw
tri 10692 0 10712 20 se
rect 10712 0 10822 3100
tri 10822 3080 10842 3100 nw
tri 11104 3080 11124 3100 ne
tri 10822 0 10842 20 sw
tri 11104 0 11124 20 se
rect 11124 0 11234 3100
tri 11234 3080 11254 3100 nw
tri 11516 3080 11536 3100 ne
tri 11234 0 11254 20 sw
tri 11516 0 11536 20 se
rect 11536 0 11646 3100
tri 11646 3080 11666 3100 nw
tri 11928 3080 11948 3100 ne
tri 11646 0 11666 20 sw
tri 11928 0 11948 20 se
rect 11948 0 12058 3100
tri 12058 3080 12078 3100 nw
tri 12340 3080 12360 3100 ne
tri 12058 0 12078 20 sw
tri 12340 0 12360 20 se
rect 12360 0 12470 3100
tri 12470 3080 12490 3100 nw
tri 12752 3080 12772 3100 ne
tri 12470 0 12490 20 sw
tri 12752 0 12772 20 se
rect 12772 0 12882 3100
tri 12882 3080 12902 3100 nw
tri 12882 0 12902 20 sw
<< mvpdiff >>
rect -232 3080 -20 3100
tri -20 3080 0 3100 sw
rect -232 3000 0 3080
rect -232 790 -202 3000
rect -100 790 0 3000
rect -232 755 0 790
rect -232 721 -202 755
rect -168 721 -134 755
rect -100 721 0 755
rect -232 686 0 721
rect -232 652 -202 686
rect -168 652 -134 686
rect -100 652 0 686
rect -232 617 0 652
rect -232 583 -202 617
rect -168 583 -134 617
rect -100 583 0 617
rect -232 548 0 583
rect -232 514 -202 548
rect -168 514 -134 548
rect -100 514 0 548
rect -232 479 0 514
rect -232 445 -202 479
rect -168 445 -134 479
rect -100 445 0 479
rect -232 410 0 445
rect -232 376 -202 410
rect -168 376 -134 410
rect -100 376 0 410
rect -232 341 0 376
rect -232 307 -202 341
rect -168 307 -134 341
rect -100 307 0 341
rect -232 272 0 307
rect -232 238 -202 272
rect -168 238 -134 272
rect -100 238 0 272
rect -232 203 0 238
rect -232 169 -202 203
rect -168 169 -134 203
rect -100 169 0 203
rect -232 134 0 169
rect -232 100 -202 134
rect -168 100 -134 134
rect -100 100 0 134
rect -232 20 0 100
rect -232 0 -20 20
tri -20 0 0 20 nw
tri 110 3080 130 3100 se
rect 130 3080 392 3100
tri 392 3080 412 3100 sw
rect 110 3000 412 3080
rect 110 790 210 3000
rect 312 790 412 3000
rect 110 755 412 790
rect 110 721 210 755
rect 244 721 278 755
rect 312 721 412 755
rect 110 686 412 721
rect 110 652 210 686
rect 244 652 278 686
rect 312 652 412 686
rect 110 617 412 652
rect 110 583 210 617
rect 244 583 278 617
rect 312 583 412 617
rect 110 548 412 583
rect 110 514 210 548
rect 244 514 278 548
rect 312 514 412 548
rect 110 479 412 514
rect 110 445 210 479
rect 244 445 278 479
rect 312 445 412 479
rect 110 410 412 445
rect 110 376 210 410
rect 244 376 278 410
rect 312 376 412 410
rect 110 341 412 376
rect 110 307 210 341
rect 244 307 278 341
rect 312 307 412 341
rect 110 272 412 307
rect 110 238 210 272
rect 244 238 278 272
rect 312 238 412 272
rect 110 203 412 238
rect 110 169 210 203
rect 244 169 278 203
rect 312 169 412 203
rect 110 134 412 169
rect 110 100 210 134
rect 244 100 278 134
rect 312 100 412 134
rect 110 20 412 100
tri 110 0 130 20 ne
rect 130 0 392 20
tri 392 0 412 20 nw
tri 522 3080 542 3100 se
rect 542 3080 804 3100
tri 804 3080 824 3100 sw
rect 522 3000 824 3080
rect 522 790 622 3000
rect 724 790 824 3000
rect 522 755 824 790
rect 522 721 622 755
rect 656 721 690 755
rect 724 721 824 755
rect 522 686 824 721
rect 522 652 622 686
rect 656 652 690 686
rect 724 652 824 686
rect 522 617 824 652
rect 522 583 622 617
rect 656 583 690 617
rect 724 583 824 617
rect 522 548 824 583
rect 522 514 622 548
rect 656 514 690 548
rect 724 514 824 548
rect 522 479 824 514
rect 522 445 622 479
rect 656 445 690 479
rect 724 445 824 479
rect 522 410 824 445
rect 522 376 622 410
rect 656 376 690 410
rect 724 376 824 410
rect 522 341 824 376
rect 522 307 622 341
rect 656 307 690 341
rect 724 307 824 341
rect 522 272 824 307
rect 522 238 622 272
rect 656 238 690 272
rect 724 238 824 272
rect 522 203 824 238
rect 522 169 622 203
rect 656 169 690 203
rect 724 169 824 203
rect 522 134 824 169
rect 522 100 622 134
rect 656 100 690 134
rect 724 100 824 134
rect 522 20 824 100
tri 522 0 542 20 ne
rect 542 0 804 20
tri 804 0 824 20 nw
tri 934 3080 954 3100 se
rect 954 3080 1216 3100
tri 1216 3080 1236 3100 sw
rect 934 3000 1236 3080
rect 934 790 1034 3000
rect 1136 790 1236 3000
rect 934 755 1236 790
rect 934 721 1034 755
rect 1068 721 1102 755
rect 1136 721 1236 755
rect 934 686 1236 721
rect 934 652 1034 686
rect 1068 652 1102 686
rect 1136 652 1236 686
rect 934 617 1236 652
rect 934 583 1034 617
rect 1068 583 1102 617
rect 1136 583 1236 617
rect 934 548 1236 583
rect 934 514 1034 548
rect 1068 514 1102 548
rect 1136 514 1236 548
rect 934 479 1236 514
rect 934 445 1034 479
rect 1068 445 1102 479
rect 1136 445 1236 479
rect 934 410 1236 445
rect 934 376 1034 410
rect 1068 376 1102 410
rect 1136 376 1236 410
rect 934 341 1236 376
rect 934 307 1034 341
rect 1068 307 1102 341
rect 1136 307 1236 341
rect 934 272 1236 307
rect 934 238 1034 272
rect 1068 238 1102 272
rect 1136 238 1236 272
rect 934 203 1236 238
rect 934 169 1034 203
rect 1068 169 1102 203
rect 1136 169 1236 203
rect 934 134 1236 169
rect 934 100 1034 134
rect 1068 100 1102 134
rect 1136 100 1236 134
rect 934 20 1236 100
tri 934 0 954 20 ne
rect 954 0 1216 20
tri 1216 0 1236 20 nw
tri 1346 3080 1366 3100 se
rect 1366 3080 1628 3100
tri 1628 3080 1648 3100 sw
rect 1346 3000 1648 3080
rect 1346 790 1446 3000
rect 1548 790 1648 3000
rect 1346 755 1648 790
rect 1346 721 1446 755
rect 1480 721 1514 755
rect 1548 721 1648 755
rect 1346 686 1648 721
rect 1346 652 1446 686
rect 1480 652 1514 686
rect 1548 652 1648 686
rect 1346 617 1648 652
rect 1346 583 1446 617
rect 1480 583 1514 617
rect 1548 583 1648 617
rect 1346 548 1648 583
rect 1346 514 1446 548
rect 1480 514 1514 548
rect 1548 514 1648 548
rect 1346 479 1648 514
rect 1346 445 1446 479
rect 1480 445 1514 479
rect 1548 445 1648 479
rect 1346 410 1648 445
rect 1346 376 1446 410
rect 1480 376 1514 410
rect 1548 376 1648 410
rect 1346 341 1648 376
rect 1346 307 1446 341
rect 1480 307 1514 341
rect 1548 307 1648 341
rect 1346 272 1648 307
rect 1346 238 1446 272
rect 1480 238 1514 272
rect 1548 238 1648 272
rect 1346 203 1648 238
rect 1346 169 1446 203
rect 1480 169 1514 203
rect 1548 169 1648 203
rect 1346 134 1648 169
rect 1346 100 1446 134
rect 1480 100 1514 134
rect 1548 100 1648 134
rect 1346 20 1648 100
tri 1346 0 1366 20 ne
rect 1366 0 1628 20
tri 1628 0 1648 20 nw
tri 1758 3080 1778 3100 se
rect 1778 3080 2040 3100
tri 2040 3080 2060 3100 sw
rect 1758 3000 2060 3080
rect 1758 790 1858 3000
rect 1960 790 2060 3000
rect 1758 755 2060 790
rect 1758 721 1858 755
rect 1892 721 1926 755
rect 1960 721 2060 755
rect 1758 686 2060 721
rect 1758 652 1858 686
rect 1892 652 1926 686
rect 1960 652 2060 686
rect 1758 617 2060 652
rect 1758 583 1858 617
rect 1892 583 1926 617
rect 1960 583 2060 617
rect 1758 548 2060 583
rect 1758 514 1858 548
rect 1892 514 1926 548
rect 1960 514 2060 548
rect 1758 479 2060 514
rect 1758 445 1858 479
rect 1892 445 1926 479
rect 1960 445 2060 479
rect 1758 410 2060 445
rect 1758 376 1858 410
rect 1892 376 1926 410
rect 1960 376 2060 410
rect 1758 341 2060 376
rect 1758 307 1858 341
rect 1892 307 1926 341
rect 1960 307 2060 341
rect 1758 272 2060 307
rect 1758 238 1858 272
rect 1892 238 1926 272
rect 1960 238 2060 272
rect 1758 203 2060 238
rect 1758 169 1858 203
rect 1892 169 1926 203
rect 1960 169 2060 203
rect 1758 134 2060 169
rect 1758 100 1858 134
rect 1892 100 1926 134
rect 1960 100 2060 134
rect 1758 20 2060 100
tri 1758 0 1778 20 ne
rect 1778 0 2040 20
tri 2040 0 2060 20 nw
tri 2170 3080 2190 3100 se
rect 2190 3080 2452 3100
tri 2452 3080 2472 3100 sw
rect 2170 3000 2472 3080
rect 2170 790 2270 3000
rect 2372 790 2472 3000
rect 2170 755 2472 790
rect 2170 721 2270 755
rect 2304 721 2338 755
rect 2372 721 2472 755
rect 2170 686 2472 721
rect 2170 652 2270 686
rect 2304 652 2338 686
rect 2372 652 2472 686
rect 2170 617 2472 652
rect 2170 583 2270 617
rect 2304 583 2338 617
rect 2372 583 2472 617
rect 2170 548 2472 583
rect 2170 514 2270 548
rect 2304 514 2338 548
rect 2372 514 2472 548
rect 2170 479 2472 514
rect 2170 445 2270 479
rect 2304 445 2338 479
rect 2372 445 2472 479
rect 2170 410 2472 445
rect 2170 376 2270 410
rect 2304 376 2338 410
rect 2372 376 2472 410
rect 2170 341 2472 376
rect 2170 307 2270 341
rect 2304 307 2338 341
rect 2372 307 2472 341
rect 2170 272 2472 307
rect 2170 238 2270 272
rect 2304 238 2338 272
rect 2372 238 2472 272
rect 2170 203 2472 238
rect 2170 169 2270 203
rect 2304 169 2338 203
rect 2372 169 2472 203
rect 2170 134 2472 169
rect 2170 100 2270 134
rect 2304 100 2338 134
rect 2372 100 2472 134
rect 2170 20 2472 100
tri 2170 0 2190 20 ne
rect 2190 0 2452 20
tri 2452 0 2472 20 nw
tri 2582 3080 2602 3100 se
rect 2602 3080 2864 3100
tri 2864 3080 2884 3100 sw
rect 2582 3000 2884 3080
rect 2582 790 2682 3000
rect 2784 790 2884 3000
rect 2582 755 2884 790
rect 2582 721 2682 755
rect 2716 721 2750 755
rect 2784 721 2884 755
rect 2582 686 2884 721
rect 2582 652 2682 686
rect 2716 652 2750 686
rect 2784 652 2884 686
rect 2582 617 2884 652
rect 2582 583 2682 617
rect 2716 583 2750 617
rect 2784 583 2884 617
rect 2582 548 2884 583
rect 2582 514 2682 548
rect 2716 514 2750 548
rect 2784 514 2884 548
rect 2582 479 2884 514
rect 2582 445 2682 479
rect 2716 445 2750 479
rect 2784 445 2884 479
rect 2582 410 2884 445
rect 2582 376 2682 410
rect 2716 376 2750 410
rect 2784 376 2884 410
rect 2582 341 2884 376
rect 2582 307 2682 341
rect 2716 307 2750 341
rect 2784 307 2884 341
rect 2582 272 2884 307
rect 2582 238 2682 272
rect 2716 238 2750 272
rect 2784 238 2884 272
rect 2582 203 2884 238
rect 2582 169 2682 203
rect 2716 169 2750 203
rect 2784 169 2884 203
rect 2582 134 2884 169
rect 2582 100 2682 134
rect 2716 100 2750 134
rect 2784 100 2884 134
rect 2582 20 2884 100
tri 2582 0 2602 20 ne
rect 2602 0 2864 20
tri 2864 0 2884 20 nw
tri 2994 3080 3014 3100 se
rect 3014 3080 3276 3100
tri 3276 3080 3296 3100 sw
rect 2994 3000 3296 3080
rect 2994 790 3094 3000
rect 3196 790 3296 3000
rect 2994 755 3296 790
rect 2994 721 3094 755
rect 3128 721 3162 755
rect 3196 721 3296 755
rect 2994 686 3296 721
rect 2994 652 3094 686
rect 3128 652 3162 686
rect 3196 652 3296 686
rect 2994 617 3296 652
rect 2994 583 3094 617
rect 3128 583 3162 617
rect 3196 583 3296 617
rect 2994 548 3296 583
rect 2994 514 3094 548
rect 3128 514 3162 548
rect 3196 514 3296 548
rect 2994 479 3296 514
rect 2994 445 3094 479
rect 3128 445 3162 479
rect 3196 445 3296 479
rect 2994 410 3296 445
rect 2994 376 3094 410
rect 3128 376 3162 410
rect 3196 376 3296 410
rect 2994 341 3296 376
rect 2994 307 3094 341
rect 3128 307 3162 341
rect 3196 307 3296 341
rect 2994 272 3296 307
rect 2994 238 3094 272
rect 3128 238 3162 272
rect 3196 238 3296 272
rect 2994 203 3296 238
rect 2994 169 3094 203
rect 3128 169 3162 203
rect 3196 169 3296 203
rect 2994 134 3296 169
rect 2994 100 3094 134
rect 3128 100 3162 134
rect 3196 100 3296 134
rect 2994 20 3296 100
tri 2994 0 3014 20 ne
rect 3014 0 3276 20
tri 3276 0 3296 20 nw
tri 3406 3080 3426 3100 se
rect 3426 3080 3688 3100
tri 3688 3080 3708 3100 sw
rect 3406 3000 3708 3080
rect 3406 790 3506 3000
rect 3608 790 3708 3000
rect 3406 755 3708 790
rect 3406 721 3506 755
rect 3540 721 3574 755
rect 3608 721 3708 755
rect 3406 686 3708 721
rect 3406 652 3506 686
rect 3540 652 3574 686
rect 3608 652 3708 686
rect 3406 617 3708 652
rect 3406 583 3506 617
rect 3540 583 3574 617
rect 3608 583 3708 617
rect 3406 548 3708 583
rect 3406 514 3506 548
rect 3540 514 3574 548
rect 3608 514 3708 548
rect 3406 479 3708 514
rect 3406 445 3506 479
rect 3540 445 3574 479
rect 3608 445 3708 479
rect 3406 410 3708 445
rect 3406 376 3506 410
rect 3540 376 3574 410
rect 3608 376 3708 410
rect 3406 341 3708 376
rect 3406 307 3506 341
rect 3540 307 3574 341
rect 3608 307 3708 341
rect 3406 272 3708 307
rect 3406 238 3506 272
rect 3540 238 3574 272
rect 3608 238 3708 272
rect 3406 203 3708 238
rect 3406 169 3506 203
rect 3540 169 3574 203
rect 3608 169 3708 203
rect 3406 134 3708 169
rect 3406 100 3506 134
rect 3540 100 3574 134
rect 3608 100 3708 134
rect 3406 20 3708 100
tri 3406 0 3426 20 ne
rect 3426 0 3688 20
tri 3688 0 3708 20 nw
tri 3818 3080 3838 3100 se
rect 3838 3080 4100 3100
tri 4100 3080 4120 3100 sw
rect 3818 3000 4120 3080
rect 3818 790 3918 3000
rect 4020 790 4120 3000
rect 3818 755 4120 790
rect 3818 721 3918 755
rect 3952 721 3986 755
rect 4020 721 4120 755
rect 3818 686 4120 721
rect 3818 652 3918 686
rect 3952 652 3986 686
rect 4020 652 4120 686
rect 3818 617 4120 652
rect 3818 583 3918 617
rect 3952 583 3986 617
rect 4020 583 4120 617
rect 3818 548 4120 583
rect 3818 514 3918 548
rect 3952 514 3986 548
rect 4020 514 4120 548
rect 3818 479 4120 514
rect 3818 445 3918 479
rect 3952 445 3986 479
rect 4020 445 4120 479
rect 3818 410 4120 445
rect 3818 376 3918 410
rect 3952 376 3986 410
rect 4020 376 4120 410
rect 3818 341 4120 376
rect 3818 307 3918 341
rect 3952 307 3986 341
rect 4020 307 4120 341
rect 3818 272 4120 307
rect 3818 238 3918 272
rect 3952 238 3986 272
rect 4020 238 4120 272
rect 3818 203 4120 238
rect 3818 169 3918 203
rect 3952 169 3986 203
rect 4020 169 4120 203
rect 3818 134 4120 169
rect 3818 100 3918 134
rect 3952 100 3986 134
rect 4020 100 4120 134
rect 3818 20 4120 100
tri 3818 0 3838 20 ne
rect 3838 0 4100 20
tri 4100 0 4120 20 nw
tri 4230 3080 4250 3100 se
rect 4250 3080 4512 3100
tri 4512 3080 4532 3100 sw
rect 4230 3000 4532 3080
rect 4230 790 4330 3000
rect 4432 790 4532 3000
rect 4230 755 4532 790
rect 4230 721 4330 755
rect 4364 721 4398 755
rect 4432 721 4532 755
rect 4230 686 4532 721
rect 4230 652 4330 686
rect 4364 652 4398 686
rect 4432 652 4532 686
rect 4230 617 4532 652
rect 4230 583 4330 617
rect 4364 583 4398 617
rect 4432 583 4532 617
rect 4230 548 4532 583
rect 4230 514 4330 548
rect 4364 514 4398 548
rect 4432 514 4532 548
rect 4230 479 4532 514
rect 4230 445 4330 479
rect 4364 445 4398 479
rect 4432 445 4532 479
rect 4230 410 4532 445
rect 4230 376 4330 410
rect 4364 376 4398 410
rect 4432 376 4532 410
rect 4230 341 4532 376
rect 4230 307 4330 341
rect 4364 307 4398 341
rect 4432 307 4532 341
rect 4230 272 4532 307
rect 4230 238 4330 272
rect 4364 238 4398 272
rect 4432 238 4532 272
rect 4230 203 4532 238
rect 4230 169 4330 203
rect 4364 169 4398 203
rect 4432 169 4532 203
rect 4230 134 4532 169
rect 4230 100 4330 134
rect 4364 100 4398 134
rect 4432 100 4532 134
rect 4230 20 4532 100
tri 4230 0 4250 20 ne
rect 4250 0 4512 20
tri 4512 0 4532 20 nw
tri 4642 3080 4662 3100 se
rect 4662 3080 4924 3100
tri 4924 3080 4944 3100 sw
rect 4642 3000 4944 3080
rect 4642 790 4742 3000
rect 4844 790 4944 3000
rect 4642 755 4944 790
rect 4642 721 4742 755
rect 4776 721 4810 755
rect 4844 721 4944 755
rect 4642 686 4944 721
rect 4642 652 4742 686
rect 4776 652 4810 686
rect 4844 652 4944 686
rect 4642 617 4944 652
rect 4642 583 4742 617
rect 4776 583 4810 617
rect 4844 583 4944 617
rect 4642 548 4944 583
rect 4642 514 4742 548
rect 4776 514 4810 548
rect 4844 514 4944 548
rect 4642 479 4944 514
rect 4642 445 4742 479
rect 4776 445 4810 479
rect 4844 445 4944 479
rect 4642 410 4944 445
rect 4642 376 4742 410
rect 4776 376 4810 410
rect 4844 376 4944 410
rect 4642 341 4944 376
rect 4642 307 4742 341
rect 4776 307 4810 341
rect 4844 307 4944 341
rect 4642 272 4944 307
rect 4642 238 4742 272
rect 4776 238 4810 272
rect 4844 238 4944 272
rect 4642 203 4944 238
rect 4642 169 4742 203
rect 4776 169 4810 203
rect 4844 169 4944 203
rect 4642 134 4944 169
rect 4642 100 4742 134
rect 4776 100 4810 134
rect 4844 100 4944 134
rect 4642 20 4944 100
tri 4642 0 4662 20 ne
rect 4662 0 4924 20
tri 4924 0 4944 20 nw
tri 5054 3080 5074 3100 se
rect 5074 3080 5336 3100
tri 5336 3080 5356 3100 sw
rect 5054 3000 5356 3080
rect 5054 790 5154 3000
rect 5256 790 5356 3000
rect 5054 755 5356 790
rect 5054 721 5154 755
rect 5188 721 5222 755
rect 5256 721 5356 755
rect 5054 686 5356 721
rect 5054 652 5154 686
rect 5188 652 5222 686
rect 5256 652 5356 686
rect 5054 617 5356 652
rect 5054 583 5154 617
rect 5188 583 5222 617
rect 5256 583 5356 617
rect 5054 548 5356 583
rect 5054 514 5154 548
rect 5188 514 5222 548
rect 5256 514 5356 548
rect 5054 479 5356 514
rect 5054 445 5154 479
rect 5188 445 5222 479
rect 5256 445 5356 479
rect 5054 410 5356 445
rect 5054 376 5154 410
rect 5188 376 5222 410
rect 5256 376 5356 410
rect 5054 341 5356 376
rect 5054 307 5154 341
rect 5188 307 5222 341
rect 5256 307 5356 341
rect 5054 272 5356 307
rect 5054 238 5154 272
rect 5188 238 5222 272
rect 5256 238 5356 272
rect 5054 203 5356 238
rect 5054 169 5154 203
rect 5188 169 5222 203
rect 5256 169 5356 203
rect 5054 134 5356 169
rect 5054 100 5154 134
rect 5188 100 5222 134
rect 5256 100 5356 134
rect 5054 20 5356 100
tri 5054 0 5074 20 ne
rect 5074 0 5336 20
tri 5336 0 5356 20 nw
tri 5466 3080 5486 3100 se
rect 5486 3080 5748 3100
tri 5748 3080 5768 3100 sw
rect 5466 3000 5768 3080
rect 5466 790 5566 3000
rect 5668 790 5768 3000
rect 5466 755 5768 790
rect 5466 721 5566 755
rect 5600 721 5634 755
rect 5668 721 5768 755
rect 5466 686 5768 721
rect 5466 652 5566 686
rect 5600 652 5634 686
rect 5668 652 5768 686
rect 5466 617 5768 652
rect 5466 583 5566 617
rect 5600 583 5634 617
rect 5668 583 5768 617
rect 5466 548 5768 583
rect 5466 514 5566 548
rect 5600 514 5634 548
rect 5668 514 5768 548
rect 5466 479 5768 514
rect 5466 445 5566 479
rect 5600 445 5634 479
rect 5668 445 5768 479
rect 5466 410 5768 445
rect 5466 376 5566 410
rect 5600 376 5634 410
rect 5668 376 5768 410
rect 5466 341 5768 376
rect 5466 307 5566 341
rect 5600 307 5634 341
rect 5668 307 5768 341
rect 5466 272 5768 307
rect 5466 238 5566 272
rect 5600 238 5634 272
rect 5668 238 5768 272
rect 5466 203 5768 238
rect 5466 169 5566 203
rect 5600 169 5634 203
rect 5668 169 5768 203
rect 5466 134 5768 169
rect 5466 100 5566 134
rect 5600 100 5634 134
rect 5668 100 5768 134
rect 5466 20 5768 100
tri 5466 0 5486 20 ne
rect 5486 0 5748 20
tri 5748 0 5768 20 nw
tri 5878 3080 5898 3100 se
rect 5898 3080 6160 3100
tri 6160 3080 6180 3100 sw
rect 5878 3000 6180 3080
rect 5878 790 5978 3000
rect 6080 790 6180 3000
rect 5878 755 6180 790
rect 5878 721 5978 755
rect 6012 721 6046 755
rect 6080 721 6180 755
rect 5878 686 6180 721
rect 5878 652 5978 686
rect 6012 652 6046 686
rect 6080 652 6180 686
rect 5878 617 6180 652
rect 5878 583 5978 617
rect 6012 583 6046 617
rect 6080 583 6180 617
rect 5878 548 6180 583
rect 5878 514 5978 548
rect 6012 514 6046 548
rect 6080 514 6180 548
rect 5878 479 6180 514
rect 5878 445 5978 479
rect 6012 445 6046 479
rect 6080 445 6180 479
rect 5878 410 6180 445
rect 5878 376 5978 410
rect 6012 376 6046 410
rect 6080 376 6180 410
rect 5878 341 6180 376
rect 5878 307 5978 341
rect 6012 307 6046 341
rect 6080 307 6180 341
rect 5878 272 6180 307
rect 5878 238 5978 272
rect 6012 238 6046 272
rect 6080 238 6180 272
rect 5878 203 6180 238
rect 5878 169 5978 203
rect 6012 169 6046 203
rect 6080 169 6180 203
rect 5878 134 6180 169
rect 5878 100 5978 134
rect 6012 100 6046 134
rect 6080 100 6180 134
rect 5878 20 6180 100
tri 5878 0 5898 20 ne
rect 5898 0 6160 20
tri 6160 0 6180 20 nw
tri 6290 3080 6310 3100 se
rect 6310 3080 6572 3100
tri 6572 3080 6592 3100 sw
rect 6290 3000 6592 3080
rect 6290 790 6390 3000
rect 6492 790 6592 3000
rect 6290 755 6592 790
rect 6290 721 6390 755
rect 6424 721 6458 755
rect 6492 721 6592 755
rect 6290 686 6592 721
rect 6290 652 6390 686
rect 6424 652 6458 686
rect 6492 652 6592 686
rect 6290 617 6592 652
rect 6290 583 6390 617
rect 6424 583 6458 617
rect 6492 583 6592 617
rect 6290 548 6592 583
rect 6290 514 6390 548
rect 6424 514 6458 548
rect 6492 514 6592 548
rect 6290 479 6592 514
rect 6290 445 6390 479
rect 6424 445 6458 479
rect 6492 445 6592 479
rect 6290 410 6592 445
rect 6290 376 6390 410
rect 6424 376 6458 410
rect 6492 376 6592 410
rect 6290 341 6592 376
rect 6290 307 6390 341
rect 6424 307 6458 341
rect 6492 307 6592 341
rect 6290 272 6592 307
rect 6290 238 6390 272
rect 6424 238 6458 272
rect 6492 238 6592 272
rect 6290 203 6592 238
rect 6290 169 6390 203
rect 6424 169 6458 203
rect 6492 169 6592 203
rect 6290 134 6592 169
rect 6290 100 6390 134
rect 6424 100 6458 134
rect 6492 100 6592 134
rect 6290 20 6592 100
tri 6290 0 6310 20 ne
rect 6310 0 6572 20
tri 6572 0 6592 20 nw
tri 6702 3080 6722 3100 se
rect 6722 3080 6984 3100
tri 6984 3080 7004 3100 sw
rect 6702 3000 7004 3080
rect 6702 790 6802 3000
rect 6904 790 7004 3000
rect 6702 755 7004 790
rect 6702 721 6802 755
rect 6836 721 6870 755
rect 6904 721 7004 755
rect 6702 686 7004 721
rect 6702 652 6802 686
rect 6836 652 6870 686
rect 6904 652 7004 686
rect 6702 617 7004 652
rect 6702 583 6802 617
rect 6836 583 6870 617
rect 6904 583 7004 617
rect 6702 548 7004 583
rect 6702 514 6802 548
rect 6836 514 6870 548
rect 6904 514 7004 548
rect 6702 479 7004 514
rect 6702 445 6802 479
rect 6836 445 6870 479
rect 6904 445 7004 479
rect 6702 410 7004 445
rect 6702 376 6802 410
rect 6836 376 6870 410
rect 6904 376 7004 410
rect 6702 341 7004 376
rect 6702 307 6802 341
rect 6836 307 6870 341
rect 6904 307 7004 341
rect 6702 272 7004 307
rect 6702 238 6802 272
rect 6836 238 6870 272
rect 6904 238 7004 272
rect 6702 203 7004 238
rect 6702 169 6802 203
rect 6836 169 6870 203
rect 6904 169 7004 203
rect 6702 134 7004 169
rect 6702 100 6802 134
rect 6836 100 6870 134
rect 6904 100 7004 134
rect 6702 20 7004 100
tri 6702 0 6722 20 ne
rect 6722 0 6984 20
tri 6984 0 7004 20 nw
tri 7114 3080 7134 3100 se
rect 7134 3080 7396 3100
tri 7396 3080 7416 3100 sw
rect 7114 3000 7416 3080
rect 7114 790 7214 3000
rect 7316 790 7416 3000
rect 7114 755 7416 790
rect 7114 721 7214 755
rect 7248 721 7282 755
rect 7316 721 7416 755
rect 7114 686 7416 721
rect 7114 652 7214 686
rect 7248 652 7282 686
rect 7316 652 7416 686
rect 7114 617 7416 652
rect 7114 583 7214 617
rect 7248 583 7282 617
rect 7316 583 7416 617
rect 7114 548 7416 583
rect 7114 514 7214 548
rect 7248 514 7282 548
rect 7316 514 7416 548
rect 7114 479 7416 514
rect 7114 445 7214 479
rect 7248 445 7282 479
rect 7316 445 7416 479
rect 7114 410 7416 445
rect 7114 376 7214 410
rect 7248 376 7282 410
rect 7316 376 7416 410
rect 7114 341 7416 376
rect 7114 307 7214 341
rect 7248 307 7282 341
rect 7316 307 7416 341
rect 7114 272 7416 307
rect 7114 238 7214 272
rect 7248 238 7282 272
rect 7316 238 7416 272
rect 7114 203 7416 238
rect 7114 169 7214 203
rect 7248 169 7282 203
rect 7316 169 7416 203
rect 7114 134 7416 169
rect 7114 100 7214 134
rect 7248 100 7282 134
rect 7316 100 7416 134
rect 7114 20 7416 100
tri 7114 0 7134 20 ne
rect 7134 0 7396 20
tri 7396 0 7416 20 nw
tri 7526 3080 7546 3100 se
rect 7546 3080 7808 3100
tri 7808 3080 7828 3100 sw
rect 7526 3000 7828 3080
rect 7526 790 7626 3000
rect 7728 790 7828 3000
rect 7526 755 7828 790
rect 7526 721 7626 755
rect 7660 721 7694 755
rect 7728 721 7828 755
rect 7526 686 7828 721
rect 7526 652 7626 686
rect 7660 652 7694 686
rect 7728 652 7828 686
rect 7526 617 7828 652
rect 7526 583 7626 617
rect 7660 583 7694 617
rect 7728 583 7828 617
rect 7526 548 7828 583
rect 7526 514 7626 548
rect 7660 514 7694 548
rect 7728 514 7828 548
rect 7526 479 7828 514
rect 7526 445 7626 479
rect 7660 445 7694 479
rect 7728 445 7828 479
rect 7526 410 7828 445
rect 7526 376 7626 410
rect 7660 376 7694 410
rect 7728 376 7828 410
rect 7526 341 7828 376
rect 7526 307 7626 341
rect 7660 307 7694 341
rect 7728 307 7828 341
rect 7526 272 7828 307
rect 7526 238 7626 272
rect 7660 238 7694 272
rect 7728 238 7828 272
rect 7526 203 7828 238
rect 7526 169 7626 203
rect 7660 169 7694 203
rect 7728 169 7828 203
rect 7526 134 7828 169
rect 7526 100 7626 134
rect 7660 100 7694 134
rect 7728 100 7828 134
rect 7526 20 7828 100
tri 7526 0 7546 20 ne
rect 7546 0 7808 20
tri 7808 0 7828 20 nw
tri 7938 3080 7958 3100 se
rect 7958 3080 8220 3100
tri 8220 3080 8240 3100 sw
rect 7938 3000 8240 3080
rect 7938 790 8038 3000
rect 8140 790 8240 3000
rect 7938 755 8240 790
rect 7938 721 8038 755
rect 8072 721 8106 755
rect 8140 721 8240 755
rect 7938 686 8240 721
rect 7938 652 8038 686
rect 8072 652 8106 686
rect 8140 652 8240 686
rect 7938 617 8240 652
rect 7938 583 8038 617
rect 8072 583 8106 617
rect 8140 583 8240 617
rect 7938 548 8240 583
rect 7938 514 8038 548
rect 8072 514 8106 548
rect 8140 514 8240 548
rect 7938 479 8240 514
rect 7938 445 8038 479
rect 8072 445 8106 479
rect 8140 445 8240 479
rect 7938 410 8240 445
rect 7938 376 8038 410
rect 8072 376 8106 410
rect 8140 376 8240 410
rect 7938 341 8240 376
rect 7938 307 8038 341
rect 8072 307 8106 341
rect 8140 307 8240 341
rect 7938 272 8240 307
rect 7938 238 8038 272
rect 8072 238 8106 272
rect 8140 238 8240 272
rect 7938 203 8240 238
rect 7938 169 8038 203
rect 8072 169 8106 203
rect 8140 169 8240 203
rect 7938 134 8240 169
rect 7938 100 8038 134
rect 8072 100 8106 134
rect 8140 100 8240 134
rect 7938 20 8240 100
tri 7938 0 7958 20 ne
rect 7958 0 8220 20
tri 8220 0 8240 20 nw
tri 8350 3080 8370 3100 se
rect 8370 3080 8632 3100
tri 8632 3080 8652 3100 sw
rect 8350 3000 8652 3080
rect 8350 790 8450 3000
rect 8552 790 8652 3000
rect 8350 755 8652 790
rect 8350 721 8450 755
rect 8484 721 8518 755
rect 8552 721 8652 755
rect 8350 686 8652 721
rect 8350 652 8450 686
rect 8484 652 8518 686
rect 8552 652 8652 686
rect 8350 617 8652 652
rect 8350 583 8450 617
rect 8484 583 8518 617
rect 8552 583 8652 617
rect 8350 548 8652 583
rect 8350 514 8450 548
rect 8484 514 8518 548
rect 8552 514 8652 548
rect 8350 479 8652 514
rect 8350 445 8450 479
rect 8484 445 8518 479
rect 8552 445 8652 479
rect 8350 410 8652 445
rect 8350 376 8450 410
rect 8484 376 8518 410
rect 8552 376 8652 410
rect 8350 341 8652 376
rect 8350 307 8450 341
rect 8484 307 8518 341
rect 8552 307 8652 341
rect 8350 272 8652 307
rect 8350 238 8450 272
rect 8484 238 8518 272
rect 8552 238 8652 272
rect 8350 203 8652 238
rect 8350 169 8450 203
rect 8484 169 8518 203
rect 8552 169 8652 203
rect 8350 134 8652 169
rect 8350 100 8450 134
rect 8484 100 8518 134
rect 8552 100 8652 134
rect 8350 20 8652 100
tri 8350 0 8370 20 ne
rect 8370 0 8632 20
tri 8632 0 8652 20 nw
tri 8762 3080 8782 3100 se
rect 8782 3080 9044 3100
tri 9044 3080 9064 3100 sw
rect 8762 3000 9064 3080
rect 8762 790 8862 3000
rect 8964 790 9064 3000
rect 8762 755 9064 790
rect 8762 721 8862 755
rect 8896 721 8930 755
rect 8964 721 9064 755
rect 8762 686 9064 721
rect 8762 652 8862 686
rect 8896 652 8930 686
rect 8964 652 9064 686
rect 8762 617 9064 652
rect 8762 583 8862 617
rect 8896 583 8930 617
rect 8964 583 9064 617
rect 8762 548 9064 583
rect 8762 514 8862 548
rect 8896 514 8930 548
rect 8964 514 9064 548
rect 8762 479 9064 514
rect 8762 445 8862 479
rect 8896 445 8930 479
rect 8964 445 9064 479
rect 8762 410 9064 445
rect 8762 376 8862 410
rect 8896 376 8930 410
rect 8964 376 9064 410
rect 8762 341 9064 376
rect 8762 307 8862 341
rect 8896 307 8930 341
rect 8964 307 9064 341
rect 8762 272 9064 307
rect 8762 238 8862 272
rect 8896 238 8930 272
rect 8964 238 9064 272
rect 8762 203 9064 238
rect 8762 169 8862 203
rect 8896 169 8930 203
rect 8964 169 9064 203
rect 8762 134 9064 169
rect 8762 100 8862 134
rect 8896 100 8930 134
rect 8964 100 9064 134
rect 8762 20 9064 100
tri 8762 0 8782 20 ne
rect 8782 0 9044 20
tri 9044 0 9064 20 nw
tri 9174 3080 9194 3100 se
rect 9194 3080 9456 3100
tri 9456 3080 9476 3100 sw
rect 9174 3000 9476 3080
rect 9174 790 9274 3000
rect 9376 790 9476 3000
rect 9174 755 9476 790
rect 9174 721 9274 755
rect 9308 721 9342 755
rect 9376 721 9476 755
rect 9174 686 9476 721
rect 9174 652 9274 686
rect 9308 652 9342 686
rect 9376 652 9476 686
rect 9174 617 9476 652
rect 9174 583 9274 617
rect 9308 583 9342 617
rect 9376 583 9476 617
rect 9174 548 9476 583
rect 9174 514 9274 548
rect 9308 514 9342 548
rect 9376 514 9476 548
rect 9174 479 9476 514
rect 9174 445 9274 479
rect 9308 445 9342 479
rect 9376 445 9476 479
rect 9174 410 9476 445
rect 9174 376 9274 410
rect 9308 376 9342 410
rect 9376 376 9476 410
rect 9174 341 9476 376
rect 9174 307 9274 341
rect 9308 307 9342 341
rect 9376 307 9476 341
rect 9174 272 9476 307
rect 9174 238 9274 272
rect 9308 238 9342 272
rect 9376 238 9476 272
rect 9174 203 9476 238
rect 9174 169 9274 203
rect 9308 169 9342 203
rect 9376 169 9476 203
rect 9174 134 9476 169
rect 9174 100 9274 134
rect 9308 100 9342 134
rect 9376 100 9476 134
rect 9174 20 9476 100
tri 9174 0 9194 20 ne
rect 9194 0 9456 20
tri 9456 0 9476 20 nw
tri 9586 3080 9606 3100 se
rect 9606 3080 9868 3100
tri 9868 3080 9888 3100 sw
rect 9586 3000 9888 3080
rect 9586 790 9686 3000
rect 9788 790 9888 3000
rect 9586 755 9888 790
rect 9586 721 9686 755
rect 9720 721 9754 755
rect 9788 721 9888 755
rect 9586 686 9888 721
rect 9586 652 9686 686
rect 9720 652 9754 686
rect 9788 652 9888 686
rect 9586 617 9888 652
rect 9586 583 9686 617
rect 9720 583 9754 617
rect 9788 583 9888 617
rect 9586 548 9888 583
rect 9586 514 9686 548
rect 9720 514 9754 548
rect 9788 514 9888 548
rect 9586 479 9888 514
rect 9586 445 9686 479
rect 9720 445 9754 479
rect 9788 445 9888 479
rect 9586 410 9888 445
rect 9586 376 9686 410
rect 9720 376 9754 410
rect 9788 376 9888 410
rect 9586 341 9888 376
rect 9586 307 9686 341
rect 9720 307 9754 341
rect 9788 307 9888 341
rect 9586 272 9888 307
rect 9586 238 9686 272
rect 9720 238 9754 272
rect 9788 238 9888 272
rect 9586 203 9888 238
rect 9586 169 9686 203
rect 9720 169 9754 203
rect 9788 169 9888 203
rect 9586 134 9888 169
rect 9586 100 9686 134
rect 9720 100 9754 134
rect 9788 100 9888 134
rect 9586 20 9888 100
tri 9586 0 9606 20 ne
rect 9606 0 9868 20
tri 9868 0 9888 20 nw
tri 9998 3080 10018 3100 se
rect 10018 3080 10280 3100
tri 10280 3080 10300 3100 sw
rect 9998 3000 10300 3080
rect 9998 790 10098 3000
rect 10200 790 10300 3000
rect 9998 755 10300 790
rect 9998 721 10098 755
rect 10132 721 10166 755
rect 10200 721 10300 755
rect 9998 686 10300 721
rect 9998 652 10098 686
rect 10132 652 10166 686
rect 10200 652 10300 686
rect 9998 617 10300 652
rect 9998 583 10098 617
rect 10132 583 10166 617
rect 10200 583 10300 617
rect 9998 548 10300 583
rect 9998 514 10098 548
rect 10132 514 10166 548
rect 10200 514 10300 548
rect 9998 479 10300 514
rect 9998 445 10098 479
rect 10132 445 10166 479
rect 10200 445 10300 479
rect 9998 410 10300 445
rect 9998 376 10098 410
rect 10132 376 10166 410
rect 10200 376 10300 410
rect 9998 341 10300 376
rect 9998 307 10098 341
rect 10132 307 10166 341
rect 10200 307 10300 341
rect 9998 272 10300 307
rect 9998 238 10098 272
rect 10132 238 10166 272
rect 10200 238 10300 272
rect 9998 203 10300 238
rect 9998 169 10098 203
rect 10132 169 10166 203
rect 10200 169 10300 203
rect 9998 134 10300 169
rect 9998 100 10098 134
rect 10132 100 10166 134
rect 10200 100 10300 134
rect 9998 20 10300 100
tri 9998 0 10018 20 ne
rect 10018 0 10280 20
tri 10280 0 10300 20 nw
tri 10410 3080 10430 3100 se
rect 10430 3080 10692 3100
tri 10692 3080 10712 3100 sw
rect 10410 3000 10712 3080
rect 10410 790 10510 3000
rect 10612 790 10712 3000
rect 10410 755 10712 790
rect 10410 721 10510 755
rect 10544 721 10578 755
rect 10612 721 10712 755
rect 10410 686 10712 721
rect 10410 652 10510 686
rect 10544 652 10578 686
rect 10612 652 10712 686
rect 10410 617 10712 652
rect 10410 583 10510 617
rect 10544 583 10578 617
rect 10612 583 10712 617
rect 10410 548 10712 583
rect 10410 514 10510 548
rect 10544 514 10578 548
rect 10612 514 10712 548
rect 10410 479 10712 514
rect 10410 445 10510 479
rect 10544 445 10578 479
rect 10612 445 10712 479
rect 10410 410 10712 445
rect 10410 376 10510 410
rect 10544 376 10578 410
rect 10612 376 10712 410
rect 10410 341 10712 376
rect 10410 307 10510 341
rect 10544 307 10578 341
rect 10612 307 10712 341
rect 10410 272 10712 307
rect 10410 238 10510 272
rect 10544 238 10578 272
rect 10612 238 10712 272
rect 10410 203 10712 238
rect 10410 169 10510 203
rect 10544 169 10578 203
rect 10612 169 10712 203
rect 10410 134 10712 169
rect 10410 100 10510 134
rect 10544 100 10578 134
rect 10612 100 10712 134
rect 10410 20 10712 100
tri 10410 0 10430 20 ne
rect 10430 0 10692 20
tri 10692 0 10712 20 nw
tri 10822 3080 10842 3100 se
rect 10842 3080 11104 3100
tri 11104 3080 11124 3100 sw
rect 10822 3000 11124 3080
rect 10822 790 10922 3000
rect 11024 790 11124 3000
rect 10822 755 11124 790
rect 10822 721 10922 755
rect 10956 721 10990 755
rect 11024 721 11124 755
rect 10822 686 11124 721
rect 10822 652 10922 686
rect 10956 652 10990 686
rect 11024 652 11124 686
rect 10822 617 11124 652
rect 10822 583 10922 617
rect 10956 583 10990 617
rect 11024 583 11124 617
rect 10822 548 11124 583
rect 10822 514 10922 548
rect 10956 514 10990 548
rect 11024 514 11124 548
rect 10822 479 11124 514
rect 10822 445 10922 479
rect 10956 445 10990 479
rect 11024 445 11124 479
rect 10822 410 11124 445
rect 10822 376 10922 410
rect 10956 376 10990 410
rect 11024 376 11124 410
rect 10822 341 11124 376
rect 10822 307 10922 341
rect 10956 307 10990 341
rect 11024 307 11124 341
rect 10822 272 11124 307
rect 10822 238 10922 272
rect 10956 238 10990 272
rect 11024 238 11124 272
rect 10822 203 11124 238
rect 10822 169 10922 203
rect 10956 169 10990 203
rect 11024 169 11124 203
rect 10822 134 11124 169
rect 10822 100 10922 134
rect 10956 100 10990 134
rect 11024 100 11124 134
rect 10822 20 11124 100
tri 10822 0 10842 20 ne
rect 10842 0 11104 20
tri 11104 0 11124 20 nw
tri 11234 3080 11254 3100 se
rect 11254 3080 11516 3100
tri 11516 3080 11536 3100 sw
rect 11234 3000 11536 3080
rect 11234 790 11334 3000
rect 11436 790 11536 3000
rect 11234 755 11536 790
rect 11234 721 11334 755
rect 11368 721 11402 755
rect 11436 721 11536 755
rect 11234 686 11536 721
rect 11234 652 11334 686
rect 11368 652 11402 686
rect 11436 652 11536 686
rect 11234 617 11536 652
rect 11234 583 11334 617
rect 11368 583 11402 617
rect 11436 583 11536 617
rect 11234 548 11536 583
rect 11234 514 11334 548
rect 11368 514 11402 548
rect 11436 514 11536 548
rect 11234 479 11536 514
rect 11234 445 11334 479
rect 11368 445 11402 479
rect 11436 445 11536 479
rect 11234 410 11536 445
rect 11234 376 11334 410
rect 11368 376 11402 410
rect 11436 376 11536 410
rect 11234 341 11536 376
rect 11234 307 11334 341
rect 11368 307 11402 341
rect 11436 307 11536 341
rect 11234 272 11536 307
rect 11234 238 11334 272
rect 11368 238 11402 272
rect 11436 238 11536 272
rect 11234 203 11536 238
rect 11234 169 11334 203
rect 11368 169 11402 203
rect 11436 169 11536 203
rect 11234 134 11536 169
rect 11234 100 11334 134
rect 11368 100 11402 134
rect 11436 100 11536 134
rect 11234 20 11536 100
tri 11234 0 11254 20 ne
rect 11254 0 11516 20
tri 11516 0 11536 20 nw
tri 11646 3080 11666 3100 se
rect 11666 3080 11928 3100
tri 11928 3080 11948 3100 sw
rect 11646 3000 11948 3080
rect 11646 790 11746 3000
rect 11848 790 11948 3000
rect 11646 755 11948 790
rect 11646 721 11746 755
rect 11780 721 11814 755
rect 11848 721 11948 755
rect 11646 686 11948 721
rect 11646 652 11746 686
rect 11780 652 11814 686
rect 11848 652 11948 686
rect 11646 617 11948 652
rect 11646 583 11746 617
rect 11780 583 11814 617
rect 11848 583 11948 617
rect 11646 548 11948 583
rect 11646 514 11746 548
rect 11780 514 11814 548
rect 11848 514 11948 548
rect 11646 479 11948 514
rect 11646 445 11746 479
rect 11780 445 11814 479
rect 11848 445 11948 479
rect 11646 410 11948 445
rect 11646 376 11746 410
rect 11780 376 11814 410
rect 11848 376 11948 410
rect 11646 341 11948 376
rect 11646 307 11746 341
rect 11780 307 11814 341
rect 11848 307 11948 341
rect 11646 272 11948 307
rect 11646 238 11746 272
rect 11780 238 11814 272
rect 11848 238 11948 272
rect 11646 203 11948 238
rect 11646 169 11746 203
rect 11780 169 11814 203
rect 11848 169 11948 203
rect 11646 134 11948 169
rect 11646 100 11746 134
rect 11780 100 11814 134
rect 11848 100 11948 134
rect 11646 20 11948 100
tri 11646 0 11666 20 ne
rect 11666 0 11928 20
tri 11928 0 11948 20 nw
tri 12058 3080 12078 3100 se
rect 12078 3080 12340 3100
tri 12340 3080 12360 3100 sw
rect 12058 3000 12360 3080
rect 12058 790 12158 3000
rect 12260 790 12360 3000
rect 12058 755 12360 790
rect 12058 721 12158 755
rect 12192 721 12226 755
rect 12260 721 12360 755
rect 12058 686 12360 721
rect 12058 652 12158 686
rect 12192 652 12226 686
rect 12260 652 12360 686
rect 12058 617 12360 652
rect 12058 583 12158 617
rect 12192 583 12226 617
rect 12260 583 12360 617
rect 12058 548 12360 583
rect 12058 514 12158 548
rect 12192 514 12226 548
rect 12260 514 12360 548
rect 12058 479 12360 514
rect 12058 445 12158 479
rect 12192 445 12226 479
rect 12260 445 12360 479
rect 12058 410 12360 445
rect 12058 376 12158 410
rect 12192 376 12226 410
rect 12260 376 12360 410
rect 12058 341 12360 376
rect 12058 307 12158 341
rect 12192 307 12226 341
rect 12260 307 12360 341
rect 12058 272 12360 307
rect 12058 238 12158 272
rect 12192 238 12226 272
rect 12260 238 12360 272
rect 12058 203 12360 238
rect 12058 169 12158 203
rect 12192 169 12226 203
rect 12260 169 12360 203
rect 12058 134 12360 169
rect 12058 100 12158 134
rect 12192 100 12226 134
rect 12260 100 12360 134
rect 12058 20 12360 100
tri 12058 0 12078 20 ne
rect 12078 0 12340 20
tri 12340 0 12360 20 nw
tri 12470 3080 12490 3100 se
rect 12490 3080 12752 3100
tri 12752 3080 12772 3100 sw
rect 12470 3000 12772 3080
rect 12470 790 12570 3000
rect 12672 790 12772 3000
rect 12470 755 12772 790
rect 12470 721 12570 755
rect 12604 721 12638 755
rect 12672 721 12772 755
rect 12470 686 12772 721
rect 12470 652 12570 686
rect 12604 652 12638 686
rect 12672 652 12772 686
rect 12470 617 12772 652
rect 12470 583 12570 617
rect 12604 583 12638 617
rect 12672 583 12772 617
rect 12470 548 12772 583
rect 12470 514 12570 548
rect 12604 514 12638 548
rect 12672 514 12772 548
rect 12470 479 12772 514
rect 12470 445 12570 479
rect 12604 445 12638 479
rect 12672 445 12772 479
rect 12470 410 12772 445
rect 12470 376 12570 410
rect 12604 376 12638 410
rect 12672 376 12772 410
rect 12470 341 12772 376
rect 12470 307 12570 341
rect 12604 307 12638 341
rect 12672 307 12772 341
rect 12470 272 12772 307
rect 12470 238 12570 272
rect 12604 238 12638 272
rect 12672 238 12772 272
rect 12470 203 12772 238
rect 12470 169 12570 203
rect 12604 169 12638 203
rect 12672 169 12772 203
rect 12470 134 12772 169
rect 12470 100 12570 134
rect 12604 100 12638 134
rect 12672 100 12772 134
rect 12470 20 12772 100
tri 12470 0 12490 20 ne
rect 12490 0 12752 20
tri 12752 0 12772 20 nw
tri 12882 3080 12902 3100 se
rect 12902 3080 13114 3100
rect 12882 3000 13114 3080
rect 12882 790 12982 3000
rect 13084 790 13114 3000
rect 12882 755 13114 790
rect 12882 721 12982 755
rect 13016 721 13050 755
rect 13084 721 13114 755
rect 12882 686 13114 721
rect 12882 652 12982 686
rect 13016 652 13050 686
rect 13084 652 13114 686
rect 12882 617 13114 652
rect 12882 583 12982 617
rect 13016 583 13050 617
rect 13084 583 13114 617
rect 12882 548 13114 583
rect 12882 514 12982 548
rect 13016 514 13050 548
rect 13084 514 13114 548
rect 12882 479 13114 514
rect 12882 445 12982 479
rect 13016 445 13050 479
rect 13084 445 13114 479
rect 12882 410 13114 445
rect 12882 376 12982 410
rect 13016 376 13050 410
rect 13084 376 13114 410
rect 12882 341 13114 376
rect 12882 307 12982 341
rect 13016 307 13050 341
rect 13084 307 13114 341
rect 12882 272 13114 307
rect 12882 238 12982 272
rect 13016 238 13050 272
rect 13084 238 13114 272
rect 12882 203 13114 238
rect 12882 169 12982 203
rect 13016 169 13050 203
rect 13084 169 13114 203
rect 12882 134 13114 169
rect 12882 100 12982 134
rect 13016 100 13050 134
rect 13084 100 13114 134
rect 12882 20 13114 100
tri 12882 0 12902 20 ne
rect 12902 0 13114 20
<< mvpdiffc >>
rect -202 790 -100 3000
rect -202 721 -168 755
rect -134 721 -100 755
rect -202 652 -168 686
rect -134 652 -100 686
rect -202 583 -168 617
rect -134 583 -100 617
rect -202 514 -168 548
rect -134 514 -100 548
rect -202 445 -168 479
rect -134 445 -100 479
rect -202 376 -168 410
rect -134 376 -100 410
rect -202 307 -168 341
rect -134 307 -100 341
rect -202 238 -168 272
rect -134 238 -100 272
rect -202 169 -168 203
rect -134 169 -100 203
rect -202 100 -168 134
rect -134 100 -100 134
rect 210 790 312 3000
rect 210 721 244 755
rect 278 721 312 755
rect 210 652 244 686
rect 278 652 312 686
rect 210 583 244 617
rect 278 583 312 617
rect 210 514 244 548
rect 278 514 312 548
rect 210 445 244 479
rect 278 445 312 479
rect 210 376 244 410
rect 278 376 312 410
rect 210 307 244 341
rect 278 307 312 341
rect 210 238 244 272
rect 278 238 312 272
rect 210 169 244 203
rect 278 169 312 203
rect 210 100 244 134
rect 278 100 312 134
rect 622 790 724 3000
rect 622 721 656 755
rect 690 721 724 755
rect 622 652 656 686
rect 690 652 724 686
rect 622 583 656 617
rect 690 583 724 617
rect 622 514 656 548
rect 690 514 724 548
rect 622 445 656 479
rect 690 445 724 479
rect 622 376 656 410
rect 690 376 724 410
rect 622 307 656 341
rect 690 307 724 341
rect 622 238 656 272
rect 690 238 724 272
rect 622 169 656 203
rect 690 169 724 203
rect 622 100 656 134
rect 690 100 724 134
rect 1034 790 1136 3000
rect 1034 721 1068 755
rect 1102 721 1136 755
rect 1034 652 1068 686
rect 1102 652 1136 686
rect 1034 583 1068 617
rect 1102 583 1136 617
rect 1034 514 1068 548
rect 1102 514 1136 548
rect 1034 445 1068 479
rect 1102 445 1136 479
rect 1034 376 1068 410
rect 1102 376 1136 410
rect 1034 307 1068 341
rect 1102 307 1136 341
rect 1034 238 1068 272
rect 1102 238 1136 272
rect 1034 169 1068 203
rect 1102 169 1136 203
rect 1034 100 1068 134
rect 1102 100 1136 134
rect 1446 790 1548 3000
rect 1446 721 1480 755
rect 1514 721 1548 755
rect 1446 652 1480 686
rect 1514 652 1548 686
rect 1446 583 1480 617
rect 1514 583 1548 617
rect 1446 514 1480 548
rect 1514 514 1548 548
rect 1446 445 1480 479
rect 1514 445 1548 479
rect 1446 376 1480 410
rect 1514 376 1548 410
rect 1446 307 1480 341
rect 1514 307 1548 341
rect 1446 238 1480 272
rect 1514 238 1548 272
rect 1446 169 1480 203
rect 1514 169 1548 203
rect 1446 100 1480 134
rect 1514 100 1548 134
rect 1858 790 1960 3000
rect 1858 721 1892 755
rect 1926 721 1960 755
rect 1858 652 1892 686
rect 1926 652 1960 686
rect 1858 583 1892 617
rect 1926 583 1960 617
rect 1858 514 1892 548
rect 1926 514 1960 548
rect 1858 445 1892 479
rect 1926 445 1960 479
rect 1858 376 1892 410
rect 1926 376 1960 410
rect 1858 307 1892 341
rect 1926 307 1960 341
rect 1858 238 1892 272
rect 1926 238 1960 272
rect 1858 169 1892 203
rect 1926 169 1960 203
rect 1858 100 1892 134
rect 1926 100 1960 134
rect 2270 790 2372 3000
rect 2270 721 2304 755
rect 2338 721 2372 755
rect 2270 652 2304 686
rect 2338 652 2372 686
rect 2270 583 2304 617
rect 2338 583 2372 617
rect 2270 514 2304 548
rect 2338 514 2372 548
rect 2270 445 2304 479
rect 2338 445 2372 479
rect 2270 376 2304 410
rect 2338 376 2372 410
rect 2270 307 2304 341
rect 2338 307 2372 341
rect 2270 238 2304 272
rect 2338 238 2372 272
rect 2270 169 2304 203
rect 2338 169 2372 203
rect 2270 100 2304 134
rect 2338 100 2372 134
rect 2682 790 2784 3000
rect 2682 721 2716 755
rect 2750 721 2784 755
rect 2682 652 2716 686
rect 2750 652 2784 686
rect 2682 583 2716 617
rect 2750 583 2784 617
rect 2682 514 2716 548
rect 2750 514 2784 548
rect 2682 445 2716 479
rect 2750 445 2784 479
rect 2682 376 2716 410
rect 2750 376 2784 410
rect 2682 307 2716 341
rect 2750 307 2784 341
rect 2682 238 2716 272
rect 2750 238 2784 272
rect 2682 169 2716 203
rect 2750 169 2784 203
rect 2682 100 2716 134
rect 2750 100 2784 134
rect 3094 790 3196 3000
rect 3094 721 3128 755
rect 3162 721 3196 755
rect 3094 652 3128 686
rect 3162 652 3196 686
rect 3094 583 3128 617
rect 3162 583 3196 617
rect 3094 514 3128 548
rect 3162 514 3196 548
rect 3094 445 3128 479
rect 3162 445 3196 479
rect 3094 376 3128 410
rect 3162 376 3196 410
rect 3094 307 3128 341
rect 3162 307 3196 341
rect 3094 238 3128 272
rect 3162 238 3196 272
rect 3094 169 3128 203
rect 3162 169 3196 203
rect 3094 100 3128 134
rect 3162 100 3196 134
rect 3506 790 3608 3000
rect 3506 721 3540 755
rect 3574 721 3608 755
rect 3506 652 3540 686
rect 3574 652 3608 686
rect 3506 583 3540 617
rect 3574 583 3608 617
rect 3506 514 3540 548
rect 3574 514 3608 548
rect 3506 445 3540 479
rect 3574 445 3608 479
rect 3506 376 3540 410
rect 3574 376 3608 410
rect 3506 307 3540 341
rect 3574 307 3608 341
rect 3506 238 3540 272
rect 3574 238 3608 272
rect 3506 169 3540 203
rect 3574 169 3608 203
rect 3506 100 3540 134
rect 3574 100 3608 134
rect 3918 790 4020 3000
rect 3918 721 3952 755
rect 3986 721 4020 755
rect 3918 652 3952 686
rect 3986 652 4020 686
rect 3918 583 3952 617
rect 3986 583 4020 617
rect 3918 514 3952 548
rect 3986 514 4020 548
rect 3918 445 3952 479
rect 3986 445 4020 479
rect 3918 376 3952 410
rect 3986 376 4020 410
rect 3918 307 3952 341
rect 3986 307 4020 341
rect 3918 238 3952 272
rect 3986 238 4020 272
rect 3918 169 3952 203
rect 3986 169 4020 203
rect 3918 100 3952 134
rect 3986 100 4020 134
rect 4330 790 4432 3000
rect 4330 721 4364 755
rect 4398 721 4432 755
rect 4330 652 4364 686
rect 4398 652 4432 686
rect 4330 583 4364 617
rect 4398 583 4432 617
rect 4330 514 4364 548
rect 4398 514 4432 548
rect 4330 445 4364 479
rect 4398 445 4432 479
rect 4330 376 4364 410
rect 4398 376 4432 410
rect 4330 307 4364 341
rect 4398 307 4432 341
rect 4330 238 4364 272
rect 4398 238 4432 272
rect 4330 169 4364 203
rect 4398 169 4432 203
rect 4330 100 4364 134
rect 4398 100 4432 134
rect 4742 790 4844 3000
rect 4742 721 4776 755
rect 4810 721 4844 755
rect 4742 652 4776 686
rect 4810 652 4844 686
rect 4742 583 4776 617
rect 4810 583 4844 617
rect 4742 514 4776 548
rect 4810 514 4844 548
rect 4742 445 4776 479
rect 4810 445 4844 479
rect 4742 376 4776 410
rect 4810 376 4844 410
rect 4742 307 4776 341
rect 4810 307 4844 341
rect 4742 238 4776 272
rect 4810 238 4844 272
rect 4742 169 4776 203
rect 4810 169 4844 203
rect 4742 100 4776 134
rect 4810 100 4844 134
rect 5154 790 5256 3000
rect 5154 721 5188 755
rect 5222 721 5256 755
rect 5154 652 5188 686
rect 5222 652 5256 686
rect 5154 583 5188 617
rect 5222 583 5256 617
rect 5154 514 5188 548
rect 5222 514 5256 548
rect 5154 445 5188 479
rect 5222 445 5256 479
rect 5154 376 5188 410
rect 5222 376 5256 410
rect 5154 307 5188 341
rect 5222 307 5256 341
rect 5154 238 5188 272
rect 5222 238 5256 272
rect 5154 169 5188 203
rect 5222 169 5256 203
rect 5154 100 5188 134
rect 5222 100 5256 134
rect 5566 790 5668 3000
rect 5566 721 5600 755
rect 5634 721 5668 755
rect 5566 652 5600 686
rect 5634 652 5668 686
rect 5566 583 5600 617
rect 5634 583 5668 617
rect 5566 514 5600 548
rect 5634 514 5668 548
rect 5566 445 5600 479
rect 5634 445 5668 479
rect 5566 376 5600 410
rect 5634 376 5668 410
rect 5566 307 5600 341
rect 5634 307 5668 341
rect 5566 238 5600 272
rect 5634 238 5668 272
rect 5566 169 5600 203
rect 5634 169 5668 203
rect 5566 100 5600 134
rect 5634 100 5668 134
rect 5978 790 6080 3000
rect 5978 721 6012 755
rect 6046 721 6080 755
rect 5978 652 6012 686
rect 6046 652 6080 686
rect 5978 583 6012 617
rect 6046 583 6080 617
rect 5978 514 6012 548
rect 6046 514 6080 548
rect 5978 445 6012 479
rect 6046 445 6080 479
rect 5978 376 6012 410
rect 6046 376 6080 410
rect 5978 307 6012 341
rect 6046 307 6080 341
rect 5978 238 6012 272
rect 6046 238 6080 272
rect 5978 169 6012 203
rect 6046 169 6080 203
rect 5978 100 6012 134
rect 6046 100 6080 134
rect 6390 790 6492 3000
rect 6390 721 6424 755
rect 6458 721 6492 755
rect 6390 652 6424 686
rect 6458 652 6492 686
rect 6390 583 6424 617
rect 6458 583 6492 617
rect 6390 514 6424 548
rect 6458 514 6492 548
rect 6390 445 6424 479
rect 6458 445 6492 479
rect 6390 376 6424 410
rect 6458 376 6492 410
rect 6390 307 6424 341
rect 6458 307 6492 341
rect 6390 238 6424 272
rect 6458 238 6492 272
rect 6390 169 6424 203
rect 6458 169 6492 203
rect 6390 100 6424 134
rect 6458 100 6492 134
rect 6802 790 6904 3000
rect 6802 721 6836 755
rect 6870 721 6904 755
rect 6802 652 6836 686
rect 6870 652 6904 686
rect 6802 583 6836 617
rect 6870 583 6904 617
rect 6802 514 6836 548
rect 6870 514 6904 548
rect 6802 445 6836 479
rect 6870 445 6904 479
rect 6802 376 6836 410
rect 6870 376 6904 410
rect 6802 307 6836 341
rect 6870 307 6904 341
rect 6802 238 6836 272
rect 6870 238 6904 272
rect 6802 169 6836 203
rect 6870 169 6904 203
rect 6802 100 6836 134
rect 6870 100 6904 134
rect 7214 790 7316 3000
rect 7214 721 7248 755
rect 7282 721 7316 755
rect 7214 652 7248 686
rect 7282 652 7316 686
rect 7214 583 7248 617
rect 7282 583 7316 617
rect 7214 514 7248 548
rect 7282 514 7316 548
rect 7214 445 7248 479
rect 7282 445 7316 479
rect 7214 376 7248 410
rect 7282 376 7316 410
rect 7214 307 7248 341
rect 7282 307 7316 341
rect 7214 238 7248 272
rect 7282 238 7316 272
rect 7214 169 7248 203
rect 7282 169 7316 203
rect 7214 100 7248 134
rect 7282 100 7316 134
rect 7626 790 7728 3000
rect 7626 721 7660 755
rect 7694 721 7728 755
rect 7626 652 7660 686
rect 7694 652 7728 686
rect 7626 583 7660 617
rect 7694 583 7728 617
rect 7626 514 7660 548
rect 7694 514 7728 548
rect 7626 445 7660 479
rect 7694 445 7728 479
rect 7626 376 7660 410
rect 7694 376 7728 410
rect 7626 307 7660 341
rect 7694 307 7728 341
rect 7626 238 7660 272
rect 7694 238 7728 272
rect 7626 169 7660 203
rect 7694 169 7728 203
rect 7626 100 7660 134
rect 7694 100 7728 134
rect 8038 790 8140 3000
rect 8038 721 8072 755
rect 8106 721 8140 755
rect 8038 652 8072 686
rect 8106 652 8140 686
rect 8038 583 8072 617
rect 8106 583 8140 617
rect 8038 514 8072 548
rect 8106 514 8140 548
rect 8038 445 8072 479
rect 8106 445 8140 479
rect 8038 376 8072 410
rect 8106 376 8140 410
rect 8038 307 8072 341
rect 8106 307 8140 341
rect 8038 238 8072 272
rect 8106 238 8140 272
rect 8038 169 8072 203
rect 8106 169 8140 203
rect 8038 100 8072 134
rect 8106 100 8140 134
rect 8450 790 8552 3000
rect 8450 721 8484 755
rect 8518 721 8552 755
rect 8450 652 8484 686
rect 8518 652 8552 686
rect 8450 583 8484 617
rect 8518 583 8552 617
rect 8450 514 8484 548
rect 8518 514 8552 548
rect 8450 445 8484 479
rect 8518 445 8552 479
rect 8450 376 8484 410
rect 8518 376 8552 410
rect 8450 307 8484 341
rect 8518 307 8552 341
rect 8450 238 8484 272
rect 8518 238 8552 272
rect 8450 169 8484 203
rect 8518 169 8552 203
rect 8450 100 8484 134
rect 8518 100 8552 134
rect 8862 790 8964 3000
rect 8862 721 8896 755
rect 8930 721 8964 755
rect 8862 652 8896 686
rect 8930 652 8964 686
rect 8862 583 8896 617
rect 8930 583 8964 617
rect 8862 514 8896 548
rect 8930 514 8964 548
rect 8862 445 8896 479
rect 8930 445 8964 479
rect 8862 376 8896 410
rect 8930 376 8964 410
rect 8862 307 8896 341
rect 8930 307 8964 341
rect 8862 238 8896 272
rect 8930 238 8964 272
rect 8862 169 8896 203
rect 8930 169 8964 203
rect 8862 100 8896 134
rect 8930 100 8964 134
rect 9274 790 9376 3000
rect 9274 721 9308 755
rect 9342 721 9376 755
rect 9274 652 9308 686
rect 9342 652 9376 686
rect 9274 583 9308 617
rect 9342 583 9376 617
rect 9274 514 9308 548
rect 9342 514 9376 548
rect 9274 445 9308 479
rect 9342 445 9376 479
rect 9274 376 9308 410
rect 9342 376 9376 410
rect 9274 307 9308 341
rect 9342 307 9376 341
rect 9274 238 9308 272
rect 9342 238 9376 272
rect 9274 169 9308 203
rect 9342 169 9376 203
rect 9274 100 9308 134
rect 9342 100 9376 134
rect 9686 790 9788 3000
rect 9686 721 9720 755
rect 9754 721 9788 755
rect 9686 652 9720 686
rect 9754 652 9788 686
rect 9686 583 9720 617
rect 9754 583 9788 617
rect 9686 514 9720 548
rect 9754 514 9788 548
rect 9686 445 9720 479
rect 9754 445 9788 479
rect 9686 376 9720 410
rect 9754 376 9788 410
rect 9686 307 9720 341
rect 9754 307 9788 341
rect 9686 238 9720 272
rect 9754 238 9788 272
rect 9686 169 9720 203
rect 9754 169 9788 203
rect 9686 100 9720 134
rect 9754 100 9788 134
rect 10098 790 10200 3000
rect 10098 721 10132 755
rect 10166 721 10200 755
rect 10098 652 10132 686
rect 10166 652 10200 686
rect 10098 583 10132 617
rect 10166 583 10200 617
rect 10098 514 10132 548
rect 10166 514 10200 548
rect 10098 445 10132 479
rect 10166 445 10200 479
rect 10098 376 10132 410
rect 10166 376 10200 410
rect 10098 307 10132 341
rect 10166 307 10200 341
rect 10098 238 10132 272
rect 10166 238 10200 272
rect 10098 169 10132 203
rect 10166 169 10200 203
rect 10098 100 10132 134
rect 10166 100 10200 134
rect 10510 790 10612 3000
rect 10510 721 10544 755
rect 10578 721 10612 755
rect 10510 652 10544 686
rect 10578 652 10612 686
rect 10510 583 10544 617
rect 10578 583 10612 617
rect 10510 514 10544 548
rect 10578 514 10612 548
rect 10510 445 10544 479
rect 10578 445 10612 479
rect 10510 376 10544 410
rect 10578 376 10612 410
rect 10510 307 10544 341
rect 10578 307 10612 341
rect 10510 238 10544 272
rect 10578 238 10612 272
rect 10510 169 10544 203
rect 10578 169 10612 203
rect 10510 100 10544 134
rect 10578 100 10612 134
rect 10922 790 11024 3000
rect 10922 721 10956 755
rect 10990 721 11024 755
rect 10922 652 10956 686
rect 10990 652 11024 686
rect 10922 583 10956 617
rect 10990 583 11024 617
rect 10922 514 10956 548
rect 10990 514 11024 548
rect 10922 445 10956 479
rect 10990 445 11024 479
rect 10922 376 10956 410
rect 10990 376 11024 410
rect 10922 307 10956 341
rect 10990 307 11024 341
rect 10922 238 10956 272
rect 10990 238 11024 272
rect 10922 169 10956 203
rect 10990 169 11024 203
rect 10922 100 10956 134
rect 10990 100 11024 134
rect 11334 790 11436 3000
rect 11334 721 11368 755
rect 11402 721 11436 755
rect 11334 652 11368 686
rect 11402 652 11436 686
rect 11334 583 11368 617
rect 11402 583 11436 617
rect 11334 514 11368 548
rect 11402 514 11436 548
rect 11334 445 11368 479
rect 11402 445 11436 479
rect 11334 376 11368 410
rect 11402 376 11436 410
rect 11334 307 11368 341
rect 11402 307 11436 341
rect 11334 238 11368 272
rect 11402 238 11436 272
rect 11334 169 11368 203
rect 11402 169 11436 203
rect 11334 100 11368 134
rect 11402 100 11436 134
rect 11746 790 11848 3000
rect 11746 721 11780 755
rect 11814 721 11848 755
rect 11746 652 11780 686
rect 11814 652 11848 686
rect 11746 583 11780 617
rect 11814 583 11848 617
rect 11746 514 11780 548
rect 11814 514 11848 548
rect 11746 445 11780 479
rect 11814 445 11848 479
rect 11746 376 11780 410
rect 11814 376 11848 410
rect 11746 307 11780 341
rect 11814 307 11848 341
rect 11746 238 11780 272
rect 11814 238 11848 272
rect 11746 169 11780 203
rect 11814 169 11848 203
rect 11746 100 11780 134
rect 11814 100 11848 134
rect 12158 790 12260 3000
rect 12158 721 12192 755
rect 12226 721 12260 755
rect 12158 652 12192 686
rect 12226 652 12260 686
rect 12158 583 12192 617
rect 12226 583 12260 617
rect 12158 514 12192 548
rect 12226 514 12260 548
rect 12158 445 12192 479
rect 12226 445 12260 479
rect 12158 376 12192 410
rect 12226 376 12260 410
rect 12158 307 12192 341
rect 12226 307 12260 341
rect 12158 238 12192 272
rect 12226 238 12260 272
rect 12158 169 12192 203
rect 12226 169 12260 203
rect 12158 100 12192 134
rect 12226 100 12260 134
rect 12570 790 12672 3000
rect 12570 721 12604 755
rect 12638 721 12672 755
rect 12570 652 12604 686
rect 12638 652 12672 686
rect 12570 583 12604 617
rect 12638 583 12672 617
rect 12570 514 12604 548
rect 12638 514 12672 548
rect 12570 445 12604 479
rect 12638 445 12672 479
rect 12570 376 12604 410
rect 12638 376 12672 410
rect 12570 307 12604 341
rect 12638 307 12672 341
rect 12570 238 12604 272
rect 12638 238 12672 272
rect 12570 169 12604 203
rect 12638 169 12672 203
rect 12570 100 12604 134
rect 12638 100 12672 134
rect 12982 790 13084 3000
rect 12982 721 13016 755
rect 13050 721 13084 755
rect 12982 652 13016 686
rect 13050 652 13084 686
rect 12982 583 13016 617
rect 13050 583 13084 617
rect 12982 514 13016 548
rect 13050 514 13084 548
rect 12982 445 13016 479
rect 13050 445 13084 479
rect 12982 376 13016 410
rect 13050 376 13084 410
rect 12982 307 13016 341
rect 13050 307 13084 341
rect 12982 238 13016 272
rect 13050 238 13084 272
rect 12982 169 13016 203
rect 13050 169 13084 203
rect 12982 100 13016 134
rect 13050 100 13084 134
<< mvpsubdiff >>
rect -1458 3880 -1390 3914
rect -1356 3880 -1321 3914
rect -1287 3880 -1252 3914
rect -1218 3880 -1183 3914
rect -1149 3880 -1114 3914
rect -1080 3880 -1045 3914
rect -1011 3880 -976 3914
rect -942 3880 -907 3914
rect -873 3880 -838 3914
rect -804 3880 -769 3914
rect -735 3880 -700 3914
rect -666 3880 -631 3914
rect -597 3880 -562 3914
rect -528 3880 -493 3914
rect -459 3880 -424 3914
rect -390 3880 -355 3914
rect -321 3880 -286 3914
rect -252 3880 -217 3914
rect -183 3880 -148 3914
rect -114 3880 -79 3914
rect -45 3880 -10 3914
rect 24 3880 59 3914
rect 93 3880 128 3914
rect 162 3880 197 3914
rect 231 3880 266 3914
rect 300 3880 335 3914
rect 369 3880 404 3914
rect 438 3880 473 3914
rect 507 3880 542 3914
rect 576 3880 611 3914
rect 645 3880 680 3914
rect 714 3880 749 3914
rect 783 3880 818 3914
rect 852 3880 887 3914
rect 921 3880 956 3914
rect 990 3880 1025 3914
rect 1059 3880 1094 3914
rect 1128 3880 1163 3914
rect 1197 3880 1232 3914
rect 1266 3880 1301 3914
rect 1335 3880 1370 3914
rect 1404 3880 1439 3914
rect 1473 3880 1508 3914
rect 1542 3880 1577 3914
rect 1611 3880 1646 3914
rect 1680 3880 1715 3914
rect 1749 3880 1784 3914
rect 1818 3880 1853 3914
rect 1887 3880 1922 3914
rect 1956 3880 1991 3914
rect 2025 3880 2060 3914
rect 2094 3880 2129 3914
rect 2163 3880 2198 3914
rect 2232 3880 2267 3914
rect 2301 3880 2336 3914
rect 2370 3880 2405 3914
rect 2439 3880 2474 3914
rect -1458 3846 2474 3880
rect -1458 3812 -1390 3846
rect -1356 3812 -1321 3846
rect -1287 3812 -1252 3846
rect -1218 3812 -1183 3846
rect -1149 3812 -1114 3846
rect -1080 3812 -1045 3846
rect -1011 3812 -976 3846
rect -942 3812 -907 3846
rect -873 3812 -838 3846
rect -804 3812 -769 3846
rect -735 3812 -700 3846
rect -666 3812 -631 3846
rect -597 3812 -562 3846
rect -528 3812 -493 3846
rect -459 3812 -424 3846
rect -390 3812 -355 3846
rect -321 3812 -286 3846
rect -252 3812 -217 3846
rect -183 3812 -148 3846
rect -114 3812 -79 3846
rect -45 3812 -10 3846
rect 24 3812 59 3846
rect 93 3812 128 3846
rect 162 3812 197 3846
rect 231 3812 266 3846
rect 300 3812 335 3846
rect 369 3812 404 3846
rect 438 3812 473 3846
rect 507 3812 542 3846
rect 576 3812 611 3846
rect 645 3812 680 3846
rect 714 3812 749 3846
rect 783 3812 818 3846
rect 852 3812 887 3846
rect 921 3812 956 3846
rect 990 3812 1025 3846
rect 1059 3812 1094 3846
rect 1128 3812 1163 3846
rect 1197 3812 1232 3846
rect 1266 3812 1301 3846
rect 1335 3812 1370 3846
rect 1404 3812 1439 3846
rect 1473 3812 1508 3846
rect 1542 3812 1577 3846
rect 1611 3812 1646 3846
rect 1680 3812 1715 3846
rect 1749 3812 1784 3846
rect 1818 3812 1853 3846
rect 1887 3812 1922 3846
rect 1956 3812 1991 3846
rect 2025 3812 2060 3846
rect 2094 3812 2129 3846
rect 2163 3812 2198 3846
rect 2232 3812 2267 3846
rect 2301 3812 2336 3846
rect 2370 3812 2405 3846
rect 2439 3812 2474 3846
rect -1458 3778 2474 3812
rect -1458 3744 -1390 3778
rect -1356 3744 -1321 3778
rect -1287 3744 -1252 3778
rect -1218 3744 -1183 3778
rect -1149 3744 -1114 3778
rect -1080 3744 -1045 3778
rect -1011 3744 -976 3778
rect -942 3744 -907 3778
rect -873 3744 -838 3778
rect -804 3744 -769 3778
rect -735 3744 -700 3778
rect -666 3744 -631 3778
rect -597 3744 -562 3778
rect -528 3744 -493 3778
rect -459 3744 -424 3778
rect -390 3744 -355 3778
rect -321 3744 -286 3778
rect -252 3744 -217 3778
rect -183 3744 -148 3778
rect -114 3744 -79 3778
rect -45 3744 -10 3778
rect 24 3744 59 3778
rect 93 3744 128 3778
rect 162 3744 197 3778
rect 231 3744 266 3778
rect 300 3744 335 3778
rect 369 3744 404 3778
rect 438 3744 473 3778
rect 507 3744 542 3778
rect 576 3744 611 3778
rect 645 3744 680 3778
rect 714 3744 749 3778
rect 783 3744 818 3778
rect 852 3744 887 3778
rect 921 3744 956 3778
rect 990 3744 1025 3778
rect 1059 3744 1094 3778
rect 1128 3744 1163 3778
rect 1197 3744 1232 3778
rect 1266 3744 1301 3778
rect 1335 3744 1370 3778
rect 1404 3744 1439 3778
rect 1473 3744 1508 3778
rect 1542 3744 1577 3778
rect 1611 3744 1646 3778
rect 1680 3744 1715 3778
rect 1749 3744 1784 3778
rect 1818 3744 1853 3778
rect 1887 3744 1922 3778
rect 1956 3744 1991 3778
rect 2025 3744 2060 3778
rect 2094 3744 2129 3778
rect 2163 3744 2198 3778
rect 2232 3744 2267 3778
rect 2301 3744 2336 3778
rect 2370 3744 2405 3778
rect 2439 3744 2474 3778
rect 14272 3744 14340 3914
rect -1458 3676 -1288 3744
rect 14170 3676 14340 3744
rect -1458 -473 -1288 -438
rect -1424 -507 -1390 -473
rect -1356 -507 -1322 -473
rect -1458 -542 -1288 -507
rect -1424 -576 -1390 -542
rect -1356 -576 -1322 -542
rect -1458 -644 -1288 -576
rect 14170 -473 14340 -438
rect 14204 -507 14238 -473
rect 14272 -507 14306 -473
rect 14170 -542 14340 -507
rect 14204 -576 14238 -542
rect 14272 -576 14306 -542
rect 14170 -644 14340 -576
rect -1458 -678 -1390 -644
rect -1356 -678 -1321 -644
rect -1287 -678 -1252 -644
rect -1218 -678 -1183 -644
rect -1149 -678 -1114 -644
rect -1080 -678 -1045 -644
rect -1011 -678 -976 -644
rect -942 -678 -907 -644
rect -873 -678 -838 -644
rect -804 -678 -769 -644
rect -735 -678 -700 -644
rect -666 -678 -631 -644
rect -597 -678 -562 -644
rect -528 -678 -493 -644
rect -459 -678 -424 -644
rect -390 -678 -355 -644
rect -321 -678 -286 -644
rect -252 -678 -217 -644
rect -183 -678 -148 -644
rect -114 -678 -79 -644
rect -45 -678 -10 -644
rect 24 -678 59 -644
rect 93 -678 128 -644
rect 162 -678 197 -644
rect 231 -678 266 -644
rect 300 -678 335 -644
rect 369 -678 404 -644
rect 438 -678 473 -644
rect 507 -678 542 -644
rect 576 -678 611 -644
rect 645 -678 680 -644
rect 714 -678 749 -644
rect 783 -678 818 -644
rect 852 -678 887 -644
rect 921 -678 956 -644
rect 990 -678 1025 -644
rect 1059 -678 1094 -644
rect 1128 -678 1163 -644
rect 1197 -678 1232 -644
rect 1266 -678 1301 -644
rect 1335 -678 1370 -644
rect 1404 -678 1439 -644
rect 1473 -678 1508 -644
rect 1542 -678 1577 -644
rect 1611 -678 1646 -644
rect 1680 -678 1715 -644
rect 1749 -678 1784 -644
rect 1818 -678 1853 -644
rect 1887 -678 1922 -644
rect 1956 -678 1991 -644
rect 2025 -678 2060 -644
rect 2094 -678 2129 -644
rect 2163 -678 2198 -644
rect 2232 -678 2267 -644
rect 2301 -678 2336 -644
rect 2370 -678 2405 -644
rect 2439 -678 2474 -644
rect -1458 -712 2474 -678
rect -1458 -746 -1390 -712
rect -1356 -746 -1321 -712
rect -1287 -746 -1252 -712
rect -1218 -746 -1183 -712
rect -1149 -746 -1114 -712
rect -1080 -746 -1045 -712
rect -1011 -746 -976 -712
rect -942 -746 -907 -712
rect -873 -746 -838 -712
rect -804 -746 -769 -712
rect -735 -746 -700 -712
rect -666 -746 -631 -712
rect -597 -746 -562 -712
rect -528 -746 -493 -712
rect -459 -746 -424 -712
rect -390 -746 -355 -712
rect -321 -746 -286 -712
rect -252 -746 -217 -712
rect -183 -746 -148 -712
rect -114 -746 -79 -712
rect -45 -746 -10 -712
rect 24 -746 59 -712
rect 93 -746 128 -712
rect 162 -746 197 -712
rect 231 -746 266 -712
rect 300 -746 335 -712
rect 369 -746 404 -712
rect 438 -746 473 -712
rect 507 -746 542 -712
rect 576 -746 611 -712
rect 645 -746 680 -712
rect 714 -746 749 -712
rect 783 -746 818 -712
rect 852 -746 887 -712
rect 921 -746 956 -712
rect 990 -746 1025 -712
rect 1059 -746 1094 -712
rect 1128 -746 1163 -712
rect 1197 -746 1232 -712
rect 1266 -746 1301 -712
rect 1335 -746 1370 -712
rect 1404 -746 1439 -712
rect 1473 -746 1508 -712
rect 1542 -746 1577 -712
rect 1611 -746 1646 -712
rect 1680 -746 1715 -712
rect 1749 -746 1784 -712
rect 1818 -746 1853 -712
rect 1887 -746 1922 -712
rect 1956 -746 1991 -712
rect 2025 -746 2060 -712
rect 2094 -746 2129 -712
rect 2163 -746 2198 -712
rect 2232 -746 2267 -712
rect 2301 -746 2336 -712
rect 2370 -746 2405 -712
rect 2439 -746 2474 -712
rect -1458 -780 2474 -746
rect -1458 -814 -1390 -780
rect -1356 -814 -1321 -780
rect -1287 -814 -1252 -780
rect -1218 -814 -1183 -780
rect -1149 -814 -1114 -780
rect -1080 -814 -1045 -780
rect -1011 -814 -976 -780
rect -942 -814 -907 -780
rect -873 -814 -838 -780
rect -804 -814 -769 -780
rect -735 -814 -700 -780
rect -666 -814 -631 -780
rect -597 -814 -562 -780
rect -528 -814 -493 -780
rect -459 -814 -424 -780
rect -390 -814 -355 -780
rect -321 -814 -286 -780
rect -252 -814 -217 -780
rect -183 -814 -148 -780
rect -114 -814 -79 -780
rect -45 -814 -10 -780
rect 24 -814 59 -780
rect 93 -814 128 -780
rect 162 -814 197 -780
rect 231 -814 266 -780
rect 300 -814 335 -780
rect 369 -814 404 -780
rect 438 -814 473 -780
rect 507 -814 542 -780
rect 576 -814 611 -780
rect 645 -814 680 -780
rect 714 -814 749 -780
rect 783 -814 818 -780
rect 852 -814 887 -780
rect 921 -814 956 -780
rect 990 -814 1025 -780
rect 1059 -814 1094 -780
rect 1128 -814 1163 -780
rect 1197 -814 1232 -780
rect 1266 -814 1301 -780
rect 1335 -814 1370 -780
rect 1404 -814 1439 -780
rect 1473 -814 1508 -780
rect 1542 -814 1577 -780
rect 1611 -814 1646 -780
rect 1680 -814 1715 -780
rect 1749 -814 1784 -780
rect 1818 -814 1853 -780
rect 1887 -814 1922 -780
rect 1956 -814 1991 -780
rect 2025 -814 2060 -780
rect 2094 -814 2129 -780
rect 2163 -814 2198 -780
rect 2232 -814 2267 -780
rect 2301 -814 2336 -780
rect 2370 -814 2405 -780
rect 2439 -814 2474 -780
rect 14272 -814 14340 -644
<< mvnsubdiff >>
rect -1088 3510 -1020 3544
rect -986 3510 -951 3544
rect -917 3510 -882 3544
rect -848 3510 -813 3544
rect -779 3510 -744 3544
rect -710 3510 -675 3544
rect -641 3510 -606 3544
rect -572 3510 -537 3544
rect -503 3510 -468 3544
rect -434 3510 -399 3544
rect -365 3510 -330 3544
rect -296 3510 -261 3544
rect -227 3510 -192 3544
rect -158 3510 -123 3544
rect -89 3510 -54 3544
rect -20 3510 15 3544
rect 49 3510 84 3544
rect 118 3510 153 3544
rect 187 3510 222 3544
rect 256 3510 291 3544
rect 325 3510 360 3544
rect 394 3510 429 3544
rect 463 3510 498 3544
rect 532 3510 567 3544
rect 601 3510 636 3544
rect 670 3510 705 3544
rect 739 3510 774 3544
rect 808 3510 843 3544
rect 877 3510 912 3544
rect 946 3510 981 3544
rect 1015 3510 1050 3544
rect 1084 3510 1119 3544
rect 1153 3510 1188 3544
rect 1222 3510 1257 3544
rect 1291 3510 1326 3544
rect 1360 3510 1395 3544
rect 1429 3510 1464 3544
rect 1498 3510 1533 3544
rect 1567 3510 1602 3544
rect 1636 3510 1671 3544
rect 1705 3510 1740 3544
rect 1774 3510 1809 3544
rect 1843 3510 1878 3544
rect 1912 3510 1947 3544
rect 1981 3510 2016 3544
rect 2050 3510 2085 3544
rect 2119 3510 2154 3544
rect 2188 3510 2223 3544
rect 2257 3510 2292 3544
rect 2326 3510 2361 3544
rect 2395 3510 2430 3544
rect 2464 3510 2499 3544
rect 2533 3510 2568 3544
rect 2602 3510 2637 3544
rect 2671 3510 2706 3544
rect 2740 3510 2775 3544
rect 2809 3510 2844 3544
rect 2878 3510 2913 3544
rect 2947 3510 2982 3544
rect 3016 3510 3051 3544
rect 3085 3510 3120 3544
rect 3154 3510 3189 3544
rect 3223 3510 3258 3544
rect 3292 3510 3327 3544
rect 3361 3510 3396 3544
rect -1088 3476 3396 3510
rect -1088 3442 -1020 3476
rect -986 3442 -951 3476
rect -917 3442 -882 3476
rect -848 3442 -813 3476
rect -779 3442 -744 3476
rect -710 3442 -675 3476
rect -641 3442 -606 3476
rect -572 3442 -537 3476
rect -503 3442 -468 3476
rect -434 3442 -399 3476
rect -365 3442 -330 3476
rect -296 3442 -261 3476
rect -227 3442 -192 3476
rect -158 3442 -123 3476
rect -89 3442 -54 3476
rect -20 3442 15 3476
rect 49 3442 84 3476
rect 118 3442 153 3476
rect 187 3442 222 3476
rect 256 3442 291 3476
rect 325 3442 360 3476
rect 394 3442 429 3476
rect 463 3442 498 3476
rect 532 3442 567 3476
rect 601 3442 636 3476
rect 670 3442 705 3476
rect 739 3442 774 3476
rect 808 3442 843 3476
rect 877 3442 912 3476
rect 946 3442 981 3476
rect 1015 3442 1050 3476
rect 1084 3442 1119 3476
rect 1153 3442 1188 3476
rect 1222 3442 1257 3476
rect 1291 3442 1326 3476
rect 1360 3442 1395 3476
rect 1429 3442 1464 3476
rect 1498 3442 1533 3476
rect 1567 3442 1602 3476
rect 1636 3442 1671 3476
rect 1705 3442 1740 3476
rect 1774 3442 1809 3476
rect 1843 3442 1878 3476
rect 1912 3442 1947 3476
rect 1981 3442 2016 3476
rect 2050 3442 2085 3476
rect 2119 3442 2154 3476
rect 2188 3442 2223 3476
rect 2257 3442 2292 3476
rect 2326 3442 2361 3476
rect 2395 3442 2430 3476
rect 2464 3442 2499 3476
rect 2533 3442 2568 3476
rect 2602 3442 2637 3476
rect 2671 3442 2706 3476
rect 2740 3442 2775 3476
rect 2809 3442 2844 3476
rect 2878 3442 2913 3476
rect 2947 3442 2982 3476
rect 3016 3442 3051 3476
rect 3085 3442 3120 3476
rect 3154 3442 3189 3476
rect 3223 3442 3258 3476
rect 3292 3442 3327 3476
rect 3361 3442 3396 3476
rect -1088 3408 3396 3442
rect -1088 3374 -1020 3408
rect -986 3374 -951 3408
rect -917 3374 -882 3408
rect -848 3374 -813 3408
rect -779 3374 -744 3408
rect -710 3374 -675 3408
rect -641 3374 -606 3408
rect -572 3374 -537 3408
rect -503 3374 -468 3408
rect -434 3374 -399 3408
rect -365 3374 -330 3408
rect -296 3374 -261 3408
rect -227 3374 -192 3408
rect -158 3374 -123 3408
rect -89 3374 -54 3408
rect -20 3374 15 3408
rect 49 3374 84 3408
rect 118 3374 153 3408
rect 187 3374 222 3408
rect 256 3374 291 3408
rect 325 3374 360 3408
rect 394 3374 429 3408
rect 463 3374 498 3408
rect 532 3374 567 3408
rect 601 3374 636 3408
rect 670 3374 705 3408
rect 739 3374 774 3408
rect 808 3374 843 3408
rect 877 3374 912 3408
rect 946 3374 981 3408
rect 1015 3374 1050 3408
rect 1084 3374 1119 3408
rect 1153 3374 1188 3408
rect 1222 3374 1257 3408
rect 1291 3374 1326 3408
rect 1360 3374 1395 3408
rect 1429 3374 1464 3408
rect 1498 3374 1533 3408
rect 1567 3374 1602 3408
rect 1636 3374 1671 3408
rect 1705 3374 1740 3408
rect 1774 3374 1809 3408
rect 1843 3374 1878 3408
rect 1912 3374 1947 3408
rect 1981 3374 2016 3408
rect 2050 3374 2085 3408
rect 2119 3374 2154 3408
rect 2188 3374 2223 3408
rect 2257 3374 2292 3408
rect 2326 3374 2361 3408
rect 2395 3374 2430 3408
rect 2464 3374 2499 3408
rect 2533 3374 2568 3408
rect 2602 3374 2637 3408
rect 2671 3374 2706 3408
rect 2740 3374 2775 3408
rect 2809 3374 2844 3408
rect 2878 3374 2913 3408
rect 2947 3374 2982 3408
rect 3016 3374 3051 3408
rect 3085 3374 3120 3408
rect 3154 3374 3189 3408
rect 3223 3374 3258 3408
rect 3292 3374 3327 3408
rect 3361 3374 3396 3408
rect 13902 3374 13970 3544
rect -1088 3306 -306 3374
rect 13188 3306 13970 3374
rect -1088 449 -306 484
rect -1054 415 -1020 449
rect -986 415 -952 449
rect -918 415 -884 449
rect -850 415 -816 449
rect -782 415 -748 449
rect -714 415 -680 449
rect -646 415 -612 449
rect -578 415 -544 449
rect -510 415 -476 449
rect -442 415 -408 449
rect -374 415 -340 449
rect -1088 380 -306 415
rect -1054 346 -1020 380
rect -986 346 -952 380
rect -918 346 -884 380
rect -850 346 -816 380
rect -782 346 -748 380
rect -714 346 -680 380
rect -646 346 -612 380
rect -578 346 -544 380
rect -510 346 -476 380
rect -442 346 -408 380
rect -374 346 -340 380
rect -1088 311 -306 346
rect -1054 277 -1020 311
rect -986 277 -952 311
rect -918 277 -884 311
rect -850 277 -816 311
rect -782 277 -748 311
rect -714 277 -680 311
rect -646 277 -612 311
rect -578 277 -544 311
rect -510 277 -476 311
rect -442 277 -408 311
rect -374 277 -340 311
rect -1088 242 -306 277
rect -1054 208 -1020 242
rect -986 208 -952 242
rect -918 208 -884 242
rect -850 208 -816 242
rect -782 208 -748 242
rect -714 208 -680 242
rect -646 208 -612 242
rect -578 208 -544 242
rect -510 208 -476 242
rect -442 208 -408 242
rect -374 208 -340 242
rect -1088 173 -306 208
rect -1054 139 -1020 173
rect -986 139 -952 173
rect -918 139 -884 173
rect -850 139 -816 173
rect -782 139 -748 173
rect -714 139 -680 173
rect -646 139 -612 173
rect -578 139 -544 173
rect -510 139 -476 173
rect -442 139 -408 173
rect -374 139 -340 173
rect -1088 104 -306 139
rect -1054 70 -1020 104
rect -986 70 -952 104
rect -918 70 -884 104
rect -850 70 -816 104
rect -782 70 -748 104
rect -714 70 -680 104
rect -646 70 -612 104
rect -578 70 -544 104
rect -510 70 -476 104
rect -442 70 -408 104
rect -374 70 -340 104
rect -1088 35 -306 70
rect -1054 1 -1020 35
rect -986 1 -952 35
rect -918 1 -884 35
rect -850 1 -816 35
rect -782 1 -748 35
rect -714 1 -680 35
rect -646 1 -612 35
rect -578 1 -544 35
rect -510 1 -476 35
rect -442 1 -408 35
rect -374 1 -340 35
rect -1088 -34 -306 1
rect 13188 449 13970 484
rect 13222 415 13256 449
rect 13290 415 13324 449
rect 13358 415 13392 449
rect 13426 415 13460 449
rect 13494 415 13528 449
rect 13562 415 13596 449
rect 13630 415 13664 449
rect 13698 415 13732 449
rect 13766 415 13800 449
rect 13834 415 13868 449
rect 13902 415 13936 449
rect 13188 380 13970 415
rect 13222 346 13256 380
rect 13290 346 13324 380
rect 13358 346 13392 380
rect 13426 346 13460 380
rect 13494 346 13528 380
rect 13562 346 13596 380
rect 13630 346 13664 380
rect 13698 346 13732 380
rect 13766 346 13800 380
rect 13834 346 13868 380
rect 13902 346 13936 380
rect 13188 311 13970 346
rect 13222 277 13256 311
rect 13290 277 13324 311
rect 13358 277 13392 311
rect 13426 277 13460 311
rect 13494 277 13528 311
rect 13562 277 13596 311
rect 13630 277 13664 311
rect 13698 277 13732 311
rect 13766 277 13800 311
rect 13834 277 13868 311
rect 13902 277 13936 311
rect 13188 242 13970 277
rect 13222 208 13256 242
rect 13290 208 13324 242
rect 13358 208 13392 242
rect 13426 208 13460 242
rect 13494 208 13528 242
rect 13562 208 13596 242
rect 13630 208 13664 242
rect 13698 208 13732 242
rect 13766 208 13800 242
rect 13834 208 13868 242
rect 13902 208 13936 242
rect 13188 173 13970 208
rect 13222 139 13256 173
rect 13290 139 13324 173
rect 13358 139 13392 173
rect 13426 139 13460 173
rect 13494 139 13528 173
rect 13562 139 13596 173
rect 13630 139 13664 173
rect 13698 139 13732 173
rect 13766 139 13800 173
rect 13834 139 13868 173
rect 13902 139 13936 173
rect 13188 104 13970 139
rect 13222 70 13256 104
rect 13290 70 13324 104
rect 13358 70 13392 104
rect 13426 70 13460 104
rect 13494 70 13528 104
rect 13562 70 13596 104
rect 13630 70 13664 104
rect 13698 70 13732 104
rect 13766 70 13800 104
rect 13834 70 13868 104
rect 13902 70 13936 104
rect 13188 35 13970 70
rect 13222 1 13256 35
rect 13290 1 13324 35
rect 13358 1 13392 35
rect 13426 1 13460 35
rect 13494 1 13528 35
rect 13562 1 13596 35
rect 13630 1 13664 35
rect 13698 1 13732 35
rect 13766 1 13800 35
rect 13834 1 13868 35
rect 13902 1 13936 35
rect -1054 -68 -1020 -34
rect -986 -68 -952 -34
rect -918 -68 -884 -34
rect -850 -68 -816 -34
rect -782 -68 -748 -34
rect -714 -68 -680 -34
rect -646 -68 -612 -34
rect -578 -68 -544 -34
rect -510 -68 -476 -34
rect -442 -68 -408 -34
rect -374 -68 -340 -34
rect -1088 -103 -306 -68
rect 13188 -34 13970 1
rect 13222 -68 13256 -34
rect 13290 -68 13324 -34
rect 13358 -68 13392 -34
rect 13426 -68 13460 -34
rect 13494 -68 13528 -34
rect 13562 -68 13596 -34
rect 13630 -68 13664 -34
rect 13698 -68 13732 -34
rect 13766 -68 13800 -34
rect 13834 -68 13868 -34
rect 13902 -68 13936 -34
rect -1054 -137 -1020 -103
rect -986 -137 -952 -103
rect -918 -137 -884 -103
rect -850 -137 -816 -103
rect -782 -137 -748 -103
rect -714 -137 -680 -103
rect -646 -137 -612 -103
rect -578 -137 -544 -103
rect -510 -137 -476 -103
rect -442 -137 -408 -103
rect -374 -137 -340 -103
rect -1088 -172 -306 -137
rect -1054 -206 -1020 -172
rect -986 -206 -952 -172
rect -918 -206 -884 -172
rect -850 -206 -816 -172
rect -782 -206 -748 -172
rect -714 -206 -680 -172
rect -646 -206 -612 -172
rect -578 -206 -544 -172
rect -510 -206 -476 -172
rect -442 -206 -408 -172
rect -374 -206 -340 -172
rect -1088 -274 -306 -206
rect 13188 -103 13970 -68
rect 13222 -137 13256 -103
rect 13290 -137 13324 -103
rect 13358 -137 13392 -103
rect 13426 -137 13460 -103
rect 13494 -137 13528 -103
rect 13562 -137 13596 -103
rect 13630 -137 13664 -103
rect 13698 -137 13732 -103
rect 13766 -137 13800 -103
rect 13834 -137 13868 -103
rect 13902 -137 13936 -103
rect 13188 -172 13970 -137
rect 13222 -206 13256 -172
rect 13290 -206 13324 -172
rect 13358 -206 13392 -172
rect 13426 -206 13460 -172
rect 13494 -206 13528 -172
rect 13562 -206 13596 -172
rect 13630 -206 13664 -172
rect 13698 -206 13732 -172
rect 13766 -206 13800 -172
rect 13834 -206 13868 -172
rect 13902 -206 13936 -172
rect 13188 -274 13970 -206
rect -1088 -308 -1020 -274
rect -986 -308 -951 -274
rect -917 -308 -882 -274
rect -848 -308 -813 -274
rect -779 -308 -744 -274
rect -710 -308 -675 -274
rect -641 -308 -606 -274
rect -572 -308 -537 -274
rect -503 -308 -468 -274
rect -434 -308 -399 -274
rect -365 -308 -330 -274
rect -296 -308 -261 -274
rect -227 -308 -192 -274
rect -158 -308 -123 -274
rect -89 -308 -54 -274
rect -20 -308 15 -274
rect 49 -308 84 -274
rect 118 -308 153 -274
rect 187 -308 222 -274
rect 256 -308 291 -274
rect 325 -308 360 -274
rect 394 -308 429 -274
rect 463 -308 498 -274
rect 532 -308 567 -274
rect 601 -308 636 -274
rect 670 -308 705 -274
rect 739 -308 774 -274
rect 808 -308 843 -274
rect 877 -308 912 -274
rect 946 -308 981 -274
rect 1015 -308 1050 -274
rect 1084 -308 1119 -274
rect 1153 -308 1188 -274
rect 1222 -308 1257 -274
rect 1291 -308 1326 -274
rect 1360 -308 1395 -274
rect 1429 -308 1464 -274
rect 1498 -308 1533 -274
rect 1567 -308 1602 -274
rect 1636 -308 1671 -274
rect 1705 -308 1740 -274
rect 1774 -308 1809 -274
rect 1843 -308 1878 -274
rect 1912 -308 1947 -274
rect 1981 -308 2016 -274
rect 2050 -308 2085 -274
rect 2119 -308 2154 -274
rect 2188 -308 2223 -274
rect 2257 -308 2292 -274
rect 2326 -308 2361 -274
rect 2395 -308 2430 -274
rect 2464 -308 2499 -274
rect 2533 -308 2568 -274
rect 2602 -308 2637 -274
rect 2671 -308 2706 -274
rect 2740 -308 2775 -274
rect 2809 -308 2844 -274
rect 2878 -308 2913 -274
rect 2947 -308 2982 -274
rect 3016 -308 3051 -274
rect 3085 -308 3120 -274
rect 3154 -308 3189 -274
rect 3223 -308 3258 -274
rect 3292 -308 3327 -274
rect 3361 -308 3396 -274
rect -1088 -342 3396 -308
rect -1088 -376 -1020 -342
rect -986 -376 -951 -342
rect -917 -376 -882 -342
rect -848 -376 -813 -342
rect -779 -376 -744 -342
rect -710 -376 -675 -342
rect -641 -376 -606 -342
rect -572 -376 -537 -342
rect -503 -376 -468 -342
rect -434 -376 -399 -342
rect -365 -376 -330 -342
rect -296 -376 -261 -342
rect -227 -376 -192 -342
rect -158 -376 -123 -342
rect -89 -376 -54 -342
rect -20 -376 15 -342
rect 49 -376 84 -342
rect 118 -376 153 -342
rect 187 -376 222 -342
rect 256 -376 291 -342
rect 325 -376 360 -342
rect 394 -376 429 -342
rect 463 -376 498 -342
rect 532 -376 567 -342
rect 601 -376 636 -342
rect 670 -376 705 -342
rect 739 -376 774 -342
rect 808 -376 843 -342
rect 877 -376 912 -342
rect 946 -376 981 -342
rect 1015 -376 1050 -342
rect 1084 -376 1119 -342
rect 1153 -376 1188 -342
rect 1222 -376 1257 -342
rect 1291 -376 1326 -342
rect 1360 -376 1395 -342
rect 1429 -376 1464 -342
rect 1498 -376 1533 -342
rect 1567 -376 1602 -342
rect 1636 -376 1671 -342
rect 1705 -376 1740 -342
rect 1774 -376 1809 -342
rect 1843 -376 1878 -342
rect 1912 -376 1947 -342
rect 1981 -376 2016 -342
rect 2050 -376 2085 -342
rect 2119 -376 2154 -342
rect 2188 -376 2223 -342
rect 2257 -376 2292 -342
rect 2326 -376 2361 -342
rect 2395 -376 2430 -342
rect 2464 -376 2499 -342
rect 2533 -376 2568 -342
rect 2602 -376 2637 -342
rect 2671 -376 2706 -342
rect 2740 -376 2775 -342
rect 2809 -376 2844 -342
rect 2878 -376 2913 -342
rect 2947 -376 2982 -342
rect 3016 -376 3051 -342
rect 3085 -376 3120 -342
rect 3154 -376 3189 -342
rect 3223 -376 3258 -342
rect 3292 -376 3327 -342
rect 3361 -376 3396 -342
rect -1088 -410 3396 -376
rect -1088 -444 -1020 -410
rect -986 -444 -951 -410
rect -917 -444 -882 -410
rect -848 -444 -813 -410
rect -779 -444 -744 -410
rect -710 -444 -675 -410
rect -641 -444 -606 -410
rect -572 -444 -537 -410
rect -503 -444 -468 -410
rect -434 -444 -399 -410
rect -365 -444 -330 -410
rect -296 -444 -261 -410
rect -227 -444 -192 -410
rect -158 -444 -123 -410
rect -89 -444 -54 -410
rect -20 -444 15 -410
rect 49 -444 84 -410
rect 118 -444 153 -410
rect 187 -444 222 -410
rect 256 -444 291 -410
rect 325 -444 360 -410
rect 394 -444 429 -410
rect 463 -444 498 -410
rect 532 -444 567 -410
rect 601 -444 636 -410
rect 670 -444 705 -410
rect 739 -444 774 -410
rect 808 -444 843 -410
rect 877 -444 912 -410
rect 946 -444 981 -410
rect 1015 -444 1050 -410
rect 1084 -444 1119 -410
rect 1153 -444 1188 -410
rect 1222 -444 1257 -410
rect 1291 -444 1326 -410
rect 1360 -444 1395 -410
rect 1429 -444 1464 -410
rect 1498 -444 1533 -410
rect 1567 -444 1602 -410
rect 1636 -444 1671 -410
rect 1705 -444 1740 -410
rect 1774 -444 1809 -410
rect 1843 -444 1878 -410
rect 1912 -444 1947 -410
rect 1981 -444 2016 -410
rect 2050 -444 2085 -410
rect 2119 -444 2154 -410
rect 2188 -444 2223 -410
rect 2257 -444 2292 -410
rect 2326 -444 2361 -410
rect 2395 -444 2430 -410
rect 2464 -444 2499 -410
rect 2533 -444 2568 -410
rect 2602 -444 2637 -410
rect 2671 -444 2706 -410
rect 2740 -444 2775 -410
rect 2809 -444 2844 -410
rect 2878 -444 2913 -410
rect 2947 -444 2982 -410
rect 3016 -444 3051 -410
rect 3085 -444 3120 -410
rect 3154 -444 3189 -410
rect 3223 -444 3258 -410
rect 3292 -444 3327 -410
rect 3361 -444 3396 -410
rect 13902 -444 13970 -274
<< mvpsubdiffcont >>
rect -1390 3880 -1356 3914
rect -1321 3880 -1287 3914
rect -1252 3880 -1218 3914
rect -1183 3880 -1149 3914
rect -1114 3880 -1080 3914
rect -1045 3880 -1011 3914
rect -976 3880 -942 3914
rect -907 3880 -873 3914
rect -838 3880 -804 3914
rect -769 3880 -735 3914
rect -700 3880 -666 3914
rect -631 3880 -597 3914
rect -562 3880 -528 3914
rect -493 3880 -459 3914
rect -424 3880 -390 3914
rect -355 3880 -321 3914
rect -286 3880 -252 3914
rect -217 3880 -183 3914
rect -148 3880 -114 3914
rect -79 3880 -45 3914
rect -10 3880 24 3914
rect 59 3880 93 3914
rect 128 3880 162 3914
rect 197 3880 231 3914
rect 266 3880 300 3914
rect 335 3880 369 3914
rect 404 3880 438 3914
rect 473 3880 507 3914
rect 542 3880 576 3914
rect 611 3880 645 3914
rect 680 3880 714 3914
rect 749 3880 783 3914
rect 818 3880 852 3914
rect 887 3880 921 3914
rect 956 3880 990 3914
rect 1025 3880 1059 3914
rect 1094 3880 1128 3914
rect 1163 3880 1197 3914
rect 1232 3880 1266 3914
rect 1301 3880 1335 3914
rect 1370 3880 1404 3914
rect 1439 3880 1473 3914
rect 1508 3880 1542 3914
rect 1577 3880 1611 3914
rect 1646 3880 1680 3914
rect 1715 3880 1749 3914
rect 1784 3880 1818 3914
rect 1853 3880 1887 3914
rect 1922 3880 1956 3914
rect 1991 3880 2025 3914
rect 2060 3880 2094 3914
rect 2129 3880 2163 3914
rect 2198 3880 2232 3914
rect 2267 3880 2301 3914
rect 2336 3880 2370 3914
rect 2405 3880 2439 3914
rect -1390 3812 -1356 3846
rect -1321 3812 -1287 3846
rect -1252 3812 -1218 3846
rect -1183 3812 -1149 3846
rect -1114 3812 -1080 3846
rect -1045 3812 -1011 3846
rect -976 3812 -942 3846
rect -907 3812 -873 3846
rect -838 3812 -804 3846
rect -769 3812 -735 3846
rect -700 3812 -666 3846
rect -631 3812 -597 3846
rect -562 3812 -528 3846
rect -493 3812 -459 3846
rect -424 3812 -390 3846
rect -355 3812 -321 3846
rect -286 3812 -252 3846
rect -217 3812 -183 3846
rect -148 3812 -114 3846
rect -79 3812 -45 3846
rect -10 3812 24 3846
rect 59 3812 93 3846
rect 128 3812 162 3846
rect 197 3812 231 3846
rect 266 3812 300 3846
rect 335 3812 369 3846
rect 404 3812 438 3846
rect 473 3812 507 3846
rect 542 3812 576 3846
rect 611 3812 645 3846
rect 680 3812 714 3846
rect 749 3812 783 3846
rect 818 3812 852 3846
rect 887 3812 921 3846
rect 956 3812 990 3846
rect 1025 3812 1059 3846
rect 1094 3812 1128 3846
rect 1163 3812 1197 3846
rect 1232 3812 1266 3846
rect 1301 3812 1335 3846
rect 1370 3812 1404 3846
rect 1439 3812 1473 3846
rect 1508 3812 1542 3846
rect 1577 3812 1611 3846
rect 1646 3812 1680 3846
rect 1715 3812 1749 3846
rect 1784 3812 1818 3846
rect 1853 3812 1887 3846
rect 1922 3812 1956 3846
rect 1991 3812 2025 3846
rect 2060 3812 2094 3846
rect 2129 3812 2163 3846
rect 2198 3812 2232 3846
rect 2267 3812 2301 3846
rect 2336 3812 2370 3846
rect 2405 3812 2439 3846
rect -1390 3744 -1356 3778
rect -1321 3744 -1287 3778
rect -1252 3744 -1218 3778
rect -1183 3744 -1149 3778
rect -1114 3744 -1080 3778
rect -1045 3744 -1011 3778
rect -976 3744 -942 3778
rect -907 3744 -873 3778
rect -838 3744 -804 3778
rect -769 3744 -735 3778
rect -700 3744 -666 3778
rect -631 3744 -597 3778
rect -562 3744 -528 3778
rect -493 3744 -459 3778
rect -424 3744 -390 3778
rect -355 3744 -321 3778
rect -286 3744 -252 3778
rect -217 3744 -183 3778
rect -148 3744 -114 3778
rect -79 3744 -45 3778
rect -10 3744 24 3778
rect 59 3744 93 3778
rect 128 3744 162 3778
rect 197 3744 231 3778
rect 266 3744 300 3778
rect 335 3744 369 3778
rect 404 3744 438 3778
rect 473 3744 507 3778
rect 542 3744 576 3778
rect 611 3744 645 3778
rect 680 3744 714 3778
rect 749 3744 783 3778
rect 818 3744 852 3778
rect 887 3744 921 3778
rect 956 3744 990 3778
rect 1025 3744 1059 3778
rect 1094 3744 1128 3778
rect 1163 3744 1197 3778
rect 1232 3744 1266 3778
rect 1301 3744 1335 3778
rect 1370 3744 1404 3778
rect 1439 3744 1473 3778
rect 1508 3744 1542 3778
rect 1577 3744 1611 3778
rect 1646 3744 1680 3778
rect 1715 3744 1749 3778
rect 1784 3744 1818 3778
rect 1853 3744 1887 3778
rect 1922 3744 1956 3778
rect 1991 3744 2025 3778
rect 2060 3744 2094 3778
rect 2129 3744 2163 3778
rect 2198 3744 2232 3778
rect 2267 3744 2301 3778
rect 2336 3744 2370 3778
rect 2405 3744 2439 3778
rect 2474 3744 14272 3914
rect -1458 -438 -1288 3676
rect 14170 -438 14340 3676
rect -1458 -507 -1424 -473
rect -1390 -507 -1356 -473
rect -1322 -507 -1288 -473
rect -1458 -576 -1424 -542
rect -1390 -576 -1356 -542
rect -1322 -576 -1288 -542
rect 14170 -507 14204 -473
rect 14238 -507 14272 -473
rect 14306 -507 14340 -473
rect 14170 -576 14204 -542
rect 14238 -576 14272 -542
rect 14306 -576 14340 -542
rect -1390 -678 -1356 -644
rect -1321 -678 -1287 -644
rect -1252 -678 -1218 -644
rect -1183 -678 -1149 -644
rect -1114 -678 -1080 -644
rect -1045 -678 -1011 -644
rect -976 -678 -942 -644
rect -907 -678 -873 -644
rect -838 -678 -804 -644
rect -769 -678 -735 -644
rect -700 -678 -666 -644
rect -631 -678 -597 -644
rect -562 -678 -528 -644
rect -493 -678 -459 -644
rect -424 -678 -390 -644
rect -355 -678 -321 -644
rect -286 -678 -252 -644
rect -217 -678 -183 -644
rect -148 -678 -114 -644
rect -79 -678 -45 -644
rect -10 -678 24 -644
rect 59 -678 93 -644
rect 128 -678 162 -644
rect 197 -678 231 -644
rect 266 -678 300 -644
rect 335 -678 369 -644
rect 404 -678 438 -644
rect 473 -678 507 -644
rect 542 -678 576 -644
rect 611 -678 645 -644
rect 680 -678 714 -644
rect 749 -678 783 -644
rect 818 -678 852 -644
rect 887 -678 921 -644
rect 956 -678 990 -644
rect 1025 -678 1059 -644
rect 1094 -678 1128 -644
rect 1163 -678 1197 -644
rect 1232 -678 1266 -644
rect 1301 -678 1335 -644
rect 1370 -678 1404 -644
rect 1439 -678 1473 -644
rect 1508 -678 1542 -644
rect 1577 -678 1611 -644
rect 1646 -678 1680 -644
rect 1715 -678 1749 -644
rect 1784 -678 1818 -644
rect 1853 -678 1887 -644
rect 1922 -678 1956 -644
rect 1991 -678 2025 -644
rect 2060 -678 2094 -644
rect 2129 -678 2163 -644
rect 2198 -678 2232 -644
rect 2267 -678 2301 -644
rect 2336 -678 2370 -644
rect 2405 -678 2439 -644
rect -1390 -746 -1356 -712
rect -1321 -746 -1287 -712
rect -1252 -746 -1218 -712
rect -1183 -746 -1149 -712
rect -1114 -746 -1080 -712
rect -1045 -746 -1011 -712
rect -976 -746 -942 -712
rect -907 -746 -873 -712
rect -838 -746 -804 -712
rect -769 -746 -735 -712
rect -700 -746 -666 -712
rect -631 -746 -597 -712
rect -562 -746 -528 -712
rect -493 -746 -459 -712
rect -424 -746 -390 -712
rect -355 -746 -321 -712
rect -286 -746 -252 -712
rect -217 -746 -183 -712
rect -148 -746 -114 -712
rect -79 -746 -45 -712
rect -10 -746 24 -712
rect 59 -746 93 -712
rect 128 -746 162 -712
rect 197 -746 231 -712
rect 266 -746 300 -712
rect 335 -746 369 -712
rect 404 -746 438 -712
rect 473 -746 507 -712
rect 542 -746 576 -712
rect 611 -746 645 -712
rect 680 -746 714 -712
rect 749 -746 783 -712
rect 818 -746 852 -712
rect 887 -746 921 -712
rect 956 -746 990 -712
rect 1025 -746 1059 -712
rect 1094 -746 1128 -712
rect 1163 -746 1197 -712
rect 1232 -746 1266 -712
rect 1301 -746 1335 -712
rect 1370 -746 1404 -712
rect 1439 -746 1473 -712
rect 1508 -746 1542 -712
rect 1577 -746 1611 -712
rect 1646 -746 1680 -712
rect 1715 -746 1749 -712
rect 1784 -746 1818 -712
rect 1853 -746 1887 -712
rect 1922 -746 1956 -712
rect 1991 -746 2025 -712
rect 2060 -746 2094 -712
rect 2129 -746 2163 -712
rect 2198 -746 2232 -712
rect 2267 -746 2301 -712
rect 2336 -746 2370 -712
rect 2405 -746 2439 -712
rect -1390 -814 -1356 -780
rect -1321 -814 -1287 -780
rect -1252 -814 -1218 -780
rect -1183 -814 -1149 -780
rect -1114 -814 -1080 -780
rect -1045 -814 -1011 -780
rect -976 -814 -942 -780
rect -907 -814 -873 -780
rect -838 -814 -804 -780
rect -769 -814 -735 -780
rect -700 -814 -666 -780
rect -631 -814 -597 -780
rect -562 -814 -528 -780
rect -493 -814 -459 -780
rect -424 -814 -390 -780
rect -355 -814 -321 -780
rect -286 -814 -252 -780
rect -217 -814 -183 -780
rect -148 -814 -114 -780
rect -79 -814 -45 -780
rect -10 -814 24 -780
rect 59 -814 93 -780
rect 128 -814 162 -780
rect 197 -814 231 -780
rect 266 -814 300 -780
rect 335 -814 369 -780
rect 404 -814 438 -780
rect 473 -814 507 -780
rect 542 -814 576 -780
rect 611 -814 645 -780
rect 680 -814 714 -780
rect 749 -814 783 -780
rect 818 -814 852 -780
rect 887 -814 921 -780
rect 956 -814 990 -780
rect 1025 -814 1059 -780
rect 1094 -814 1128 -780
rect 1163 -814 1197 -780
rect 1232 -814 1266 -780
rect 1301 -814 1335 -780
rect 1370 -814 1404 -780
rect 1439 -814 1473 -780
rect 1508 -814 1542 -780
rect 1577 -814 1611 -780
rect 1646 -814 1680 -780
rect 1715 -814 1749 -780
rect 1784 -814 1818 -780
rect 1853 -814 1887 -780
rect 1922 -814 1956 -780
rect 1991 -814 2025 -780
rect 2060 -814 2094 -780
rect 2129 -814 2163 -780
rect 2198 -814 2232 -780
rect 2267 -814 2301 -780
rect 2336 -814 2370 -780
rect 2405 -814 2439 -780
rect 2474 -814 14272 -644
<< mvnsubdiffcont >>
rect -1020 3510 -986 3544
rect -951 3510 -917 3544
rect -882 3510 -848 3544
rect -813 3510 -779 3544
rect -744 3510 -710 3544
rect -675 3510 -641 3544
rect -606 3510 -572 3544
rect -537 3510 -503 3544
rect -468 3510 -434 3544
rect -399 3510 -365 3544
rect -330 3510 -296 3544
rect -261 3510 -227 3544
rect -192 3510 -158 3544
rect -123 3510 -89 3544
rect -54 3510 -20 3544
rect 15 3510 49 3544
rect 84 3510 118 3544
rect 153 3510 187 3544
rect 222 3510 256 3544
rect 291 3510 325 3544
rect 360 3510 394 3544
rect 429 3510 463 3544
rect 498 3510 532 3544
rect 567 3510 601 3544
rect 636 3510 670 3544
rect 705 3510 739 3544
rect 774 3510 808 3544
rect 843 3510 877 3544
rect 912 3510 946 3544
rect 981 3510 1015 3544
rect 1050 3510 1084 3544
rect 1119 3510 1153 3544
rect 1188 3510 1222 3544
rect 1257 3510 1291 3544
rect 1326 3510 1360 3544
rect 1395 3510 1429 3544
rect 1464 3510 1498 3544
rect 1533 3510 1567 3544
rect 1602 3510 1636 3544
rect 1671 3510 1705 3544
rect 1740 3510 1774 3544
rect 1809 3510 1843 3544
rect 1878 3510 1912 3544
rect 1947 3510 1981 3544
rect 2016 3510 2050 3544
rect 2085 3510 2119 3544
rect 2154 3510 2188 3544
rect 2223 3510 2257 3544
rect 2292 3510 2326 3544
rect 2361 3510 2395 3544
rect 2430 3510 2464 3544
rect 2499 3510 2533 3544
rect 2568 3510 2602 3544
rect 2637 3510 2671 3544
rect 2706 3510 2740 3544
rect 2775 3510 2809 3544
rect 2844 3510 2878 3544
rect 2913 3510 2947 3544
rect 2982 3510 3016 3544
rect 3051 3510 3085 3544
rect 3120 3510 3154 3544
rect 3189 3510 3223 3544
rect 3258 3510 3292 3544
rect 3327 3510 3361 3544
rect -1020 3442 -986 3476
rect -951 3442 -917 3476
rect -882 3442 -848 3476
rect -813 3442 -779 3476
rect -744 3442 -710 3476
rect -675 3442 -641 3476
rect -606 3442 -572 3476
rect -537 3442 -503 3476
rect -468 3442 -434 3476
rect -399 3442 -365 3476
rect -330 3442 -296 3476
rect -261 3442 -227 3476
rect -192 3442 -158 3476
rect -123 3442 -89 3476
rect -54 3442 -20 3476
rect 15 3442 49 3476
rect 84 3442 118 3476
rect 153 3442 187 3476
rect 222 3442 256 3476
rect 291 3442 325 3476
rect 360 3442 394 3476
rect 429 3442 463 3476
rect 498 3442 532 3476
rect 567 3442 601 3476
rect 636 3442 670 3476
rect 705 3442 739 3476
rect 774 3442 808 3476
rect 843 3442 877 3476
rect 912 3442 946 3476
rect 981 3442 1015 3476
rect 1050 3442 1084 3476
rect 1119 3442 1153 3476
rect 1188 3442 1222 3476
rect 1257 3442 1291 3476
rect 1326 3442 1360 3476
rect 1395 3442 1429 3476
rect 1464 3442 1498 3476
rect 1533 3442 1567 3476
rect 1602 3442 1636 3476
rect 1671 3442 1705 3476
rect 1740 3442 1774 3476
rect 1809 3442 1843 3476
rect 1878 3442 1912 3476
rect 1947 3442 1981 3476
rect 2016 3442 2050 3476
rect 2085 3442 2119 3476
rect 2154 3442 2188 3476
rect 2223 3442 2257 3476
rect 2292 3442 2326 3476
rect 2361 3442 2395 3476
rect 2430 3442 2464 3476
rect 2499 3442 2533 3476
rect 2568 3442 2602 3476
rect 2637 3442 2671 3476
rect 2706 3442 2740 3476
rect 2775 3442 2809 3476
rect 2844 3442 2878 3476
rect 2913 3442 2947 3476
rect 2982 3442 3016 3476
rect 3051 3442 3085 3476
rect 3120 3442 3154 3476
rect 3189 3442 3223 3476
rect 3258 3442 3292 3476
rect 3327 3442 3361 3476
rect -1020 3374 -986 3408
rect -951 3374 -917 3408
rect -882 3374 -848 3408
rect -813 3374 -779 3408
rect -744 3374 -710 3408
rect -675 3374 -641 3408
rect -606 3374 -572 3408
rect -537 3374 -503 3408
rect -468 3374 -434 3408
rect -399 3374 -365 3408
rect -330 3374 -296 3408
rect -261 3374 -227 3408
rect -192 3374 -158 3408
rect -123 3374 -89 3408
rect -54 3374 -20 3408
rect 15 3374 49 3408
rect 84 3374 118 3408
rect 153 3374 187 3408
rect 222 3374 256 3408
rect 291 3374 325 3408
rect 360 3374 394 3408
rect 429 3374 463 3408
rect 498 3374 532 3408
rect 567 3374 601 3408
rect 636 3374 670 3408
rect 705 3374 739 3408
rect 774 3374 808 3408
rect 843 3374 877 3408
rect 912 3374 946 3408
rect 981 3374 1015 3408
rect 1050 3374 1084 3408
rect 1119 3374 1153 3408
rect 1188 3374 1222 3408
rect 1257 3374 1291 3408
rect 1326 3374 1360 3408
rect 1395 3374 1429 3408
rect 1464 3374 1498 3408
rect 1533 3374 1567 3408
rect 1602 3374 1636 3408
rect 1671 3374 1705 3408
rect 1740 3374 1774 3408
rect 1809 3374 1843 3408
rect 1878 3374 1912 3408
rect 1947 3374 1981 3408
rect 2016 3374 2050 3408
rect 2085 3374 2119 3408
rect 2154 3374 2188 3408
rect 2223 3374 2257 3408
rect 2292 3374 2326 3408
rect 2361 3374 2395 3408
rect 2430 3374 2464 3408
rect 2499 3374 2533 3408
rect 2568 3374 2602 3408
rect 2637 3374 2671 3408
rect 2706 3374 2740 3408
rect 2775 3374 2809 3408
rect 2844 3374 2878 3408
rect 2913 3374 2947 3408
rect 2982 3374 3016 3408
rect 3051 3374 3085 3408
rect 3120 3374 3154 3408
rect 3189 3374 3223 3408
rect 3258 3374 3292 3408
rect 3327 3374 3361 3408
rect 3396 3374 13902 3544
rect -1088 484 -306 3306
rect -1088 415 -1054 449
rect -1020 415 -986 449
rect -952 415 -918 449
rect -884 415 -850 449
rect -816 415 -782 449
rect -748 415 -714 449
rect -680 415 -646 449
rect -612 415 -578 449
rect -544 415 -510 449
rect -476 415 -442 449
rect -408 415 -374 449
rect -340 415 -306 449
rect -1088 346 -1054 380
rect -1020 346 -986 380
rect -952 346 -918 380
rect -884 346 -850 380
rect -816 346 -782 380
rect -748 346 -714 380
rect -680 346 -646 380
rect -612 346 -578 380
rect -544 346 -510 380
rect -476 346 -442 380
rect -408 346 -374 380
rect -340 346 -306 380
rect -1088 277 -1054 311
rect -1020 277 -986 311
rect -952 277 -918 311
rect -884 277 -850 311
rect -816 277 -782 311
rect -748 277 -714 311
rect -680 277 -646 311
rect -612 277 -578 311
rect -544 277 -510 311
rect -476 277 -442 311
rect -408 277 -374 311
rect -340 277 -306 311
rect -1088 208 -1054 242
rect -1020 208 -986 242
rect -952 208 -918 242
rect -884 208 -850 242
rect -816 208 -782 242
rect -748 208 -714 242
rect -680 208 -646 242
rect -612 208 -578 242
rect -544 208 -510 242
rect -476 208 -442 242
rect -408 208 -374 242
rect -340 208 -306 242
rect -1088 139 -1054 173
rect -1020 139 -986 173
rect -952 139 -918 173
rect -884 139 -850 173
rect -816 139 -782 173
rect -748 139 -714 173
rect -680 139 -646 173
rect -612 139 -578 173
rect -544 139 -510 173
rect -476 139 -442 173
rect -408 139 -374 173
rect -340 139 -306 173
rect -1088 70 -1054 104
rect -1020 70 -986 104
rect -952 70 -918 104
rect -884 70 -850 104
rect -816 70 -782 104
rect -748 70 -714 104
rect -680 70 -646 104
rect -612 70 -578 104
rect -544 70 -510 104
rect -476 70 -442 104
rect -408 70 -374 104
rect -340 70 -306 104
rect -1088 1 -1054 35
rect -1020 1 -986 35
rect -952 1 -918 35
rect -884 1 -850 35
rect -816 1 -782 35
rect -748 1 -714 35
rect -680 1 -646 35
rect -612 1 -578 35
rect -544 1 -510 35
rect -476 1 -442 35
rect -408 1 -374 35
rect -340 1 -306 35
rect 13188 484 13970 3306
rect 13188 415 13222 449
rect 13256 415 13290 449
rect 13324 415 13358 449
rect 13392 415 13426 449
rect 13460 415 13494 449
rect 13528 415 13562 449
rect 13596 415 13630 449
rect 13664 415 13698 449
rect 13732 415 13766 449
rect 13800 415 13834 449
rect 13868 415 13902 449
rect 13936 415 13970 449
rect 13188 346 13222 380
rect 13256 346 13290 380
rect 13324 346 13358 380
rect 13392 346 13426 380
rect 13460 346 13494 380
rect 13528 346 13562 380
rect 13596 346 13630 380
rect 13664 346 13698 380
rect 13732 346 13766 380
rect 13800 346 13834 380
rect 13868 346 13902 380
rect 13936 346 13970 380
rect 13188 277 13222 311
rect 13256 277 13290 311
rect 13324 277 13358 311
rect 13392 277 13426 311
rect 13460 277 13494 311
rect 13528 277 13562 311
rect 13596 277 13630 311
rect 13664 277 13698 311
rect 13732 277 13766 311
rect 13800 277 13834 311
rect 13868 277 13902 311
rect 13936 277 13970 311
rect 13188 208 13222 242
rect 13256 208 13290 242
rect 13324 208 13358 242
rect 13392 208 13426 242
rect 13460 208 13494 242
rect 13528 208 13562 242
rect 13596 208 13630 242
rect 13664 208 13698 242
rect 13732 208 13766 242
rect 13800 208 13834 242
rect 13868 208 13902 242
rect 13936 208 13970 242
rect 13188 139 13222 173
rect 13256 139 13290 173
rect 13324 139 13358 173
rect 13392 139 13426 173
rect 13460 139 13494 173
rect 13528 139 13562 173
rect 13596 139 13630 173
rect 13664 139 13698 173
rect 13732 139 13766 173
rect 13800 139 13834 173
rect 13868 139 13902 173
rect 13936 139 13970 173
rect 13188 70 13222 104
rect 13256 70 13290 104
rect 13324 70 13358 104
rect 13392 70 13426 104
rect 13460 70 13494 104
rect 13528 70 13562 104
rect 13596 70 13630 104
rect 13664 70 13698 104
rect 13732 70 13766 104
rect 13800 70 13834 104
rect 13868 70 13902 104
rect 13936 70 13970 104
rect 13188 1 13222 35
rect 13256 1 13290 35
rect 13324 1 13358 35
rect 13392 1 13426 35
rect 13460 1 13494 35
rect 13528 1 13562 35
rect 13596 1 13630 35
rect 13664 1 13698 35
rect 13732 1 13766 35
rect 13800 1 13834 35
rect 13868 1 13902 35
rect 13936 1 13970 35
rect -1088 -68 -1054 -34
rect -1020 -68 -986 -34
rect -952 -68 -918 -34
rect -884 -68 -850 -34
rect -816 -68 -782 -34
rect -748 -68 -714 -34
rect -680 -68 -646 -34
rect -612 -68 -578 -34
rect -544 -68 -510 -34
rect -476 -68 -442 -34
rect -408 -68 -374 -34
rect -340 -68 -306 -34
rect 13188 -68 13222 -34
rect 13256 -68 13290 -34
rect 13324 -68 13358 -34
rect 13392 -68 13426 -34
rect 13460 -68 13494 -34
rect 13528 -68 13562 -34
rect 13596 -68 13630 -34
rect 13664 -68 13698 -34
rect 13732 -68 13766 -34
rect 13800 -68 13834 -34
rect 13868 -68 13902 -34
rect 13936 -68 13970 -34
rect -1088 -137 -1054 -103
rect -1020 -137 -986 -103
rect -952 -137 -918 -103
rect -884 -137 -850 -103
rect -816 -137 -782 -103
rect -748 -137 -714 -103
rect -680 -137 -646 -103
rect -612 -137 -578 -103
rect -544 -137 -510 -103
rect -476 -137 -442 -103
rect -408 -137 -374 -103
rect -340 -137 -306 -103
rect -1088 -206 -1054 -172
rect -1020 -206 -986 -172
rect -952 -206 -918 -172
rect -884 -206 -850 -172
rect -816 -206 -782 -172
rect -748 -206 -714 -172
rect -680 -206 -646 -172
rect -612 -206 -578 -172
rect -544 -206 -510 -172
rect -476 -206 -442 -172
rect -408 -206 -374 -172
rect -340 -206 -306 -172
rect 13188 -137 13222 -103
rect 13256 -137 13290 -103
rect 13324 -137 13358 -103
rect 13392 -137 13426 -103
rect 13460 -137 13494 -103
rect 13528 -137 13562 -103
rect 13596 -137 13630 -103
rect 13664 -137 13698 -103
rect 13732 -137 13766 -103
rect 13800 -137 13834 -103
rect 13868 -137 13902 -103
rect 13936 -137 13970 -103
rect 13188 -206 13222 -172
rect 13256 -206 13290 -172
rect 13324 -206 13358 -172
rect 13392 -206 13426 -172
rect 13460 -206 13494 -172
rect 13528 -206 13562 -172
rect 13596 -206 13630 -172
rect 13664 -206 13698 -172
rect 13732 -206 13766 -172
rect 13800 -206 13834 -172
rect 13868 -206 13902 -172
rect 13936 -206 13970 -172
rect -1020 -308 -986 -274
rect -951 -308 -917 -274
rect -882 -308 -848 -274
rect -813 -308 -779 -274
rect -744 -308 -710 -274
rect -675 -308 -641 -274
rect -606 -308 -572 -274
rect -537 -308 -503 -274
rect -468 -308 -434 -274
rect -399 -308 -365 -274
rect -330 -308 -296 -274
rect -261 -308 -227 -274
rect -192 -308 -158 -274
rect -123 -308 -89 -274
rect -54 -308 -20 -274
rect 15 -308 49 -274
rect 84 -308 118 -274
rect 153 -308 187 -274
rect 222 -308 256 -274
rect 291 -308 325 -274
rect 360 -308 394 -274
rect 429 -308 463 -274
rect 498 -308 532 -274
rect 567 -308 601 -274
rect 636 -308 670 -274
rect 705 -308 739 -274
rect 774 -308 808 -274
rect 843 -308 877 -274
rect 912 -308 946 -274
rect 981 -308 1015 -274
rect 1050 -308 1084 -274
rect 1119 -308 1153 -274
rect 1188 -308 1222 -274
rect 1257 -308 1291 -274
rect 1326 -308 1360 -274
rect 1395 -308 1429 -274
rect 1464 -308 1498 -274
rect 1533 -308 1567 -274
rect 1602 -308 1636 -274
rect 1671 -308 1705 -274
rect 1740 -308 1774 -274
rect 1809 -308 1843 -274
rect 1878 -308 1912 -274
rect 1947 -308 1981 -274
rect 2016 -308 2050 -274
rect 2085 -308 2119 -274
rect 2154 -308 2188 -274
rect 2223 -308 2257 -274
rect 2292 -308 2326 -274
rect 2361 -308 2395 -274
rect 2430 -308 2464 -274
rect 2499 -308 2533 -274
rect 2568 -308 2602 -274
rect 2637 -308 2671 -274
rect 2706 -308 2740 -274
rect 2775 -308 2809 -274
rect 2844 -308 2878 -274
rect 2913 -308 2947 -274
rect 2982 -308 3016 -274
rect 3051 -308 3085 -274
rect 3120 -308 3154 -274
rect 3189 -308 3223 -274
rect 3258 -308 3292 -274
rect 3327 -308 3361 -274
rect -1020 -376 -986 -342
rect -951 -376 -917 -342
rect -882 -376 -848 -342
rect -813 -376 -779 -342
rect -744 -376 -710 -342
rect -675 -376 -641 -342
rect -606 -376 -572 -342
rect -537 -376 -503 -342
rect -468 -376 -434 -342
rect -399 -376 -365 -342
rect -330 -376 -296 -342
rect -261 -376 -227 -342
rect -192 -376 -158 -342
rect -123 -376 -89 -342
rect -54 -376 -20 -342
rect 15 -376 49 -342
rect 84 -376 118 -342
rect 153 -376 187 -342
rect 222 -376 256 -342
rect 291 -376 325 -342
rect 360 -376 394 -342
rect 429 -376 463 -342
rect 498 -376 532 -342
rect 567 -376 601 -342
rect 636 -376 670 -342
rect 705 -376 739 -342
rect 774 -376 808 -342
rect 843 -376 877 -342
rect 912 -376 946 -342
rect 981 -376 1015 -342
rect 1050 -376 1084 -342
rect 1119 -376 1153 -342
rect 1188 -376 1222 -342
rect 1257 -376 1291 -342
rect 1326 -376 1360 -342
rect 1395 -376 1429 -342
rect 1464 -376 1498 -342
rect 1533 -376 1567 -342
rect 1602 -376 1636 -342
rect 1671 -376 1705 -342
rect 1740 -376 1774 -342
rect 1809 -376 1843 -342
rect 1878 -376 1912 -342
rect 1947 -376 1981 -342
rect 2016 -376 2050 -342
rect 2085 -376 2119 -342
rect 2154 -376 2188 -342
rect 2223 -376 2257 -342
rect 2292 -376 2326 -342
rect 2361 -376 2395 -342
rect 2430 -376 2464 -342
rect 2499 -376 2533 -342
rect 2568 -376 2602 -342
rect 2637 -376 2671 -342
rect 2706 -376 2740 -342
rect 2775 -376 2809 -342
rect 2844 -376 2878 -342
rect 2913 -376 2947 -342
rect 2982 -376 3016 -342
rect 3051 -376 3085 -342
rect 3120 -376 3154 -342
rect 3189 -376 3223 -342
rect 3258 -376 3292 -342
rect 3327 -376 3361 -342
rect -1020 -444 -986 -410
rect -951 -444 -917 -410
rect -882 -444 -848 -410
rect -813 -444 -779 -410
rect -744 -444 -710 -410
rect -675 -444 -641 -410
rect -606 -444 -572 -410
rect -537 -444 -503 -410
rect -468 -444 -434 -410
rect -399 -444 -365 -410
rect -330 -444 -296 -410
rect -261 -444 -227 -410
rect -192 -444 -158 -410
rect -123 -444 -89 -410
rect -54 -444 -20 -410
rect 15 -444 49 -410
rect 84 -444 118 -410
rect 153 -444 187 -410
rect 222 -444 256 -410
rect 291 -444 325 -410
rect 360 -444 394 -410
rect 429 -444 463 -410
rect 498 -444 532 -410
rect 567 -444 601 -410
rect 636 -444 670 -410
rect 705 -444 739 -410
rect 774 -444 808 -410
rect 843 -444 877 -410
rect 912 -444 946 -410
rect 981 -444 1015 -410
rect 1050 -444 1084 -410
rect 1119 -444 1153 -410
rect 1188 -444 1222 -410
rect 1257 -444 1291 -410
rect 1326 -444 1360 -410
rect 1395 -444 1429 -410
rect 1464 -444 1498 -410
rect 1533 -444 1567 -410
rect 1602 -444 1636 -410
rect 1671 -444 1705 -410
rect 1740 -444 1774 -410
rect 1809 -444 1843 -410
rect 1878 -444 1912 -410
rect 1947 -444 1981 -410
rect 2016 -444 2050 -410
rect 2085 -444 2119 -410
rect 2154 -444 2188 -410
rect 2223 -444 2257 -410
rect 2292 -444 2326 -410
rect 2361 -444 2395 -410
rect 2430 -444 2464 -410
rect 2499 -444 2533 -410
rect 2568 -444 2602 -410
rect 2637 -444 2671 -410
rect 2706 -444 2740 -410
rect 2775 -444 2809 -410
rect 2844 -444 2878 -410
rect 2913 -444 2947 -410
rect 2982 -444 3016 -410
rect 3051 -444 3085 -410
rect 3120 -444 3154 -410
rect 3189 -444 3223 -410
rect 3258 -444 3292 -410
rect 3327 -444 3361 -410
rect 3396 -444 13902 -274
<< poly >>
rect -40 3120 150 3198
tri -40 3100 -20 3120 ne
rect -20 3100 130 3120
tri 130 3100 150 3120 nw
rect 372 3120 562 3198
tri 372 3100 392 3120 ne
rect 392 3100 542 3120
tri 542 3100 562 3120 nw
rect 784 3120 974 3198
tri 784 3100 804 3120 ne
rect 804 3100 954 3120
tri 954 3100 974 3120 nw
rect 1196 3120 1386 3198
tri 1196 3100 1216 3120 ne
rect 1216 3100 1366 3120
tri 1366 3100 1386 3120 nw
rect 1608 3120 1798 3198
tri 1608 3100 1628 3120 ne
rect 1628 3100 1778 3120
tri 1778 3100 1798 3120 nw
rect 2020 3120 2210 3198
tri 2020 3100 2040 3120 ne
rect 2040 3100 2190 3120
tri 2190 3100 2210 3120 nw
rect 2432 3120 2622 3198
tri 2432 3100 2452 3120 ne
rect 2452 3100 2602 3120
tri 2602 3100 2622 3120 nw
rect 2844 3120 3034 3198
tri 2844 3100 2864 3120 ne
rect 2864 3100 3014 3120
tri 3014 3100 3034 3120 nw
rect 3256 3120 3446 3198
tri 3256 3100 3276 3120 ne
rect 3276 3100 3426 3120
tri 3426 3100 3446 3120 nw
rect 3668 3120 3858 3198
tri 3668 3100 3688 3120 ne
rect 3688 3100 3838 3120
tri 3838 3100 3858 3120 nw
rect 4080 3120 4270 3198
tri 4080 3100 4100 3120 ne
rect 4100 3100 4250 3120
tri 4250 3100 4270 3120 nw
rect 4492 3120 4682 3198
tri 4492 3100 4512 3120 ne
rect 4512 3100 4662 3120
tri 4662 3100 4682 3120 nw
rect 4904 3120 5094 3198
tri 4904 3100 4924 3120 ne
rect 4924 3100 5074 3120
tri 5074 3100 5094 3120 nw
rect 5316 3120 5506 3198
tri 5316 3100 5336 3120 ne
rect 5336 3100 5486 3120
tri 5486 3100 5506 3120 nw
rect 5728 3120 5918 3198
tri 5728 3100 5748 3120 ne
rect 5748 3100 5898 3120
tri 5898 3100 5918 3120 nw
rect 6140 3120 6330 3198
tri 6140 3100 6160 3120 ne
rect 6160 3100 6310 3120
tri 6310 3100 6330 3120 nw
rect 6552 3120 6742 3198
tri 6552 3100 6572 3120 ne
rect 6572 3100 6722 3120
tri 6722 3100 6742 3120 nw
rect 6964 3120 7154 3198
tri 6964 3100 6984 3120 ne
rect 6984 3100 7134 3120
tri 7134 3100 7154 3120 nw
rect 7376 3120 7566 3198
tri 7376 3100 7396 3120 ne
rect 7396 3100 7546 3120
tri 7546 3100 7566 3120 nw
rect 7788 3120 7978 3198
tri 7788 3100 7808 3120 ne
rect 7808 3100 7958 3120
tri 7958 3100 7978 3120 nw
rect 8200 3120 8390 3198
tri 8200 3100 8220 3120 ne
rect 8220 3100 8370 3120
tri 8370 3100 8390 3120 nw
rect 8612 3120 8802 3198
tri 8612 3100 8632 3120 ne
rect 8632 3100 8782 3120
tri 8782 3100 8802 3120 nw
rect 9024 3120 9214 3198
tri 9024 3100 9044 3120 ne
rect 9044 3100 9194 3120
tri 9194 3100 9214 3120 nw
rect 9436 3120 9626 3198
tri 9436 3100 9456 3120 ne
rect 9456 3100 9606 3120
tri 9606 3100 9626 3120 nw
rect 9848 3120 10038 3198
tri 9848 3100 9868 3120 ne
rect 9868 3100 10018 3120
tri 10018 3100 10038 3120 nw
rect 10260 3120 10450 3198
tri 10260 3100 10280 3120 ne
rect 10280 3100 10430 3120
tri 10430 3100 10450 3120 nw
rect 10672 3120 10862 3198
tri 10672 3100 10692 3120 ne
rect 10692 3100 10842 3120
tri 10842 3100 10862 3120 nw
rect 11084 3120 11274 3198
tri 11084 3100 11104 3120 ne
rect 11104 3100 11254 3120
tri 11254 3100 11274 3120 nw
rect 11496 3120 11686 3198
tri 11496 3100 11516 3120 ne
rect 11516 3100 11666 3120
tri 11666 3100 11686 3120 nw
rect 11908 3120 12098 3198
tri 11908 3100 11928 3120 ne
rect 11928 3100 12078 3120
tri 12078 3100 12098 3120 nw
rect 12320 3120 12510 3198
tri 12320 3100 12340 3120 ne
rect 12340 3100 12490 3120
tri 12490 3100 12510 3120 nw
rect 12732 3120 12922 3198
tri 12732 3100 12752 3120 ne
rect 12752 3100 12902 3120
tri 12902 3100 12922 3120 nw
tri -40 -20 -20 0 se
rect -20 -20 130 0
tri 130 -20 150 0 sw
rect -40 -98 150 -20
tri 372 -20 392 0 se
rect 392 -20 542 0
tri 542 -20 562 0 sw
rect 372 -98 562 -20
tri 784 -20 804 0 se
rect 804 -20 954 0
tri 954 -20 974 0 sw
rect 784 -98 974 -20
tri 1196 -20 1216 0 se
rect 1216 -20 1366 0
tri 1366 -20 1386 0 sw
rect 1196 -98 1386 -20
tri 1608 -20 1628 0 se
rect 1628 -20 1778 0
tri 1778 -20 1798 0 sw
rect 1608 -98 1798 -20
tri 2020 -20 2040 0 se
rect 2040 -20 2190 0
tri 2190 -20 2210 0 sw
rect 2020 -98 2210 -20
tri 2432 -20 2452 0 se
rect 2452 -20 2602 0
tri 2602 -20 2622 0 sw
rect 2432 -98 2622 -20
tri 2844 -20 2864 0 se
rect 2864 -20 3014 0
tri 3014 -20 3034 0 sw
rect 2844 -98 3034 -20
tri 3256 -20 3276 0 se
rect 3276 -20 3426 0
tri 3426 -20 3446 0 sw
rect 3256 -98 3446 -20
tri 3668 -20 3688 0 se
rect 3688 -20 3838 0
tri 3838 -20 3858 0 sw
rect 3668 -98 3858 -20
tri 4080 -20 4100 0 se
rect 4100 -20 4250 0
tri 4250 -20 4270 0 sw
rect 4080 -98 4270 -20
tri 4492 -20 4512 0 se
rect 4512 -20 4662 0
tri 4662 -20 4682 0 sw
rect 4492 -98 4682 -20
tri 4904 -20 4924 0 se
rect 4924 -20 5074 0
tri 5074 -20 5094 0 sw
rect 4904 -98 5094 -20
tri 5316 -20 5336 0 se
rect 5336 -20 5486 0
tri 5486 -20 5506 0 sw
rect 5316 -98 5506 -20
tri 5728 -20 5748 0 se
rect 5748 -20 5898 0
tri 5898 -20 5918 0 sw
rect 5728 -98 5918 -20
tri 6140 -20 6160 0 se
rect 6160 -20 6310 0
tri 6310 -20 6330 0 sw
rect 6140 -98 6330 -20
tri 6552 -20 6572 0 se
rect 6572 -20 6722 0
tri 6722 -20 6742 0 sw
rect 6552 -98 6742 -20
tri 6964 -20 6984 0 se
rect 6984 -20 7134 0
tri 7134 -20 7154 0 sw
rect 6964 -98 7154 -20
tri 7376 -20 7396 0 se
rect 7396 -20 7546 0
tri 7546 -20 7566 0 sw
rect 7376 -98 7566 -20
tri 7788 -20 7808 0 se
rect 7808 -20 7958 0
tri 7958 -20 7978 0 sw
rect 7788 -98 7978 -20
tri 8200 -20 8220 0 se
rect 8220 -20 8370 0
tri 8370 -20 8390 0 sw
rect 8200 -98 8390 -20
tri 8612 -20 8632 0 se
rect 8632 -20 8782 0
tri 8782 -20 8802 0 sw
rect 8612 -98 8802 -20
tri 9024 -20 9044 0 se
rect 9044 -20 9194 0
tri 9194 -20 9214 0 sw
rect 9024 -98 9214 -20
tri 9436 -20 9456 0 se
rect 9456 -20 9606 0
tri 9606 -20 9626 0 sw
rect 9436 -98 9626 -20
tri 9848 -20 9868 0 se
rect 9868 -20 10018 0
tri 10018 -20 10038 0 sw
rect 9848 -98 10038 -20
tri 10260 -20 10280 0 se
rect 10280 -20 10430 0
tri 10430 -20 10450 0 sw
rect 10260 -98 10450 -20
tri 10672 -20 10692 0 se
rect 10692 -20 10842 0
tri 10842 -20 10862 0 sw
rect 10672 -98 10862 -20
tri 11084 -20 11104 0 se
rect 11104 -20 11254 0
tri 11254 -20 11274 0 sw
rect 11084 -98 11274 -20
tri 11496 -20 11516 0 se
rect 11516 -20 11666 0
tri 11666 -20 11686 0 sw
rect 11496 -98 11686 -20
tri 11908 -20 11928 0 se
rect 11928 -20 12078 0
tri 12078 -20 12098 0 sw
rect 11908 -98 12098 -20
tri 12320 -20 12340 0 se
rect 12340 -20 12490 0
tri 12490 -20 12510 0 sw
rect 12320 -98 12510 -20
tri 12732 -20 12752 0 se
rect 12752 -20 12902 0
tri 12902 -20 12922 0 sw
rect 12732 -98 12922 -20
<< locali >>
rect -1458 3880 -1390 3914
rect -1356 3880 -1321 3914
rect -1287 3880 -1252 3914
rect -1218 3882 -1183 3914
rect -1149 3882 -1114 3914
rect -1218 3880 -1191 3882
rect -1149 3880 -1118 3882
rect -1080 3880 -1045 3914
rect -1011 3880 -976 3914
rect -942 3882 -907 3914
rect -873 3882 -838 3914
rect -804 3882 -769 3914
rect -735 3882 -700 3914
rect -666 3882 -631 3914
rect -597 3882 -562 3914
rect -528 3882 -493 3914
rect -459 3882 -424 3914
rect -938 3880 -907 3882
rect -865 3880 -838 3882
rect -792 3880 -769 3882
rect -719 3880 -700 3882
rect -646 3880 -631 3882
rect -573 3880 -562 3882
rect -500 3880 -493 3882
rect -427 3880 -424 3882
rect -390 3882 -355 3914
rect -321 3882 -286 3914
rect -252 3882 -217 3914
rect -183 3882 -148 3914
rect -114 3882 -79 3914
rect -45 3882 -10 3914
rect 24 3882 59 3914
rect 93 3882 128 3914
rect 162 3882 197 3914
rect -390 3880 -388 3882
rect -321 3880 -315 3882
rect -252 3880 -242 3882
rect -183 3880 -169 3882
rect -114 3880 -96 3882
rect -45 3880 -23 3882
rect 24 3880 50 3882
rect 93 3880 123 3882
rect 162 3880 196 3882
rect 231 3880 266 3914
rect 300 3882 335 3914
rect 369 3882 404 3914
rect 438 3882 473 3914
rect 507 3882 542 3914
rect 576 3882 611 3914
rect 645 3882 680 3914
rect 714 3882 749 3914
rect 783 3882 818 3914
rect 303 3880 335 3882
rect 376 3880 404 3882
rect 449 3880 473 3882
rect 522 3880 542 3882
rect 595 3880 611 3882
rect 668 3880 680 3882
rect 741 3880 749 3882
rect 814 3880 818 3882
rect 852 3882 887 3914
rect 852 3880 853 3882
rect -1458 3848 -1191 3880
rect -1157 3848 -1118 3880
rect -1084 3848 -1045 3880
rect -1011 3848 -972 3880
rect -938 3848 -899 3880
rect -865 3848 -826 3880
rect -792 3848 -753 3880
rect -719 3848 -680 3880
rect -646 3848 -607 3880
rect -573 3848 -534 3880
rect -500 3848 -461 3880
rect -427 3848 -388 3880
rect -354 3848 -315 3880
rect -281 3848 -242 3880
rect -208 3848 -169 3880
rect -135 3848 -96 3880
rect -62 3848 -23 3880
rect 11 3848 50 3880
rect 84 3848 123 3880
rect 157 3848 196 3880
rect 230 3848 269 3880
rect 303 3848 342 3880
rect 376 3848 415 3880
rect 449 3848 488 3880
rect 522 3848 561 3880
rect 595 3848 634 3880
rect 668 3848 707 3880
rect 741 3848 780 3880
rect 814 3848 853 3880
rect 921 3882 956 3914
rect 990 3882 1025 3914
rect 1059 3882 1094 3914
rect 1128 3882 1163 3914
rect 1197 3882 1232 3914
rect 1266 3882 1301 3914
rect 1335 3882 1370 3914
rect 1404 3882 1439 3914
rect 921 3880 926 3882
rect 990 3880 999 3882
rect 1059 3880 1072 3882
rect 1128 3880 1145 3882
rect 1197 3880 1218 3882
rect 1266 3880 1291 3882
rect 1335 3880 1364 3882
rect 1404 3880 1437 3882
rect 1473 3880 1508 3914
rect 1542 3882 1577 3914
rect 1611 3882 1646 3914
rect 1680 3882 1715 3914
rect 1749 3882 1784 3914
rect 1818 3882 1853 3914
rect 1887 3882 1922 3914
rect 1956 3882 1991 3914
rect 2025 3882 2060 3914
rect 2094 3882 2129 3914
rect 2163 3882 2198 3914
rect 2232 3882 2267 3914
rect 2301 3882 2336 3914
rect 2370 3882 2405 3914
rect 2439 3882 2474 3914
rect 1544 3880 1577 3882
rect 887 3848 926 3880
rect 960 3848 999 3880
rect 1033 3848 1072 3880
rect 1106 3848 1145 3880
rect 1179 3848 1218 3880
rect 1252 3848 1291 3880
rect 1325 3848 1364 3880
rect 1398 3848 1437 3880
rect 1471 3848 1510 3880
rect 1544 3848 1583 3880
rect -1458 3846 1583 3848
rect -1458 3812 -1390 3846
rect -1356 3812 -1321 3846
rect -1287 3812 -1252 3846
rect -1218 3812 -1183 3846
rect -1149 3812 -1114 3846
rect -1080 3812 -1045 3846
rect -1011 3812 -976 3846
rect -942 3812 -907 3846
rect -873 3812 -838 3846
rect -804 3812 -769 3846
rect -735 3812 -700 3846
rect -666 3812 -631 3846
rect -597 3812 -562 3846
rect -528 3812 -493 3846
rect -459 3812 -424 3846
rect -390 3812 -355 3846
rect -321 3812 -286 3846
rect -252 3812 -217 3846
rect -183 3812 -148 3846
rect -114 3812 -79 3846
rect -45 3812 -10 3846
rect 24 3812 59 3846
rect 93 3812 128 3846
rect 162 3812 197 3846
rect 231 3812 266 3846
rect 300 3812 335 3846
rect 369 3812 404 3846
rect 438 3812 473 3846
rect 507 3812 542 3846
rect 576 3812 611 3846
rect 645 3812 680 3846
rect 714 3812 749 3846
rect 783 3812 818 3846
rect 852 3812 887 3846
rect 921 3812 956 3846
rect 990 3812 1025 3846
rect 1059 3812 1094 3846
rect 1128 3812 1163 3846
rect 1197 3812 1232 3846
rect 1266 3812 1301 3846
rect 1335 3812 1370 3846
rect 1404 3812 1439 3846
rect 1473 3812 1508 3846
rect 1542 3812 1577 3846
rect -1458 3810 1583 3812
rect -1458 3778 -1191 3810
rect -1157 3778 -1118 3810
rect -1084 3778 -1045 3810
rect -1011 3778 -972 3810
rect -938 3778 -899 3810
rect -865 3778 -826 3810
rect -792 3778 -753 3810
rect -719 3778 -680 3810
rect -646 3778 -607 3810
rect -573 3778 -534 3810
rect -500 3778 -461 3810
rect -427 3778 -388 3810
rect -354 3778 -315 3810
rect -281 3778 -242 3810
rect -208 3778 -169 3810
rect -135 3778 -96 3810
rect -62 3778 -23 3810
rect 11 3778 50 3810
rect 84 3778 123 3810
rect 157 3778 196 3810
rect 230 3778 269 3810
rect 303 3778 342 3810
rect 376 3778 415 3810
rect 449 3778 488 3810
rect 522 3778 561 3810
rect 595 3778 634 3810
rect 668 3778 707 3810
rect 741 3778 780 3810
rect 814 3778 853 3810
rect -1458 3744 -1390 3778
rect -1356 3744 -1321 3778
rect -1287 3744 -1252 3778
rect -1218 3776 -1191 3778
rect -1149 3776 -1118 3778
rect -1218 3744 -1183 3776
rect -1149 3744 -1114 3776
rect -1080 3744 -1045 3778
rect -1011 3744 -976 3778
rect -938 3776 -907 3778
rect -865 3776 -838 3778
rect -792 3776 -769 3778
rect -719 3776 -700 3778
rect -646 3776 -631 3778
rect -573 3776 -562 3778
rect -500 3776 -493 3778
rect -427 3776 -424 3778
rect -942 3744 -907 3776
rect -873 3744 -838 3776
rect -804 3744 -769 3776
rect -735 3744 -700 3776
rect -666 3744 -631 3776
rect -597 3744 -562 3776
rect -528 3744 -493 3776
rect -459 3744 -424 3776
rect -390 3776 -388 3778
rect -321 3776 -315 3778
rect -252 3776 -242 3778
rect -183 3776 -169 3778
rect -114 3776 -96 3778
rect -45 3776 -23 3778
rect 24 3776 50 3778
rect 93 3776 123 3778
rect 162 3776 196 3778
rect -390 3744 -355 3776
rect -321 3744 -286 3776
rect -252 3744 -217 3776
rect -183 3744 -148 3776
rect -114 3744 -79 3776
rect -45 3744 -10 3776
rect 24 3744 59 3776
rect 93 3744 128 3776
rect 162 3744 197 3776
rect 231 3744 266 3778
rect 303 3776 335 3778
rect 376 3776 404 3778
rect 449 3776 473 3778
rect 522 3776 542 3778
rect 595 3776 611 3778
rect 668 3776 680 3778
rect 741 3776 749 3778
rect 814 3776 818 3778
rect 300 3744 335 3776
rect 369 3744 404 3776
rect 438 3744 473 3776
rect 507 3744 542 3776
rect 576 3744 611 3776
rect 645 3744 680 3776
rect 714 3744 749 3776
rect 783 3744 818 3776
rect 852 3776 853 3778
rect 887 3778 926 3810
rect 960 3778 999 3810
rect 1033 3778 1072 3810
rect 1106 3778 1145 3810
rect 1179 3778 1218 3810
rect 1252 3778 1291 3810
rect 1325 3778 1364 3810
rect 1398 3778 1437 3810
rect 1471 3778 1510 3810
rect 1544 3778 1583 3810
rect 852 3744 887 3776
rect 921 3776 926 3778
rect 990 3776 999 3778
rect 1059 3776 1072 3778
rect 1128 3776 1145 3778
rect 1197 3776 1218 3778
rect 1266 3776 1291 3778
rect 1335 3776 1364 3778
rect 1404 3776 1437 3778
rect 921 3744 956 3776
rect 990 3744 1025 3776
rect 1059 3744 1094 3776
rect 1128 3744 1163 3776
rect 1197 3744 1232 3776
rect 1266 3744 1301 3776
rect 1335 3744 1370 3776
rect 1404 3744 1439 3776
rect 1473 3744 1508 3778
rect 1544 3776 1577 3778
rect 1542 3744 1577 3776
rect 1611 3744 1646 3776
rect 1680 3744 1715 3776
rect 1749 3744 1784 3776
rect 1818 3744 1853 3776
rect 1887 3744 1922 3776
rect 1956 3744 1991 3776
rect 2025 3744 2060 3776
rect 2094 3744 2129 3776
rect 2163 3744 2198 3776
rect 2232 3744 2267 3776
rect 2301 3744 2336 3776
rect 2370 3744 2405 3776
rect 2439 3744 2474 3776
rect 14272 3744 14340 3914
rect -1458 3676 -1288 3744
rect 14170 3676 14340 3744
rect -1458 -440 -1288 -438
rect -1458 -473 -1426 -440
rect -1392 -473 -1354 -440
rect -1320 -473 -1288 -440
rect -1088 3510 -1020 3544
rect -986 3510 -951 3544
rect -917 3512 -882 3544
rect -917 3510 -886 3512
rect -848 3510 -813 3544
rect -779 3510 -744 3544
rect -710 3512 -675 3544
rect -641 3512 -606 3544
rect -572 3512 -537 3544
rect -503 3512 -468 3544
rect -434 3512 -399 3544
rect -365 3512 -330 3544
rect -296 3512 -261 3544
rect -227 3512 -192 3544
rect -158 3512 -123 3544
rect -89 3512 -54 3544
rect -20 3512 15 3544
rect 49 3512 84 3544
rect 118 3512 153 3544
rect 187 3512 222 3544
rect 256 3512 291 3544
rect 325 3512 360 3544
rect 394 3512 429 3544
rect 463 3512 498 3544
rect 532 3512 567 3544
rect 601 3512 636 3544
rect 670 3512 705 3544
rect 739 3512 774 3544
rect 808 3512 843 3544
rect 877 3512 912 3544
rect 946 3512 981 3544
rect 1015 3512 1050 3544
rect 1084 3512 1119 3544
rect 1153 3512 1188 3544
rect 1222 3512 1257 3544
rect 1291 3512 1326 3544
rect 1360 3512 1395 3544
rect 1429 3512 1464 3544
rect 1498 3512 1533 3544
rect 1567 3512 1602 3544
rect 1636 3512 1671 3544
rect 1705 3512 1740 3544
rect 1774 3512 1809 3544
rect 1843 3512 1878 3544
rect 1912 3512 1947 3544
rect 1981 3512 2016 3544
rect 2050 3512 2085 3544
rect 2119 3512 2154 3544
rect 2188 3512 2223 3544
rect 2257 3512 2292 3544
rect 2326 3512 2361 3544
rect 2395 3512 2430 3544
rect 2464 3512 2499 3544
rect 2533 3512 2568 3544
rect 2602 3512 2637 3544
rect 2671 3512 2706 3544
rect 2740 3512 2775 3544
rect 2809 3512 2844 3544
rect 2878 3512 2913 3544
rect 2947 3512 2982 3544
rect 3016 3512 3051 3544
rect 3085 3512 3120 3544
rect 3154 3512 3189 3544
rect 3223 3512 3258 3544
rect 3292 3512 3327 3544
rect 3361 3512 3396 3544
rect -706 3510 -675 3512
rect -633 3510 -606 3512
rect -1088 3478 -886 3510
rect -852 3478 -813 3510
rect -779 3478 -740 3510
rect -706 3478 -667 3510
rect -633 3478 -594 3510
rect -1088 3476 -594 3478
rect -1088 3442 -1020 3476
rect -986 3442 -951 3476
rect -917 3442 -882 3476
rect -848 3442 -813 3476
rect -779 3442 -744 3476
rect -710 3442 -675 3476
rect -641 3442 -606 3476
rect -1088 3440 -594 3442
rect -1088 3408 -886 3440
rect -852 3408 -813 3440
rect -779 3408 -740 3440
rect -706 3408 -667 3440
rect -633 3408 -594 3440
rect -1088 3374 -1020 3408
rect -986 3374 -951 3408
rect -917 3406 -886 3408
rect -917 3374 -882 3406
rect -848 3374 -813 3408
rect -779 3374 -744 3408
rect -706 3406 -675 3408
rect -633 3406 -606 3408
rect -710 3374 -675 3406
rect -641 3374 -606 3406
rect -572 3374 -537 3406
rect -503 3374 -468 3406
rect -434 3374 -399 3406
rect -365 3374 -330 3406
rect -296 3374 -261 3406
rect -227 3374 -192 3406
rect -158 3374 -123 3406
rect -89 3374 -54 3406
rect -20 3374 15 3406
rect 49 3374 84 3406
rect 118 3374 153 3406
rect 187 3374 222 3406
rect 256 3374 291 3406
rect 325 3374 360 3406
rect 394 3374 429 3406
rect 463 3374 498 3406
rect 532 3374 567 3406
rect 601 3374 636 3406
rect 670 3374 705 3406
rect 739 3374 774 3406
rect 808 3374 843 3406
rect 877 3374 912 3406
rect 946 3374 981 3406
rect 1015 3374 1050 3406
rect 1084 3374 1119 3406
rect 1153 3374 1188 3406
rect 1222 3374 1257 3406
rect 1291 3374 1326 3406
rect 1360 3374 1395 3406
rect 1429 3374 1464 3406
rect 1498 3374 1533 3406
rect 1567 3374 1602 3406
rect 1636 3374 1671 3406
rect 1705 3374 1740 3406
rect 1774 3374 1809 3406
rect 1843 3374 1878 3406
rect 1912 3374 1947 3406
rect 1981 3374 2016 3406
rect 2050 3374 2085 3406
rect 2119 3374 2154 3406
rect 2188 3374 2223 3406
rect 2257 3374 2292 3406
rect 2326 3374 2361 3406
rect 2395 3374 2430 3406
rect 2464 3374 2499 3406
rect 2533 3374 2568 3406
rect 2602 3374 2637 3406
rect 2671 3374 2706 3406
rect 2740 3374 2775 3406
rect 2809 3374 2844 3406
rect 2878 3374 2913 3406
rect 2947 3374 2982 3406
rect 3016 3374 3051 3406
rect 3085 3374 3120 3406
rect 3154 3374 3189 3406
rect 3223 3374 3258 3406
rect 3292 3374 3327 3406
rect 3361 3374 3396 3406
rect 13902 3374 13970 3544
rect -1088 3306 -306 3374
rect 13188 3306 13970 3374
rect -1088 480 -1074 484
rect -1040 480 -1002 484
rect -968 480 -930 484
rect -896 480 -858 484
rect -824 480 -786 484
rect -752 480 -714 484
rect -680 480 -642 484
rect -608 480 -570 484
rect -536 480 -498 484
rect -464 480 -426 484
rect -392 480 -354 484
rect -320 480 -306 484
rect -1088 449 -306 480
rect -1054 441 -1020 449
rect -986 441 -952 449
rect -918 441 -884 449
rect -850 441 -816 449
rect -782 441 -748 449
rect -1040 415 -1020 441
rect -968 415 -952 441
rect -896 415 -884 441
rect -824 415 -816 441
rect -752 415 -748 441
rect -714 441 -680 449
rect -1088 407 -1074 415
rect -1040 407 -1002 415
rect -968 407 -930 415
rect -896 407 -858 415
rect -824 407 -786 415
rect -752 407 -714 415
rect -646 441 -612 449
rect -578 441 -544 449
rect -510 441 -476 449
rect -442 441 -408 449
rect -374 441 -340 449
rect -646 415 -642 441
rect -578 415 -570 441
rect -510 415 -498 441
rect -442 415 -426 441
rect -374 415 -354 441
rect -680 407 -642 415
rect -608 407 -570 415
rect -536 407 -498 415
rect -464 407 -426 415
rect -392 407 -354 415
rect -320 407 -306 415
rect -1088 380 -306 407
rect -1054 368 -1020 380
rect -986 368 -952 380
rect -918 368 -884 380
rect -850 368 -816 380
rect -782 368 -748 380
rect -1040 346 -1020 368
rect -968 346 -952 368
rect -896 346 -884 368
rect -824 346 -816 368
rect -752 346 -748 368
rect -714 368 -680 380
rect -1088 334 -1074 346
rect -1040 334 -1002 346
rect -968 334 -930 346
rect -896 334 -858 346
rect -824 334 -786 346
rect -752 334 -714 346
rect -646 368 -612 380
rect -578 368 -544 380
rect -510 368 -476 380
rect -442 368 -408 380
rect -374 368 -340 380
rect -646 346 -642 368
rect -578 346 -570 368
rect -510 346 -498 368
rect -442 346 -426 368
rect -374 346 -354 368
rect -680 334 -642 346
rect -608 334 -570 346
rect -536 334 -498 346
rect -464 334 -426 346
rect -392 334 -354 346
rect -320 334 -306 346
rect -1088 311 -306 334
rect -1054 295 -1020 311
rect -986 295 -952 311
rect -918 295 -884 311
rect -850 295 -816 311
rect -782 295 -748 311
rect -1040 277 -1020 295
rect -968 277 -952 295
rect -896 277 -884 295
rect -824 277 -816 295
rect -752 277 -748 295
rect -714 295 -680 311
rect -1088 261 -1074 277
rect -1040 261 -1002 277
rect -968 261 -930 277
rect -896 261 -858 277
rect -824 261 -786 277
rect -752 261 -714 277
rect -646 295 -612 311
rect -578 295 -544 311
rect -510 295 -476 311
rect -442 295 -408 311
rect -374 295 -340 311
rect -646 277 -642 295
rect -578 277 -570 295
rect -510 277 -498 295
rect -442 277 -426 295
rect -374 277 -354 295
rect -680 261 -642 277
rect -608 261 -570 277
rect -536 261 -498 277
rect -464 261 -426 277
rect -392 261 -354 277
rect -320 261 -306 277
rect -1088 242 -306 261
rect -1054 222 -1020 242
rect -986 222 -952 242
rect -918 222 -884 242
rect -850 222 -816 242
rect -782 222 -748 242
rect -1040 208 -1020 222
rect -968 208 -952 222
rect -896 208 -884 222
rect -824 208 -816 222
rect -752 208 -748 222
rect -714 222 -680 242
rect -1088 188 -1074 208
rect -1040 188 -1002 208
rect -968 188 -930 208
rect -896 188 -858 208
rect -824 188 -786 208
rect -752 188 -714 208
rect -646 222 -612 242
rect -578 222 -544 242
rect -510 222 -476 242
rect -442 222 -408 242
rect -374 222 -340 242
rect -646 208 -642 222
rect -578 208 -570 222
rect -510 208 -498 222
rect -442 208 -426 222
rect -374 208 -354 222
rect -680 188 -642 208
rect -608 188 -570 208
rect -536 188 -498 208
rect -464 188 -426 208
rect -392 188 -354 208
rect -320 188 -306 208
rect -1088 173 -306 188
rect -1054 149 -1020 173
rect -986 149 -952 173
rect -918 149 -884 173
rect -850 149 -816 173
rect -782 149 -748 173
rect -1040 139 -1020 149
rect -968 139 -952 149
rect -896 139 -884 149
rect -824 139 -816 149
rect -752 139 -748 149
rect -714 149 -680 173
rect -1088 115 -1074 139
rect -1040 115 -1002 139
rect -968 115 -930 139
rect -896 115 -858 139
rect -824 115 -786 139
rect -752 115 -714 139
rect -646 149 -612 173
rect -578 149 -544 173
rect -510 149 -476 173
rect -442 149 -408 173
rect -374 149 -340 173
rect -646 139 -642 149
rect -578 139 -570 149
rect -510 139 -498 149
rect -442 139 -426 149
rect -374 139 -354 149
rect -680 115 -642 139
rect -608 115 -570 139
rect -536 115 -498 139
rect -464 115 -426 139
rect -392 115 -354 139
rect -320 115 -306 139
rect -1088 104 -306 115
rect -1054 76 -1020 104
rect -986 76 -952 104
rect -918 76 -884 104
rect -850 76 -816 104
rect -782 76 -748 104
rect -1040 70 -1020 76
rect -968 70 -952 76
rect -896 70 -884 76
rect -824 70 -816 76
rect -752 70 -748 76
rect -714 76 -680 104
rect -1088 42 -1074 70
rect -1040 42 -1002 70
rect -968 42 -930 70
rect -896 42 -858 70
rect -824 42 -786 70
rect -752 42 -714 70
rect -646 76 -612 104
rect -578 76 -544 104
rect -510 76 -476 104
rect -442 76 -408 104
rect -374 76 -340 104
rect -646 70 -642 76
rect -578 70 -570 76
rect -510 70 -498 76
rect -442 70 -426 76
rect -374 70 -354 76
rect -680 42 -642 70
rect -608 42 -570 70
rect -536 42 -498 70
rect -464 42 -426 70
rect -392 42 -354 70
rect -320 42 -306 70
rect -1088 35 -306 42
rect -1054 3 -1020 35
rect -986 3 -952 35
rect -918 3 -884 35
rect -850 3 -816 35
rect -782 3 -748 35
rect -1040 1 -1020 3
rect -968 1 -952 3
rect -896 1 -884 3
rect -824 1 -816 3
rect -752 1 -748 3
rect -714 3 -680 35
rect -1088 -31 -1074 1
rect -1040 -31 -1002 1
rect -968 -31 -930 1
rect -896 -31 -858 1
rect -824 -31 -786 1
rect -752 -31 -714 1
rect -646 3 -612 35
rect -578 3 -544 35
rect -510 3 -476 35
rect -442 3 -408 35
rect -374 3 -340 35
rect -646 1 -642 3
rect -578 1 -570 3
rect -510 1 -498 3
rect -442 1 -426 3
rect -374 1 -354 3
rect -680 -31 -642 1
rect -608 -31 -570 1
rect -536 -31 -498 1
rect -464 -31 -426 1
rect -392 -31 -354 1
rect -320 -31 -306 1
rect -204 3000 -98 3100
rect -204 2927 -202 2966
rect -100 2927 -98 2966
rect -204 2854 -202 2893
rect -100 2854 -98 2893
rect -204 2781 -202 2820
rect -100 2781 -98 2820
rect -204 2708 -202 2747
rect -100 2708 -98 2747
rect -204 2635 -202 2674
rect -100 2635 -98 2674
rect -204 2562 -202 2601
rect -100 2562 -98 2601
rect -204 2489 -202 2528
rect -100 2489 -98 2528
rect -204 2416 -202 2455
rect -100 2416 -98 2455
rect -204 2343 -202 2382
rect -100 2343 -98 2382
rect -204 2270 -202 2309
rect -100 2270 -98 2309
rect -204 2197 -202 2236
rect -100 2197 -98 2236
rect -204 2124 -202 2163
rect -100 2124 -98 2163
rect -204 2051 -202 2090
rect -100 2051 -98 2090
rect -204 1978 -202 2017
rect -100 1978 -98 2017
rect -204 1905 -202 1944
rect -100 1905 -98 1944
rect -204 1832 -202 1871
rect -100 1832 -98 1871
rect -204 1759 -202 1798
rect -100 1759 -98 1798
rect -204 1686 -202 1725
rect -100 1686 -98 1725
rect -204 1613 -202 1652
rect -100 1613 -98 1652
rect -204 1540 -202 1579
rect -100 1540 -98 1579
rect -204 1466 -202 1506
rect -100 1466 -98 1506
rect -204 1392 -202 1432
rect -100 1392 -98 1432
rect -204 1318 -202 1358
rect -100 1318 -98 1358
rect -204 1244 -202 1284
rect -100 1244 -98 1284
rect -204 1170 -202 1210
rect -100 1170 -98 1210
rect -204 1096 -202 1136
rect -100 1096 -98 1136
rect -204 1022 -202 1062
rect -100 1022 -98 1062
rect -204 948 -202 988
rect -100 948 -98 988
rect -204 874 -202 914
rect -100 874 -98 914
rect -204 800 -202 840
rect -100 800 -98 840
rect -170 766 -132 790
rect -204 755 -98 766
rect -204 726 -202 755
rect -168 721 -134 755
rect -100 726 -98 755
rect -170 692 -132 721
rect -204 686 -98 692
rect -204 652 -202 686
rect -168 652 -134 686
rect -100 652 -98 686
rect -170 618 -132 652
rect -204 617 -98 618
rect -204 583 -202 617
rect -168 583 -134 617
rect -100 583 -98 617
rect -204 578 -98 583
rect -170 548 -132 578
rect -204 514 -202 544
rect -168 514 -134 548
rect -100 514 -98 544
rect -204 504 -98 514
rect -170 479 -132 504
rect -204 445 -202 470
rect -168 445 -134 479
rect -100 445 -98 470
rect -204 430 -98 445
rect -170 410 -132 430
rect -204 376 -202 396
rect -168 376 -134 410
rect -100 376 -98 396
rect -204 356 -98 376
rect -170 341 -132 356
rect -204 307 -202 322
rect -168 307 -134 341
rect -100 307 -98 322
rect -204 282 -98 307
rect -170 272 -132 282
rect -204 238 -202 248
rect -168 238 -134 272
rect -100 238 -98 248
rect -204 208 -98 238
rect -170 203 -132 208
rect -204 169 -202 174
rect -168 169 -134 203
rect -100 169 -98 174
rect -204 134 -98 169
rect -168 100 -134 134
rect -204 0 -98 100
rect 208 3000 314 3100
rect 208 2927 210 2966
rect 312 2927 314 2966
rect 208 2854 210 2893
rect 312 2854 314 2893
rect 208 2781 210 2820
rect 312 2781 314 2820
rect 208 2708 210 2747
rect 312 2708 314 2747
rect 208 2635 210 2674
rect 312 2635 314 2674
rect 208 2562 210 2601
rect 312 2562 314 2601
rect 208 2489 210 2528
rect 312 2489 314 2528
rect 208 2416 210 2455
rect 312 2416 314 2455
rect 208 2343 210 2382
rect 312 2343 314 2382
rect 208 2270 210 2309
rect 312 2270 314 2309
rect 208 2197 210 2236
rect 312 2197 314 2236
rect 208 2124 210 2163
rect 312 2124 314 2163
rect 208 2051 210 2090
rect 312 2051 314 2090
rect 208 1978 210 2017
rect 312 1978 314 2017
rect 208 1905 210 1944
rect 312 1905 314 1944
rect 208 1832 210 1871
rect 312 1832 314 1871
rect 208 1759 210 1798
rect 312 1759 314 1798
rect 208 1686 210 1725
rect 312 1686 314 1725
rect 208 1613 210 1652
rect 312 1613 314 1652
rect 208 1540 210 1579
rect 312 1540 314 1579
rect 208 1466 210 1506
rect 312 1466 314 1506
rect 208 1392 210 1432
rect 312 1392 314 1432
rect 208 1318 210 1358
rect 312 1318 314 1358
rect 208 1244 210 1284
rect 312 1244 314 1284
rect 208 1170 210 1210
rect 312 1170 314 1210
rect 208 1096 210 1136
rect 312 1096 314 1136
rect 208 1022 210 1062
rect 312 1022 314 1062
rect 208 948 210 988
rect 312 948 314 988
rect 208 874 210 914
rect 312 874 314 914
rect 208 800 210 840
rect 312 800 314 840
rect 242 766 280 790
rect 208 755 314 766
rect 208 726 210 755
rect 244 721 278 755
rect 312 726 314 755
rect 242 692 280 721
rect 208 686 314 692
rect 208 652 210 686
rect 244 652 278 686
rect 312 652 314 686
rect 242 618 280 652
rect 208 617 314 618
rect 208 583 210 617
rect 244 583 278 617
rect 312 583 314 617
rect 208 578 314 583
rect 242 548 280 578
rect 208 514 210 544
rect 244 514 278 548
rect 312 514 314 544
rect 208 504 314 514
rect 242 479 280 504
rect 208 445 210 470
rect 244 445 278 479
rect 312 445 314 470
rect 208 430 314 445
rect 242 410 280 430
rect 208 376 210 396
rect 244 376 278 410
rect 312 376 314 396
rect 208 356 314 376
rect 242 341 280 356
rect 208 307 210 322
rect 244 307 278 341
rect 312 307 314 322
rect 208 282 314 307
rect 242 272 280 282
rect 208 238 210 248
rect 244 238 278 272
rect 312 238 314 248
rect 208 208 314 238
rect 242 203 280 208
rect 208 169 210 174
rect 244 169 278 203
rect 312 169 314 174
rect 208 134 314 169
rect 244 100 278 134
rect 208 0 314 100
rect 620 3000 726 3100
rect 620 2927 622 2966
rect 724 2927 726 2966
rect 620 2854 622 2893
rect 724 2854 726 2893
rect 620 2781 622 2820
rect 724 2781 726 2820
rect 620 2708 622 2747
rect 724 2708 726 2747
rect 620 2635 622 2674
rect 724 2635 726 2674
rect 620 2562 622 2601
rect 724 2562 726 2601
rect 620 2489 622 2528
rect 724 2489 726 2528
rect 620 2416 622 2455
rect 724 2416 726 2455
rect 620 2343 622 2382
rect 724 2343 726 2382
rect 620 2270 622 2309
rect 724 2270 726 2309
rect 620 2197 622 2236
rect 724 2197 726 2236
rect 620 2124 622 2163
rect 724 2124 726 2163
rect 620 2051 622 2090
rect 724 2051 726 2090
rect 620 1978 622 2017
rect 724 1978 726 2017
rect 620 1905 622 1944
rect 724 1905 726 1944
rect 620 1832 622 1871
rect 724 1832 726 1871
rect 620 1759 622 1798
rect 724 1759 726 1798
rect 620 1686 622 1725
rect 724 1686 726 1725
rect 620 1613 622 1652
rect 724 1613 726 1652
rect 620 1540 622 1579
rect 724 1540 726 1579
rect 620 1466 622 1506
rect 724 1466 726 1506
rect 620 1392 622 1432
rect 724 1392 726 1432
rect 620 1318 622 1358
rect 724 1318 726 1358
rect 620 1244 622 1284
rect 724 1244 726 1284
rect 620 1170 622 1210
rect 724 1170 726 1210
rect 620 1096 622 1136
rect 724 1096 726 1136
rect 620 1022 622 1062
rect 724 1022 726 1062
rect 620 948 622 988
rect 724 948 726 988
rect 620 874 622 914
rect 724 874 726 914
rect 620 800 622 840
rect 724 800 726 840
rect 654 766 692 790
rect 620 755 726 766
rect 620 726 622 755
rect 656 721 690 755
rect 724 726 726 755
rect 654 692 692 721
rect 620 686 726 692
rect 620 652 622 686
rect 656 652 690 686
rect 724 652 726 686
rect 654 618 692 652
rect 620 617 726 618
rect 620 583 622 617
rect 656 583 690 617
rect 724 583 726 617
rect 620 578 726 583
rect 654 548 692 578
rect 620 514 622 544
rect 656 514 690 548
rect 724 514 726 544
rect 620 504 726 514
rect 654 479 692 504
rect 620 445 622 470
rect 656 445 690 479
rect 724 445 726 470
rect 620 430 726 445
rect 654 410 692 430
rect 620 376 622 396
rect 656 376 690 410
rect 724 376 726 396
rect 620 356 726 376
rect 654 341 692 356
rect 620 307 622 322
rect 656 307 690 341
rect 724 307 726 322
rect 620 282 726 307
rect 654 272 692 282
rect 620 238 622 248
rect 656 238 690 272
rect 724 238 726 248
rect 620 208 726 238
rect 654 203 692 208
rect 620 169 622 174
rect 656 169 690 203
rect 724 169 726 174
rect 620 134 726 169
rect 656 100 690 134
rect 620 0 726 100
rect 1032 3000 1138 3100
rect 1032 2927 1034 2966
rect 1136 2927 1138 2966
rect 1032 2854 1034 2893
rect 1136 2854 1138 2893
rect 1032 2781 1034 2820
rect 1136 2781 1138 2820
rect 1032 2708 1034 2747
rect 1136 2708 1138 2747
rect 1032 2635 1034 2674
rect 1136 2635 1138 2674
rect 1032 2562 1034 2601
rect 1136 2562 1138 2601
rect 1032 2489 1034 2528
rect 1136 2489 1138 2528
rect 1032 2416 1034 2455
rect 1136 2416 1138 2455
rect 1032 2343 1034 2382
rect 1136 2343 1138 2382
rect 1032 2270 1034 2309
rect 1136 2270 1138 2309
rect 1032 2197 1034 2236
rect 1136 2197 1138 2236
rect 1032 2124 1034 2163
rect 1136 2124 1138 2163
rect 1032 2051 1034 2090
rect 1136 2051 1138 2090
rect 1032 1978 1034 2017
rect 1136 1978 1138 2017
rect 1032 1905 1034 1944
rect 1136 1905 1138 1944
rect 1032 1832 1034 1871
rect 1136 1832 1138 1871
rect 1032 1759 1034 1798
rect 1136 1759 1138 1798
rect 1032 1686 1034 1725
rect 1136 1686 1138 1725
rect 1032 1613 1034 1652
rect 1136 1613 1138 1652
rect 1032 1540 1034 1579
rect 1136 1540 1138 1579
rect 1032 1466 1034 1506
rect 1136 1466 1138 1506
rect 1032 1392 1034 1432
rect 1136 1392 1138 1432
rect 1032 1318 1034 1358
rect 1136 1318 1138 1358
rect 1032 1244 1034 1284
rect 1136 1244 1138 1284
rect 1032 1170 1034 1210
rect 1136 1170 1138 1210
rect 1032 1096 1034 1136
rect 1136 1096 1138 1136
rect 1032 1022 1034 1062
rect 1136 1022 1138 1062
rect 1032 948 1034 988
rect 1136 948 1138 988
rect 1032 874 1034 914
rect 1136 874 1138 914
rect 1032 800 1034 840
rect 1136 800 1138 840
rect 1066 766 1104 790
rect 1032 755 1138 766
rect 1032 726 1034 755
rect 1068 721 1102 755
rect 1136 726 1138 755
rect 1066 692 1104 721
rect 1032 686 1138 692
rect 1032 652 1034 686
rect 1068 652 1102 686
rect 1136 652 1138 686
rect 1066 618 1104 652
rect 1032 617 1138 618
rect 1032 583 1034 617
rect 1068 583 1102 617
rect 1136 583 1138 617
rect 1032 578 1138 583
rect 1066 548 1104 578
rect 1032 514 1034 544
rect 1068 514 1102 548
rect 1136 514 1138 544
rect 1032 504 1138 514
rect 1066 479 1104 504
rect 1032 445 1034 470
rect 1068 445 1102 479
rect 1136 445 1138 470
rect 1032 430 1138 445
rect 1066 410 1104 430
rect 1032 376 1034 396
rect 1068 376 1102 410
rect 1136 376 1138 396
rect 1032 356 1138 376
rect 1066 341 1104 356
rect 1032 307 1034 322
rect 1068 307 1102 341
rect 1136 307 1138 322
rect 1032 282 1138 307
rect 1066 272 1104 282
rect 1032 238 1034 248
rect 1068 238 1102 272
rect 1136 238 1138 248
rect 1032 208 1138 238
rect 1066 203 1104 208
rect 1032 169 1034 174
rect 1068 169 1102 203
rect 1136 169 1138 174
rect 1032 134 1138 169
rect 1068 100 1102 134
rect 1032 0 1138 100
rect 1444 3000 1550 3100
rect 1444 2927 1446 2966
rect 1548 2927 1550 2966
rect 1444 2854 1446 2893
rect 1548 2854 1550 2893
rect 1444 2781 1446 2820
rect 1548 2781 1550 2820
rect 1444 2708 1446 2747
rect 1548 2708 1550 2747
rect 1444 2635 1446 2674
rect 1548 2635 1550 2674
rect 1444 2562 1446 2601
rect 1548 2562 1550 2601
rect 1444 2489 1446 2528
rect 1548 2489 1550 2528
rect 1444 2416 1446 2455
rect 1548 2416 1550 2455
rect 1444 2343 1446 2382
rect 1548 2343 1550 2382
rect 1444 2270 1446 2309
rect 1548 2270 1550 2309
rect 1444 2197 1446 2236
rect 1548 2197 1550 2236
rect 1444 2124 1446 2163
rect 1548 2124 1550 2163
rect 1444 2051 1446 2090
rect 1548 2051 1550 2090
rect 1444 1978 1446 2017
rect 1548 1978 1550 2017
rect 1444 1905 1446 1944
rect 1548 1905 1550 1944
rect 1444 1832 1446 1871
rect 1548 1832 1550 1871
rect 1444 1759 1446 1798
rect 1548 1759 1550 1798
rect 1444 1686 1446 1725
rect 1548 1686 1550 1725
rect 1444 1613 1446 1652
rect 1548 1613 1550 1652
rect 1444 1540 1446 1579
rect 1548 1540 1550 1579
rect 1444 1466 1446 1506
rect 1548 1466 1550 1506
rect 1444 1392 1446 1432
rect 1548 1392 1550 1432
rect 1444 1318 1446 1358
rect 1548 1318 1550 1358
rect 1444 1244 1446 1284
rect 1548 1244 1550 1284
rect 1444 1170 1446 1210
rect 1548 1170 1550 1210
rect 1444 1096 1446 1136
rect 1548 1096 1550 1136
rect 1444 1022 1446 1062
rect 1548 1022 1550 1062
rect 1444 948 1446 988
rect 1548 948 1550 988
rect 1444 874 1446 914
rect 1548 874 1550 914
rect 1444 800 1446 840
rect 1548 800 1550 840
rect 1478 766 1516 790
rect 1444 755 1550 766
rect 1444 726 1446 755
rect 1480 721 1514 755
rect 1548 726 1550 755
rect 1478 692 1516 721
rect 1444 686 1550 692
rect 1444 652 1446 686
rect 1480 652 1514 686
rect 1548 652 1550 686
rect 1478 618 1516 652
rect 1444 617 1550 618
rect 1444 583 1446 617
rect 1480 583 1514 617
rect 1548 583 1550 617
rect 1444 578 1550 583
rect 1478 548 1516 578
rect 1444 514 1446 544
rect 1480 514 1514 548
rect 1548 514 1550 544
rect 1444 504 1550 514
rect 1478 479 1516 504
rect 1444 445 1446 470
rect 1480 445 1514 479
rect 1548 445 1550 470
rect 1444 430 1550 445
rect 1478 410 1516 430
rect 1444 376 1446 396
rect 1480 376 1514 410
rect 1548 376 1550 396
rect 1444 356 1550 376
rect 1478 341 1516 356
rect 1444 307 1446 322
rect 1480 307 1514 341
rect 1548 307 1550 322
rect 1444 282 1550 307
rect 1478 272 1516 282
rect 1444 238 1446 248
rect 1480 238 1514 272
rect 1548 238 1550 248
rect 1444 208 1550 238
rect 1478 203 1516 208
rect 1444 169 1446 174
rect 1480 169 1514 203
rect 1548 169 1550 174
rect 1444 134 1550 169
rect 1480 100 1514 134
rect 1444 0 1550 100
rect 1856 3000 1962 3100
rect 1856 2927 1858 2966
rect 1960 2927 1962 2966
rect 1856 2854 1858 2893
rect 1960 2854 1962 2893
rect 1856 2781 1858 2820
rect 1960 2781 1962 2820
rect 1856 2708 1858 2747
rect 1960 2708 1962 2747
rect 1856 2635 1858 2674
rect 1960 2635 1962 2674
rect 1856 2562 1858 2601
rect 1960 2562 1962 2601
rect 1856 2489 1858 2528
rect 1960 2489 1962 2528
rect 1856 2416 1858 2455
rect 1960 2416 1962 2455
rect 1856 2343 1858 2382
rect 1960 2343 1962 2382
rect 1856 2270 1858 2309
rect 1960 2270 1962 2309
rect 1856 2197 1858 2236
rect 1960 2197 1962 2236
rect 1856 2124 1858 2163
rect 1960 2124 1962 2163
rect 1856 2051 1858 2090
rect 1960 2051 1962 2090
rect 1856 1978 1858 2017
rect 1960 1978 1962 2017
rect 1856 1905 1858 1944
rect 1960 1905 1962 1944
rect 1856 1832 1858 1871
rect 1960 1832 1962 1871
rect 1856 1759 1858 1798
rect 1960 1759 1962 1798
rect 1856 1686 1858 1725
rect 1960 1686 1962 1725
rect 1856 1613 1858 1652
rect 1960 1613 1962 1652
rect 1856 1540 1858 1579
rect 1960 1540 1962 1579
rect 1856 1466 1858 1506
rect 1960 1466 1962 1506
rect 1856 1392 1858 1432
rect 1960 1392 1962 1432
rect 1856 1318 1858 1358
rect 1960 1318 1962 1358
rect 1856 1244 1858 1284
rect 1960 1244 1962 1284
rect 1856 1170 1858 1210
rect 1960 1170 1962 1210
rect 1856 1096 1858 1136
rect 1960 1096 1962 1136
rect 1856 1022 1858 1062
rect 1960 1022 1962 1062
rect 1856 948 1858 988
rect 1960 948 1962 988
rect 1856 874 1858 914
rect 1960 874 1962 914
rect 1856 800 1858 840
rect 1960 800 1962 840
rect 1890 766 1928 790
rect 1856 755 1962 766
rect 1856 726 1858 755
rect 1892 721 1926 755
rect 1960 726 1962 755
rect 1890 692 1928 721
rect 1856 686 1962 692
rect 1856 652 1858 686
rect 1892 652 1926 686
rect 1960 652 1962 686
rect 1890 618 1928 652
rect 1856 617 1962 618
rect 1856 583 1858 617
rect 1892 583 1926 617
rect 1960 583 1962 617
rect 1856 578 1962 583
rect 1890 548 1928 578
rect 1856 514 1858 544
rect 1892 514 1926 548
rect 1960 514 1962 544
rect 1856 504 1962 514
rect 1890 479 1928 504
rect 1856 445 1858 470
rect 1892 445 1926 479
rect 1960 445 1962 470
rect 1856 430 1962 445
rect 1890 410 1928 430
rect 1856 376 1858 396
rect 1892 376 1926 410
rect 1960 376 1962 396
rect 1856 356 1962 376
rect 1890 341 1928 356
rect 1856 307 1858 322
rect 1892 307 1926 341
rect 1960 307 1962 322
rect 1856 282 1962 307
rect 1890 272 1928 282
rect 1856 238 1858 248
rect 1892 238 1926 272
rect 1960 238 1962 248
rect 1856 208 1962 238
rect 1890 203 1928 208
rect 1856 169 1858 174
rect 1892 169 1926 203
rect 1960 169 1962 174
rect 1856 134 1962 169
rect 1892 100 1926 134
rect 1856 0 1962 100
rect 2268 3000 2374 3100
rect 2268 2927 2270 2966
rect 2372 2927 2374 2966
rect 2268 2854 2270 2893
rect 2372 2854 2374 2893
rect 2268 2781 2270 2820
rect 2372 2781 2374 2820
rect 2268 2708 2270 2747
rect 2372 2708 2374 2747
rect 2268 2635 2270 2674
rect 2372 2635 2374 2674
rect 2268 2562 2270 2601
rect 2372 2562 2374 2601
rect 2268 2489 2270 2528
rect 2372 2489 2374 2528
rect 2268 2416 2270 2455
rect 2372 2416 2374 2455
rect 2268 2343 2270 2382
rect 2372 2343 2374 2382
rect 2268 2270 2270 2309
rect 2372 2270 2374 2309
rect 2268 2197 2270 2236
rect 2372 2197 2374 2236
rect 2268 2124 2270 2163
rect 2372 2124 2374 2163
rect 2268 2051 2270 2090
rect 2372 2051 2374 2090
rect 2268 1978 2270 2017
rect 2372 1978 2374 2017
rect 2268 1905 2270 1944
rect 2372 1905 2374 1944
rect 2268 1832 2270 1871
rect 2372 1832 2374 1871
rect 2268 1759 2270 1798
rect 2372 1759 2374 1798
rect 2268 1686 2270 1725
rect 2372 1686 2374 1725
rect 2268 1613 2270 1652
rect 2372 1613 2374 1652
rect 2268 1540 2270 1579
rect 2372 1540 2374 1579
rect 2268 1466 2270 1506
rect 2372 1466 2374 1506
rect 2268 1392 2270 1432
rect 2372 1392 2374 1432
rect 2268 1318 2270 1358
rect 2372 1318 2374 1358
rect 2268 1244 2270 1284
rect 2372 1244 2374 1284
rect 2268 1170 2270 1210
rect 2372 1170 2374 1210
rect 2268 1096 2270 1136
rect 2372 1096 2374 1136
rect 2268 1022 2270 1062
rect 2372 1022 2374 1062
rect 2268 948 2270 988
rect 2372 948 2374 988
rect 2268 874 2270 914
rect 2372 874 2374 914
rect 2268 800 2270 840
rect 2372 800 2374 840
rect 2302 766 2340 790
rect 2268 755 2374 766
rect 2268 726 2270 755
rect 2304 721 2338 755
rect 2372 726 2374 755
rect 2302 692 2340 721
rect 2268 686 2374 692
rect 2268 652 2270 686
rect 2304 652 2338 686
rect 2372 652 2374 686
rect 2302 618 2340 652
rect 2268 617 2374 618
rect 2268 583 2270 617
rect 2304 583 2338 617
rect 2372 583 2374 617
rect 2268 578 2374 583
rect 2302 548 2340 578
rect 2268 514 2270 544
rect 2304 514 2338 548
rect 2372 514 2374 544
rect 2268 504 2374 514
rect 2302 479 2340 504
rect 2268 445 2270 470
rect 2304 445 2338 479
rect 2372 445 2374 470
rect 2268 430 2374 445
rect 2302 410 2340 430
rect 2268 376 2270 396
rect 2304 376 2338 410
rect 2372 376 2374 396
rect 2268 356 2374 376
rect 2302 341 2340 356
rect 2268 307 2270 322
rect 2304 307 2338 341
rect 2372 307 2374 322
rect 2268 282 2374 307
rect 2302 272 2340 282
rect 2268 238 2270 248
rect 2304 238 2338 272
rect 2372 238 2374 248
rect 2268 208 2374 238
rect 2302 203 2340 208
rect 2268 169 2270 174
rect 2304 169 2338 203
rect 2372 169 2374 174
rect 2268 134 2374 169
rect 2304 100 2338 134
rect 2268 0 2374 100
rect 2680 3000 2786 3100
rect 2680 2927 2682 2966
rect 2784 2927 2786 2966
rect 2680 2854 2682 2893
rect 2784 2854 2786 2893
rect 2680 2781 2682 2820
rect 2784 2781 2786 2820
rect 2680 2708 2682 2747
rect 2784 2708 2786 2747
rect 2680 2635 2682 2674
rect 2784 2635 2786 2674
rect 2680 2562 2682 2601
rect 2784 2562 2786 2601
rect 2680 2489 2682 2528
rect 2784 2489 2786 2528
rect 2680 2416 2682 2455
rect 2784 2416 2786 2455
rect 2680 2343 2682 2382
rect 2784 2343 2786 2382
rect 2680 2270 2682 2309
rect 2784 2270 2786 2309
rect 2680 2197 2682 2236
rect 2784 2197 2786 2236
rect 2680 2124 2682 2163
rect 2784 2124 2786 2163
rect 2680 2051 2682 2090
rect 2784 2051 2786 2090
rect 2680 1978 2682 2017
rect 2784 1978 2786 2017
rect 2680 1905 2682 1944
rect 2784 1905 2786 1944
rect 2680 1832 2682 1871
rect 2784 1832 2786 1871
rect 2680 1759 2682 1798
rect 2784 1759 2786 1798
rect 2680 1686 2682 1725
rect 2784 1686 2786 1725
rect 2680 1613 2682 1652
rect 2784 1613 2786 1652
rect 2680 1540 2682 1579
rect 2784 1540 2786 1579
rect 2680 1466 2682 1506
rect 2784 1466 2786 1506
rect 2680 1392 2682 1432
rect 2784 1392 2786 1432
rect 2680 1318 2682 1358
rect 2784 1318 2786 1358
rect 2680 1244 2682 1284
rect 2784 1244 2786 1284
rect 2680 1170 2682 1210
rect 2784 1170 2786 1210
rect 2680 1096 2682 1136
rect 2784 1096 2786 1136
rect 2680 1022 2682 1062
rect 2784 1022 2786 1062
rect 2680 948 2682 988
rect 2784 948 2786 988
rect 2680 874 2682 914
rect 2784 874 2786 914
rect 2680 800 2682 840
rect 2784 800 2786 840
rect 2714 766 2752 790
rect 2680 755 2786 766
rect 2680 726 2682 755
rect 2716 721 2750 755
rect 2784 726 2786 755
rect 2714 692 2752 721
rect 2680 686 2786 692
rect 2680 652 2682 686
rect 2716 652 2750 686
rect 2784 652 2786 686
rect 2714 618 2752 652
rect 2680 617 2786 618
rect 2680 583 2682 617
rect 2716 583 2750 617
rect 2784 583 2786 617
rect 2680 578 2786 583
rect 2714 548 2752 578
rect 2680 514 2682 544
rect 2716 514 2750 548
rect 2784 514 2786 544
rect 2680 504 2786 514
rect 2714 479 2752 504
rect 2680 445 2682 470
rect 2716 445 2750 479
rect 2784 445 2786 470
rect 2680 430 2786 445
rect 2714 410 2752 430
rect 2680 376 2682 396
rect 2716 376 2750 410
rect 2784 376 2786 396
rect 2680 356 2786 376
rect 2714 341 2752 356
rect 2680 307 2682 322
rect 2716 307 2750 341
rect 2784 307 2786 322
rect 2680 282 2786 307
rect 2714 272 2752 282
rect 2680 238 2682 248
rect 2716 238 2750 272
rect 2784 238 2786 248
rect 2680 208 2786 238
rect 2714 203 2752 208
rect 2680 169 2682 174
rect 2716 169 2750 203
rect 2784 169 2786 174
rect 2680 134 2786 169
rect 2716 100 2750 134
rect 2680 0 2786 100
rect 3092 3000 3198 3100
rect 3092 2927 3094 2966
rect 3196 2927 3198 2966
rect 3092 2854 3094 2893
rect 3196 2854 3198 2893
rect 3092 2781 3094 2820
rect 3196 2781 3198 2820
rect 3092 2708 3094 2747
rect 3196 2708 3198 2747
rect 3092 2635 3094 2674
rect 3196 2635 3198 2674
rect 3092 2562 3094 2601
rect 3196 2562 3198 2601
rect 3092 2489 3094 2528
rect 3196 2489 3198 2528
rect 3092 2416 3094 2455
rect 3196 2416 3198 2455
rect 3092 2343 3094 2382
rect 3196 2343 3198 2382
rect 3092 2270 3094 2309
rect 3196 2270 3198 2309
rect 3092 2197 3094 2236
rect 3196 2197 3198 2236
rect 3092 2124 3094 2163
rect 3196 2124 3198 2163
rect 3092 2051 3094 2090
rect 3196 2051 3198 2090
rect 3092 1978 3094 2017
rect 3196 1978 3198 2017
rect 3092 1905 3094 1944
rect 3196 1905 3198 1944
rect 3092 1832 3094 1871
rect 3196 1832 3198 1871
rect 3092 1759 3094 1798
rect 3196 1759 3198 1798
rect 3092 1686 3094 1725
rect 3196 1686 3198 1725
rect 3092 1613 3094 1652
rect 3196 1613 3198 1652
rect 3092 1540 3094 1579
rect 3196 1540 3198 1579
rect 3092 1466 3094 1506
rect 3196 1466 3198 1506
rect 3092 1392 3094 1432
rect 3196 1392 3198 1432
rect 3092 1318 3094 1358
rect 3196 1318 3198 1358
rect 3092 1244 3094 1284
rect 3196 1244 3198 1284
rect 3092 1170 3094 1210
rect 3196 1170 3198 1210
rect 3092 1096 3094 1136
rect 3196 1096 3198 1136
rect 3092 1022 3094 1062
rect 3196 1022 3198 1062
rect 3092 948 3094 988
rect 3196 948 3198 988
rect 3092 874 3094 914
rect 3196 874 3198 914
rect 3092 800 3094 840
rect 3196 800 3198 840
rect 3126 766 3164 790
rect 3092 755 3198 766
rect 3092 726 3094 755
rect 3128 721 3162 755
rect 3196 726 3198 755
rect 3126 692 3164 721
rect 3092 686 3198 692
rect 3092 652 3094 686
rect 3128 652 3162 686
rect 3196 652 3198 686
rect 3126 618 3164 652
rect 3092 617 3198 618
rect 3092 583 3094 617
rect 3128 583 3162 617
rect 3196 583 3198 617
rect 3092 578 3198 583
rect 3126 548 3164 578
rect 3092 514 3094 544
rect 3128 514 3162 548
rect 3196 514 3198 544
rect 3092 504 3198 514
rect 3126 479 3164 504
rect 3092 445 3094 470
rect 3128 445 3162 479
rect 3196 445 3198 470
rect 3092 430 3198 445
rect 3126 410 3164 430
rect 3092 376 3094 396
rect 3128 376 3162 410
rect 3196 376 3198 396
rect 3092 356 3198 376
rect 3126 341 3164 356
rect 3092 307 3094 322
rect 3128 307 3162 341
rect 3196 307 3198 322
rect 3092 282 3198 307
rect 3126 272 3164 282
rect 3092 238 3094 248
rect 3128 238 3162 272
rect 3196 238 3198 248
rect 3092 208 3198 238
rect 3126 203 3164 208
rect 3092 169 3094 174
rect 3128 169 3162 203
rect 3196 169 3198 174
rect 3092 134 3198 169
rect 3128 100 3162 134
rect 3092 0 3198 100
rect 3504 3000 3610 3100
rect 3504 2927 3506 2966
rect 3608 2927 3610 2966
rect 3504 2854 3506 2893
rect 3608 2854 3610 2893
rect 3504 2781 3506 2820
rect 3608 2781 3610 2820
rect 3504 2708 3506 2747
rect 3608 2708 3610 2747
rect 3504 2635 3506 2674
rect 3608 2635 3610 2674
rect 3504 2562 3506 2601
rect 3608 2562 3610 2601
rect 3504 2489 3506 2528
rect 3608 2489 3610 2528
rect 3504 2416 3506 2455
rect 3608 2416 3610 2455
rect 3504 2343 3506 2382
rect 3608 2343 3610 2382
rect 3504 2270 3506 2309
rect 3608 2270 3610 2309
rect 3504 2197 3506 2236
rect 3608 2197 3610 2236
rect 3504 2124 3506 2163
rect 3608 2124 3610 2163
rect 3504 2051 3506 2090
rect 3608 2051 3610 2090
rect 3504 1978 3506 2017
rect 3608 1978 3610 2017
rect 3504 1905 3506 1944
rect 3608 1905 3610 1944
rect 3504 1832 3506 1871
rect 3608 1832 3610 1871
rect 3504 1759 3506 1798
rect 3608 1759 3610 1798
rect 3504 1686 3506 1725
rect 3608 1686 3610 1725
rect 3504 1613 3506 1652
rect 3608 1613 3610 1652
rect 3504 1540 3506 1579
rect 3608 1540 3610 1579
rect 3504 1466 3506 1506
rect 3608 1466 3610 1506
rect 3504 1392 3506 1432
rect 3608 1392 3610 1432
rect 3504 1318 3506 1358
rect 3608 1318 3610 1358
rect 3504 1244 3506 1284
rect 3608 1244 3610 1284
rect 3504 1170 3506 1210
rect 3608 1170 3610 1210
rect 3504 1096 3506 1136
rect 3608 1096 3610 1136
rect 3504 1022 3506 1062
rect 3608 1022 3610 1062
rect 3504 948 3506 988
rect 3608 948 3610 988
rect 3504 874 3506 914
rect 3608 874 3610 914
rect 3504 800 3506 840
rect 3608 800 3610 840
rect 3538 766 3576 790
rect 3504 755 3610 766
rect 3504 726 3506 755
rect 3540 721 3574 755
rect 3608 726 3610 755
rect 3538 692 3576 721
rect 3504 686 3610 692
rect 3504 652 3506 686
rect 3540 652 3574 686
rect 3608 652 3610 686
rect 3538 618 3576 652
rect 3504 617 3610 618
rect 3504 583 3506 617
rect 3540 583 3574 617
rect 3608 583 3610 617
rect 3504 578 3610 583
rect 3538 548 3576 578
rect 3504 514 3506 544
rect 3540 514 3574 548
rect 3608 514 3610 544
rect 3504 504 3610 514
rect 3538 479 3576 504
rect 3504 445 3506 470
rect 3540 445 3574 479
rect 3608 445 3610 470
rect 3504 430 3610 445
rect 3538 410 3576 430
rect 3504 376 3506 396
rect 3540 376 3574 410
rect 3608 376 3610 396
rect 3504 356 3610 376
rect 3538 341 3576 356
rect 3504 307 3506 322
rect 3540 307 3574 341
rect 3608 307 3610 322
rect 3504 282 3610 307
rect 3538 272 3576 282
rect 3504 238 3506 248
rect 3540 238 3574 272
rect 3608 238 3610 248
rect 3504 208 3610 238
rect 3538 203 3576 208
rect 3504 169 3506 174
rect 3540 169 3574 203
rect 3608 169 3610 174
rect 3504 134 3610 169
rect 3540 100 3574 134
rect 3504 0 3610 100
rect 3916 3000 4022 3100
rect 3916 2927 3918 2966
rect 4020 2927 4022 2966
rect 3916 2854 3918 2893
rect 4020 2854 4022 2893
rect 3916 2781 3918 2820
rect 4020 2781 4022 2820
rect 3916 2708 3918 2747
rect 4020 2708 4022 2747
rect 3916 2635 3918 2674
rect 4020 2635 4022 2674
rect 3916 2562 3918 2601
rect 4020 2562 4022 2601
rect 3916 2489 3918 2528
rect 4020 2489 4022 2528
rect 3916 2416 3918 2455
rect 4020 2416 4022 2455
rect 3916 2343 3918 2382
rect 4020 2343 4022 2382
rect 3916 2270 3918 2309
rect 4020 2270 4022 2309
rect 3916 2197 3918 2236
rect 4020 2197 4022 2236
rect 3916 2124 3918 2163
rect 4020 2124 4022 2163
rect 3916 2051 3918 2090
rect 4020 2051 4022 2090
rect 3916 1978 3918 2017
rect 4020 1978 4022 2017
rect 3916 1905 3918 1944
rect 4020 1905 4022 1944
rect 3916 1832 3918 1871
rect 4020 1832 4022 1871
rect 3916 1759 3918 1798
rect 4020 1759 4022 1798
rect 3916 1686 3918 1725
rect 4020 1686 4022 1725
rect 3916 1613 3918 1652
rect 4020 1613 4022 1652
rect 3916 1540 3918 1579
rect 4020 1540 4022 1579
rect 3916 1466 3918 1506
rect 4020 1466 4022 1506
rect 3916 1392 3918 1432
rect 4020 1392 4022 1432
rect 3916 1318 3918 1358
rect 4020 1318 4022 1358
rect 3916 1244 3918 1284
rect 4020 1244 4022 1284
rect 3916 1170 3918 1210
rect 4020 1170 4022 1210
rect 3916 1096 3918 1136
rect 4020 1096 4022 1136
rect 3916 1022 3918 1062
rect 4020 1022 4022 1062
rect 3916 948 3918 988
rect 4020 948 4022 988
rect 3916 874 3918 914
rect 4020 874 4022 914
rect 3916 800 3918 840
rect 4020 800 4022 840
rect 3950 766 3988 790
rect 3916 755 4022 766
rect 3916 726 3918 755
rect 3952 721 3986 755
rect 4020 726 4022 755
rect 3950 692 3988 721
rect 3916 686 4022 692
rect 3916 652 3918 686
rect 3952 652 3986 686
rect 4020 652 4022 686
rect 3950 618 3988 652
rect 3916 617 4022 618
rect 3916 583 3918 617
rect 3952 583 3986 617
rect 4020 583 4022 617
rect 3916 578 4022 583
rect 3950 548 3988 578
rect 3916 514 3918 544
rect 3952 514 3986 548
rect 4020 514 4022 544
rect 3916 504 4022 514
rect 3950 479 3988 504
rect 3916 445 3918 470
rect 3952 445 3986 479
rect 4020 445 4022 470
rect 3916 430 4022 445
rect 3950 410 3988 430
rect 3916 376 3918 396
rect 3952 376 3986 410
rect 4020 376 4022 396
rect 3916 356 4022 376
rect 3950 341 3988 356
rect 3916 307 3918 322
rect 3952 307 3986 341
rect 4020 307 4022 322
rect 3916 282 4022 307
rect 3950 272 3988 282
rect 3916 238 3918 248
rect 3952 238 3986 272
rect 4020 238 4022 248
rect 3916 208 4022 238
rect 3950 203 3988 208
rect 3916 169 3918 174
rect 3952 169 3986 203
rect 4020 169 4022 174
rect 3916 134 4022 169
rect 3952 100 3986 134
rect 3916 0 4022 100
rect 4328 3000 4434 3100
rect 4328 2927 4330 2966
rect 4432 2927 4434 2966
rect 4328 2854 4330 2893
rect 4432 2854 4434 2893
rect 4328 2781 4330 2820
rect 4432 2781 4434 2820
rect 4328 2708 4330 2747
rect 4432 2708 4434 2747
rect 4328 2635 4330 2674
rect 4432 2635 4434 2674
rect 4328 2562 4330 2601
rect 4432 2562 4434 2601
rect 4328 2489 4330 2528
rect 4432 2489 4434 2528
rect 4328 2416 4330 2455
rect 4432 2416 4434 2455
rect 4328 2343 4330 2382
rect 4432 2343 4434 2382
rect 4328 2270 4330 2309
rect 4432 2270 4434 2309
rect 4328 2197 4330 2236
rect 4432 2197 4434 2236
rect 4328 2124 4330 2163
rect 4432 2124 4434 2163
rect 4328 2051 4330 2090
rect 4432 2051 4434 2090
rect 4328 1978 4330 2017
rect 4432 1978 4434 2017
rect 4328 1905 4330 1944
rect 4432 1905 4434 1944
rect 4328 1832 4330 1871
rect 4432 1832 4434 1871
rect 4328 1759 4330 1798
rect 4432 1759 4434 1798
rect 4328 1686 4330 1725
rect 4432 1686 4434 1725
rect 4328 1613 4330 1652
rect 4432 1613 4434 1652
rect 4328 1540 4330 1579
rect 4432 1540 4434 1579
rect 4328 1466 4330 1506
rect 4432 1466 4434 1506
rect 4328 1392 4330 1432
rect 4432 1392 4434 1432
rect 4328 1318 4330 1358
rect 4432 1318 4434 1358
rect 4328 1244 4330 1284
rect 4432 1244 4434 1284
rect 4328 1170 4330 1210
rect 4432 1170 4434 1210
rect 4328 1096 4330 1136
rect 4432 1096 4434 1136
rect 4328 1022 4330 1062
rect 4432 1022 4434 1062
rect 4328 948 4330 988
rect 4432 948 4434 988
rect 4328 874 4330 914
rect 4432 874 4434 914
rect 4328 800 4330 840
rect 4432 800 4434 840
rect 4362 766 4400 790
rect 4328 755 4434 766
rect 4328 726 4330 755
rect 4364 721 4398 755
rect 4432 726 4434 755
rect 4362 692 4400 721
rect 4328 686 4434 692
rect 4328 652 4330 686
rect 4364 652 4398 686
rect 4432 652 4434 686
rect 4362 618 4400 652
rect 4328 617 4434 618
rect 4328 583 4330 617
rect 4364 583 4398 617
rect 4432 583 4434 617
rect 4328 578 4434 583
rect 4362 548 4400 578
rect 4328 514 4330 544
rect 4364 514 4398 548
rect 4432 514 4434 544
rect 4328 504 4434 514
rect 4362 479 4400 504
rect 4328 445 4330 470
rect 4364 445 4398 479
rect 4432 445 4434 470
rect 4328 430 4434 445
rect 4362 410 4400 430
rect 4328 376 4330 396
rect 4364 376 4398 410
rect 4432 376 4434 396
rect 4328 356 4434 376
rect 4362 341 4400 356
rect 4328 307 4330 322
rect 4364 307 4398 341
rect 4432 307 4434 322
rect 4328 282 4434 307
rect 4362 272 4400 282
rect 4328 238 4330 248
rect 4364 238 4398 272
rect 4432 238 4434 248
rect 4328 208 4434 238
rect 4362 203 4400 208
rect 4328 169 4330 174
rect 4364 169 4398 203
rect 4432 169 4434 174
rect 4328 134 4434 169
rect 4364 100 4398 134
rect 4328 0 4434 100
rect 4740 3000 4846 3100
rect 4740 2927 4742 2966
rect 4844 2927 4846 2966
rect 4740 2854 4742 2893
rect 4844 2854 4846 2893
rect 4740 2781 4742 2820
rect 4844 2781 4846 2820
rect 4740 2708 4742 2747
rect 4844 2708 4846 2747
rect 4740 2635 4742 2674
rect 4844 2635 4846 2674
rect 4740 2562 4742 2601
rect 4844 2562 4846 2601
rect 4740 2489 4742 2528
rect 4844 2489 4846 2528
rect 4740 2416 4742 2455
rect 4844 2416 4846 2455
rect 4740 2343 4742 2382
rect 4844 2343 4846 2382
rect 4740 2270 4742 2309
rect 4844 2270 4846 2309
rect 4740 2197 4742 2236
rect 4844 2197 4846 2236
rect 4740 2124 4742 2163
rect 4844 2124 4846 2163
rect 4740 2051 4742 2090
rect 4844 2051 4846 2090
rect 4740 1978 4742 2017
rect 4844 1978 4846 2017
rect 4740 1905 4742 1944
rect 4844 1905 4846 1944
rect 4740 1832 4742 1871
rect 4844 1832 4846 1871
rect 4740 1759 4742 1798
rect 4844 1759 4846 1798
rect 4740 1686 4742 1725
rect 4844 1686 4846 1725
rect 4740 1613 4742 1652
rect 4844 1613 4846 1652
rect 4740 1540 4742 1579
rect 4844 1540 4846 1579
rect 4740 1466 4742 1506
rect 4844 1466 4846 1506
rect 4740 1392 4742 1432
rect 4844 1392 4846 1432
rect 4740 1318 4742 1358
rect 4844 1318 4846 1358
rect 4740 1244 4742 1284
rect 4844 1244 4846 1284
rect 4740 1170 4742 1210
rect 4844 1170 4846 1210
rect 4740 1096 4742 1136
rect 4844 1096 4846 1136
rect 4740 1022 4742 1062
rect 4844 1022 4846 1062
rect 4740 948 4742 988
rect 4844 948 4846 988
rect 4740 874 4742 914
rect 4844 874 4846 914
rect 4740 800 4742 840
rect 4844 800 4846 840
rect 4774 766 4812 790
rect 4740 755 4846 766
rect 4740 726 4742 755
rect 4776 721 4810 755
rect 4844 726 4846 755
rect 4774 692 4812 721
rect 4740 686 4846 692
rect 4740 652 4742 686
rect 4776 652 4810 686
rect 4844 652 4846 686
rect 4774 618 4812 652
rect 4740 617 4846 618
rect 4740 583 4742 617
rect 4776 583 4810 617
rect 4844 583 4846 617
rect 4740 578 4846 583
rect 4774 548 4812 578
rect 4740 514 4742 544
rect 4776 514 4810 548
rect 4844 514 4846 544
rect 4740 504 4846 514
rect 4774 479 4812 504
rect 4740 445 4742 470
rect 4776 445 4810 479
rect 4844 445 4846 470
rect 4740 430 4846 445
rect 4774 410 4812 430
rect 4740 376 4742 396
rect 4776 376 4810 410
rect 4844 376 4846 396
rect 4740 356 4846 376
rect 4774 341 4812 356
rect 4740 307 4742 322
rect 4776 307 4810 341
rect 4844 307 4846 322
rect 4740 282 4846 307
rect 4774 272 4812 282
rect 4740 238 4742 248
rect 4776 238 4810 272
rect 4844 238 4846 248
rect 4740 208 4846 238
rect 4774 203 4812 208
rect 4740 169 4742 174
rect 4776 169 4810 203
rect 4844 169 4846 174
rect 4740 134 4846 169
rect 4776 100 4810 134
rect 4740 0 4846 100
rect 5152 3000 5258 3100
rect 5152 2927 5154 2966
rect 5256 2927 5258 2966
rect 5152 2854 5154 2893
rect 5256 2854 5258 2893
rect 5152 2781 5154 2820
rect 5256 2781 5258 2820
rect 5152 2708 5154 2747
rect 5256 2708 5258 2747
rect 5152 2635 5154 2674
rect 5256 2635 5258 2674
rect 5152 2562 5154 2601
rect 5256 2562 5258 2601
rect 5152 2489 5154 2528
rect 5256 2489 5258 2528
rect 5152 2416 5154 2455
rect 5256 2416 5258 2455
rect 5152 2343 5154 2382
rect 5256 2343 5258 2382
rect 5152 2270 5154 2309
rect 5256 2270 5258 2309
rect 5152 2197 5154 2236
rect 5256 2197 5258 2236
rect 5152 2124 5154 2163
rect 5256 2124 5258 2163
rect 5152 2051 5154 2090
rect 5256 2051 5258 2090
rect 5152 1978 5154 2017
rect 5256 1978 5258 2017
rect 5152 1905 5154 1944
rect 5256 1905 5258 1944
rect 5152 1832 5154 1871
rect 5256 1832 5258 1871
rect 5152 1759 5154 1798
rect 5256 1759 5258 1798
rect 5152 1686 5154 1725
rect 5256 1686 5258 1725
rect 5152 1613 5154 1652
rect 5256 1613 5258 1652
rect 5152 1540 5154 1579
rect 5256 1540 5258 1579
rect 5152 1466 5154 1506
rect 5256 1466 5258 1506
rect 5152 1392 5154 1432
rect 5256 1392 5258 1432
rect 5152 1318 5154 1358
rect 5256 1318 5258 1358
rect 5152 1244 5154 1284
rect 5256 1244 5258 1284
rect 5152 1170 5154 1210
rect 5256 1170 5258 1210
rect 5152 1096 5154 1136
rect 5256 1096 5258 1136
rect 5152 1022 5154 1062
rect 5256 1022 5258 1062
rect 5152 948 5154 988
rect 5256 948 5258 988
rect 5152 874 5154 914
rect 5256 874 5258 914
rect 5152 800 5154 840
rect 5256 800 5258 840
rect 5186 766 5224 790
rect 5152 755 5258 766
rect 5152 726 5154 755
rect 5188 721 5222 755
rect 5256 726 5258 755
rect 5186 692 5224 721
rect 5152 686 5258 692
rect 5152 652 5154 686
rect 5188 652 5222 686
rect 5256 652 5258 686
rect 5186 618 5224 652
rect 5152 617 5258 618
rect 5152 583 5154 617
rect 5188 583 5222 617
rect 5256 583 5258 617
rect 5152 578 5258 583
rect 5186 548 5224 578
rect 5152 514 5154 544
rect 5188 514 5222 548
rect 5256 514 5258 544
rect 5152 504 5258 514
rect 5186 479 5224 504
rect 5152 445 5154 470
rect 5188 445 5222 479
rect 5256 445 5258 470
rect 5152 430 5258 445
rect 5186 410 5224 430
rect 5152 376 5154 396
rect 5188 376 5222 410
rect 5256 376 5258 396
rect 5152 356 5258 376
rect 5186 341 5224 356
rect 5152 307 5154 322
rect 5188 307 5222 341
rect 5256 307 5258 322
rect 5152 282 5258 307
rect 5186 272 5224 282
rect 5152 238 5154 248
rect 5188 238 5222 272
rect 5256 238 5258 248
rect 5152 208 5258 238
rect 5186 203 5224 208
rect 5152 169 5154 174
rect 5188 169 5222 203
rect 5256 169 5258 174
rect 5152 134 5258 169
rect 5188 100 5222 134
rect 5152 0 5258 100
rect 5564 3000 5670 3100
rect 5564 2927 5566 2966
rect 5668 2927 5670 2966
rect 5564 2854 5566 2893
rect 5668 2854 5670 2893
rect 5564 2781 5566 2820
rect 5668 2781 5670 2820
rect 5564 2708 5566 2747
rect 5668 2708 5670 2747
rect 5564 2635 5566 2674
rect 5668 2635 5670 2674
rect 5564 2562 5566 2601
rect 5668 2562 5670 2601
rect 5564 2489 5566 2528
rect 5668 2489 5670 2528
rect 5564 2416 5566 2455
rect 5668 2416 5670 2455
rect 5564 2343 5566 2382
rect 5668 2343 5670 2382
rect 5564 2270 5566 2309
rect 5668 2270 5670 2309
rect 5564 2197 5566 2236
rect 5668 2197 5670 2236
rect 5564 2124 5566 2163
rect 5668 2124 5670 2163
rect 5564 2051 5566 2090
rect 5668 2051 5670 2090
rect 5564 1978 5566 2017
rect 5668 1978 5670 2017
rect 5564 1905 5566 1944
rect 5668 1905 5670 1944
rect 5564 1832 5566 1871
rect 5668 1832 5670 1871
rect 5564 1759 5566 1798
rect 5668 1759 5670 1798
rect 5564 1686 5566 1725
rect 5668 1686 5670 1725
rect 5564 1613 5566 1652
rect 5668 1613 5670 1652
rect 5564 1540 5566 1579
rect 5668 1540 5670 1579
rect 5564 1466 5566 1506
rect 5668 1466 5670 1506
rect 5564 1392 5566 1432
rect 5668 1392 5670 1432
rect 5564 1318 5566 1358
rect 5668 1318 5670 1358
rect 5564 1244 5566 1284
rect 5668 1244 5670 1284
rect 5564 1170 5566 1210
rect 5668 1170 5670 1210
rect 5564 1096 5566 1136
rect 5668 1096 5670 1136
rect 5564 1022 5566 1062
rect 5668 1022 5670 1062
rect 5564 948 5566 988
rect 5668 948 5670 988
rect 5564 874 5566 914
rect 5668 874 5670 914
rect 5564 800 5566 840
rect 5668 800 5670 840
rect 5598 766 5636 790
rect 5564 755 5670 766
rect 5564 726 5566 755
rect 5600 721 5634 755
rect 5668 726 5670 755
rect 5598 692 5636 721
rect 5564 686 5670 692
rect 5564 652 5566 686
rect 5600 652 5634 686
rect 5668 652 5670 686
rect 5598 618 5636 652
rect 5564 617 5670 618
rect 5564 583 5566 617
rect 5600 583 5634 617
rect 5668 583 5670 617
rect 5564 578 5670 583
rect 5598 548 5636 578
rect 5564 514 5566 544
rect 5600 514 5634 548
rect 5668 514 5670 544
rect 5564 504 5670 514
rect 5598 479 5636 504
rect 5564 445 5566 470
rect 5600 445 5634 479
rect 5668 445 5670 470
rect 5564 430 5670 445
rect 5598 410 5636 430
rect 5564 376 5566 396
rect 5600 376 5634 410
rect 5668 376 5670 396
rect 5564 356 5670 376
rect 5598 341 5636 356
rect 5564 307 5566 322
rect 5600 307 5634 341
rect 5668 307 5670 322
rect 5564 282 5670 307
rect 5598 272 5636 282
rect 5564 238 5566 248
rect 5600 238 5634 272
rect 5668 238 5670 248
rect 5564 208 5670 238
rect 5598 203 5636 208
rect 5564 169 5566 174
rect 5600 169 5634 203
rect 5668 169 5670 174
rect 5564 134 5670 169
rect 5600 100 5634 134
rect 5564 0 5670 100
rect 5976 3000 6082 3100
rect 5976 2927 5978 2966
rect 6080 2927 6082 2966
rect 5976 2854 5978 2893
rect 6080 2854 6082 2893
rect 5976 2781 5978 2820
rect 6080 2781 6082 2820
rect 5976 2708 5978 2747
rect 6080 2708 6082 2747
rect 5976 2635 5978 2674
rect 6080 2635 6082 2674
rect 5976 2562 5978 2601
rect 6080 2562 6082 2601
rect 5976 2489 5978 2528
rect 6080 2489 6082 2528
rect 5976 2416 5978 2455
rect 6080 2416 6082 2455
rect 5976 2343 5978 2382
rect 6080 2343 6082 2382
rect 5976 2270 5978 2309
rect 6080 2270 6082 2309
rect 5976 2197 5978 2236
rect 6080 2197 6082 2236
rect 5976 2124 5978 2163
rect 6080 2124 6082 2163
rect 5976 2051 5978 2090
rect 6080 2051 6082 2090
rect 5976 1978 5978 2017
rect 6080 1978 6082 2017
rect 5976 1905 5978 1944
rect 6080 1905 6082 1944
rect 5976 1832 5978 1871
rect 6080 1832 6082 1871
rect 5976 1759 5978 1798
rect 6080 1759 6082 1798
rect 5976 1686 5978 1725
rect 6080 1686 6082 1725
rect 5976 1613 5978 1652
rect 6080 1613 6082 1652
rect 5976 1540 5978 1579
rect 6080 1540 6082 1579
rect 5976 1466 5978 1506
rect 6080 1466 6082 1506
rect 5976 1392 5978 1432
rect 6080 1392 6082 1432
rect 5976 1318 5978 1358
rect 6080 1318 6082 1358
rect 5976 1244 5978 1284
rect 6080 1244 6082 1284
rect 5976 1170 5978 1210
rect 6080 1170 6082 1210
rect 5976 1096 5978 1136
rect 6080 1096 6082 1136
rect 5976 1022 5978 1062
rect 6080 1022 6082 1062
rect 5976 948 5978 988
rect 6080 948 6082 988
rect 5976 874 5978 914
rect 6080 874 6082 914
rect 5976 800 5978 840
rect 6080 800 6082 840
rect 6010 766 6048 790
rect 5976 755 6082 766
rect 5976 726 5978 755
rect 6012 721 6046 755
rect 6080 726 6082 755
rect 6010 692 6048 721
rect 5976 686 6082 692
rect 5976 652 5978 686
rect 6012 652 6046 686
rect 6080 652 6082 686
rect 6010 618 6048 652
rect 5976 617 6082 618
rect 5976 583 5978 617
rect 6012 583 6046 617
rect 6080 583 6082 617
rect 5976 578 6082 583
rect 6010 548 6048 578
rect 5976 514 5978 544
rect 6012 514 6046 548
rect 6080 514 6082 544
rect 5976 504 6082 514
rect 6010 479 6048 504
rect 5976 445 5978 470
rect 6012 445 6046 479
rect 6080 445 6082 470
rect 5976 430 6082 445
rect 6010 410 6048 430
rect 5976 376 5978 396
rect 6012 376 6046 410
rect 6080 376 6082 396
rect 5976 356 6082 376
rect 6010 341 6048 356
rect 5976 307 5978 322
rect 6012 307 6046 341
rect 6080 307 6082 322
rect 5976 282 6082 307
rect 6010 272 6048 282
rect 5976 238 5978 248
rect 6012 238 6046 272
rect 6080 238 6082 248
rect 5976 208 6082 238
rect 6010 203 6048 208
rect 5976 169 5978 174
rect 6012 169 6046 203
rect 6080 169 6082 174
rect 5976 134 6082 169
rect 6012 100 6046 134
rect 5976 0 6082 100
rect 6388 3000 6494 3100
rect 6388 2927 6390 2966
rect 6492 2927 6494 2966
rect 6388 2854 6390 2893
rect 6492 2854 6494 2893
rect 6388 2781 6390 2820
rect 6492 2781 6494 2820
rect 6388 2708 6390 2747
rect 6492 2708 6494 2747
rect 6388 2635 6390 2674
rect 6492 2635 6494 2674
rect 6388 2562 6390 2601
rect 6492 2562 6494 2601
rect 6388 2489 6390 2528
rect 6492 2489 6494 2528
rect 6388 2416 6390 2455
rect 6492 2416 6494 2455
rect 6388 2343 6390 2382
rect 6492 2343 6494 2382
rect 6388 2270 6390 2309
rect 6492 2270 6494 2309
rect 6388 2197 6390 2236
rect 6492 2197 6494 2236
rect 6388 2124 6390 2163
rect 6492 2124 6494 2163
rect 6388 2051 6390 2090
rect 6492 2051 6494 2090
rect 6388 1978 6390 2017
rect 6492 1978 6494 2017
rect 6388 1905 6390 1944
rect 6492 1905 6494 1944
rect 6388 1832 6390 1871
rect 6492 1832 6494 1871
rect 6388 1759 6390 1798
rect 6492 1759 6494 1798
rect 6388 1686 6390 1725
rect 6492 1686 6494 1725
rect 6388 1613 6390 1652
rect 6492 1613 6494 1652
rect 6388 1540 6390 1579
rect 6492 1540 6494 1579
rect 6388 1466 6390 1506
rect 6492 1466 6494 1506
rect 6388 1392 6390 1432
rect 6492 1392 6494 1432
rect 6388 1318 6390 1358
rect 6492 1318 6494 1358
rect 6388 1244 6390 1284
rect 6492 1244 6494 1284
rect 6388 1170 6390 1210
rect 6492 1170 6494 1210
rect 6388 1096 6390 1136
rect 6492 1096 6494 1136
rect 6388 1022 6390 1062
rect 6492 1022 6494 1062
rect 6388 948 6390 988
rect 6492 948 6494 988
rect 6388 874 6390 914
rect 6492 874 6494 914
rect 6388 800 6390 840
rect 6492 800 6494 840
rect 6422 766 6460 790
rect 6388 755 6494 766
rect 6388 726 6390 755
rect 6424 721 6458 755
rect 6492 726 6494 755
rect 6422 692 6460 721
rect 6388 686 6494 692
rect 6388 652 6390 686
rect 6424 652 6458 686
rect 6492 652 6494 686
rect 6422 618 6460 652
rect 6388 617 6494 618
rect 6388 583 6390 617
rect 6424 583 6458 617
rect 6492 583 6494 617
rect 6388 578 6494 583
rect 6422 548 6460 578
rect 6388 514 6390 544
rect 6424 514 6458 548
rect 6492 514 6494 544
rect 6388 504 6494 514
rect 6422 479 6460 504
rect 6388 445 6390 470
rect 6424 445 6458 479
rect 6492 445 6494 470
rect 6388 430 6494 445
rect 6422 410 6460 430
rect 6388 376 6390 396
rect 6424 376 6458 410
rect 6492 376 6494 396
rect 6388 356 6494 376
rect 6422 341 6460 356
rect 6388 307 6390 322
rect 6424 307 6458 341
rect 6492 307 6494 322
rect 6388 282 6494 307
rect 6422 272 6460 282
rect 6388 238 6390 248
rect 6424 238 6458 272
rect 6492 238 6494 248
rect 6388 208 6494 238
rect 6422 203 6460 208
rect 6388 169 6390 174
rect 6424 169 6458 203
rect 6492 169 6494 174
rect 6388 134 6494 169
rect 6424 100 6458 134
rect 6388 0 6494 100
rect 6800 3000 6906 3100
rect 6800 2927 6802 2966
rect 6904 2927 6906 2966
rect 6800 2854 6802 2893
rect 6904 2854 6906 2893
rect 6800 2781 6802 2820
rect 6904 2781 6906 2820
rect 6800 2708 6802 2747
rect 6904 2708 6906 2747
rect 6800 2635 6802 2674
rect 6904 2635 6906 2674
rect 6800 2562 6802 2601
rect 6904 2562 6906 2601
rect 6800 2489 6802 2528
rect 6904 2489 6906 2528
rect 6800 2416 6802 2455
rect 6904 2416 6906 2455
rect 6800 2343 6802 2382
rect 6904 2343 6906 2382
rect 6800 2270 6802 2309
rect 6904 2270 6906 2309
rect 6800 2197 6802 2236
rect 6904 2197 6906 2236
rect 6800 2124 6802 2163
rect 6904 2124 6906 2163
rect 6800 2051 6802 2090
rect 6904 2051 6906 2090
rect 6800 1978 6802 2017
rect 6904 1978 6906 2017
rect 6800 1905 6802 1944
rect 6904 1905 6906 1944
rect 6800 1832 6802 1871
rect 6904 1832 6906 1871
rect 6800 1759 6802 1798
rect 6904 1759 6906 1798
rect 6800 1686 6802 1725
rect 6904 1686 6906 1725
rect 6800 1613 6802 1652
rect 6904 1613 6906 1652
rect 6800 1540 6802 1579
rect 6904 1540 6906 1579
rect 6800 1466 6802 1506
rect 6904 1466 6906 1506
rect 6800 1392 6802 1432
rect 6904 1392 6906 1432
rect 6800 1318 6802 1358
rect 6904 1318 6906 1358
rect 6800 1244 6802 1284
rect 6904 1244 6906 1284
rect 6800 1170 6802 1210
rect 6904 1170 6906 1210
rect 6800 1096 6802 1136
rect 6904 1096 6906 1136
rect 6800 1022 6802 1062
rect 6904 1022 6906 1062
rect 6800 948 6802 988
rect 6904 948 6906 988
rect 6800 874 6802 914
rect 6904 874 6906 914
rect 6800 800 6802 840
rect 6904 800 6906 840
rect 6834 766 6872 790
rect 6800 755 6906 766
rect 6800 726 6802 755
rect 6836 721 6870 755
rect 6904 726 6906 755
rect 6834 692 6872 721
rect 6800 686 6906 692
rect 6800 652 6802 686
rect 6836 652 6870 686
rect 6904 652 6906 686
rect 6834 618 6872 652
rect 6800 617 6906 618
rect 6800 583 6802 617
rect 6836 583 6870 617
rect 6904 583 6906 617
rect 6800 578 6906 583
rect 6834 548 6872 578
rect 6800 514 6802 544
rect 6836 514 6870 548
rect 6904 514 6906 544
rect 6800 504 6906 514
rect 6834 479 6872 504
rect 6800 445 6802 470
rect 6836 445 6870 479
rect 6904 445 6906 470
rect 6800 430 6906 445
rect 6834 410 6872 430
rect 6800 376 6802 396
rect 6836 376 6870 410
rect 6904 376 6906 396
rect 6800 356 6906 376
rect 6834 341 6872 356
rect 6800 307 6802 322
rect 6836 307 6870 341
rect 6904 307 6906 322
rect 6800 282 6906 307
rect 6834 272 6872 282
rect 6800 238 6802 248
rect 6836 238 6870 272
rect 6904 238 6906 248
rect 6800 208 6906 238
rect 6834 203 6872 208
rect 6800 169 6802 174
rect 6836 169 6870 203
rect 6904 169 6906 174
rect 6800 134 6906 169
rect 6836 100 6870 134
rect 6800 0 6906 100
rect 7212 3000 7318 3100
rect 7212 2927 7214 2966
rect 7316 2927 7318 2966
rect 7212 2854 7214 2893
rect 7316 2854 7318 2893
rect 7212 2781 7214 2820
rect 7316 2781 7318 2820
rect 7212 2708 7214 2747
rect 7316 2708 7318 2747
rect 7212 2635 7214 2674
rect 7316 2635 7318 2674
rect 7212 2562 7214 2601
rect 7316 2562 7318 2601
rect 7212 2489 7214 2528
rect 7316 2489 7318 2528
rect 7212 2416 7214 2455
rect 7316 2416 7318 2455
rect 7212 2343 7214 2382
rect 7316 2343 7318 2382
rect 7212 2270 7214 2309
rect 7316 2270 7318 2309
rect 7212 2197 7214 2236
rect 7316 2197 7318 2236
rect 7212 2124 7214 2163
rect 7316 2124 7318 2163
rect 7212 2051 7214 2090
rect 7316 2051 7318 2090
rect 7212 1978 7214 2017
rect 7316 1978 7318 2017
rect 7212 1905 7214 1944
rect 7316 1905 7318 1944
rect 7212 1832 7214 1871
rect 7316 1832 7318 1871
rect 7212 1759 7214 1798
rect 7316 1759 7318 1798
rect 7212 1686 7214 1725
rect 7316 1686 7318 1725
rect 7212 1613 7214 1652
rect 7316 1613 7318 1652
rect 7212 1540 7214 1579
rect 7316 1540 7318 1579
rect 7212 1466 7214 1506
rect 7316 1466 7318 1506
rect 7212 1392 7214 1432
rect 7316 1392 7318 1432
rect 7212 1318 7214 1358
rect 7316 1318 7318 1358
rect 7212 1244 7214 1284
rect 7316 1244 7318 1284
rect 7212 1170 7214 1210
rect 7316 1170 7318 1210
rect 7212 1096 7214 1136
rect 7316 1096 7318 1136
rect 7212 1022 7214 1062
rect 7316 1022 7318 1062
rect 7212 948 7214 988
rect 7316 948 7318 988
rect 7212 874 7214 914
rect 7316 874 7318 914
rect 7212 800 7214 840
rect 7316 800 7318 840
rect 7246 766 7284 790
rect 7212 755 7318 766
rect 7212 726 7214 755
rect 7248 721 7282 755
rect 7316 726 7318 755
rect 7246 692 7284 721
rect 7212 686 7318 692
rect 7212 652 7214 686
rect 7248 652 7282 686
rect 7316 652 7318 686
rect 7246 618 7284 652
rect 7212 617 7318 618
rect 7212 583 7214 617
rect 7248 583 7282 617
rect 7316 583 7318 617
rect 7212 578 7318 583
rect 7246 548 7284 578
rect 7212 514 7214 544
rect 7248 514 7282 548
rect 7316 514 7318 544
rect 7212 504 7318 514
rect 7246 479 7284 504
rect 7212 445 7214 470
rect 7248 445 7282 479
rect 7316 445 7318 470
rect 7212 430 7318 445
rect 7246 410 7284 430
rect 7212 376 7214 396
rect 7248 376 7282 410
rect 7316 376 7318 396
rect 7212 356 7318 376
rect 7246 341 7284 356
rect 7212 307 7214 322
rect 7248 307 7282 341
rect 7316 307 7318 322
rect 7212 282 7318 307
rect 7246 272 7284 282
rect 7212 238 7214 248
rect 7248 238 7282 272
rect 7316 238 7318 248
rect 7212 208 7318 238
rect 7246 203 7284 208
rect 7212 169 7214 174
rect 7248 169 7282 203
rect 7316 169 7318 174
rect 7212 134 7318 169
rect 7248 100 7282 134
rect 7212 0 7318 100
rect 7624 3000 7730 3100
rect 7624 2927 7626 2966
rect 7728 2927 7730 2966
rect 7624 2854 7626 2893
rect 7728 2854 7730 2893
rect 7624 2781 7626 2820
rect 7728 2781 7730 2820
rect 7624 2708 7626 2747
rect 7728 2708 7730 2747
rect 7624 2635 7626 2674
rect 7728 2635 7730 2674
rect 7624 2562 7626 2601
rect 7728 2562 7730 2601
rect 7624 2489 7626 2528
rect 7728 2489 7730 2528
rect 7624 2416 7626 2455
rect 7728 2416 7730 2455
rect 7624 2343 7626 2382
rect 7728 2343 7730 2382
rect 7624 2270 7626 2309
rect 7728 2270 7730 2309
rect 7624 2197 7626 2236
rect 7728 2197 7730 2236
rect 7624 2124 7626 2163
rect 7728 2124 7730 2163
rect 7624 2051 7626 2090
rect 7728 2051 7730 2090
rect 7624 1978 7626 2017
rect 7728 1978 7730 2017
rect 7624 1905 7626 1944
rect 7728 1905 7730 1944
rect 7624 1832 7626 1871
rect 7728 1832 7730 1871
rect 7624 1759 7626 1798
rect 7728 1759 7730 1798
rect 7624 1686 7626 1725
rect 7728 1686 7730 1725
rect 7624 1613 7626 1652
rect 7728 1613 7730 1652
rect 7624 1540 7626 1579
rect 7728 1540 7730 1579
rect 7624 1466 7626 1506
rect 7728 1466 7730 1506
rect 7624 1392 7626 1432
rect 7728 1392 7730 1432
rect 7624 1318 7626 1358
rect 7728 1318 7730 1358
rect 7624 1244 7626 1284
rect 7728 1244 7730 1284
rect 7624 1170 7626 1210
rect 7728 1170 7730 1210
rect 7624 1096 7626 1136
rect 7728 1096 7730 1136
rect 7624 1022 7626 1062
rect 7728 1022 7730 1062
rect 7624 948 7626 988
rect 7728 948 7730 988
rect 7624 874 7626 914
rect 7728 874 7730 914
rect 7624 800 7626 840
rect 7728 800 7730 840
rect 7658 766 7696 790
rect 7624 755 7730 766
rect 7624 726 7626 755
rect 7660 721 7694 755
rect 7728 726 7730 755
rect 7658 692 7696 721
rect 7624 686 7730 692
rect 7624 652 7626 686
rect 7660 652 7694 686
rect 7728 652 7730 686
rect 7658 618 7696 652
rect 7624 617 7730 618
rect 7624 583 7626 617
rect 7660 583 7694 617
rect 7728 583 7730 617
rect 7624 578 7730 583
rect 7658 548 7696 578
rect 7624 514 7626 544
rect 7660 514 7694 548
rect 7728 514 7730 544
rect 7624 504 7730 514
rect 7658 479 7696 504
rect 7624 445 7626 470
rect 7660 445 7694 479
rect 7728 445 7730 470
rect 7624 430 7730 445
rect 7658 410 7696 430
rect 7624 376 7626 396
rect 7660 376 7694 410
rect 7728 376 7730 396
rect 7624 356 7730 376
rect 7658 341 7696 356
rect 7624 307 7626 322
rect 7660 307 7694 341
rect 7728 307 7730 322
rect 7624 282 7730 307
rect 7658 272 7696 282
rect 7624 238 7626 248
rect 7660 238 7694 272
rect 7728 238 7730 248
rect 7624 208 7730 238
rect 7658 203 7696 208
rect 7624 169 7626 174
rect 7660 169 7694 203
rect 7728 169 7730 174
rect 7624 134 7730 169
rect 7660 100 7694 134
rect 7624 0 7730 100
rect 8036 3000 8142 3100
rect 8036 2927 8038 2966
rect 8140 2927 8142 2966
rect 8036 2854 8038 2893
rect 8140 2854 8142 2893
rect 8036 2781 8038 2820
rect 8140 2781 8142 2820
rect 8036 2708 8038 2747
rect 8140 2708 8142 2747
rect 8036 2635 8038 2674
rect 8140 2635 8142 2674
rect 8036 2562 8038 2601
rect 8140 2562 8142 2601
rect 8036 2489 8038 2528
rect 8140 2489 8142 2528
rect 8036 2416 8038 2455
rect 8140 2416 8142 2455
rect 8036 2343 8038 2382
rect 8140 2343 8142 2382
rect 8036 2270 8038 2309
rect 8140 2270 8142 2309
rect 8036 2197 8038 2236
rect 8140 2197 8142 2236
rect 8036 2124 8038 2163
rect 8140 2124 8142 2163
rect 8036 2051 8038 2090
rect 8140 2051 8142 2090
rect 8036 1978 8038 2017
rect 8140 1978 8142 2017
rect 8036 1905 8038 1944
rect 8140 1905 8142 1944
rect 8036 1832 8038 1871
rect 8140 1832 8142 1871
rect 8036 1759 8038 1798
rect 8140 1759 8142 1798
rect 8036 1686 8038 1725
rect 8140 1686 8142 1725
rect 8036 1613 8038 1652
rect 8140 1613 8142 1652
rect 8036 1540 8038 1579
rect 8140 1540 8142 1579
rect 8036 1466 8038 1506
rect 8140 1466 8142 1506
rect 8036 1392 8038 1432
rect 8140 1392 8142 1432
rect 8036 1318 8038 1358
rect 8140 1318 8142 1358
rect 8036 1244 8038 1284
rect 8140 1244 8142 1284
rect 8036 1170 8038 1210
rect 8140 1170 8142 1210
rect 8036 1096 8038 1136
rect 8140 1096 8142 1136
rect 8036 1022 8038 1062
rect 8140 1022 8142 1062
rect 8036 948 8038 988
rect 8140 948 8142 988
rect 8036 874 8038 914
rect 8140 874 8142 914
rect 8036 800 8038 840
rect 8140 800 8142 840
rect 8070 766 8108 790
rect 8036 755 8142 766
rect 8036 726 8038 755
rect 8072 721 8106 755
rect 8140 726 8142 755
rect 8070 692 8108 721
rect 8036 686 8142 692
rect 8036 652 8038 686
rect 8072 652 8106 686
rect 8140 652 8142 686
rect 8070 618 8108 652
rect 8036 617 8142 618
rect 8036 583 8038 617
rect 8072 583 8106 617
rect 8140 583 8142 617
rect 8036 578 8142 583
rect 8070 548 8108 578
rect 8036 514 8038 544
rect 8072 514 8106 548
rect 8140 514 8142 544
rect 8036 504 8142 514
rect 8070 479 8108 504
rect 8036 445 8038 470
rect 8072 445 8106 479
rect 8140 445 8142 470
rect 8036 430 8142 445
rect 8070 410 8108 430
rect 8036 376 8038 396
rect 8072 376 8106 410
rect 8140 376 8142 396
rect 8036 356 8142 376
rect 8070 341 8108 356
rect 8036 307 8038 322
rect 8072 307 8106 341
rect 8140 307 8142 322
rect 8036 282 8142 307
rect 8070 272 8108 282
rect 8036 238 8038 248
rect 8072 238 8106 272
rect 8140 238 8142 248
rect 8036 208 8142 238
rect 8070 203 8108 208
rect 8036 169 8038 174
rect 8072 169 8106 203
rect 8140 169 8142 174
rect 8036 134 8142 169
rect 8072 100 8106 134
rect 8036 0 8142 100
rect 8448 3000 8554 3100
rect 8448 2927 8450 2966
rect 8552 2927 8554 2966
rect 8448 2854 8450 2893
rect 8552 2854 8554 2893
rect 8448 2781 8450 2820
rect 8552 2781 8554 2820
rect 8448 2708 8450 2747
rect 8552 2708 8554 2747
rect 8448 2635 8450 2674
rect 8552 2635 8554 2674
rect 8448 2562 8450 2601
rect 8552 2562 8554 2601
rect 8448 2489 8450 2528
rect 8552 2489 8554 2528
rect 8448 2416 8450 2455
rect 8552 2416 8554 2455
rect 8448 2343 8450 2382
rect 8552 2343 8554 2382
rect 8448 2270 8450 2309
rect 8552 2270 8554 2309
rect 8448 2197 8450 2236
rect 8552 2197 8554 2236
rect 8448 2124 8450 2163
rect 8552 2124 8554 2163
rect 8448 2051 8450 2090
rect 8552 2051 8554 2090
rect 8448 1978 8450 2017
rect 8552 1978 8554 2017
rect 8448 1905 8450 1944
rect 8552 1905 8554 1944
rect 8448 1832 8450 1871
rect 8552 1832 8554 1871
rect 8448 1759 8450 1798
rect 8552 1759 8554 1798
rect 8448 1686 8450 1725
rect 8552 1686 8554 1725
rect 8448 1613 8450 1652
rect 8552 1613 8554 1652
rect 8448 1540 8450 1579
rect 8552 1540 8554 1579
rect 8448 1466 8450 1506
rect 8552 1466 8554 1506
rect 8448 1392 8450 1432
rect 8552 1392 8554 1432
rect 8448 1318 8450 1358
rect 8552 1318 8554 1358
rect 8448 1244 8450 1284
rect 8552 1244 8554 1284
rect 8448 1170 8450 1210
rect 8552 1170 8554 1210
rect 8448 1096 8450 1136
rect 8552 1096 8554 1136
rect 8448 1022 8450 1062
rect 8552 1022 8554 1062
rect 8448 948 8450 988
rect 8552 948 8554 988
rect 8448 874 8450 914
rect 8552 874 8554 914
rect 8448 800 8450 840
rect 8552 800 8554 840
rect 8482 766 8520 790
rect 8448 755 8554 766
rect 8448 726 8450 755
rect 8484 721 8518 755
rect 8552 726 8554 755
rect 8482 692 8520 721
rect 8448 686 8554 692
rect 8448 652 8450 686
rect 8484 652 8518 686
rect 8552 652 8554 686
rect 8482 618 8520 652
rect 8448 617 8554 618
rect 8448 583 8450 617
rect 8484 583 8518 617
rect 8552 583 8554 617
rect 8448 578 8554 583
rect 8482 548 8520 578
rect 8448 514 8450 544
rect 8484 514 8518 548
rect 8552 514 8554 544
rect 8448 504 8554 514
rect 8482 479 8520 504
rect 8448 445 8450 470
rect 8484 445 8518 479
rect 8552 445 8554 470
rect 8448 430 8554 445
rect 8482 410 8520 430
rect 8448 376 8450 396
rect 8484 376 8518 410
rect 8552 376 8554 396
rect 8448 356 8554 376
rect 8482 341 8520 356
rect 8448 307 8450 322
rect 8484 307 8518 341
rect 8552 307 8554 322
rect 8448 282 8554 307
rect 8482 272 8520 282
rect 8448 238 8450 248
rect 8484 238 8518 272
rect 8552 238 8554 248
rect 8448 208 8554 238
rect 8482 203 8520 208
rect 8448 169 8450 174
rect 8484 169 8518 203
rect 8552 169 8554 174
rect 8448 134 8554 169
rect 8484 100 8518 134
rect 8448 0 8554 100
rect 8860 3000 8966 3100
rect 8860 2927 8862 2966
rect 8964 2927 8966 2966
rect 8860 2854 8862 2893
rect 8964 2854 8966 2893
rect 8860 2781 8862 2820
rect 8964 2781 8966 2820
rect 8860 2708 8862 2747
rect 8964 2708 8966 2747
rect 8860 2635 8862 2674
rect 8964 2635 8966 2674
rect 8860 2562 8862 2601
rect 8964 2562 8966 2601
rect 8860 2489 8862 2528
rect 8964 2489 8966 2528
rect 8860 2416 8862 2455
rect 8964 2416 8966 2455
rect 8860 2343 8862 2382
rect 8964 2343 8966 2382
rect 8860 2270 8862 2309
rect 8964 2270 8966 2309
rect 8860 2197 8862 2236
rect 8964 2197 8966 2236
rect 8860 2124 8862 2163
rect 8964 2124 8966 2163
rect 8860 2051 8862 2090
rect 8964 2051 8966 2090
rect 8860 1978 8862 2017
rect 8964 1978 8966 2017
rect 8860 1905 8862 1944
rect 8964 1905 8966 1944
rect 8860 1832 8862 1871
rect 8964 1832 8966 1871
rect 8860 1759 8862 1798
rect 8964 1759 8966 1798
rect 8860 1686 8862 1725
rect 8964 1686 8966 1725
rect 8860 1613 8862 1652
rect 8964 1613 8966 1652
rect 8860 1540 8862 1579
rect 8964 1540 8966 1579
rect 8860 1466 8862 1506
rect 8964 1466 8966 1506
rect 8860 1392 8862 1432
rect 8964 1392 8966 1432
rect 8860 1318 8862 1358
rect 8964 1318 8966 1358
rect 8860 1244 8862 1284
rect 8964 1244 8966 1284
rect 8860 1170 8862 1210
rect 8964 1170 8966 1210
rect 8860 1096 8862 1136
rect 8964 1096 8966 1136
rect 8860 1022 8862 1062
rect 8964 1022 8966 1062
rect 8860 948 8862 988
rect 8964 948 8966 988
rect 8860 874 8862 914
rect 8964 874 8966 914
rect 8860 800 8862 840
rect 8964 800 8966 840
rect 8894 766 8932 790
rect 8860 755 8966 766
rect 8860 726 8862 755
rect 8896 721 8930 755
rect 8964 726 8966 755
rect 8894 692 8932 721
rect 8860 686 8966 692
rect 8860 652 8862 686
rect 8896 652 8930 686
rect 8964 652 8966 686
rect 8894 618 8932 652
rect 8860 617 8966 618
rect 8860 583 8862 617
rect 8896 583 8930 617
rect 8964 583 8966 617
rect 8860 578 8966 583
rect 8894 548 8932 578
rect 8860 514 8862 544
rect 8896 514 8930 548
rect 8964 514 8966 544
rect 8860 504 8966 514
rect 8894 479 8932 504
rect 8860 445 8862 470
rect 8896 445 8930 479
rect 8964 445 8966 470
rect 8860 430 8966 445
rect 8894 410 8932 430
rect 8860 376 8862 396
rect 8896 376 8930 410
rect 8964 376 8966 396
rect 8860 356 8966 376
rect 8894 341 8932 356
rect 8860 307 8862 322
rect 8896 307 8930 341
rect 8964 307 8966 322
rect 8860 282 8966 307
rect 8894 272 8932 282
rect 8860 238 8862 248
rect 8896 238 8930 272
rect 8964 238 8966 248
rect 8860 208 8966 238
rect 8894 203 8932 208
rect 8860 169 8862 174
rect 8896 169 8930 203
rect 8964 169 8966 174
rect 8860 134 8966 169
rect 8896 100 8930 134
rect 8860 0 8966 100
rect 9272 3000 9378 3100
rect 9272 2927 9274 2966
rect 9376 2927 9378 2966
rect 9272 2854 9274 2893
rect 9376 2854 9378 2893
rect 9272 2781 9274 2820
rect 9376 2781 9378 2820
rect 9272 2708 9274 2747
rect 9376 2708 9378 2747
rect 9272 2635 9274 2674
rect 9376 2635 9378 2674
rect 9272 2562 9274 2601
rect 9376 2562 9378 2601
rect 9272 2489 9274 2528
rect 9376 2489 9378 2528
rect 9272 2416 9274 2455
rect 9376 2416 9378 2455
rect 9272 2343 9274 2382
rect 9376 2343 9378 2382
rect 9272 2270 9274 2309
rect 9376 2270 9378 2309
rect 9272 2197 9274 2236
rect 9376 2197 9378 2236
rect 9272 2124 9274 2163
rect 9376 2124 9378 2163
rect 9272 2051 9274 2090
rect 9376 2051 9378 2090
rect 9272 1978 9274 2017
rect 9376 1978 9378 2017
rect 9272 1905 9274 1944
rect 9376 1905 9378 1944
rect 9272 1832 9274 1871
rect 9376 1832 9378 1871
rect 9272 1759 9274 1798
rect 9376 1759 9378 1798
rect 9272 1686 9274 1725
rect 9376 1686 9378 1725
rect 9272 1613 9274 1652
rect 9376 1613 9378 1652
rect 9272 1540 9274 1579
rect 9376 1540 9378 1579
rect 9272 1466 9274 1506
rect 9376 1466 9378 1506
rect 9272 1392 9274 1432
rect 9376 1392 9378 1432
rect 9272 1318 9274 1358
rect 9376 1318 9378 1358
rect 9272 1244 9274 1284
rect 9376 1244 9378 1284
rect 9272 1170 9274 1210
rect 9376 1170 9378 1210
rect 9272 1096 9274 1136
rect 9376 1096 9378 1136
rect 9272 1022 9274 1062
rect 9376 1022 9378 1062
rect 9272 948 9274 988
rect 9376 948 9378 988
rect 9272 874 9274 914
rect 9376 874 9378 914
rect 9272 800 9274 840
rect 9376 800 9378 840
rect 9306 766 9344 790
rect 9272 755 9378 766
rect 9272 726 9274 755
rect 9308 721 9342 755
rect 9376 726 9378 755
rect 9306 692 9344 721
rect 9272 686 9378 692
rect 9272 652 9274 686
rect 9308 652 9342 686
rect 9376 652 9378 686
rect 9306 618 9344 652
rect 9272 617 9378 618
rect 9272 583 9274 617
rect 9308 583 9342 617
rect 9376 583 9378 617
rect 9272 578 9378 583
rect 9306 548 9344 578
rect 9272 514 9274 544
rect 9308 514 9342 548
rect 9376 514 9378 544
rect 9272 504 9378 514
rect 9306 479 9344 504
rect 9272 445 9274 470
rect 9308 445 9342 479
rect 9376 445 9378 470
rect 9272 430 9378 445
rect 9306 410 9344 430
rect 9272 376 9274 396
rect 9308 376 9342 410
rect 9376 376 9378 396
rect 9272 356 9378 376
rect 9306 341 9344 356
rect 9272 307 9274 322
rect 9308 307 9342 341
rect 9376 307 9378 322
rect 9272 282 9378 307
rect 9306 272 9344 282
rect 9272 238 9274 248
rect 9308 238 9342 272
rect 9376 238 9378 248
rect 9272 208 9378 238
rect 9306 203 9344 208
rect 9272 169 9274 174
rect 9308 169 9342 203
rect 9376 169 9378 174
rect 9272 134 9378 169
rect 9308 100 9342 134
rect 9272 0 9378 100
rect 9684 3000 9790 3100
rect 9684 2927 9686 2966
rect 9788 2927 9790 2966
rect 9684 2854 9686 2893
rect 9788 2854 9790 2893
rect 9684 2781 9686 2820
rect 9788 2781 9790 2820
rect 9684 2708 9686 2747
rect 9788 2708 9790 2747
rect 9684 2635 9686 2674
rect 9788 2635 9790 2674
rect 9684 2562 9686 2601
rect 9788 2562 9790 2601
rect 9684 2489 9686 2528
rect 9788 2489 9790 2528
rect 9684 2416 9686 2455
rect 9788 2416 9790 2455
rect 9684 2343 9686 2382
rect 9788 2343 9790 2382
rect 9684 2270 9686 2309
rect 9788 2270 9790 2309
rect 9684 2197 9686 2236
rect 9788 2197 9790 2236
rect 9684 2124 9686 2163
rect 9788 2124 9790 2163
rect 9684 2051 9686 2090
rect 9788 2051 9790 2090
rect 9684 1978 9686 2017
rect 9788 1978 9790 2017
rect 9684 1905 9686 1944
rect 9788 1905 9790 1944
rect 9684 1832 9686 1871
rect 9788 1832 9790 1871
rect 9684 1759 9686 1798
rect 9788 1759 9790 1798
rect 9684 1686 9686 1725
rect 9788 1686 9790 1725
rect 9684 1613 9686 1652
rect 9788 1613 9790 1652
rect 9684 1540 9686 1579
rect 9788 1540 9790 1579
rect 9684 1466 9686 1506
rect 9788 1466 9790 1506
rect 9684 1392 9686 1432
rect 9788 1392 9790 1432
rect 9684 1318 9686 1358
rect 9788 1318 9790 1358
rect 9684 1244 9686 1284
rect 9788 1244 9790 1284
rect 9684 1170 9686 1210
rect 9788 1170 9790 1210
rect 9684 1096 9686 1136
rect 9788 1096 9790 1136
rect 9684 1022 9686 1062
rect 9788 1022 9790 1062
rect 9684 948 9686 988
rect 9788 948 9790 988
rect 9684 874 9686 914
rect 9788 874 9790 914
rect 9684 800 9686 840
rect 9788 800 9790 840
rect 9718 766 9756 790
rect 9684 755 9790 766
rect 9684 726 9686 755
rect 9720 721 9754 755
rect 9788 726 9790 755
rect 9718 692 9756 721
rect 9684 686 9790 692
rect 9684 652 9686 686
rect 9720 652 9754 686
rect 9788 652 9790 686
rect 9718 618 9756 652
rect 9684 617 9790 618
rect 9684 583 9686 617
rect 9720 583 9754 617
rect 9788 583 9790 617
rect 9684 578 9790 583
rect 9718 548 9756 578
rect 9684 514 9686 544
rect 9720 514 9754 548
rect 9788 514 9790 544
rect 9684 504 9790 514
rect 9718 479 9756 504
rect 9684 445 9686 470
rect 9720 445 9754 479
rect 9788 445 9790 470
rect 9684 430 9790 445
rect 9718 410 9756 430
rect 9684 376 9686 396
rect 9720 376 9754 410
rect 9788 376 9790 396
rect 9684 356 9790 376
rect 9718 341 9756 356
rect 9684 307 9686 322
rect 9720 307 9754 341
rect 9788 307 9790 322
rect 9684 282 9790 307
rect 9718 272 9756 282
rect 9684 238 9686 248
rect 9720 238 9754 272
rect 9788 238 9790 248
rect 9684 208 9790 238
rect 9718 203 9756 208
rect 9684 169 9686 174
rect 9720 169 9754 203
rect 9788 169 9790 174
rect 9684 134 9790 169
rect 9720 100 9754 134
rect 9684 0 9790 100
rect 10096 3000 10202 3100
rect 10096 2927 10098 2966
rect 10200 2927 10202 2966
rect 10096 2854 10098 2893
rect 10200 2854 10202 2893
rect 10096 2781 10098 2820
rect 10200 2781 10202 2820
rect 10096 2708 10098 2747
rect 10200 2708 10202 2747
rect 10096 2635 10098 2674
rect 10200 2635 10202 2674
rect 10096 2562 10098 2601
rect 10200 2562 10202 2601
rect 10096 2489 10098 2528
rect 10200 2489 10202 2528
rect 10096 2416 10098 2455
rect 10200 2416 10202 2455
rect 10096 2343 10098 2382
rect 10200 2343 10202 2382
rect 10096 2270 10098 2309
rect 10200 2270 10202 2309
rect 10096 2197 10098 2236
rect 10200 2197 10202 2236
rect 10096 2124 10098 2163
rect 10200 2124 10202 2163
rect 10096 2051 10098 2090
rect 10200 2051 10202 2090
rect 10096 1978 10098 2017
rect 10200 1978 10202 2017
rect 10096 1905 10098 1944
rect 10200 1905 10202 1944
rect 10096 1832 10098 1871
rect 10200 1832 10202 1871
rect 10096 1759 10098 1798
rect 10200 1759 10202 1798
rect 10096 1686 10098 1725
rect 10200 1686 10202 1725
rect 10096 1613 10098 1652
rect 10200 1613 10202 1652
rect 10096 1540 10098 1579
rect 10200 1540 10202 1579
rect 10096 1466 10098 1506
rect 10200 1466 10202 1506
rect 10096 1392 10098 1432
rect 10200 1392 10202 1432
rect 10096 1318 10098 1358
rect 10200 1318 10202 1358
rect 10096 1244 10098 1284
rect 10200 1244 10202 1284
rect 10096 1170 10098 1210
rect 10200 1170 10202 1210
rect 10096 1096 10098 1136
rect 10200 1096 10202 1136
rect 10096 1022 10098 1062
rect 10200 1022 10202 1062
rect 10096 948 10098 988
rect 10200 948 10202 988
rect 10096 874 10098 914
rect 10200 874 10202 914
rect 10096 800 10098 840
rect 10200 800 10202 840
rect 10130 766 10168 790
rect 10096 755 10202 766
rect 10096 726 10098 755
rect 10132 721 10166 755
rect 10200 726 10202 755
rect 10130 692 10168 721
rect 10096 686 10202 692
rect 10096 652 10098 686
rect 10132 652 10166 686
rect 10200 652 10202 686
rect 10130 618 10168 652
rect 10096 617 10202 618
rect 10096 583 10098 617
rect 10132 583 10166 617
rect 10200 583 10202 617
rect 10096 578 10202 583
rect 10130 548 10168 578
rect 10096 514 10098 544
rect 10132 514 10166 548
rect 10200 514 10202 544
rect 10096 504 10202 514
rect 10130 479 10168 504
rect 10096 445 10098 470
rect 10132 445 10166 479
rect 10200 445 10202 470
rect 10096 430 10202 445
rect 10130 410 10168 430
rect 10096 376 10098 396
rect 10132 376 10166 410
rect 10200 376 10202 396
rect 10096 356 10202 376
rect 10130 341 10168 356
rect 10096 307 10098 322
rect 10132 307 10166 341
rect 10200 307 10202 322
rect 10096 282 10202 307
rect 10130 272 10168 282
rect 10096 238 10098 248
rect 10132 238 10166 272
rect 10200 238 10202 248
rect 10096 208 10202 238
rect 10130 203 10168 208
rect 10096 169 10098 174
rect 10132 169 10166 203
rect 10200 169 10202 174
rect 10096 134 10202 169
rect 10132 100 10166 134
rect 10096 0 10202 100
rect 10508 3000 10614 3100
rect 10508 2927 10510 2966
rect 10612 2927 10614 2966
rect 10508 2854 10510 2893
rect 10612 2854 10614 2893
rect 10508 2781 10510 2820
rect 10612 2781 10614 2820
rect 10508 2708 10510 2747
rect 10612 2708 10614 2747
rect 10508 2635 10510 2674
rect 10612 2635 10614 2674
rect 10508 2562 10510 2601
rect 10612 2562 10614 2601
rect 10508 2489 10510 2528
rect 10612 2489 10614 2528
rect 10508 2416 10510 2455
rect 10612 2416 10614 2455
rect 10508 2343 10510 2382
rect 10612 2343 10614 2382
rect 10508 2270 10510 2309
rect 10612 2270 10614 2309
rect 10508 2197 10510 2236
rect 10612 2197 10614 2236
rect 10508 2124 10510 2163
rect 10612 2124 10614 2163
rect 10508 2051 10510 2090
rect 10612 2051 10614 2090
rect 10508 1978 10510 2017
rect 10612 1978 10614 2017
rect 10508 1905 10510 1944
rect 10612 1905 10614 1944
rect 10508 1832 10510 1871
rect 10612 1832 10614 1871
rect 10508 1759 10510 1798
rect 10612 1759 10614 1798
rect 10508 1686 10510 1725
rect 10612 1686 10614 1725
rect 10508 1613 10510 1652
rect 10612 1613 10614 1652
rect 10508 1540 10510 1579
rect 10612 1540 10614 1579
rect 10508 1466 10510 1506
rect 10612 1466 10614 1506
rect 10508 1392 10510 1432
rect 10612 1392 10614 1432
rect 10508 1318 10510 1358
rect 10612 1318 10614 1358
rect 10508 1244 10510 1284
rect 10612 1244 10614 1284
rect 10508 1170 10510 1210
rect 10612 1170 10614 1210
rect 10508 1096 10510 1136
rect 10612 1096 10614 1136
rect 10508 1022 10510 1062
rect 10612 1022 10614 1062
rect 10508 948 10510 988
rect 10612 948 10614 988
rect 10508 874 10510 914
rect 10612 874 10614 914
rect 10508 800 10510 840
rect 10612 800 10614 840
rect 10542 766 10580 790
rect 10508 755 10614 766
rect 10508 726 10510 755
rect 10544 721 10578 755
rect 10612 726 10614 755
rect 10542 692 10580 721
rect 10508 686 10614 692
rect 10508 652 10510 686
rect 10544 652 10578 686
rect 10612 652 10614 686
rect 10542 618 10580 652
rect 10508 617 10614 618
rect 10508 583 10510 617
rect 10544 583 10578 617
rect 10612 583 10614 617
rect 10508 578 10614 583
rect 10542 548 10580 578
rect 10508 514 10510 544
rect 10544 514 10578 548
rect 10612 514 10614 544
rect 10508 504 10614 514
rect 10542 479 10580 504
rect 10508 445 10510 470
rect 10544 445 10578 479
rect 10612 445 10614 470
rect 10508 430 10614 445
rect 10542 410 10580 430
rect 10508 376 10510 396
rect 10544 376 10578 410
rect 10612 376 10614 396
rect 10508 356 10614 376
rect 10542 341 10580 356
rect 10508 307 10510 322
rect 10544 307 10578 341
rect 10612 307 10614 322
rect 10508 282 10614 307
rect 10542 272 10580 282
rect 10508 238 10510 248
rect 10544 238 10578 272
rect 10612 238 10614 248
rect 10508 208 10614 238
rect 10542 203 10580 208
rect 10508 169 10510 174
rect 10544 169 10578 203
rect 10612 169 10614 174
rect 10508 134 10614 169
rect 10544 100 10578 134
rect 10508 0 10614 100
rect 10920 3000 11026 3100
rect 10920 2927 10922 2966
rect 11024 2927 11026 2966
rect 10920 2854 10922 2893
rect 11024 2854 11026 2893
rect 10920 2781 10922 2820
rect 11024 2781 11026 2820
rect 10920 2708 10922 2747
rect 11024 2708 11026 2747
rect 10920 2635 10922 2674
rect 11024 2635 11026 2674
rect 10920 2562 10922 2601
rect 11024 2562 11026 2601
rect 10920 2489 10922 2528
rect 11024 2489 11026 2528
rect 10920 2416 10922 2455
rect 11024 2416 11026 2455
rect 10920 2343 10922 2382
rect 11024 2343 11026 2382
rect 10920 2270 10922 2309
rect 11024 2270 11026 2309
rect 10920 2197 10922 2236
rect 11024 2197 11026 2236
rect 10920 2124 10922 2163
rect 11024 2124 11026 2163
rect 10920 2051 10922 2090
rect 11024 2051 11026 2090
rect 10920 1978 10922 2017
rect 11024 1978 11026 2017
rect 10920 1905 10922 1944
rect 11024 1905 11026 1944
rect 10920 1832 10922 1871
rect 11024 1832 11026 1871
rect 10920 1759 10922 1798
rect 11024 1759 11026 1798
rect 10920 1686 10922 1725
rect 11024 1686 11026 1725
rect 10920 1613 10922 1652
rect 11024 1613 11026 1652
rect 10920 1540 10922 1579
rect 11024 1540 11026 1579
rect 10920 1466 10922 1506
rect 11024 1466 11026 1506
rect 10920 1392 10922 1432
rect 11024 1392 11026 1432
rect 10920 1318 10922 1358
rect 11024 1318 11026 1358
rect 10920 1244 10922 1284
rect 11024 1244 11026 1284
rect 10920 1170 10922 1210
rect 11024 1170 11026 1210
rect 10920 1096 10922 1136
rect 11024 1096 11026 1136
rect 10920 1022 10922 1062
rect 11024 1022 11026 1062
rect 10920 948 10922 988
rect 11024 948 11026 988
rect 10920 874 10922 914
rect 11024 874 11026 914
rect 10920 800 10922 840
rect 11024 800 11026 840
rect 10954 766 10992 790
rect 10920 755 11026 766
rect 10920 726 10922 755
rect 10956 721 10990 755
rect 11024 726 11026 755
rect 10954 692 10992 721
rect 10920 686 11026 692
rect 10920 652 10922 686
rect 10956 652 10990 686
rect 11024 652 11026 686
rect 10954 618 10992 652
rect 10920 617 11026 618
rect 10920 583 10922 617
rect 10956 583 10990 617
rect 11024 583 11026 617
rect 10920 578 11026 583
rect 10954 548 10992 578
rect 10920 514 10922 544
rect 10956 514 10990 548
rect 11024 514 11026 544
rect 10920 504 11026 514
rect 10954 479 10992 504
rect 10920 445 10922 470
rect 10956 445 10990 479
rect 11024 445 11026 470
rect 10920 430 11026 445
rect 10954 410 10992 430
rect 10920 376 10922 396
rect 10956 376 10990 410
rect 11024 376 11026 396
rect 10920 356 11026 376
rect 10954 341 10992 356
rect 10920 307 10922 322
rect 10956 307 10990 341
rect 11024 307 11026 322
rect 10920 282 11026 307
rect 10954 272 10992 282
rect 10920 238 10922 248
rect 10956 238 10990 272
rect 11024 238 11026 248
rect 10920 208 11026 238
rect 10954 203 10992 208
rect 10920 169 10922 174
rect 10956 169 10990 203
rect 11024 169 11026 174
rect 10920 134 11026 169
rect 10956 100 10990 134
rect 10920 0 11026 100
rect 11332 3000 11438 3100
rect 11332 2927 11334 2966
rect 11436 2927 11438 2966
rect 11332 2854 11334 2893
rect 11436 2854 11438 2893
rect 11332 2781 11334 2820
rect 11436 2781 11438 2820
rect 11332 2708 11334 2747
rect 11436 2708 11438 2747
rect 11332 2635 11334 2674
rect 11436 2635 11438 2674
rect 11332 2562 11334 2601
rect 11436 2562 11438 2601
rect 11332 2489 11334 2528
rect 11436 2489 11438 2528
rect 11332 2416 11334 2455
rect 11436 2416 11438 2455
rect 11332 2343 11334 2382
rect 11436 2343 11438 2382
rect 11332 2270 11334 2309
rect 11436 2270 11438 2309
rect 11332 2197 11334 2236
rect 11436 2197 11438 2236
rect 11332 2124 11334 2163
rect 11436 2124 11438 2163
rect 11332 2051 11334 2090
rect 11436 2051 11438 2090
rect 11332 1978 11334 2017
rect 11436 1978 11438 2017
rect 11332 1905 11334 1944
rect 11436 1905 11438 1944
rect 11332 1832 11334 1871
rect 11436 1832 11438 1871
rect 11332 1759 11334 1798
rect 11436 1759 11438 1798
rect 11332 1686 11334 1725
rect 11436 1686 11438 1725
rect 11332 1613 11334 1652
rect 11436 1613 11438 1652
rect 11332 1540 11334 1579
rect 11436 1540 11438 1579
rect 11332 1466 11334 1506
rect 11436 1466 11438 1506
rect 11332 1392 11334 1432
rect 11436 1392 11438 1432
rect 11332 1318 11334 1358
rect 11436 1318 11438 1358
rect 11332 1244 11334 1284
rect 11436 1244 11438 1284
rect 11332 1170 11334 1210
rect 11436 1170 11438 1210
rect 11332 1096 11334 1136
rect 11436 1096 11438 1136
rect 11332 1022 11334 1062
rect 11436 1022 11438 1062
rect 11332 948 11334 988
rect 11436 948 11438 988
rect 11332 874 11334 914
rect 11436 874 11438 914
rect 11332 800 11334 840
rect 11436 800 11438 840
rect 11366 766 11404 790
rect 11332 755 11438 766
rect 11332 726 11334 755
rect 11368 721 11402 755
rect 11436 726 11438 755
rect 11366 692 11404 721
rect 11332 686 11438 692
rect 11332 652 11334 686
rect 11368 652 11402 686
rect 11436 652 11438 686
rect 11366 618 11404 652
rect 11332 617 11438 618
rect 11332 583 11334 617
rect 11368 583 11402 617
rect 11436 583 11438 617
rect 11332 578 11438 583
rect 11366 548 11404 578
rect 11332 514 11334 544
rect 11368 514 11402 548
rect 11436 514 11438 544
rect 11332 504 11438 514
rect 11366 479 11404 504
rect 11332 445 11334 470
rect 11368 445 11402 479
rect 11436 445 11438 470
rect 11332 430 11438 445
rect 11366 410 11404 430
rect 11332 376 11334 396
rect 11368 376 11402 410
rect 11436 376 11438 396
rect 11332 356 11438 376
rect 11366 341 11404 356
rect 11332 307 11334 322
rect 11368 307 11402 341
rect 11436 307 11438 322
rect 11332 282 11438 307
rect 11366 272 11404 282
rect 11332 238 11334 248
rect 11368 238 11402 272
rect 11436 238 11438 248
rect 11332 208 11438 238
rect 11366 203 11404 208
rect 11332 169 11334 174
rect 11368 169 11402 203
rect 11436 169 11438 174
rect 11332 134 11438 169
rect 11368 100 11402 134
rect 11332 0 11438 100
rect 11744 3000 11850 3100
rect 11744 2927 11746 2966
rect 11848 2927 11850 2966
rect 11744 2854 11746 2893
rect 11848 2854 11850 2893
rect 11744 2781 11746 2820
rect 11848 2781 11850 2820
rect 11744 2708 11746 2747
rect 11848 2708 11850 2747
rect 11744 2635 11746 2674
rect 11848 2635 11850 2674
rect 11744 2562 11746 2601
rect 11848 2562 11850 2601
rect 11744 2489 11746 2528
rect 11848 2489 11850 2528
rect 11744 2416 11746 2455
rect 11848 2416 11850 2455
rect 11744 2343 11746 2382
rect 11848 2343 11850 2382
rect 11744 2270 11746 2309
rect 11848 2270 11850 2309
rect 11744 2197 11746 2236
rect 11848 2197 11850 2236
rect 11744 2124 11746 2163
rect 11848 2124 11850 2163
rect 11744 2051 11746 2090
rect 11848 2051 11850 2090
rect 11744 1978 11746 2017
rect 11848 1978 11850 2017
rect 11744 1905 11746 1944
rect 11848 1905 11850 1944
rect 11744 1832 11746 1871
rect 11848 1832 11850 1871
rect 11744 1759 11746 1798
rect 11848 1759 11850 1798
rect 11744 1686 11746 1725
rect 11848 1686 11850 1725
rect 11744 1613 11746 1652
rect 11848 1613 11850 1652
rect 11744 1540 11746 1579
rect 11848 1540 11850 1579
rect 11744 1466 11746 1506
rect 11848 1466 11850 1506
rect 11744 1392 11746 1432
rect 11848 1392 11850 1432
rect 11744 1318 11746 1358
rect 11848 1318 11850 1358
rect 11744 1244 11746 1284
rect 11848 1244 11850 1284
rect 11744 1170 11746 1210
rect 11848 1170 11850 1210
rect 11744 1096 11746 1136
rect 11848 1096 11850 1136
rect 11744 1022 11746 1062
rect 11848 1022 11850 1062
rect 11744 948 11746 988
rect 11848 948 11850 988
rect 11744 874 11746 914
rect 11848 874 11850 914
rect 11744 800 11746 840
rect 11848 800 11850 840
rect 11778 766 11816 790
rect 11744 755 11850 766
rect 11744 726 11746 755
rect 11780 721 11814 755
rect 11848 726 11850 755
rect 11778 692 11816 721
rect 11744 686 11850 692
rect 11744 652 11746 686
rect 11780 652 11814 686
rect 11848 652 11850 686
rect 11778 618 11816 652
rect 11744 617 11850 618
rect 11744 583 11746 617
rect 11780 583 11814 617
rect 11848 583 11850 617
rect 11744 578 11850 583
rect 11778 548 11816 578
rect 11744 514 11746 544
rect 11780 514 11814 548
rect 11848 514 11850 544
rect 11744 504 11850 514
rect 11778 479 11816 504
rect 11744 445 11746 470
rect 11780 445 11814 479
rect 11848 445 11850 470
rect 11744 430 11850 445
rect 11778 410 11816 430
rect 11744 376 11746 396
rect 11780 376 11814 410
rect 11848 376 11850 396
rect 11744 356 11850 376
rect 11778 341 11816 356
rect 11744 307 11746 322
rect 11780 307 11814 341
rect 11848 307 11850 322
rect 11744 282 11850 307
rect 11778 272 11816 282
rect 11744 238 11746 248
rect 11780 238 11814 272
rect 11848 238 11850 248
rect 11744 208 11850 238
rect 11778 203 11816 208
rect 11744 169 11746 174
rect 11780 169 11814 203
rect 11848 169 11850 174
rect 11744 134 11850 169
rect 11780 100 11814 134
rect 11744 0 11850 100
rect 12156 3000 12262 3100
rect 12156 2927 12158 2966
rect 12260 2927 12262 2966
rect 12156 2854 12158 2893
rect 12260 2854 12262 2893
rect 12156 2781 12158 2820
rect 12260 2781 12262 2820
rect 12156 2708 12158 2747
rect 12260 2708 12262 2747
rect 12156 2635 12158 2674
rect 12260 2635 12262 2674
rect 12156 2562 12158 2601
rect 12260 2562 12262 2601
rect 12156 2489 12158 2528
rect 12260 2489 12262 2528
rect 12156 2416 12158 2455
rect 12260 2416 12262 2455
rect 12156 2343 12158 2382
rect 12260 2343 12262 2382
rect 12156 2270 12158 2309
rect 12260 2270 12262 2309
rect 12156 2197 12158 2236
rect 12260 2197 12262 2236
rect 12156 2124 12158 2163
rect 12260 2124 12262 2163
rect 12156 2051 12158 2090
rect 12260 2051 12262 2090
rect 12156 1978 12158 2017
rect 12260 1978 12262 2017
rect 12156 1905 12158 1944
rect 12260 1905 12262 1944
rect 12156 1832 12158 1871
rect 12260 1832 12262 1871
rect 12156 1759 12158 1798
rect 12260 1759 12262 1798
rect 12156 1686 12158 1725
rect 12260 1686 12262 1725
rect 12156 1613 12158 1652
rect 12260 1613 12262 1652
rect 12156 1540 12158 1579
rect 12260 1540 12262 1579
rect 12156 1466 12158 1506
rect 12260 1466 12262 1506
rect 12156 1392 12158 1432
rect 12260 1392 12262 1432
rect 12156 1318 12158 1358
rect 12260 1318 12262 1358
rect 12156 1244 12158 1284
rect 12260 1244 12262 1284
rect 12156 1170 12158 1210
rect 12260 1170 12262 1210
rect 12156 1096 12158 1136
rect 12260 1096 12262 1136
rect 12156 1022 12158 1062
rect 12260 1022 12262 1062
rect 12156 948 12158 988
rect 12260 948 12262 988
rect 12156 874 12158 914
rect 12260 874 12262 914
rect 12156 800 12158 840
rect 12260 800 12262 840
rect 12190 766 12228 790
rect 12156 755 12262 766
rect 12156 726 12158 755
rect 12192 721 12226 755
rect 12260 726 12262 755
rect 12190 692 12228 721
rect 12156 686 12262 692
rect 12156 652 12158 686
rect 12192 652 12226 686
rect 12260 652 12262 686
rect 12190 618 12228 652
rect 12156 617 12262 618
rect 12156 583 12158 617
rect 12192 583 12226 617
rect 12260 583 12262 617
rect 12156 578 12262 583
rect 12190 548 12228 578
rect 12156 514 12158 544
rect 12192 514 12226 548
rect 12260 514 12262 544
rect 12156 504 12262 514
rect 12190 479 12228 504
rect 12156 445 12158 470
rect 12192 445 12226 479
rect 12260 445 12262 470
rect 12156 430 12262 445
rect 12190 410 12228 430
rect 12156 376 12158 396
rect 12192 376 12226 410
rect 12260 376 12262 396
rect 12156 356 12262 376
rect 12190 341 12228 356
rect 12156 307 12158 322
rect 12192 307 12226 341
rect 12260 307 12262 322
rect 12156 282 12262 307
rect 12190 272 12228 282
rect 12156 238 12158 248
rect 12192 238 12226 272
rect 12260 238 12262 248
rect 12156 208 12262 238
rect 12190 203 12228 208
rect 12156 169 12158 174
rect 12192 169 12226 203
rect 12260 169 12262 174
rect 12156 134 12262 169
rect 12192 100 12226 134
rect 12156 0 12262 100
rect 12568 3000 12674 3100
rect 12568 2927 12570 2966
rect 12672 2927 12674 2966
rect 12568 2854 12570 2893
rect 12672 2854 12674 2893
rect 12568 2781 12570 2820
rect 12672 2781 12674 2820
rect 12568 2708 12570 2747
rect 12672 2708 12674 2747
rect 12568 2635 12570 2674
rect 12672 2635 12674 2674
rect 12568 2562 12570 2601
rect 12672 2562 12674 2601
rect 12568 2489 12570 2528
rect 12672 2489 12674 2528
rect 12568 2416 12570 2455
rect 12672 2416 12674 2455
rect 12568 2343 12570 2382
rect 12672 2343 12674 2382
rect 12568 2270 12570 2309
rect 12672 2270 12674 2309
rect 12568 2197 12570 2236
rect 12672 2197 12674 2236
rect 12568 2124 12570 2163
rect 12672 2124 12674 2163
rect 12568 2051 12570 2090
rect 12672 2051 12674 2090
rect 12568 1978 12570 2017
rect 12672 1978 12674 2017
rect 12568 1905 12570 1944
rect 12672 1905 12674 1944
rect 12568 1832 12570 1871
rect 12672 1832 12674 1871
rect 12568 1759 12570 1798
rect 12672 1759 12674 1798
rect 12568 1686 12570 1725
rect 12672 1686 12674 1725
rect 12568 1613 12570 1652
rect 12672 1613 12674 1652
rect 12568 1540 12570 1579
rect 12672 1540 12674 1579
rect 12568 1466 12570 1506
rect 12672 1466 12674 1506
rect 12568 1392 12570 1432
rect 12672 1392 12674 1432
rect 12568 1318 12570 1358
rect 12672 1318 12674 1358
rect 12568 1244 12570 1284
rect 12672 1244 12674 1284
rect 12568 1170 12570 1210
rect 12672 1170 12674 1210
rect 12568 1096 12570 1136
rect 12672 1096 12674 1136
rect 12568 1022 12570 1062
rect 12672 1022 12674 1062
rect 12568 948 12570 988
rect 12672 948 12674 988
rect 12568 874 12570 914
rect 12672 874 12674 914
rect 12568 800 12570 840
rect 12672 800 12674 840
rect 12602 766 12640 790
rect 12568 755 12674 766
rect 12568 726 12570 755
rect 12604 721 12638 755
rect 12672 726 12674 755
rect 12602 692 12640 721
rect 12568 686 12674 692
rect 12568 652 12570 686
rect 12604 652 12638 686
rect 12672 652 12674 686
rect 12602 618 12640 652
rect 12568 617 12674 618
rect 12568 583 12570 617
rect 12604 583 12638 617
rect 12672 583 12674 617
rect 12568 578 12674 583
rect 12602 548 12640 578
rect 12568 514 12570 544
rect 12604 514 12638 548
rect 12672 514 12674 544
rect 12568 504 12674 514
rect 12602 479 12640 504
rect 12568 445 12570 470
rect 12604 445 12638 479
rect 12672 445 12674 470
rect 12568 430 12674 445
rect 12602 410 12640 430
rect 12568 376 12570 396
rect 12604 376 12638 410
rect 12672 376 12674 396
rect 12568 356 12674 376
rect 12602 341 12640 356
rect 12568 307 12570 322
rect 12604 307 12638 341
rect 12672 307 12674 322
rect 12568 282 12674 307
rect 12602 272 12640 282
rect 12568 238 12570 248
rect 12604 238 12638 272
rect 12672 238 12674 248
rect 12568 208 12674 238
rect 12602 203 12640 208
rect 12568 169 12570 174
rect 12604 169 12638 203
rect 12672 169 12674 174
rect 12568 134 12674 169
rect 12604 100 12638 134
rect 12568 0 12674 100
rect 12980 3000 13086 3100
rect 12980 2927 12982 2966
rect 13084 2927 13086 2966
rect 12980 2854 12982 2893
rect 13084 2854 13086 2893
rect 12980 2781 12982 2820
rect 13084 2781 13086 2820
rect 12980 2708 12982 2747
rect 13084 2708 13086 2747
rect 12980 2635 12982 2674
rect 13084 2635 13086 2674
rect 12980 2562 12982 2601
rect 13084 2562 13086 2601
rect 12980 2489 12982 2528
rect 13084 2489 13086 2528
rect 12980 2416 12982 2455
rect 13084 2416 13086 2455
rect 12980 2343 12982 2382
rect 13084 2343 13086 2382
rect 12980 2270 12982 2309
rect 13084 2270 13086 2309
rect 12980 2197 12982 2236
rect 13084 2197 13086 2236
rect 12980 2124 12982 2163
rect 13084 2124 13086 2163
rect 12980 2051 12982 2090
rect 13084 2051 13086 2090
rect 12980 1978 12982 2017
rect 13084 1978 13086 2017
rect 12980 1905 12982 1944
rect 13084 1905 13086 1944
rect 12980 1832 12982 1871
rect 13084 1832 13086 1871
rect 12980 1759 12982 1798
rect 13084 1759 13086 1798
rect 12980 1686 12982 1725
rect 13084 1686 13086 1725
rect 12980 1613 12982 1652
rect 13084 1613 13086 1652
rect 12980 1540 12982 1579
rect 13084 1540 13086 1579
rect 12980 1466 12982 1506
rect 13084 1466 13086 1506
rect 12980 1392 12982 1432
rect 13084 1392 13086 1432
rect 12980 1318 12982 1358
rect 13084 1318 13086 1358
rect 12980 1244 12982 1284
rect 13084 1244 13086 1284
rect 12980 1170 12982 1210
rect 13084 1170 13086 1210
rect 12980 1096 12982 1136
rect 13084 1096 13086 1136
rect 12980 1022 12982 1062
rect 13084 1022 13086 1062
rect 12980 948 12982 988
rect 13084 948 13086 988
rect 12980 874 12982 914
rect 13084 874 13086 914
rect 12980 800 12982 840
rect 13084 800 13086 840
rect 13014 766 13052 790
rect 12980 755 13086 766
rect 12980 726 12982 755
rect 13016 721 13050 755
rect 13084 726 13086 755
rect 13014 692 13052 721
rect 12980 686 13086 692
rect 12980 652 12982 686
rect 13016 652 13050 686
rect 13084 652 13086 686
rect 13014 618 13052 652
rect 12980 617 13086 618
rect 12980 583 12982 617
rect 13016 583 13050 617
rect 13084 583 13086 617
rect 12980 578 13086 583
rect 13014 548 13052 578
rect 12980 514 12982 544
rect 13016 514 13050 548
rect 13084 514 13086 544
rect 12980 504 13086 514
rect 13014 479 13052 504
rect 12980 445 12982 470
rect 13016 445 13050 479
rect 13084 445 13086 470
rect 12980 430 13086 445
rect 13014 410 13052 430
rect 12980 376 12982 396
rect 13016 376 13050 410
rect 13084 376 13086 396
rect 12980 356 13086 376
rect 13014 341 13052 356
rect 12980 307 12982 322
rect 13016 307 13050 341
rect 13084 307 13086 322
rect 12980 282 13086 307
rect 13014 272 13052 282
rect 12980 238 12982 248
rect 13016 238 13050 272
rect 13084 238 13086 248
rect 12980 208 13086 238
rect 13014 203 13052 208
rect 12980 169 12982 174
rect 13016 169 13050 203
rect 13084 169 13086 174
rect 12980 134 13086 169
rect 13016 100 13050 134
rect 12980 0 13086 100
rect 13188 480 13202 484
rect 13236 480 13274 484
rect 13308 480 13346 484
rect 13380 480 13418 484
rect 13452 480 13490 484
rect 13524 480 13562 484
rect 13596 480 13634 484
rect 13668 480 13706 484
rect 13740 480 13778 484
rect 13812 480 13850 484
rect 13884 480 13922 484
rect 13956 480 13970 484
rect 13188 449 13970 480
rect 13222 441 13256 449
rect 13290 441 13324 449
rect 13358 441 13392 449
rect 13426 441 13460 449
rect 13494 441 13528 449
rect 13236 415 13256 441
rect 13308 415 13324 441
rect 13380 415 13392 441
rect 13452 415 13460 441
rect 13524 415 13528 441
rect 13562 441 13596 449
rect 13188 407 13202 415
rect 13236 407 13274 415
rect 13308 407 13346 415
rect 13380 407 13418 415
rect 13452 407 13490 415
rect 13524 407 13562 415
rect 13630 441 13664 449
rect 13698 441 13732 449
rect 13766 441 13800 449
rect 13834 441 13868 449
rect 13902 441 13936 449
rect 13630 415 13634 441
rect 13698 415 13706 441
rect 13766 415 13778 441
rect 13834 415 13850 441
rect 13902 415 13922 441
rect 13596 407 13634 415
rect 13668 407 13706 415
rect 13740 407 13778 415
rect 13812 407 13850 415
rect 13884 407 13922 415
rect 13956 407 13970 415
rect 13188 380 13970 407
rect 13222 368 13256 380
rect 13290 368 13324 380
rect 13358 368 13392 380
rect 13426 368 13460 380
rect 13494 368 13528 380
rect 13236 346 13256 368
rect 13308 346 13324 368
rect 13380 346 13392 368
rect 13452 346 13460 368
rect 13524 346 13528 368
rect 13562 368 13596 380
rect 13188 334 13202 346
rect 13236 334 13274 346
rect 13308 334 13346 346
rect 13380 334 13418 346
rect 13452 334 13490 346
rect 13524 334 13562 346
rect 13630 368 13664 380
rect 13698 368 13732 380
rect 13766 368 13800 380
rect 13834 368 13868 380
rect 13902 368 13936 380
rect 13630 346 13634 368
rect 13698 346 13706 368
rect 13766 346 13778 368
rect 13834 346 13850 368
rect 13902 346 13922 368
rect 13596 334 13634 346
rect 13668 334 13706 346
rect 13740 334 13778 346
rect 13812 334 13850 346
rect 13884 334 13922 346
rect 13956 334 13970 346
rect 13188 311 13970 334
rect 13222 295 13256 311
rect 13290 295 13324 311
rect 13358 295 13392 311
rect 13426 295 13460 311
rect 13494 295 13528 311
rect 13236 277 13256 295
rect 13308 277 13324 295
rect 13380 277 13392 295
rect 13452 277 13460 295
rect 13524 277 13528 295
rect 13562 295 13596 311
rect 13188 261 13202 277
rect 13236 261 13274 277
rect 13308 261 13346 277
rect 13380 261 13418 277
rect 13452 261 13490 277
rect 13524 261 13562 277
rect 13630 295 13664 311
rect 13698 295 13732 311
rect 13766 295 13800 311
rect 13834 295 13868 311
rect 13902 295 13936 311
rect 13630 277 13634 295
rect 13698 277 13706 295
rect 13766 277 13778 295
rect 13834 277 13850 295
rect 13902 277 13922 295
rect 13596 261 13634 277
rect 13668 261 13706 277
rect 13740 261 13778 277
rect 13812 261 13850 277
rect 13884 261 13922 277
rect 13956 261 13970 277
rect 13188 242 13970 261
rect 13222 222 13256 242
rect 13290 222 13324 242
rect 13358 222 13392 242
rect 13426 222 13460 242
rect 13494 222 13528 242
rect 13236 208 13256 222
rect 13308 208 13324 222
rect 13380 208 13392 222
rect 13452 208 13460 222
rect 13524 208 13528 222
rect 13562 222 13596 242
rect 13188 188 13202 208
rect 13236 188 13274 208
rect 13308 188 13346 208
rect 13380 188 13418 208
rect 13452 188 13490 208
rect 13524 188 13562 208
rect 13630 222 13664 242
rect 13698 222 13732 242
rect 13766 222 13800 242
rect 13834 222 13868 242
rect 13902 222 13936 242
rect 13630 208 13634 222
rect 13698 208 13706 222
rect 13766 208 13778 222
rect 13834 208 13850 222
rect 13902 208 13922 222
rect 13596 188 13634 208
rect 13668 188 13706 208
rect 13740 188 13778 208
rect 13812 188 13850 208
rect 13884 188 13922 208
rect 13956 188 13970 208
rect 13188 173 13970 188
rect 13222 149 13256 173
rect 13290 149 13324 173
rect 13358 149 13392 173
rect 13426 149 13460 173
rect 13494 149 13528 173
rect 13236 139 13256 149
rect 13308 139 13324 149
rect 13380 139 13392 149
rect 13452 139 13460 149
rect 13524 139 13528 149
rect 13562 149 13596 173
rect 13188 115 13202 139
rect 13236 115 13274 139
rect 13308 115 13346 139
rect 13380 115 13418 139
rect 13452 115 13490 139
rect 13524 115 13562 139
rect 13630 149 13664 173
rect 13698 149 13732 173
rect 13766 149 13800 173
rect 13834 149 13868 173
rect 13902 149 13936 173
rect 13630 139 13634 149
rect 13698 139 13706 149
rect 13766 139 13778 149
rect 13834 139 13850 149
rect 13902 139 13922 149
rect 13596 115 13634 139
rect 13668 115 13706 139
rect 13740 115 13778 139
rect 13812 115 13850 139
rect 13884 115 13922 139
rect 13956 115 13970 139
rect 13188 104 13970 115
rect 13222 76 13256 104
rect 13290 76 13324 104
rect 13358 76 13392 104
rect 13426 76 13460 104
rect 13494 76 13528 104
rect 13236 70 13256 76
rect 13308 70 13324 76
rect 13380 70 13392 76
rect 13452 70 13460 76
rect 13524 70 13528 76
rect 13562 76 13596 104
rect 13188 42 13202 70
rect 13236 42 13274 70
rect 13308 42 13346 70
rect 13380 42 13418 70
rect 13452 42 13490 70
rect 13524 42 13562 70
rect 13630 76 13664 104
rect 13698 76 13732 104
rect 13766 76 13800 104
rect 13834 76 13868 104
rect 13902 76 13936 104
rect 13630 70 13634 76
rect 13698 70 13706 76
rect 13766 70 13778 76
rect 13834 70 13850 76
rect 13902 70 13922 76
rect 13596 42 13634 70
rect 13668 42 13706 70
rect 13740 42 13778 70
rect 13812 42 13850 70
rect 13884 42 13922 70
rect 13956 42 13970 70
rect 13188 35 13970 42
rect 13222 3 13256 35
rect 13290 3 13324 35
rect 13358 3 13392 35
rect 13426 3 13460 35
rect 13494 3 13528 35
rect 13236 1 13256 3
rect 13308 1 13324 3
rect 13380 1 13392 3
rect 13452 1 13460 3
rect 13524 1 13528 3
rect 13562 3 13596 35
rect -1088 -34 -306 -31
rect -1054 -68 -1020 -34
rect -986 -68 -952 -34
rect -918 -68 -884 -34
rect -850 -68 -816 -34
rect -782 -68 -748 -34
rect -714 -68 -680 -34
rect -646 -68 -612 -34
rect -578 -68 -544 -34
rect -510 -68 -476 -34
rect -442 -68 -408 -34
rect -374 -68 -340 -34
rect -1088 -70 -306 -68
rect -1088 -103 -1074 -70
rect -1040 -103 -1002 -70
rect -968 -103 -930 -70
rect -896 -103 -858 -70
rect -824 -103 -786 -70
rect -752 -103 -714 -70
rect -1040 -104 -1020 -103
rect -968 -104 -952 -103
rect -896 -104 -884 -103
rect -824 -104 -816 -103
rect -752 -104 -748 -103
rect -1054 -137 -1020 -104
rect -986 -137 -952 -104
rect -918 -137 -884 -104
rect -850 -137 -816 -104
rect -782 -137 -748 -104
rect -680 -103 -642 -70
rect -608 -103 -570 -70
rect -536 -103 -498 -70
rect -464 -103 -426 -70
rect -392 -103 -354 -70
rect -320 -103 -306 -70
rect -714 -137 -680 -104
rect -646 -104 -642 -103
rect -578 -104 -570 -103
rect -510 -104 -498 -103
rect -442 -104 -426 -103
rect -374 -104 -354 -103
rect -646 -137 -612 -104
rect -578 -137 -544 -104
rect -510 -137 -476 -104
rect -442 -137 -408 -104
rect -374 -137 -340 -104
rect -1088 -143 -306 -137
rect -1088 -172 -1074 -143
rect -1040 -172 -1002 -143
rect -968 -172 -930 -143
rect -896 -172 -858 -143
rect -824 -172 -786 -143
rect -752 -172 -714 -143
rect -1040 -177 -1020 -172
rect -968 -177 -952 -172
rect -896 -177 -884 -172
rect -824 -177 -816 -172
rect -752 -177 -748 -172
rect -1054 -206 -1020 -177
rect -986 -206 -952 -177
rect -918 -206 -884 -177
rect -850 -206 -816 -177
rect -782 -206 -748 -177
rect -680 -172 -642 -143
rect -608 -172 -570 -143
rect -536 -172 -498 -143
rect -464 -172 -426 -143
rect -392 -172 -354 -143
rect -320 -172 -306 -143
rect -714 -206 -680 -177
rect -646 -177 -642 -172
rect -578 -177 -570 -172
rect -510 -177 -498 -172
rect -442 -177 -426 -172
rect -374 -177 -354 -172
rect -646 -206 -612 -177
rect -578 -206 -544 -177
rect -510 -206 -476 -177
rect -442 -206 -408 -177
rect -374 -206 -340 -177
rect -1088 -274 -306 -206
rect 13188 -31 13202 1
rect 13236 -31 13274 1
rect 13308 -31 13346 1
rect 13380 -31 13418 1
rect 13452 -31 13490 1
rect 13524 -31 13562 1
rect 13630 3 13664 35
rect 13698 3 13732 35
rect 13766 3 13800 35
rect 13834 3 13868 35
rect 13902 3 13936 35
rect 13630 1 13634 3
rect 13698 1 13706 3
rect 13766 1 13778 3
rect 13834 1 13850 3
rect 13902 1 13922 3
rect 13596 -31 13634 1
rect 13668 -31 13706 1
rect 13740 -31 13778 1
rect 13812 -31 13850 1
rect 13884 -31 13922 1
rect 13956 -31 13970 1
rect 13188 -34 13970 -31
rect 13222 -68 13256 -34
rect 13290 -68 13324 -34
rect 13358 -68 13392 -34
rect 13426 -68 13460 -34
rect 13494 -68 13528 -34
rect 13562 -68 13596 -34
rect 13630 -68 13664 -34
rect 13698 -68 13732 -34
rect 13766 -68 13800 -34
rect 13834 -68 13868 -34
rect 13902 -68 13936 -34
rect 13188 -70 13970 -68
rect 13188 -103 13202 -70
rect 13236 -103 13274 -70
rect 13308 -103 13346 -70
rect 13380 -103 13418 -70
rect 13452 -103 13490 -70
rect 13524 -103 13562 -70
rect 13236 -104 13256 -103
rect 13308 -104 13324 -103
rect 13380 -104 13392 -103
rect 13452 -104 13460 -103
rect 13524 -104 13528 -103
rect 13222 -137 13256 -104
rect 13290 -137 13324 -104
rect 13358 -137 13392 -104
rect 13426 -137 13460 -104
rect 13494 -137 13528 -104
rect 13596 -103 13634 -70
rect 13668 -103 13706 -70
rect 13740 -103 13778 -70
rect 13812 -103 13850 -70
rect 13884 -103 13922 -70
rect 13956 -103 13970 -70
rect 13562 -137 13596 -104
rect 13630 -104 13634 -103
rect 13698 -104 13706 -103
rect 13766 -104 13778 -103
rect 13834 -104 13850 -103
rect 13902 -104 13922 -103
rect 13630 -137 13664 -104
rect 13698 -137 13732 -104
rect 13766 -137 13800 -104
rect 13834 -137 13868 -104
rect 13902 -137 13936 -104
rect 13188 -143 13970 -137
rect 13188 -172 13202 -143
rect 13236 -172 13274 -143
rect 13308 -172 13346 -143
rect 13380 -172 13418 -143
rect 13452 -172 13490 -143
rect 13524 -172 13562 -143
rect 13236 -177 13256 -172
rect 13308 -177 13324 -172
rect 13380 -177 13392 -172
rect 13452 -177 13460 -172
rect 13524 -177 13528 -172
rect 13222 -206 13256 -177
rect 13290 -206 13324 -177
rect 13358 -206 13392 -177
rect 13426 -206 13460 -177
rect 13494 -206 13528 -177
rect 13596 -172 13634 -143
rect 13668 -172 13706 -143
rect 13740 -172 13778 -143
rect 13812 -172 13850 -143
rect 13884 -172 13922 -143
rect 13956 -172 13970 -143
rect 13562 -206 13596 -177
rect 13630 -177 13634 -172
rect 13698 -177 13706 -172
rect 13766 -177 13778 -172
rect 13834 -177 13850 -172
rect 13902 -177 13922 -172
rect 13630 -206 13664 -177
rect 13698 -206 13732 -177
rect 13766 -206 13800 -177
rect 13834 -206 13868 -177
rect 13902 -206 13936 -177
rect 13188 -274 13970 -206
rect -1088 -308 -1020 -274
rect -986 -308 -951 -274
rect -917 -306 -882 -274
rect -917 -308 -886 -306
rect -848 -308 -813 -274
rect -779 -308 -744 -274
rect -710 -306 -675 -274
rect -641 -306 -606 -274
rect -572 -306 -537 -274
rect -503 -306 -468 -274
rect -434 -306 -399 -274
rect -365 -306 -330 -274
rect -296 -306 -261 -274
rect -227 -306 -192 -274
rect -158 -306 -123 -274
rect -89 -306 -54 -274
rect -20 -306 15 -274
rect 49 -306 84 -274
rect 118 -306 153 -274
rect 187 -306 222 -274
rect 256 -306 291 -274
rect 325 -306 360 -274
rect 394 -306 429 -274
rect 463 -306 498 -274
rect 532 -306 567 -274
rect 601 -306 636 -274
rect 670 -306 705 -274
rect 739 -306 774 -274
rect 808 -306 843 -274
rect 877 -306 912 -274
rect 946 -306 981 -274
rect 1015 -306 1050 -274
rect 1084 -306 1119 -274
rect 1153 -306 1188 -274
rect 1222 -306 1257 -274
rect 1291 -306 1326 -274
rect 1360 -306 1395 -274
rect 1429 -306 1464 -274
rect 1498 -306 1533 -274
rect 1567 -306 1602 -274
rect 1636 -306 1671 -274
rect 1705 -306 1740 -274
rect 1774 -306 1809 -274
rect 1843 -306 1878 -274
rect 1912 -306 1947 -274
rect 1981 -306 2016 -274
rect 2050 -306 2085 -274
rect 2119 -306 2154 -274
rect 2188 -306 2223 -274
rect 2257 -306 2292 -274
rect 2326 -306 2361 -274
rect 2395 -306 2430 -274
rect 2464 -306 2499 -274
rect 2533 -306 2568 -274
rect 2602 -306 2637 -274
rect 2671 -306 2706 -274
rect 2740 -306 2775 -274
rect 2809 -306 2844 -274
rect 2878 -306 2913 -274
rect 2947 -306 2982 -274
rect 3016 -306 3051 -274
rect 3085 -306 3120 -274
rect 3154 -306 3189 -274
rect 3223 -306 3258 -274
rect 3292 -306 3327 -274
rect 3361 -306 3396 -274
rect -706 -308 -675 -306
rect -633 -308 -606 -306
rect -1088 -340 -886 -308
rect -852 -340 -813 -308
rect -779 -340 -740 -308
rect -706 -340 -667 -308
rect -633 -340 -594 -308
rect -1088 -342 -594 -340
rect -1088 -376 -1020 -342
rect -986 -376 -951 -342
rect -917 -376 -882 -342
rect -848 -376 -813 -342
rect -779 -376 -744 -342
rect -710 -376 -675 -342
rect -641 -376 -606 -342
rect -1088 -378 -594 -376
rect -1088 -410 -886 -378
rect -852 -410 -813 -378
rect -779 -410 -740 -378
rect -706 -410 -667 -378
rect -633 -410 -594 -378
rect -1088 -444 -1020 -410
rect -986 -444 -951 -410
rect -917 -412 -886 -410
rect -917 -444 -882 -412
rect -848 -444 -813 -410
rect -779 -444 -744 -410
rect -706 -412 -675 -410
rect -633 -412 -606 -410
rect -710 -444 -675 -412
rect -641 -444 -606 -412
rect -572 -444 -537 -412
rect -503 -444 -468 -412
rect -434 -444 -399 -412
rect -365 -444 -330 -412
rect -296 -444 -261 -412
rect -227 -444 -192 -412
rect -158 -444 -123 -412
rect -89 -444 -54 -412
rect -20 -444 15 -412
rect 49 -444 84 -412
rect 118 -444 153 -412
rect 187 -444 222 -412
rect 256 -444 291 -412
rect 325 -444 360 -412
rect 394 -444 429 -412
rect 463 -444 498 -412
rect 532 -444 567 -412
rect 601 -444 636 -412
rect 670 -444 705 -412
rect 739 -444 774 -412
rect 808 -444 843 -412
rect 877 -444 912 -412
rect 946 -444 981 -412
rect 1015 -444 1050 -412
rect 1084 -444 1119 -412
rect 1153 -444 1188 -412
rect 1222 -444 1257 -412
rect 1291 -444 1326 -412
rect 1360 -444 1395 -412
rect 1429 -444 1464 -412
rect 1498 -444 1533 -412
rect 1567 -444 1602 -412
rect 1636 -444 1671 -412
rect 1705 -444 1740 -412
rect 1774 -444 1809 -412
rect 1843 -444 1878 -412
rect 1912 -444 1947 -412
rect 1981 -444 2016 -412
rect 2050 -444 2085 -412
rect 2119 -444 2154 -412
rect 2188 -444 2223 -412
rect 2257 -444 2292 -412
rect 2326 -444 2361 -412
rect 2395 -444 2430 -412
rect 2464 -444 2499 -412
rect 2533 -444 2568 -412
rect 2602 -444 2637 -412
rect 2671 -444 2706 -412
rect 2740 -444 2775 -412
rect 2809 -444 2844 -412
rect 2878 -444 2913 -412
rect 2947 -444 2982 -412
rect 3016 -444 3051 -412
rect 3085 -444 3120 -412
rect 3154 -444 3189 -412
rect 3223 -444 3258 -412
rect 3292 -444 3327 -412
rect 3361 -444 3396 -412
rect 13902 -444 13970 -274
rect 14170 -440 14340 -438
rect -1392 -474 -1390 -473
rect -1424 -507 -1390 -474
rect -1356 -474 -1354 -473
rect -1356 -507 -1322 -474
rect -1458 -513 -1288 -507
rect -1458 -542 -1426 -513
rect -1392 -542 -1354 -513
rect -1320 -542 -1288 -513
rect -1392 -547 -1390 -542
rect -1424 -576 -1390 -547
rect -1356 -547 -1354 -542
rect -1356 -576 -1322 -547
rect -1458 -644 -1288 -576
rect 14170 -473 14202 -440
rect 14236 -473 14274 -440
rect 14308 -473 14340 -440
rect 14236 -474 14238 -473
rect 14204 -507 14238 -474
rect 14272 -474 14274 -473
rect 14272 -507 14306 -474
rect 14170 -513 14340 -507
rect 14170 -542 14202 -513
rect 14236 -542 14274 -513
rect 14308 -542 14340 -513
rect 14236 -547 14238 -542
rect 14204 -576 14238 -547
rect 14272 -547 14274 -542
rect 14272 -576 14306 -547
rect 14170 -644 14340 -576
rect -1458 -678 -1390 -644
rect -1356 -678 -1321 -644
rect -1287 -678 -1252 -644
rect -1218 -676 -1183 -644
rect -1149 -676 -1114 -644
rect -1218 -678 -1191 -676
rect -1149 -678 -1118 -676
rect -1080 -678 -1045 -644
rect -1011 -678 -976 -644
rect -942 -676 -907 -644
rect -873 -676 -838 -644
rect -804 -676 -769 -644
rect -735 -676 -700 -644
rect -666 -676 -631 -644
rect -597 -676 -562 -644
rect -528 -676 -493 -644
rect -459 -676 -424 -644
rect -938 -678 -907 -676
rect -865 -678 -838 -676
rect -792 -678 -769 -676
rect -719 -678 -700 -676
rect -646 -678 -631 -676
rect -573 -678 -562 -676
rect -500 -678 -493 -676
rect -427 -678 -424 -676
rect -390 -676 -355 -644
rect -321 -676 -286 -644
rect -252 -676 -217 -644
rect -183 -676 -148 -644
rect -114 -676 -79 -644
rect -45 -676 -10 -644
rect 24 -676 59 -644
rect 93 -676 128 -644
rect 162 -676 197 -644
rect -390 -678 -388 -676
rect -321 -678 -315 -676
rect -252 -678 -242 -676
rect -183 -678 -169 -676
rect -114 -678 -96 -676
rect -45 -678 -23 -676
rect 24 -678 50 -676
rect 93 -678 123 -676
rect 162 -678 196 -676
rect 231 -678 266 -644
rect 300 -676 335 -644
rect 369 -676 404 -644
rect 438 -676 473 -644
rect 507 -676 542 -644
rect 576 -676 611 -644
rect 645 -676 680 -644
rect 714 -676 749 -644
rect 783 -676 818 -644
rect 303 -678 335 -676
rect 376 -678 404 -676
rect 449 -678 473 -676
rect 522 -678 542 -676
rect 595 -678 611 -676
rect 668 -678 680 -676
rect 741 -678 749 -676
rect 814 -678 818 -676
rect 852 -676 887 -644
rect 852 -678 853 -676
rect -1458 -710 -1191 -678
rect -1157 -710 -1118 -678
rect -1084 -710 -1045 -678
rect -1011 -710 -972 -678
rect -938 -710 -899 -678
rect -865 -710 -826 -678
rect -792 -710 -753 -678
rect -719 -710 -680 -678
rect -646 -710 -607 -678
rect -573 -710 -534 -678
rect -500 -710 -461 -678
rect -427 -710 -388 -678
rect -354 -710 -315 -678
rect -281 -710 -242 -678
rect -208 -710 -169 -678
rect -135 -710 -96 -678
rect -62 -710 -23 -678
rect 11 -710 50 -678
rect 84 -710 123 -678
rect 157 -710 196 -678
rect 230 -710 269 -678
rect 303 -710 342 -678
rect 376 -710 415 -678
rect 449 -710 488 -678
rect 522 -710 561 -678
rect 595 -710 634 -678
rect 668 -710 707 -678
rect 741 -710 780 -678
rect 814 -710 853 -678
rect 921 -676 956 -644
rect 990 -676 1025 -644
rect 1059 -676 1094 -644
rect 1128 -676 1163 -644
rect 1197 -676 1232 -644
rect 1266 -676 1301 -644
rect 1335 -676 1370 -644
rect 1404 -676 1439 -644
rect 921 -678 926 -676
rect 990 -678 999 -676
rect 1059 -678 1072 -676
rect 1128 -678 1145 -676
rect 1197 -678 1218 -676
rect 1266 -678 1291 -676
rect 1335 -678 1364 -676
rect 1404 -678 1437 -676
rect 1473 -678 1508 -644
rect 1542 -676 1577 -644
rect 1611 -676 1646 -644
rect 1680 -676 1715 -644
rect 1749 -676 1784 -644
rect 1818 -676 1853 -644
rect 1887 -676 1922 -644
rect 1956 -676 1991 -644
rect 2025 -676 2060 -644
rect 2094 -676 2129 -644
rect 2163 -676 2198 -644
rect 2232 -676 2267 -644
rect 2301 -676 2336 -644
rect 2370 -676 2405 -644
rect 2439 -676 2474 -644
rect 1544 -678 1577 -676
rect 887 -710 926 -678
rect 960 -710 999 -678
rect 1033 -710 1072 -678
rect 1106 -710 1145 -678
rect 1179 -710 1218 -678
rect 1252 -710 1291 -678
rect 1325 -710 1364 -678
rect 1398 -710 1437 -678
rect 1471 -710 1510 -678
rect 1544 -710 1583 -678
rect -1458 -712 1583 -710
rect -1458 -746 -1390 -712
rect -1356 -746 -1321 -712
rect -1287 -746 -1252 -712
rect -1218 -746 -1183 -712
rect -1149 -746 -1114 -712
rect -1080 -746 -1045 -712
rect -1011 -746 -976 -712
rect -942 -746 -907 -712
rect -873 -746 -838 -712
rect -804 -746 -769 -712
rect -735 -746 -700 -712
rect -666 -746 -631 -712
rect -597 -746 -562 -712
rect -528 -746 -493 -712
rect -459 -746 -424 -712
rect -390 -746 -355 -712
rect -321 -746 -286 -712
rect -252 -746 -217 -712
rect -183 -746 -148 -712
rect -114 -746 -79 -712
rect -45 -746 -10 -712
rect 24 -746 59 -712
rect 93 -746 128 -712
rect 162 -746 197 -712
rect 231 -746 266 -712
rect 300 -746 335 -712
rect 369 -746 404 -712
rect 438 -746 473 -712
rect 507 -746 542 -712
rect 576 -746 611 -712
rect 645 -746 680 -712
rect 714 -746 749 -712
rect 783 -746 818 -712
rect 852 -746 887 -712
rect 921 -746 956 -712
rect 990 -746 1025 -712
rect 1059 -746 1094 -712
rect 1128 -746 1163 -712
rect 1197 -746 1232 -712
rect 1266 -746 1301 -712
rect 1335 -746 1370 -712
rect 1404 -746 1439 -712
rect 1473 -746 1508 -712
rect 1542 -746 1577 -712
rect -1458 -748 1583 -746
rect -1458 -780 -1191 -748
rect -1157 -780 -1118 -748
rect -1084 -780 -1045 -748
rect -1011 -780 -972 -748
rect -938 -780 -899 -748
rect -865 -780 -826 -748
rect -792 -780 -753 -748
rect -719 -780 -680 -748
rect -646 -780 -607 -748
rect -573 -780 -534 -748
rect -500 -780 -461 -748
rect -427 -780 -388 -748
rect -354 -780 -315 -748
rect -281 -780 -242 -748
rect -208 -780 -169 -748
rect -135 -780 -96 -748
rect -62 -780 -23 -748
rect 11 -780 50 -748
rect 84 -780 123 -748
rect 157 -780 196 -748
rect 230 -780 269 -748
rect 303 -780 342 -748
rect 376 -780 415 -748
rect 449 -780 488 -748
rect 522 -780 561 -748
rect 595 -780 634 -748
rect 668 -780 707 -748
rect 741 -780 780 -748
rect 814 -780 853 -748
rect -1458 -814 -1390 -780
rect -1356 -814 -1321 -780
rect -1287 -814 -1252 -780
rect -1218 -782 -1191 -780
rect -1149 -782 -1118 -780
rect -1218 -814 -1183 -782
rect -1149 -814 -1114 -782
rect -1080 -814 -1045 -780
rect -1011 -814 -976 -780
rect -938 -782 -907 -780
rect -865 -782 -838 -780
rect -792 -782 -769 -780
rect -719 -782 -700 -780
rect -646 -782 -631 -780
rect -573 -782 -562 -780
rect -500 -782 -493 -780
rect -427 -782 -424 -780
rect -942 -814 -907 -782
rect -873 -814 -838 -782
rect -804 -814 -769 -782
rect -735 -814 -700 -782
rect -666 -814 -631 -782
rect -597 -814 -562 -782
rect -528 -814 -493 -782
rect -459 -814 -424 -782
rect -390 -782 -388 -780
rect -321 -782 -315 -780
rect -252 -782 -242 -780
rect -183 -782 -169 -780
rect -114 -782 -96 -780
rect -45 -782 -23 -780
rect 24 -782 50 -780
rect 93 -782 123 -780
rect 162 -782 196 -780
rect -390 -814 -355 -782
rect -321 -814 -286 -782
rect -252 -814 -217 -782
rect -183 -814 -148 -782
rect -114 -814 -79 -782
rect -45 -814 -10 -782
rect 24 -814 59 -782
rect 93 -814 128 -782
rect 162 -814 197 -782
rect 231 -814 266 -780
rect 303 -782 335 -780
rect 376 -782 404 -780
rect 449 -782 473 -780
rect 522 -782 542 -780
rect 595 -782 611 -780
rect 668 -782 680 -780
rect 741 -782 749 -780
rect 814 -782 818 -780
rect 300 -814 335 -782
rect 369 -814 404 -782
rect 438 -814 473 -782
rect 507 -814 542 -782
rect 576 -814 611 -782
rect 645 -814 680 -782
rect 714 -814 749 -782
rect 783 -814 818 -782
rect 852 -782 853 -780
rect 887 -780 926 -748
rect 960 -780 999 -748
rect 1033 -780 1072 -748
rect 1106 -780 1145 -748
rect 1179 -780 1218 -748
rect 1252 -780 1291 -748
rect 1325 -780 1364 -748
rect 1398 -780 1437 -748
rect 1471 -780 1510 -748
rect 1544 -780 1583 -748
rect 852 -814 887 -782
rect 921 -782 926 -780
rect 990 -782 999 -780
rect 1059 -782 1072 -780
rect 1128 -782 1145 -780
rect 1197 -782 1218 -780
rect 1266 -782 1291 -780
rect 1335 -782 1364 -780
rect 1404 -782 1437 -780
rect 921 -814 956 -782
rect 990 -814 1025 -782
rect 1059 -814 1094 -782
rect 1128 -814 1163 -782
rect 1197 -814 1232 -782
rect 1266 -814 1301 -782
rect 1335 -814 1370 -782
rect 1404 -814 1439 -782
rect 1473 -814 1508 -780
rect 1544 -782 1577 -780
rect 1542 -814 1577 -782
rect 1611 -814 1646 -782
rect 1680 -814 1715 -782
rect 1749 -814 1784 -782
rect 1818 -814 1853 -782
rect 1887 -814 1922 -782
rect 1956 -814 1991 -782
rect 2025 -814 2060 -782
rect 2094 -814 2129 -782
rect 2163 -814 2198 -782
rect 2232 -814 2267 -782
rect 2301 -814 2336 -782
rect 2370 -814 2405 -782
rect 2439 -814 2474 -782
rect 14272 -814 14340 -644
<< viali >>
rect -1191 3880 -1183 3882
rect -1183 3880 -1157 3882
rect -1118 3880 -1114 3882
rect -1114 3880 -1084 3882
rect -1045 3880 -1011 3882
rect -972 3880 -942 3882
rect -942 3880 -938 3882
rect -899 3880 -873 3882
rect -873 3880 -865 3882
rect -826 3880 -804 3882
rect -804 3880 -792 3882
rect -753 3880 -735 3882
rect -735 3880 -719 3882
rect -680 3880 -666 3882
rect -666 3880 -646 3882
rect -607 3880 -597 3882
rect -597 3880 -573 3882
rect -534 3880 -528 3882
rect -528 3880 -500 3882
rect -461 3880 -459 3882
rect -459 3880 -427 3882
rect -388 3880 -355 3882
rect -355 3880 -354 3882
rect -315 3880 -286 3882
rect -286 3880 -281 3882
rect -242 3880 -217 3882
rect -217 3880 -208 3882
rect -169 3880 -148 3882
rect -148 3880 -135 3882
rect -96 3880 -79 3882
rect -79 3880 -62 3882
rect -23 3880 -10 3882
rect -10 3880 11 3882
rect 50 3880 59 3882
rect 59 3880 84 3882
rect 123 3880 128 3882
rect 128 3880 157 3882
rect 196 3880 197 3882
rect 197 3880 230 3882
rect 269 3880 300 3882
rect 300 3880 303 3882
rect 342 3880 369 3882
rect 369 3880 376 3882
rect 415 3880 438 3882
rect 438 3880 449 3882
rect 488 3880 507 3882
rect 507 3880 522 3882
rect 561 3880 576 3882
rect 576 3880 595 3882
rect 634 3880 645 3882
rect 645 3880 668 3882
rect 707 3880 714 3882
rect 714 3880 741 3882
rect 780 3880 783 3882
rect 783 3880 814 3882
rect -1191 3848 -1157 3880
rect -1118 3848 -1084 3880
rect -1045 3848 -1011 3880
rect -972 3848 -938 3880
rect -899 3848 -865 3880
rect -826 3848 -792 3880
rect -753 3848 -719 3880
rect -680 3848 -646 3880
rect -607 3848 -573 3880
rect -534 3848 -500 3880
rect -461 3848 -427 3880
rect -388 3848 -354 3880
rect -315 3848 -281 3880
rect -242 3848 -208 3880
rect -169 3848 -135 3880
rect -96 3848 -62 3880
rect -23 3848 11 3880
rect 50 3848 84 3880
rect 123 3848 157 3880
rect 196 3848 230 3880
rect 269 3848 303 3880
rect 342 3848 376 3880
rect 415 3848 449 3880
rect 488 3848 522 3880
rect 561 3848 595 3880
rect 634 3848 668 3880
rect 707 3848 741 3880
rect 780 3848 814 3880
rect 853 3848 887 3882
rect 926 3880 956 3882
rect 956 3880 960 3882
rect 999 3880 1025 3882
rect 1025 3880 1033 3882
rect 1072 3880 1094 3882
rect 1094 3880 1106 3882
rect 1145 3880 1163 3882
rect 1163 3880 1179 3882
rect 1218 3880 1232 3882
rect 1232 3880 1252 3882
rect 1291 3880 1301 3882
rect 1301 3880 1325 3882
rect 1364 3880 1370 3882
rect 1370 3880 1398 3882
rect 1437 3880 1439 3882
rect 1439 3880 1471 3882
rect 1510 3880 1542 3882
rect 1542 3880 1544 3882
rect 1583 3880 1611 3882
rect 1611 3880 1646 3882
rect 1646 3880 1680 3882
rect 1680 3880 1715 3882
rect 1715 3880 1749 3882
rect 1749 3880 1784 3882
rect 1784 3880 1818 3882
rect 1818 3880 1853 3882
rect 1853 3880 1887 3882
rect 1887 3880 1922 3882
rect 1922 3880 1956 3882
rect 1956 3880 1991 3882
rect 1991 3880 2025 3882
rect 2025 3880 2060 3882
rect 2060 3880 2094 3882
rect 2094 3880 2129 3882
rect 2129 3880 2163 3882
rect 2163 3880 2198 3882
rect 2198 3880 2232 3882
rect 2232 3880 2267 3882
rect 2267 3880 2301 3882
rect 2301 3880 2336 3882
rect 2336 3880 2370 3882
rect 2370 3880 2405 3882
rect 2405 3880 2439 3882
rect 2439 3880 2474 3882
rect 926 3848 960 3880
rect 999 3848 1033 3880
rect 1072 3848 1106 3880
rect 1145 3848 1179 3880
rect 1218 3848 1252 3880
rect 1291 3848 1325 3880
rect 1364 3848 1398 3880
rect 1437 3848 1471 3880
rect 1510 3848 1544 3880
rect 1583 3846 2474 3880
rect 1583 3812 1611 3846
rect 1611 3812 1646 3846
rect 1646 3812 1680 3846
rect 1680 3812 1715 3846
rect 1715 3812 1749 3846
rect 1749 3812 1784 3846
rect 1784 3812 1818 3846
rect 1818 3812 1853 3846
rect 1853 3812 1887 3846
rect 1887 3812 1922 3846
rect 1922 3812 1956 3846
rect 1956 3812 1991 3846
rect 1991 3812 2025 3846
rect 2025 3812 2060 3846
rect 2060 3812 2094 3846
rect 2094 3812 2129 3846
rect 2129 3812 2163 3846
rect 2163 3812 2198 3846
rect 2198 3812 2232 3846
rect 2232 3812 2267 3846
rect 2267 3812 2301 3846
rect 2301 3812 2336 3846
rect 2336 3812 2370 3846
rect 2370 3812 2405 3846
rect 2405 3812 2439 3846
rect 2439 3812 2474 3846
rect -1191 3778 -1157 3810
rect -1118 3778 -1084 3810
rect -1045 3778 -1011 3810
rect -972 3778 -938 3810
rect -899 3778 -865 3810
rect -826 3778 -792 3810
rect -753 3778 -719 3810
rect -680 3778 -646 3810
rect -607 3778 -573 3810
rect -534 3778 -500 3810
rect -461 3778 -427 3810
rect -388 3778 -354 3810
rect -315 3778 -281 3810
rect -242 3778 -208 3810
rect -169 3778 -135 3810
rect -96 3778 -62 3810
rect -23 3778 11 3810
rect 50 3778 84 3810
rect 123 3778 157 3810
rect 196 3778 230 3810
rect 269 3778 303 3810
rect 342 3778 376 3810
rect 415 3778 449 3810
rect 488 3778 522 3810
rect 561 3778 595 3810
rect 634 3778 668 3810
rect 707 3778 741 3810
rect 780 3778 814 3810
rect -1191 3776 -1183 3778
rect -1183 3776 -1157 3778
rect -1118 3776 -1114 3778
rect -1114 3776 -1084 3778
rect -1045 3776 -1011 3778
rect -972 3776 -942 3778
rect -942 3776 -938 3778
rect -899 3776 -873 3778
rect -873 3776 -865 3778
rect -826 3776 -804 3778
rect -804 3776 -792 3778
rect -753 3776 -735 3778
rect -735 3776 -719 3778
rect -680 3776 -666 3778
rect -666 3776 -646 3778
rect -607 3776 -597 3778
rect -597 3776 -573 3778
rect -534 3776 -528 3778
rect -528 3776 -500 3778
rect -461 3776 -459 3778
rect -459 3776 -427 3778
rect -388 3776 -355 3778
rect -355 3776 -354 3778
rect -315 3776 -286 3778
rect -286 3776 -281 3778
rect -242 3776 -217 3778
rect -217 3776 -208 3778
rect -169 3776 -148 3778
rect -148 3776 -135 3778
rect -96 3776 -79 3778
rect -79 3776 -62 3778
rect -23 3776 -10 3778
rect -10 3776 11 3778
rect 50 3776 59 3778
rect 59 3776 84 3778
rect 123 3776 128 3778
rect 128 3776 157 3778
rect 196 3776 197 3778
rect 197 3776 230 3778
rect 269 3776 300 3778
rect 300 3776 303 3778
rect 342 3776 369 3778
rect 369 3776 376 3778
rect 415 3776 438 3778
rect 438 3776 449 3778
rect 488 3776 507 3778
rect 507 3776 522 3778
rect 561 3776 576 3778
rect 576 3776 595 3778
rect 634 3776 645 3778
rect 645 3776 668 3778
rect 707 3776 714 3778
rect 714 3776 741 3778
rect 780 3776 783 3778
rect 783 3776 814 3778
rect 853 3776 887 3810
rect 926 3778 960 3810
rect 999 3778 1033 3810
rect 1072 3778 1106 3810
rect 1145 3778 1179 3810
rect 1218 3778 1252 3810
rect 1291 3778 1325 3810
rect 1364 3778 1398 3810
rect 1437 3778 1471 3810
rect 1510 3778 1544 3810
rect 1583 3778 2474 3812
rect 926 3776 956 3778
rect 956 3776 960 3778
rect 999 3776 1025 3778
rect 1025 3776 1033 3778
rect 1072 3776 1094 3778
rect 1094 3776 1106 3778
rect 1145 3776 1163 3778
rect 1163 3776 1179 3778
rect 1218 3776 1232 3778
rect 1232 3776 1252 3778
rect 1291 3776 1301 3778
rect 1301 3776 1325 3778
rect 1364 3776 1370 3778
rect 1370 3776 1398 3778
rect 1437 3776 1439 3778
rect 1439 3776 1471 3778
rect 1510 3776 1542 3778
rect 1542 3776 1544 3778
rect 1583 3776 1611 3778
rect 1611 3776 1646 3778
rect 1646 3776 1680 3778
rect 1680 3776 1715 3778
rect 1715 3776 1749 3778
rect 1749 3776 1784 3778
rect 1784 3776 1818 3778
rect 1818 3776 1853 3778
rect 1853 3776 1887 3778
rect 1887 3776 1922 3778
rect 1922 3776 1956 3778
rect 1956 3776 1991 3778
rect 1991 3776 2025 3778
rect 2025 3776 2060 3778
rect 2060 3776 2094 3778
rect 2094 3776 2129 3778
rect 2129 3776 2163 3778
rect 2163 3776 2198 3778
rect 2198 3776 2232 3778
rect 2232 3776 2267 3778
rect 2267 3776 2301 3778
rect 2301 3776 2336 3778
rect 2336 3776 2370 3778
rect 2370 3776 2405 3778
rect 2405 3776 2439 3778
rect 2439 3776 2474 3778
rect 2474 3776 14073 3882
rect -1426 3541 -1320 3647
rect -1426 3468 -1392 3502
rect -1354 3468 -1320 3502
rect -1426 3395 -1392 3429
rect -1354 3395 -1320 3429
rect -1426 3322 -1392 3356
rect -1354 3322 -1320 3356
rect -1426 3249 -1392 3283
rect -1354 3249 -1320 3283
rect -1426 3176 -1392 3210
rect -1354 3176 -1320 3210
rect -1426 3103 -1392 3137
rect -1354 3103 -1320 3137
rect -1426 3030 -1392 3064
rect -1354 3030 -1320 3064
rect -1426 2957 -1392 2991
rect -1354 2957 -1320 2991
rect -1426 2884 -1392 2918
rect -1354 2884 -1320 2918
rect -1426 2811 -1392 2845
rect -1354 2811 -1320 2845
rect -1426 2738 -1392 2772
rect -1354 2738 -1320 2772
rect -1426 2665 -1392 2699
rect -1354 2665 -1320 2699
rect -1426 2592 -1392 2626
rect -1354 2592 -1320 2626
rect -1426 2519 -1392 2553
rect -1354 2519 -1320 2553
rect -1426 2446 -1392 2480
rect -1354 2446 -1320 2480
rect -1426 2373 -1392 2407
rect -1354 2373 -1320 2407
rect -1426 2300 -1392 2334
rect -1354 2300 -1320 2334
rect -1426 2227 -1392 2261
rect -1354 2227 -1320 2261
rect -1426 2154 -1392 2188
rect -1354 2154 -1320 2188
rect -1426 2081 -1392 2115
rect -1354 2081 -1320 2115
rect -1426 2008 -1392 2042
rect -1354 2008 -1320 2042
rect -1426 1935 -1392 1969
rect -1354 1935 -1320 1969
rect -1426 1862 -1392 1896
rect -1354 1862 -1320 1896
rect -1426 1789 -1392 1823
rect -1354 1789 -1320 1823
rect -1426 1716 -1392 1750
rect -1354 1716 -1320 1750
rect -1426 1643 -1392 1677
rect -1354 1643 -1320 1677
rect -1426 1570 -1392 1604
rect -1354 1570 -1320 1604
rect -1426 1497 -1392 1531
rect -1354 1497 -1320 1531
rect -1426 1424 -1392 1458
rect -1354 1424 -1320 1458
rect -1426 1351 -1392 1385
rect -1354 1351 -1320 1385
rect -1426 1278 -1392 1312
rect -1354 1278 -1320 1312
rect -1426 1205 -1392 1239
rect -1354 1205 -1320 1239
rect -1426 1132 -1392 1166
rect -1354 1132 -1320 1166
rect -1426 1059 -1392 1093
rect -1354 1059 -1320 1093
rect -1426 986 -1392 1020
rect -1354 986 -1320 1020
rect -1426 913 -1392 947
rect -1354 913 -1320 947
rect -1426 840 -1392 874
rect -1354 840 -1320 874
rect -1426 767 -1392 801
rect -1354 767 -1320 801
rect -1426 694 -1392 728
rect -1354 694 -1320 728
rect -1426 621 -1392 655
rect -1354 621 -1320 655
rect -1426 548 -1392 582
rect -1354 548 -1320 582
rect -1426 475 -1392 509
rect -1354 475 -1320 509
rect -1426 402 -1392 436
rect -1354 402 -1320 436
rect -1426 329 -1392 363
rect -1354 329 -1320 363
rect -1426 256 -1392 290
rect -1354 256 -1320 290
rect -1426 183 -1392 217
rect -1354 183 -1320 217
rect -1426 110 -1392 144
rect -1354 110 -1320 144
rect -1426 37 -1392 71
rect -1354 37 -1320 71
rect -1426 -36 -1392 -2
rect -1354 -36 -1320 -2
rect -1426 -109 -1392 -75
rect -1354 -109 -1320 -75
rect -1426 -182 -1392 -148
rect -1354 -182 -1320 -148
rect -1426 -255 -1392 -221
rect -1354 -255 -1320 -221
rect -1426 -328 -1392 -294
rect -1354 -328 -1320 -294
rect -1426 -401 -1392 -367
rect -1354 -401 -1320 -367
rect -1426 -473 -1392 -440
rect -1354 -473 -1320 -440
rect -886 3510 -882 3512
rect -882 3510 -852 3512
rect -813 3510 -779 3512
rect -740 3510 -710 3512
rect -710 3510 -706 3512
rect -667 3510 -641 3512
rect -641 3510 -633 3512
rect -594 3510 -572 3512
rect -572 3510 -537 3512
rect -537 3510 -503 3512
rect -503 3510 -468 3512
rect -468 3510 -434 3512
rect -434 3510 -399 3512
rect -399 3510 -365 3512
rect -365 3510 -330 3512
rect -330 3510 -296 3512
rect -296 3510 -261 3512
rect -261 3510 -227 3512
rect -227 3510 -192 3512
rect -192 3510 -158 3512
rect -158 3510 -123 3512
rect -123 3510 -89 3512
rect -89 3510 -54 3512
rect -54 3510 -20 3512
rect -20 3510 15 3512
rect 15 3510 49 3512
rect 49 3510 84 3512
rect 84 3510 118 3512
rect 118 3510 153 3512
rect 153 3510 187 3512
rect 187 3510 222 3512
rect 222 3510 256 3512
rect 256 3510 291 3512
rect 291 3510 325 3512
rect 325 3510 360 3512
rect 360 3510 394 3512
rect 394 3510 429 3512
rect 429 3510 463 3512
rect 463 3510 498 3512
rect 498 3510 532 3512
rect 532 3510 567 3512
rect 567 3510 601 3512
rect 601 3510 636 3512
rect 636 3510 670 3512
rect 670 3510 705 3512
rect 705 3510 739 3512
rect 739 3510 774 3512
rect 774 3510 808 3512
rect 808 3510 843 3512
rect 843 3510 877 3512
rect 877 3510 912 3512
rect 912 3510 946 3512
rect 946 3510 981 3512
rect 981 3510 1015 3512
rect 1015 3510 1050 3512
rect 1050 3510 1084 3512
rect 1084 3510 1119 3512
rect 1119 3510 1153 3512
rect 1153 3510 1188 3512
rect 1188 3510 1222 3512
rect 1222 3510 1257 3512
rect 1257 3510 1291 3512
rect 1291 3510 1326 3512
rect 1326 3510 1360 3512
rect 1360 3510 1395 3512
rect 1395 3510 1429 3512
rect 1429 3510 1464 3512
rect 1464 3510 1498 3512
rect 1498 3510 1533 3512
rect 1533 3510 1567 3512
rect 1567 3510 1602 3512
rect 1602 3510 1636 3512
rect 1636 3510 1671 3512
rect 1671 3510 1705 3512
rect 1705 3510 1740 3512
rect 1740 3510 1774 3512
rect 1774 3510 1809 3512
rect 1809 3510 1843 3512
rect 1843 3510 1878 3512
rect 1878 3510 1912 3512
rect 1912 3510 1947 3512
rect 1947 3510 1981 3512
rect 1981 3510 2016 3512
rect 2016 3510 2050 3512
rect 2050 3510 2085 3512
rect 2085 3510 2119 3512
rect 2119 3510 2154 3512
rect 2154 3510 2188 3512
rect 2188 3510 2223 3512
rect 2223 3510 2257 3512
rect 2257 3510 2292 3512
rect 2292 3510 2326 3512
rect 2326 3510 2361 3512
rect 2361 3510 2395 3512
rect 2395 3510 2430 3512
rect 2430 3510 2464 3512
rect 2464 3510 2499 3512
rect 2499 3510 2533 3512
rect 2533 3510 2568 3512
rect 2568 3510 2602 3512
rect 2602 3510 2637 3512
rect 2637 3510 2671 3512
rect 2671 3510 2706 3512
rect 2706 3510 2740 3512
rect 2740 3510 2775 3512
rect 2775 3510 2809 3512
rect 2809 3510 2844 3512
rect 2844 3510 2878 3512
rect 2878 3510 2913 3512
rect 2913 3510 2947 3512
rect 2947 3510 2982 3512
rect 2982 3510 3016 3512
rect 3016 3510 3051 3512
rect 3051 3510 3085 3512
rect 3085 3510 3120 3512
rect 3120 3510 3154 3512
rect 3154 3510 3189 3512
rect 3189 3510 3223 3512
rect 3223 3510 3258 3512
rect 3258 3510 3292 3512
rect 3292 3510 3327 3512
rect 3327 3510 3361 3512
rect 3361 3510 3396 3512
rect -886 3478 -852 3510
rect -813 3478 -779 3510
rect -740 3478 -706 3510
rect -667 3478 -633 3510
rect -594 3476 3396 3510
rect -594 3442 -572 3476
rect -572 3442 -537 3476
rect -537 3442 -503 3476
rect -503 3442 -468 3476
rect -468 3442 -434 3476
rect -434 3442 -399 3476
rect -399 3442 -365 3476
rect -365 3442 -330 3476
rect -330 3442 -296 3476
rect -296 3442 -261 3476
rect -261 3442 -227 3476
rect -227 3442 -192 3476
rect -192 3442 -158 3476
rect -158 3442 -123 3476
rect -123 3442 -89 3476
rect -89 3442 -54 3476
rect -54 3442 -20 3476
rect -20 3442 15 3476
rect 15 3442 49 3476
rect 49 3442 84 3476
rect 84 3442 118 3476
rect 118 3442 153 3476
rect 153 3442 187 3476
rect 187 3442 222 3476
rect 222 3442 256 3476
rect 256 3442 291 3476
rect 291 3442 325 3476
rect 325 3442 360 3476
rect 360 3442 394 3476
rect 394 3442 429 3476
rect 429 3442 463 3476
rect 463 3442 498 3476
rect 498 3442 532 3476
rect 532 3442 567 3476
rect 567 3442 601 3476
rect 601 3442 636 3476
rect 636 3442 670 3476
rect 670 3442 705 3476
rect 705 3442 739 3476
rect 739 3442 774 3476
rect 774 3442 808 3476
rect 808 3442 843 3476
rect 843 3442 877 3476
rect 877 3442 912 3476
rect 912 3442 946 3476
rect 946 3442 981 3476
rect 981 3442 1015 3476
rect 1015 3442 1050 3476
rect 1050 3442 1084 3476
rect 1084 3442 1119 3476
rect 1119 3442 1153 3476
rect 1153 3442 1188 3476
rect 1188 3442 1222 3476
rect 1222 3442 1257 3476
rect 1257 3442 1291 3476
rect 1291 3442 1326 3476
rect 1326 3442 1360 3476
rect 1360 3442 1395 3476
rect 1395 3442 1429 3476
rect 1429 3442 1464 3476
rect 1464 3442 1498 3476
rect 1498 3442 1533 3476
rect 1533 3442 1567 3476
rect 1567 3442 1602 3476
rect 1602 3442 1636 3476
rect 1636 3442 1671 3476
rect 1671 3442 1705 3476
rect 1705 3442 1740 3476
rect 1740 3442 1774 3476
rect 1774 3442 1809 3476
rect 1809 3442 1843 3476
rect 1843 3442 1878 3476
rect 1878 3442 1912 3476
rect 1912 3442 1947 3476
rect 1947 3442 1981 3476
rect 1981 3442 2016 3476
rect 2016 3442 2050 3476
rect 2050 3442 2085 3476
rect 2085 3442 2119 3476
rect 2119 3442 2154 3476
rect 2154 3442 2188 3476
rect 2188 3442 2223 3476
rect 2223 3442 2257 3476
rect 2257 3442 2292 3476
rect 2292 3442 2326 3476
rect 2326 3442 2361 3476
rect 2361 3442 2395 3476
rect 2395 3442 2430 3476
rect 2430 3442 2464 3476
rect 2464 3442 2499 3476
rect 2499 3442 2533 3476
rect 2533 3442 2568 3476
rect 2568 3442 2602 3476
rect 2602 3442 2637 3476
rect 2637 3442 2671 3476
rect 2671 3442 2706 3476
rect 2706 3442 2740 3476
rect 2740 3442 2775 3476
rect 2775 3442 2809 3476
rect 2809 3442 2844 3476
rect 2844 3442 2878 3476
rect 2878 3442 2913 3476
rect 2913 3442 2947 3476
rect 2947 3442 2982 3476
rect 2982 3442 3016 3476
rect 3016 3442 3051 3476
rect 3051 3442 3085 3476
rect 3085 3442 3120 3476
rect 3120 3442 3154 3476
rect 3154 3442 3189 3476
rect 3189 3442 3223 3476
rect 3223 3442 3258 3476
rect 3258 3442 3292 3476
rect 3292 3442 3327 3476
rect 3327 3442 3361 3476
rect 3361 3442 3396 3476
rect -886 3408 -852 3440
rect -813 3408 -779 3440
rect -740 3408 -706 3440
rect -667 3408 -633 3440
rect -594 3408 3396 3442
rect -886 3406 -882 3408
rect -882 3406 -852 3408
rect -813 3406 -779 3408
rect -740 3406 -710 3408
rect -710 3406 -706 3408
rect -667 3406 -641 3408
rect -641 3406 -633 3408
rect -594 3406 -572 3408
rect -572 3406 -537 3408
rect -537 3406 -503 3408
rect -503 3406 -468 3408
rect -468 3406 -434 3408
rect -434 3406 -399 3408
rect -399 3406 -365 3408
rect -365 3406 -330 3408
rect -330 3406 -296 3408
rect -296 3406 -261 3408
rect -261 3406 -227 3408
rect -227 3406 -192 3408
rect -192 3406 -158 3408
rect -158 3406 -123 3408
rect -123 3406 -89 3408
rect -89 3406 -54 3408
rect -54 3406 -20 3408
rect -20 3406 15 3408
rect 15 3406 49 3408
rect 49 3406 84 3408
rect 84 3406 118 3408
rect 118 3406 153 3408
rect 153 3406 187 3408
rect 187 3406 222 3408
rect 222 3406 256 3408
rect 256 3406 291 3408
rect 291 3406 325 3408
rect 325 3406 360 3408
rect 360 3406 394 3408
rect 394 3406 429 3408
rect 429 3406 463 3408
rect 463 3406 498 3408
rect 498 3406 532 3408
rect 532 3406 567 3408
rect 567 3406 601 3408
rect 601 3406 636 3408
rect 636 3406 670 3408
rect 670 3406 705 3408
rect 705 3406 739 3408
rect 739 3406 774 3408
rect 774 3406 808 3408
rect 808 3406 843 3408
rect 843 3406 877 3408
rect 877 3406 912 3408
rect 912 3406 946 3408
rect 946 3406 981 3408
rect 981 3406 1015 3408
rect 1015 3406 1050 3408
rect 1050 3406 1084 3408
rect 1084 3406 1119 3408
rect 1119 3406 1153 3408
rect 1153 3406 1188 3408
rect 1188 3406 1222 3408
rect 1222 3406 1257 3408
rect 1257 3406 1291 3408
rect 1291 3406 1326 3408
rect 1326 3406 1360 3408
rect 1360 3406 1395 3408
rect 1395 3406 1429 3408
rect 1429 3406 1464 3408
rect 1464 3406 1498 3408
rect 1498 3406 1533 3408
rect 1533 3406 1567 3408
rect 1567 3406 1602 3408
rect 1602 3406 1636 3408
rect 1636 3406 1671 3408
rect 1671 3406 1705 3408
rect 1705 3406 1740 3408
rect 1740 3406 1774 3408
rect 1774 3406 1809 3408
rect 1809 3406 1843 3408
rect 1843 3406 1878 3408
rect 1878 3406 1912 3408
rect 1912 3406 1947 3408
rect 1947 3406 1981 3408
rect 1981 3406 2016 3408
rect 2016 3406 2050 3408
rect 2050 3406 2085 3408
rect 2085 3406 2119 3408
rect 2119 3406 2154 3408
rect 2154 3406 2188 3408
rect 2188 3406 2223 3408
rect 2223 3406 2257 3408
rect 2257 3406 2292 3408
rect 2292 3406 2326 3408
rect 2326 3406 2361 3408
rect 2361 3406 2395 3408
rect 2395 3406 2430 3408
rect 2430 3406 2464 3408
rect 2464 3406 2499 3408
rect 2499 3406 2533 3408
rect 2533 3406 2568 3408
rect 2568 3406 2602 3408
rect 2602 3406 2637 3408
rect 2637 3406 2671 3408
rect 2671 3406 2706 3408
rect 2706 3406 2740 3408
rect 2740 3406 2775 3408
rect 2775 3406 2809 3408
rect 2809 3406 2844 3408
rect 2844 3406 2878 3408
rect 2878 3406 2913 3408
rect 2913 3406 2947 3408
rect 2947 3406 2982 3408
rect 2982 3406 3016 3408
rect 3016 3406 3051 3408
rect 3051 3406 3085 3408
rect 3085 3406 3120 3408
rect 3120 3406 3154 3408
rect 3154 3406 3189 3408
rect 3189 3406 3223 3408
rect 3223 3406 3258 3408
rect 3258 3406 3292 3408
rect 3292 3406 3327 3408
rect 3327 3406 3361 3408
rect 3361 3406 3396 3408
rect 3396 3406 13768 3512
rect -1074 2451 -320 3277
rect -1074 2378 -1040 2412
rect -1002 2378 -968 2412
rect -930 2378 -896 2412
rect -858 2378 -824 2412
rect -786 2378 -752 2412
rect -714 2378 -680 2412
rect -642 2378 -608 2412
rect -570 2378 -536 2412
rect -498 2378 -464 2412
rect -426 2378 -392 2412
rect -354 2378 -320 2412
rect -1074 2305 -1040 2339
rect -1002 2305 -968 2339
rect -930 2305 -896 2339
rect -858 2305 -824 2339
rect -786 2305 -752 2339
rect -714 2305 -680 2339
rect -642 2305 -608 2339
rect -570 2305 -536 2339
rect -498 2305 -464 2339
rect -426 2305 -392 2339
rect -354 2305 -320 2339
rect -1074 2232 -1040 2266
rect -1002 2232 -968 2266
rect -930 2232 -896 2266
rect -858 2232 -824 2266
rect -786 2232 -752 2266
rect -714 2232 -680 2266
rect -642 2232 -608 2266
rect -570 2232 -536 2266
rect -498 2232 -464 2266
rect -426 2232 -392 2266
rect -354 2232 -320 2266
rect -1074 2159 -1040 2193
rect -1002 2159 -968 2193
rect -930 2159 -896 2193
rect -858 2159 -824 2193
rect -786 2159 -752 2193
rect -714 2159 -680 2193
rect -642 2159 -608 2193
rect -570 2159 -536 2193
rect -498 2159 -464 2193
rect -426 2159 -392 2193
rect -354 2159 -320 2193
rect -1074 2086 -1040 2120
rect -1002 2086 -968 2120
rect -930 2086 -896 2120
rect -858 2086 -824 2120
rect -786 2086 -752 2120
rect -714 2086 -680 2120
rect -642 2086 -608 2120
rect -570 2086 -536 2120
rect -498 2086 -464 2120
rect -426 2086 -392 2120
rect -354 2086 -320 2120
rect -1074 2013 -1040 2047
rect -1002 2013 -968 2047
rect -930 2013 -896 2047
rect -858 2013 -824 2047
rect -786 2013 -752 2047
rect -714 2013 -680 2047
rect -642 2013 -608 2047
rect -570 2013 -536 2047
rect -498 2013 -464 2047
rect -426 2013 -392 2047
rect -354 2013 -320 2047
rect -1074 1940 -1040 1974
rect -1002 1940 -968 1974
rect -930 1940 -896 1974
rect -858 1940 -824 1974
rect -786 1940 -752 1974
rect -714 1940 -680 1974
rect -642 1940 -608 1974
rect -570 1940 -536 1974
rect -498 1940 -464 1974
rect -426 1940 -392 1974
rect -354 1940 -320 1974
rect -1074 1867 -1040 1901
rect -1002 1867 -968 1901
rect -930 1867 -896 1901
rect -858 1867 -824 1901
rect -786 1867 -752 1901
rect -714 1867 -680 1901
rect -642 1867 -608 1901
rect -570 1867 -536 1901
rect -498 1867 -464 1901
rect -426 1867 -392 1901
rect -354 1867 -320 1901
rect -1074 1794 -1040 1828
rect -1002 1794 -968 1828
rect -930 1794 -896 1828
rect -858 1794 -824 1828
rect -786 1794 -752 1828
rect -714 1794 -680 1828
rect -642 1794 -608 1828
rect -570 1794 -536 1828
rect -498 1794 -464 1828
rect -426 1794 -392 1828
rect -354 1794 -320 1828
rect -1074 1721 -1040 1755
rect -1002 1721 -968 1755
rect -930 1721 -896 1755
rect -858 1721 -824 1755
rect -786 1721 -752 1755
rect -714 1721 -680 1755
rect -642 1721 -608 1755
rect -570 1721 -536 1755
rect -498 1721 -464 1755
rect -426 1721 -392 1755
rect -354 1721 -320 1755
rect -1074 1648 -1040 1682
rect -1002 1648 -968 1682
rect -930 1648 -896 1682
rect -858 1648 -824 1682
rect -786 1648 -752 1682
rect -714 1648 -680 1682
rect -642 1648 -608 1682
rect -570 1648 -536 1682
rect -498 1648 -464 1682
rect -426 1648 -392 1682
rect -354 1648 -320 1682
rect -1074 1575 -1040 1609
rect -1002 1575 -968 1609
rect -930 1575 -896 1609
rect -858 1575 -824 1609
rect -786 1575 -752 1609
rect -714 1575 -680 1609
rect -642 1575 -608 1609
rect -570 1575 -536 1609
rect -498 1575 -464 1609
rect -426 1575 -392 1609
rect -354 1575 -320 1609
rect -1074 1502 -1040 1536
rect -1002 1502 -968 1536
rect -930 1502 -896 1536
rect -858 1502 -824 1536
rect -786 1502 -752 1536
rect -714 1502 -680 1536
rect -642 1502 -608 1536
rect -570 1502 -536 1536
rect -498 1502 -464 1536
rect -426 1502 -392 1536
rect -354 1502 -320 1536
rect -1074 1429 -1040 1463
rect -1002 1429 -968 1463
rect -930 1429 -896 1463
rect -858 1429 -824 1463
rect -786 1429 -752 1463
rect -714 1429 -680 1463
rect -642 1429 -608 1463
rect -570 1429 -536 1463
rect -498 1429 -464 1463
rect -426 1429 -392 1463
rect -354 1429 -320 1463
rect -1074 1356 -1040 1390
rect -1002 1356 -968 1390
rect -930 1356 -896 1390
rect -858 1356 -824 1390
rect -786 1356 -752 1390
rect -714 1356 -680 1390
rect -642 1356 -608 1390
rect -570 1356 -536 1390
rect -498 1356 -464 1390
rect -426 1356 -392 1390
rect -354 1356 -320 1390
rect -1074 1283 -1040 1317
rect -1002 1283 -968 1317
rect -930 1283 -896 1317
rect -858 1283 -824 1317
rect -786 1283 -752 1317
rect -714 1283 -680 1317
rect -642 1283 -608 1317
rect -570 1283 -536 1317
rect -498 1283 -464 1317
rect -426 1283 -392 1317
rect -354 1283 -320 1317
rect -1074 1210 -1040 1244
rect -1002 1210 -968 1244
rect -930 1210 -896 1244
rect -858 1210 -824 1244
rect -786 1210 -752 1244
rect -714 1210 -680 1244
rect -642 1210 -608 1244
rect -570 1210 -536 1244
rect -498 1210 -464 1244
rect -426 1210 -392 1244
rect -354 1210 -320 1244
rect -1074 1137 -1040 1171
rect -1002 1137 -968 1171
rect -930 1137 -896 1171
rect -858 1137 -824 1171
rect -786 1137 -752 1171
rect -714 1137 -680 1171
rect -642 1137 -608 1171
rect -570 1137 -536 1171
rect -498 1137 -464 1171
rect -426 1137 -392 1171
rect -354 1137 -320 1171
rect -1074 1064 -1040 1098
rect -1002 1064 -968 1098
rect -930 1064 -896 1098
rect -858 1064 -824 1098
rect -786 1064 -752 1098
rect -714 1064 -680 1098
rect -642 1064 -608 1098
rect -570 1064 -536 1098
rect -498 1064 -464 1098
rect -426 1064 -392 1098
rect -354 1064 -320 1098
rect -1074 991 -1040 1025
rect -1002 991 -968 1025
rect -930 991 -896 1025
rect -858 991 -824 1025
rect -786 991 -752 1025
rect -714 991 -680 1025
rect -642 991 -608 1025
rect -570 991 -536 1025
rect -498 991 -464 1025
rect -426 991 -392 1025
rect -354 991 -320 1025
rect -1074 918 -1040 952
rect -1002 918 -968 952
rect -930 918 -896 952
rect -858 918 -824 952
rect -786 918 -752 952
rect -714 918 -680 952
rect -642 918 -608 952
rect -570 918 -536 952
rect -498 918 -464 952
rect -426 918 -392 952
rect -354 918 -320 952
rect -1074 845 -1040 879
rect -1002 845 -968 879
rect -930 845 -896 879
rect -858 845 -824 879
rect -786 845 -752 879
rect -714 845 -680 879
rect -642 845 -608 879
rect -570 845 -536 879
rect -498 845 -464 879
rect -426 845 -392 879
rect -354 845 -320 879
rect -1074 772 -1040 806
rect -1002 772 -968 806
rect -930 772 -896 806
rect -858 772 -824 806
rect -786 772 -752 806
rect -714 772 -680 806
rect -642 772 -608 806
rect -570 772 -536 806
rect -498 772 -464 806
rect -426 772 -392 806
rect -354 772 -320 806
rect -1074 699 -1040 733
rect -1002 699 -968 733
rect -930 699 -896 733
rect -858 699 -824 733
rect -786 699 -752 733
rect -714 699 -680 733
rect -642 699 -608 733
rect -570 699 -536 733
rect -498 699 -464 733
rect -426 699 -392 733
rect -354 699 -320 733
rect -1074 626 -1040 660
rect -1002 626 -968 660
rect -930 626 -896 660
rect -858 626 -824 660
rect -786 626 -752 660
rect -714 626 -680 660
rect -642 626 -608 660
rect -570 626 -536 660
rect -498 626 -464 660
rect -426 626 -392 660
rect -354 626 -320 660
rect -1074 553 -1040 587
rect -1002 553 -968 587
rect -930 553 -896 587
rect -858 553 -824 587
rect -786 553 -752 587
rect -714 553 -680 587
rect -642 553 -608 587
rect -570 553 -536 587
rect -498 553 -464 587
rect -426 553 -392 587
rect -354 553 -320 587
rect -1074 484 -1040 514
rect -1002 484 -968 514
rect -930 484 -896 514
rect -858 484 -824 514
rect -786 484 -752 514
rect -714 484 -680 514
rect -642 484 -608 514
rect -570 484 -536 514
rect -498 484 -464 514
rect -426 484 -392 514
rect -354 484 -320 514
rect -1074 480 -1040 484
rect -1002 480 -968 484
rect -930 480 -896 484
rect -858 480 -824 484
rect -786 480 -752 484
rect -714 480 -680 484
rect -642 480 -608 484
rect -570 480 -536 484
rect -498 480 -464 484
rect -426 480 -392 484
rect -354 480 -320 484
rect -1074 415 -1054 441
rect -1054 415 -1040 441
rect -1002 415 -986 441
rect -986 415 -968 441
rect -930 415 -918 441
rect -918 415 -896 441
rect -858 415 -850 441
rect -850 415 -824 441
rect -786 415 -782 441
rect -782 415 -752 441
rect -1074 407 -1040 415
rect -1002 407 -968 415
rect -930 407 -896 415
rect -858 407 -824 415
rect -786 407 -752 415
rect -714 407 -680 441
rect -642 415 -612 441
rect -612 415 -608 441
rect -570 415 -544 441
rect -544 415 -536 441
rect -498 415 -476 441
rect -476 415 -464 441
rect -426 415 -408 441
rect -408 415 -392 441
rect -354 415 -340 441
rect -340 415 -320 441
rect -642 407 -608 415
rect -570 407 -536 415
rect -498 407 -464 415
rect -426 407 -392 415
rect -354 407 -320 415
rect -1074 346 -1054 368
rect -1054 346 -1040 368
rect -1002 346 -986 368
rect -986 346 -968 368
rect -930 346 -918 368
rect -918 346 -896 368
rect -858 346 -850 368
rect -850 346 -824 368
rect -786 346 -782 368
rect -782 346 -752 368
rect -1074 334 -1040 346
rect -1002 334 -968 346
rect -930 334 -896 346
rect -858 334 -824 346
rect -786 334 -752 346
rect -714 334 -680 368
rect -642 346 -612 368
rect -612 346 -608 368
rect -570 346 -544 368
rect -544 346 -536 368
rect -498 346 -476 368
rect -476 346 -464 368
rect -426 346 -408 368
rect -408 346 -392 368
rect -354 346 -340 368
rect -340 346 -320 368
rect -642 334 -608 346
rect -570 334 -536 346
rect -498 334 -464 346
rect -426 334 -392 346
rect -354 334 -320 346
rect -1074 277 -1054 295
rect -1054 277 -1040 295
rect -1002 277 -986 295
rect -986 277 -968 295
rect -930 277 -918 295
rect -918 277 -896 295
rect -858 277 -850 295
rect -850 277 -824 295
rect -786 277 -782 295
rect -782 277 -752 295
rect -1074 261 -1040 277
rect -1002 261 -968 277
rect -930 261 -896 277
rect -858 261 -824 277
rect -786 261 -752 277
rect -714 261 -680 295
rect -642 277 -612 295
rect -612 277 -608 295
rect -570 277 -544 295
rect -544 277 -536 295
rect -498 277 -476 295
rect -476 277 -464 295
rect -426 277 -408 295
rect -408 277 -392 295
rect -354 277 -340 295
rect -340 277 -320 295
rect -642 261 -608 277
rect -570 261 -536 277
rect -498 261 -464 277
rect -426 261 -392 277
rect -354 261 -320 277
rect -1074 208 -1054 222
rect -1054 208 -1040 222
rect -1002 208 -986 222
rect -986 208 -968 222
rect -930 208 -918 222
rect -918 208 -896 222
rect -858 208 -850 222
rect -850 208 -824 222
rect -786 208 -782 222
rect -782 208 -752 222
rect -1074 188 -1040 208
rect -1002 188 -968 208
rect -930 188 -896 208
rect -858 188 -824 208
rect -786 188 -752 208
rect -714 188 -680 222
rect -642 208 -612 222
rect -612 208 -608 222
rect -570 208 -544 222
rect -544 208 -536 222
rect -498 208 -476 222
rect -476 208 -464 222
rect -426 208 -408 222
rect -408 208 -392 222
rect -354 208 -340 222
rect -340 208 -320 222
rect -642 188 -608 208
rect -570 188 -536 208
rect -498 188 -464 208
rect -426 188 -392 208
rect -354 188 -320 208
rect -1074 139 -1054 149
rect -1054 139 -1040 149
rect -1002 139 -986 149
rect -986 139 -968 149
rect -930 139 -918 149
rect -918 139 -896 149
rect -858 139 -850 149
rect -850 139 -824 149
rect -786 139 -782 149
rect -782 139 -752 149
rect -1074 115 -1040 139
rect -1002 115 -968 139
rect -930 115 -896 139
rect -858 115 -824 139
rect -786 115 -752 139
rect -714 115 -680 149
rect -642 139 -612 149
rect -612 139 -608 149
rect -570 139 -544 149
rect -544 139 -536 149
rect -498 139 -476 149
rect -476 139 -464 149
rect -426 139 -408 149
rect -408 139 -392 149
rect -354 139 -340 149
rect -340 139 -320 149
rect -642 115 -608 139
rect -570 115 -536 139
rect -498 115 -464 139
rect -426 115 -392 139
rect -354 115 -320 139
rect -1074 70 -1054 76
rect -1054 70 -1040 76
rect -1002 70 -986 76
rect -986 70 -968 76
rect -930 70 -918 76
rect -918 70 -896 76
rect -858 70 -850 76
rect -850 70 -824 76
rect -786 70 -782 76
rect -782 70 -752 76
rect -1074 42 -1040 70
rect -1002 42 -968 70
rect -930 42 -896 70
rect -858 42 -824 70
rect -786 42 -752 70
rect -714 42 -680 76
rect -642 70 -612 76
rect -612 70 -608 76
rect -570 70 -544 76
rect -544 70 -536 76
rect -498 70 -476 76
rect -476 70 -464 76
rect -426 70 -408 76
rect -408 70 -392 76
rect -354 70 -340 76
rect -340 70 -320 76
rect -642 42 -608 70
rect -570 42 -536 70
rect -498 42 -464 70
rect -426 42 -392 70
rect -354 42 -320 70
rect -1074 1 -1054 3
rect -1054 1 -1040 3
rect -1002 1 -986 3
rect -986 1 -968 3
rect -930 1 -918 3
rect -918 1 -896 3
rect -858 1 -850 3
rect -850 1 -824 3
rect -786 1 -782 3
rect -782 1 -752 3
rect -1074 -31 -1040 1
rect -1002 -31 -968 1
rect -930 -31 -896 1
rect -858 -31 -824 1
rect -786 -31 -752 1
rect -714 -31 -680 3
rect -642 1 -612 3
rect -612 1 -608 3
rect -570 1 -544 3
rect -544 1 -536 3
rect -498 1 -476 3
rect -476 1 -464 3
rect -426 1 -408 3
rect -408 1 -392 3
rect -354 1 -340 3
rect -340 1 -320 3
rect -642 -31 -608 1
rect -570 -31 -536 1
rect -498 -31 -464 1
rect -426 -31 -392 1
rect -354 -31 -320 1
rect -204 2966 -202 3000
rect -202 2966 -170 3000
rect -132 2966 -100 3000
rect -100 2966 -98 3000
rect -204 2893 -202 2927
rect -202 2893 -170 2927
rect -132 2893 -100 2927
rect -100 2893 -98 2927
rect -204 2820 -202 2854
rect -202 2820 -170 2854
rect -132 2820 -100 2854
rect -100 2820 -98 2854
rect -204 2747 -202 2781
rect -202 2747 -170 2781
rect -132 2747 -100 2781
rect -100 2747 -98 2781
rect -204 2674 -202 2708
rect -202 2674 -170 2708
rect -132 2674 -100 2708
rect -100 2674 -98 2708
rect -204 2601 -202 2635
rect -202 2601 -170 2635
rect -132 2601 -100 2635
rect -100 2601 -98 2635
rect -204 2528 -202 2562
rect -202 2528 -170 2562
rect -132 2528 -100 2562
rect -100 2528 -98 2562
rect -204 2455 -202 2489
rect -202 2455 -170 2489
rect -132 2455 -100 2489
rect -100 2455 -98 2489
rect -204 2382 -202 2416
rect -202 2382 -170 2416
rect -132 2382 -100 2416
rect -100 2382 -98 2416
rect -204 2309 -202 2343
rect -202 2309 -170 2343
rect -132 2309 -100 2343
rect -100 2309 -98 2343
rect -204 2236 -202 2270
rect -202 2236 -170 2270
rect -132 2236 -100 2270
rect -100 2236 -98 2270
rect -204 2163 -202 2197
rect -202 2163 -170 2197
rect -132 2163 -100 2197
rect -100 2163 -98 2197
rect -204 2090 -202 2124
rect -202 2090 -170 2124
rect -132 2090 -100 2124
rect -100 2090 -98 2124
rect -204 2017 -202 2051
rect -202 2017 -170 2051
rect -132 2017 -100 2051
rect -100 2017 -98 2051
rect -204 1944 -202 1978
rect -202 1944 -170 1978
rect -132 1944 -100 1978
rect -100 1944 -98 1978
rect -204 1871 -202 1905
rect -202 1871 -170 1905
rect -132 1871 -100 1905
rect -100 1871 -98 1905
rect -204 1798 -202 1832
rect -202 1798 -170 1832
rect -132 1798 -100 1832
rect -100 1798 -98 1832
rect -204 1725 -202 1759
rect -202 1725 -170 1759
rect -132 1725 -100 1759
rect -100 1725 -98 1759
rect -204 1652 -202 1686
rect -202 1652 -170 1686
rect -132 1652 -100 1686
rect -100 1652 -98 1686
rect -204 1579 -202 1613
rect -202 1579 -170 1613
rect -132 1579 -100 1613
rect -100 1579 -98 1613
rect -204 1506 -202 1540
rect -202 1506 -170 1540
rect -132 1506 -100 1540
rect -100 1506 -98 1540
rect -204 1432 -202 1466
rect -202 1432 -170 1466
rect -132 1432 -100 1466
rect -100 1432 -98 1466
rect -204 1358 -202 1392
rect -202 1358 -170 1392
rect -132 1358 -100 1392
rect -100 1358 -98 1392
rect -204 1284 -202 1318
rect -202 1284 -170 1318
rect -132 1284 -100 1318
rect -100 1284 -98 1318
rect -204 1210 -202 1244
rect -202 1210 -170 1244
rect -132 1210 -100 1244
rect -100 1210 -98 1244
rect -204 1136 -202 1170
rect -202 1136 -170 1170
rect -132 1136 -100 1170
rect -100 1136 -98 1170
rect -204 1062 -202 1096
rect -202 1062 -170 1096
rect -132 1062 -100 1096
rect -100 1062 -98 1096
rect -204 988 -202 1022
rect -202 988 -170 1022
rect -132 988 -100 1022
rect -100 988 -98 1022
rect -204 914 -202 948
rect -202 914 -170 948
rect -132 914 -100 948
rect -100 914 -98 948
rect -204 840 -202 874
rect -202 840 -170 874
rect -132 840 -100 874
rect -100 840 -98 874
rect -204 790 -202 800
rect -202 790 -170 800
rect -132 790 -100 800
rect -100 790 -98 800
rect -204 766 -170 790
rect -132 766 -98 790
rect -204 721 -202 726
rect -202 721 -170 726
rect -132 721 -100 726
rect -100 721 -98 726
rect -204 692 -170 721
rect -132 692 -98 721
rect -204 618 -170 652
rect -132 618 -98 652
rect -204 548 -170 578
rect -132 548 -98 578
rect -204 544 -202 548
rect -202 544 -170 548
rect -132 544 -100 548
rect -100 544 -98 548
rect -204 479 -170 504
rect -132 479 -98 504
rect -204 470 -202 479
rect -202 470 -170 479
rect -132 470 -100 479
rect -100 470 -98 479
rect -204 410 -170 430
rect -132 410 -98 430
rect -204 396 -202 410
rect -202 396 -170 410
rect -132 396 -100 410
rect -100 396 -98 410
rect -204 341 -170 356
rect -132 341 -98 356
rect -204 322 -202 341
rect -202 322 -170 341
rect -132 322 -100 341
rect -100 322 -98 341
rect -204 272 -170 282
rect -132 272 -98 282
rect -204 248 -202 272
rect -202 248 -170 272
rect -132 248 -100 272
rect -100 248 -98 272
rect -204 203 -170 208
rect -132 203 -98 208
rect -204 174 -202 203
rect -202 174 -170 203
rect -132 174 -100 203
rect -100 174 -98 203
rect -204 100 -202 134
rect -202 100 -170 134
rect -132 100 -100 134
rect -100 100 -98 134
rect 208 2966 210 3000
rect 210 2966 242 3000
rect 280 2966 312 3000
rect 312 2966 314 3000
rect 208 2893 210 2927
rect 210 2893 242 2927
rect 280 2893 312 2927
rect 312 2893 314 2927
rect 208 2820 210 2854
rect 210 2820 242 2854
rect 280 2820 312 2854
rect 312 2820 314 2854
rect 208 2747 210 2781
rect 210 2747 242 2781
rect 280 2747 312 2781
rect 312 2747 314 2781
rect 208 2674 210 2708
rect 210 2674 242 2708
rect 280 2674 312 2708
rect 312 2674 314 2708
rect 208 2601 210 2635
rect 210 2601 242 2635
rect 280 2601 312 2635
rect 312 2601 314 2635
rect 208 2528 210 2562
rect 210 2528 242 2562
rect 280 2528 312 2562
rect 312 2528 314 2562
rect 208 2455 210 2489
rect 210 2455 242 2489
rect 280 2455 312 2489
rect 312 2455 314 2489
rect 208 2382 210 2416
rect 210 2382 242 2416
rect 280 2382 312 2416
rect 312 2382 314 2416
rect 208 2309 210 2343
rect 210 2309 242 2343
rect 280 2309 312 2343
rect 312 2309 314 2343
rect 208 2236 210 2270
rect 210 2236 242 2270
rect 280 2236 312 2270
rect 312 2236 314 2270
rect 208 2163 210 2197
rect 210 2163 242 2197
rect 280 2163 312 2197
rect 312 2163 314 2197
rect 208 2090 210 2124
rect 210 2090 242 2124
rect 280 2090 312 2124
rect 312 2090 314 2124
rect 208 2017 210 2051
rect 210 2017 242 2051
rect 280 2017 312 2051
rect 312 2017 314 2051
rect 208 1944 210 1978
rect 210 1944 242 1978
rect 280 1944 312 1978
rect 312 1944 314 1978
rect 208 1871 210 1905
rect 210 1871 242 1905
rect 280 1871 312 1905
rect 312 1871 314 1905
rect 208 1798 210 1832
rect 210 1798 242 1832
rect 280 1798 312 1832
rect 312 1798 314 1832
rect 208 1725 210 1759
rect 210 1725 242 1759
rect 280 1725 312 1759
rect 312 1725 314 1759
rect 208 1652 210 1686
rect 210 1652 242 1686
rect 280 1652 312 1686
rect 312 1652 314 1686
rect 208 1579 210 1613
rect 210 1579 242 1613
rect 280 1579 312 1613
rect 312 1579 314 1613
rect 208 1506 210 1540
rect 210 1506 242 1540
rect 280 1506 312 1540
rect 312 1506 314 1540
rect 208 1432 210 1466
rect 210 1432 242 1466
rect 280 1432 312 1466
rect 312 1432 314 1466
rect 208 1358 210 1392
rect 210 1358 242 1392
rect 280 1358 312 1392
rect 312 1358 314 1392
rect 208 1284 210 1318
rect 210 1284 242 1318
rect 280 1284 312 1318
rect 312 1284 314 1318
rect 208 1210 210 1244
rect 210 1210 242 1244
rect 280 1210 312 1244
rect 312 1210 314 1244
rect 208 1136 210 1170
rect 210 1136 242 1170
rect 280 1136 312 1170
rect 312 1136 314 1170
rect 208 1062 210 1096
rect 210 1062 242 1096
rect 280 1062 312 1096
rect 312 1062 314 1096
rect 208 988 210 1022
rect 210 988 242 1022
rect 280 988 312 1022
rect 312 988 314 1022
rect 208 914 210 948
rect 210 914 242 948
rect 280 914 312 948
rect 312 914 314 948
rect 208 840 210 874
rect 210 840 242 874
rect 280 840 312 874
rect 312 840 314 874
rect 208 790 210 800
rect 210 790 242 800
rect 280 790 312 800
rect 312 790 314 800
rect 208 766 242 790
rect 280 766 314 790
rect 208 721 210 726
rect 210 721 242 726
rect 280 721 312 726
rect 312 721 314 726
rect 208 692 242 721
rect 280 692 314 721
rect 208 618 242 652
rect 280 618 314 652
rect 208 548 242 578
rect 280 548 314 578
rect 208 544 210 548
rect 210 544 242 548
rect 280 544 312 548
rect 312 544 314 548
rect 208 479 242 504
rect 280 479 314 504
rect 208 470 210 479
rect 210 470 242 479
rect 280 470 312 479
rect 312 470 314 479
rect 208 410 242 430
rect 280 410 314 430
rect 208 396 210 410
rect 210 396 242 410
rect 280 396 312 410
rect 312 396 314 410
rect 208 341 242 356
rect 280 341 314 356
rect 208 322 210 341
rect 210 322 242 341
rect 280 322 312 341
rect 312 322 314 341
rect 208 272 242 282
rect 280 272 314 282
rect 208 248 210 272
rect 210 248 242 272
rect 280 248 312 272
rect 312 248 314 272
rect 208 203 242 208
rect 280 203 314 208
rect 208 174 210 203
rect 210 174 242 203
rect 280 174 312 203
rect 312 174 314 203
rect 208 100 210 134
rect 210 100 242 134
rect 280 100 312 134
rect 312 100 314 134
rect 620 2966 622 3000
rect 622 2966 654 3000
rect 692 2966 724 3000
rect 724 2966 726 3000
rect 620 2893 622 2927
rect 622 2893 654 2927
rect 692 2893 724 2927
rect 724 2893 726 2927
rect 620 2820 622 2854
rect 622 2820 654 2854
rect 692 2820 724 2854
rect 724 2820 726 2854
rect 620 2747 622 2781
rect 622 2747 654 2781
rect 692 2747 724 2781
rect 724 2747 726 2781
rect 620 2674 622 2708
rect 622 2674 654 2708
rect 692 2674 724 2708
rect 724 2674 726 2708
rect 620 2601 622 2635
rect 622 2601 654 2635
rect 692 2601 724 2635
rect 724 2601 726 2635
rect 620 2528 622 2562
rect 622 2528 654 2562
rect 692 2528 724 2562
rect 724 2528 726 2562
rect 620 2455 622 2489
rect 622 2455 654 2489
rect 692 2455 724 2489
rect 724 2455 726 2489
rect 620 2382 622 2416
rect 622 2382 654 2416
rect 692 2382 724 2416
rect 724 2382 726 2416
rect 620 2309 622 2343
rect 622 2309 654 2343
rect 692 2309 724 2343
rect 724 2309 726 2343
rect 620 2236 622 2270
rect 622 2236 654 2270
rect 692 2236 724 2270
rect 724 2236 726 2270
rect 620 2163 622 2197
rect 622 2163 654 2197
rect 692 2163 724 2197
rect 724 2163 726 2197
rect 620 2090 622 2124
rect 622 2090 654 2124
rect 692 2090 724 2124
rect 724 2090 726 2124
rect 620 2017 622 2051
rect 622 2017 654 2051
rect 692 2017 724 2051
rect 724 2017 726 2051
rect 620 1944 622 1978
rect 622 1944 654 1978
rect 692 1944 724 1978
rect 724 1944 726 1978
rect 620 1871 622 1905
rect 622 1871 654 1905
rect 692 1871 724 1905
rect 724 1871 726 1905
rect 620 1798 622 1832
rect 622 1798 654 1832
rect 692 1798 724 1832
rect 724 1798 726 1832
rect 620 1725 622 1759
rect 622 1725 654 1759
rect 692 1725 724 1759
rect 724 1725 726 1759
rect 620 1652 622 1686
rect 622 1652 654 1686
rect 692 1652 724 1686
rect 724 1652 726 1686
rect 620 1579 622 1613
rect 622 1579 654 1613
rect 692 1579 724 1613
rect 724 1579 726 1613
rect 620 1506 622 1540
rect 622 1506 654 1540
rect 692 1506 724 1540
rect 724 1506 726 1540
rect 620 1432 622 1466
rect 622 1432 654 1466
rect 692 1432 724 1466
rect 724 1432 726 1466
rect 620 1358 622 1392
rect 622 1358 654 1392
rect 692 1358 724 1392
rect 724 1358 726 1392
rect 620 1284 622 1318
rect 622 1284 654 1318
rect 692 1284 724 1318
rect 724 1284 726 1318
rect 620 1210 622 1244
rect 622 1210 654 1244
rect 692 1210 724 1244
rect 724 1210 726 1244
rect 620 1136 622 1170
rect 622 1136 654 1170
rect 692 1136 724 1170
rect 724 1136 726 1170
rect 620 1062 622 1096
rect 622 1062 654 1096
rect 692 1062 724 1096
rect 724 1062 726 1096
rect 620 988 622 1022
rect 622 988 654 1022
rect 692 988 724 1022
rect 724 988 726 1022
rect 620 914 622 948
rect 622 914 654 948
rect 692 914 724 948
rect 724 914 726 948
rect 620 840 622 874
rect 622 840 654 874
rect 692 840 724 874
rect 724 840 726 874
rect 620 790 622 800
rect 622 790 654 800
rect 692 790 724 800
rect 724 790 726 800
rect 620 766 654 790
rect 692 766 726 790
rect 620 721 622 726
rect 622 721 654 726
rect 692 721 724 726
rect 724 721 726 726
rect 620 692 654 721
rect 692 692 726 721
rect 620 618 654 652
rect 692 618 726 652
rect 620 548 654 578
rect 692 548 726 578
rect 620 544 622 548
rect 622 544 654 548
rect 692 544 724 548
rect 724 544 726 548
rect 620 479 654 504
rect 692 479 726 504
rect 620 470 622 479
rect 622 470 654 479
rect 692 470 724 479
rect 724 470 726 479
rect 620 410 654 430
rect 692 410 726 430
rect 620 396 622 410
rect 622 396 654 410
rect 692 396 724 410
rect 724 396 726 410
rect 620 341 654 356
rect 692 341 726 356
rect 620 322 622 341
rect 622 322 654 341
rect 692 322 724 341
rect 724 322 726 341
rect 620 272 654 282
rect 692 272 726 282
rect 620 248 622 272
rect 622 248 654 272
rect 692 248 724 272
rect 724 248 726 272
rect 620 203 654 208
rect 692 203 726 208
rect 620 174 622 203
rect 622 174 654 203
rect 692 174 724 203
rect 724 174 726 203
rect 620 100 622 134
rect 622 100 654 134
rect 692 100 724 134
rect 724 100 726 134
rect 1032 2966 1034 3000
rect 1034 2966 1066 3000
rect 1104 2966 1136 3000
rect 1136 2966 1138 3000
rect 1032 2893 1034 2927
rect 1034 2893 1066 2927
rect 1104 2893 1136 2927
rect 1136 2893 1138 2927
rect 1032 2820 1034 2854
rect 1034 2820 1066 2854
rect 1104 2820 1136 2854
rect 1136 2820 1138 2854
rect 1032 2747 1034 2781
rect 1034 2747 1066 2781
rect 1104 2747 1136 2781
rect 1136 2747 1138 2781
rect 1032 2674 1034 2708
rect 1034 2674 1066 2708
rect 1104 2674 1136 2708
rect 1136 2674 1138 2708
rect 1032 2601 1034 2635
rect 1034 2601 1066 2635
rect 1104 2601 1136 2635
rect 1136 2601 1138 2635
rect 1032 2528 1034 2562
rect 1034 2528 1066 2562
rect 1104 2528 1136 2562
rect 1136 2528 1138 2562
rect 1032 2455 1034 2489
rect 1034 2455 1066 2489
rect 1104 2455 1136 2489
rect 1136 2455 1138 2489
rect 1032 2382 1034 2416
rect 1034 2382 1066 2416
rect 1104 2382 1136 2416
rect 1136 2382 1138 2416
rect 1032 2309 1034 2343
rect 1034 2309 1066 2343
rect 1104 2309 1136 2343
rect 1136 2309 1138 2343
rect 1032 2236 1034 2270
rect 1034 2236 1066 2270
rect 1104 2236 1136 2270
rect 1136 2236 1138 2270
rect 1032 2163 1034 2197
rect 1034 2163 1066 2197
rect 1104 2163 1136 2197
rect 1136 2163 1138 2197
rect 1032 2090 1034 2124
rect 1034 2090 1066 2124
rect 1104 2090 1136 2124
rect 1136 2090 1138 2124
rect 1032 2017 1034 2051
rect 1034 2017 1066 2051
rect 1104 2017 1136 2051
rect 1136 2017 1138 2051
rect 1032 1944 1034 1978
rect 1034 1944 1066 1978
rect 1104 1944 1136 1978
rect 1136 1944 1138 1978
rect 1032 1871 1034 1905
rect 1034 1871 1066 1905
rect 1104 1871 1136 1905
rect 1136 1871 1138 1905
rect 1032 1798 1034 1832
rect 1034 1798 1066 1832
rect 1104 1798 1136 1832
rect 1136 1798 1138 1832
rect 1032 1725 1034 1759
rect 1034 1725 1066 1759
rect 1104 1725 1136 1759
rect 1136 1725 1138 1759
rect 1032 1652 1034 1686
rect 1034 1652 1066 1686
rect 1104 1652 1136 1686
rect 1136 1652 1138 1686
rect 1032 1579 1034 1613
rect 1034 1579 1066 1613
rect 1104 1579 1136 1613
rect 1136 1579 1138 1613
rect 1032 1506 1034 1540
rect 1034 1506 1066 1540
rect 1104 1506 1136 1540
rect 1136 1506 1138 1540
rect 1032 1432 1034 1466
rect 1034 1432 1066 1466
rect 1104 1432 1136 1466
rect 1136 1432 1138 1466
rect 1032 1358 1034 1392
rect 1034 1358 1066 1392
rect 1104 1358 1136 1392
rect 1136 1358 1138 1392
rect 1032 1284 1034 1318
rect 1034 1284 1066 1318
rect 1104 1284 1136 1318
rect 1136 1284 1138 1318
rect 1032 1210 1034 1244
rect 1034 1210 1066 1244
rect 1104 1210 1136 1244
rect 1136 1210 1138 1244
rect 1032 1136 1034 1170
rect 1034 1136 1066 1170
rect 1104 1136 1136 1170
rect 1136 1136 1138 1170
rect 1032 1062 1034 1096
rect 1034 1062 1066 1096
rect 1104 1062 1136 1096
rect 1136 1062 1138 1096
rect 1032 988 1034 1022
rect 1034 988 1066 1022
rect 1104 988 1136 1022
rect 1136 988 1138 1022
rect 1032 914 1034 948
rect 1034 914 1066 948
rect 1104 914 1136 948
rect 1136 914 1138 948
rect 1032 840 1034 874
rect 1034 840 1066 874
rect 1104 840 1136 874
rect 1136 840 1138 874
rect 1032 790 1034 800
rect 1034 790 1066 800
rect 1104 790 1136 800
rect 1136 790 1138 800
rect 1032 766 1066 790
rect 1104 766 1138 790
rect 1032 721 1034 726
rect 1034 721 1066 726
rect 1104 721 1136 726
rect 1136 721 1138 726
rect 1032 692 1066 721
rect 1104 692 1138 721
rect 1032 618 1066 652
rect 1104 618 1138 652
rect 1032 548 1066 578
rect 1104 548 1138 578
rect 1032 544 1034 548
rect 1034 544 1066 548
rect 1104 544 1136 548
rect 1136 544 1138 548
rect 1032 479 1066 504
rect 1104 479 1138 504
rect 1032 470 1034 479
rect 1034 470 1066 479
rect 1104 470 1136 479
rect 1136 470 1138 479
rect 1032 410 1066 430
rect 1104 410 1138 430
rect 1032 396 1034 410
rect 1034 396 1066 410
rect 1104 396 1136 410
rect 1136 396 1138 410
rect 1032 341 1066 356
rect 1104 341 1138 356
rect 1032 322 1034 341
rect 1034 322 1066 341
rect 1104 322 1136 341
rect 1136 322 1138 341
rect 1032 272 1066 282
rect 1104 272 1138 282
rect 1032 248 1034 272
rect 1034 248 1066 272
rect 1104 248 1136 272
rect 1136 248 1138 272
rect 1032 203 1066 208
rect 1104 203 1138 208
rect 1032 174 1034 203
rect 1034 174 1066 203
rect 1104 174 1136 203
rect 1136 174 1138 203
rect 1032 100 1034 134
rect 1034 100 1066 134
rect 1104 100 1136 134
rect 1136 100 1138 134
rect 1444 2966 1446 3000
rect 1446 2966 1478 3000
rect 1516 2966 1548 3000
rect 1548 2966 1550 3000
rect 1444 2893 1446 2927
rect 1446 2893 1478 2927
rect 1516 2893 1548 2927
rect 1548 2893 1550 2927
rect 1444 2820 1446 2854
rect 1446 2820 1478 2854
rect 1516 2820 1548 2854
rect 1548 2820 1550 2854
rect 1444 2747 1446 2781
rect 1446 2747 1478 2781
rect 1516 2747 1548 2781
rect 1548 2747 1550 2781
rect 1444 2674 1446 2708
rect 1446 2674 1478 2708
rect 1516 2674 1548 2708
rect 1548 2674 1550 2708
rect 1444 2601 1446 2635
rect 1446 2601 1478 2635
rect 1516 2601 1548 2635
rect 1548 2601 1550 2635
rect 1444 2528 1446 2562
rect 1446 2528 1478 2562
rect 1516 2528 1548 2562
rect 1548 2528 1550 2562
rect 1444 2455 1446 2489
rect 1446 2455 1478 2489
rect 1516 2455 1548 2489
rect 1548 2455 1550 2489
rect 1444 2382 1446 2416
rect 1446 2382 1478 2416
rect 1516 2382 1548 2416
rect 1548 2382 1550 2416
rect 1444 2309 1446 2343
rect 1446 2309 1478 2343
rect 1516 2309 1548 2343
rect 1548 2309 1550 2343
rect 1444 2236 1446 2270
rect 1446 2236 1478 2270
rect 1516 2236 1548 2270
rect 1548 2236 1550 2270
rect 1444 2163 1446 2197
rect 1446 2163 1478 2197
rect 1516 2163 1548 2197
rect 1548 2163 1550 2197
rect 1444 2090 1446 2124
rect 1446 2090 1478 2124
rect 1516 2090 1548 2124
rect 1548 2090 1550 2124
rect 1444 2017 1446 2051
rect 1446 2017 1478 2051
rect 1516 2017 1548 2051
rect 1548 2017 1550 2051
rect 1444 1944 1446 1978
rect 1446 1944 1478 1978
rect 1516 1944 1548 1978
rect 1548 1944 1550 1978
rect 1444 1871 1446 1905
rect 1446 1871 1478 1905
rect 1516 1871 1548 1905
rect 1548 1871 1550 1905
rect 1444 1798 1446 1832
rect 1446 1798 1478 1832
rect 1516 1798 1548 1832
rect 1548 1798 1550 1832
rect 1444 1725 1446 1759
rect 1446 1725 1478 1759
rect 1516 1725 1548 1759
rect 1548 1725 1550 1759
rect 1444 1652 1446 1686
rect 1446 1652 1478 1686
rect 1516 1652 1548 1686
rect 1548 1652 1550 1686
rect 1444 1579 1446 1613
rect 1446 1579 1478 1613
rect 1516 1579 1548 1613
rect 1548 1579 1550 1613
rect 1444 1506 1446 1540
rect 1446 1506 1478 1540
rect 1516 1506 1548 1540
rect 1548 1506 1550 1540
rect 1444 1432 1446 1466
rect 1446 1432 1478 1466
rect 1516 1432 1548 1466
rect 1548 1432 1550 1466
rect 1444 1358 1446 1392
rect 1446 1358 1478 1392
rect 1516 1358 1548 1392
rect 1548 1358 1550 1392
rect 1444 1284 1446 1318
rect 1446 1284 1478 1318
rect 1516 1284 1548 1318
rect 1548 1284 1550 1318
rect 1444 1210 1446 1244
rect 1446 1210 1478 1244
rect 1516 1210 1548 1244
rect 1548 1210 1550 1244
rect 1444 1136 1446 1170
rect 1446 1136 1478 1170
rect 1516 1136 1548 1170
rect 1548 1136 1550 1170
rect 1444 1062 1446 1096
rect 1446 1062 1478 1096
rect 1516 1062 1548 1096
rect 1548 1062 1550 1096
rect 1444 988 1446 1022
rect 1446 988 1478 1022
rect 1516 988 1548 1022
rect 1548 988 1550 1022
rect 1444 914 1446 948
rect 1446 914 1478 948
rect 1516 914 1548 948
rect 1548 914 1550 948
rect 1444 840 1446 874
rect 1446 840 1478 874
rect 1516 840 1548 874
rect 1548 840 1550 874
rect 1444 790 1446 800
rect 1446 790 1478 800
rect 1516 790 1548 800
rect 1548 790 1550 800
rect 1444 766 1478 790
rect 1516 766 1550 790
rect 1444 721 1446 726
rect 1446 721 1478 726
rect 1516 721 1548 726
rect 1548 721 1550 726
rect 1444 692 1478 721
rect 1516 692 1550 721
rect 1444 618 1478 652
rect 1516 618 1550 652
rect 1444 548 1478 578
rect 1516 548 1550 578
rect 1444 544 1446 548
rect 1446 544 1478 548
rect 1516 544 1548 548
rect 1548 544 1550 548
rect 1444 479 1478 504
rect 1516 479 1550 504
rect 1444 470 1446 479
rect 1446 470 1478 479
rect 1516 470 1548 479
rect 1548 470 1550 479
rect 1444 410 1478 430
rect 1516 410 1550 430
rect 1444 396 1446 410
rect 1446 396 1478 410
rect 1516 396 1548 410
rect 1548 396 1550 410
rect 1444 341 1478 356
rect 1516 341 1550 356
rect 1444 322 1446 341
rect 1446 322 1478 341
rect 1516 322 1548 341
rect 1548 322 1550 341
rect 1444 272 1478 282
rect 1516 272 1550 282
rect 1444 248 1446 272
rect 1446 248 1478 272
rect 1516 248 1548 272
rect 1548 248 1550 272
rect 1444 203 1478 208
rect 1516 203 1550 208
rect 1444 174 1446 203
rect 1446 174 1478 203
rect 1516 174 1548 203
rect 1548 174 1550 203
rect 1444 100 1446 134
rect 1446 100 1478 134
rect 1516 100 1548 134
rect 1548 100 1550 134
rect 1856 2966 1858 3000
rect 1858 2966 1890 3000
rect 1928 2966 1960 3000
rect 1960 2966 1962 3000
rect 1856 2893 1858 2927
rect 1858 2893 1890 2927
rect 1928 2893 1960 2927
rect 1960 2893 1962 2927
rect 1856 2820 1858 2854
rect 1858 2820 1890 2854
rect 1928 2820 1960 2854
rect 1960 2820 1962 2854
rect 1856 2747 1858 2781
rect 1858 2747 1890 2781
rect 1928 2747 1960 2781
rect 1960 2747 1962 2781
rect 1856 2674 1858 2708
rect 1858 2674 1890 2708
rect 1928 2674 1960 2708
rect 1960 2674 1962 2708
rect 1856 2601 1858 2635
rect 1858 2601 1890 2635
rect 1928 2601 1960 2635
rect 1960 2601 1962 2635
rect 1856 2528 1858 2562
rect 1858 2528 1890 2562
rect 1928 2528 1960 2562
rect 1960 2528 1962 2562
rect 1856 2455 1858 2489
rect 1858 2455 1890 2489
rect 1928 2455 1960 2489
rect 1960 2455 1962 2489
rect 1856 2382 1858 2416
rect 1858 2382 1890 2416
rect 1928 2382 1960 2416
rect 1960 2382 1962 2416
rect 1856 2309 1858 2343
rect 1858 2309 1890 2343
rect 1928 2309 1960 2343
rect 1960 2309 1962 2343
rect 1856 2236 1858 2270
rect 1858 2236 1890 2270
rect 1928 2236 1960 2270
rect 1960 2236 1962 2270
rect 1856 2163 1858 2197
rect 1858 2163 1890 2197
rect 1928 2163 1960 2197
rect 1960 2163 1962 2197
rect 1856 2090 1858 2124
rect 1858 2090 1890 2124
rect 1928 2090 1960 2124
rect 1960 2090 1962 2124
rect 1856 2017 1858 2051
rect 1858 2017 1890 2051
rect 1928 2017 1960 2051
rect 1960 2017 1962 2051
rect 1856 1944 1858 1978
rect 1858 1944 1890 1978
rect 1928 1944 1960 1978
rect 1960 1944 1962 1978
rect 1856 1871 1858 1905
rect 1858 1871 1890 1905
rect 1928 1871 1960 1905
rect 1960 1871 1962 1905
rect 1856 1798 1858 1832
rect 1858 1798 1890 1832
rect 1928 1798 1960 1832
rect 1960 1798 1962 1832
rect 1856 1725 1858 1759
rect 1858 1725 1890 1759
rect 1928 1725 1960 1759
rect 1960 1725 1962 1759
rect 1856 1652 1858 1686
rect 1858 1652 1890 1686
rect 1928 1652 1960 1686
rect 1960 1652 1962 1686
rect 1856 1579 1858 1613
rect 1858 1579 1890 1613
rect 1928 1579 1960 1613
rect 1960 1579 1962 1613
rect 1856 1506 1858 1540
rect 1858 1506 1890 1540
rect 1928 1506 1960 1540
rect 1960 1506 1962 1540
rect 1856 1432 1858 1466
rect 1858 1432 1890 1466
rect 1928 1432 1960 1466
rect 1960 1432 1962 1466
rect 1856 1358 1858 1392
rect 1858 1358 1890 1392
rect 1928 1358 1960 1392
rect 1960 1358 1962 1392
rect 1856 1284 1858 1318
rect 1858 1284 1890 1318
rect 1928 1284 1960 1318
rect 1960 1284 1962 1318
rect 1856 1210 1858 1244
rect 1858 1210 1890 1244
rect 1928 1210 1960 1244
rect 1960 1210 1962 1244
rect 1856 1136 1858 1170
rect 1858 1136 1890 1170
rect 1928 1136 1960 1170
rect 1960 1136 1962 1170
rect 1856 1062 1858 1096
rect 1858 1062 1890 1096
rect 1928 1062 1960 1096
rect 1960 1062 1962 1096
rect 1856 988 1858 1022
rect 1858 988 1890 1022
rect 1928 988 1960 1022
rect 1960 988 1962 1022
rect 1856 914 1858 948
rect 1858 914 1890 948
rect 1928 914 1960 948
rect 1960 914 1962 948
rect 1856 840 1858 874
rect 1858 840 1890 874
rect 1928 840 1960 874
rect 1960 840 1962 874
rect 1856 790 1858 800
rect 1858 790 1890 800
rect 1928 790 1960 800
rect 1960 790 1962 800
rect 1856 766 1890 790
rect 1928 766 1962 790
rect 1856 721 1858 726
rect 1858 721 1890 726
rect 1928 721 1960 726
rect 1960 721 1962 726
rect 1856 692 1890 721
rect 1928 692 1962 721
rect 1856 618 1890 652
rect 1928 618 1962 652
rect 1856 548 1890 578
rect 1928 548 1962 578
rect 1856 544 1858 548
rect 1858 544 1890 548
rect 1928 544 1960 548
rect 1960 544 1962 548
rect 1856 479 1890 504
rect 1928 479 1962 504
rect 1856 470 1858 479
rect 1858 470 1890 479
rect 1928 470 1960 479
rect 1960 470 1962 479
rect 1856 410 1890 430
rect 1928 410 1962 430
rect 1856 396 1858 410
rect 1858 396 1890 410
rect 1928 396 1960 410
rect 1960 396 1962 410
rect 1856 341 1890 356
rect 1928 341 1962 356
rect 1856 322 1858 341
rect 1858 322 1890 341
rect 1928 322 1960 341
rect 1960 322 1962 341
rect 1856 272 1890 282
rect 1928 272 1962 282
rect 1856 248 1858 272
rect 1858 248 1890 272
rect 1928 248 1960 272
rect 1960 248 1962 272
rect 1856 203 1890 208
rect 1928 203 1962 208
rect 1856 174 1858 203
rect 1858 174 1890 203
rect 1928 174 1960 203
rect 1960 174 1962 203
rect 1856 100 1858 134
rect 1858 100 1890 134
rect 1928 100 1960 134
rect 1960 100 1962 134
rect 2268 2966 2270 3000
rect 2270 2966 2302 3000
rect 2340 2966 2372 3000
rect 2372 2966 2374 3000
rect 2268 2893 2270 2927
rect 2270 2893 2302 2927
rect 2340 2893 2372 2927
rect 2372 2893 2374 2927
rect 2268 2820 2270 2854
rect 2270 2820 2302 2854
rect 2340 2820 2372 2854
rect 2372 2820 2374 2854
rect 2268 2747 2270 2781
rect 2270 2747 2302 2781
rect 2340 2747 2372 2781
rect 2372 2747 2374 2781
rect 2268 2674 2270 2708
rect 2270 2674 2302 2708
rect 2340 2674 2372 2708
rect 2372 2674 2374 2708
rect 2268 2601 2270 2635
rect 2270 2601 2302 2635
rect 2340 2601 2372 2635
rect 2372 2601 2374 2635
rect 2268 2528 2270 2562
rect 2270 2528 2302 2562
rect 2340 2528 2372 2562
rect 2372 2528 2374 2562
rect 2268 2455 2270 2489
rect 2270 2455 2302 2489
rect 2340 2455 2372 2489
rect 2372 2455 2374 2489
rect 2268 2382 2270 2416
rect 2270 2382 2302 2416
rect 2340 2382 2372 2416
rect 2372 2382 2374 2416
rect 2268 2309 2270 2343
rect 2270 2309 2302 2343
rect 2340 2309 2372 2343
rect 2372 2309 2374 2343
rect 2268 2236 2270 2270
rect 2270 2236 2302 2270
rect 2340 2236 2372 2270
rect 2372 2236 2374 2270
rect 2268 2163 2270 2197
rect 2270 2163 2302 2197
rect 2340 2163 2372 2197
rect 2372 2163 2374 2197
rect 2268 2090 2270 2124
rect 2270 2090 2302 2124
rect 2340 2090 2372 2124
rect 2372 2090 2374 2124
rect 2268 2017 2270 2051
rect 2270 2017 2302 2051
rect 2340 2017 2372 2051
rect 2372 2017 2374 2051
rect 2268 1944 2270 1978
rect 2270 1944 2302 1978
rect 2340 1944 2372 1978
rect 2372 1944 2374 1978
rect 2268 1871 2270 1905
rect 2270 1871 2302 1905
rect 2340 1871 2372 1905
rect 2372 1871 2374 1905
rect 2268 1798 2270 1832
rect 2270 1798 2302 1832
rect 2340 1798 2372 1832
rect 2372 1798 2374 1832
rect 2268 1725 2270 1759
rect 2270 1725 2302 1759
rect 2340 1725 2372 1759
rect 2372 1725 2374 1759
rect 2268 1652 2270 1686
rect 2270 1652 2302 1686
rect 2340 1652 2372 1686
rect 2372 1652 2374 1686
rect 2268 1579 2270 1613
rect 2270 1579 2302 1613
rect 2340 1579 2372 1613
rect 2372 1579 2374 1613
rect 2268 1506 2270 1540
rect 2270 1506 2302 1540
rect 2340 1506 2372 1540
rect 2372 1506 2374 1540
rect 2268 1432 2270 1466
rect 2270 1432 2302 1466
rect 2340 1432 2372 1466
rect 2372 1432 2374 1466
rect 2268 1358 2270 1392
rect 2270 1358 2302 1392
rect 2340 1358 2372 1392
rect 2372 1358 2374 1392
rect 2268 1284 2270 1318
rect 2270 1284 2302 1318
rect 2340 1284 2372 1318
rect 2372 1284 2374 1318
rect 2268 1210 2270 1244
rect 2270 1210 2302 1244
rect 2340 1210 2372 1244
rect 2372 1210 2374 1244
rect 2268 1136 2270 1170
rect 2270 1136 2302 1170
rect 2340 1136 2372 1170
rect 2372 1136 2374 1170
rect 2268 1062 2270 1096
rect 2270 1062 2302 1096
rect 2340 1062 2372 1096
rect 2372 1062 2374 1096
rect 2268 988 2270 1022
rect 2270 988 2302 1022
rect 2340 988 2372 1022
rect 2372 988 2374 1022
rect 2268 914 2270 948
rect 2270 914 2302 948
rect 2340 914 2372 948
rect 2372 914 2374 948
rect 2268 840 2270 874
rect 2270 840 2302 874
rect 2340 840 2372 874
rect 2372 840 2374 874
rect 2268 790 2270 800
rect 2270 790 2302 800
rect 2340 790 2372 800
rect 2372 790 2374 800
rect 2268 766 2302 790
rect 2340 766 2374 790
rect 2268 721 2270 726
rect 2270 721 2302 726
rect 2340 721 2372 726
rect 2372 721 2374 726
rect 2268 692 2302 721
rect 2340 692 2374 721
rect 2268 618 2302 652
rect 2340 618 2374 652
rect 2268 548 2302 578
rect 2340 548 2374 578
rect 2268 544 2270 548
rect 2270 544 2302 548
rect 2340 544 2372 548
rect 2372 544 2374 548
rect 2268 479 2302 504
rect 2340 479 2374 504
rect 2268 470 2270 479
rect 2270 470 2302 479
rect 2340 470 2372 479
rect 2372 470 2374 479
rect 2268 410 2302 430
rect 2340 410 2374 430
rect 2268 396 2270 410
rect 2270 396 2302 410
rect 2340 396 2372 410
rect 2372 396 2374 410
rect 2268 341 2302 356
rect 2340 341 2374 356
rect 2268 322 2270 341
rect 2270 322 2302 341
rect 2340 322 2372 341
rect 2372 322 2374 341
rect 2268 272 2302 282
rect 2340 272 2374 282
rect 2268 248 2270 272
rect 2270 248 2302 272
rect 2340 248 2372 272
rect 2372 248 2374 272
rect 2268 203 2302 208
rect 2340 203 2374 208
rect 2268 174 2270 203
rect 2270 174 2302 203
rect 2340 174 2372 203
rect 2372 174 2374 203
rect 2268 100 2270 134
rect 2270 100 2302 134
rect 2340 100 2372 134
rect 2372 100 2374 134
rect 2680 2966 2682 3000
rect 2682 2966 2714 3000
rect 2752 2966 2784 3000
rect 2784 2966 2786 3000
rect 2680 2893 2682 2927
rect 2682 2893 2714 2927
rect 2752 2893 2784 2927
rect 2784 2893 2786 2927
rect 2680 2820 2682 2854
rect 2682 2820 2714 2854
rect 2752 2820 2784 2854
rect 2784 2820 2786 2854
rect 2680 2747 2682 2781
rect 2682 2747 2714 2781
rect 2752 2747 2784 2781
rect 2784 2747 2786 2781
rect 2680 2674 2682 2708
rect 2682 2674 2714 2708
rect 2752 2674 2784 2708
rect 2784 2674 2786 2708
rect 2680 2601 2682 2635
rect 2682 2601 2714 2635
rect 2752 2601 2784 2635
rect 2784 2601 2786 2635
rect 2680 2528 2682 2562
rect 2682 2528 2714 2562
rect 2752 2528 2784 2562
rect 2784 2528 2786 2562
rect 2680 2455 2682 2489
rect 2682 2455 2714 2489
rect 2752 2455 2784 2489
rect 2784 2455 2786 2489
rect 2680 2382 2682 2416
rect 2682 2382 2714 2416
rect 2752 2382 2784 2416
rect 2784 2382 2786 2416
rect 2680 2309 2682 2343
rect 2682 2309 2714 2343
rect 2752 2309 2784 2343
rect 2784 2309 2786 2343
rect 2680 2236 2682 2270
rect 2682 2236 2714 2270
rect 2752 2236 2784 2270
rect 2784 2236 2786 2270
rect 2680 2163 2682 2197
rect 2682 2163 2714 2197
rect 2752 2163 2784 2197
rect 2784 2163 2786 2197
rect 2680 2090 2682 2124
rect 2682 2090 2714 2124
rect 2752 2090 2784 2124
rect 2784 2090 2786 2124
rect 2680 2017 2682 2051
rect 2682 2017 2714 2051
rect 2752 2017 2784 2051
rect 2784 2017 2786 2051
rect 2680 1944 2682 1978
rect 2682 1944 2714 1978
rect 2752 1944 2784 1978
rect 2784 1944 2786 1978
rect 2680 1871 2682 1905
rect 2682 1871 2714 1905
rect 2752 1871 2784 1905
rect 2784 1871 2786 1905
rect 2680 1798 2682 1832
rect 2682 1798 2714 1832
rect 2752 1798 2784 1832
rect 2784 1798 2786 1832
rect 2680 1725 2682 1759
rect 2682 1725 2714 1759
rect 2752 1725 2784 1759
rect 2784 1725 2786 1759
rect 2680 1652 2682 1686
rect 2682 1652 2714 1686
rect 2752 1652 2784 1686
rect 2784 1652 2786 1686
rect 2680 1579 2682 1613
rect 2682 1579 2714 1613
rect 2752 1579 2784 1613
rect 2784 1579 2786 1613
rect 2680 1506 2682 1540
rect 2682 1506 2714 1540
rect 2752 1506 2784 1540
rect 2784 1506 2786 1540
rect 2680 1432 2682 1466
rect 2682 1432 2714 1466
rect 2752 1432 2784 1466
rect 2784 1432 2786 1466
rect 2680 1358 2682 1392
rect 2682 1358 2714 1392
rect 2752 1358 2784 1392
rect 2784 1358 2786 1392
rect 2680 1284 2682 1318
rect 2682 1284 2714 1318
rect 2752 1284 2784 1318
rect 2784 1284 2786 1318
rect 2680 1210 2682 1244
rect 2682 1210 2714 1244
rect 2752 1210 2784 1244
rect 2784 1210 2786 1244
rect 2680 1136 2682 1170
rect 2682 1136 2714 1170
rect 2752 1136 2784 1170
rect 2784 1136 2786 1170
rect 2680 1062 2682 1096
rect 2682 1062 2714 1096
rect 2752 1062 2784 1096
rect 2784 1062 2786 1096
rect 2680 988 2682 1022
rect 2682 988 2714 1022
rect 2752 988 2784 1022
rect 2784 988 2786 1022
rect 2680 914 2682 948
rect 2682 914 2714 948
rect 2752 914 2784 948
rect 2784 914 2786 948
rect 2680 840 2682 874
rect 2682 840 2714 874
rect 2752 840 2784 874
rect 2784 840 2786 874
rect 2680 790 2682 800
rect 2682 790 2714 800
rect 2752 790 2784 800
rect 2784 790 2786 800
rect 2680 766 2714 790
rect 2752 766 2786 790
rect 2680 721 2682 726
rect 2682 721 2714 726
rect 2752 721 2784 726
rect 2784 721 2786 726
rect 2680 692 2714 721
rect 2752 692 2786 721
rect 2680 618 2714 652
rect 2752 618 2786 652
rect 2680 548 2714 578
rect 2752 548 2786 578
rect 2680 544 2682 548
rect 2682 544 2714 548
rect 2752 544 2784 548
rect 2784 544 2786 548
rect 2680 479 2714 504
rect 2752 479 2786 504
rect 2680 470 2682 479
rect 2682 470 2714 479
rect 2752 470 2784 479
rect 2784 470 2786 479
rect 2680 410 2714 430
rect 2752 410 2786 430
rect 2680 396 2682 410
rect 2682 396 2714 410
rect 2752 396 2784 410
rect 2784 396 2786 410
rect 2680 341 2714 356
rect 2752 341 2786 356
rect 2680 322 2682 341
rect 2682 322 2714 341
rect 2752 322 2784 341
rect 2784 322 2786 341
rect 2680 272 2714 282
rect 2752 272 2786 282
rect 2680 248 2682 272
rect 2682 248 2714 272
rect 2752 248 2784 272
rect 2784 248 2786 272
rect 2680 203 2714 208
rect 2752 203 2786 208
rect 2680 174 2682 203
rect 2682 174 2714 203
rect 2752 174 2784 203
rect 2784 174 2786 203
rect 2680 100 2682 134
rect 2682 100 2714 134
rect 2752 100 2784 134
rect 2784 100 2786 134
rect 3092 2966 3094 3000
rect 3094 2966 3126 3000
rect 3164 2966 3196 3000
rect 3196 2966 3198 3000
rect 3092 2893 3094 2927
rect 3094 2893 3126 2927
rect 3164 2893 3196 2927
rect 3196 2893 3198 2927
rect 3092 2820 3094 2854
rect 3094 2820 3126 2854
rect 3164 2820 3196 2854
rect 3196 2820 3198 2854
rect 3092 2747 3094 2781
rect 3094 2747 3126 2781
rect 3164 2747 3196 2781
rect 3196 2747 3198 2781
rect 3092 2674 3094 2708
rect 3094 2674 3126 2708
rect 3164 2674 3196 2708
rect 3196 2674 3198 2708
rect 3092 2601 3094 2635
rect 3094 2601 3126 2635
rect 3164 2601 3196 2635
rect 3196 2601 3198 2635
rect 3092 2528 3094 2562
rect 3094 2528 3126 2562
rect 3164 2528 3196 2562
rect 3196 2528 3198 2562
rect 3092 2455 3094 2489
rect 3094 2455 3126 2489
rect 3164 2455 3196 2489
rect 3196 2455 3198 2489
rect 3092 2382 3094 2416
rect 3094 2382 3126 2416
rect 3164 2382 3196 2416
rect 3196 2382 3198 2416
rect 3092 2309 3094 2343
rect 3094 2309 3126 2343
rect 3164 2309 3196 2343
rect 3196 2309 3198 2343
rect 3092 2236 3094 2270
rect 3094 2236 3126 2270
rect 3164 2236 3196 2270
rect 3196 2236 3198 2270
rect 3092 2163 3094 2197
rect 3094 2163 3126 2197
rect 3164 2163 3196 2197
rect 3196 2163 3198 2197
rect 3092 2090 3094 2124
rect 3094 2090 3126 2124
rect 3164 2090 3196 2124
rect 3196 2090 3198 2124
rect 3092 2017 3094 2051
rect 3094 2017 3126 2051
rect 3164 2017 3196 2051
rect 3196 2017 3198 2051
rect 3092 1944 3094 1978
rect 3094 1944 3126 1978
rect 3164 1944 3196 1978
rect 3196 1944 3198 1978
rect 3092 1871 3094 1905
rect 3094 1871 3126 1905
rect 3164 1871 3196 1905
rect 3196 1871 3198 1905
rect 3092 1798 3094 1832
rect 3094 1798 3126 1832
rect 3164 1798 3196 1832
rect 3196 1798 3198 1832
rect 3092 1725 3094 1759
rect 3094 1725 3126 1759
rect 3164 1725 3196 1759
rect 3196 1725 3198 1759
rect 3092 1652 3094 1686
rect 3094 1652 3126 1686
rect 3164 1652 3196 1686
rect 3196 1652 3198 1686
rect 3092 1579 3094 1613
rect 3094 1579 3126 1613
rect 3164 1579 3196 1613
rect 3196 1579 3198 1613
rect 3092 1506 3094 1540
rect 3094 1506 3126 1540
rect 3164 1506 3196 1540
rect 3196 1506 3198 1540
rect 3092 1432 3094 1466
rect 3094 1432 3126 1466
rect 3164 1432 3196 1466
rect 3196 1432 3198 1466
rect 3092 1358 3094 1392
rect 3094 1358 3126 1392
rect 3164 1358 3196 1392
rect 3196 1358 3198 1392
rect 3092 1284 3094 1318
rect 3094 1284 3126 1318
rect 3164 1284 3196 1318
rect 3196 1284 3198 1318
rect 3092 1210 3094 1244
rect 3094 1210 3126 1244
rect 3164 1210 3196 1244
rect 3196 1210 3198 1244
rect 3092 1136 3094 1170
rect 3094 1136 3126 1170
rect 3164 1136 3196 1170
rect 3196 1136 3198 1170
rect 3092 1062 3094 1096
rect 3094 1062 3126 1096
rect 3164 1062 3196 1096
rect 3196 1062 3198 1096
rect 3092 988 3094 1022
rect 3094 988 3126 1022
rect 3164 988 3196 1022
rect 3196 988 3198 1022
rect 3092 914 3094 948
rect 3094 914 3126 948
rect 3164 914 3196 948
rect 3196 914 3198 948
rect 3092 840 3094 874
rect 3094 840 3126 874
rect 3164 840 3196 874
rect 3196 840 3198 874
rect 3092 790 3094 800
rect 3094 790 3126 800
rect 3164 790 3196 800
rect 3196 790 3198 800
rect 3092 766 3126 790
rect 3164 766 3198 790
rect 3092 721 3094 726
rect 3094 721 3126 726
rect 3164 721 3196 726
rect 3196 721 3198 726
rect 3092 692 3126 721
rect 3164 692 3198 721
rect 3092 618 3126 652
rect 3164 618 3198 652
rect 3092 548 3126 578
rect 3164 548 3198 578
rect 3092 544 3094 548
rect 3094 544 3126 548
rect 3164 544 3196 548
rect 3196 544 3198 548
rect 3092 479 3126 504
rect 3164 479 3198 504
rect 3092 470 3094 479
rect 3094 470 3126 479
rect 3164 470 3196 479
rect 3196 470 3198 479
rect 3092 410 3126 430
rect 3164 410 3198 430
rect 3092 396 3094 410
rect 3094 396 3126 410
rect 3164 396 3196 410
rect 3196 396 3198 410
rect 3092 341 3126 356
rect 3164 341 3198 356
rect 3092 322 3094 341
rect 3094 322 3126 341
rect 3164 322 3196 341
rect 3196 322 3198 341
rect 3092 272 3126 282
rect 3164 272 3198 282
rect 3092 248 3094 272
rect 3094 248 3126 272
rect 3164 248 3196 272
rect 3196 248 3198 272
rect 3092 203 3126 208
rect 3164 203 3198 208
rect 3092 174 3094 203
rect 3094 174 3126 203
rect 3164 174 3196 203
rect 3196 174 3198 203
rect 3092 100 3094 134
rect 3094 100 3126 134
rect 3164 100 3196 134
rect 3196 100 3198 134
rect 3504 2966 3506 3000
rect 3506 2966 3538 3000
rect 3576 2966 3608 3000
rect 3608 2966 3610 3000
rect 3504 2893 3506 2927
rect 3506 2893 3538 2927
rect 3576 2893 3608 2927
rect 3608 2893 3610 2927
rect 3504 2820 3506 2854
rect 3506 2820 3538 2854
rect 3576 2820 3608 2854
rect 3608 2820 3610 2854
rect 3504 2747 3506 2781
rect 3506 2747 3538 2781
rect 3576 2747 3608 2781
rect 3608 2747 3610 2781
rect 3504 2674 3506 2708
rect 3506 2674 3538 2708
rect 3576 2674 3608 2708
rect 3608 2674 3610 2708
rect 3504 2601 3506 2635
rect 3506 2601 3538 2635
rect 3576 2601 3608 2635
rect 3608 2601 3610 2635
rect 3504 2528 3506 2562
rect 3506 2528 3538 2562
rect 3576 2528 3608 2562
rect 3608 2528 3610 2562
rect 3504 2455 3506 2489
rect 3506 2455 3538 2489
rect 3576 2455 3608 2489
rect 3608 2455 3610 2489
rect 3504 2382 3506 2416
rect 3506 2382 3538 2416
rect 3576 2382 3608 2416
rect 3608 2382 3610 2416
rect 3504 2309 3506 2343
rect 3506 2309 3538 2343
rect 3576 2309 3608 2343
rect 3608 2309 3610 2343
rect 3504 2236 3506 2270
rect 3506 2236 3538 2270
rect 3576 2236 3608 2270
rect 3608 2236 3610 2270
rect 3504 2163 3506 2197
rect 3506 2163 3538 2197
rect 3576 2163 3608 2197
rect 3608 2163 3610 2197
rect 3504 2090 3506 2124
rect 3506 2090 3538 2124
rect 3576 2090 3608 2124
rect 3608 2090 3610 2124
rect 3504 2017 3506 2051
rect 3506 2017 3538 2051
rect 3576 2017 3608 2051
rect 3608 2017 3610 2051
rect 3504 1944 3506 1978
rect 3506 1944 3538 1978
rect 3576 1944 3608 1978
rect 3608 1944 3610 1978
rect 3504 1871 3506 1905
rect 3506 1871 3538 1905
rect 3576 1871 3608 1905
rect 3608 1871 3610 1905
rect 3504 1798 3506 1832
rect 3506 1798 3538 1832
rect 3576 1798 3608 1832
rect 3608 1798 3610 1832
rect 3504 1725 3506 1759
rect 3506 1725 3538 1759
rect 3576 1725 3608 1759
rect 3608 1725 3610 1759
rect 3504 1652 3506 1686
rect 3506 1652 3538 1686
rect 3576 1652 3608 1686
rect 3608 1652 3610 1686
rect 3504 1579 3506 1613
rect 3506 1579 3538 1613
rect 3576 1579 3608 1613
rect 3608 1579 3610 1613
rect 3504 1506 3506 1540
rect 3506 1506 3538 1540
rect 3576 1506 3608 1540
rect 3608 1506 3610 1540
rect 3504 1432 3506 1466
rect 3506 1432 3538 1466
rect 3576 1432 3608 1466
rect 3608 1432 3610 1466
rect 3504 1358 3506 1392
rect 3506 1358 3538 1392
rect 3576 1358 3608 1392
rect 3608 1358 3610 1392
rect 3504 1284 3506 1318
rect 3506 1284 3538 1318
rect 3576 1284 3608 1318
rect 3608 1284 3610 1318
rect 3504 1210 3506 1244
rect 3506 1210 3538 1244
rect 3576 1210 3608 1244
rect 3608 1210 3610 1244
rect 3504 1136 3506 1170
rect 3506 1136 3538 1170
rect 3576 1136 3608 1170
rect 3608 1136 3610 1170
rect 3504 1062 3506 1096
rect 3506 1062 3538 1096
rect 3576 1062 3608 1096
rect 3608 1062 3610 1096
rect 3504 988 3506 1022
rect 3506 988 3538 1022
rect 3576 988 3608 1022
rect 3608 988 3610 1022
rect 3504 914 3506 948
rect 3506 914 3538 948
rect 3576 914 3608 948
rect 3608 914 3610 948
rect 3504 840 3506 874
rect 3506 840 3538 874
rect 3576 840 3608 874
rect 3608 840 3610 874
rect 3504 790 3506 800
rect 3506 790 3538 800
rect 3576 790 3608 800
rect 3608 790 3610 800
rect 3504 766 3538 790
rect 3576 766 3610 790
rect 3504 721 3506 726
rect 3506 721 3538 726
rect 3576 721 3608 726
rect 3608 721 3610 726
rect 3504 692 3538 721
rect 3576 692 3610 721
rect 3504 618 3538 652
rect 3576 618 3610 652
rect 3504 548 3538 578
rect 3576 548 3610 578
rect 3504 544 3506 548
rect 3506 544 3538 548
rect 3576 544 3608 548
rect 3608 544 3610 548
rect 3504 479 3538 504
rect 3576 479 3610 504
rect 3504 470 3506 479
rect 3506 470 3538 479
rect 3576 470 3608 479
rect 3608 470 3610 479
rect 3504 410 3538 430
rect 3576 410 3610 430
rect 3504 396 3506 410
rect 3506 396 3538 410
rect 3576 396 3608 410
rect 3608 396 3610 410
rect 3504 341 3538 356
rect 3576 341 3610 356
rect 3504 322 3506 341
rect 3506 322 3538 341
rect 3576 322 3608 341
rect 3608 322 3610 341
rect 3504 272 3538 282
rect 3576 272 3610 282
rect 3504 248 3506 272
rect 3506 248 3538 272
rect 3576 248 3608 272
rect 3608 248 3610 272
rect 3504 203 3538 208
rect 3576 203 3610 208
rect 3504 174 3506 203
rect 3506 174 3538 203
rect 3576 174 3608 203
rect 3608 174 3610 203
rect 3504 100 3506 134
rect 3506 100 3538 134
rect 3576 100 3608 134
rect 3608 100 3610 134
rect 3916 2966 3918 3000
rect 3918 2966 3950 3000
rect 3988 2966 4020 3000
rect 4020 2966 4022 3000
rect 3916 2893 3918 2927
rect 3918 2893 3950 2927
rect 3988 2893 4020 2927
rect 4020 2893 4022 2927
rect 3916 2820 3918 2854
rect 3918 2820 3950 2854
rect 3988 2820 4020 2854
rect 4020 2820 4022 2854
rect 3916 2747 3918 2781
rect 3918 2747 3950 2781
rect 3988 2747 4020 2781
rect 4020 2747 4022 2781
rect 3916 2674 3918 2708
rect 3918 2674 3950 2708
rect 3988 2674 4020 2708
rect 4020 2674 4022 2708
rect 3916 2601 3918 2635
rect 3918 2601 3950 2635
rect 3988 2601 4020 2635
rect 4020 2601 4022 2635
rect 3916 2528 3918 2562
rect 3918 2528 3950 2562
rect 3988 2528 4020 2562
rect 4020 2528 4022 2562
rect 3916 2455 3918 2489
rect 3918 2455 3950 2489
rect 3988 2455 4020 2489
rect 4020 2455 4022 2489
rect 3916 2382 3918 2416
rect 3918 2382 3950 2416
rect 3988 2382 4020 2416
rect 4020 2382 4022 2416
rect 3916 2309 3918 2343
rect 3918 2309 3950 2343
rect 3988 2309 4020 2343
rect 4020 2309 4022 2343
rect 3916 2236 3918 2270
rect 3918 2236 3950 2270
rect 3988 2236 4020 2270
rect 4020 2236 4022 2270
rect 3916 2163 3918 2197
rect 3918 2163 3950 2197
rect 3988 2163 4020 2197
rect 4020 2163 4022 2197
rect 3916 2090 3918 2124
rect 3918 2090 3950 2124
rect 3988 2090 4020 2124
rect 4020 2090 4022 2124
rect 3916 2017 3918 2051
rect 3918 2017 3950 2051
rect 3988 2017 4020 2051
rect 4020 2017 4022 2051
rect 3916 1944 3918 1978
rect 3918 1944 3950 1978
rect 3988 1944 4020 1978
rect 4020 1944 4022 1978
rect 3916 1871 3918 1905
rect 3918 1871 3950 1905
rect 3988 1871 4020 1905
rect 4020 1871 4022 1905
rect 3916 1798 3918 1832
rect 3918 1798 3950 1832
rect 3988 1798 4020 1832
rect 4020 1798 4022 1832
rect 3916 1725 3918 1759
rect 3918 1725 3950 1759
rect 3988 1725 4020 1759
rect 4020 1725 4022 1759
rect 3916 1652 3918 1686
rect 3918 1652 3950 1686
rect 3988 1652 4020 1686
rect 4020 1652 4022 1686
rect 3916 1579 3918 1613
rect 3918 1579 3950 1613
rect 3988 1579 4020 1613
rect 4020 1579 4022 1613
rect 3916 1506 3918 1540
rect 3918 1506 3950 1540
rect 3988 1506 4020 1540
rect 4020 1506 4022 1540
rect 3916 1432 3918 1466
rect 3918 1432 3950 1466
rect 3988 1432 4020 1466
rect 4020 1432 4022 1466
rect 3916 1358 3918 1392
rect 3918 1358 3950 1392
rect 3988 1358 4020 1392
rect 4020 1358 4022 1392
rect 3916 1284 3918 1318
rect 3918 1284 3950 1318
rect 3988 1284 4020 1318
rect 4020 1284 4022 1318
rect 3916 1210 3918 1244
rect 3918 1210 3950 1244
rect 3988 1210 4020 1244
rect 4020 1210 4022 1244
rect 3916 1136 3918 1170
rect 3918 1136 3950 1170
rect 3988 1136 4020 1170
rect 4020 1136 4022 1170
rect 3916 1062 3918 1096
rect 3918 1062 3950 1096
rect 3988 1062 4020 1096
rect 4020 1062 4022 1096
rect 3916 988 3918 1022
rect 3918 988 3950 1022
rect 3988 988 4020 1022
rect 4020 988 4022 1022
rect 3916 914 3918 948
rect 3918 914 3950 948
rect 3988 914 4020 948
rect 4020 914 4022 948
rect 3916 840 3918 874
rect 3918 840 3950 874
rect 3988 840 4020 874
rect 4020 840 4022 874
rect 3916 790 3918 800
rect 3918 790 3950 800
rect 3988 790 4020 800
rect 4020 790 4022 800
rect 3916 766 3950 790
rect 3988 766 4022 790
rect 3916 721 3918 726
rect 3918 721 3950 726
rect 3988 721 4020 726
rect 4020 721 4022 726
rect 3916 692 3950 721
rect 3988 692 4022 721
rect 3916 618 3950 652
rect 3988 618 4022 652
rect 3916 548 3950 578
rect 3988 548 4022 578
rect 3916 544 3918 548
rect 3918 544 3950 548
rect 3988 544 4020 548
rect 4020 544 4022 548
rect 3916 479 3950 504
rect 3988 479 4022 504
rect 3916 470 3918 479
rect 3918 470 3950 479
rect 3988 470 4020 479
rect 4020 470 4022 479
rect 3916 410 3950 430
rect 3988 410 4022 430
rect 3916 396 3918 410
rect 3918 396 3950 410
rect 3988 396 4020 410
rect 4020 396 4022 410
rect 3916 341 3950 356
rect 3988 341 4022 356
rect 3916 322 3918 341
rect 3918 322 3950 341
rect 3988 322 4020 341
rect 4020 322 4022 341
rect 3916 272 3950 282
rect 3988 272 4022 282
rect 3916 248 3918 272
rect 3918 248 3950 272
rect 3988 248 4020 272
rect 4020 248 4022 272
rect 3916 203 3950 208
rect 3988 203 4022 208
rect 3916 174 3918 203
rect 3918 174 3950 203
rect 3988 174 4020 203
rect 4020 174 4022 203
rect 3916 100 3918 134
rect 3918 100 3950 134
rect 3988 100 4020 134
rect 4020 100 4022 134
rect 4328 2966 4330 3000
rect 4330 2966 4362 3000
rect 4400 2966 4432 3000
rect 4432 2966 4434 3000
rect 4328 2893 4330 2927
rect 4330 2893 4362 2927
rect 4400 2893 4432 2927
rect 4432 2893 4434 2927
rect 4328 2820 4330 2854
rect 4330 2820 4362 2854
rect 4400 2820 4432 2854
rect 4432 2820 4434 2854
rect 4328 2747 4330 2781
rect 4330 2747 4362 2781
rect 4400 2747 4432 2781
rect 4432 2747 4434 2781
rect 4328 2674 4330 2708
rect 4330 2674 4362 2708
rect 4400 2674 4432 2708
rect 4432 2674 4434 2708
rect 4328 2601 4330 2635
rect 4330 2601 4362 2635
rect 4400 2601 4432 2635
rect 4432 2601 4434 2635
rect 4328 2528 4330 2562
rect 4330 2528 4362 2562
rect 4400 2528 4432 2562
rect 4432 2528 4434 2562
rect 4328 2455 4330 2489
rect 4330 2455 4362 2489
rect 4400 2455 4432 2489
rect 4432 2455 4434 2489
rect 4328 2382 4330 2416
rect 4330 2382 4362 2416
rect 4400 2382 4432 2416
rect 4432 2382 4434 2416
rect 4328 2309 4330 2343
rect 4330 2309 4362 2343
rect 4400 2309 4432 2343
rect 4432 2309 4434 2343
rect 4328 2236 4330 2270
rect 4330 2236 4362 2270
rect 4400 2236 4432 2270
rect 4432 2236 4434 2270
rect 4328 2163 4330 2197
rect 4330 2163 4362 2197
rect 4400 2163 4432 2197
rect 4432 2163 4434 2197
rect 4328 2090 4330 2124
rect 4330 2090 4362 2124
rect 4400 2090 4432 2124
rect 4432 2090 4434 2124
rect 4328 2017 4330 2051
rect 4330 2017 4362 2051
rect 4400 2017 4432 2051
rect 4432 2017 4434 2051
rect 4328 1944 4330 1978
rect 4330 1944 4362 1978
rect 4400 1944 4432 1978
rect 4432 1944 4434 1978
rect 4328 1871 4330 1905
rect 4330 1871 4362 1905
rect 4400 1871 4432 1905
rect 4432 1871 4434 1905
rect 4328 1798 4330 1832
rect 4330 1798 4362 1832
rect 4400 1798 4432 1832
rect 4432 1798 4434 1832
rect 4328 1725 4330 1759
rect 4330 1725 4362 1759
rect 4400 1725 4432 1759
rect 4432 1725 4434 1759
rect 4328 1652 4330 1686
rect 4330 1652 4362 1686
rect 4400 1652 4432 1686
rect 4432 1652 4434 1686
rect 4328 1579 4330 1613
rect 4330 1579 4362 1613
rect 4400 1579 4432 1613
rect 4432 1579 4434 1613
rect 4328 1506 4330 1540
rect 4330 1506 4362 1540
rect 4400 1506 4432 1540
rect 4432 1506 4434 1540
rect 4328 1432 4330 1466
rect 4330 1432 4362 1466
rect 4400 1432 4432 1466
rect 4432 1432 4434 1466
rect 4328 1358 4330 1392
rect 4330 1358 4362 1392
rect 4400 1358 4432 1392
rect 4432 1358 4434 1392
rect 4328 1284 4330 1318
rect 4330 1284 4362 1318
rect 4400 1284 4432 1318
rect 4432 1284 4434 1318
rect 4328 1210 4330 1244
rect 4330 1210 4362 1244
rect 4400 1210 4432 1244
rect 4432 1210 4434 1244
rect 4328 1136 4330 1170
rect 4330 1136 4362 1170
rect 4400 1136 4432 1170
rect 4432 1136 4434 1170
rect 4328 1062 4330 1096
rect 4330 1062 4362 1096
rect 4400 1062 4432 1096
rect 4432 1062 4434 1096
rect 4328 988 4330 1022
rect 4330 988 4362 1022
rect 4400 988 4432 1022
rect 4432 988 4434 1022
rect 4328 914 4330 948
rect 4330 914 4362 948
rect 4400 914 4432 948
rect 4432 914 4434 948
rect 4328 840 4330 874
rect 4330 840 4362 874
rect 4400 840 4432 874
rect 4432 840 4434 874
rect 4328 790 4330 800
rect 4330 790 4362 800
rect 4400 790 4432 800
rect 4432 790 4434 800
rect 4328 766 4362 790
rect 4400 766 4434 790
rect 4328 721 4330 726
rect 4330 721 4362 726
rect 4400 721 4432 726
rect 4432 721 4434 726
rect 4328 692 4362 721
rect 4400 692 4434 721
rect 4328 618 4362 652
rect 4400 618 4434 652
rect 4328 548 4362 578
rect 4400 548 4434 578
rect 4328 544 4330 548
rect 4330 544 4362 548
rect 4400 544 4432 548
rect 4432 544 4434 548
rect 4328 479 4362 504
rect 4400 479 4434 504
rect 4328 470 4330 479
rect 4330 470 4362 479
rect 4400 470 4432 479
rect 4432 470 4434 479
rect 4328 410 4362 430
rect 4400 410 4434 430
rect 4328 396 4330 410
rect 4330 396 4362 410
rect 4400 396 4432 410
rect 4432 396 4434 410
rect 4328 341 4362 356
rect 4400 341 4434 356
rect 4328 322 4330 341
rect 4330 322 4362 341
rect 4400 322 4432 341
rect 4432 322 4434 341
rect 4328 272 4362 282
rect 4400 272 4434 282
rect 4328 248 4330 272
rect 4330 248 4362 272
rect 4400 248 4432 272
rect 4432 248 4434 272
rect 4328 203 4362 208
rect 4400 203 4434 208
rect 4328 174 4330 203
rect 4330 174 4362 203
rect 4400 174 4432 203
rect 4432 174 4434 203
rect 4328 100 4330 134
rect 4330 100 4362 134
rect 4400 100 4432 134
rect 4432 100 4434 134
rect 4740 2966 4742 3000
rect 4742 2966 4774 3000
rect 4812 2966 4844 3000
rect 4844 2966 4846 3000
rect 4740 2893 4742 2927
rect 4742 2893 4774 2927
rect 4812 2893 4844 2927
rect 4844 2893 4846 2927
rect 4740 2820 4742 2854
rect 4742 2820 4774 2854
rect 4812 2820 4844 2854
rect 4844 2820 4846 2854
rect 4740 2747 4742 2781
rect 4742 2747 4774 2781
rect 4812 2747 4844 2781
rect 4844 2747 4846 2781
rect 4740 2674 4742 2708
rect 4742 2674 4774 2708
rect 4812 2674 4844 2708
rect 4844 2674 4846 2708
rect 4740 2601 4742 2635
rect 4742 2601 4774 2635
rect 4812 2601 4844 2635
rect 4844 2601 4846 2635
rect 4740 2528 4742 2562
rect 4742 2528 4774 2562
rect 4812 2528 4844 2562
rect 4844 2528 4846 2562
rect 4740 2455 4742 2489
rect 4742 2455 4774 2489
rect 4812 2455 4844 2489
rect 4844 2455 4846 2489
rect 4740 2382 4742 2416
rect 4742 2382 4774 2416
rect 4812 2382 4844 2416
rect 4844 2382 4846 2416
rect 4740 2309 4742 2343
rect 4742 2309 4774 2343
rect 4812 2309 4844 2343
rect 4844 2309 4846 2343
rect 4740 2236 4742 2270
rect 4742 2236 4774 2270
rect 4812 2236 4844 2270
rect 4844 2236 4846 2270
rect 4740 2163 4742 2197
rect 4742 2163 4774 2197
rect 4812 2163 4844 2197
rect 4844 2163 4846 2197
rect 4740 2090 4742 2124
rect 4742 2090 4774 2124
rect 4812 2090 4844 2124
rect 4844 2090 4846 2124
rect 4740 2017 4742 2051
rect 4742 2017 4774 2051
rect 4812 2017 4844 2051
rect 4844 2017 4846 2051
rect 4740 1944 4742 1978
rect 4742 1944 4774 1978
rect 4812 1944 4844 1978
rect 4844 1944 4846 1978
rect 4740 1871 4742 1905
rect 4742 1871 4774 1905
rect 4812 1871 4844 1905
rect 4844 1871 4846 1905
rect 4740 1798 4742 1832
rect 4742 1798 4774 1832
rect 4812 1798 4844 1832
rect 4844 1798 4846 1832
rect 4740 1725 4742 1759
rect 4742 1725 4774 1759
rect 4812 1725 4844 1759
rect 4844 1725 4846 1759
rect 4740 1652 4742 1686
rect 4742 1652 4774 1686
rect 4812 1652 4844 1686
rect 4844 1652 4846 1686
rect 4740 1579 4742 1613
rect 4742 1579 4774 1613
rect 4812 1579 4844 1613
rect 4844 1579 4846 1613
rect 4740 1506 4742 1540
rect 4742 1506 4774 1540
rect 4812 1506 4844 1540
rect 4844 1506 4846 1540
rect 4740 1432 4742 1466
rect 4742 1432 4774 1466
rect 4812 1432 4844 1466
rect 4844 1432 4846 1466
rect 4740 1358 4742 1392
rect 4742 1358 4774 1392
rect 4812 1358 4844 1392
rect 4844 1358 4846 1392
rect 4740 1284 4742 1318
rect 4742 1284 4774 1318
rect 4812 1284 4844 1318
rect 4844 1284 4846 1318
rect 4740 1210 4742 1244
rect 4742 1210 4774 1244
rect 4812 1210 4844 1244
rect 4844 1210 4846 1244
rect 4740 1136 4742 1170
rect 4742 1136 4774 1170
rect 4812 1136 4844 1170
rect 4844 1136 4846 1170
rect 4740 1062 4742 1096
rect 4742 1062 4774 1096
rect 4812 1062 4844 1096
rect 4844 1062 4846 1096
rect 4740 988 4742 1022
rect 4742 988 4774 1022
rect 4812 988 4844 1022
rect 4844 988 4846 1022
rect 4740 914 4742 948
rect 4742 914 4774 948
rect 4812 914 4844 948
rect 4844 914 4846 948
rect 4740 840 4742 874
rect 4742 840 4774 874
rect 4812 840 4844 874
rect 4844 840 4846 874
rect 4740 790 4742 800
rect 4742 790 4774 800
rect 4812 790 4844 800
rect 4844 790 4846 800
rect 4740 766 4774 790
rect 4812 766 4846 790
rect 4740 721 4742 726
rect 4742 721 4774 726
rect 4812 721 4844 726
rect 4844 721 4846 726
rect 4740 692 4774 721
rect 4812 692 4846 721
rect 4740 618 4774 652
rect 4812 618 4846 652
rect 4740 548 4774 578
rect 4812 548 4846 578
rect 4740 544 4742 548
rect 4742 544 4774 548
rect 4812 544 4844 548
rect 4844 544 4846 548
rect 4740 479 4774 504
rect 4812 479 4846 504
rect 4740 470 4742 479
rect 4742 470 4774 479
rect 4812 470 4844 479
rect 4844 470 4846 479
rect 4740 410 4774 430
rect 4812 410 4846 430
rect 4740 396 4742 410
rect 4742 396 4774 410
rect 4812 396 4844 410
rect 4844 396 4846 410
rect 4740 341 4774 356
rect 4812 341 4846 356
rect 4740 322 4742 341
rect 4742 322 4774 341
rect 4812 322 4844 341
rect 4844 322 4846 341
rect 4740 272 4774 282
rect 4812 272 4846 282
rect 4740 248 4742 272
rect 4742 248 4774 272
rect 4812 248 4844 272
rect 4844 248 4846 272
rect 4740 203 4774 208
rect 4812 203 4846 208
rect 4740 174 4742 203
rect 4742 174 4774 203
rect 4812 174 4844 203
rect 4844 174 4846 203
rect 4740 100 4742 134
rect 4742 100 4774 134
rect 4812 100 4844 134
rect 4844 100 4846 134
rect 5152 2966 5154 3000
rect 5154 2966 5186 3000
rect 5224 2966 5256 3000
rect 5256 2966 5258 3000
rect 5152 2893 5154 2927
rect 5154 2893 5186 2927
rect 5224 2893 5256 2927
rect 5256 2893 5258 2927
rect 5152 2820 5154 2854
rect 5154 2820 5186 2854
rect 5224 2820 5256 2854
rect 5256 2820 5258 2854
rect 5152 2747 5154 2781
rect 5154 2747 5186 2781
rect 5224 2747 5256 2781
rect 5256 2747 5258 2781
rect 5152 2674 5154 2708
rect 5154 2674 5186 2708
rect 5224 2674 5256 2708
rect 5256 2674 5258 2708
rect 5152 2601 5154 2635
rect 5154 2601 5186 2635
rect 5224 2601 5256 2635
rect 5256 2601 5258 2635
rect 5152 2528 5154 2562
rect 5154 2528 5186 2562
rect 5224 2528 5256 2562
rect 5256 2528 5258 2562
rect 5152 2455 5154 2489
rect 5154 2455 5186 2489
rect 5224 2455 5256 2489
rect 5256 2455 5258 2489
rect 5152 2382 5154 2416
rect 5154 2382 5186 2416
rect 5224 2382 5256 2416
rect 5256 2382 5258 2416
rect 5152 2309 5154 2343
rect 5154 2309 5186 2343
rect 5224 2309 5256 2343
rect 5256 2309 5258 2343
rect 5152 2236 5154 2270
rect 5154 2236 5186 2270
rect 5224 2236 5256 2270
rect 5256 2236 5258 2270
rect 5152 2163 5154 2197
rect 5154 2163 5186 2197
rect 5224 2163 5256 2197
rect 5256 2163 5258 2197
rect 5152 2090 5154 2124
rect 5154 2090 5186 2124
rect 5224 2090 5256 2124
rect 5256 2090 5258 2124
rect 5152 2017 5154 2051
rect 5154 2017 5186 2051
rect 5224 2017 5256 2051
rect 5256 2017 5258 2051
rect 5152 1944 5154 1978
rect 5154 1944 5186 1978
rect 5224 1944 5256 1978
rect 5256 1944 5258 1978
rect 5152 1871 5154 1905
rect 5154 1871 5186 1905
rect 5224 1871 5256 1905
rect 5256 1871 5258 1905
rect 5152 1798 5154 1832
rect 5154 1798 5186 1832
rect 5224 1798 5256 1832
rect 5256 1798 5258 1832
rect 5152 1725 5154 1759
rect 5154 1725 5186 1759
rect 5224 1725 5256 1759
rect 5256 1725 5258 1759
rect 5152 1652 5154 1686
rect 5154 1652 5186 1686
rect 5224 1652 5256 1686
rect 5256 1652 5258 1686
rect 5152 1579 5154 1613
rect 5154 1579 5186 1613
rect 5224 1579 5256 1613
rect 5256 1579 5258 1613
rect 5152 1506 5154 1540
rect 5154 1506 5186 1540
rect 5224 1506 5256 1540
rect 5256 1506 5258 1540
rect 5152 1432 5154 1466
rect 5154 1432 5186 1466
rect 5224 1432 5256 1466
rect 5256 1432 5258 1466
rect 5152 1358 5154 1392
rect 5154 1358 5186 1392
rect 5224 1358 5256 1392
rect 5256 1358 5258 1392
rect 5152 1284 5154 1318
rect 5154 1284 5186 1318
rect 5224 1284 5256 1318
rect 5256 1284 5258 1318
rect 5152 1210 5154 1244
rect 5154 1210 5186 1244
rect 5224 1210 5256 1244
rect 5256 1210 5258 1244
rect 5152 1136 5154 1170
rect 5154 1136 5186 1170
rect 5224 1136 5256 1170
rect 5256 1136 5258 1170
rect 5152 1062 5154 1096
rect 5154 1062 5186 1096
rect 5224 1062 5256 1096
rect 5256 1062 5258 1096
rect 5152 988 5154 1022
rect 5154 988 5186 1022
rect 5224 988 5256 1022
rect 5256 988 5258 1022
rect 5152 914 5154 948
rect 5154 914 5186 948
rect 5224 914 5256 948
rect 5256 914 5258 948
rect 5152 840 5154 874
rect 5154 840 5186 874
rect 5224 840 5256 874
rect 5256 840 5258 874
rect 5152 790 5154 800
rect 5154 790 5186 800
rect 5224 790 5256 800
rect 5256 790 5258 800
rect 5152 766 5186 790
rect 5224 766 5258 790
rect 5152 721 5154 726
rect 5154 721 5186 726
rect 5224 721 5256 726
rect 5256 721 5258 726
rect 5152 692 5186 721
rect 5224 692 5258 721
rect 5152 618 5186 652
rect 5224 618 5258 652
rect 5152 548 5186 578
rect 5224 548 5258 578
rect 5152 544 5154 548
rect 5154 544 5186 548
rect 5224 544 5256 548
rect 5256 544 5258 548
rect 5152 479 5186 504
rect 5224 479 5258 504
rect 5152 470 5154 479
rect 5154 470 5186 479
rect 5224 470 5256 479
rect 5256 470 5258 479
rect 5152 410 5186 430
rect 5224 410 5258 430
rect 5152 396 5154 410
rect 5154 396 5186 410
rect 5224 396 5256 410
rect 5256 396 5258 410
rect 5152 341 5186 356
rect 5224 341 5258 356
rect 5152 322 5154 341
rect 5154 322 5186 341
rect 5224 322 5256 341
rect 5256 322 5258 341
rect 5152 272 5186 282
rect 5224 272 5258 282
rect 5152 248 5154 272
rect 5154 248 5186 272
rect 5224 248 5256 272
rect 5256 248 5258 272
rect 5152 203 5186 208
rect 5224 203 5258 208
rect 5152 174 5154 203
rect 5154 174 5186 203
rect 5224 174 5256 203
rect 5256 174 5258 203
rect 5152 100 5154 134
rect 5154 100 5186 134
rect 5224 100 5256 134
rect 5256 100 5258 134
rect 5564 2966 5566 3000
rect 5566 2966 5598 3000
rect 5636 2966 5668 3000
rect 5668 2966 5670 3000
rect 5564 2893 5566 2927
rect 5566 2893 5598 2927
rect 5636 2893 5668 2927
rect 5668 2893 5670 2927
rect 5564 2820 5566 2854
rect 5566 2820 5598 2854
rect 5636 2820 5668 2854
rect 5668 2820 5670 2854
rect 5564 2747 5566 2781
rect 5566 2747 5598 2781
rect 5636 2747 5668 2781
rect 5668 2747 5670 2781
rect 5564 2674 5566 2708
rect 5566 2674 5598 2708
rect 5636 2674 5668 2708
rect 5668 2674 5670 2708
rect 5564 2601 5566 2635
rect 5566 2601 5598 2635
rect 5636 2601 5668 2635
rect 5668 2601 5670 2635
rect 5564 2528 5566 2562
rect 5566 2528 5598 2562
rect 5636 2528 5668 2562
rect 5668 2528 5670 2562
rect 5564 2455 5566 2489
rect 5566 2455 5598 2489
rect 5636 2455 5668 2489
rect 5668 2455 5670 2489
rect 5564 2382 5566 2416
rect 5566 2382 5598 2416
rect 5636 2382 5668 2416
rect 5668 2382 5670 2416
rect 5564 2309 5566 2343
rect 5566 2309 5598 2343
rect 5636 2309 5668 2343
rect 5668 2309 5670 2343
rect 5564 2236 5566 2270
rect 5566 2236 5598 2270
rect 5636 2236 5668 2270
rect 5668 2236 5670 2270
rect 5564 2163 5566 2197
rect 5566 2163 5598 2197
rect 5636 2163 5668 2197
rect 5668 2163 5670 2197
rect 5564 2090 5566 2124
rect 5566 2090 5598 2124
rect 5636 2090 5668 2124
rect 5668 2090 5670 2124
rect 5564 2017 5566 2051
rect 5566 2017 5598 2051
rect 5636 2017 5668 2051
rect 5668 2017 5670 2051
rect 5564 1944 5566 1978
rect 5566 1944 5598 1978
rect 5636 1944 5668 1978
rect 5668 1944 5670 1978
rect 5564 1871 5566 1905
rect 5566 1871 5598 1905
rect 5636 1871 5668 1905
rect 5668 1871 5670 1905
rect 5564 1798 5566 1832
rect 5566 1798 5598 1832
rect 5636 1798 5668 1832
rect 5668 1798 5670 1832
rect 5564 1725 5566 1759
rect 5566 1725 5598 1759
rect 5636 1725 5668 1759
rect 5668 1725 5670 1759
rect 5564 1652 5566 1686
rect 5566 1652 5598 1686
rect 5636 1652 5668 1686
rect 5668 1652 5670 1686
rect 5564 1579 5566 1613
rect 5566 1579 5598 1613
rect 5636 1579 5668 1613
rect 5668 1579 5670 1613
rect 5564 1506 5566 1540
rect 5566 1506 5598 1540
rect 5636 1506 5668 1540
rect 5668 1506 5670 1540
rect 5564 1432 5566 1466
rect 5566 1432 5598 1466
rect 5636 1432 5668 1466
rect 5668 1432 5670 1466
rect 5564 1358 5566 1392
rect 5566 1358 5598 1392
rect 5636 1358 5668 1392
rect 5668 1358 5670 1392
rect 5564 1284 5566 1318
rect 5566 1284 5598 1318
rect 5636 1284 5668 1318
rect 5668 1284 5670 1318
rect 5564 1210 5566 1244
rect 5566 1210 5598 1244
rect 5636 1210 5668 1244
rect 5668 1210 5670 1244
rect 5564 1136 5566 1170
rect 5566 1136 5598 1170
rect 5636 1136 5668 1170
rect 5668 1136 5670 1170
rect 5564 1062 5566 1096
rect 5566 1062 5598 1096
rect 5636 1062 5668 1096
rect 5668 1062 5670 1096
rect 5564 988 5566 1022
rect 5566 988 5598 1022
rect 5636 988 5668 1022
rect 5668 988 5670 1022
rect 5564 914 5566 948
rect 5566 914 5598 948
rect 5636 914 5668 948
rect 5668 914 5670 948
rect 5564 840 5566 874
rect 5566 840 5598 874
rect 5636 840 5668 874
rect 5668 840 5670 874
rect 5564 790 5566 800
rect 5566 790 5598 800
rect 5636 790 5668 800
rect 5668 790 5670 800
rect 5564 766 5598 790
rect 5636 766 5670 790
rect 5564 721 5566 726
rect 5566 721 5598 726
rect 5636 721 5668 726
rect 5668 721 5670 726
rect 5564 692 5598 721
rect 5636 692 5670 721
rect 5564 618 5598 652
rect 5636 618 5670 652
rect 5564 548 5598 578
rect 5636 548 5670 578
rect 5564 544 5566 548
rect 5566 544 5598 548
rect 5636 544 5668 548
rect 5668 544 5670 548
rect 5564 479 5598 504
rect 5636 479 5670 504
rect 5564 470 5566 479
rect 5566 470 5598 479
rect 5636 470 5668 479
rect 5668 470 5670 479
rect 5564 410 5598 430
rect 5636 410 5670 430
rect 5564 396 5566 410
rect 5566 396 5598 410
rect 5636 396 5668 410
rect 5668 396 5670 410
rect 5564 341 5598 356
rect 5636 341 5670 356
rect 5564 322 5566 341
rect 5566 322 5598 341
rect 5636 322 5668 341
rect 5668 322 5670 341
rect 5564 272 5598 282
rect 5636 272 5670 282
rect 5564 248 5566 272
rect 5566 248 5598 272
rect 5636 248 5668 272
rect 5668 248 5670 272
rect 5564 203 5598 208
rect 5636 203 5670 208
rect 5564 174 5566 203
rect 5566 174 5598 203
rect 5636 174 5668 203
rect 5668 174 5670 203
rect 5564 100 5566 134
rect 5566 100 5598 134
rect 5636 100 5668 134
rect 5668 100 5670 134
rect 5976 2966 5978 3000
rect 5978 2966 6010 3000
rect 6048 2966 6080 3000
rect 6080 2966 6082 3000
rect 5976 2893 5978 2927
rect 5978 2893 6010 2927
rect 6048 2893 6080 2927
rect 6080 2893 6082 2927
rect 5976 2820 5978 2854
rect 5978 2820 6010 2854
rect 6048 2820 6080 2854
rect 6080 2820 6082 2854
rect 5976 2747 5978 2781
rect 5978 2747 6010 2781
rect 6048 2747 6080 2781
rect 6080 2747 6082 2781
rect 5976 2674 5978 2708
rect 5978 2674 6010 2708
rect 6048 2674 6080 2708
rect 6080 2674 6082 2708
rect 5976 2601 5978 2635
rect 5978 2601 6010 2635
rect 6048 2601 6080 2635
rect 6080 2601 6082 2635
rect 5976 2528 5978 2562
rect 5978 2528 6010 2562
rect 6048 2528 6080 2562
rect 6080 2528 6082 2562
rect 5976 2455 5978 2489
rect 5978 2455 6010 2489
rect 6048 2455 6080 2489
rect 6080 2455 6082 2489
rect 5976 2382 5978 2416
rect 5978 2382 6010 2416
rect 6048 2382 6080 2416
rect 6080 2382 6082 2416
rect 5976 2309 5978 2343
rect 5978 2309 6010 2343
rect 6048 2309 6080 2343
rect 6080 2309 6082 2343
rect 5976 2236 5978 2270
rect 5978 2236 6010 2270
rect 6048 2236 6080 2270
rect 6080 2236 6082 2270
rect 5976 2163 5978 2197
rect 5978 2163 6010 2197
rect 6048 2163 6080 2197
rect 6080 2163 6082 2197
rect 5976 2090 5978 2124
rect 5978 2090 6010 2124
rect 6048 2090 6080 2124
rect 6080 2090 6082 2124
rect 5976 2017 5978 2051
rect 5978 2017 6010 2051
rect 6048 2017 6080 2051
rect 6080 2017 6082 2051
rect 5976 1944 5978 1978
rect 5978 1944 6010 1978
rect 6048 1944 6080 1978
rect 6080 1944 6082 1978
rect 5976 1871 5978 1905
rect 5978 1871 6010 1905
rect 6048 1871 6080 1905
rect 6080 1871 6082 1905
rect 5976 1798 5978 1832
rect 5978 1798 6010 1832
rect 6048 1798 6080 1832
rect 6080 1798 6082 1832
rect 5976 1725 5978 1759
rect 5978 1725 6010 1759
rect 6048 1725 6080 1759
rect 6080 1725 6082 1759
rect 5976 1652 5978 1686
rect 5978 1652 6010 1686
rect 6048 1652 6080 1686
rect 6080 1652 6082 1686
rect 5976 1579 5978 1613
rect 5978 1579 6010 1613
rect 6048 1579 6080 1613
rect 6080 1579 6082 1613
rect 5976 1506 5978 1540
rect 5978 1506 6010 1540
rect 6048 1506 6080 1540
rect 6080 1506 6082 1540
rect 5976 1432 5978 1466
rect 5978 1432 6010 1466
rect 6048 1432 6080 1466
rect 6080 1432 6082 1466
rect 5976 1358 5978 1392
rect 5978 1358 6010 1392
rect 6048 1358 6080 1392
rect 6080 1358 6082 1392
rect 5976 1284 5978 1318
rect 5978 1284 6010 1318
rect 6048 1284 6080 1318
rect 6080 1284 6082 1318
rect 5976 1210 5978 1244
rect 5978 1210 6010 1244
rect 6048 1210 6080 1244
rect 6080 1210 6082 1244
rect 5976 1136 5978 1170
rect 5978 1136 6010 1170
rect 6048 1136 6080 1170
rect 6080 1136 6082 1170
rect 5976 1062 5978 1096
rect 5978 1062 6010 1096
rect 6048 1062 6080 1096
rect 6080 1062 6082 1096
rect 5976 988 5978 1022
rect 5978 988 6010 1022
rect 6048 988 6080 1022
rect 6080 988 6082 1022
rect 5976 914 5978 948
rect 5978 914 6010 948
rect 6048 914 6080 948
rect 6080 914 6082 948
rect 5976 840 5978 874
rect 5978 840 6010 874
rect 6048 840 6080 874
rect 6080 840 6082 874
rect 5976 790 5978 800
rect 5978 790 6010 800
rect 6048 790 6080 800
rect 6080 790 6082 800
rect 5976 766 6010 790
rect 6048 766 6082 790
rect 5976 721 5978 726
rect 5978 721 6010 726
rect 6048 721 6080 726
rect 6080 721 6082 726
rect 5976 692 6010 721
rect 6048 692 6082 721
rect 5976 618 6010 652
rect 6048 618 6082 652
rect 5976 548 6010 578
rect 6048 548 6082 578
rect 5976 544 5978 548
rect 5978 544 6010 548
rect 6048 544 6080 548
rect 6080 544 6082 548
rect 5976 479 6010 504
rect 6048 479 6082 504
rect 5976 470 5978 479
rect 5978 470 6010 479
rect 6048 470 6080 479
rect 6080 470 6082 479
rect 5976 410 6010 430
rect 6048 410 6082 430
rect 5976 396 5978 410
rect 5978 396 6010 410
rect 6048 396 6080 410
rect 6080 396 6082 410
rect 5976 341 6010 356
rect 6048 341 6082 356
rect 5976 322 5978 341
rect 5978 322 6010 341
rect 6048 322 6080 341
rect 6080 322 6082 341
rect 5976 272 6010 282
rect 6048 272 6082 282
rect 5976 248 5978 272
rect 5978 248 6010 272
rect 6048 248 6080 272
rect 6080 248 6082 272
rect 5976 203 6010 208
rect 6048 203 6082 208
rect 5976 174 5978 203
rect 5978 174 6010 203
rect 6048 174 6080 203
rect 6080 174 6082 203
rect 5976 100 5978 134
rect 5978 100 6010 134
rect 6048 100 6080 134
rect 6080 100 6082 134
rect 6388 2966 6390 3000
rect 6390 2966 6422 3000
rect 6460 2966 6492 3000
rect 6492 2966 6494 3000
rect 6388 2893 6390 2927
rect 6390 2893 6422 2927
rect 6460 2893 6492 2927
rect 6492 2893 6494 2927
rect 6388 2820 6390 2854
rect 6390 2820 6422 2854
rect 6460 2820 6492 2854
rect 6492 2820 6494 2854
rect 6388 2747 6390 2781
rect 6390 2747 6422 2781
rect 6460 2747 6492 2781
rect 6492 2747 6494 2781
rect 6388 2674 6390 2708
rect 6390 2674 6422 2708
rect 6460 2674 6492 2708
rect 6492 2674 6494 2708
rect 6388 2601 6390 2635
rect 6390 2601 6422 2635
rect 6460 2601 6492 2635
rect 6492 2601 6494 2635
rect 6388 2528 6390 2562
rect 6390 2528 6422 2562
rect 6460 2528 6492 2562
rect 6492 2528 6494 2562
rect 6388 2455 6390 2489
rect 6390 2455 6422 2489
rect 6460 2455 6492 2489
rect 6492 2455 6494 2489
rect 6388 2382 6390 2416
rect 6390 2382 6422 2416
rect 6460 2382 6492 2416
rect 6492 2382 6494 2416
rect 6388 2309 6390 2343
rect 6390 2309 6422 2343
rect 6460 2309 6492 2343
rect 6492 2309 6494 2343
rect 6388 2236 6390 2270
rect 6390 2236 6422 2270
rect 6460 2236 6492 2270
rect 6492 2236 6494 2270
rect 6388 2163 6390 2197
rect 6390 2163 6422 2197
rect 6460 2163 6492 2197
rect 6492 2163 6494 2197
rect 6388 2090 6390 2124
rect 6390 2090 6422 2124
rect 6460 2090 6492 2124
rect 6492 2090 6494 2124
rect 6388 2017 6390 2051
rect 6390 2017 6422 2051
rect 6460 2017 6492 2051
rect 6492 2017 6494 2051
rect 6388 1944 6390 1978
rect 6390 1944 6422 1978
rect 6460 1944 6492 1978
rect 6492 1944 6494 1978
rect 6388 1871 6390 1905
rect 6390 1871 6422 1905
rect 6460 1871 6492 1905
rect 6492 1871 6494 1905
rect 6388 1798 6390 1832
rect 6390 1798 6422 1832
rect 6460 1798 6492 1832
rect 6492 1798 6494 1832
rect 6388 1725 6390 1759
rect 6390 1725 6422 1759
rect 6460 1725 6492 1759
rect 6492 1725 6494 1759
rect 6388 1652 6390 1686
rect 6390 1652 6422 1686
rect 6460 1652 6492 1686
rect 6492 1652 6494 1686
rect 6388 1579 6390 1613
rect 6390 1579 6422 1613
rect 6460 1579 6492 1613
rect 6492 1579 6494 1613
rect 6388 1506 6390 1540
rect 6390 1506 6422 1540
rect 6460 1506 6492 1540
rect 6492 1506 6494 1540
rect 6388 1432 6390 1466
rect 6390 1432 6422 1466
rect 6460 1432 6492 1466
rect 6492 1432 6494 1466
rect 6388 1358 6390 1392
rect 6390 1358 6422 1392
rect 6460 1358 6492 1392
rect 6492 1358 6494 1392
rect 6388 1284 6390 1318
rect 6390 1284 6422 1318
rect 6460 1284 6492 1318
rect 6492 1284 6494 1318
rect 6388 1210 6390 1244
rect 6390 1210 6422 1244
rect 6460 1210 6492 1244
rect 6492 1210 6494 1244
rect 6388 1136 6390 1170
rect 6390 1136 6422 1170
rect 6460 1136 6492 1170
rect 6492 1136 6494 1170
rect 6388 1062 6390 1096
rect 6390 1062 6422 1096
rect 6460 1062 6492 1096
rect 6492 1062 6494 1096
rect 6388 988 6390 1022
rect 6390 988 6422 1022
rect 6460 988 6492 1022
rect 6492 988 6494 1022
rect 6388 914 6390 948
rect 6390 914 6422 948
rect 6460 914 6492 948
rect 6492 914 6494 948
rect 6388 840 6390 874
rect 6390 840 6422 874
rect 6460 840 6492 874
rect 6492 840 6494 874
rect 6388 790 6390 800
rect 6390 790 6422 800
rect 6460 790 6492 800
rect 6492 790 6494 800
rect 6388 766 6422 790
rect 6460 766 6494 790
rect 6388 721 6390 726
rect 6390 721 6422 726
rect 6460 721 6492 726
rect 6492 721 6494 726
rect 6388 692 6422 721
rect 6460 692 6494 721
rect 6388 618 6422 652
rect 6460 618 6494 652
rect 6388 548 6422 578
rect 6460 548 6494 578
rect 6388 544 6390 548
rect 6390 544 6422 548
rect 6460 544 6492 548
rect 6492 544 6494 548
rect 6388 479 6422 504
rect 6460 479 6494 504
rect 6388 470 6390 479
rect 6390 470 6422 479
rect 6460 470 6492 479
rect 6492 470 6494 479
rect 6388 410 6422 430
rect 6460 410 6494 430
rect 6388 396 6390 410
rect 6390 396 6422 410
rect 6460 396 6492 410
rect 6492 396 6494 410
rect 6388 341 6422 356
rect 6460 341 6494 356
rect 6388 322 6390 341
rect 6390 322 6422 341
rect 6460 322 6492 341
rect 6492 322 6494 341
rect 6388 272 6422 282
rect 6460 272 6494 282
rect 6388 248 6390 272
rect 6390 248 6422 272
rect 6460 248 6492 272
rect 6492 248 6494 272
rect 6388 203 6422 208
rect 6460 203 6494 208
rect 6388 174 6390 203
rect 6390 174 6422 203
rect 6460 174 6492 203
rect 6492 174 6494 203
rect 6388 100 6390 134
rect 6390 100 6422 134
rect 6460 100 6492 134
rect 6492 100 6494 134
rect 6800 2966 6802 3000
rect 6802 2966 6834 3000
rect 6872 2966 6904 3000
rect 6904 2966 6906 3000
rect 6800 2893 6802 2927
rect 6802 2893 6834 2927
rect 6872 2893 6904 2927
rect 6904 2893 6906 2927
rect 6800 2820 6802 2854
rect 6802 2820 6834 2854
rect 6872 2820 6904 2854
rect 6904 2820 6906 2854
rect 6800 2747 6802 2781
rect 6802 2747 6834 2781
rect 6872 2747 6904 2781
rect 6904 2747 6906 2781
rect 6800 2674 6802 2708
rect 6802 2674 6834 2708
rect 6872 2674 6904 2708
rect 6904 2674 6906 2708
rect 6800 2601 6802 2635
rect 6802 2601 6834 2635
rect 6872 2601 6904 2635
rect 6904 2601 6906 2635
rect 6800 2528 6802 2562
rect 6802 2528 6834 2562
rect 6872 2528 6904 2562
rect 6904 2528 6906 2562
rect 6800 2455 6802 2489
rect 6802 2455 6834 2489
rect 6872 2455 6904 2489
rect 6904 2455 6906 2489
rect 6800 2382 6802 2416
rect 6802 2382 6834 2416
rect 6872 2382 6904 2416
rect 6904 2382 6906 2416
rect 6800 2309 6802 2343
rect 6802 2309 6834 2343
rect 6872 2309 6904 2343
rect 6904 2309 6906 2343
rect 6800 2236 6802 2270
rect 6802 2236 6834 2270
rect 6872 2236 6904 2270
rect 6904 2236 6906 2270
rect 6800 2163 6802 2197
rect 6802 2163 6834 2197
rect 6872 2163 6904 2197
rect 6904 2163 6906 2197
rect 6800 2090 6802 2124
rect 6802 2090 6834 2124
rect 6872 2090 6904 2124
rect 6904 2090 6906 2124
rect 6800 2017 6802 2051
rect 6802 2017 6834 2051
rect 6872 2017 6904 2051
rect 6904 2017 6906 2051
rect 6800 1944 6802 1978
rect 6802 1944 6834 1978
rect 6872 1944 6904 1978
rect 6904 1944 6906 1978
rect 6800 1871 6802 1905
rect 6802 1871 6834 1905
rect 6872 1871 6904 1905
rect 6904 1871 6906 1905
rect 6800 1798 6802 1832
rect 6802 1798 6834 1832
rect 6872 1798 6904 1832
rect 6904 1798 6906 1832
rect 6800 1725 6802 1759
rect 6802 1725 6834 1759
rect 6872 1725 6904 1759
rect 6904 1725 6906 1759
rect 6800 1652 6802 1686
rect 6802 1652 6834 1686
rect 6872 1652 6904 1686
rect 6904 1652 6906 1686
rect 6800 1579 6802 1613
rect 6802 1579 6834 1613
rect 6872 1579 6904 1613
rect 6904 1579 6906 1613
rect 6800 1506 6802 1540
rect 6802 1506 6834 1540
rect 6872 1506 6904 1540
rect 6904 1506 6906 1540
rect 6800 1432 6802 1466
rect 6802 1432 6834 1466
rect 6872 1432 6904 1466
rect 6904 1432 6906 1466
rect 6800 1358 6802 1392
rect 6802 1358 6834 1392
rect 6872 1358 6904 1392
rect 6904 1358 6906 1392
rect 6800 1284 6802 1318
rect 6802 1284 6834 1318
rect 6872 1284 6904 1318
rect 6904 1284 6906 1318
rect 6800 1210 6802 1244
rect 6802 1210 6834 1244
rect 6872 1210 6904 1244
rect 6904 1210 6906 1244
rect 6800 1136 6802 1170
rect 6802 1136 6834 1170
rect 6872 1136 6904 1170
rect 6904 1136 6906 1170
rect 6800 1062 6802 1096
rect 6802 1062 6834 1096
rect 6872 1062 6904 1096
rect 6904 1062 6906 1096
rect 6800 988 6802 1022
rect 6802 988 6834 1022
rect 6872 988 6904 1022
rect 6904 988 6906 1022
rect 6800 914 6802 948
rect 6802 914 6834 948
rect 6872 914 6904 948
rect 6904 914 6906 948
rect 6800 840 6802 874
rect 6802 840 6834 874
rect 6872 840 6904 874
rect 6904 840 6906 874
rect 6800 790 6802 800
rect 6802 790 6834 800
rect 6872 790 6904 800
rect 6904 790 6906 800
rect 6800 766 6834 790
rect 6872 766 6906 790
rect 6800 721 6802 726
rect 6802 721 6834 726
rect 6872 721 6904 726
rect 6904 721 6906 726
rect 6800 692 6834 721
rect 6872 692 6906 721
rect 6800 618 6834 652
rect 6872 618 6906 652
rect 6800 548 6834 578
rect 6872 548 6906 578
rect 6800 544 6802 548
rect 6802 544 6834 548
rect 6872 544 6904 548
rect 6904 544 6906 548
rect 6800 479 6834 504
rect 6872 479 6906 504
rect 6800 470 6802 479
rect 6802 470 6834 479
rect 6872 470 6904 479
rect 6904 470 6906 479
rect 6800 410 6834 430
rect 6872 410 6906 430
rect 6800 396 6802 410
rect 6802 396 6834 410
rect 6872 396 6904 410
rect 6904 396 6906 410
rect 6800 341 6834 356
rect 6872 341 6906 356
rect 6800 322 6802 341
rect 6802 322 6834 341
rect 6872 322 6904 341
rect 6904 322 6906 341
rect 6800 272 6834 282
rect 6872 272 6906 282
rect 6800 248 6802 272
rect 6802 248 6834 272
rect 6872 248 6904 272
rect 6904 248 6906 272
rect 6800 203 6834 208
rect 6872 203 6906 208
rect 6800 174 6802 203
rect 6802 174 6834 203
rect 6872 174 6904 203
rect 6904 174 6906 203
rect 6800 100 6802 134
rect 6802 100 6834 134
rect 6872 100 6904 134
rect 6904 100 6906 134
rect 7212 2966 7214 3000
rect 7214 2966 7246 3000
rect 7284 2966 7316 3000
rect 7316 2966 7318 3000
rect 7212 2893 7214 2927
rect 7214 2893 7246 2927
rect 7284 2893 7316 2927
rect 7316 2893 7318 2927
rect 7212 2820 7214 2854
rect 7214 2820 7246 2854
rect 7284 2820 7316 2854
rect 7316 2820 7318 2854
rect 7212 2747 7214 2781
rect 7214 2747 7246 2781
rect 7284 2747 7316 2781
rect 7316 2747 7318 2781
rect 7212 2674 7214 2708
rect 7214 2674 7246 2708
rect 7284 2674 7316 2708
rect 7316 2674 7318 2708
rect 7212 2601 7214 2635
rect 7214 2601 7246 2635
rect 7284 2601 7316 2635
rect 7316 2601 7318 2635
rect 7212 2528 7214 2562
rect 7214 2528 7246 2562
rect 7284 2528 7316 2562
rect 7316 2528 7318 2562
rect 7212 2455 7214 2489
rect 7214 2455 7246 2489
rect 7284 2455 7316 2489
rect 7316 2455 7318 2489
rect 7212 2382 7214 2416
rect 7214 2382 7246 2416
rect 7284 2382 7316 2416
rect 7316 2382 7318 2416
rect 7212 2309 7214 2343
rect 7214 2309 7246 2343
rect 7284 2309 7316 2343
rect 7316 2309 7318 2343
rect 7212 2236 7214 2270
rect 7214 2236 7246 2270
rect 7284 2236 7316 2270
rect 7316 2236 7318 2270
rect 7212 2163 7214 2197
rect 7214 2163 7246 2197
rect 7284 2163 7316 2197
rect 7316 2163 7318 2197
rect 7212 2090 7214 2124
rect 7214 2090 7246 2124
rect 7284 2090 7316 2124
rect 7316 2090 7318 2124
rect 7212 2017 7214 2051
rect 7214 2017 7246 2051
rect 7284 2017 7316 2051
rect 7316 2017 7318 2051
rect 7212 1944 7214 1978
rect 7214 1944 7246 1978
rect 7284 1944 7316 1978
rect 7316 1944 7318 1978
rect 7212 1871 7214 1905
rect 7214 1871 7246 1905
rect 7284 1871 7316 1905
rect 7316 1871 7318 1905
rect 7212 1798 7214 1832
rect 7214 1798 7246 1832
rect 7284 1798 7316 1832
rect 7316 1798 7318 1832
rect 7212 1725 7214 1759
rect 7214 1725 7246 1759
rect 7284 1725 7316 1759
rect 7316 1725 7318 1759
rect 7212 1652 7214 1686
rect 7214 1652 7246 1686
rect 7284 1652 7316 1686
rect 7316 1652 7318 1686
rect 7212 1579 7214 1613
rect 7214 1579 7246 1613
rect 7284 1579 7316 1613
rect 7316 1579 7318 1613
rect 7212 1506 7214 1540
rect 7214 1506 7246 1540
rect 7284 1506 7316 1540
rect 7316 1506 7318 1540
rect 7212 1432 7214 1466
rect 7214 1432 7246 1466
rect 7284 1432 7316 1466
rect 7316 1432 7318 1466
rect 7212 1358 7214 1392
rect 7214 1358 7246 1392
rect 7284 1358 7316 1392
rect 7316 1358 7318 1392
rect 7212 1284 7214 1318
rect 7214 1284 7246 1318
rect 7284 1284 7316 1318
rect 7316 1284 7318 1318
rect 7212 1210 7214 1244
rect 7214 1210 7246 1244
rect 7284 1210 7316 1244
rect 7316 1210 7318 1244
rect 7212 1136 7214 1170
rect 7214 1136 7246 1170
rect 7284 1136 7316 1170
rect 7316 1136 7318 1170
rect 7212 1062 7214 1096
rect 7214 1062 7246 1096
rect 7284 1062 7316 1096
rect 7316 1062 7318 1096
rect 7212 988 7214 1022
rect 7214 988 7246 1022
rect 7284 988 7316 1022
rect 7316 988 7318 1022
rect 7212 914 7214 948
rect 7214 914 7246 948
rect 7284 914 7316 948
rect 7316 914 7318 948
rect 7212 840 7214 874
rect 7214 840 7246 874
rect 7284 840 7316 874
rect 7316 840 7318 874
rect 7212 790 7214 800
rect 7214 790 7246 800
rect 7284 790 7316 800
rect 7316 790 7318 800
rect 7212 766 7246 790
rect 7284 766 7318 790
rect 7212 721 7214 726
rect 7214 721 7246 726
rect 7284 721 7316 726
rect 7316 721 7318 726
rect 7212 692 7246 721
rect 7284 692 7318 721
rect 7212 618 7246 652
rect 7284 618 7318 652
rect 7212 548 7246 578
rect 7284 548 7318 578
rect 7212 544 7214 548
rect 7214 544 7246 548
rect 7284 544 7316 548
rect 7316 544 7318 548
rect 7212 479 7246 504
rect 7284 479 7318 504
rect 7212 470 7214 479
rect 7214 470 7246 479
rect 7284 470 7316 479
rect 7316 470 7318 479
rect 7212 410 7246 430
rect 7284 410 7318 430
rect 7212 396 7214 410
rect 7214 396 7246 410
rect 7284 396 7316 410
rect 7316 396 7318 410
rect 7212 341 7246 356
rect 7284 341 7318 356
rect 7212 322 7214 341
rect 7214 322 7246 341
rect 7284 322 7316 341
rect 7316 322 7318 341
rect 7212 272 7246 282
rect 7284 272 7318 282
rect 7212 248 7214 272
rect 7214 248 7246 272
rect 7284 248 7316 272
rect 7316 248 7318 272
rect 7212 203 7246 208
rect 7284 203 7318 208
rect 7212 174 7214 203
rect 7214 174 7246 203
rect 7284 174 7316 203
rect 7316 174 7318 203
rect 7212 100 7214 134
rect 7214 100 7246 134
rect 7284 100 7316 134
rect 7316 100 7318 134
rect 7624 2966 7626 3000
rect 7626 2966 7658 3000
rect 7696 2966 7728 3000
rect 7728 2966 7730 3000
rect 7624 2893 7626 2927
rect 7626 2893 7658 2927
rect 7696 2893 7728 2927
rect 7728 2893 7730 2927
rect 7624 2820 7626 2854
rect 7626 2820 7658 2854
rect 7696 2820 7728 2854
rect 7728 2820 7730 2854
rect 7624 2747 7626 2781
rect 7626 2747 7658 2781
rect 7696 2747 7728 2781
rect 7728 2747 7730 2781
rect 7624 2674 7626 2708
rect 7626 2674 7658 2708
rect 7696 2674 7728 2708
rect 7728 2674 7730 2708
rect 7624 2601 7626 2635
rect 7626 2601 7658 2635
rect 7696 2601 7728 2635
rect 7728 2601 7730 2635
rect 7624 2528 7626 2562
rect 7626 2528 7658 2562
rect 7696 2528 7728 2562
rect 7728 2528 7730 2562
rect 7624 2455 7626 2489
rect 7626 2455 7658 2489
rect 7696 2455 7728 2489
rect 7728 2455 7730 2489
rect 7624 2382 7626 2416
rect 7626 2382 7658 2416
rect 7696 2382 7728 2416
rect 7728 2382 7730 2416
rect 7624 2309 7626 2343
rect 7626 2309 7658 2343
rect 7696 2309 7728 2343
rect 7728 2309 7730 2343
rect 7624 2236 7626 2270
rect 7626 2236 7658 2270
rect 7696 2236 7728 2270
rect 7728 2236 7730 2270
rect 7624 2163 7626 2197
rect 7626 2163 7658 2197
rect 7696 2163 7728 2197
rect 7728 2163 7730 2197
rect 7624 2090 7626 2124
rect 7626 2090 7658 2124
rect 7696 2090 7728 2124
rect 7728 2090 7730 2124
rect 7624 2017 7626 2051
rect 7626 2017 7658 2051
rect 7696 2017 7728 2051
rect 7728 2017 7730 2051
rect 7624 1944 7626 1978
rect 7626 1944 7658 1978
rect 7696 1944 7728 1978
rect 7728 1944 7730 1978
rect 7624 1871 7626 1905
rect 7626 1871 7658 1905
rect 7696 1871 7728 1905
rect 7728 1871 7730 1905
rect 7624 1798 7626 1832
rect 7626 1798 7658 1832
rect 7696 1798 7728 1832
rect 7728 1798 7730 1832
rect 7624 1725 7626 1759
rect 7626 1725 7658 1759
rect 7696 1725 7728 1759
rect 7728 1725 7730 1759
rect 7624 1652 7626 1686
rect 7626 1652 7658 1686
rect 7696 1652 7728 1686
rect 7728 1652 7730 1686
rect 7624 1579 7626 1613
rect 7626 1579 7658 1613
rect 7696 1579 7728 1613
rect 7728 1579 7730 1613
rect 7624 1506 7626 1540
rect 7626 1506 7658 1540
rect 7696 1506 7728 1540
rect 7728 1506 7730 1540
rect 7624 1432 7626 1466
rect 7626 1432 7658 1466
rect 7696 1432 7728 1466
rect 7728 1432 7730 1466
rect 7624 1358 7626 1392
rect 7626 1358 7658 1392
rect 7696 1358 7728 1392
rect 7728 1358 7730 1392
rect 7624 1284 7626 1318
rect 7626 1284 7658 1318
rect 7696 1284 7728 1318
rect 7728 1284 7730 1318
rect 7624 1210 7626 1244
rect 7626 1210 7658 1244
rect 7696 1210 7728 1244
rect 7728 1210 7730 1244
rect 7624 1136 7626 1170
rect 7626 1136 7658 1170
rect 7696 1136 7728 1170
rect 7728 1136 7730 1170
rect 7624 1062 7626 1096
rect 7626 1062 7658 1096
rect 7696 1062 7728 1096
rect 7728 1062 7730 1096
rect 7624 988 7626 1022
rect 7626 988 7658 1022
rect 7696 988 7728 1022
rect 7728 988 7730 1022
rect 7624 914 7626 948
rect 7626 914 7658 948
rect 7696 914 7728 948
rect 7728 914 7730 948
rect 7624 840 7626 874
rect 7626 840 7658 874
rect 7696 840 7728 874
rect 7728 840 7730 874
rect 7624 790 7626 800
rect 7626 790 7658 800
rect 7696 790 7728 800
rect 7728 790 7730 800
rect 7624 766 7658 790
rect 7696 766 7730 790
rect 7624 721 7626 726
rect 7626 721 7658 726
rect 7696 721 7728 726
rect 7728 721 7730 726
rect 7624 692 7658 721
rect 7696 692 7730 721
rect 7624 618 7658 652
rect 7696 618 7730 652
rect 7624 548 7658 578
rect 7696 548 7730 578
rect 7624 544 7626 548
rect 7626 544 7658 548
rect 7696 544 7728 548
rect 7728 544 7730 548
rect 7624 479 7658 504
rect 7696 479 7730 504
rect 7624 470 7626 479
rect 7626 470 7658 479
rect 7696 470 7728 479
rect 7728 470 7730 479
rect 7624 410 7658 430
rect 7696 410 7730 430
rect 7624 396 7626 410
rect 7626 396 7658 410
rect 7696 396 7728 410
rect 7728 396 7730 410
rect 7624 341 7658 356
rect 7696 341 7730 356
rect 7624 322 7626 341
rect 7626 322 7658 341
rect 7696 322 7728 341
rect 7728 322 7730 341
rect 7624 272 7658 282
rect 7696 272 7730 282
rect 7624 248 7626 272
rect 7626 248 7658 272
rect 7696 248 7728 272
rect 7728 248 7730 272
rect 7624 203 7658 208
rect 7696 203 7730 208
rect 7624 174 7626 203
rect 7626 174 7658 203
rect 7696 174 7728 203
rect 7728 174 7730 203
rect 7624 100 7626 134
rect 7626 100 7658 134
rect 7696 100 7728 134
rect 7728 100 7730 134
rect 8036 2966 8038 3000
rect 8038 2966 8070 3000
rect 8108 2966 8140 3000
rect 8140 2966 8142 3000
rect 8036 2893 8038 2927
rect 8038 2893 8070 2927
rect 8108 2893 8140 2927
rect 8140 2893 8142 2927
rect 8036 2820 8038 2854
rect 8038 2820 8070 2854
rect 8108 2820 8140 2854
rect 8140 2820 8142 2854
rect 8036 2747 8038 2781
rect 8038 2747 8070 2781
rect 8108 2747 8140 2781
rect 8140 2747 8142 2781
rect 8036 2674 8038 2708
rect 8038 2674 8070 2708
rect 8108 2674 8140 2708
rect 8140 2674 8142 2708
rect 8036 2601 8038 2635
rect 8038 2601 8070 2635
rect 8108 2601 8140 2635
rect 8140 2601 8142 2635
rect 8036 2528 8038 2562
rect 8038 2528 8070 2562
rect 8108 2528 8140 2562
rect 8140 2528 8142 2562
rect 8036 2455 8038 2489
rect 8038 2455 8070 2489
rect 8108 2455 8140 2489
rect 8140 2455 8142 2489
rect 8036 2382 8038 2416
rect 8038 2382 8070 2416
rect 8108 2382 8140 2416
rect 8140 2382 8142 2416
rect 8036 2309 8038 2343
rect 8038 2309 8070 2343
rect 8108 2309 8140 2343
rect 8140 2309 8142 2343
rect 8036 2236 8038 2270
rect 8038 2236 8070 2270
rect 8108 2236 8140 2270
rect 8140 2236 8142 2270
rect 8036 2163 8038 2197
rect 8038 2163 8070 2197
rect 8108 2163 8140 2197
rect 8140 2163 8142 2197
rect 8036 2090 8038 2124
rect 8038 2090 8070 2124
rect 8108 2090 8140 2124
rect 8140 2090 8142 2124
rect 8036 2017 8038 2051
rect 8038 2017 8070 2051
rect 8108 2017 8140 2051
rect 8140 2017 8142 2051
rect 8036 1944 8038 1978
rect 8038 1944 8070 1978
rect 8108 1944 8140 1978
rect 8140 1944 8142 1978
rect 8036 1871 8038 1905
rect 8038 1871 8070 1905
rect 8108 1871 8140 1905
rect 8140 1871 8142 1905
rect 8036 1798 8038 1832
rect 8038 1798 8070 1832
rect 8108 1798 8140 1832
rect 8140 1798 8142 1832
rect 8036 1725 8038 1759
rect 8038 1725 8070 1759
rect 8108 1725 8140 1759
rect 8140 1725 8142 1759
rect 8036 1652 8038 1686
rect 8038 1652 8070 1686
rect 8108 1652 8140 1686
rect 8140 1652 8142 1686
rect 8036 1579 8038 1613
rect 8038 1579 8070 1613
rect 8108 1579 8140 1613
rect 8140 1579 8142 1613
rect 8036 1506 8038 1540
rect 8038 1506 8070 1540
rect 8108 1506 8140 1540
rect 8140 1506 8142 1540
rect 8036 1432 8038 1466
rect 8038 1432 8070 1466
rect 8108 1432 8140 1466
rect 8140 1432 8142 1466
rect 8036 1358 8038 1392
rect 8038 1358 8070 1392
rect 8108 1358 8140 1392
rect 8140 1358 8142 1392
rect 8036 1284 8038 1318
rect 8038 1284 8070 1318
rect 8108 1284 8140 1318
rect 8140 1284 8142 1318
rect 8036 1210 8038 1244
rect 8038 1210 8070 1244
rect 8108 1210 8140 1244
rect 8140 1210 8142 1244
rect 8036 1136 8038 1170
rect 8038 1136 8070 1170
rect 8108 1136 8140 1170
rect 8140 1136 8142 1170
rect 8036 1062 8038 1096
rect 8038 1062 8070 1096
rect 8108 1062 8140 1096
rect 8140 1062 8142 1096
rect 8036 988 8038 1022
rect 8038 988 8070 1022
rect 8108 988 8140 1022
rect 8140 988 8142 1022
rect 8036 914 8038 948
rect 8038 914 8070 948
rect 8108 914 8140 948
rect 8140 914 8142 948
rect 8036 840 8038 874
rect 8038 840 8070 874
rect 8108 840 8140 874
rect 8140 840 8142 874
rect 8036 790 8038 800
rect 8038 790 8070 800
rect 8108 790 8140 800
rect 8140 790 8142 800
rect 8036 766 8070 790
rect 8108 766 8142 790
rect 8036 721 8038 726
rect 8038 721 8070 726
rect 8108 721 8140 726
rect 8140 721 8142 726
rect 8036 692 8070 721
rect 8108 692 8142 721
rect 8036 618 8070 652
rect 8108 618 8142 652
rect 8036 548 8070 578
rect 8108 548 8142 578
rect 8036 544 8038 548
rect 8038 544 8070 548
rect 8108 544 8140 548
rect 8140 544 8142 548
rect 8036 479 8070 504
rect 8108 479 8142 504
rect 8036 470 8038 479
rect 8038 470 8070 479
rect 8108 470 8140 479
rect 8140 470 8142 479
rect 8036 410 8070 430
rect 8108 410 8142 430
rect 8036 396 8038 410
rect 8038 396 8070 410
rect 8108 396 8140 410
rect 8140 396 8142 410
rect 8036 341 8070 356
rect 8108 341 8142 356
rect 8036 322 8038 341
rect 8038 322 8070 341
rect 8108 322 8140 341
rect 8140 322 8142 341
rect 8036 272 8070 282
rect 8108 272 8142 282
rect 8036 248 8038 272
rect 8038 248 8070 272
rect 8108 248 8140 272
rect 8140 248 8142 272
rect 8036 203 8070 208
rect 8108 203 8142 208
rect 8036 174 8038 203
rect 8038 174 8070 203
rect 8108 174 8140 203
rect 8140 174 8142 203
rect 8036 100 8038 134
rect 8038 100 8070 134
rect 8108 100 8140 134
rect 8140 100 8142 134
rect 8448 2966 8450 3000
rect 8450 2966 8482 3000
rect 8520 2966 8552 3000
rect 8552 2966 8554 3000
rect 8448 2893 8450 2927
rect 8450 2893 8482 2927
rect 8520 2893 8552 2927
rect 8552 2893 8554 2927
rect 8448 2820 8450 2854
rect 8450 2820 8482 2854
rect 8520 2820 8552 2854
rect 8552 2820 8554 2854
rect 8448 2747 8450 2781
rect 8450 2747 8482 2781
rect 8520 2747 8552 2781
rect 8552 2747 8554 2781
rect 8448 2674 8450 2708
rect 8450 2674 8482 2708
rect 8520 2674 8552 2708
rect 8552 2674 8554 2708
rect 8448 2601 8450 2635
rect 8450 2601 8482 2635
rect 8520 2601 8552 2635
rect 8552 2601 8554 2635
rect 8448 2528 8450 2562
rect 8450 2528 8482 2562
rect 8520 2528 8552 2562
rect 8552 2528 8554 2562
rect 8448 2455 8450 2489
rect 8450 2455 8482 2489
rect 8520 2455 8552 2489
rect 8552 2455 8554 2489
rect 8448 2382 8450 2416
rect 8450 2382 8482 2416
rect 8520 2382 8552 2416
rect 8552 2382 8554 2416
rect 8448 2309 8450 2343
rect 8450 2309 8482 2343
rect 8520 2309 8552 2343
rect 8552 2309 8554 2343
rect 8448 2236 8450 2270
rect 8450 2236 8482 2270
rect 8520 2236 8552 2270
rect 8552 2236 8554 2270
rect 8448 2163 8450 2197
rect 8450 2163 8482 2197
rect 8520 2163 8552 2197
rect 8552 2163 8554 2197
rect 8448 2090 8450 2124
rect 8450 2090 8482 2124
rect 8520 2090 8552 2124
rect 8552 2090 8554 2124
rect 8448 2017 8450 2051
rect 8450 2017 8482 2051
rect 8520 2017 8552 2051
rect 8552 2017 8554 2051
rect 8448 1944 8450 1978
rect 8450 1944 8482 1978
rect 8520 1944 8552 1978
rect 8552 1944 8554 1978
rect 8448 1871 8450 1905
rect 8450 1871 8482 1905
rect 8520 1871 8552 1905
rect 8552 1871 8554 1905
rect 8448 1798 8450 1832
rect 8450 1798 8482 1832
rect 8520 1798 8552 1832
rect 8552 1798 8554 1832
rect 8448 1725 8450 1759
rect 8450 1725 8482 1759
rect 8520 1725 8552 1759
rect 8552 1725 8554 1759
rect 8448 1652 8450 1686
rect 8450 1652 8482 1686
rect 8520 1652 8552 1686
rect 8552 1652 8554 1686
rect 8448 1579 8450 1613
rect 8450 1579 8482 1613
rect 8520 1579 8552 1613
rect 8552 1579 8554 1613
rect 8448 1506 8450 1540
rect 8450 1506 8482 1540
rect 8520 1506 8552 1540
rect 8552 1506 8554 1540
rect 8448 1432 8450 1466
rect 8450 1432 8482 1466
rect 8520 1432 8552 1466
rect 8552 1432 8554 1466
rect 8448 1358 8450 1392
rect 8450 1358 8482 1392
rect 8520 1358 8552 1392
rect 8552 1358 8554 1392
rect 8448 1284 8450 1318
rect 8450 1284 8482 1318
rect 8520 1284 8552 1318
rect 8552 1284 8554 1318
rect 8448 1210 8450 1244
rect 8450 1210 8482 1244
rect 8520 1210 8552 1244
rect 8552 1210 8554 1244
rect 8448 1136 8450 1170
rect 8450 1136 8482 1170
rect 8520 1136 8552 1170
rect 8552 1136 8554 1170
rect 8448 1062 8450 1096
rect 8450 1062 8482 1096
rect 8520 1062 8552 1096
rect 8552 1062 8554 1096
rect 8448 988 8450 1022
rect 8450 988 8482 1022
rect 8520 988 8552 1022
rect 8552 988 8554 1022
rect 8448 914 8450 948
rect 8450 914 8482 948
rect 8520 914 8552 948
rect 8552 914 8554 948
rect 8448 840 8450 874
rect 8450 840 8482 874
rect 8520 840 8552 874
rect 8552 840 8554 874
rect 8448 790 8450 800
rect 8450 790 8482 800
rect 8520 790 8552 800
rect 8552 790 8554 800
rect 8448 766 8482 790
rect 8520 766 8554 790
rect 8448 721 8450 726
rect 8450 721 8482 726
rect 8520 721 8552 726
rect 8552 721 8554 726
rect 8448 692 8482 721
rect 8520 692 8554 721
rect 8448 618 8482 652
rect 8520 618 8554 652
rect 8448 548 8482 578
rect 8520 548 8554 578
rect 8448 544 8450 548
rect 8450 544 8482 548
rect 8520 544 8552 548
rect 8552 544 8554 548
rect 8448 479 8482 504
rect 8520 479 8554 504
rect 8448 470 8450 479
rect 8450 470 8482 479
rect 8520 470 8552 479
rect 8552 470 8554 479
rect 8448 410 8482 430
rect 8520 410 8554 430
rect 8448 396 8450 410
rect 8450 396 8482 410
rect 8520 396 8552 410
rect 8552 396 8554 410
rect 8448 341 8482 356
rect 8520 341 8554 356
rect 8448 322 8450 341
rect 8450 322 8482 341
rect 8520 322 8552 341
rect 8552 322 8554 341
rect 8448 272 8482 282
rect 8520 272 8554 282
rect 8448 248 8450 272
rect 8450 248 8482 272
rect 8520 248 8552 272
rect 8552 248 8554 272
rect 8448 203 8482 208
rect 8520 203 8554 208
rect 8448 174 8450 203
rect 8450 174 8482 203
rect 8520 174 8552 203
rect 8552 174 8554 203
rect 8448 100 8450 134
rect 8450 100 8482 134
rect 8520 100 8552 134
rect 8552 100 8554 134
rect 8860 2966 8862 3000
rect 8862 2966 8894 3000
rect 8932 2966 8964 3000
rect 8964 2966 8966 3000
rect 8860 2893 8862 2927
rect 8862 2893 8894 2927
rect 8932 2893 8964 2927
rect 8964 2893 8966 2927
rect 8860 2820 8862 2854
rect 8862 2820 8894 2854
rect 8932 2820 8964 2854
rect 8964 2820 8966 2854
rect 8860 2747 8862 2781
rect 8862 2747 8894 2781
rect 8932 2747 8964 2781
rect 8964 2747 8966 2781
rect 8860 2674 8862 2708
rect 8862 2674 8894 2708
rect 8932 2674 8964 2708
rect 8964 2674 8966 2708
rect 8860 2601 8862 2635
rect 8862 2601 8894 2635
rect 8932 2601 8964 2635
rect 8964 2601 8966 2635
rect 8860 2528 8862 2562
rect 8862 2528 8894 2562
rect 8932 2528 8964 2562
rect 8964 2528 8966 2562
rect 8860 2455 8862 2489
rect 8862 2455 8894 2489
rect 8932 2455 8964 2489
rect 8964 2455 8966 2489
rect 8860 2382 8862 2416
rect 8862 2382 8894 2416
rect 8932 2382 8964 2416
rect 8964 2382 8966 2416
rect 8860 2309 8862 2343
rect 8862 2309 8894 2343
rect 8932 2309 8964 2343
rect 8964 2309 8966 2343
rect 8860 2236 8862 2270
rect 8862 2236 8894 2270
rect 8932 2236 8964 2270
rect 8964 2236 8966 2270
rect 8860 2163 8862 2197
rect 8862 2163 8894 2197
rect 8932 2163 8964 2197
rect 8964 2163 8966 2197
rect 8860 2090 8862 2124
rect 8862 2090 8894 2124
rect 8932 2090 8964 2124
rect 8964 2090 8966 2124
rect 8860 2017 8862 2051
rect 8862 2017 8894 2051
rect 8932 2017 8964 2051
rect 8964 2017 8966 2051
rect 8860 1944 8862 1978
rect 8862 1944 8894 1978
rect 8932 1944 8964 1978
rect 8964 1944 8966 1978
rect 8860 1871 8862 1905
rect 8862 1871 8894 1905
rect 8932 1871 8964 1905
rect 8964 1871 8966 1905
rect 8860 1798 8862 1832
rect 8862 1798 8894 1832
rect 8932 1798 8964 1832
rect 8964 1798 8966 1832
rect 8860 1725 8862 1759
rect 8862 1725 8894 1759
rect 8932 1725 8964 1759
rect 8964 1725 8966 1759
rect 8860 1652 8862 1686
rect 8862 1652 8894 1686
rect 8932 1652 8964 1686
rect 8964 1652 8966 1686
rect 8860 1579 8862 1613
rect 8862 1579 8894 1613
rect 8932 1579 8964 1613
rect 8964 1579 8966 1613
rect 8860 1506 8862 1540
rect 8862 1506 8894 1540
rect 8932 1506 8964 1540
rect 8964 1506 8966 1540
rect 8860 1432 8862 1466
rect 8862 1432 8894 1466
rect 8932 1432 8964 1466
rect 8964 1432 8966 1466
rect 8860 1358 8862 1392
rect 8862 1358 8894 1392
rect 8932 1358 8964 1392
rect 8964 1358 8966 1392
rect 8860 1284 8862 1318
rect 8862 1284 8894 1318
rect 8932 1284 8964 1318
rect 8964 1284 8966 1318
rect 8860 1210 8862 1244
rect 8862 1210 8894 1244
rect 8932 1210 8964 1244
rect 8964 1210 8966 1244
rect 8860 1136 8862 1170
rect 8862 1136 8894 1170
rect 8932 1136 8964 1170
rect 8964 1136 8966 1170
rect 8860 1062 8862 1096
rect 8862 1062 8894 1096
rect 8932 1062 8964 1096
rect 8964 1062 8966 1096
rect 8860 988 8862 1022
rect 8862 988 8894 1022
rect 8932 988 8964 1022
rect 8964 988 8966 1022
rect 8860 914 8862 948
rect 8862 914 8894 948
rect 8932 914 8964 948
rect 8964 914 8966 948
rect 8860 840 8862 874
rect 8862 840 8894 874
rect 8932 840 8964 874
rect 8964 840 8966 874
rect 8860 790 8862 800
rect 8862 790 8894 800
rect 8932 790 8964 800
rect 8964 790 8966 800
rect 8860 766 8894 790
rect 8932 766 8966 790
rect 8860 721 8862 726
rect 8862 721 8894 726
rect 8932 721 8964 726
rect 8964 721 8966 726
rect 8860 692 8894 721
rect 8932 692 8966 721
rect 8860 618 8894 652
rect 8932 618 8966 652
rect 8860 548 8894 578
rect 8932 548 8966 578
rect 8860 544 8862 548
rect 8862 544 8894 548
rect 8932 544 8964 548
rect 8964 544 8966 548
rect 8860 479 8894 504
rect 8932 479 8966 504
rect 8860 470 8862 479
rect 8862 470 8894 479
rect 8932 470 8964 479
rect 8964 470 8966 479
rect 8860 410 8894 430
rect 8932 410 8966 430
rect 8860 396 8862 410
rect 8862 396 8894 410
rect 8932 396 8964 410
rect 8964 396 8966 410
rect 8860 341 8894 356
rect 8932 341 8966 356
rect 8860 322 8862 341
rect 8862 322 8894 341
rect 8932 322 8964 341
rect 8964 322 8966 341
rect 8860 272 8894 282
rect 8932 272 8966 282
rect 8860 248 8862 272
rect 8862 248 8894 272
rect 8932 248 8964 272
rect 8964 248 8966 272
rect 8860 203 8894 208
rect 8932 203 8966 208
rect 8860 174 8862 203
rect 8862 174 8894 203
rect 8932 174 8964 203
rect 8964 174 8966 203
rect 8860 100 8862 134
rect 8862 100 8894 134
rect 8932 100 8964 134
rect 8964 100 8966 134
rect 9272 2966 9274 3000
rect 9274 2966 9306 3000
rect 9344 2966 9376 3000
rect 9376 2966 9378 3000
rect 9272 2893 9274 2927
rect 9274 2893 9306 2927
rect 9344 2893 9376 2927
rect 9376 2893 9378 2927
rect 9272 2820 9274 2854
rect 9274 2820 9306 2854
rect 9344 2820 9376 2854
rect 9376 2820 9378 2854
rect 9272 2747 9274 2781
rect 9274 2747 9306 2781
rect 9344 2747 9376 2781
rect 9376 2747 9378 2781
rect 9272 2674 9274 2708
rect 9274 2674 9306 2708
rect 9344 2674 9376 2708
rect 9376 2674 9378 2708
rect 9272 2601 9274 2635
rect 9274 2601 9306 2635
rect 9344 2601 9376 2635
rect 9376 2601 9378 2635
rect 9272 2528 9274 2562
rect 9274 2528 9306 2562
rect 9344 2528 9376 2562
rect 9376 2528 9378 2562
rect 9272 2455 9274 2489
rect 9274 2455 9306 2489
rect 9344 2455 9376 2489
rect 9376 2455 9378 2489
rect 9272 2382 9274 2416
rect 9274 2382 9306 2416
rect 9344 2382 9376 2416
rect 9376 2382 9378 2416
rect 9272 2309 9274 2343
rect 9274 2309 9306 2343
rect 9344 2309 9376 2343
rect 9376 2309 9378 2343
rect 9272 2236 9274 2270
rect 9274 2236 9306 2270
rect 9344 2236 9376 2270
rect 9376 2236 9378 2270
rect 9272 2163 9274 2197
rect 9274 2163 9306 2197
rect 9344 2163 9376 2197
rect 9376 2163 9378 2197
rect 9272 2090 9274 2124
rect 9274 2090 9306 2124
rect 9344 2090 9376 2124
rect 9376 2090 9378 2124
rect 9272 2017 9274 2051
rect 9274 2017 9306 2051
rect 9344 2017 9376 2051
rect 9376 2017 9378 2051
rect 9272 1944 9274 1978
rect 9274 1944 9306 1978
rect 9344 1944 9376 1978
rect 9376 1944 9378 1978
rect 9272 1871 9274 1905
rect 9274 1871 9306 1905
rect 9344 1871 9376 1905
rect 9376 1871 9378 1905
rect 9272 1798 9274 1832
rect 9274 1798 9306 1832
rect 9344 1798 9376 1832
rect 9376 1798 9378 1832
rect 9272 1725 9274 1759
rect 9274 1725 9306 1759
rect 9344 1725 9376 1759
rect 9376 1725 9378 1759
rect 9272 1652 9274 1686
rect 9274 1652 9306 1686
rect 9344 1652 9376 1686
rect 9376 1652 9378 1686
rect 9272 1579 9274 1613
rect 9274 1579 9306 1613
rect 9344 1579 9376 1613
rect 9376 1579 9378 1613
rect 9272 1506 9274 1540
rect 9274 1506 9306 1540
rect 9344 1506 9376 1540
rect 9376 1506 9378 1540
rect 9272 1432 9274 1466
rect 9274 1432 9306 1466
rect 9344 1432 9376 1466
rect 9376 1432 9378 1466
rect 9272 1358 9274 1392
rect 9274 1358 9306 1392
rect 9344 1358 9376 1392
rect 9376 1358 9378 1392
rect 9272 1284 9274 1318
rect 9274 1284 9306 1318
rect 9344 1284 9376 1318
rect 9376 1284 9378 1318
rect 9272 1210 9274 1244
rect 9274 1210 9306 1244
rect 9344 1210 9376 1244
rect 9376 1210 9378 1244
rect 9272 1136 9274 1170
rect 9274 1136 9306 1170
rect 9344 1136 9376 1170
rect 9376 1136 9378 1170
rect 9272 1062 9274 1096
rect 9274 1062 9306 1096
rect 9344 1062 9376 1096
rect 9376 1062 9378 1096
rect 9272 988 9274 1022
rect 9274 988 9306 1022
rect 9344 988 9376 1022
rect 9376 988 9378 1022
rect 9272 914 9274 948
rect 9274 914 9306 948
rect 9344 914 9376 948
rect 9376 914 9378 948
rect 9272 840 9274 874
rect 9274 840 9306 874
rect 9344 840 9376 874
rect 9376 840 9378 874
rect 9272 790 9274 800
rect 9274 790 9306 800
rect 9344 790 9376 800
rect 9376 790 9378 800
rect 9272 766 9306 790
rect 9344 766 9378 790
rect 9272 721 9274 726
rect 9274 721 9306 726
rect 9344 721 9376 726
rect 9376 721 9378 726
rect 9272 692 9306 721
rect 9344 692 9378 721
rect 9272 618 9306 652
rect 9344 618 9378 652
rect 9272 548 9306 578
rect 9344 548 9378 578
rect 9272 544 9274 548
rect 9274 544 9306 548
rect 9344 544 9376 548
rect 9376 544 9378 548
rect 9272 479 9306 504
rect 9344 479 9378 504
rect 9272 470 9274 479
rect 9274 470 9306 479
rect 9344 470 9376 479
rect 9376 470 9378 479
rect 9272 410 9306 430
rect 9344 410 9378 430
rect 9272 396 9274 410
rect 9274 396 9306 410
rect 9344 396 9376 410
rect 9376 396 9378 410
rect 9272 341 9306 356
rect 9344 341 9378 356
rect 9272 322 9274 341
rect 9274 322 9306 341
rect 9344 322 9376 341
rect 9376 322 9378 341
rect 9272 272 9306 282
rect 9344 272 9378 282
rect 9272 248 9274 272
rect 9274 248 9306 272
rect 9344 248 9376 272
rect 9376 248 9378 272
rect 9272 203 9306 208
rect 9344 203 9378 208
rect 9272 174 9274 203
rect 9274 174 9306 203
rect 9344 174 9376 203
rect 9376 174 9378 203
rect 9272 100 9274 134
rect 9274 100 9306 134
rect 9344 100 9376 134
rect 9376 100 9378 134
rect 9684 2966 9686 3000
rect 9686 2966 9718 3000
rect 9756 2966 9788 3000
rect 9788 2966 9790 3000
rect 9684 2893 9686 2927
rect 9686 2893 9718 2927
rect 9756 2893 9788 2927
rect 9788 2893 9790 2927
rect 9684 2820 9686 2854
rect 9686 2820 9718 2854
rect 9756 2820 9788 2854
rect 9788 2820 9790 2854
rect 9684 2747 9686 2781
rect 9686 2747 9718 2781
rect 9756 2747 9788 2781
rect 9788 2747 9790 2781
rect 9684 2674 9686 2708
rect 9686 2674 9718 2708
rect 9756 2674 9788 2708
rect 9788 2674 9790 2708
rect 9684 2601 9686 2635
rect 9686 2601 9718 2635
rect 9756 2601 9788 2635
rect 9788 2601 9790 2635
rect 9684 2528 9686 2562
rect 9686 2528 9718 2562
rect 9756 2528 9788 2562
rect 9788 2528 9790 2562
rect 9684 2455 9686 2489
rect 9686 2455 9718 2489
rect 9756 2455 9788 2489
rect 9788 2455 9790 2489
rect 9684 2382 9686 2416
rect 9686 2382 9718 2416
rect 9756 2382 9788 2416
rect 9788 2382 9790 2416
rect 9684 2309 9686 2343
rect 9686 2309 9718 2343
rect 9756 2309 9788 2343
rect 9788 2309 9790 2343
rect 9684 2236 9686 2270
rect 9686 2236 9718 2270
rect 9756 2236 9788 2270
rect 9788 2236 9790 2270
rect 9684 2163 9686 2197
rect 9686 2163 9718 2197
rect 9756 2163 9788 2197
rect 9788 2163 9790 2197
rect 9684 2090 9686 2124
rect 9686 2090 9718 2124
rect 9756 2090 9788 2124
rect 9788 2090 9790 2124
rect 9684 2017 9686 2051
rect 9686 2017 9718 2051
rect 9756 2017 9788 2051
rect 9788 2017 9790 2051
rect 9684 1944 9686 1978
rect 9686 1944 9718 1978
rect 9756 1944 9788 1978
rect 9788 1944 9790 1978
rect 9684 1871 9686 1905
rect 9686 1871 9718 1905
rect 9756 1871 9788 1905
rect 9788 1871 9790 1905
rect 9684 1798 9686 1832
rect 9686 1798 9718 1832
rect 9756 1798 9788 1832
rect 9788 1798 9790 1832
rect 9684 1725 9686 1759
rect 9686 1725 9718 1759
rect 9756 1725 9788 1759
rect 9788 1725 9790 1759
rect 9684 1652 9686 1686
rect 9686 1652 9718 1686
rect 9756 1652 9788 1686
rect 9788 1652 9790 1686
rect 9684 1579 9686 1613
rect 9686 1579 9718 1613
rect 9756 1579 9788 1613
rect 9788 1579 9790 1613
rect 9684 1506 9686 1540
rect 9686 1506 9718 1540
rect 9756 1506 9788 1540
rect 9788 1506 9790 1540
rect 9684 1432 9686 1466
rect 9686 1432 9718 1466
rect 9756 1432 9788 1466
rect 9788 1432 9790 1466
rect 9684 1358 9686 1392
rect 9686 1358 9718 1392
rect 9756 1358 9788 1392
rect 9788 1358 9790 1392
rect 9684 1284 9686 1318
rect 9686 1284 9718 1318
rect 9756 1284 9788 1318
rect 9788 1284 9790 1318
rect 9684 1210 9686 1244
rect 9686 1210 9718 1244
rect 9756 1210 9788 1244
rect 9788 1210 9790 1244
rect 9684 1136 9686 1170
rect 9686 1136 9718 1170
rect 9756 1136 9788 1170
rect 9788 1136 9790 1170
rect 9684 1062 9686 1096
rect 9686 1062 9718 1096
rect 9756 1062 9788 1096
rect 9788 1062 9790 1096
rect 9684 988 9686 1022
rect 9686 988 9718 1022
rect 9756 988 9788 1022
rect 9788 988 9790 1022
rect 9684 914 9686 948
rect 9686 914 9718 948
rect 9756 914 9788 948
rect 9788 914 9790 948
rect 9684 840 9686 874
rect 9686 840 9718 874
rect 9756 840 9788 874
rect 9788 840 9790 874
rect 9684 790 9686 800
rect 9686 790 9718 800
rect 9756 790 9788 800
rect 9788 790 9790 800
rect 9684 766 9718 790
rect 9756 766 9790 790
rect 9684 721 9686 726
rect 9686 721 9718 726
rect 9756 721 9788 726
rect 9788 721 9790 726
rect 9684 692 9718 721
rect 9756 692 9790 721
rect 9684 618 9718 652
rect 9756 618 9790 652
rect 9684 548 9718 578
rect 9756 548 9790 578
rect 9684 544 9686 548
rect 9686 544 9718 548
rect 9756 544 9788 548
rect 9788 544 9790 548
rect 9684 479 9718 504
rect 9756 479 9790 504
rect 9684 470 9686 479
rect 9686 470 9718 479
rect 9756 470 9788 479
rect 9788 470 9790 479
rect 9684 410 9718 430
rect 9756 410 9790 430
rect 9684 396 9686 410
rect 9686 396 9718 410
rect 9756 396 9788 410
rect 9788 396 9790 410
rect 9684 341 9718 356
rect 9756 341 9790 356
rect 9684 322 9686 341
rect 9686 322 9718 341
rect 9756 322 9788 341
rect 9788 322 9790 341
rect 9684 272 9718 282
rect 9756 272 9790 282
rect 9684 248 9686 272
rect 9686 248 9718 272
rect 9756 248 9788 272
rect 9788 248 9790 272
rect 9684 203 9718 208
rect 9756 203 9790 208
rect 9684 174 9686 203
rect 9686 174 9718 203
rect 9756 174 9788 203
rect 9788 174 9790 203
rect 9684 100 9686 134
rect 9686 100 9718 134
rect 9756 100 9788 134
rect 9788 100 9790 134
rect 10096 2966 10098 3000
rect 10098 2966 10130 3000
rect 10168 2966 10200 3000
rect 10200 2966 10202 3000
rect 10096 2893 10098 2927
rect 10098 2893 10130 2927
rect 10168 2893 10200 2927
rect 10200 2893 10202 2927
rect 10096 2820 10098 2854
rect 10098 2820 10130 2854
rect 10168 2820 10200 2854
rect 10200 2820 10202 2854
rect 10096 2747 10098 2781
rect 10098 2747 10130 2781
rect 10168 2747 10200 2781
rect 10200 2747 10202 2781
rect 10096 2674 10098 2708
rect 10098 2674 10130 2708
rect 10168 2674 10200 2708
rect 10200 2674 10202 2708
rect 10096 2601 10098 2635
rect 10098 2601 10130 2635
rect 10168 2601 10200 2635
rect 10200 2601 10202 2635
rect 10096 2528 10098 2562
rect 10098 2528 10130 2562
rect 10168 2528 10200 2562
rect 10200 2528 10202 2562
rect 10096 2455 10098 2489
rect 10098 2455 10130 2489
rect 10168 2455 10200 2489
rect 10200 2455 10202 2489
rect 10096 2382 10098 2416
rect 10098 2382 10130 2416
rect 10168 2382 10200 2416
rect 10200 2382 10202 2416
rect 10096 2309 10098 2343
rect 10098 2309 10130 2343
rect 10168 2309 10200 2343
rect 10200 2309 10202 2343
rect 10096 2236 10098 2270
rect 10098 2236 10130 2270
rect 10168 2236 10200 2270
rect 10200 2236 10202 2270
rect 10096 2163 10098 2197
rect 10098 2163 10130 2197
rect 10168 2163 10200 2197
rect 10200 2163 10202 2197
rect 10096 2090 10098 2124
rect 10098 2090 10130 2124
rect 10168 2090 10200 2124
rect 10200 2090 10202 2124
rect 10096 2017 10098 2051
rect 10098 2017 10130 2051
rect 10168 2017 10200 2051
rect 10200 2017 10202 2051
rect 10096 1944 10098 1978
rect 10098 1944 10130 1978
rect 10168 1944 10200 1978
rect 10200 1944 10202 1978
rect 10096 1871 10098 1905
rect 10098 1871 10130 1905
rect 10168 1871 10200 1905
rect 10200 1871 10202 1905
rect 10096 1798 10098 1832
rect 10098 1798 10130 1832
rect 10168 1798 10200 1832
rect 10200 1798 10202 1832
rect 10096 1725 10098 1759
rect 10098 1725 10130 1759
rect 10168 1725 10200 1759
rect 10200 1725 10202 1759
rect 10096 1652 10098 1686
rect 10098 1652 10130 1686
rect 10168 1652 10200 1686
rect 10200 1652 10202 1686
rect 10096 1579 10098 1613
rect 10098 1579 10130 1613
rect 10168 1579 10200 1613
rect 10200 1579 10202 1613
rect 10096 1506 10098 1540
rect 10098 1506 10130 1540
rect 10168 1506 10200 1540
rect 10200 1506 10202 1540
rect 10096 1432 10098 1466
rect 10098 1432 10130 1466
rect 10168 1432 10200 1466
rect 10200 1432 10202 1466
rect 10096 1358 10098 1392
rect 10098 1358 10130 1392
rect 10168 1358 10200 1392
rect 10200 1358 10202 1392
rect 10096 1284 10098 1318
rect 10098 1284 10130 1318
rect 10168 1284 10200 1318
rect 10200 1284 10202 1318
rect 10096 1210 10098 1244
rect 10098 1210 10130 1244
rect 10168 1210 10200 1244
rect 10200 1210 10202 1244
rect 10096 1136 10098 1170
rect 10098 1136 10130 1170
rect 10168 1136 10200 1170
rect 10200 1136 10202 1170
rect 10096 1062 10098 1096
rect 10098 1062 10130 1096
rect 10168 1062 10200 1096
rect 10200 1062 10202 1096
rect 10096 988 10098 1022
rect 10098 988 10130 1022
rect 10168 988 10200 1022
rect 10200 988 10202 1022
rect 10096 914 10098 948
rect 10098 914 10130 948
rect 10168 914 10200 948
rect 10200 914 10202 948
rect 10096 840 10098 874
rect 10098 840 10130 874
rect 10168 840 10200 874
rect 10200 840 10202 874
rect 10096 790 10098 800
rect 10098 790 10130 800
rect 10168 790 10200 800
rect 10200 790 10202 800
rect 10096 766 10130 790
rect 10168 766 10202 790
rect 10096 721 10098 726
rect 10098 721 10130 726
rect 10168 721 10200 726
rect 10200 721 10202 726
rect 10096 692 10130 721
rect 10168 692 10202 721
rect 10096 618 10130 652
rect 10168 618 10202 652
rect 10096 548 10130 578
rect 10168 548 10202 578
rect 10096 544 10098 548
rect 10098 544 10130 548
rect 10168 544 10200 548
rect 10200 544 10202 548
rect 10096 479 10130 504
rect 10168 479 10202 504
rect 10096 470 10098 479
rect 10098 470 10130 479
rect 10168 470 10200 479
rect 10200 470 10202 479
rect 10096 410 10130 430
rect 10168 410 10202 430
rect 10096 396 10098 410
rect 10098 396 10130 410
rect 10168 396 10200 410
rect 10200 396 10202 410
rect 10096 341 10130 356
rect 10168 341 10202 356
rect 10096 322 10098 341
rect 10098 322 10130 341
rect 10168 322 10200 341
rect 10200 322 10202 341
rect 10096 272 10130 282
rect 10168 272 10202 282
rect 10096 248 10098 272
rect 10098 248 10130 272
rect 10168 248 10200 272
rect 10200 248 10202 272
rect 10096 203 10130 208
rect 10168 203 10202 208
rect 10096 174 10098 203
rect 10098 174 10130 203
rect 10168 174 10200 203
rect 10200 174 10202 203
rect 10096 100 10098 134
rect 10098 100 10130 134
rect 10168 100 10200 134
rect 10200 100 10202 134
rect 10508 2966 10510 3000
rect 10510 2966 10542 3000
rect 10580 2966 10612 3000
rect 10612 2966 10614 3000
rect 10508 2893 10510 2927
rect 10510 2893 10542 2927
rect 10580 2893 10612 2927
rect 10612 2893 10614 2927
rect 10508 2820 10510 2854
rect 10510 2820 10542 2854
rect 10580 2820 10612 2854
rect 10612 2820 10614 2854
rect 10508 2747 10510 2781
rect 10510 2747 10542 2781
rect 10580 2747 10612 2781
rect 10612 2747 10614 2781
rect 10508 2674 10510 2708
rect 10510 2674 10542 2708
rect 10580 2674 10612 2708
rect 10612 2674 10614 2708
rect 10508 2601 10510 2635
rect 10510 2601 10542 2635
rect 10580 2601 10612 2635
rect 10612 2601 10614 2635
rect 10508 2528 10510 2562
rect 10510 2528 10542 2562
rect 10580 2528 10612 2562
rect 10612 2528 10614 2562
rect 10508 2455 10510 2489
rect 10510 2455 10542 2489
rect 10580 2455 10612 2489
rect 10612 2455 10614 2489
rect 10508 2382 10510 2416
rect 10510 2382 10542 2416
rect 10580 2382 10612 2416
rect 10612 2382 10614 2416
rect 10508 2309 10510 2343
rect 10510 2309 10542 2343
rect 10580 2309 10612 2343
rect 10612 2309 10614 2343
rect 10508 2236 10510 2270
rect 10510 2236 10542 2270
rect 10580 2236 10612 2270
rect 10612 2236 10614 2270
rect 10508 2163 10510 2197
rect 10510 2163 10542 2197
rect 10580 2163 10612 2197
rect 10612 2163 10614 2197
rect 10508 2090 10510 2124
rect 10510 2090 10542 2124
rect 10580 2090 10612 2124
rect 10612 2090 10614 2124
rect 10508 2017 10510 2051
rect 10510 2017 10542 2051
rect 10580 2017 10612 2051
rect 10612 2017 10614 2051
rect 10508 1944 10510 1978
rect 10510 1944 10542 1978
rect 10580 1944 10612 1978
rect 10612 1944 10614 1978
rect 10508 1871 10510 1905
rect 10510 1871 10542 1905
rect 10580 1871 10612 1905
rect 10612 1871 10614 1905
rect 10508 1798 10510 1832
rect 10510 1798 10542 1832
rect 10580 1798 10612 1832
rect 10612 1798 10614 1832
rect 10508 1725 10510 1759
rect 10510 1725 10542 1759
rect 10580 1725 10612 1759
rect 10612 1725 10614 1759
rect 10508 1652 10510 1686
rect 10510 1652 10542 1686
rect 10580 1652 10612 1686
rect 10612 1652 10614 1686
rect 10508 1579 10510 1613
rect 10510 1579 10542 1613
rect 10580 1579 10612 1613
rect 10612 1579 10614 1613
rect 10508 1506 10510 1540
rect 10510 1506 10542 1540
rect 10580 1506 10612 1540
rect 10612 1506 10614 1540
rect 10508 1432 10510 1466
rect 10510 1432 10542 1466
rect 10580 1432 10612 1466
rect 10612 1432 10614 1466
rect 10508 1358 10510 1392
rect 10510 1358 10542 1392
rect 10580 1358 10612 1392
rect 10612 1358 10614 1392
rect 10508 1284 10510 1318
rect 10510 1284 10542 1318
rect 10580 1284 10612 1318
rect 10612 1284 10614 1318
rect 10508 1210 10510 1244
rect 10510 1210 10542 1244
rect 10580 1210 10612 1244
rect 10612 1210 10614 1244
rect 10508 1136 10510 1170
rect 10510 1136 10542 1170
rect 10580 1136 10612 1170
rect 10612 1136 10614 1170
rect 10508 1062 10510 1096
rect 10510 1062 10542 1096
rect 10580 1062 10612 1096
rect 10612 1062 10614 1096
rect 10508 988 10510 1022
rect 10510 988 10542 1022
rect 10580 988 10612 1022
rect 10612 988 10614 1022
rect 10508 914 10510 948
rect 10510 914 10542 948
rect 10580 914 10612 948
rect 10612 914 10614 948
rect 10508 840 10510 874
rect 10510 840 10542 874
rect 10580 840 10612 874
rect 10612 840 10614 874
rect 10508 790 10510 800
rect 10510 790 10542 800
rect 10580 790 10612 800
rect 10612 790 10614 800
rect 10508 766 10542 790
rect 10580 766 10614 790
rect 10508 721 10510 726
rect 10510 721 10542 726
rect 10580 721 10612 726
rect 10612 721 10614 726
rect 10508 692 10542 721
rect 10580 692 10614 721
rect 10508 618 10542 652
rect 10580 618 10614 652
rect 10508 548 10542 578
rect 10580 548 10614 578
rect 10508 544 10510 548
rect 10510 544 10542 548
rect 10580 544 10612 548
rect 10612 544 10614 548
rect 10508 479 10542 504
rect 10580 479 10614 504
rect 10508 470 10510 479
rect 10510 470 10542 479
rect 10580 470 10612 479
rect 10612 470 10614 479
rect 10508 410 10542 430
rect 10580 410 10614 430
rect 10508 396 10510 410
rect 10510 396 10542 410
rect 10580 396 10612 410
rect 10612 396 10614 410
rect 10508 341 10542 356
rect 10580 341 10614 356
rect 10508 322 10510 341
rect 10510 322 10542 341
rect 10580 322 10612 341
rect 10612 322 10614 341
rect 10508 272 10542 282
rect 10580 272 10614 282
rect 10508 248 10510 272
rect 10510 248 10542 272
rect 10580 248 10612 272
rect 10612 248 10614 272
rect 10508 203 10542 208
rect 10580 203 10614 208
rect 10508 174 10510 203
rect 10510 174 10542 203
rect 10580 174 10612 203
rect 10612 174 10614 203
rect 10508 100 10510 134
rect 10510 100 10542 134
rect 10580 100 10612 134
rect 10612 100 10614 134
rect 10920 2966 10922 3000
rect 10922 2966 10954 3000
rect 10992 2966 11024 3000
rect 11024 2966 11026 3000
rect 10920 2893 10922 2927
rect 10922 2893 10954 2927
rect 10992 2893 11024 2927
rect 11024 2893 11026 2927
rect 10920 2820 10922 2854
rect 10922 2820 10954 2854
rect 10992 2820 11024 2854
rect 11024 2820 11026 2854
rect 10920 2747 10922 2781
rect 10922 2747 10954 2781
rect 10992 2747 11024 2781
rect 11024 2747 11026 2781
rect 10920 2674 10922 2708
rect 10922 2674 10954 2708
rect 10992 2674 11024 2708
rect 11024 2674 11026 2708
rect 10920 2601 10922 2635
rect 10922 2601 10954 2635
rect 10992 2601 11024 2635
rect 11024 2601 11026 2635
rect 10920 2528 10922 2562
rect 10922 2528 10954 2562
rect 10992 2528 11024 2562
rect 11024 2528 11026 2562
rect 10920 2455 10922 2489
rect 10922 2455 10954 2489
rect 10992 2455 11024 2489
rect 11024 2455 11026 2489
rect 10920 2382 10922 2416
rect 10922 2382 10954 2416
rect 10992 2382 11024 2416
rect 11024 2382 11026 2416
rect 10920 2309 10922 2343
rect 10922 2309 10954 2343
rect 10992 2309 11024 2343
rect 11024 2309 11026 2343
rect 10920 2236 10922 2270
rect 10922 2236 10954 2270
rect 10992 2236 11024 2270
rect 11024 2236 11026 2270
rect 10920 2163 10922 2197
rect 10922 2163 10954 2197
rect 10992 2163 11024 2197
rect 11024 2163 11026 2197
rect 10920 2090 10922 2124
rect 10922 2090 10954 2124
rect 10992 2090 11024 2124
rect 11024 2090 11026 2124
rect 10920 2017 10922 2051
rect 10922 2017 10954 2051
rect 10992 2017 11024 2051
rect 11024 2017 11026 2051
rect 10920 1944 10922 1978
rect 10922 1944 10954 1978
rect 10992 1944 11024 1978
rect 11024 1944 11026 1978
rect 10920 1871 10922 1905
rect 10922 1871 10954 1905
rect 10992 1871 11024 1905
rect 11024 1871 11026 1905
rect 10920 1798 10922 1832
rect 10922 1798 10954 1832
rect 10992 1798 11024 1832
rect 11024 1798 11026 1832
rect 10920 1725 10922 1759
rect 10922 1725 10954 1759
rect 10992 1725 11024 1759
rect 11024 1725 11026 1759
rect 10920 1652 10922 1686
rect 10922 1652 10954 1686
rect 10992 1652 11024 1686
rect 11024 1652 11026 1686
rect 10920 1579 10922 1613
rect 10922 1579 10954 1613
rect 10992 1579 11024 1613
rect 11024 1579 11026 1613
rect 10920 1506 10922 1540
rect 10922 1506 10954 1540
rect 10992 1506 11024 1540
rect 11024 1506 11026 1540
rect 10920 1432 10922 1466
rect 10922 1432 10954 1466
rect 10992 1432 11024 1466
rect 11024 1432 11026 1466
rect 10920 1358 10922 1392
rect 10922 1358 10954 1392
rect 10992 1358 11024 1392
rect 11024 1358 11026 1392
rect 10920 1284 10922 1318
rect 10922 1284 10954 1318
rect 10992 1284 11024 1318
rect 11024 1284 11026 1318
rect 10920 1210 10922 1244
rect 10922 1210 10954 1244
rect 10992 1210 11024 1244
rect 11024 1210 11026 1244
rect 10920 1136 10922 1170
rect 10922 1136 10954 1170
rect 10992 1136 11024 1170
rect 11024 1136 11026 1170
rect 10920 1062 10922 1096
rect 10922 1062 10954 1096
rect 10992 1062 11024 1096
rect 11024 1062 11026 1096
rect 10920 988 10922 1022
rect 10922 988 10954 1022
rect 10992 988 11024 1022
rect 11024 988 11026 1022
rect 10920 914 10922 948
rect 10922 914 10954 948
rect 10992 914 11024 948
rect 11024 914 11026 948
rect 10920 840 10922 874
rect 10922 840 10954 874
rect 10992 840 11024 874
rect 11024 840 11026 874
rect 10920 790 10922 800
rect 10922 790 10954 800
rect 10992 790 11024 800
rect 11024 790 11026 800
rect 10920 766 10954 790
rect 10992 766 11026 790
rect 10920 721 10922 726
rect 10922 721 10954 726
rect 10992 721 11024 726
rect 11024 721 11026 726
rect 10920 692 10954 721
rect 10992 692 11026 721
rect 10920 618 10954 652
rect 10992 618 11026 652
rect 10920 548 10954 578
rect 10992 548 11026 578
rect 10920 544 10922 548
rect 10922 544 10954 548
rect 10992 544 11024 548
rect 11024 544 11026 548
rect 10920 479 10954 504
rect 10992 479 11026 504
rect 10920 470 10922 479
rect 10922 470 10954 479
rect 10992 470 11024 479
rect 11024 470 11026 479
rect 10920 410 10954 430
rect 10992 410 11026 430
rect 10920 396 10922 410
rect 10922 396 10954 410
rect 10992 396 11024 410
rect 11024 396 11026 410
rect 10920 341 10954 356
rect 10992 341 11026 356
rect 10920 322 10922 341
rect 10922 322 10954 341
rect 10992 322 11024 341
rect 11024 322 11026 341
rect 10920 272 10954 282
rect 10992 272 11026 282
rect 10920 248 10922 272
rect 10922 248 10954 272
rect 10992 248 11024 272
rect 11024 248 11026 272
rect 10920 203 10954 208
rect 10992 203 11026 208
rect 10920 174 10922 203
rect 10922 174 10954 203
rect 10992 174 11024 203
rect 11024 174 11026 203
rect 10920 100 10922 134
rect 10922 100 10954 134
rect 10992 100 11024 134
rect 11024 100 11026 134
rect 11332 2966 11334 3000
rect 11334 2966 11366 3000
rect 11404 2966 11436 3000
rect 11436 2966 11438 3000
rect 11332 2893 11334 2927
rect 11334 2893 11366 2927
rect 11404 2893 11436 2927
rect 11436 2893 11438 2927
rect 11332 2820 11334 2854
rect 11334 2820 11366 2854
rect 11404 2820 11436 2854
rect 11436 2820 11438 2854
rect 11332 2747 11334 2781
rect 11334 2747 11366 2781
rect 11404 2747 11436 2781
rect 11436 2747 11438 2781
rect 11332 2674 11334 2708
rect 11334 2674 11366 2708
rect 11404 2674 11436 2708
rect 11436 2674 11438 2708
rect 11332 2601 11334 2635
rect 11334 2601 11366 2635
rect 11404 2601 11436 2635
rect 11436 2601 11438 2635
rect 11332 2528 11334 2562
rect 11334 2528 11366 2562
rect 11404 2528 11436 2562
rect 11436 2528 11438 2562
rect 11332 2455 11334 2489
rect 11334 2455 11366 2489
rect 11404 2455 11436 2489
rect 11436 2455 11438 2489
rect 11332 2382 11334 2416
rect 11334 2382 11366 2416
rect 11404 2382 11436 2416
rect 11436 2382 11438 2416
rect 11332 2309 11334 2343
rect 11334 2309 11366 2343
rect 11404 2309 11436 2343
rect 11436 2309 11438 2343
rect 11332 2236 11334 2270
rect 11334 2236 11366 2270
rect 11404 2236 11436 2270
rect 11436 2236 11438 2270
rect 11332 2163 11334 2197
rect 11334 2163 11366 2197
rect 11404 2163 11436 2197
rect 11436 2163 11438 2197
rect 11332 2090 11334 2124
rect 11334 2090 11366 2124
rect 11404 2090 11436 2124
rect 11436 2090 11438 2124
rect 11332 2017 11334 2051
rect 11334 2017 11366 2051
rect 11404 2017 11436 2051
rect 11436 2017 11438 2051
rect 11332 1944 11334 1978
rect 11334 1944 11366 1978
rect 11404 1944 11436 1978
rect 11436 1944 11438 1978
rect 11332 1871 11334 1905
rect 11334 1871 11366 1905
rect 11404 1871 11436 1905
rect 11436 1871 11438 1905
rect 11332 1798 11334 1832
rect 11334 1798 11366 1832
rect 11404 1798 11436 1832
rect 11436 1798 11438 1832
rect 11332 1725 11334 1759
rect 11334 1725 11366 1759
rect 11404 1725 11436 1759
rect 11436 1725 11438 1759
rect 11332 1652 11334 1686
rect 11334 1652 11366 1686
rect 11404 1652 11436 1686
rect 11436 1652 11438 1686
rect 11332 1579 11334 1613
rect 11334 1579 11366 1613
rect 11404 1579 11436 1613
rect 11436 1579 11438 1613
rect 11332 1506 11334 1540
rect 11334 1506 11366 1540
rect 11404 1506 11436 1540
rect 11436 1506 11438 1540
rect 11332 1432 11334 1466
rect 11334 1432 11366 1466
rect 11404 1432 11436 1466
rect 11436 1432 11438 1466
rect 11332 1358 11334 1392
rect 11334 1358 11366 1392
rect 11404 1358 11436 1392
rect 11436 1358 11438 1392
rect 11332 1284 11334 1318
rect 11334 1284 11366 1318
rect 11404 1284 11436 1318
rect 11436 1284 11438 1318
rect 11332 1210 11334 1244
rect 11334 1210 11366 1244
rect 11404 1210 11436 1244
rect 11436 1210 11438 1244
rect 11332 1136 11334 1170
rect 11334 1136 11366 1170
rect 11404 1136 11436 1170
rect 11436 1136 11438 1170
rect 11332 1062 11334 1096
rect 11334 1062 11366 1096
rect 11404 1062 11436 1096
rect 11436 1062 11438 1096
rect 11332 988 11334 1022
rect 11334 988 11366 1022
rect 11404 988 11436 1022
rect 11436 988 11438 1022
rect 11332 914 11334 948
rect 11334 914 11366 948
rect 11404 914 11436 948
rect 11436 914 11438 948
rect 11332 840 11334 874
rect 11334 840 11366 874
rect 11404 840 11436 874
rect 11436 840 11438 874
rect 11332 790 11334 800
rect 11334 790 11366 800
rect 11404 790 11436 800
rect 11436 790 11438 800
rect 11332 766 11366 790
rect 11404 766 11438 790
rect 11332 721 11334 726
rect 11334 721 11366 726
rect 11404 721 11436 726
rect 11436 721 11438 726
rect 11332 692 11366 721
rect 11404 692 11438 721
rect 11332 618 11366 652
rect 11404 618 11438 652
rect 11332 548 11366 578
rect 11404 548 11438 578
rect 11332 544 11334 548
rect 11334 544 11366 548
rect 11404 544 11436 548
rect 11436 544 11438 548
rect 11332 479 11366 504
rect 11404 479 11438 504
rect 11332 470 11334 479
rect 11334 470 11366 479
rect 11404 470 11436 479
rect 11436 470 11438 479
rect 11332 410 11366 430
rect 11404 410 11438 430
rect 11332 396 11334 410
rect 11334 396 11366 410
rect 11404 396 11436 410
rect 11436 396 11438 410
rect 11332 341 11366 356
rect 11404 341 11438 356
rect 11332 322 11334 341
rect 11334 322 11366 341
rect 11404 322 11436 341
rect 11436 322 11438 341
rect 11332 272 11366 282
rect 11404 272 11438 282
rect 11332 248 11334 272
rect 11334 248 11366 272
rect 11404 248 11436 272
rect 11436 248 11438 272
rect 11332 203 11366 208
rect 11404 203 11438 208
rect 11332 174 11334 203
rect 11334 174 11366 203
rect 11404 174 11436 203
rect 11436 174 11438 203
rect 11332 100 11334 134
rect 11334 100 11366 134
rect 11404 100 11436 134
rect 11436 100 11438 134
rect 11744 2966 11746 3000
rect 11746 2966 11778 3000
rect 11816 2966 11848 3000
rect 11848 2966 11850 3000
rect 11744 2893 11746 2927
rect 11746 2893 11778 2927
rect 11816 2893 11848 2927
rect 11848 2893 11850 2927
rect 11744 2820 11746 2854
rect 11746 2820 11778 2854
rect 11816 2820 11848 2854
rect 11848 2820 11850 2854
rect 11744 2747 11746 2781
rect 11746 2747 11778 2781
rect 11816 2747 11848 2781
rect 11848 2747 11850 2781
rect 11744 2674 11746 2708
rect 11746 2674 11778 2708
rect 11816 2674 11848 2708
rect 11848 2674 11850 2708
rect 11744 2601 11746 2635
rect 11746 2601 11778 2635
rect 11816 2601 11848 2635
rect 11848 2601 11850 2635
rect 11744 2528 11746 2562
rect 11746 2528 11778 2562
rect 11816 2528 11848 2562
rect 11848 2528 11850 2562
rect 11744 2455 11746 2489
rect 11746 2455 11778 2489
rect 11816 2455 11848 2489
rect 11848 2455 11850 2489
rect 11744 2382 11746 2416
rect 11746 2382 11778 2416
rect 11816 2382 11848 2416
rect 11848 2382 11850 2416
rect 11744 2309 11746 2343
rect 11746 2309 11778 2343
rect 11816 2309 11848 2343
rect 11848 2309 11850 2343
rect 11744 2236 11746 2270
rect 11746 2236 11778 2270
rect 11816 2236 11848 2270
rect 11848 2236 11850 2270
rect 11744 2163 11746 2197
rect 11746 2163 11778 2197
rect 11816 2163 11848 2197
rect 11848 2163 11850 2197
rect 11744 2090 11746 2124
rect 11746 2090 11778 2124
rect 11816 2090 11848 2124
rect 11848 2090 11850 2124
rect 11744 2017 11746 2051
rect 11746 2017 11778 2051
rect 11816 2017 11848 2051
rect 11848 2017 11850 2051
rect 11744 1944 11746 1978
rect 11746 1944 11778 1978
rect 11816 1944 11848 1978
rect 11848 1944 11850 1978
rect 11744 1871 11746 1905
rect 11746 1871 11778 1905
rect 11816 1871 11848 1905
rect 11848 1871 11850 1905
rect 11744 1798 11746 1832
rect 11746 1798 11778 1832
rect 11816 1798 11848 1832
rect 11848 1798 11850 1832
rect 11744 1725 11746 1759
rect 11746 1725 11778 1759
rect 11816 1725 11848 1759
rect 11848 1725 11850 1759
rect 11744 1652 11746 1686
rect 11746 1652 11778 1686
rect 11816 1652 11848 1686
rect 11848 1652 11850 1686
rect 11744 1579 11746 1613
rect 11746 1579 11778 1613
rect 11816 1579 11848 1613
rect 11848 1579 11850 1613
rect 11744 1506 11746 1540
rect 11746 1506 11778 1540
rect 11816 1506 11848 1540
rect 11848 1506 11850 1540
rect 11744 1432 11746 1466
rect 11746 1432 11778 1466
rect 11816 1432 11848 1466
rect 11848 1432 11850 1466
rect 11744 1358 11746 1392
rect 11746 1358 11778 1392
rect 11816 1358 11848 1392
rect 11848 1358 11850 1392
rect 11744 1284 11746 1318
rect 11746 1284 11778 1318
rect 11816 1284 11848 1318
rect 11848 1284 11850 1318
rect 11744 1210 11746 1244
rect 11746 1210 11778 1244
rect 11816 1210 11848 1244
rect 11848 1210 11850 1244
rect 11744 1136 11746 1170
rect 11746 1136 11778 1170
rect 11816 1136 11848 1170
rect 11848 1136 11850 1170
rect 11744 1062 11746 1096
rect 11746 1062 11778 1096
rect 11816 1062 11848 1096
rect 11848 1062 11850 1096
rect 11744 988 11746 1022
rect 11746 988 11778 1022
rect 11816 988 11848 1022
rect 11848 988 11850 1022
rect 11744 914 11746 948
rect 11746 914 11778 948
rect 11816 914 11848 948
rect 11848 914 11850 948
rect 11744 840 11746 874
rect 11746 840 11778 874
rect 11816 840 11848 874
rect 11848 840 11850 874
rect 11744 790 11746 800
rect 11746 790 11778 800
rect 11816 790 11848 800
rect 11848 790 11850 800
rect 11744 766 11778 790
rect 11816 766 11850 790
rect 11744 721 11746 726
rect 11746 721 11778 726
rect 11816 721 11848 726
rect 11848 721 11850 726
rect 11744 692 11778 721
rect 11816 692 11850 721
rect 11744 618 11778 652
rect 11816 618 11850 652
rect 11744 548 11778 578
rect 11816 548 11850 578
rect 11744 544 11746 548
rect 11746 544 11778 548
rect 11816 544 11848 548
rect 11848 544 11850 548
rect 11744 479 11778 504
rect 11816 479 11850 504
rect 11744 470 11746 479
rect 11746 470 11778 479
rect 11816 470 11848 479
rect 11848 470 11850 479
rect 11744 410 11778 430
rect 11816 410 11850 430
rect 11744 396 11746 410
rect 11746 396 11778 410
rect 11816 396 11848 410
rect 11848 396 11850 410
rect 11744 341 11778 356
rect 11816 341 11850 356
rect 11744 322 11746 341
rect 11746 322 11778 341
rect 11816 322 11848 341
rect 11848 322 11850 341
rect 11744 272 11778 282
rect 11816 272 11850 282
rect 11744 248 11746 272
rect 11746 248 11778 272
rect 11816 248 11848 272
rect 11848 248 11850 272
rect 11744 203 11778 208
rect 11816 203 11850 208
rect 11744 174 11746 203
rect 11746 174 11778 203
rect 11816 174 11848 203
rect 11848 174 11850 203
rect 11744 100 11746 134
rect 11746 100 11778 134
rect 11816 100 11848 134
rect 11848 100 11850 134
rect 12156 2966 12158 3000
rect 12158 2966 12190 3000
rect 12228 2966 12260 3000
rect 12260 2966 12262 3000
rect 12156 2893 12158 2927
rect 12158 2893 12190 2927
rect 12228 2893 12260 2927
rect 12260 2893 12262 2927
rect 12156 2820 12158 2854
rect 12158 2820 12190 2854
rect 12228 2820 12260 2854
rect 12260 2820 12262 2854
rect 12156 2747 12158 2781
rect 12158 2747 12190 2781
rect 12228 2747 12260 2781
rect 12260 2747 12262 2781
rect 12156 2674 12158 2708
rect 12158 2674 12190 2708
rect 12228 2674 12260 2708
rect 12260 2674 12262 2708
rect 12156 2601 12158 2635
rect 12158 2601 12190 2635
rect 12228 2601 12260 2635
rect 12260 2601 12262 2635
rect 12156 2528 12158 2562
rect 12158 2528 12190 2562
rect 12228 2528 12260 2562
rect 12260 2528 12262 2562
rect 12156 2455 12158 2489
rect 12158 2455 12190 2489
rect 12228 2455 12260 2489
rect 12260 2455 12262 2489
rect 12156 2382 12158 2416
rect 12158 2382 12190 2416
rect 12228 2382 12260 2416
rect 12260 2382 12262 2416
rect 12156 2309 12158 2343
rect 12158 2309 12190 2343
rect 12228 2309 12260 2343
rect 12260 2309 12262 2343
rect 12156 2236 12158 2270
rect 12158 2236 12190 2270
rect 12228 2236 12260 2270
rect 12260 2236 12262 2270
rect 12156 2163 12158 2197
rect 12158 2163 12190 2197
rect 12228 2163 12260 2197
rect 12260 2163 12262 2197
rect 12156 2090 12158 2124
rect 12158 2090 12190 2124
rect 12228 2090 12260 2124
rect 12260 2090 12262 2124
rect 12156 2017 12158 2051
rect 12158 2017 12190 2051
rect 12228 2017 12260 2051
rect 12260 2017 12262 2051
rect 12156 1944 12158 1978
rect 12158 1944 12190 1978
rect 12228 1944 12260 1978
rect 12260 1944 12262 1978
rect 12156 1871 12158 1905
rect 12158 1871 12190 1905
rect 12228 1871 12260 1905
rect 12260 1871 12262 1905
rect 12156 1798 12158 1832
rect 12158 1798 12190 1832
rect 12228 1798 12260 1832
rect 12260 1798 12262 1832
rect 12156 1725 12158 1759
rect 12158 1725 12190 1759
rect 12228 1725 12260 1759
rect 12260 1725 12262 1759
rect 12156 1652 12158 1686
rect 12158 1652 12190 1686
rect 12228 1652 12260 1686
rect 12260 1652 12262 1686
rect 12156 1579 12158 1613
rect 12158 1579 12190 1613
rect 12228 1579 12260 1613
rect 12260 1579 12262 1613
rect 12156 1506 12158 1540
rect 12158 1506 12190 1540
rect 12228 1506 12260 1540
rect 12260 1506 12262 1540
rect 12156 1432 12158 1466
rect 12158 1432 12190 1466
rect 12228 1432 12260 1466
rect 12260 1432 12262 1466
rect 12156 1358 12158 1392
rect 12158 1358 12190 1392
rect 12228 1358 12260 1392
rect 12260 1358 12262 1392
rect 12156 1284 12158 1318
rect 12158 1284 12190 1318
rect 12228 1284 12260 1318
rect 12260 1284 12262 1318
rect 12156 1210 12158 1244
rect 12158 1210 12190 1244
rect 12228 1210 12260 1244
rect 12260 1210 12262 1244
rect 12156 1136 12158 1170
rect 12158 1136 12190 1170
rect 12228 1136 12260 1170
rect 12260 1136 12262 1170
rect 12156 1062 12158 1096
rect 12158 1062 12190 1096
rect 12228 1062 12260 1096
rect 12260 1062 12262 1096
rect 12156 988 12158 1022
rect 12158 988 12190 1022
rect 12228 988 12260 1022
rect 12260 988 12262 1022
rect 12156 914 12158 948
rect 12158 914 12190 948
rect 12228 914 12260 948
rect 12260 914 12262 948
rect 12156 840 12158 874
rect 12158 840 12190 874
rect 12228 840 12260 874
rect 12260 840 12262 874
rect 12156 790 12158 800
rect 12158 790 12190 800
rect 12228 790 12260 800
rect 12260 790 12262 800
rect 12156 766 12190 790
rect 12228 766 12262 790
rect 12156 721 12158 726
rect 12158 721 12190 726
rect 12228 721 12260 726
rect 12260 721 12262 726
rect 12156 692 12190 721
rect 12228 692 12262 721
rect 12156 618 12190 652
rect 12228 618 12262 652
rect 12156 548 12190 578
rect 12228 548 12262 578
rect 12156 544 12158 548
rect 12158 544 12190 548
rect 12228 544 12260 548
rect 12260 544 12262 548
rect 12156 479 12190 504
rect 12228 479 12262 504
rect 12156 470 12158 479
rect 12158 470 12190 479
rect 12228 470 12260 479
rect 12260 470 12262 479
rect 12156 410 12190 430
rect 12228 410 12262 430
rect 12156 396 12158 410
rect 12158 396 12190 410
rect 12228 396 12260 410
rect 12260 396 12262 410
rect 12156 341 12190 356
rect 12228 341 12262 356
rect 12156 322 12158 341
rect 12158 322 12190 341
rect 12228 322 12260 341
rect 12260 322 12262 341
rect 12156 272 12190 282
rect 12228 272 12262 282
rect 12156 248 12158 272
rect 12158 248 12190 272
rect 12228 248 12260 272
rect 12260 248 12262 272
rect 12156 203 12190 208
rect 12228 203 12262 208
rect 12156 174 12158 203
rect 12158 174 12190 203
rect 12228 174 12260 203
rect 12260 174 12262 203
rect 12156 100 12158 134
rect 12158 100 12190 134
rect 12228 100 12260 134
rect 12260 100 12262 134
rect 12568 2966 12570 3000
rect 12570 2966 12602 3000
rect 12640 2966 12672 3000
rect 12672 2966 12674 3000
rect 12568 2893 12570 2927
rect 12570 2893 12602 2927
rect 12640 2893 12672 2927
rect 12672 2893 12674 2927
rect 12568 2820 12570 2854
rect 12570 2820 12602 2854
rect 12640 2820 12672 2854
rect 12672 2820 12674 2854
rect 12568 2747 12570 2781
rect 12570 2747 12602 2781
rect 12640 2747 12672 2781
rect 12672 2747 12674 2781
rect 12568 2674 12570 2708
rect 12570 2674 12602 2708
rect 12640 2674 12672 2708
rect 12672 2674 12674 2708
rect 12568 2601 12570 2635
rect 12570 2601 12602 2635
rect 12640 2601 12672 2635
rect 12672 2601 12674 2635
rect 12568 2528 12570 2562
rect 12570 2528 12602 2562
rect 12640 2528 12672 2562
rect 12672 2528 12674 2562
rect 12568 2455 12570 2489
rect 12570 2455 12602 2489
rect 12640 2455 12672 2489
rect 12672 2455 12674 2489
rect 12568 2382 12570 2416
rect 12570 2382 12602 2416
rect 12640 2382 12672 2416
rect 12672 2382 12674 2416
rect 12568 2309 12570 2343
rect 12570 2309 12602 2343
rect 12640 2309 12672 2343
rect 12672 2309 12674 2343
rect 12568 2236 12570 2270
rect 12570 2236 12602 2270
rect 12640 2236 12672 2270
rect 12672 2236 12674 2270
rect 12568 2163 12570 2197
rect 12570 2163 12602 2197
rect 12640 2163 12672 2197
rect 12672 2163 12674 2197
rect 12568 2090 12570 2124
rect 12570 2090 12602 2124
rect 12640 2090 12672 2124
rect 12672 2090 12674 2124
rect 12568 2017 12570 2051
rect 12570 2017 12602 2051
rect 12640 2017 12672 2051
rect 12672 2017 12674 2051
rect 12568 1944 12570 1978
rect 12570 1944 12602 1978
rect 12640 1944 12672 1978
rect 12672 1944 12674 1978
rect 12568 1871 12570 1905
rect 12570 1871 12602 1905
rect 12640 1871 12672 1905
rect 12672 1871 12674 1905
rect 12568 1798 12570 1832
rect 12570 1798 12602 1832
rect 12640 1798 12672 1832
rect 12672 1798 12674 1832
rect 12568 1725 12570 1759
rect 12570 1725 12602 1759
rect 12640 1725 12672 1759
rect 12672 1725 12674 1759
rect 12568 1652 12570 1686
rect 12570 1652 12602 1686
rect 12640 1652 12672 1686
rect 12672 1652 12674 1686
rect 12568 1579 12570 1613
rect 12570 1579 12602 1613
rect 12640 1579 12672 1613
rect 12672 1579 12674 1613
rect 12568 1506 12570 1540
rect 12570 1506 12602 1540
rect 12640 1506 12672 1540
rect 12672 1506 12674 1540
rect 12568 1432 12570 1466
rect 12570 1432 12602 1466
rect 12640 1432 12672 1466
rect 12672 1432 12674 1466
rect 12568 1358 12570 1392
rect 12570 1358 12602 1392
rect 12640 1358 12672 1392
rect 12672 1358 12674 1392
rect 12568 1284 12570 1318
rect 12570 1284 12602 1318
rect 12640 1284 12672 1318
rect 12672 1284 12674 1318
rect 12568 1210 12570 1244
rect 12570 1210 12602 1244
rect 12640 1210 12672 1244
rect 12672 1210 12674 1244
rect 12568 1136 12570 1170
rect 12570 1136 12602 1170
rect 12640 1136 12672 1170
rect 12672 1136 12674 1170
rect 12568 1062 12570 1096
rect 12570 1062 12602 1096
rect 12640 1062 12672 1096
rect 12672 1062 12674 1096
rect 12568 988 12570 1022
rect 12570 988 12602 1022
rect 12640 988 12672 1022
rect 12672 988 12674 1022
rect 12568 914 12570 948
rect 12570 914 12602 948
rect 12640 914 12672 948
rect 12672 914 12674 948
rect 12568 840 12570 874
rect 12570 840 12602 874
rect 12640 840 12672 874
rect 12672 840 12674 874
rect 12568 790 12570 800
rect 12570 790 12602 800
rect 12640 790 12672 800
rect 12672 790 12674 800
rect 12568 766 12602 790
rect 12640 766 12674 790
rect 12568 721 12570 726
rect 12570 721 12602 726
rect 12640 721 12672 726
rect 12672 721 12674 726
rect 12568 692 12602 721
rect 12640 692 12674 721
rect 12568 618 12602 652
rect 12640 618 12674 652
rect 12568 548 12602 578
rect 12640 548 12674 578
rect 12568 544 12570 548
rect 12570 544 12602 548
rect 12640 544 12672 548
rect 12672 544 12674 548
rect 12568 479 12602 504
rect 12640 479 12674 504
rect 12568 470 12570 479
rect 12570 470 12602 479
rect 12640 470 12672 479
rect 12672 470 12674 479
rect 12568 410 12602 430
rect 12640 410 12674 430
rect 12568 396 12570 410
rect 12570 396 12602 410
rect 12640 396 12672 410
rect 12672 396 12674 410
rect 12568 341 12602 356
rect 12640 341 12674 356
rect 12568 322 12570 341
rect 12570 322 12602 341
rect 12640 322 12672 341
rect 12672 322 12674 341
rect 12568 272 12602 282
rect 12640 272 12674 282
rect 12568 248 12570 272
rect 12570 248 12602 272
rect 12640 248 12672 272
rect 12672 248 12674 272
rect 12568 203 12602 208
rect 12640 203 12674 208
rect 12568 174 12570 203
rect 12570 174 12602 203
rect 12640 174 12672 203
rect 12672 174 12674 203
rect 12568 100 12570 134
rect 12570 100 12602 134
rect 12640 100 12672 134
rect 12672 100 12674 134
rect 12980 2966 12982 3000
rect 12982 2966 13014 3000
rect 13052 2966 13084 3000
rect 13084 2966 13086 3000
rect 12980 2893 12982 2927
rect 12982 2893 13014 2927
rect 13052 2893 13084 2927
rect 13084 2893 13086 2927
rect 12980 2820 12982 2854
rect 12982 2820 13014 2854
rect 13052 2820 13084 2854
rect 13084 2820 13086 2854
rect 12980 2747 12982 2781
rect 12982 2747 13014 2781
rect 13052 2747 13084 2781
rect 13084 2747 13086 2781
rect 12980 2674 12982 2708
rect 12982 2674 13014 2708
rect 13052 2674 13084 2708
rect 13084 2674 13086 2708
rect 12980 2601 12982 2635
rect 12982 2601 13014 2635
rect 13052 2601 13084 2635
rect 13084 2601 13086 2635
rect 12980 2528 12982 2562
rect 12982 2528 13014 2562
rect 13052 2528 13084 2562
rect 13084 2528 13086 2562
rect 12980 2455 12982 2489
rect 12982 2455 13014 2489
rect 13052 2455 13084 2489
rect 13084 2455 13086 2489
rect 12980 2382 12982 2416
rect 12982 2382 13014 2416
rect 13052 2382 13084 2416
rect 13084 2382 13086 2416
rect 12980 2309 12982 2343
rect 12982 2309 13014 2343
rect 13052 2309 13084 2343
rect 13084 2309 13086 2343
rect 12980 2236 12982 2270
rect 12982 2236 13014 2270
rect 13052 2236 13084 2270
rect 13084 2236 13086 2270
rect 12980 2163 12982 2197
rect 12982 2163 13014 2197
rect 13052 2163 13084 2197
rect 13084 2163 13086 2197
rect 12980 2090 12982 2124
rect 12982 2090 13014 2124
rect 13052 2090 13084 2124
rect 13084 2090 13086 2124
rect 12980 2017 12982 2051
rect 12982 2017 13014 2051
rect 13052 2017 13084 2051
rect 13084 2017 13086 2051
rect 12980 1944 12982 1978
rect 12982 1944 13014 1978
rect 13052 1944 13084 1978
rect 13084 1944 13086 1978
rect 12980 1871 12982 1905
rect 12982 1871 13014 1905
rect 13052 1871 13084 1905
rect 13084 1871 13086 1905
rect 12980 1798 12982 1832
rect 12982 1798 13014 1832
rect 13052 1798 13084 1832
rect 13084 1798 13086 1832
rect 12980 1725 12982 1759
rect 12982 1725 13014 1759
rect 13052 1725 13084 1759
rect 13084 1725 13086 1759
rect 12980 1652 12982 1686
rect 12982 1652 13014 1686
rect 13052 1652 13084 1686
rect 13084 1652 13086 1686
rect 12980 1579 12982 1613
rect 12982 1579 13014 1613
rect 13052 1579 13084 1613
rect 13084 1579 13086 1613
rect 12980 1506 12982 1540
rect 12982 1506 13014 1540
rect 13052 1506 13084 1540
rect 13084 1506 13086 1540
rect 12980 1432 12982 1466
rect 12982 1432 13014 1466
rect 13052 1432 13084 1466
rect 13084 1432 13086 1466
rect 12980 1358 12982 1392
rect 12982 1358 13014 1392
rect 13052 1358 13084 1392
rect 13084 1358 13086 1392
rect 12980 1284 12982 1318
rect 12982 1284 13014 1318
rect 13052 1284 13084 1318
rect 13084 1284 13086 1318
rect 12980 1210 12982 1244
rect 12982 1210 13014 1244
rect 13052 1210 13084 1244
rect 13084 1210 13086 1244
rect 12980 1136 12982 1170
rect 12982 1136 13014 1170
rect 13052 1136 13084 1170
rect 13084 1136 13086 1170
rect 12980 1062 12982 1096
rect 12982 1062 13014 1096
rect 13052 1062 13084 1096
rect 13084 1062 13086 1096
rect 12980 988 12982 1022
rect 12982 988 13014 1022
rect 13052 988 13084 1022
rect 13084 988 13086 1022
rect 12980 914 12982 948
rect 12982 914 13014 948
rect 13052 914 13084 948
rect 13084 914 13086 948
rect 12980 840 12982 874
rect 12982 840 13014 874
rect 13052 840 13084 874
rect 13084 840 13086 874
rect 12980 790 12982 800
rect 12982 790 13014 800
rect 13052 790 13084 800
rect 13084 790 13086 800
rect 12980 766 13014 790
rect 13052 766 13086 790
rect 12980 721 12982 726
rect 12982 721 13014 726
rect 13052 721 13084 726
rect 13084 721 13086 726
rect 12980 692 13014 721
rect 13052 692 13086 721
rect 12980 618 13014 652
rect 13052 618 13086 652
rect 12980 548 13014 578
rect 13052 548 13086 578
rect 12980 544 12982 548
rect 12982 544 13014 548
rect 13052 544 13084 548
rect 13084 544 13086 548
rect 12980 479 13014 504
rect 13052 479 13086 504
rect 12980 470 12982 479
rect 12982 470 13014 479
rect 13052 470 13084 479
rect 13084 470 13086 479
rect 12980 410 13014 430
rect 13052 410 13086 430
rect 12980 396 12982 410
rect 12982 396 13014 410
rect 13052 396 13084 410
rect 13084 396 13086 410
rect 12980 341 13014 356
rect 13052 341 13086 356
rect 12980 322 12982 341
rect 12982 322 13014 341
rect 13052 322 13084 341
rect 13084 322 13086 341
rect 12980 272 13014 282
rect 13052 272 13086 282
rect 12980 248 12982 272
rect 12982 248 13014 272
rect 13052 248 13084 272
rect 13084 248 13086 272
rect 12980 203 13014 208
rect 13052 203 13086 208
rect 12980 174 12982 203
rect 12982 174 13014 203
rect 13052 174 13084 203
rect 13084 174 13086 203
rect 12980 100 12982 134
rect 12982 100 13014 134
rect 13052 100 13084 134
rect 13084 100 13086 134
rect 13202 2451 13956 3277
rect 13202 2378 13236 2412
rect 13274 2378 13308 2412
rect 13346 2378 13380 2412
rect 13418 2378 13452 2412
rect 13490 2378 13524 2412
rect 13562 2378 13596 2412
rect 13634 2378 13668 2412
rect 13706 2378 13740 2412
rect 13778 2378 13812 2412
rect 13850 2378 13884 2412
rect 13922 2378 13956 2412
rect 13202 2305 13236 2339
rect 13274 2305 13308 2339
rect 13346 2305 13380 2339
rect 13418 2305 13452 2339
rect 13490 2305 13524 2339
rect 13562 2305 13596 2339
rect 13634 2305 13668 2339
rect 13706 2305 13740 2339
rect 13778 2305 13812 2339
rect 13850 2305 13884 2339
rect 13922 2305 13956 2339
rect 13202 2232 13236 2266
rect 13274 2232 13308 2266
rect 13346 2232 13380 2266
rect 13418 2232 13452 2266
rect 13490 2232 13524 2266
rect 13562 2232 13596 2266
rect 13634 2232 13668 2266
rect 13706 2232 13740 2266
rect 13778 2232 13812 2266
rect 13850 2232 13884 2266
rect 13922 2232 13956 2266
rect 13202 2159 13236 2193
rect 13274 2159 13308 2193
rect 13346 2159 13380 2193
rect 13418 2159 13452 2193
rect 13490 2159 13524 2193
rect 13562 2159 13596 2193
rect 13634 2159 13668 2193
rect 13706 2159 13740 2193
rect 13778 2159 13812 2193
rect 13850 2159 13884 2193
rect 13922 2159 13956 2193
rect 13202 2086 13236 2120
rect 13274 2086 13308 2120
rect 13346 2086 13380 2120
rect 13418 2086 13452 2120
rect 13490 2086 13524 2120
rect 13562 2086 13596 2120
rect 13634 2086 13668 2120
rect 13706 2086 13740 2120
rect 13778 2086 13812 2120
rect 13850 2086 13884 2120
rect 13922 2086 13956 2120
rect 13202 2013 13236 2047
rect 13274 2013 13308 2047
rect 13346 2013 13380 2047
rect 13418 2013 13452 2047
rect 13490 2013 13524 2047
rect 13562 2013 13596 2047
rect 13634 2013 13668 2047
rect 13706 2013 13740 2047
rect 13778 2013 13812 2047
rect 13850 2013 13884 2047
rect 13922 2013 13956 2047
rect 13202 1940 13236 1974
rect 13274 1940 13308 1974
rect 13346 1940 13380 1974
rect 13418 1940 13452 1974
rect 13490 1940 13524 1974
rect 13562 1940 13596 1974
rect 13634 1940 13668 1974
rect 13706 1940 13740 1974
rect 13778 1940 13812 1974
rect 13850 1940 13884 1974
rect 13922 1940 13956 1974
rect 13202 1867 13236 1901
rect 13274 1867 13308 1901
rect 13346 1867 13380 1901
rect 13418 1867 13452 1901
rect 13490 1867 13524 1901
rect 13562 1867 13596 1901
rect 13634 1867 13668 1901
rect 13706 1867 13740 1901
rect 13778 1867 13812 1901
rect 13850 1867 13884 1901
rect 13922 1867 13956 1901
rect 13202 1794 13236 1828
rect 13274 1794 13308 1828
rect 13346 1794 13380 1828
rect 13418 1794 13452 1828
rect 13490 1794 13524 1828
rect 13562 1794 13596 1828
rect 13634 1794 13668 1828
rect 13706 1794 13740 1828
rect 13778 1794 13812 1828
rect 13850 1794 13884 1828
rect 13922 1794 13956 1828
rect 13202 1721 13236 1755
rect 13274 1721 13308 1755
rect 13346 1721 13380 1755
rect 13418 1721 13452 1755
rect 13490 1721 13524 1755
rect 13562 1721 13596 1755
rect 13634 1721 13668 1755
rect 13706 1721 13740 1755
rect 13778 1721 13812 1755
rect 13850 1721 13884 1755
rect 13922 1721 13956 1755
rect 13202 1648 13236 1682
rect 13274 1648 13308 1682
rect 13346 1648 13380 1682
rect 13418 1648 13452 1682
rect 13490 1648 13524 1682
rect 13562 1648 13596 1682
rect 13634 1648 13668 1682
rect 13706 1648 13740 1682
rect 13778 1648 13812 1682
rect 13850 1648 13884 1682
rect 13922 1648 13956 1682
rect 13202 1575 13236 1609
rect 13274 1575 13308 1609
rect 13346 1575 13380 1609
rect 13418 1575 13452 1609
rect 13490 1575 13524 1609
rect 13562 1575 13596 1609
rect 13634 1575 13668 1609
rect 13706 1575 13740 1609
rect 13778 1575 13812 1609
rect 13850 1575 13884 1609
rect 13922 1575 13956 1609
rect 13202 1502 13236 1536
rect 13274 1502 13308 1536
rect 13346 1502 13380 1536
rect 13418 1502 13452 1536
rect 13490 1502 13524 1536
rect 13562 1502 13596 1536
rect 13634 1502 13668 1536
rect 13706 1502 13740 1536
rect 13778 1502 13812 1536
rect 13850 1502 13884 1536
rect 13922 1502 13956 1536
rect 13202 1429 13236 1463
rect 13274 1429 13308 1463
rect 13346 1429 13380 1463
rect 13418 1429 13452 1463
rect 13490 1429 13524 1463
rect 13562 1429 13596 1463
rect 13634 1429 13668 1463
rect 13706 1429 13740 1463
rect 13778 1429 13812 1463
rect 13850 1429 13884 1463
rect 13922 1429 13956 1463
rect 13202 1356 13236 1390
rect 13274 1356 13308 1390
rect 13346 1356 13380 1390
rect 13418 1356 13452 1390
rect 13490 1356 13524 1390
rect 13562 1356 13596 1390
rect 13634 1356 13668 1390
rect 13706 1356 13740 1390
rect 13778 1356 13812 1390
rect 13850 1356 13884 1390
rect 13922 1356 13956 1390
rect 13202 1283 13236 1317
rect 13274 1283 13308 1317
rect 13346 1283 13380 1317
rect 13418 1283 13452 1317
rect 13490 1283 13524 1317
rect 13562 1283 13596 1317
rect 13634 1283 13668 1317
rect 13706 1283 13740 1317
rect 13778 1283 13812 1317
rect 13850 1283 13884 1317
rect 13922 1283 13956 1317
rect 13202 1210 13236 1244
rect 13274 1210 13308 1244
rect 13346 1210 13380 1244
rect 13418 1210 13452 1244
rect 13490 1210 13524 1244
rect 13562 1210 13596 1244
rect 13634 1210 13668 1244
rect 13706 1210 13740 1244
rect 13778 1210 13812 1244
rect 13850 1210 13884 1244
rect 13922 1210 13956 1244
rect 13202 1137 13236 1171
rect 13274 1137 13308 1171
rect 13346 1137 13380 1171
rect 13418 1137 13452 1171
rect 13490 1137 13524 1171
rect 13562 1137 13596 1171
rect 13634 1137 13668 1171
rect 13706 1137 13740 1171
rect 13778 1137 13812 1171
rect 13850 1137 13884 1171
rect 13922 1137 13956 1171
rect 13202 1064 13236 1098
rect 13274 1064 13308 1098
rect 13346 1064 13380 1098
rect 13418 1064 13452 1098
rect 13490 1064 13524 1098
rect 13562 1064 13596 1098
rect 13634 1064 13668 1098
rect 13706 1064 13740 1098
rect 13778 1064 13812 1098
rect 13850 1064 13884 1098
rect 13922 1064 13956 1098
rect 13202 991 13236 1025
rect 13274 991 13308 1025
rect 13346 991 13380 1025
rect 13418 991 13452 1025
rect 13490 991 13524 1025
rect 13562 991 13596 1025
rect 13634 991 13668 1025
rect 13706 991 13740 1025
rect 13778 991 13812 1025
rect 13850 991 13884 1025
rect 13922 991 13956 1025
rect 13202 918 13236 952
rect 13274 918 13308 952
rect 13346 918 13380 952
rect 13418 918 13452 952
rect 13490 918 13524 952
rect 13562 918 13596 952
rect 13634 918 13668 952
rect 13706 918 13740 952
rect 13778 918 13812 952
rect 13850 918 13884 952
rect 13922 918 13956 952
rect 13202 845 13236 879
rect 13274 845 13308 879
rect 13346 845 13380 879
rect 13418 845 13452 879
rect 13490 845 13524 879
rect 13562 845 13596 879
rect 13634 845 13668 879
rect 13706 845 13740 879
rect 13778 845 13812 879
rect 13850 845 13884 879
rect 13922 845 13956 879
rect 13202 772 13236 806
rect 13274 772 13308 806
rect 13346 772 13380 806
rect 13418 772 13452 806
rect 13490 772 13524 806
rect 13562 772 13596 806
rect 13634 772 13668 806
rect 13706 772 13740 806
rect 13778 772 13812 806
rect 13850 772 13884 806
rect 13922 772 13956 806
rect 13202 699 13236 733
rect 13274 699 13308 733
rect 13346 699 13380 733
rect 13418 699 13452 733
rect 13490 699 13524 733
rect 13562 699 13596 733
rect 13634 699 13668 733
rect 13706 699 13740 733
rect 13778 699 13812 733
rect 13850 699 13884 733
rect 13922 699 13956 733
rect 13202 626 13236 660
rect 13274 626 13308 660
rect 13346 626 13380 660
rect 13418 626 13452 660
rect 13490 626 13524 660
rect 13562 626 13596 660
rect 13634 626 13668 660
rect 13706 626 13740 660
rect 13778 626 13812 660
rect 13850 626 13884 660
rect 13922 626 13956 660
rect 13202 553 13236 587
rect 13274 553 13308 587
rect 13346 553 13380 587
rect 13418 553 13452 587
rect 13490 553 13524 587
rect 13562 553 13596 587
rect 13634 553 13668 587
rect 13706 553 13740 587
rect 13778 553 13812 587
rect 13850 553 13884 587
rect 13922 553 13956 587
rect 13202 484 13236 514
rect 13274 484 13308 514
rect 13346 484 13380 514
rect 13418 484 13452 514
rect 13490 484 13524 514
rect 13562 484 13596 514
rect 13634 484 13668 514
rect 13706 484 13740 514
rect 13778 484 13812 514
rect 13850 484 13884 514
rect 13922 484 13956 514
rect 13202 480 13236 484
rect 13274 480 13308 484
rect 13346 480 13380 484
rect 13418 480 13452 484
rect 13490 480 13524 484
rect 13562 480 13596 484
rect 13634 480 13668 484
rect 13706 480 13740 484
rect 13778 480 13812 484
rect 13850 480 13884 484
rect 13922 480 13956 484
rect 13202 415 13222 441
rect 13222 415 13236 441
rect 13274 415 13290 441
rect 13290 415 13308 441
rect 13346 415 13358 441
rect 13358 415 13380 441
rect 13418 415 13426 441
rect 13426 415 13452 441
rect 13490 415 13494 441
rect 13494 415 13524 441
rect 13202 407 13236 415
rect 13274 407 13308 415
rect 13346 407 13380 415
rect 13418 407 13452 415
rect 13490 407 13524 415
rect 13562 407 13596 441
rect 13634 415 13664 441
rect 13664 415 13668 441
rect 13706 415 13732 441
rect 13732 415 13740 441
rect 13778 415 13800 441
rect 13800 415 13812 441
rect 13850 415 13868 441
rect 13868 415 13884 441
rect 13922 415 13936 441
rect 13936 415 13956 441
rect 13634 407 13668 415
rect 13706 407 13740 415
rect 13778 407 13812 415
rect 13850 407 13884 415
rect 13922 407 13956 415
rect 13202 346 13222 368
rect 13222 346 13236 368
rect 13274 346 13290 368
rect 13290 346 13308 368
rect 13346 346 13358 368
rect 13358 346 13380 368
rect 13418 346 13426 368
rect 13426 346 13452 368
rect 13490 346 13494 368
rect 13494 346 13524 368
rect 13202 334 13236 346
rect 13274 334 13308 346
rect 13346 334 13380 346
rect 13418 334 13452 346
rect 13490 334 13524 346
rect 13562 334 13596 368
rect 13634 346 13664 368
rect 13664 346 13668 368
rect 13706 346 13732 368
rect 13732 346 13740 368
rect 13778 346 13800 368
rect 13800 346 13812 368
rect 13850 346 13868 368
rect 13868 346 13884 368
rect 13922 346 13936 368
rect 13936 346 13956 368
rect 13634 334 13668 346
rect 13706 334 13740 346
rect 13778 334 13812 346
rect 13850 334 13884 346
rect 13922 334 13956 346
rect 13202 277 13222 295
rect 13222 277 13236 295
rect 13274 277 13290 295
rect 13290 277 13308 295
rect 13346 277 13358 295
rect 13358 277 13380 295
rect 13418 277 13426 295
rect 13426 277 13452 295
rect 13490 277 13494 295
rect 13494 277 13524 295
rect 13202 261 13236 277
rect 13274 261 13308 277
rect 13346 261 13380 277
rect 13418 261 13452 277
rect 13490 261 13524 277
rect 13562 261 13596 295
rect 13634 277 13664 295
rect 13664 277 13668 295
rect 13706 277 13732 295
rect 13732 277 13740 295
rect 13778 277 13800 295
rect 13800 277 13812 295
rect 13850 277 13868 295
rect 13868 277 13884 295
rect 13922 277 13936 295
rect 13936 277 13956 295
rect 13634 261 13668 277
rect 13706 261 13740 277
rect 13778 261 13812 277
rect 13850 261 13884 277
rect 13922 261 13956 277
rect 13202 208 13222 222
rect 13222 208 13236 222
rect 13274 208 13290 222
rect 13290 208 13308 222
rect 13346 208 13358 222
rect 13358 208 13380 222
rect 13418 208 13426 222
rect 13426 208 13452 222
rect 13490 208 13494 222
rect 13494 208 13524 222
rect 13202 188 13236 208
rect 13274 188 13308 208
rect 13346 188 13380 208
rect 13418 188 13452 208
rect 13490 188 13524 208
rect 13562 188 13596 222
rect 13634 208 13664 222
rect 13664 208 13668 222
rect 13706 208 13732 222
rect 13732 208 13740 222
rect 13778 208 13800 222
rect 13800 208 13812 222
rect 13850 208 13868 222
rect 13868 208 13884 222
rect 13922 208 13936 222
rect 13936 208 13956 222
rect 13634 188 13668 208
rect 13706 188 13740 208
rect 13778 188 13812 208
rect 13850 188 13884 208
rect 13922 188 13956 208
rect 13202 139 13222 149
rect 13222 139 13236 149
rect 13274 139 13290 149
rect 13290 139 13308 149
rect 13346 139 13358 149
rect 13358 139 13380 149
rect 13418 139 13426 149
rect 13426 139 13452 149
rect 13490 139 13494 149
rect 13494 139 13524 149
rect 13202 115 13236 139
rect 13274 115 13308 139
rect 13346 115 13380 139
rect 13418 115 13452 139
rect 13490 115 13524 139
rect 13562 115 13596 149
rect 13634 139 13664 149
rect 13664 139 13668 149
rect 13706 139 13732 149
rect 13732 139 13740 149
rect 13778 139 13800 149
rect 13800 139 13812 149
rect 13850 139 13868 149
rect 13868 139 13884 149
rect 13922 139 13936 149
rect 13936 139 13956 149
rect 13634 115 13668 139
rect 13706 115 13740 139
rect 13778 115 13812 139
rect 13850 115 13884 139
rect 13922 115 13956 139
rect 13202 70 13222 76
rect 13222 70 13236 76
rect 13274 70 13290 76
rect 13290 70 13308 76
rect 13346 70 13358 76
rect 13358 70 13380 76
rect 13418 70 13426 76
rect 13426 70 13452 76
rect 13490 70 13494 76
rect 13494 70 13524 76
rect 13202 42 13236 70
rect 13274 42 13308 70
rect 13346 42 13380 70
rect 13418 42 13452 70
rect 13490 42 13524 70
rect 13562 42 13596 76
rect 13634 70 13664 76
rect 13664 70 13668 76
rect 13706 70 13732 76
rect 13732 70 13740 76
rect 13778 70 13800 76
rect 13800 70 13812 76
rect 13850 70 13868 76
rect 13868 70 13884 76
rect 13922 70 13936 76
rect 13936 70 13956 76
rect 13634 42 13668 70
rect 13706 42 13740 70
rect 13778 42 13812 70
rect 13850 42 13884 70
rect 13922 42 13956 70
rect 13202 1 13222 3
rect 13222 1 13236 3
rect 13274 1 13290 3
rect 13290 1 13308 3
rect 13346 1 13358 3
rect 13358 1 13380 3
rect 13418 1 13426 3
rect 13426 1 13452 3
rect 13490 1 13494 3
rect 13494 1 13524 3
rect -1074 -103 -1040 -70
rect -1002 -103 -968 -70
rect -930 -103 -896 -70
rect -858 -103 -824 -70
rect -786 -103 -752 -70
rect -1074 -104 -1054 -103
rect -1054 -104 -1040 -103
rect -1002 -104 -986 -103
rect -986 -104 -968 -103
rect -930 -104 -918 -103
rect -918 -104 -896 -103
rect -858 -104 -850 -103
rect -850 -104 -824 -103
rect -786 -104 -782 -103
rect -782 -104 -752 -103
rect -714 -104 -680 -70
rect -642 -103 -608 -70
rect -570 -103 -536 -70
rect -498 -103 -464 -70
rect -426 -103 -392 -70
rect -354 -103 -320 -70
rect -642 -104 -612 -103
rect -612 -104 -608 -103
rect -570 -104 -544 -103
rect -544 -104 -536 -103
rect -498 -104 -476 -103
rect -476 -104 -464 -103
rect -426 -104 -408 -103
rect -408 -104 -392 -103
rect -354 -104 -340 -103
rect -340 -104 -320 -103
rect -1074 -172 -1040 -143
rect -1002 -172 -968 -143
rect -930 -172 -896 -143
rect -858 -172 -824 -143
rect -786 -172 -752 -143
rect -1074 -177 -1054 -172
rect -1054 -177 -1040 -172
rect -1002 -177 -986 -172
rect -986 -177 -968 -172
rect -930 -177 -918 -172
rect -918 -177 -896 -172
rect -858 -177 -850 -172
rect -850 -177 -824 -172
rect -786 -177 -782 -172
rect -782 -177 -752 -172
rect -714 -177 -680 -143
rect -642 -172 -608 -143
rect -570 -172 -536 -143
rect -498 -172 -464 -143
rect -426 -172 -392 -143
rect -354 -172 -320 -143
rect -642 -177 -612 -172
rect -612 -177 -608 -172
rect -570 -177 -544 -172
rect -544 -177 -536 -172
rect -498 -177 -476 -172
rect -476 -177 -464 -172
rect -426 -177 -408 -172
rect -408 -177 -392 -172
rect -354 -177 -340 -172
rect -340 -177 -320 -172
rect 13202 -31 13236 1
rect 13274 -31 13308 1
rect 13346 -31 13380 1
rect 13418 -31 13452 1
rect 13490 -31 13524 1
rect 13562 -31 13596 3
rect 13634 1 13664 3
rect 13664 1 13668 3
rect 13706 1 13732 3
rect 13732 1 13740 3
rect 13778 1 13800 3
rect 13800 1 13812 3
rect 13850 1 13868 3
rect 13868 1 13884 3
rect 13922 1 13936 3
rect 13936 1 13956 3
rect 13634 -31 13668 1
rect 13706 -31 13740 1
rect 13778 -31 13812 1
rect 13850 -31 13884 1
rect 13922 -31 13956 1
rect 13202 -103 13236 -70
rect 13274 -103 13308 -70
rect 13346 -103 13380 -70
rect 13418 -103 13452 -70
rect 13490 -103 13524 -70
rect 13202 -104 13222 -103
rect 13222 -104 13236 -103
rect 13274 -104 13290 -103
rect 13290 -104 13308 -103
rect 13346 -104 13358 -103
rect 13358 -104 13380 -103
rect 13418 -104 13426 -103
rect 13426 -104 13452 -103
rect 13490 -104 13494 -103
rect 13494 -104 13524 -103
rect 13562 -104 13596 -70
rect 13634 -103 13668 -70
rect 13706 -103 13740 -70
rect 13778 -103 13812 -70
rect 13850 -103 13884 -70
rect 13922 -103 13956 -70
rect 13634 -104 13664 -103
rect 13664 -104 13668 -103
rect 13706 -104 13732 -103
rect 13732 -104 13740 -103
rect 13778 -104 13800 -103
rect 13800 -104 13812 -103
rect 13850 -104 13868 -103
rect 13868 -104 13884 -103
rect 13922 -104 13936 -103
rect 13936 -104 13956 -103
rect 13202 -172 13236 -143
rect 13274 -172 13308 -143
rect 13346 -172 13380 -143
rect 13418 -172 13452 -143
rect 13490 -172 13524 -143
rect 13202 -177 13222 -172
rect 13222 -177 13236 -172
rect 13274 -177 13290 -172
rect 13290 -177 13308 -172
rect 13346 -177 13358 -172
rect 13358 -177 13380 -172
rect 13418 -177 13426 -172
rect 13426 -177 13452 -172
rect 13490 -177 13494 -172
rect 13494 -177 13524 -172
rect 13562 -177 13596 -143
rect 13634 -172 13668 -143
rect 13706 -172 13740 -143
rect 13778 -172 13812 -143
rect 13850 -172 13884 -143
rect 13922 -172 13956 -143
rect 13634 -177 13664 -172
rect 13664 -177 13668 -172
rect 13706 -177 13732 -172
rect 13732 -177 13740 -172
rect 13778 -177 13800 -172
rect 13800 -177 13812 -172
rect 13850 -177 13868 -172
rect 13868 -177 13884 -172
rect 13922 -177 13936 -172
rect 13936 -177 13956 -172
rect -886 -308 -882 -306
rect -882 -308 -852 -306
rect -813 -308 -779 -306
rect -740 -308 -710 -306
rect -710 -308 -706 -306
rect -667 -308 -641 -306
rect -641 -308 -633 -306
rect -594 -308 -572 -306
rect -572 -308 -537 -306
rect -537 -308 -503 -306
rect -503 -308 -468 -306
rect -468 -308 -434 -306
rect -434 -308 -399 -306
rect -399 -308 -365 -306
rect -365 -308 -330 -306
rect -330 -308 -296 -306
rect -296 -308 -261 -306
rect -261 -308 -227 -306
rect -227 -308 -192 -306
rect -192 -308 -158 -306
rect -158 -308 -123 -306
rect -123 -308 -89 -306
rect -89 -308 -54 -306
rect -54 -308 -20 -306
rect -20 -308 15 -306
rect 15 -308 49 -306
rect 49 -308 84 -306
rect 84 -308 118 -306
rect 118 -308 153 -306
rect 153 -308 187 -306
rect 187 -308 222 -306
rect 222 -308 256 -306
rect 256 -308 291 -306
rect 291 -308 325 -306
rect 325 -308 360 -306
rect 360 -308 394 -306
rect 394 -308 429 -306
rect 429 -308 463 -306
rect 463 -308 498 -306
rect 498 -308 532 -306
rect 532 -308 567 -306
rect 567 -308 601 -306
rect 601 -308 636 -306
rect 636 -308 670 -306
rect 670 -308 705 -306
rect 705 -308 739 -306
rect 739 -308 774 -306
rect 774 -308 808 -306
rect 808 -308 843 -306
rect 843 -308 877 -306
rect 877 -308 912 -306
rect 912 -308 946 -306
rect 946 -308 981 -306
rect 981 -308 1015 -306
rect 1015 -308 1050 -306
rect 1050 -308 1084 -306
rect 1084 -308 1119 -306
rect 1119 -308 1153 -306
rect 1153 -308 1188 -306
rect 1188 -308 1222 -306
rect 1222 -308 1257 -306
rect 1257 -308 1291 -306
rect 1291 -308 1326 -306
rect 1326 -308 1360 -306
rect 1360 -308 1395 -306
rect 1395 -308 1429 -306
rect 1429 -308 1464 -306
rect 1464 -308 1498 -306
rect 1498 -308 1533 -306
rect 1533 -308 1567 -306
rect 1567 -308 1602 -306
rect 1602 -308 1636 -306
rect 1636 -308 1671 -306
rect 1671 -308 1705 -306
rect 1705 -308 1740 -306
rect 1740 -308 1774 -306
rect 1774 -308 1809 -306
rect 1809 -308 1843 -306
rect 1843 -308 1878 -306
rect 1878 -308 1912 -306
rect 1912 -308 1947 -306
rect 1947 -308 1981 -306
rect 1981 -308 2016 -306
rect 2016 -308 2050 -306
rect 2050 -308 2085 -306
rect 2085 -308 2119 -306
rect 2119 -308 2154 -306
rect 2154 -308 2188 -306
rect 2188 -308 2223 -306
rect 2223 -308 2257 -306
rect 2257 -308 2292 -306
rect 2292 -308 2326 -306
rect 2326 -308 2361 -306
rect 2361 -308 2395 -306
rect 2395 -308 2430 -306
rect 2430 -308 2464 -306
rect 2464 -308 2499 -306
rect 2499 -308 2533 -306
rect 2533 -308 2568 -306
rect 2568 -308 2602 -306
rect 2602 -308 2637 -306
rect 2637 -308 2671 -306
rect 2671 -308 2706 -306
rect 2706 -308 2740 -306
rect 2740 -308 2775 -306
rect 2775 -308 2809 -306
rect 2809 -308 2844 -306
rect 2844 -308 2878 -306
rect 2878 -308 2913 -306
rect 2913 -308 2947 -306
rect 2947 -308 2982 -306
rect 2982 -308 3016 -306
rect 3016 -308 3051 -306
rect 3051 -308 3085 -306
rect 3085 -308 3120 -306
rect 3120 -308 3154 -306
rect 3154 -308 3189 -306
rect 3189 -308 3223 -306
rect 3223 -308 3258 -306
rect 3258 -308 3292 -306
rect 3292 -308 3327 -306
rect 3327 -308 3361 -306
rect 3361 -308 3396 -306
rect -886 -340 -852 -308
rect -813 -340 -779 -308
rect -740 -340 -706 -308
rect -667 -340 -633 -308
rect -594 -342 3396 -308
rect -594 -376 -572 -342
rect -572 -376 -537 -342
rect -537 -376 -503 -342
rect -503 -376 -468 -342
rect -468 -376 -434 -342
rect -434 -376 -399 -342
rect -399 -376 -365 -342
rect -365 -376 -330 -342
rect -330 -376 -296 -342
rect -296 -376 -261 -342
rect -261 -376 -227 -342
rect -227 -376 -192 -342
rect -192 -376 -158 -342
rect -158 -376 -123 -342
rect -123 -376 -89 -342
rect -89 -376 -54 -342
rect -54 -376 -20 -342
rect -20 -376 15 -342
rect 15 -376 49 -342
rect 49 -376 84 -342
rect 84 -376 118 -342
rect 118 -376 153 -342
rect 153 -376 187 -342
rect 187 -376 222 -342
rect 222 -376 256 -342
rect 256 -376 291 -342
rect 291 -376 325 -342
rect 325 -376 360 -342
rect 360 -376 394 -342
rect 394 -376 429 -342
rect 429 -376 463 -342
rect 463 -376 498 -342
rect 498 -376 532 -342
rect 532 -376 567 -342
rect 567 -376 601 -342
rect 601 -376 636 -342
rect 636 -376 670 -342
rect 670 -376 705 -342
rect 705 -376 739 -342
rect 739 -376 774 -342
rect 774 -376 808 -342
rect 808 -376 843 -342
rect 843 -376 877 -342
rect 877 -376 912 -342
rect 912 -376 946 -342
rect 946 -376 981 -342
rect 981 -376 1015 -342
rect 1015 -376 1050 -342
rect 1050 -376 1084 -342
rect 1084 -376 1119 -342
rect 1119 -376 1153 -342
rect 1153 -376 1188 -342
rect 1188 -376 1222 -342
rect 1222 -376 1257 -342
rect 1257 -376 1291 -342
rect 1291 -376 1326 -342
rect 1326 -376 1360 -342
rect 1360 -376 1395 -342
rect 1395 -376 1429 -342
rect 1429 -376 1464 -342
rect 1464 -376 1498 -342
rect 1498 -376 1533 -342
rect 1533 -376 1567 -342
rect 1567 -376 1602 -342
rect 1602 -376 1636 -342
rect 1636 -376 1671 -342
rect 1671 -376 1705 -342
rect 1705 -376 1740 -342
rect 1740 -376 1774 -342
rect 1774 -376 1809 -342
rect 1809 -376 1843 -342
rect 1843 -376 1878 -342
rect 1878 -376 1912 -342
rect 1912 -376 1947 -342
rect 1947 -376 1981 -342
rect 1981 -376 2016 -342
rect 2016 -376 2050 -342
rect 2050 -376 2085 -342
rect 2085 -376 2119 -342
rect 2119 -376 2154 -342
rect 2154 -376 2188 -342
rect 2188 -376 2223 -342
rect 2223 -376 2257 -342
rect 2257 -376 2292 -342
rect 2292 -376 2326 -342
rect 2326 -376 2361 -342
rect 2361 -376 2395 -342
rect 2395 -376 2430 -342
rect 2430 -376 2464 -342
rect 2464 -376 2499 -342
rect 2499 -376 2533 -342
rect 2533 -376 2568 -342
rect 2568 -376 2602 -342
rect 2602 -376 2637 -342
rect 2637 -376 2671 -342
rect 2671 -376 2706 -342
rect 2706 -376 2740 -342
rect 2740 -376 2775 -342
rect 2775 -376 2809 -342
rect 2809 -376 2844 -342
rect 2844 -376 2878 -342
rect 2878 -376 2913 -342
rect 2913 -376 2947 -342
rect 2947 -376 2982 -342
rect 2982 -376 3016 -342
rect 3016 -376 3051 -342
rect 3051 -376 3085 -342
rect 3085 -376 3120 -342
rect 3120 -376 3154 -342
rect 3154 -376 3189 -342
rect 3189 -376 3223 -342
rect 3223 -376 3258 -342
rect 3258 -376 3292 -342
rect 3292 -376 3327 -342
rect 3327 -376 3361 -342
rect 3361 -376 3396 -342
rect -886 -410 -852 -378
rect -813 -410 -779 -378
rect -740 -410 -706 -378
rect -667 -410 -633 -378
rect -594 -410 3396 -376
rect -886 -412 -882 -410
rect -882 -412 -852 -410
rect -813 -412 -779 -410
rect -740 -412 -710 -410
rect -710 -412 -706 -410
rect -667 -412 -641 -410
rect -641 -412 -633 -410
rect -594 -412 -572 -410
rect -572 -412 -537 -410
rect -537 -412 -503 -410
rect -503 -412 -468 -410
rect -468 -412 -434 -410
rect -434 -412 -399 -410
rect -399 -412 -365 -410
rect -365 -412 -330 -410
rect -330 -412 -296 -410
rect -296 -412 -261 -410
rect -261 -412 -227 -410
rect -227 -412 -192 -410
rect -192 -412 -158 -410
rect -158 -412 -123 -410
rect -123 -412 -89 -410
rect -89 -412 -54 -410
rect -54 -412 -20 -410
rect -20 -412 15 -410
rect 15 -412 49 -410
rect 49 -412 84 -410
rect 84 -412 118 -410
rect 118 -412 153 -410
rect 153 -412 187 -410
rect 187 -412 222 -410
rect 222 -412 256 -410
rect 256 -412 291 -410
rect 291 -412 325 -410
rect 325 -412 360 -410
rect 360 -412 394 -410
rect 394 -412 429 -410
rect 429 -412 463 -410
rect 463 -412 498 -410
rect 498 -412 532 -410
rect 532 -412 567 -410
rect 567 -412 601 -410
rect 601 -412 636 -410
rect 636 -412 670 -410
rect 670 -412 705 -410
rect 705 -412 739 -410
rect 739 -412 774 -410
rect 774 -412 808 -410
rect 808 -412 843 -410
rect 843 -412 877 -410
rect 877 -412 912 -410
rect 912 -412 946 -410
rect 946 -412 981 -410
rect 981 -412 1015 -410
rect 1015 -412 1050 -410
rect 1050 -412 1084 -410
rect 1084 -412 1119 -410
rect 1119 -412 1153 -410
rect 1153 -412 1188 -410
rect 1188 -412 1222 -410
rect 1222 -412 1257 -410
rect 1257 -412 1291 -410
rect 1291 -412 1326 -410
rect 1326 -412 1360 -410
rect 1360 -412 1395 -410
rect 1395 -412 1429 -410
rect 1429 -412 1464 -410
rect 1464 -412 1498 -410
rect 1498 -412 1533 -410
rect 1533 -412 1567 -410
rect 1567 -412 1602 -410
rect 1602 -412 1636 -410
rect 1636 -412 1671 -410
rect 1671 -412 1705 -410
rect 1705 -412 1740 -410
rect 1740 -412 1774 -410
rect 1774 -412 1809 -410
rect 1809 -412 1843 -410
rect 1843 -412 1878 -410
rect 1878 -412 1912 -410
rect 1912 -412 1947 -410
rect 1947 -412 1981 -410
rect 1981 -412 2016 -410
rect 2016 -412 2050 -410
rect 2050 -412 2085 -410
rect 2085 -412 2119 -410
rect 2119 -412 2154 -410
rect 2154 -412 2188 -410
rect 2188 -412 2223 -410
rect 2223 -412 2257 -410
rect 2257 -412 2292 -410
rect 2292 -412 2326 -410
rect 2326 -412 2361 -410
rect 2361 -412 2395 -410
rect 2395 -412 2430 -410
rect 2430 -412 2464 -410
rect 2464 -412 2499 -410
rect 2499 -412 2533 -410
rect 2533 -412 2568 -410
rect 2568 -412 2602 -410
rect 2602 -412 2637 -410
rect 2637 -412 2671 -410
rect 2671 -412 2706 -410
rect 2706 -412 2740 -410
rect 2740 -412 2775 -410
rect 2775 -412 2809 -410
rect 2809 -412 2844 -410
rect 2844 -412 2878 -410
rect 2878 -412 2913 -410
rect 2913 -412 2947 -410
rect 2947 -412 2982 -410
rect 2982 -412 3016 -410
rect 3016 -412 3051 -410
rect 3051 -412 3085 -410
rect 3085 -412 3120 -410
rect 3120 -412 3154 -410
rect 3154 -412 3189 -410
rect 3189 -412 3223 -410
rect 3223 -412 3258 -410
rect 3258 -412 3292 -410
rect 3292 -412 3327 -410
rect 3327 -412 3361 -410
rect 3361 -412 3396 -410
rect 3396 -412 13768 -306
rect 14202 3541 14308 3647
rect 14202 3468 14236 3502
rect 14274 3468 14308 3502
rect 14202 3395 14236 3429
rect 14274 3395 14308 3429
rect 14202 3322 14236 3356
rect 14274 3322 14308 3356
rect 14202 3249 14236 3283
rect 14274 3249 14308 3283
rect 14202 3176 14236 3210
rect 14274 3176 14308 3210
rect 14202 3103 14236 3137
rect 14274 3103 14308 3137
rect 14202 3030 14236 3064
rect 14274 3030 14308 3064
rect 14202 2957 14236 2991
rect 14274 2957 14308 2991
rect 14202 2884 14236 2918
rect 14274 2884 14308 2918
rect 14202 2811 14236 2845
rect 14274 2811 14308 2845
rect 14202 2738 14236 2772
rect 14274 2738 14308 2772
rect 14202 2665 14236 2699
rect 14274 2665 14308 2699
rect 14202 2592 14236 2626
rect 14274 2592 14308 2626
rect 14202 2519 14236 2553
rect 14274 2519 14308 2553
rect 14202 2446 14236 2480
rect 14274 2446 14308 2480
rect 14202 2373 14236 2407
rect 14274 2373 14308 2407
rect 14202 2300 14236 2334
rect 14274 2300 14308 2334
rect 14202 2227 14236 2261
rect 14274 2227 14308 2261
rect 14202 2154 14236 2188
rect 14274 2154 14308 2188
rect 14202 2081 14236 2115
rect 14274 2081 14308 2115
rect 14202 2008 14236 2042
rect 14274 2008 14308 2042
rect 14202 1935 14236 1969
rect 14274 1935 14308 1969
rect 14202 1862 14236 1896
rect 14274 1862 14308 1896
rect 14202 1789 14236 1823
rect 14274 1789 14308 1823
rect 14202 1716 14236 1750
rect 14274 1716 14308 1750
rect 14202 1643 14236 1677
rect 14274 1643 14308 1677
rect 14202 1570 14236 1604
rect 14274 1570 14308 1604
rect 14202 1497 14236 1531
rect 14274 1497 14308 1531
rect 14202 1424 14236 1458
rect 14274 1424 14308 1458
rect 14202 1351 14236 1385
rect 14274 1351 14308 1385
rect 14202 1278 14236 1312
rect 14274 1278 14308 1312
rect 14202 1205 14236 1239
rect 14274 1205 14308 1239
rect 14202 1132 14236 1166
rect 14274 1132 14308 1166
rect 14202 1059 14236 1093
rect 14274 1059 14308 1093
rect 14202 986 14236 1020
rect 14274 986 14308 1020
rect 14202 913 14236 947
rect 14274 913 14308 947
rect 14202 840 14236 874
rect 14274 840 14308 874
rect 14202 767 14236 801
rect 14274 767 14308 801
rect 14202 694 14236 728
rect 14274 694 14308 728
rect 14202 621 14236 655
rect 14274 621 14308 655
rect 14202 548 14236 582
rect 14274 548 14308 582
rect 14202 475 14236 509
rect 14274 475 14308 509
rect 14202 402 14236 436
rect 14274 402 14308 436
rect 14202 329 14236 363
rect 14274 329 14308 363
rect 14202 256 14236 290
rect 14274 256 14308 290
rect 14202 183 14236 217
rect 14274 183 14308 217
rect 14202 110 14236 144
rect 14274 110 14308 144
rect 14202 37 14236 71
rect 14274 37 14308 71
rect 14202 -36 14236 -2
rect 14274 -36 14308 -2
rect 14202 -109 14236 -75
rect 14274 -109 14308 -75
rect 14202 -182 14236 -148
rect 14274 -182 14308 -148
rect 14202 -255 14236 -221
rect 14274 -255 14308 -221
rect 14202 -328 14236 -294
rect 14274 -328 14308 -294
rect 14202 -401 14236 -367
rect 14274 -401 14308 -367
rect -1426 -474 -1424 -473
rect -1424 -474 -1392 -473
rect -1354 -474 -1322 -473
rect -1322 -474 -1320 -473
rect -1426 -542 -1392 -513
rect -1354 -542 -1320 -513
rect -1426 -547 -1424 -542
rect -1424 -547 -1392 -542
rect -1354 -547 -1322 -542
rect -1322 -547 -1320 -542
rect 14202 -473 14236 -440
rect 14274 -473 14308 -440
rect 14202 -474 14204 -473
rect 14204 -474 14236 -473
rect 14274 -474 14306 -473
rect 14306 -474 14308 -473
rect 14202 -542 14236 -513
rect 14274 -542 14308 -513
rect 14202 -547 14204 -542
rect 14204 -547 14236 -542
rect 14274 -547 14306 -542
rect 14306 -547 14308 -542
rect -1191 -678 -1183 -676
rect -1183 -678 -1157 -676
rect -1118 -678 -1114 -676
rect -1114 -678 -1084 -676
rect -1045 -678 -1011 -676
rect -972 -678 -942 -676
rect -942 -678 -938 -676
rect -899 -678 -873 -676
rect -873 -678 -865 -676
rect -826 -678 -804 -676
rect -804 -678 -792 -676
rect -753 -678 -735 -676
rect -735 -678 -719 -676
rect -680 -678 -666 -676
rect -666 -678 -646 -676
rect -607 -678 -597 -676
rect -597 -678 -573 -676
rect -534 -678 -528 -676
rect -528 -678 -500 -676
rect -461 -678 -459 -676
rect -459 -678 -427 -676
rect -388 -678 -355 -676
rect -355 -678 -354 -676
rect -315 -678 -286 -676
rect -286 -678 -281 -676
rect -242 -678 -217 -676
rect -217 -678 -208 -676
rect -169 -678 -148 -676
rect -148 -678 -135 -676
rect -96 -678 -79 -676
rect -79 -678 -62 -676
rect -23 -678 -10 -676
rect -10 -678 11 -676
rect 50 -678 59 -676
rect 59 -678 84 -676
rect 123 -678 128 -676
rect 128 -678 157 -676
rect 196 -678 197 -676
rect 197 -678 230 -676
rect 269 -678 300 -676
rect 300 -678 303 -676
rect 342 -678 369 -676
rect 369 -678 376 -676
rect 415 -678 438 -676
rect 438 -678 449 -676
rect 488 -678 507 -676
rect 507 -678 522 -676
rect 561 -678 576 -676
rect 576 -678 595 -676
rect 634 -678 645 -676
rect 645 -678 668 -676
rect 707 -678 714 -676
rect 714 -678 741 -676
rect 780 -678 783 -676
rect 783 -678 814 -676
rect -1191 -710 -1157 -678
rect -1118 -710 -1084 -678
rect -1045 -710 -1011 -678
rect -972 -710 -938 -678
rect -899 -710 -865 -678
rect -826 -710 -792 -678
rect -753 -710 -719 -678
rect -680 -710 -646 -678
rect -607 -710 -573 -678
rect -534 -710 -500 -678
rect -461 -710 -427 -678
rect -388 -710 -354 -678
rect -315 -710 -281 -678
rect -242 -710 -208 -678
rect -169 -710 -135 -678
rect -96 -710 -62 -678
rect -23 -710 11 -678
rect 50 -710 84 -678
rect 123 -710 157 -678
rect 196 -710 230 -678
rect 269 -710 303 -678
rect 342 -710 376 -678
rect 415 -710 449 -678
rect 488 -710 522 -678
rect 561 -710 595 -678
rect 634 -710 668 -678
rect 707 -710 741 -678
rect 780 -710 814 -678
rect 853 -710 887 -676
rect 926 -678 956 -676
rect 956 -678 960 -676
rect 999 -678 1025 -676
rect 1025 -678 1033 -676
rect 1072 -678 1094 -676
rect 1094 -678 1106 -676
rect 1145 -678 1163 -676
rect 1163 -678 1179 -676
rect 1218 -678 1232 -676
rect 1232 -678 1252 -676
rect 1291 -678 1301 -676
rect 1301 -678 1325 -676
rect 1364 -678 1370 -676
rect 1370 -678 1398 -676
rect 1437 -678 1439 -676
rect 1439 -678 1471 -676
rect 1510 -678 1542 -676
rect 1542 -678 1544 -676
rect 1583 -678 1611 -676
rect 1611 -678 1646 -676
rect 1646 -678 1680 -676
rect 1680 -678 1715 -676
rect 1715 -678 1749 -676
rect 1749 -678 1784 -676
rect 1784 -678 1818 -676
rect 1818 -678 1853 -676
rect 1853 -678 1887 -676
rect 1887 -678 1922 -676
rect 1922 -678 1956 -676
rect 1956 -678 1991 -676
rect 1991 -678 2025 -676
rect 2025 -678 2060 -676
rect 2060 -678 2094 -676
rect 2094 -678 2129 -676
rect 2129 -678 2163 -676
rect 2163 -678 2198 -676
rect 2198 -678 2232 -676
rect 2232 -678 2267 -676
rect 2267 -678 2301 -676
rect 2301 -678 2336 -676
rect 2336 -678 2370 -676
rect 2370 -678 2405 -676
rect 2405 -678 2439 -676
rect 2439 -678 2474 -676
rect 926 -710 960 -678
rect 999 -710 1033 -678
rect 1072 -710 1106 -678
rect 1145 -710 1179 -678
rect 1218 -710 1252 -678
rect 1291 -710 1325 -678
rect 1364 -710 1398 -678
rect 1437 -710 1471 -678
rect 1510 -710 1544 -678
rect 1583 -712 2474 -678
rect 1583 -746 1611 -712
rect 1611 -746 1646 -712
rect 1646 -746 1680 -712
rect 1680 -746 1715 -712
rect 1715 -746 1749 -712
rect 1749 -746 1784 -712
rect 1784 -746 1818 -712
rect 1818 -746 1853 -712
rect 1853 -746 1887 -712
rect 1887 -746 1922 -712
rect 1922 -746 1956 -712
rect 1956 -746 1991 -712
rect 1991 -746 2025 -712
rect 2025 -746 2060 -712
rect 2060 -746 2094 -712
rect 2094 -746 2129 -712
rect 2129 -746 2163 -712
rect 2163 -746 2198 -712
rect 2198 -746 2232 -712
rect 2232 -746 2267 -712
rect 2267 -746 2301 -712
rect 2301 -746 2336 -712
rect 2336 -746 2370 -712
rect 2370 -746 2405 -712
rect 2405 -746 2439 -712
rect 2439 -746 2474 -712
rect -1191 -780 -1157 -748
rect -1118 -780 -1084 -748
rect -1045 -780 -1011 -748
rect -972 -780 -938 -748
rect -899 -780 -865 -748
rect -826 -780 -792 -748
rect -753 -780 -719 -748
rect -680 -780 -646 -748
rect -607 -780 -573 -748
rect -534 -780 -500 -748
rect -461 -780 -427 -748
rect -388 -780 -354 -748
rect -315 -780 -281 -748
rect -242 -780 -208 -748
rect -169 -780 -135 -748
rect -96 -780 -62 -748
rect -23 -780 11 -748
rect 50 -780 84 -748
rect 123 -780 157 -748
rect 196 -780 230 -748
rect 269 -780 303 -748
rect 342 -780 376 -748
rect 415 -780 449 -748
rect 488 -780 522 -748
rect 561 -780 595 -748
rect 634 -780 668 -748
rect 707 -780 741 -748
rect 780 -780 814 -748
rect -1191 -782 -1183 -780
rect -1183 -782 -1157 -780
rect -1118 -782 -1114 -780
rect -1114 -782 -1084 -780
rect -1045 -782 -1011 -780
rect -972 -782 -942 -780
rect -942 -782 -938 -780
rect -899 -782 -873 -780
rect -873 -782 -865 -780
rect -826 -782 -804 -780
rect -804 -782 -792 -780
rect -753 -782 -735 -780
rect -735 -782 -719 -780
rect -680 -782 -666 -780
rect -666 -782 -646 -780
rect -607 -782 -597 -780
rect -597 -782 -573 -780
rect -534 -782 -528 -780
rect -528 -782 -500 -780
rect -461 -782 -459 -780
rect -459 -782 -427 -780
rect -388 -782 -355 -780
rect -355 -782 -354 -780
rect -315 -782 -286 -780
rect -286 -782 -281 -780
rect -242 -782 -217 -780
rect -217 -782 -208 -780
rect -169 -782 -148 -780
rect -148 -782 -135 -780
rect -96 -782 -79 -780
rect -79 -782 -62 -780
rect -23 -782 -10 -780
rect -10 -782 11 -780
rect 50 -782 59 -780
rect 59 -782 84 -780
rect 123 -782 128 -780
rect 128 -782 157 -780
rect 196 -782 197 -780
rect 197 -782 230 -780
rect 269 -782 300 -780
rect 300 -782 303 -780
rect 342 -782 369 -780
rect 369 -782 376 -780
rect 415 -782 438 -780
rect 438 -782 449 -780
rect 488 -782 507 -780
rect 507 -782 522 -780
rect 561 -782 576 -780
rect 576 -782 595 -780
rect 634 -782 645 -780
rect 645 -782 668 -780
rect 707 -782 714 -780
rect 714 -782 741 -780
rect 780 -782 783 -780
rect 783 -782 814 -780
rect 853 -782 887 -748
rect 926 -780 960 -748
rect 999 -780 1033 -748
rect 1072 -780 1106 -748
rect 1145 -780 1179 -748
rect 1218 -780 1252 -748
rect 1291 -780 1325 -748
rect 1364 -780 1398 -748
rect 1437 -780 1471 -748
rect 1510 -780 1544 -748
rect 1583 -780 2474 -746
rect 926 -782 956 -780
rect 956 -782 960 -780
rect 999 -782 1025 -780
rect 1025 -782 1033 -780
rect 1072 -782 1094 -780
rect 1094 -782 1106 -780
rect 1145 -782 1163 -780
rect 1163 -782 1179 -780
rect 1218 -782 1232 -780
rect 1232 -782 1252 -780
rect 1291 -782 1301 -780
rect 1301 -782 1325 -780
rect 1364 -782 1370 -780
rect 1370 -782 1398 -780
rect 1437 -782 1439 -780
rect 1439 -782 1471 -780
rect 1510 -782 1542 -780
rect 1542 -782 1544 -780
rect 1583 -782 1611 -780
rect 1611 -782 1646 -780
rect 1646 -782 1680 -780
rect 1680 -782 1715 -780
rect 1715 -782 1749 -780
rect 1749 -782 1784 -780
rect 1784 -782 1818 -780
rect 1818 -782 1853 -780
rect 1853 -782 1887 -780
rect 1887 -782 1922 -780
rect 1922 -782 1956 -780
rect 1956 -782 1991 -780
rect 1991 -782 2025 -780
rect 2025 -782 2060 -780
rect 2060 -782 2094 -780
rect 2094 -782 2129 -780
rect 2129 -782 2163 -780
rect 2163 -782 2198 -780
rect 2198 -782 2232 -780
rect 2232 -782 2267 -780
rect 2267 -782 2301 -780
rect 2301 -782 2336 -780
rect 2336 -782 2370 -780
rect 2370 -782 2405 -780
rect 2405 -782 2439 -780
rect 2439 -782 2474 -780
rect 2474 -782 14073 -676
<< metal1 >>
tri -1320 3882 -1308 3894 se
rect -1308 3882 14190 3894
tri -1354 3848 -1320 3882 se
rect -1320 3848 -1191 3882
rect -1157 3848 -1118 3882
rect -1084 3848 -1045 3882
rect -1011 3848 -972 3882
rect -938 3848 -899 3882
rect -865 3848 -826 3882
rect -792 3848 -753 3882
rect -719 3848 -680 3882
rect -646 3848 -607 3882
rect -573 3848 -534 3882
rect -500 3848 -461 3882
rect -427 3848 -388 3882
rect -354 3848 -315 3882
rect -281 3848 -242 3882
rect -208 3848 -169 3882
rect -135 3848 -96 3882
rect -62 3848 -23 3882
rect 11 3848 50 3882
rect 84 3848 123 3882
rect 157 3848 196 3882
rect 230 3848 269 3882
rect 303 3848 342 3882
rect 376 3848 415 3882
rect 449 3848 488 3882
rect 522 3848 561 3882
rect 595 3848 634 3882
rect 668 3848 707 3882
rect 741 3848 780 3882
rect 814 3848 853 3882
rect 887 3848 926 3882
rect 960 3848 999 3882
rect 1033 3848 1072 3882
rect 1106 3848 1145 3882
rect 1179 3848 1218 3882
rect 1252 3848 1291 3882
rect 1325 3848 1364 3882
rect 1398 3848 1437 3882
rect 1471 3848 1510 3882
rect 1544 3848 1583 3882
tri -1392 3810 -1354 3848 se
rect -1354 3810 1583 3848
tri -1426 3776 -1392 3810 se
rect -1392 3776 -1191 3810
rect -1157 3776 -1118 3810
rect -1084 3776 -1045 3810
rect -1011 3776 -972 3810
rect -938 3776 -899 3810
rect -865 3776 -826 3810
rect -792 3776 -753 3810
rect -719 3776 -680 3810
rect -646 3776 -607 3810
rect -573 3776 -534 3810
rect -500 3776 -461 3810
rect -427 3776 -388 3810
rect -354 3776 -315 3810
rect -281 3776 -242 3810
rect -208 3776 -169 3810
rect -135 3776 -96 3810
rect -62 3776 -23 3810
rect 11 3776 50 3810
rect 84 3776 123 3810
rect 157 3776 196 3810
rect 230 3776 269 3810
rect 303 3776 342 3810
rect 376 3776 415 3810
rect 449 3776 488 3810
rect 522 3776 561 3810
rect 595 3776 634 3810
rect 668 3776 707 3810
rect 741 3776 780 3810
rect 814 3776 853 3810
rect 887 3776 926 3810
rect 960 3776 999 3810
rect 1033 3776 1072 3810
rect 1106 3776 1145 3810
rect 1179 3776 1218 3810
rect 1252 3776 1291 3810
rect 1325 3776 1364 3810
rect 1398 3776 1437 3810
rect 1471 3776 1510 3810
rect 1544 3776 1583 3810
rect 14073 3776 14190 3882
tri -1438 3764 -1426 3776 se
rect -1426 3764 14190 3776
tri 14190 3764 14320 3894 sw
rect -1438 3719 -1245 3764
tri -1245 3719 -1200 3764 nw
tri 14082 3719 14127 3764 ne
rect 14127 3719 14320 3764
rect -1438 3647 -1308 3719
tri -1308 3656 -1245 3719 nw
tri 14127 3656 14190 3719 ne
rect -1438 3541 -1426 3647
rect -1320 3541 -1308 3647
rect -1438 3502 -1308 3541
rect 14190 3647 14320 3719
rect 14190 3541 14202 3647
rect 14308 3541 14320 3647
tri -968 3512 -958 3522 se
rect -958 3512 13840 3524
rect -1438 3468 -1426 3502
rect -1392 3468 -1354 3502
rect -1320 3468 -1308 3502
tri -1002 3478 -968 3512 se
rect -968 3478 -886 3512
rect -852 3478 -813 3512
rect -779 3478 -740 3512
rect -706 3478 -667 3512
rect -633 3478 -594 3512
rect -1438 3429 -1308 3468
tri -1040 3440 -1002 3478 se
rect -1002 3440 -594 3478
rect -1438 3395 -1426 3429
rect -1392 3395 -1354 3429
rect -1320 3395 -1308 3429
tri -1074 3406 -1040 3440 se
rect -1040 3406 -886 3440
rect -852 3406 -813 3440
rect -779 3406 -740 3440
rect -706 3406 -667 3440
rect -633 3406 -594 3440
rect 13768 3502 13840 3512
tri 13840 3502 13860 3522 sw
rect 14190 3502 14320 3541
rect 13768 3468 13860 3502
tri 13860 3468 13894 3502 sw
rect 14190 3468 14202 3502
rect 14236 3468 14274 3502
rect 14308 3468 14320 3502
rect 13768 3429 13894 3468
tri 13894 3429 13933 3468 sw
rect 14190 3429 14320 3468
rect 13768 3406 13933 3429
tri -1085 3395 -1074 3406 se
rect -1074 3395 13933 3406
tri 13933 3395 13967 3429 sw
rect 14190 3395 14202 3429
rect 14236 3395 14274 3429
rect 14308 3395 14320 3429
rect -1438 3356 -1308 3395
rect -1438 3322 -1426 3356
rect -1392 3322 -1354 3356
rect -1320 3322 -1308 3356
rect -1438 3283 -1308 3322
rect -1438 3249 -1426 3283
rect -1392 3249 -1354 3283
rect -1320 3249 -1308 3283
rect -1438 3210 -1308 3249
rect -1438 3176 -1426 3210
rect -1392 3176 -1354 3210
rect -1320 3176 -1308 3210
rect -1438 3137 -1308 3176
rect -1438 3103 -1426 3137
rect -1392 3103 -1354 3137
rect -1320 3103 -1308 3137
rect -1438 3064 -1308 3103
rect -1438 3030 -1426 3064
rect -1392 3030 -1354 3064
rect -1320 3030 -1308 3064
rect -1438 2991 -1308 3030
rect -1438 2957 -1426 2991
rect -1392 2957 -1354 2991
rect -1320 2957 -1308 2991
rect -1438 2918 -1308 2957
rect -1438 2884 -1426 2918
rect -1392 2884 -1354 2918
rect -1320 2884 -1308 2918
rect -1438 2845 -1308 2884
rect -1438 2811 -1426 2845
rect -1392 2811 -1354 2845
rect -1320 2811 -1308 2845
rect -1438 2772 -1308 2811
rect -1438 2738 -1426 2772
rect -1392 2738 -1354 2772
rect -1320 2738 -1308 2772
rect -1438 2699 -1308 2738
rect -1438 2665 -1426 2699
rect -1392 2665 -1354 2699
rect -1320 2665 -1308 2699
rect -1438 2626 -1308 2665
rect -1438 2592 -1426 2626
rect -1392 2592 -1354 2626
rect -1320 2592 -1308 2626
rect -1438 2553 -1308 2592
rect -1438 2519 -1426 2553
rect -1392 2519 -1354 2553
rect -1320 2519 -1308 2553
rect -1438 2480 -1308 2519
rect -1438 2446 -1426 2480
rect -1392 2446 -1354 2480
rect -1320 2446 -1308 2480
rect -1438 2407 -1308 2446
rect -1438 2373 -1426 2407
rect -1392 2373 -1354 2407
rect -1320 2373 -1308 2407
rect -1438 2334 -1308 2373
rect -1438 2300 -1426 2334
rect -1392 2300 -1354 2334
rect -1320 2300 -1308 2334
rect -1438 2261 -1308 2300
rect -1438 2227 -1426 2261
rect -1392 2227 -1354 2261
rect -1320 2227 -1308 2261
rect -1438 2188 -1308 2227
rect -1438 2154 -1426 2188
rect -1392 2154 -1354 2188
rect -1320 2154 -1308 2188
rect -1438 2115 -1308 2154
rect -1438 2081 -1426 2115
rect -1392 2081 -1354 2115
rect -1320 2081 -1308 2115
rect -1438 2042 -1308 2081
rect -1438 2008 -1426 2042
rect -1392 2008 -1354 2042
rect -1320 2008 -1308 2042
rect -1438 1969 -1308 2008
rect -1438 1935 -1426 1969
rect -1392 1935 -1354 1969
rect -1320 1935 -1308 1969
rect -1438 1896 -1308 1935
rect -1438 1862 -1426 1896
rect -1392 1862 -1354 1896
rect -1320 1862 -1308 1896
rect -1438 1823 -1308 1862
rect -1438 1789 -1426 1823
rect -1392 1789 -1354 1823
rect -1320 1789 -1308 1823
rect -1438 1750 -1308 1789
rect -1438 1716 -1426 1750
rect -1392 1716 -1354 1750
rect -1320 1716 -1308 1750
rect -1438 1677 -1308 1716
rect -1438 1643 -1426 1677
rect -1392 1643 -1354 1677
rect -1320 1643 -1308 1677
rect -1438 1604 -1308 1643
rect -1438 1570 -1426 1604
rect -1392 1570 -1354 1604
rect -1320 1570 -1308 1604
rect -1438 1531 -1308 1570
rect -1438 1497 -1426 1531
rect -1392 1497 -1354 1531
rect -1320 1497 -1308 1531
rect -1438 1458 -1308 1497
rect -1438 1424 -1426 1458
rect -1392 1424 -1354 1458
rect -1320 1424 -1308 1458
rect -1438 1385 -1308 1424
rect -1438 1351 -1426 1385
rect -1392 1351 -1354 1385
rect -1320 1351 -1308 1385
rect -1438 1312 -1308 1351
rect -1438 1278 -1426 1312
rect -1392 1278 -1354 1312
rect -1320 1278 -1308 1312
rect -1438 1239 -1308 1278
rect -1438 1205 -1426 1239
rect -1392 1205 -1354 1239
rect -1320 1205 -1308 1239
rect -1438 1166 -1308 1205
rect -1438 1132 -1426 1166
rect -1392 1132 -1354 1166
rect -1320 1132 -1308 1166
rect -1438 1093 -1308 1132
rect -1438 1059 -1426 1093
rect -1392 1059 -1354 1093
rect -1320 1059 -1308 1093
rect -1438 1020 -1308 1059
rect -1438 986 -1426 1020
rect -1392 986 -1354 1020
rect -1320 986 -1308 1020
rect -1438 947 -1308 986
rect -1438 913 -1426 947
rect -1392 913 -1354 947
rect -1320 913 -1308 947
rect -1438 874 -1308 913
rect -1438 840 -1426 874
rect -1392 840 -1354 874
rect -1320 840 -1308 874
rect -1438 801 -1308 840
rect -1438 767 -1426 801
rect -1392 767 -1354 801
rect -1320 767 -1308 801
rect -1438 728 -1308 767
rect -1438 694 -1426 728
rect -1392 694 -1354 728
rect -1320 694 -1308 728
rect -1438 655 -1308 694
rect -1438 621 -1426 655
rect -1392 621 -1354 655
rect -1320 621 -1308 655
rect -1438 582 -1308 621
rect -1438 548 -1426 582
rect -1392 548 -1354 582
rect -1320 548 -1308 582
rect -1438 509 -1308 548
rect -1438 475 -1426 509
rect -1392 475 -1354 509
rect -1320 475 -1308 509
rect -1438 436 -1308 475
rect -1438 402 -1426 436
rect -1392 402 -1354 436
rect -1320 402 -1308 436
rect -1438 363 -1308 402
rect -1438 329 -1426 363
rect -1392 329 -1354 363
rect -1320 329 -1308 363
rect -1438 290 -1308 329
rect -1438 256 -1426 290
rect -1392 256 -1354 290
rect -1320 256 -1308 290
rect -1438 217 -1308 256
rect -1438 183 -1426 217
rect -1392 183 -1354 217
rect -1320 183 -1308 217
rect -1438 144 -1308 183
rect -1438 110 -1426 144
rect -1392 110 -1354 144
rect -1320 110 -1308 144
rect -1438 71 -1308 110
rect -1438 37 -1426 71
rect -1392 37 -1354 71
rect -1320 37 -1308 71
rect -1438 -2 -1308 37
rect -1438 -36 -1426 -2
rect -1392 -36 -1354 -2
rect -1320 -36 -1308 -2
rect -1438 -75 -1308 -36
rect -1438 -109 -1426 -75
rect -1392 -109 -1354 -75
rect -1320 -109 -1308 -75
rect -1438 -148 -1308 -109
rect -1438 -182 -1426 -148
rect -1392 -182 -1354 -148
rect -1320 -182 -1308 -148
rect -1438 -221 -1308 -182
rect -1438 -255 -1426 -221
rect -1392 -255 -1354 -221
rect -1320 -255 -1308 -221
rect -1438 -294 -1308 -255
rect -1438 -328 -1426 -294
rect -1392 -328 -1354 -294
rect -1320 -328 -1308 -294
tri -1086 3394 -1085 3395 se
rect -1085 3394 13967 3395
tri 13967 3394 13968 3395 sw
rect -1086 3356 -249 3394
tri -249 3356 -211 3394 nw
tri 13093 3356 13131 3394 ne
rect 13131 3356 13968 3394
rect -1086 3349 -256 3356
tri -256 3349 -249 3356 nw
tri 13131 3349 13138 3356 ne
rect 13138 3349 13968 3356
rect -1086 3322 -283 3349
tri -283 3322 -256 3349 nw
tri 13138 3322 13165 3349 ne
rect 13165 3322 13968 3349
rect -1086 3277 -308 3322
tri -308 3297 -283 3322 nw
tri 13165 3297 13190 3322 ne
rect -1086 2451 -1074 3277
rect -320 2451 -308 3277
rect 13190 3277 13968 3322
rect -1086 2412 -308 2451
rect -1086 2378 -1074 2412
rect -1040 2378 -1002 2412
rect -968 2378 -930 2412
rect -896 2378 -858 2412
rect -824 2378 -786 2412
rect -752 2378 -714 2412
rect -680 2378 -642 2412
rect -608 2378 -570 2412
rect -536 2378 -498 2412
rect -464 2378 -426 2412
rect -392 2378 -354 2412
rect -320 2378 -308 2412
rect -1086 2339 -308 2378
rect -1086 2305 -1074 2339
rect -1040 2305 -1002 2339
rect -968 2305 -930 2339
rect -896 2305 -858 2339
rect -824 2305 -786 2339
rect -752 2305 -714 2339
rect -680 2305 -642 2339
rect -608 2305 -570 2339
rect -536 2305 -498 2339
rect -464 2305 -426 2339
rect -392 2305 -354 2339
rect -320 2305 -308 2339
rect -1086 2266 -308 2305
rect -1086 2232 -1074 2266
rect -1040 2232 -1002 2266
rect -968 2232 -930 2266
rect -896 2232 -858 2266
rect -824 2232 -786 2266
rect -752 2232 -714 2266
rect -680 2232 -642 2266
rect -608 2232 -570 2266
rect -536 2232 -498 2266
rect -464 2232 -426 2266
rect -392 2232 -354 2266
rect -320 2232 -308 2266
rect -1086 2193 -308 2232
rect -1086 2159 -1074 2193
rect -1040 2159 -1002 2193
rect -968 2159 -930 2193
rect -896 2159 -858 2193
rect -824 2159 -786 2193
rect -752 2159 -714 2193
rect -680 2159 -642 2193
rect -608 2159 -570 2193
rect -536 2159 -498 2193
rect -464 2159 -426 2193
rect -392 2159 -354 2193
rect -320 2159 -308 2193
rect -1086 2120 -308 2159
rect -1086 2086 -1074 2120
rect -1040 2086 -1002 2120
rect -968 2086 -930 2120
rect -896 2086 -858 2120
rect -824 2086 -786 2120
rect -752 2086 -714 2120
rect -680 2086 -642 2120
rect -608 2086 -570 2120
rect -536 2086 -498 2120
rect -464 2086 -426 2120
rect -392 2086 -354 2120
rect -320 2086 -308 2120
rect -1086 2047 -308 2086
rect -1086 2013 -1074 2047
rect -1040 2013 -1002 2047
rect -968 2013 -930 2047
rect -896 2013 -858 2047
rect -824 2013 -786 2047
rect -752 2013 -714 2047
rect -680 2013 -642 2047
rect -608 2013 -570 2047
rect -536 2013 -498 2047
rect -464 2013 -426 2047
rect -392 2013 -354 2047
rect -320 2013 -308 2047
rect -1086 1974 -308 2013
rect -1086 1940 -1074 1974
rect -1040 1940 -1002 1974
rect -968 1940 -930 1974
rect -896 1940 -858 1974
rect -824 1940 -786 1974
rect -752 1940 -714 1974
rect -680 1940 -642 1974
rect -608 1940 -570 1974
rect -536 1940 -498 1974
rect -464 1940 -426 1974
rect -392 1940 -354 1974
rect -320 1940 -308 1974
rect -1086 1901 -308 1940
rect -1086 1867 -1074 1901
rect -1040 1867 -1002 1901
rect -968 1867 -930 1901
rect -896 1867 -858 1901
rect -824 1867 -786 1901
rect -752 1867 -714 1901
rect -680 1867 -642 1901
rect -608 1867 -570 1901
rect -536 1867 -498 1901
rect -464 1867 -426 1901
rect -392 1867 -354 1901
rect -320 1867 -308 1901
rect -1086 1828 -308 1867
rect -1086 1794 -1074 1828
rect -1040 1794 -1002 1828
rect -968 1794 -930 1828
rect -896 1794 -858 1828
rect -824 1794 -786 1828
rect -752 1794 -714 1828
rect -680 1794 -642 1828
rect -608 1794 -570 1828
rect -536 1794 -498 1828
rect -464 1794 -426 1828
rect -392 1794 -354 1828
rect -320 1794 -308 1828
rect -1086 1755 -308 1794
rect -1086 1721 -1074 1755
rect -1040 1721 -1002 1755
rect -968 1721 -930 1755
rect -896 1721 -858 1755
rect -824 1721 -786 1755
rect -752 1721 -714 1755
rect -680 1721 -642 1755
rect -608 1721 -570 1755
rect -536 1721 -498 1755
rect -464 1721 -426 1755
rect -392 1721 -354 1755
rect -320 1721 -308 1755
rect -1086 1682 -308 1721
rect -1086 1648 -1074 1682
rect -1040 1648 -1002 1682
rect -968 1648 -930 1682
rect -896 1648 -858 1682
rect -824 1648 -786 1682
rect -752 1648 -714 1682
rect -680 1648 -642 1682
rect -608 1648 -570 1682
rect -536 1648 -498 1682
rect -464 1648 -426 1682
rect -392 1648 -354 1682
rect -320 1648 -308 1682
rect -1086 1609 -308 1648
rect -1086 1575 -1074 1609
rect -1040 1575 -1002 1609
rect -968 1575 -930 1609
rect -896 1575 -858 1609
rect -824 1575 -786 1609
rect -752 1575 -714 1609
rect -680 1575 -642 1609
rect -608 1575 -570 1609
rect -536 1575 -498 1609
rect -464 1575 -426 1609
rect -392 1575 -354 1609
rect -320 1575 -308 1609
rect -1086 1536 -308 1575
rect -1086 1502 -1074 1536
rect -1040 1502 -1002 1536
rect -968 1502 -930 1536
rect -896 1502 -858 1536
rect -824 1502 -786 1536
rect -752 1502 -714 1536
rect -680 1502 -642 1536
rect -608 1502 -570 1536
rect -536 1502 -498 1536
rect -464 1502 -426 1536
rect -392 1502 -354 1536
rect -320 1502 -308 1536
rect -1086 1463 -308 1502
rect -1086 1429 -1074 1463
rect -1040 1429 -1002 1463
rect -968 1429 -930 1463
rect -896 1429 -858 1463
rect -824 1429 -786 1463
rect -752 1429 -714 1463
rect -680 1429 -642 1463
rect -608 1429 -570 1463
rect -536 1429 -498 1463
rect -464 1429 -426 1463
rect -392 1429 -354 1463
rect -320 1429 -308 1463
rect -1086 1390 -308 1429
rect -1086 1356 -1074 1390
rect -1040 1356 -1002 1390
rect -968 1356 -930 1390
rect -896 1356 -858 1390
rect -824 1356 -786 1390
rect -752 1356 -714 1390
rect -680 1356 -642 1390
rect -608 1356 -570 1390
rect -536 1356 -498 1390
rect -464 1356 -426 1390
rect -392 1356 -354 1390
rect -320 1356 -308 1390
rect -1086 1317 -308 1356
rect -1086 1283 -1074 1317
rect -1040 1283 -1002 1317
rect -968 1283 -930 1317
rect -896 1283 -858 1317
rect -824 1283 -786 1317
rect -752 1283 -714 1317
rect -680 1283 -642 1317
rect -608 1283 -570 1317
rect -536 1283 -498 1317
rect -464 1283 -426 1317
rect -392 1283 -354 1317
rect -320 1283 -308 1317
rect -1086 1244 -308 1283
rect -1086 1210 -1074 1244
rect -1040 1210 -1002 1244
rect -968 1210 -930 1244
rect -896 1210 -858 1244
rect -824 1210 -786 1244
rect -752 1210 -714 1244
rect -680 1210 -642 1244
rect -608 1210 -570 1244
rect -536 1210 -498 1244
rect -464 1210 -426 1244
rect -392 1210 -354 1244
rect -320 1210 -308 1244
rect -1086 1171 -308 1210
rect -1086 1137 -1074 1171
rect -1040 1137 -1002 1171
rect -968 1137 -930 1171
rect -896 1137 -858 1171
rect -824 1137 -786 1171
rect -752 1137 -714 1171
rect -680 1137 -642 1171
rect -608 1137 -570 1171
rect -536 1137 -498 1171
rect -464 1137 -426 1171
rect -392 1137 -354 1171
rect -320 1137 -308 1171
rect -1086 1098 -308 1137
rect -1086 1064 -1074 1098
rect -1040 1064 -1002 1098
rect -968 1064 -930 1098
rect -896 1064 -858 1098
rect -824 1064 -786 1098
rect -752 1064 -714 1098
rect -680 1064 -642 1098
rect -608 1064 -570 1098
rect -536 1064 -498 1098
rect -464 1064 -426 1098
rect -392 1064 -354 1098
rect -320 1064 -308 1098
rect -1086 1025 -308 1064
rect -1086 991 -1074 1025
rect -1040 991 -1002 1025
rect -968 991 -930 1025
rect -896 991 -858 1025
rect -824 991 -786 1025
rect -752 991 -714 1025
rect -680 991 -642 1025
rect -608 991 -570 1025
rect -536 991 -498 1025
rect -464 991 -426 1025
rect -392 991 -354 1025
rect -320 991 -308 1025
rect -1086 952 -308 991
rect -1086 918 -1074 952
rect -1040 918 -1002 952
rect -968 918 -930 952
rect -896 918 -858 952
rect -824 918 -786 952
rect -752 918 -714 952
rect -680 918 -642 952
rect -608 918 -570 952
rect -536 918 -498 952
rect -464 918 -426 952
rect -392 918 -354 952
rect -320 918 -308 952
rect -1086 879 -308 918
rect -1086 845 -1074 879
rect -1040 845 -1002 879
rect -968 845 -930 879
rect -896 845 -858 879
rect -824 845 -786 879
rect -752 845 -714 879
rect -680 845 -642 879
rect -608 845 -570 879
rect -536 845 -498 879
rect -464 845 -426 879
rect -392 845 -354 879
rect -320 845 -308 879
rect -1086 806 -308 845
rect -1086 772 -1074 806
rect -1040 772 -1002 806
rect -968 772 -930 806
rect -896 772 -858 806
rect -824 772 -786 806
rect -752 772 -714 806
rect -680 772 -642 806
rect -608 772 -570 806
rect -536 772 -498 806
rect -464 772 -426 806
rect -392 772 -354 806
rect -320 772 -308 806
rect -1086 733 -308 772
rect -1086 699 -1074 733
rect -1040 699 -1002 733
rect -968 699 -930 733
rect -896 699 -858 733
rect -824 699 -786 733
rect -752 699 -714 733
rect -680 699 -642 733
rect -608 699 -570 733
rect -536 699 -498 733
rect -464 699 -426 733
rect -392 699 -354 733
rect -320 699 -308 733
rect -1086 660 -308 699
rect -1086 626 -1074 660
rect -1040 626 -1002 660
rect -968 626 -930 660
rect -896 626 -858 660
rect -824 626 -786 660
rect -752 626 -714 660
rect -680 626 -642 660
rect -608 626 -570 660
rect -536 626 -498 660
rect -464 626 -426 660
rect -392 626 -354 660
rect -320 626 -308 660
rect -1086 587 -308 626
rect -1086 553 -1074 587
rect -1040 553 -1002 587
rect -968 553 -930 587
rect -896 553 -858 587
rect -824 553 -786 587
rect -752 553 -714 587
rect -680 553 -642 587
rect -608 553 -570 587
rect -536 553 -498 587
rect -464 553 -426 587
rect -392 553 -354 587
rect -320 553 -308 587
rect -1086 514 -308 553
rect -1086 480 -1074 514
rect -1040 480 -1002 514
rect -968 480 -930 514
rect -896 480 -858 514
rect -824 480 -786 514
rect -752 480 -714 514
rect -680 480 -642 514
rect -608 480 -570 514
rect -536 480 -498 514
rect -464 480 -426 514
rect -392 480 -354 514
rect -320 480 -308 514
rect -1086 441 -308 480
rect -1086 407 -1074 441
rect -1040 407 -1002 441
rect -968 407 -930 441
rect -896 407 -858 441
rect -824 407 -786 441
rect -752 407 -714 441
rect -680 407 -642 441
rect -608 407 -570 441
rect -536 407 -498 441
rect -464 407 -426 441
rect -392 407 -354 441
rect -320 407 -308 441
rect -1086 368 -308 407
rect -1086 334 -1074 368
rect -1040 334 -1002 368
rect -968 334 -930 368
rect -896 334 -858 368
rect -824 334 -786 368
rect -752 334 -714 368
rect -680 334 -642 368
rect -608 334 -570 368
rect -536 334 -498 368
rect -464 334 -426 368
rect -392 334 -354 368
rect -320 334 -308 368
rect -1086 295 -308 334
rect -1086 261 -1074 295
rect -1040 261 -1002 295
rect -968 261 -930 295
rect -896 261 -858 295
rect -824 261 -786 295
rect -752 261 -714 295
rect -680 261 -642 295
rect -608 261 -570 295
rect -536 261 -498 295
rect -464 261 -426 295
rect -392 261 -354 295
rect -320 261 -308 295
rect -1086 222 -308 261
rect -1086 188 -1074 222
rect -1040 188 -1002 222
rect -968 188 -930 222
rect -896 188 -858 222
rect -824 188 -786 222
rect -752 188 -714 222
rect -680 188 -642 222
rect -608 188 -570 222
rect -536 188 -498 222
rect -464 188 -426 222
rect -392 188 -354 222
rect -320 188 -308 222
rect -1086 149 -308 188
rect -1086 115 -1074 149
rect -1040 115 -1002 149
rect -968 115 -930 149
rect -896 115 -858 149
rect -824 115 -786 149
rect -752 115 -714 149
rect -680 115 -642 149
rect -608 115 -570 149
rect -536 115 -498 149
rect -464 115 -426 149
rect -392 115 -354 149
rect -320 115 -308 149
rect -1086 76 -308 115
rect -1086 42 -1074 76
rect -1040 42 -1002 76
rect -968 42 -930 76
rect -896 42 -858 76
rect -824 42 -786 76
rect -752 42 -714 76
rect -680 42 -642 76
rect -608 42 -570 76
rect -536 42 -498 76
rect -464 42 -426 76
rect -392 42 -354 76
rect -320 42 -308 76
tri -251 3053 -204 3100 se
rect -204 3053 -98 3100
tri -98 3053 -51 3100 sw
rect -251 3000 -51 3053
rect -251 2966 -204 3000
rect -170 2966 -132 3000
rect -98 2966 -51 3000
rect -251 2927 -51 2966
rect -251 2893 -204 2927
rect -170 2893 -132 2927
rect -98 2893 -51 2927
rect -251 2854 -51 2893
rect -251 2820 -204 2854
rect -170 2820 -132 2854
rect -98 2820 -51 2854
rect -251 2781 -51 2820
rect -251 2747 -204 2781
rect -170 2747 -132 2781
rect -98 2747 -51 2781
rect -251 2708 -51 2747
rect -251 2674 -204 2708
rect -170 2674 -132 2708
rect -98 2674 -51 2708
rect -251 2635 -51 2674
rect -251 2601 -204 2635
rect -170 2601 -132 2635
rect -98 2601 -51 2635
rect -251 2562 -51 2601
rect -251 2528 -204 2562
rect -170 2528 -132 2562
rect -98 2528 -51 2562
rect -251 2489 -51 2528
rect -251 2455 -204 2489
rect -170 2455 -132 2489
rect -98 2455 -51 2489
rect -251 2416 -51 2455
rect -251 2382 -204 2416
rect -170 2382 -132 2416
rect -98 2382 -51 2416
rect -251 2343 -51 2382
rect -251 2309 -204 2343
rect -170 2309 -132 2343
rect -98 2309 -51 2343
rect -251 2270 -51 2309
rect -251 2236 -204 2270
rect -170 2236 -132 2270
rect -98 2236 -51 2270
rect -251 2197 -51 2236
rect -251 2163 -204 2197
rect -170 2163 -132 2197
rect -98 2163 -51 2197
rect -251 2124 -51 2163
rect -251 2090 -204 2124
rect -170 2090 -132 2124
rect -98 2090 -51 2124
rect -251 2051 -51 2090
rect -251 2017 -204 2051
rect -170 2017 -132 2051
rect -98 2017 -51 2051
rect -251 1978 -51 2017
rect -251 1944 -204 1978
rect -170 1944 -132 1978
rect -98 1944 -51 1978
rect -251 1905 -51 1944
rect -251 1871 -204 1905
rect -170 1871 -132 1905
rect -98 1871 -51 1905
rect -251 1832 -51 1871
rect -251 1798 -204 1832
rect -170 1798 -132 1832
rect -98 1798 -51 1832
rect -251 1759 -51 1798
rect -251 1725 -204 1759
rect -170 1725 -132 1759
rect -98 1725 -51 1759
rect -251 1686 -51 1725
rect -251 1652 -204 1686
rect -170 1652 -132 1686
rect -98 1652 -51 1686
rect -251 1613 -51 1652
rect -251 1579 -204 1613
rect -170 1579 -132 1613
rect -98 1579 -51 1613
rect -251 1540 -51 1579
rect -251 1506 -204 1540
rect -170 1506 -132 1540
rect -98 1506 -51 1540
rect -251 1466 -51 1506
rect -251 1432 -204 1466
rect -170 1432 -132 1466
rect -98 1432 -51 1466
rect -251 1392 -51 1432
rect -251 1358 -204 1392
rect -170 1358 -132 1392
rect -98 1358 -51 1392
rect -251 1318 -51 1358
rect -251 1284 -204 1318
rect -170 1284 -132 1318
rect -98 1284 -51 1318
rect -251 1244 -51 1284
rect -251 1210 -204 1244
rect -170 1210 -132 1244
rect -98 1210 -51 1244
rect -251 1170 -51 1210
rect -251 1136 -204 1170
rect -170 1136 -132 1170
rect -98 1136 -51 1170
rect -251 1096 -51 1136
rect -251 1062 -204 1096
rect -170 1062 -132 1096
rect -98 1062 -51 1096
rect -251 1022 -51 1062
rect -251 988 -204 1022
rect -170 988 -132 1022
rect -98 988 -51 1022
rect -251 948 -51 988
rect -251 914 -204 948
rect -170 914 -132 948
rect -98 914 -51 948
rect -251 874 -51 914
rect -251 840 -204 874
rect -170 840 -132 874
rect -98 840 -51 874
rect -251 800 -51 840
rect -251 766 -204 800
rect -170 766 -132 800
rect -98 766 -51 800
rect -251 726 -51 766
rect -251 692 -204 726
rect -170 692 -132 726
rect -98 692 -51 726
rect -251 652 -51 692
rect -251 618 -204 652
rect -170 618 -132 652
rect -98 618 -51 652
rect -251 578 -51 618
rect -251 544 -204 578
rect -170 544 -132 578
rect -98 544 -51 578
rect -251 504 -51 544
rect -251 470 -204 504
rect -170 470 -132 504
rect -98 470 -51 504
rect -251 430 -51 470
rect -251 396 -204 430
rect -170 396 -132 430
rect -98 396 -51 430
rect -251 356 -51 396
rect -251 322 -204 356
rect -170 322 -132 356
rect -98 322 -51 356
rect -251 282 -51 322
rect -251 248 -204 282
rect -170 248 -132 282
rect -98 248 -51 282
rect -251 208 -51 248
rect -251 174 -204 208
rect -170 174 -132 208
rect -98 174 -51 208
rect -251 134 -51 174
rect -251 100 -204 134
rect -170 100 -132 134
rect -98 100 -51 134
rect -251 47 -51 100
tri -251 42 -246 47 ne
rect -246 42 -56 47
tri -56 42 -51 47 nw
tri 61 3053 108 3100 se
rect 108 3053 414 3100
tri 414 3053 461 3100 sw
rect 61 3000 461 3053
rect 61 2966 208 3000
rect 242 2966 280 3000
rect 314 2966 461 3000
rect 61 2927 461 2966
rect 61 2893 208 2927
rect 242 2893 280 2927
rect 314 2893 461 2927
rect 61 2854 461 2893
rect 61 2820 208 2854
rect 242 2820 280 2854
rect 314 2820 461 2854
rect 61 2781 461 2820
rect 61 2747 208 2781
rect 242 2747 280 2781
rect 314 2747 461 2781
rect 61 2708 461 2747
rect 61 2674 208 2708
rect 242 2674 280 2708
rect 314 2674 461 2708
rect 61 2635 461 2674
rect 61 2601 208 2635
rect 242 2601 280 2635
rect 314 2601 461 2635
rect 61 2562 461 2601
rect 61 2528 208 2562
rect 242 2528 280 2562
rect 314 2528 461 2562
rect 61 2489 461 2528
rect 61 2455 208 2489
rect 242 2455 280 2489
rect 314 2455 461 2489
rect 61 2416 461 2455
rect 61 2382 208 2416
rect 242 2382 280 2416
rect 314 2382 461 2416
rect 61 2343 461 2382
rect 61 2309 208 2343
rect 242 2309 280 2343
rect 314 2309 461 2343
rect 61 2270 461 2309
rect 61 2236 208 2270
rect 242 2236 280 2270
rect 314 2236 461 2270
rect 61 2197 461 2236
rect 61 2163 208 2197
rect 242 2163 280 2197
rect 314 2163 461 2197
rect 61 2124 461 2163
rect 61 2090 208 2124
rect 242 2090 280 2124
rect 314 2090 461 2124
rect 61 2051 461 2090
rect 61 2017 208 2051
rect 242 2017 280 2051
rect 314 2017 461 2051
rect 61 1978 461 2017
rect 61 1944 208 1978
rect 242 1944 280 1978
rect 314 1944 461 1978
rect 61 1905 461 1944
rect 61 1871 208 1905
rect 242 1871 280 1905
rect 314 1871 461 1905
rect 61 1832 461 1871
rect 61 1798 208 1832
rect 242 1798 280 1832
rect 314 1798 461 1832
rect 61 1759 461 1798
rect 61 1725 208 1759
rect 242 1725 280 1759
rect 314 1725 461 1759
rect 61 1686 461 1725
rect 61 1652 208 1686
rect 242 1652 280 1686
rect 314 1652 461 1686
rect 61 1613 461 1652
rect 61 1579 208 1613
rect 242 1579 280 1613
rect 314 1579 461 1613
rect 61 1540 461 1579
rect 61 1506 208 1540
rect 242 1506 280 1540
rect 314 1506 461 1540
rect 61 1466 461 1506
rect 61 1432 208 1466
rect 242 1432 280 1466
rect 314 1432 461 1466
rect 61 1392 461 1432
rect 61 1358 208 1392
rect 242 1358 280 1392
rect 314 1358 461 1392
rect 61 1318 461 1358
rect 61 1284 208 1318
rect 242 1284 280 1318
rect 314 1284 461 1318
rect 61 1244 461 1284
rect 61 1210 208 1244
rect 242 1210 280 1244
rect 314 1210 461 1244
rect 61 1170 461 1210
rect 61 1136 208 1170
rect 242 1136 280 1170
rect 314 1136 461 1170
rect 61 1096 461 1136
rect 61 1062 208 1096
rect 242 1062 280 1096
rect 314 1062 461 1096
rect 61 1022 461 1062
rect 61 988 208 1022
rect 242 988 280 1022
rect 314 988 461 1022
rect 61 948 461 988
rect 61 914 208 948
rect 242 914 280 948
rect 314 914 461 948
rect 61 874 461 914
rect 61 840 208 874
rect 242 840 280 874
rect 314 840 461 874
rect 61 800 461 840
rect 61 766 208 800
rect 242 766 280 800
rect 314 766 461 800
rect 61 726 461 766
rect 61 692 208 726
rect 242 692 280 726
rect 314 692 461 726
rect 61 652 461 692
rect 61 618 208 652
rect 242 618 280 652
rect 314 618 461 652
rect 61 578 461 618
rect 61 544 208 578
rect 242 544 280 578
rect 314 544 461 578
rect 61 504 461 544
rect 61 470 208 504
rect 242 470 280 504
rect 314 470 461 504
rect 61 430 461 470
rect 61 396 208 430
rect 242 396 280 430
rect 314 396 461 430
rect 61 356 461 396
rect 61 322 208 356
rect 242 322 280 356
rect 314 322 461 356
rect 61 282 461 322
rect 61 248 208 282
rect 242 248 280 282
rect 314 248 461 282
rect 61 208 461 248
rect 61 174 208 208
rect 242 174 280 208
rect 314 174 461 208
rect 61 134 461 174
rect 61 100 208 134
rect 242 100 280 134
rect 314 100 461 134
rect 61 47 461 100
tri 61 42 66 47 ne
rect 66 42 456 47
tri 456 42 461 47 nw
tri 573 3053 620 3100 se
rect 620 3053 726 3100
tri 726 3053 773 3100 sw
rect 573 3000 773 3053
rect 573 2966 620 3000
rect 654 2966 692 3000
rect 726 2966 773 3000
rect 573 2927 773 2966
rect 573 2893 620 2927
rect 654 2893 692 2927
rect 726 2893 773 2927
rect 573 2854 773 2893
rect 573 2820 620 2854
rect 654 2820 692 2854
rect 726 2820 773 2854
rect 573 2781 773 2820
rect 573 2747 620 2781
rect 654 2747 692 2781
rect 726 2747 773 2781
rect 573 2708 773 2747
rect 573 2674 620 2708
rect 654 2674 692 2708
rect 726 2674 773 2708
rect 573 2635 773 2674
rect 573 2601 620 2635
rect 654 2601 692 2635
rect 726 2601 773 2635
rect 573 2562 773 2601
rect 573 2528 620 2562
rect 654 2528 692 2562
rect 726 2528 773 2562
rect 573 2489 773 2528
rect 573 2455 620 2489
rect 654 2455 692 2489
rect 726 2455 773 2489
rect 573 2416 773 2455
rect 573 2382 620 2416
rect 654 2382 692 2416
rect 726 2382 773 2416
rect 573 2343 773 2382
rect 573 2309 620 2343
rect 654 2309 692 2343
rect 726 2309 773 2343
rect 573 2270 773 2309
rect 573 2236 620 2270
rect 654 2236 692 2270
rect 726 2236 773 2270
rect 573 2197 773 2236
rect 573 2163 620 2197
rect 654 2163 692 2197
rect 726 2163 773 2197
rect 573 2124 773 2163
rect 573 2090 620 2124
rect 654 2090 692 2124
rect 726 2090 773 2124
rect 573 2051 773 2090
rect 573 2017 620 2051
rect 654 2017 692 2051
rect 726 2017 773 2051
rect 573 1978 773 2017
rect 573 1944 620 1978
rect 654 1944 692 1978
rect 726 1944 773 1978
rect 573 1905 773 1944
rect 573 1871 620 1905
rect 654 1871 692 1905
rect 726 1871 773 1905
rect 573 1832 773 1871
rect 573 1798 620 1832
rect 654 1798 692 1832
rect 726 1798 773 1832
rect 573 1759 773 1798
rect 573 1725 620 1759
rect 654 1725 692 1759
rect 726 1725 773 1759
rect 573 1686 773 1725
rect 573 1652 620 1686
rect 654 1652 692 1686
rect 726 1652 773 1686
rect 573 1613 773 1652
rect 573 1579 620 1613
rect 654 1579 692 1613
rect 726 1579 773 1613
rect 573 1540 773 1579
rect 573 1506 620 1540
rect 654 1506 692 1540
rect 726 1506 773 1540
rect 573 1466 773 1506
rect 573 1432 620 1466
rect 654 1432 692 1466
rect 726 1432 773 1466
rect 573 1392 773 1432
rect 573 1358 620 1392
rect 654 1358 692 1392
rect 726 1358 773 1392
rect 573 1318 773 1358
rect 573 1284 620 1318
rect 654 1284 692 1318
rect 726 1284 773 1318
rect 573 1244 773 1284
rect 573 1210 620 1244
rect 654 1210 692 1244
rect 726 1210 773 1244
rect 573 1170 773 1210
rect 573 1136 620 1170
rect 654 1136 692 1170
rect 726 1136 773 1170
rect 573 1096 773 1136
rect 573 1062 620 1096
rect 654 1062 692 1096
rect 726 1062 773 1096
rect 573 1022 773 1062
rect 573 988 620 1022
rect 654 988 692 1022
rect 726 988 773 1022
rect 573 948 773 988
rect 573 914 620 948
rect 654 914 692 948
rect 726 914 773 948
rect 573 874 773 914
rect 573 840 620 874
rect 654 840 692 874
rect 726 840 773 874
rect 573 800 773 840
rect 573 766 620 800
rect 654 766 692 800
rect 726 766 773 800
rect 573 726 773 766
rect 573 692 620 726
rect 654 692 692 726
rect 726 692 773 726
rect 573 652 773 692
rect 573 618 620 652
rect 654 618 692 652
rect 726 618 773 652
rect 573 578 773 618
rect 573 544 620 578
rect 654 544 692 578
rect 726 544 773 578
rect 573 504 773 544
rect 573 470 620 504
rect 654 470 692 504
rect 726 470 773 504
rect 573 430 773 470
rect 573 396 620 430
rect 654 396 692 430
rect 726 396 773 430
rect 573 356 773 396
rect 573 322 620 356
rect 654 322 692 356
rect 726 322 773 356
rect 573 282 773 322
rect 573 248 620 282
rect 654 248 692 282
rect 726 248 773 282
rect 573 208 773 248
rect 573 174 620 208
rect 654 174 692 208
rect 726 174 773 208
rect 573 134 773 174
rect 573 100 620 134
rect 654 100 692 134
rect 726 100 773 134
rect 573 47 773 100
tri 573 42 578 47 ne
rect 578 42 768 47
tri 768 42 773 47 nw
tri 885 3053 932 3100 se
rect 932 3053 1238 3100
tri 1238 3053 1285 3100 sw
rect 885 3000 1285 3053
rect 885 2966 1032 3000
rect 1066 2966 1104 3000
rect 1138 2966 1285 3000
rect 885 2927 1285 2966
rect 885 2893 1032 2927
rect 1066 2893 1104 2927
rect 1138 2893 1285 2927
rect 885 2854 1285 2893
rect 885 2820 1032 2854
rect 1066 2820 1104 2854
rect 1138 2820 1285 2854
rect 885 2781 1285 2820
rect 885 2747 1032 2781
rect 1066 2747 1104 2781
rect 1138 2747 1285 2781
rect 885 2708 1285 2747
rect 885 2674 1032 2708
rect 1066 2674 1104 2708
rect 1138 2674 1285 2708
rect 885 2635 1285 2674
rect 885 2601 1032 2635
rect 1066 2601 1104 2635
rect 1138 2601 1285 2635
rect 885 2562 1285 2601
rect 885 2528 1032 2562
rect 1066 2528 1104 2562
rect 1138 2528 1285 2562
rect 885 2489 1285 2528
rect 885 2455 1032 2489
rect 1066 2455 1104 2489
rect 1138 2455 1285 2489
rect 885 2416 1285 2455
rect 885 2382 1032 2416
rect 1066 2382 1104 2416
rect 1138 2382 1285 2416
rect 885 2343 1285 2382
rect 885 2309 1032 2343
rect 1066 2309 1104 2343
rect 1138 2309 1285 2343
rect 885 2270 1285 2309
rect 885 2236 1032 2270
rect 1066 2236 1104 2270
rect 1138 2236 1285 2270
rect 885 2197 1285 2236
rect 885 2163 1032 2197
rect 1066 2163 1104 2197
rect 1138 2163 1285 2197
rect 885 2124 1285 2163
rect 885 2090 1032 2124
rect 1066 2090 1104 2124
rect 1138 2090 1285 2124
rect 885 2051 1285 2090
rect 885 2017 1032 2051
rect 1066 2017 1104 2051
rect 1138 2017 1285 2051
rect 885 1978 1285 2017
rect 885 1944 1032 1978
rect 1066 1944 1104 1978
rect 1138 1944 1285 1978
rect 885 1905 1285 1944
rect 885 1871 1032 1905
rect 1066 1871 1104 1905
rect 1138 1871 1285 1905
rect 885 1832 1285 1871
rect 885 1798 1032 1832
rect 1066 1798 1104 1832
rect 1138 1798 1285 1832
rect 885 1759 1285 1798
rect 885 1725 1032 1759
rect 1066 1725 1104 1759
rect 1138 1725 1285 1759
rect 885 1686 1285 1725
rect 885 1652 1032 1686
rect 1066 1652 1104 1686
rect 1138 1652 1285 1686
rect 885 1613 1285 1652
rect 885 1579 1032 1613
rect 1066 1579 1104 1613
rect 1138 1579 1285 1613
rect 885 1540 1285 1579
rect 885 1506 1032 1540
rect 1066 1506 1104 1540
rect 1138 1506 1285 1540
rect 885 1466 1285 1506
rect 885 1432 1032 1466
rect 1066 1432 1104 1466
rect 1138 1432 1285 1466
rect 885 1392 1285 1432
rect 885 1358 1032 1392
rect 1066 1358 1104 1392
rect 1138 1358 1285 1392
rect 885 1318 1285 1358
rect 885 1284 1032 1318
rect 1066 1284 1104 1318
rect 1138 1284 1285 1318
rect 885 1244 1285 1284
rect 885 1210 1032 1244
rect 1066 1210 1104 1244
rect 1138 1210 1285 1244
rect 885 1170 1285 1210
rect 885 1136 1032 1170
rect 1066 1136 1104 1170
rect 1138 1136 1285 1170
rect 885 1096 1285 1136
rect 885 1062 1032 1096
rect 1066 1062 1104 1096
rect 1138 1062 1285 1096
rect 885 1022 1285 1062
rect 885 988 1032 1022
rect 1066 988 1104 1022
rect 1138 988 1285 1022
rect 885 948 1285 988
rect 885 914 1032 948
rect 1066 914 1104 948
rect 1138 914 1285 948
rect 885 874 1285 914
rect 885 840 1032 874
rect 1066 840 1104 874
rect 1138 840 1285 874
rect 885 800 1285 840
rect 885 766 1032 800
rect 1066 766 1104 800
rect 1138 766 1285 800
rect 885 726 1285 766
rect 885 692 1032 726
rect 1066 692 1104 726
rect 1138 692 1285 726
rect 885 652 1285 692
rect 885 618 1032 652
rect 1066 618 1104 652
rect 1138 618 1285 652
rect 885 578 1285 618
rect 885 544 1032 578
rect 1066 544 1104 578
rect 1138 544 1285 578
rect 885 504 1285 544
rect 885 470 1032 504
rect 1066 470 1104 504
rect 1138 470 1285 504
rect 885 430 1285 470
rect 885 396 1032 430
rect 1066 396 1104 430
rect 1138 396 1285 430
rect 885 356 1285 396
rect 885 322 1032 356
rect 1066 322 1104 356
rect 1138 322 1285 356
rect 885 282 1285 322
rect 885 248 1032 282
rect 1066 248 1104 282
rect 1138 248 1285 282
rect 885 208 1285 248
rect 885 174 1032 208
rect 1066 174 1104 208
rect 1138 174 1285 208
rect 885 134 1285 174
rect 885 100 1032 134
rect 1066 100 1104 134
rect 1138 100 1285 134
rect 885 47 1285 100
tri 885 42 890 47 ne
rect 890 42 1280 47
tri 1280 42 1285 47 nw
tri 1397 3053 1444 3100 se
rect 1444 3053 1550 3100
tri 1550 3053 1597 3100 sw
rect 1397 3000 1597 3053
rect 1397 2966 1444 3000
rect 1478 2966 1516 3000
rect 1550 2966 1597 3000
rect 1397 2927 1597 2966
rect 1397 2893 1444 2927
rect 1478 2893 1516 2927
rect 1550 2893 1597 2927
rect 1397 2854 1597 2893
rect 1397 2820 1444 2854
rect 1478 2820 1516 2854
rect 1550 2820 1597 2854
rect 1397 2781 1597 2820
rect 1397 2747 1444 2781
rect 1478 2747 1516 2781
rect 1550 2747 1597 2781
rect 1397 2708 1597 2747
rect 1397 2674 1444 2708
rect 1478 2674 1516 2708
rect 1550 2674 1597 2708
rect 1397 2635 1597 2674
rect 1397 2601 1444 2635
rect 1478 2601 1516 2635
rect 1550 2601 1597 2635
rect 1397 2562 1597 2601
rect 1397 2528 1444 2562
rect 1478 2528 1516 2562
rect 1550 2528 1597 2562
rect 1397 2489 1597 2528
rect 1397 2455 1444 2489
rect 1478 2455 1516 2489
rect 1550 2455 1597 2489
rect 1397 2416 1597 2455
rect 1397 2382 1444 2416
rect 1478 2382 1516 2416
rect 1550 2382 1597 2416
rect 1397 2343 1597 2382
rect 1397 2309 1444 2343
rect 1478 2309 1516 2343
rect 1550 2309 1597 2343
rect 1397 2270 1597 2309
rect 1397 2236 1444 2270
rect 1478 2236 1516 2270
rect 1550 2236 1597 2270
rect 1397 2197 1597 2236
rect 1397 2163 1444 2197
rect 1478 2163 1516 2197
rect 1550 2163 1597 2197
rect 1397 2124 1597 2163
rect 1397 2090 1444 2124
rect 1478 2090 1516 2124
rect 1550 2090 1597 2124
rect 1397 2051 1597 2090
rect 1397 2017 1444 2051
rect 1478 2017 1516 2051
rect 1550 2017 1597 2051
rect 1397 1978 1597 2017
rect 1397 1944 1444 1978
rect 1478 1944 1516 1978
rect 1550 1944 1597 1978
rect 1397 1905 1597 1944
rect 1397 1871 1444 1905
rect 1478 1871 1516 1905
rect 1550 1871 1597 1905
rect 1397 1832 1597 1871
rect 1397 1798 1444 1832
rect 1478 1798 1516 1832
rect 1550 1798 1597 1832
rect 1397 1759 1597 1798
rect 1397 1725 1444 1759
rect 1478 1725 1516 1759
rect 1550 1725 1597 1759
rect 1397 1686 1597 1725
rect 1397 1652 1444 1686
rect 1478 1652 1516 1686
rect 1550 1652 1597 1686
rect 1397 1613 1597 1652
rect 1397 1579 1444 1613
rect 1478 1579 1516 1613
rect 1550 1579 1597 1613
rect 1397 1540 1597 1579
rect 1397 1506 1444 1540
rect 1478 1506 1516 1540
rect 1550 1506 1597 1540
rect 1397 1466 1597 1506
rect 1397 1432 1444 1466
rect 1478 1432 1516 1466
rect 1550 1432 1597 1466
rect 1397 1392 1597 1432
rect 1397 1358 1444 1392
rect 1478 1358 1516 1392
rect 1550 1358 1597 1392
rect 1397 1318 1597 1358
rect 1397 1284 1444 1318
rect 1478 1284 1516 1318
rect 1550 1284 1597 1318
rect 1397 1244 1597 1284
rect 1397 1210 1444 1244
rect 1478 1210 1516 1244
rect 1550 1210 1597 1244
rect 1397 1170 1597 1210
rect 1397 1136 1444 1170
rect 1478 1136 1516 1170
rect 1550 1136 1597 1170
rect 1397 1096 1597 1136
rect 1397 1062 1444 1096
rect 1478 1062 1516 1096
rect 1550 1062 1597 1096
rect 1397 1022 1597 1062
rect 1397 988 1444 1022
rect 1478 988 1516 1022
rect 1550 988 1597 1022
rect 1397 948 1597 988
rect 1397 914 1444 948
rect 1478 914 1516 948
rect 1550 914 1597 948
rect 1397 874 1597 914
rect 1397 840 1444 874
rect 1478 840 1516 874
rect 1550 840 1597 874
rect 1397 800 1597 840
rect 1397 766 1444 800
rect 1478 766 1516 800
rect 1550 766 1597 800
rect 1397 726 1597 766
rect 1397 692 1444 726
rect 1478 692 1516 726
rect 1550 692 1597 726
rect 1397 652 1597 692
rect 1397 618 1444 652
rect 1478 618 1516 652
rect 1550 618 1597 652
rect 1397 578 1597 618
rect 1397 544 1444 578
rect 1478 544 1516 578
rect 1550 544 1597 578
rect 1397 504 1597 544
rect 1397 470 1444 504
rect 1478 470 1516 504
rect 1550 470 1597 504
rect 1397 430 1597 470
rect 1397 396 1444 430
rect 1478 396 1516 430
rect 1550 396 1597 430
rect 1397 356 1597 396
rect 1397 322 1444 356
rect 1478 322 1516 356
rect 1550 322 1597 356
rect 1397 282 1597 322
rect 1397 248 1444 282
rect 1478 248 1516 282
rect 1550 248 1597 282
rect 1397 208 1597 248
rect 1397 174 1444 208
rect 1478 174 1516 208
rect 1550 174 1597 208
rect 1397 134 1597 174
rect 1397 100 1444 134
rect 1478 100 1516 134
rect 1550 100 1597 134
rect 1397 47 1597 100
tri 1397 42 1402 47 ne
rect 1402 42 1592 47
tri 1592 42 1597 47 nw
tri 1709 3053 1756 3100 se
rect 1756 3053 2062 3100
tri 2062 3053 2109 3100 sw
rect 1709 3000 2109 3053
rect 1709 2966 1856 3000
rect 1890 2966 1928 3000
rect 1962 2966 2109 3000
rect 1709 2927 2109 2966
rect 1709 2893 1856 2927
rect 1890 2893 1928 2927
rect 1962 2893 2109 2927
rect 1709 2854 2109 2893
rect 1709 2820 1856 2854
rect 1890 2820 1928 2854
rect 1962 2820 2109 2854
rect 1709 2781 2109 2820
rect 1709 2747 1856 2781
rect 1890 2747 1928 2781
rect 1962 2747 2109 2781
rect 1709 2708 2109 2747
rect 1709 2674 1856 2708
rect 1890 2674 1928 2708
rect 1962 2674 2109 2708
rect 1709 2635 2109 2674
rect 1709 2601 1856 2635
rect 1890 2601 1928 2635
rect 1962 2601 2109 2635
rect 1709 2562 2109 2601
rect 1709 2528 1856 2562
rect 1890 2528 1928 2562
rect 1962 2528 2109 2562
rect 1709 2489 2109 2528
rect 1709 2455 1856 2489
rect 1890 2455 1928 2489
rect 1962 2455 2109 2489
rect 1709 2416 2109 2455
rect 1709 2382 1856 2416
rect 1890 2382 1928 2416
rect 1962 2382 2109 2416
rect 1709 2343 2109 2382
rect 1709 2309 1856 2343
rect 1890 2309 1928 2343
rect 1962 2309 2109 2343
rect 1709 2270 2109 2309
rect 1709 2236 1856 2270
rect 1890 2236 1928 2270
rect 1962 2236 2109 2270
rect 1709 2197 2109 2236
rect 1709 2163 1856 2197
rect 1890 2163 1928 2197
rect 1962 2163 2109 2197
rect 1709 2124 2109 2163
rect 1709 2090 1856 2124
rect 1890 2090 1928 2124
rect 1962 2090 2109 2124
rect 1709 2051 2109 2090
rect 1709 2017 1856 2051
rect 1890 2017 1928 2051
rect 1962 2017 2109 2051
rect 1709 1978 2109 2017
rect 1709 1944 1856 1978
rect 1890 1944 1928 1978
rect 1962 1944 2109 1978
rect 1709 1905 2109 1944
rect 1709 1871 1856 1905
rect 1890 1871 1928 1905
rect 1962 1871 2109 1905
rect 1709 1832 2109 1871
rect 1709 1798 1856 1832
rect 1890 1798 1928 1832
rect 1962 1798 2109 1832
rect 1709 1759 2109 1798
rect 1709 1725 1856 1759
rect 1890 1725 1928 1759
rect 1962 1725 2109 1759
rect 1709 1686 2109 1725
rect 1709 1652 1856 1686
rect 1890 1652 1928 1686
rect 1962 1652 2109 1686
rect 1709 1613 2109 1652
rect 1709 1579 1856 1613
rect 1890 1579 1928 1613
rect 1962 1579 2109 1613
rect 1709 1540 2109 1579
rect 1709 1506 1856 1540
rect 1890 1506 1928 1540
rect 1962 1506 2109 1540
rect 1709 1466 2109 1506
rect 1709 1432 1856 1466
rect 1890 1432 1928 1466
rect 1962 1432 2109 1466
rect 1709 1392 2109 1432
rect 1709 1358 1856 1392
rect 1890 1358 1928 1392
rect 1962 1358 2109 1392
rect 1709 1318 2109 1358
rect 1709 1284 1856 1318
rect 1890 1284 1928 1318
rect 1962 1284 2109 1318
rect 1709 1244 2109 1284
rect 1709 1210 1856 1244
rect 1890 1210 1928 1244
rect 1962 1210 2109 1244
rect 1709 1170 2109 1210
rect 1709 1136 1856 1170
rect 1890 1136 1928 1170
rect 1962 1136 2109 1170
rect 1709 1096 2109 1136
rect 1709 1062 1856 1096
rect 1890 1062 1928 1096
rect 1962 1062 2109 1096
rect 1709 1022 2109 1062
rect 1709 988 1856 1022
rect 1890 988 1928 1022
rect 1962 988 2109 1022
rect 1709 948 2109 988
rect 1709 914 1856 948
rect 1890 914 1928 948
rect 1962 914 2109 948
rect 1709 874 2109 914
rect 1709 840 1856 874
rect 1890 840 1928 874
rect 1962 840 2109 874
rect 1709 800 2109 840
rect 1709 766 1856 800
rect 1890 766 1928 800
rect 1962 766 2109 800
rect 1709 726 2109 766
rect 1709 692 1856 726
rect 1890 692 1928 726
rect 1962 692 2109 726
rect 1709 652 2109 692
rect 1709 618 1856 652
rect 1890 618 1928 652
rect 1962 618 2109 652
rect 1709 578 2109 618
rect 1709 544 1856 578
rect 1890 544 1928 578
rect 1962 544 2109 578
rect 1709 504 2109 544
rect 1709 470 1856 504
rect 1890 470 1928 504
rect 1962 470 2109 504
rect 1709 430 2109 470
rect 1709 396 1856 430
rect 1890 396 1928 430
rect 1962 396 2109 430
rect 1709 356 2109 396
rect 1709 322 1856 356
rect 1890 322 1928 356
rect 1962 322 2109 356
rect 1709 282 2109 322
rect 1709 248 1856 282
rect 1890 248 1928 282
rect 1962 248 2109 282
rect 1709 208 2109 248
rect 1709 174 1856 208
rect 1890 174 1928 208
rect 1962 174 2109 208
rect 1709 134 2109 174
rect 1709 100 1856 134
rect 1890 100 1928 134
rect 1962 100 2109 134
rect 1709 47 2109 100
tri 1709 42 1714 47 ne
rect 1714 42 2104 47
tri 2104 42 2109 47 nw
tri 2221 3053 2268 3100 se
rect 2268 3053 2374 3100
tri 2374 3053 2421 3100 sw
rect 2221 3000 2421 3053
rect 2221 2966 2268 3000
rect 2302 2966 2340 3000
rect 2374 2966 2421 3000
rect 2221 2927 2421 2966
rect 2221 2893 2268 2927
rect 2302 2893 2340 2927
rect 2374 2893 2421 2927
rect 2221 2854 2421 2893
rect 2221 2820 2268 2854
rect 2302 2820 2340 2854
rect 2374 2820 2421 2854
rect 2221 2781 2421 2820
rect 2221 2747 2268 2781
rect 2302 2747 2340 2781
rect 2374 2747 2421 2781
rect 2221 2708 2421 2747
rect 2221 2674 2268 2708
rect 2302 2674 2340 2708
rect 2374 2674 2421 2708
rect 2221 2635 2421 2674
rect 2221 2601 2268 2635
rect 2302 2601 2340 2635
rect 2374 2601 2421 2635
rect 2221 2562 2421 2601
rect 2221 2528 2268 2562
rect 2302 2528 2340 2562
rect 2374 2528 2421 2562
rect 2221 2489 2421 2528
rect 2221 2455 2268 2489
rect 2302 2455 2340 2489
rect 2374 2455 2421 2489
rect 2221 2416 2421 2455
rect 2221 2382 2268 2416
rect 2302 2382 2340 2416
rect 2374 2382 2421 2416
rect 2221 2343 2421 2382
rect 2221 2309 2268 2343
rect 2302 2309 2340 2343
rect 2374 2309 2421 2343
rect 2221 2270 2421 2309
rect 2221 2236 2268 2270
rect 2302 2236 2340 2270
rect 2374 2236 2421 2270
rect 2221 2197 2421 2236
rect 2221 2163 2268 2197
rect 2302 2163 2340 2197
rect 2374 2163 2421 2197
rect 2221 2124 2421 2163
rect 2221 2090 2268 2124
rect 2302 2090 2340 2124
rect 2374 2090 2421 2124
rect 2221 2051 2421 2090
rect 2221 2017 2268 2051
rect 2302 2017 2340 2051
rect 2374 2017 2421 2051
rect 2221 1978 2421 2017
rect 2221 1944 2268 1978
rect 2302 1944 2340 1978
rect 2374 1944 2421 1978
rect 2221 1905 2421 1944
rect 2221 1871 2268 1905
rect 2302 1871 2340 1905
rect 2374 1871 2421 1905
rect 2221 1832 2421 1871
rect 2221 1798 2268 1832
rect 2302 1798 2340 1832
rect 2374 1798 2421 1832
rect 2221 1759 2421 1798
rect 2221 1725 2268 1759
rect 2302 1725 2340 1759
rect 2374 1725 2421 1759
rect 2221 1686 2421 1725
rect 2221 1652 2268 1686
rect 2302 1652 2340 1686
rect 2374 1652 2421 1686
rect 2221 1613 2421 1652
rect 2221 1579 2268 1613
rect 2302 1579 2340 1613
rect 2374 1579 2421 1613
rect 2221 1540 2421 1579
rect 2221 1506 2268 1540
rect 2302 1506 2340 1540
rect 2374 1506 2421 1540
rect 2221 1466 2421 1506
rect 2221 1432 2268 1466
rect 2302 1432 2340 1466
rect 2374 1432 2421 1466
rect 2221 1392 2421 1432
rect 2221 1358 2268 1392
rect 2302 1358 2340 1392
rect 2374 1358 2421 1392
rect 2221 1318 2421 1358
rect 2221 1284 2268 1318
rect 2302 1284 2340 1318
rect 2374 1284 2421 1318
rect 2221 1244 2421 1284
rect 2221 1210 2268 1244
rect 2302 1210 2340 1244
rect 2374 1210 2421 1244
rect 2221 1170 2421 1210
rect 2221 1136 2268 1170
rect 2302 1136 2340 1170
rect 2374 1136 2421 1170
rect 2221 1096 2421 1136
rect 2221 1062 2268 1096
rect 2302 1062 2340 1096
rect 2374 1062 2421 1096
rect 2221 1022 2421 1062
rect 2221 988 2268 1022
rect 2302 988 2340 1022
rect 2374 988 2421 1022
rect 2221 948 2421 988
rect 2221 914 2268 948
rect 2302 914 2340 948
rect 2374 914 2421 948
rect 2221 874 2421 914
rect 2221 840 2268 874
rect 2302 840 2340 874
rect 2374 840 2421 874
rect 2221 800 2421 840
rect 2221 766 2268 800
rect 2302 766 2340 800
rect 2374 766 2421 800
rect 2221 726 2421 766
rect 2221 692 2268 726
rect 2302 692 2340 726
rect 2374 692 2421 726
rect 2221 652 2421 692
rect 2221 618 2268 652
rect 2302 618 2340 652
rect 2374 618 2421 652
rect 2221 578 2421 618
rect 2221 544 2268 578
rect 2302 544 2340 578
rect 2374 544 2421 578
rect 2221 504 2421 544
rect 2221 470 2268 504
rect 2302 470 2340 504
rect 2374 470 2421 504
rect 2221 430 2421 470
rect 2221 396 2268 430
rect 2302 396 2340 430
rect 2374 396 2421 430
rect 2221 356 2421 396
rect 2221 322 2268 356
rect 2302 322 2340 356
rect 2374 322 2421 356
rect 2221 282 2421 322
rect 2221 248 2268 282
rect 2302 248 2340 282
rect 2374 248 2421 282
rect 2221 208 2421 248
rect 2221 174 2268 208
rect 2302 174 2340 208
rect 2374 174 2421 208
rect 2221 134 2421 174
rect 2221 100 2268 134
rect 2302 100 2340 134
rect 2374 100 2421 134
rect 2221 47 2421 100
tri 2221 42 2226 47 ne
rect 2226 42 2416 47
tri 2416 42 2421 47 nw
tri 2533 3053 2580 3100 se
rect 2580 3053 2886 3100
tri 2886 3053 2933 3100 sw
rect 2533 3000 2933 3053
rect 2533 2966 2680 3000
rect 2714 2966 2752 3000
rect 2786 2966 2933 3000
rect 2533 2927 2933 2966
rect 2533 2893 2680 2927
rect 2714 2893 2752 2927
rect 2786 2893 2933 2927
rect 2533 2854 2933 2893
rect 2533 2820 2680 2854
rect 2714 2820 2752 2854
rect 2786 2820 2933 2854
rect 2533 2781 2933 2820
rect 2533 2747 2680 2781
rect 2714 2747 2752 2781
rect 2786 2747 2933 2781
rect 2533 2708 2933 2747
rect 2533 2674 2680 2708
rect 2714 2674 2752 2708
rect 2786 2674 2933 2708
rect 2533 2635 2933 2674
rect 2533 2601 2680 2635
rect 2714 2601 2752 2635
rect 2786 2601 2933 2635
rect 2533 2562 2933 2601
rect 2533 2528 2680 2562
rect 2714 2528 2752 2562
rect 2786 2528 2933 2562
rect 2533 2489 2933 2528
rect 2533 2455 2680 2489
rect 2714 2455 2752 2489
rect 2786 2455 2933 2489
rect 2533 2416 2933 2455
rect 2533 2382 2680 2416
rect 2714 2382 2752 2416
rect 2786 2382 2933 2416
rect 2533 2343 2933 2382
rect 2533 2309 2680 2343
rect 2714 2309 2752 2343
rect 2786 2309 2933 2343
rect 2533 2270 2933 2309
rect 2533 2236 2680 2270
rect 2714 2236 2752 2270
rect 2786 2236 2933 2270
rect 2533 2197 2933 2236
rect 2533 2163 2680 2197
rect 2714 2163 2752 2197
rect 2786 2163 2933 2197
rect 2533 2124 2933 2163
rect 2533 2090 2680 2124
rect 2714 2090 2752 2124
rect 2786 2090 2933 2124
rect 2533 2051 2933 2090
rect 2533 2017 2680 2051
rect 2714 2017 2752 2051
rect 2786 2017 2933 2051
rect 2533 1978 2933 2017
rect 2533 1944 2680 1978
rect 2714 1944 2752 1978
rect 2786 1944 2933 1978
rect 2533 1905 2933 1944
rect 2533 1871 2680 1905
rect 2714 1871 2752 1905
rect 2786 1871 2933 1905
rect 2533 1832 2933 1871
rect 2533 1798 2680 1832
rect 2714 1798 2752 1832
rect 2786 1798 2933 1832
rect 2533 1759 2933 1798
rect 2533 1725 2680 1759
rect 2714 1725 2752 1759
rect 2786 1725 2933 1759
rect 2533 1686 2933 1725
rect 2533 1652 2680 1686
rect 2714 1652 2752 1686
rect 2786 1652 2933 1686
rect 2533 1613 2933 1652
rect 2533 1579 2680 1613
rect 2714 1579 2752 1613
rect 2786 1579 2933 1613
rect 2533 1540 2933 1579
rect 2533 1506 2680 1540
rect 2714 1506 2752 1540
rect 2786 1506 2933 1540
rect 2533 1466 2933 1506
rect 2533 1432 2680 1466
rect 2714 1432 2752 1466
rect 2786 1432 2933 1466
rect 2533 1392 2933 1432
rect 2533 1358 2680 1392
rect 2714 1358 2752 1392
rect 2786 1358 2933 1392
rect 2533 1318 2933 1358
rect 2533 1284 2680 1318
rect 2714 1284 2752 1318
rect 2786 1284 2933 1318
rect 2533 1244 2933 1284
rect 2533 1210 2680 1244
rect 2714 1210 2752 1244
rect 2786 1210 2933 1244
rect 2533 1170 2933 1210
rect 2533 1136 2680 1170
rect 2714 1136 2752 1170
rect 2786 1136 2933 1170
rect 2533 1096 2933 1136
rect 2533 1062 2680 1096
rect 2714 1062 2752 1096
rect 2786 1062 2933 1096
rect 2533 1022 2933 1062
rect 2533 988 2680 1022
rect 2714 988 2752 1022
rect 2786 988 2933 1022
rect 2533 948 2933 988
rect 2533 914 2680 948
rect 2714 914 2752 948
rect 2786 914 2933 948
rect 2533 874 2933 914
rect 2533 840 2680 874
rect 2714 840 2752 874
rect 2786 840 2933 874
rect 2533 800 2933 840
rect 2533 766 2680 800
rect 2714 766 2752 800
rect 2786 766 2933 800
rect 2533 726 2933 766
rect 2533 692 2680 726
rect 2714 692 2752 726
rect 2786 692 2933 726
rect 2533 652 2933 692
rect 2533 618 2680 652
rect 2714 618 2752 652
rect 2786 618 2933 652
rect 2533 578 2933 618
rect 2533 544 2680 578
rect 2714 544 2752 578
rect 2786 544 2933 578
rect 2533 504 2933 544
rect 2533 470 2680 504
rect 2714 470 2752 504
rect 2786 470 2933 504
rect 2533 430 2933 470
rect 2533 396 2680 430
rect 2714 396 2752 430
rect 2786 396 2933 430
rect 2533 356 2933 396
rect 2533 322 2680 356
rect 2714 322 2752 356
rect 2786 322 2933 356
rect 2533 282 2933 322
rect 2533 248 2680 282
rect 2714 248 2752 282
rect 2786 248 2933 282
rect 2533 208 2933 248
rect 2533 174 2680 208
rect 2714 174 2752 208
rect 2786 174 2933 208
rect 2533 134 2933 174
rect 2533 100 2680 134
rect 2714 100 2752 134
rect 2786 100 2933 134
rect 2533 47 2933 100
tri 2533 42 2538 47 ne
rect 2538 42 2928 47
tri 2928 42 2933 47 nw
tri 3045 3053 3092 3100 se
rect 3092 3053 3198 3100
tri 3198 3053 3245 3100 sw
rect 3045 3000 3245 3053
rect 3045 2966 3092 3000
rect 3126 2966 3164 3000
rect 3198 2966 3245 3000
rect 3045 2927 3245 2966
rect 3045 2893 3092 2927
rect 3126 2893 3164 2927
rect 3198 2893 3245 2927
rect 3045 2854 3245 2893
rect 3045 2820 3092 2854
rect 3126 2820 3164 2854
rect 3198 2820 3245 2854
rect 3045 2781 3245 2820
rect 3045 2747 3092 2781
rect 3126 2747 3164 2781
rect 3198 2747 3245 2781
rect 3045 2708 3245 2747
rect 3045 2674 3092 2708
rect 3126 2674 3164 2708
rect 3198 2674 3245 2708
rect 3045 2635 3245 2674
rect 3045 2601 3092 2635
rect 3126 2601 3164 2635
rect 3198 2601 3245 2635
rect 3045 2562 3245 2601
rect 3045 2528 3092 2562
rect 3126 2528 3164 2562
rect 3198 2528 3245 2562
rect 3045 2489 3245 2528
rect 3045 2455 3092 2489
rect 3126 2455 3164 2489
rect 3198 2455 3245 2489
rect 3045 2416 3245 2455
rect 3045 2382 3092 2416
rect 3126 2382 3164 2416
rect 3198 2382 3245 2416
rect 3045 2343 3245 2382
rect 3045 2309 3092 2343
rect 3126 2309 3164 2343
rect 3198 2309 3245 2343
rect 3045 2270 3245 2309
rect 3045 2236 3092 2270
rect 3126 2236 3164 2270
rect 3198 2236 3245 2270
rect 3045 2197 3245 2236
rect 3045 2163 3092 2197
rect 3126 2163 3164 2197
rect 3198 2163 3245 2197
rect 3045 2124 3245 2163
rect 3045 2090 3092 2124
rect 3126 2090 3164 2124
rect 3198 2090 3245 2124
rect 3045 2051 3245 2090
rect 3045 2017 3092 2051
rect 3126 2017 3164 2051
rect 3198 2017 3245 2051
rect 3045 1978 3245 2017
rect 3045 1944 3092 1978
rect 3126 1944 3164 1978
rect 3198 1944 3245 1978
rect 3045 1905 3245 1944
rect 3045 1871 3092 1905
rect 3126 1871 3164 1905
rect 3198 1871 3245 1905
rect 3045 1832 3245 1871
rect 3045 1798 3092 1832
rect 3126 1798 3164 1832
rect 3198 1798 3245 1832
rect 3045 1759 3245 1798
rect 3045 1725 3092 1759
rect 3126 1725 3164 1759
rect 3198 1725 3245 1759
rect 3045 1686 3245 1725
rect 3045 1652 3092 1686
rect 3126 1652 3164 1686
rect 3198 1652 3245 1686
rect 3045 1613 3245 1652
rect 3045 1579 3092 1613
rect 3126 1579 3164 1613
rect 3198 1579 3245 1613
rect 3045 1540 3245 1579
rect 3045 1506 3092 1540
rect 3126 1506 3164 1540
rect 3198 1506 3245 1540
rect 3045 1466 3245 1506
rect 3045 1432 3092 1466
rect 3126 1432 3164 1466
rect 3198 1432 3245 1466
rect 3045 1392 3245 1432
rect 3045 1358 3092 1392
rect 3126 1358 3164 1392
rect 3198 1358 3245 1392
rect 3045 1318 3245 1358
rect 3045 1284 3092 1318
rect 3126 1284 3164 1318
rect 3198 1284 3245 1318
rect 3045 1244 3245 1284
rect 3045 1210 3092 1244
rect 3126 1210 3164 1244
rect 3198 1210 3245 1244
rect 3045 1170 3245 1210
rect 3045 1136 3092 1170
rect 3126 1136 3164 1170
rect 3198 1136 3245 1170
rect 3045 1096 3245 1136
rect 3045 1062 3092 1096
rect 3126 1062 3164 1096
rect 3198 1062 3245 1096
rect 3045 1022 3245 1062
rect 3045 988 3092 1022
rect 3126 988 3164 1022
rect 3198 988 3245 1022
rect 3045 948 3245 988
rect 3045 914 3092 948
rect 3126 914 3164 948
rect 3198 914 3245 948
rect 3045 874 3245 914
rect 3045 840 3092 874
rect 3126 840 3164 874
rect 3198 840 3245 874
rect 3045 800 3245 840
rect 3045 766 3092 800
rect 3126 766 3164 800
rect 3198 766 3245 800
rect 3045 726 3245 766
rect 3045 692 3092 726
rect 3126 692 3164 726
rect 3198 692 3245 726
rect 3045 652 3245 692
rect 3045 618 3092 652
rect 3126 618 3164 652
rect 3198 618 3245 652
rect 3045 578 3245 618
rect 3045 544 3092 578
rect 3126 544 3164 578
rect 3198 544 3245 578
rect 3045 504 3245 544
rect 3045 470 3092 504
rect 3126 470 3164 504
rect 3198 470 3245 504
rect 3045 430 3245 470
rect 3045 396 3092 430
rect 3126 396 3164 430
rect 3198 396 3245 430
rect 3045 356 3245 396
rect 3045 322 3092 356
rect 3126 322 3164 356
rect 3198 322 3245 356
rect 3045 282 3245 322
rect 3045 248 3092 282
rect 3126 248 3164 282
rect 3198 248 3245 282
rect 3045 208 3245 248
rect 3045 174 3092 208
rect 3126 174 3164 208
rect 3198 174 3245 208
rect 3045 134 3245 174
rect 3045 100 3092 134
rect 3126 100 3164 134
rect 3198 100 3245 134
rect 3045 47 3245 100
tri 3045 42 3050 47 ne
rect 3050 42 3240 47
tri 3240 42 3245 47 nw
tri 3357 3053 3404 3100 se
rect 3404 3053 3710 3100
tri 3710 3053 3757 3100 sw
rect 3357 3000 3757 3053
rect 3357 2966 3504 3000
rect 3538 2966 3576 3000
rect 3610 2966 3757 3000
rect 3357 2927 3757 2966
rect 3357 2893 3504 2927
rect 3538 2893 3576 2927
rect 3610 2893 3757 2927
rect 3357 2854 3757 2893
rect 3357 2820 3504 2854
rect 3538 2820 3576 2854
rect 3610 2820 3757 2854
rect 3357 2781 3757 2820
rect 3357 2747 3504 2781
rect 3538 2747 3576 2781
rect 3610 2747 3757 2781
rect 3357 2708 3757 2747
rect 3357 2674 3504 2708
rect 3538 2674 3576 2708
rect 3610 2674 3757 2708
rect 3357 2635 3757 2674
rect 3357 2601 3504 2635
rect 3538 2601 3576 2635
rect 3610 2601 3757 2635
rect 3357 2562 3757 2601
rect 3357 2528 3504 2562
rect 3538 2528 3576 2562
rect 3610 2528 3757 2562
rect 3357 2489 3757 2528
rect 3357 2455 3504 2489
rect 3538 2455 3576 2489
rect 3610 2455 3757 2489
rect 3357 2416 3757 2455
rect 3357 2382 3504 2416
rect 3538 2382 3576 2416
rect 3610 2382 3757 2416
rect 3357 2343 3757 2382
rect 3357 2309 3504 2343
rect 3538 2309 3576 2343
rect 3610 2309 3757 2343
rect 3357 2270 3757 2309
rect 3357 2236 3504 2270
rect 3538 2236 3576 2270
rect 3610 2236 3757 2270
rect 3357 2197 3757 2236
rect 3357 2163 3504 2197
rect 3538 2163 3576 2197
rect 3610 2163 3757 2197
rect 3357 2124 3757 2163
rect 3357 2090 3504 2124
rect 3538 2090 3576 2124
rect 3610 2090 3757 2124
rect 3357 2051 3757 2090
rect 3357 2017 3504 2051
rect 3538 2017 3576 2051
rect 3610 2017 3757 2051
rect 3357 1978 3757 2017
rect 3357 1944 3504 1978
rect 3538 1944 3576 1978
rect 3610 1944 3757 1978
rect 3357 1905 3757 1944
rect 3357 1871 3504 1905
rect 3538 1871 3576 1905
rect 3610 1871 3757 1905
rect 3357 1832 3757 1871
rect 3357 1798 3504 1832
rect 3538 1798 3576 1832
rect 3610 1798 3757 1832
rect 3357 1759 3757 1798
rect 3357 1725 3504 1759
rect 3538 1725 3576 1759
rect 3610 1725 3757 1759
rect 3357 1686 3757 1725
rect 3357 1652 3504 1686
rect 3538 1652 3576 1686
rect 3610 1652 3757 1686
rect 3357 1613 3757 1652
rect 3357 1579 3504 1613
rect 3538 1579 3576 1613
rect 3610 1579 3757 1613
rect 3357 1540 3757 1579
rect 3357 1506 3504 1540
rect 3538 1506 3576 1540
rect 3610 1506 3757 1540
rect 3357 1466 3757 1506
rect 3357 1432 3504 1466
rect 3538 1432 3576 1466
rect 3610 1432 3757 1466
rect 3357 1392 3757 1432
rect 3357 1358 3504 1392
rect 3538 1358 3576 1392
rect 3610 1358 3757 1392
rect 3357 1318 3757 1358
rect 3357 1284 3504 1318
rect 3538 1284 3576 1318
rect 3610 1284 3757 1318
rect 3357 1244 3757 1284
rect 3357 1210 3504 1244
rect 3538 1210 3576 1244
rect 3610 1210 3757 1244
rect 3357 1170 3757 1210
rect 3357 1136 3504 1170
rect 3538 1136 3576 1170
rect 3610 1136 3757 1170
rect 3357 1096 3757 1136
rect 3357 1062 3504 1096
rect 3538 1062 3576 1096
rect 3610 1062 3757 1096
rect 3357 1022 3757 1062
rect 3357 988 3504 1022
rect 3538 988 3576 1022
rect 3610 988 3757 1022
rect 3357 948 3757 988
rect 3357 914 3504 948
rect 3538 914 3576 948
rect 3610 914 3757 948
rect 3357 874 3757 914
rect 3357 840 3504 874
rect 3538 840 3576 874
rect 3610 840 3757 874
rect 3357 800 3757 840
rect 3357 766 3504 800
rect 3538 766 3576 800
rect 3610 766 3757 800
rect 3357 726 3757 766
rect 3357 692 3504 726
rect 3538 692 3576 726
rect 3610 692 3757 726
rect 3357 652 3757 692
rect 3357 618 3504 652
rect 3538 618 3576 652
rect 3610 618 3757 652
rect 3357 578 3757 618
rect 3357 544 3504 578
rect 3538 544 3576 578
rect 3610 544 3757 578
rect 3357 504 3757 544
rect 3357 470 3504 504
rect 3538 470 3576 504
rect 3610 470 3757 504
rect 3357 430 3757 470
rect 3357 396 3504 430
rect 3538 396 3576 430
rect 3610 396 3757 430
rect 3357 356 3757 396
rect 3357 322 3504 356
rect 3538 322 3576 356
rect 3610 322 3757 356
rect 3357 282 3757 322
rect 3357 248 3504 282
rect 3538 248 3576 282
rect 3610 248 3757 282
rect 3357 208 3757 248
rect 3357 174 3504 208
rect 3538 174 3576 208
rect 3610 174 3757 208
rect 3357 134 3757 174
rect 3357 100 3504 134
rect 3538 100 3576 134
rect 3610 100 3757 134
rect 3357 47 3757 100
tri 3357 42 3362 47 ne
rect 3362 42 3752 47
tri 3752 42 3757 47 nw
tri 3869 3053 3916 3100 se
rect 3916 3053 4022 3100
tri 4022 3053 4069 3100 sw
rect 3869 3000 4069 3053
rect 3869 2966 3916 3000
rect 3950 2966 3988 3000
rect 4022 2966 4069 3000
rect 3869 2927 4069 2966
rect 3869 2893 3916 2927
rect 3950 2893 3988 2927
rect 4022 2893 4069 2927
rect 3869 2854 4069 2893
rect 3869 2820 3916 2854
rect 3950 2820 3988 2854
rect 4022 2820 4069 2854
rect 3869 2781 4069 2820
rect 3869 2747 3916 2781
rect 3950 2747 3988 2781
rect 4022 2747 4069 2781
rect 3869 2708 4069 2747
rect 3869 2674 3916 2708
rect 3950 2674 3988 2708
rect 4022 2674 4069 2708
rect 3869 2635 4069 2674
rect 3869 2601 3916 2635
rect 3950 2601 3988 2635
rect 4022 2601 4069 2635
rect 3869 2562 4069 2601
rect 3869 2528 3916 2562
rect 3950 2528 3988 2562
rect 4022 2528 4069 2562
rect 3869 2489 4069 2528
rect 3869 2455 3916 2489
rect 3950 2455 3988 2489
rect 4022 2455 4069 2489
rect 3869 2416 4069 2455
rect 3869 2382 3916 2416
rect 3950 2382 3988 2416
rect 4022 2382 4069 2416
rect 3869 2343 4069 2382
rect 3869 2309 3916 2343
rect 3950 2309 3988 2343
rect 4022 2309 4069 2343
rect 3869 2270 4069 2309
rect 3869 2236 3916 2270
rect 3950 2236 3988 2270
rect 4022 2236 4069 2270
rect 3869 2197 4069 2236
rect 3869 2163 3916 2197
rect 3950 2163 3988 2197
rect 4022 2163 4069 2197
rect 3869 2124 4069 2163
rect 3869 2090 3916 2124
rect 3950 2090 3988 2124
rect 4022 2090 4069 2124
rect 3869 2051 4069 2090
rect 3869 2017 3916 2051
rect 3950 2017 3988 2051
rect 4022 2017 4069 2051
rect 3869 1978 4069 2017
rect 3869 1944 3916 1978
rect 3950 1944 3988 1978
rect 4022 1944 4069 1978
rect 3869 1905 4069 1944
rect 3869 1871 3916 1905
rect 3950 1871 3988 1905
rect 4022 1871 4069 1905
rect 3869 1832 4069 1871
rect 3869 1798 3916 1832
rect 3950 1798 3988 1832
rect 4022 1798 4069 1832
rect 3869 1759 4069 1798
rect 3869 1725 3916 1759
rect 3950 1725 3988 1759
rect 4022 1725 4069 1759
rect 3869 1686 4069 1725
rect 3869 1652 3916 1686
rect 3950 1652 3988 1686
rect 4022 1652 4069 1686
rect 3869 1613 4069 1652
rect 3869 1579 3916 1613
rect 3950 1579 3988 1613
rect 4022 1579 4069 1613
rect 3869 1540 4069 1579
rect 3869 1506 3916 1540
rect 3950 1506 3988 1540
rect 4022 1506 4069 1540
rect 3869 1466 4069 1506
rect 3869 1432 3916 1466
rect 3950 1432 3988 1466
rect 4022 1432 4069 1466
rect 3869 1392 4069 1432
rect 3869 1358 3916 1392
rect 3950 1358 3988 1392
rect 4022 1358 4069 1392
rect 3869 1318 4069 1358
rect 3869 1284 3916 1318
rect 3950 1284 3988 1318
rect 4022 1284 4069 1318
rect 3869 1244 4069 1284
rect 3869 1210 3916 1244
rect 3950 1210 3988 1244
rect 4022 1210 4069 1244
rect 3869 1170 4069 1210
rect 3869 1136 3916 1170
rect 3950 1136 3988 1170
rect 4022 1136 4069 1170
rect 3869 1096 4069 1136
rect 3869 1062 3916 1096
rect 3950 1062 3988 1096
rect 4022 1062 4069 1096
rect 3869 1022 4069 1062
rect 3869 988 3916 1022
rect 3950 988 3988 1022
rect 4022 988 4069 1022
rect 3869 948 4069 988
rect 3869 914 3916 948
rect 3950 914 3988 948
rect 4022 914 4069 948
rect 3869 874 4069 914
rect 3869 840 3916 874
rect 3950 840 3988 874
rect 4022 840 4069 874
rect 3869 800 4069 840
rect 3869 766 3916 800
rect 3950 766 3988 800
rect 4022 766 4069 800
rect 3869 726 4069 766
rect 3869 692 3916 726
rect 3950 692 3988 726
rect 4022 692 4069 726
rect 3869 652 4069 692
rect 3869 618 3916 652
rect 3950 618 3988 652
rect 4022 618 4069 652
rect 3869 578 4069 618
rect 3869 544 3916 578
rect 3950 544 3988 578
rect 4022 544 4069 578
rect 3869 504 4069 544
rect 3869 470 3916 504
rect 3950 470 3988 504
rect 4022 470 4069 504
rect 3869 430 4069 470
rect 3869 396 3916 430
rect 3950 396 3988 430
rect 4022 396 4069 430
rect 3869 356 4069 396
rect 3869 322 3916 356
rect 3950 322 3988 356
rect 4022 322 4069 356
rect 3869 282 4069 322
rect 3869 248 3916 282
rect 3950 248 3988 282
rect 4022 248 4069 282
rect 3869 208 4069 248
rect 3869 174 3916 208
rect 3950 174 3988 208
rect 4022 174 4069 208
rect 3869 134 4069 174
rect 3869 100 3916 134
rect 3950 100 3988 134
rect 4022 100 4069 134
rect 3869 47 4069 100
tri 3869 42 3874 47 ne
rect 3874 42 4064 47
tri 4064 42 4069 47 nw
tri 4181 3053 4228 3100 se
rect 4228 3053 4534 3100
tri 4534 3053 4581 3100 sw
rect 4181 3000 4581 3053
rect 4181 2966 4328 3000
rect 4362 2966 4400 3000
rect 4434 2966 4581 3000
rect 4181 2927 4581 2966
rect 4181 2893 4328 2927
rect 4362 2893 4400 2927
rect 4434 2893 4581 2927
rect 4181 2854 4581 2893
rect 4181 2820 4328 2854
rect 4362 2820 4400 2854
rect 4434 2820 4581 2854
rect 4181 2781 4581 2820
rect 4181 2747 4328 2781
rect 4362 2747 4400 2781
rect 4434 2747 4581 2781
rect 4181 2708 4581 2747
rect 4181 2674 4328 2708
rect 4362 2674 4400 2708
rect 4434 2674 4581 2708
rect 4181 2635 4581 2674
rect 4181 2601 4328 2635
rect 4362 2601 4400 2635
rect 4434 2601 4581 2635
rect 4181 2562 4581 2601
rect 4181 2528 4328 2562
rect 4362 2528 4400 2562
rect 4434 2528 4581 2562
rect 4181 2489 4581 2528
rect 4181 2455 4328 2489
rect 4362 2455 4400 2489
rect 4434 2455 4581 2489
rect 4181 2416 4581 2455
rect 4181 2382 4328 2416
rect 4362 2382 4400 2416
rect 4434 2382 4581 2416
rect 4181 2343 4581 2382
rect 4181 2309 4328 2343
rect 4362 2309 4400 2343
rect 4434 2309 4581 2343
rect 4181 2270 4581 2309
rect 4181 2236 4328 2270
rect 4362 2236 4400 2270
rect 4434 2236 4581 2270
rect 4181 2197 4581 2236
rect 4181 2163 4328 2197
rect 4362 2163 4400 2197
rect 4434 2163 4581 2197
rect 4181 2124 4581 2163
rect 4181 2090 4328 2124
rect 4362 2090 4400 2124
rect 4434 2090 4581 2124
rect 4181 2051 4581 2090
rect 4181 2017 4328 2051
rect 4362 2017 4400 2051
rect 4434 2017 4581 2051
rect 4181 1978 4581 2017
rect 4181 1944 4328 1978
rect 4362 1944 4400 1978
rect 4434 1944 4581 1978
rect 4181 1905 4581 1944
rect 4181 1871 4328 1905
rect 4362 1871 4400 1905
rect 4434 1871 4581 1905
rect 4181 1832 4581 1871
rect 4181 1798 4328 1832
rect 4362 1798 4400 1832
rect 4434 1798 4581 1832
rect 4181 1759 4581 1798
rect 4181 1725 4328 1759
rect 4362 1725 4400 1759
rect 4434 1725 4581 1759
rect 4181 1686 4581 1725
rect 4181 1652 4328 1686
rect 4362 1652 4400 1686
rect 4434 1652 4581 1686
rect 4181 1613 4581 1652
rect 4181 1579 4328 1613
rect 4362 1579 4400 1613
rect 4434 1579 4581 1613
rect 4181 1540 4581 1579
rect 4181 1506 4328 1540
rect 4362 1506 4400 1540
rect 4434 1506 4581 1540
rect 4181 1466 4581 1506
rect 4181 1432 4328 1466
rect 4362 1432 4400 1466
rect 4434 1432 4581 1466
rect 4181 1392 4581 1432
rect 4181 1358 4328 1392
rect 4362 1358 4400 1392
rect 4434 1358 4581 1392
rect 4181 1318 4581 1358
rect 4181 1284 4328 1318
rect 4362 1284 4400 1318
rect 4434 1284 4581 1318
rect 4181 1244 4581 1284
rect 4181 1210 4328 1244
rect 4362 1210 4400 1244
rect 4434 1210 4581 1244
rect 4181 1170 4581 1210
rect 4181 1136 4328 1170
rect 4362 1136 4400 1170
rect 4434 1136 4581 1170
rect 4181 1096 4581 1136
rect 4181 1062 4328 1096
rect 4362 1062 4400 1096
rect 4434 1062 4581 1096
rect 4181 1022 4581 1062
rect 4181 988 4328 1022
rect 4362 988 4400 1022
rect 4434 988 4581 1022
rect 4181 948 4581 988
rect 4181 914 4328 948
rect 4362 914 4400 948
rect 4434 914 4581 948
rect 4181 874 4581 914
rect 4181 840 4328 874
rect 4362 840 4400 874
rect 4434 840 4581 874
rect 4181 800 4581 840
rect 4181 766 4328 800
rect 4362 766 4400 800
rect 4434 766 4581 800
rect 4181 726 4581 766
rect 4181 692 4328 726
rect 4362 692 4400 726
rect 4434 692 4581 726
rect 4181 652 4581 692
rect 4181 618 4328 652
rect 4362 618 4400 652
rect 4434 618 4581 652
rect 4181 578 4581 618
rect 4181 544 4328 578
rect 4362 544 4400 578
rect 4434 544 4581 578
rect 4181 504 4581 544
rect 4181 470 4328 504
rect 4362 470 4400 504
rect 4434 470 4581 504
rect 4181 430 4581 470
rect 4181 396 4328 430
rect 4362 396 4400 430
rect 4434 396 4581 430
rect 4181 356 4581 396
rect 4181 322 4328 356
rect 4362 322 4400 356
rect 4434 322 4581 356
rect 4181 282 4581 322
rect 4181 248 4328 282
rect 4362 248 4400 282
rect 4434 248 4581 282
rect 4181 208 4581 248
rect 4181 174 4328 208
rect 4362 174 4400 208
rect 4434 174 4581 208
rect 4181 134 4581 174
rect 4181 100 4328 134
rect 4362 100 4400 134
rect 4434 100 4581 134
rect 4181 47 4581 100
tri 4181 42 4186 47 ne
rect 4186 42 4576 47
tri 4576 42 4581 47 nw
tri 4693 3053 4740 3100 se
rect 4740 3053 4846 3100
tri 4846 3053 4893 3100 sw
rect 4693 3000 4893 3053
rect 4693 2966 4740 3000
rect 4774 2966 4812 3000
rect 4846 2966 4893 3000
rect 4693 2927 4893 2966
rect 4693 2893 4740 2927
rect 4774 2893 4812 2927
rect 4846 2893 4893 2927
rect 4693 2854 4893 2893
rect 4693 2820 4740 2854
rect 4774 2820 4812 2854
rect 4846 2820 4893 2854
rect 4693 2781 4893 2820
rect 4693 2747 4740 2781
rect 4774 2747 4812 2781
rect 4846 2747 4893 2781
rect 4693 2708 4893 2747
rect 4693 2674 4740 2708
rect 4774 2674 4812 2708
rect 4846 2674 4893 2708
rect 4693 2635 4893 2674
rect 4693 2601 4740 2635
rect 4774 2601 4812 2635
rect 4846 2601 4893 2635
rect 4693 2562 4893 2601
rect 4693 2528 4740 2562
rect 4774 2528 4812 2562
rect 4846 2528 4893 2562
rect 4693 2489 4893 2528
rect 4693 2455 4740 2489
rect 4774 2455 4812 2489
rect 4846 2455 4893 2489
rect 4693 2416 4893 2455
rect 4693 2382 4740 2416
rect 4774 2382 4812 2416
rect 4846 2382 4893 2416
rect 4693 2343 4893 2382
rect 4693 2309 4740 2343
rect 4774 2309 4812 2343
rect 4846 2309 4893 2343
rect 4693 2270 4893 2309
rect 4693 2236 4740 2270
rect 4774 2236 4812 2270
rect 4846 2236 4893 2270
rect 4693 2197 4893 2236
rect 4693 2163 4740 2197
rect 4774 2163 4812 2197
rect 4846 2163 4893 2197
rect 4693 2124 4893 2163
rect 4693 2090 4740 2124
rect 4774 2090 4812 2124
rect 4846 2090 4893 2124
rect 4693 2051 4893 2090
rect 4693 2017 4740 2051
rect 4774 2017 4812 2051
rect 4846 2017 4893 2051
rect 4693 1978 4893 2017
rect 4693 1944 4740 1978
rect 4774 1944 4812 1978
rect 4846 1944 4893 1978
rect 4693 1905 4893 1944
rect 4693 1871 4740 1905
rect 4774 1871 4812 1905
rect 4846 1871 4893 1905
rect 4693 1832 4893 1871
rect 4693 1798 4740 1832
rect 4774 1798 4812 1832
rect 4846 1798 4893 1832
rect 4693 1759 4893 1798
rect 4693 1725 4740 1759
rect 4774 1725 4812 1759
rect 4846 1725 4893 1759
rect 4693 1686 4893 1725
rect 4693 1652 4740 1686
rect 4774 1652 4812 1686
rect 4846 1652 4893 1686
rect 4693 1613 4893 1652
rect 4693 1579 4740 1613
rect 4774 1579 4812 1613
rect 4846 1579 4893 1613
rect 4693 1540 4893 1579
rect 4693 1506 4740 1540
rect 4774 1506 4812 1540
rect 4846 1506 4893 1540
rect 4693 1466 4893 1506
rect 4693 1432 4740 1466
rect 4774 1432 4812 1466
rect 4846 1432 4893 1466
rect 4693 1392 4893 1432
rect 4693 1358 4740 1392
rect 4774 1358 4812 1392
rect 4846 1358 4893 1392
rect 4693 1318 4893 1358
rect 4693 1284 4740 1318
rect 4774 1284 4812 1318
rect 4846 1284 4893 1318
rect 4693 1244 4893 1284
rect 4693 1210 4740 1244
rect 4774 1210 4812 1244
rect 4846 1210 4893 1244
rect 4693 1170 4893 1210
rect 4693 1136 4740 1170
rect 4774 1136 4812 1170
rect 4846 1136 4893 1170
rect 4693 1096 4893 1136
rect 4693 1062 4740 1096
rect 4774 1062 4812 1096
rect 4846 1062 4893 1096
rect 4693 1022 4893 1062
rect 4693 988 4740 1022
rect 4774 988 4812 1022
rect 4846 988 4893 1022
rect 4693 948 4893 988
rect 4693 914 4740 948
rect 4774 914 4812 948
rect 4846 914 4893 948
rect 4693 874 4893 914
rect 4693 840 4740 874
rect 4774 840 4812 874
rect 4846 840 4893 874
rect 4693 800 4893 840
rect 4693 766 4740 800
rect 4774 766 4812 800
rect 4846 766 4893 800
rect 4693 726 4893 766
rect 4693 692 4740 726
rect 4774 692 4812 726
rect 4846 692 4893 726
rect 4693 652 4893 692
rect 4693 618 4740 652
rect 4774 618 4812 652
rect 4846 618 4893 652
rect 4693 578 4893 618
rect 4693 544 4740 578
rect 4774 544 4812 578
rect 4846 544 4893 578
rect 4693 504 4893 544
rect 4693 470 4740 504
rect 4774 470 4812 504
rect 4846 470 4893 504
rect 4693 430 4893 470
rect 4693 396 4740 430
rect 4774 396 4812 430
rect 4846 396 4893 430
rect 4693 356 4893 396
rect 4693 322 4740 356
rect 4774 322 4812 356
rect 4846 322 4893 356
rect 4693 282 4893 322
rect 4693 248 4740 282
rect 4774 248 4812 282
rect 4846 248 4893 282
rect 4693 208 4893 248
rect 4693 174 4740 208
rect 4774 174 4812 208
rect 4846 174 4893 208
rect 4693 134 4893 174
rect 4693 100 4740 134
rect 4774 100 4812 134
rect 4846 100 4893 134
rect 4693 47 4893 100
tri 4693 42 4698 47 ne
rect 4698 42 4888 47
tri 4888 42 4893 47 nw
tri 5005 3053 5052 3100 se
rect 5052 3053 5358 3100
tri 5358 3053 5405 3100 sw
rect 5005 3000 5405 3053
rect 5005 2966 5152 3000
rect 5186 2966 5224 3000
rect 5258 2966 5405 3000
rect 5005 2927 5405 2966
rect 5005 2893 5152 2927
rect 5186 2893 5224 2927
rect 5258 2893 5405 2927
rect 5005 2854 5405 2893
rect 5005 2820 5152 2854
rect 5186 2820 5224 2854
rect 5258 2820 5405 2854
rect 5005 2781 5405 2820
rect 5005 2747 5152 2781
rect 5186 2747 5224 2781
rect 5258 2747 5405 2781
rect 5005 2708 5405 2747
rect 5005 2674 5152 2708
rect 5186 2674 5224 2708
rect 5258 2674 5405 2708
rect 5005 2635 5405 2674
rect 5005 2601 5152 2635
rect 5186 2601 5224 2635
rect 5258 2601 5405 2635
rect 5005 2562 5405 2601
rect 5005 2528 5152 2562
rect 5186 2528 5224 2562
rect 5258 2528 5405 2562
rect 5005 2489 5405 2528
rect 5005 2455 5152 2489
rect 5186 2455 5224 2489
rect 5258 2455 5405 2489
rect 5005 2416 5405 2455
rect 5005 2382 5152 2416
rect 5186 2382 5224 2416
rect 5258 2382 5405 2416
rect 5005 2343 5405 2382
rect 5005 2309 5152 2343
rect 5186 2309 5224 2343
rect 5258 2309 5405 2343
rect 5005 2270 5405 2309
rect 5005 2236 5152 2270
rect 5186 2236 5224 2270
rect 5258 2236 5405 2270
rect 5005 2197 5405 2236
rect 5005 2163 5152 2197
rect 5186 2163 5224 2197
rect 5258 2163 5405 2197
rect 5005 2124 5405 2163
rect 5005 2090 5152 2124
rect 5186 2090 5224 2124
rect 5258 2090 5405 2124
rect 5005 2051 5405 2090
rect 5005 2017 5152 2051
rect 5186 2017 5224 2051
rect 5258 2017 5405 2051
rect 5005 1978 5405 2017
rect 5005 1944 5152 1978
rect 5186 1944 5224 1978
rect 5258 1944 5405 1978
rect 5005 1905 5405 1944
rect 5005 1871 5152 1905
rect 5186 1871 5224 1905
rect 5258 1871 5405 1905
rect 5005 1832 5405 1871
rect 5005 1798 5152 1832
rect 5186 1798 5224 1832
rect 5258 1798 5405 1832
rect 5005 1759 5405 1798
rect 5005 1725 5152 1759
rect 5186 1725 5224 1759
rect 5258 1725 5405 1759
rect 5005 1686 5405 1725
rect 5005 1652 5152 1686
rect 5186 1652 5224 1686
rect 5258 1652 5405 1686
rect 5005 1613 5405 1652
rect 5005 1579 5152 1613
rect 5186 1579 5224 1613
rect 5258 1579 5405 1613
rect 5005 1540 5405 1579
rect 5005 1506 5152 1540
rect 5186 1506 5224 1540
rect 5258 1506 5405 1540
rect 5005 1466 5405 1506
rect 5005 1432 5152 1466
rect 5186 1432 5224 1466
rect 5258 1432 5405 1466
rect 5005 1392 5405 1432
rect 5005 1358 5152 1392
rect 5186 1358 5224 1392
rect 5258 1358 5405 1392
rect 5005 1318 5405 1358
rect 5005 1284 5152 1318
rect 5186 1284 5224 1318
rect 5258 1284 5405 1318
rect 5005 1244 5405 1284
rect 5005 1210 5152 1244
rect 5186 1210 5224 1244
rect 5258 1210 5405 1244
rect 5005 1170 5405 1210
rect 5005 1136 5152 1170
rect 5186 1136 5224 1170
rect 5258 1136 5405 1170
rect 5005 1096 5405 1136
rect 5005 1062 5152 1096
rect 5186 1062 5224 1096
rect 5258 1062 5405 1096
rect 5005 1022 5405 1062
rect 5005 988 5152 1022
rect 5186 988 5224 1022
rect 5258 988 5405 1022
rect 5005 948 5405 988
rect 5005 914 5152 948
rect 5186 914 5224 948
rect 5258 914 5405 948
rect 5005 874 5405 914
rect 5005 840 5152 874
rect 5186 840 5224 874
rect 5258 840 5405 874
rect 5005 800 5405 840
rect 5005 766 5152 800
rect 5186 766 5224 800
rect 5258 766 5405 800
rect 5005 726 5405 766
rect 5005 692 5152 726
rect 5186 692 5224 726
rect 5258 692 5405 726
rect 5005 652 5405 692
rect 5005 618 5152 652
rect 5186 618 5224 652
rect 5258 618 5405 652
rect 5005 578 5405 618
rect 5005 544 5152 578
rect 5186 544 5224 578
rect 5258 544 5405 578
rect 5005 504 5405 544
rect 5005 470 5152 504
rect 5186 470 5224 504
rect 5258 470 5405 504
rect 5005 430 5405 470
rect 5005 396 5152 430
rect 5186 396 5224 430
rect 5258 396 5405 430
rect 5005 356 5405 396
rect 5005 322 5152 356
rect 5186 322 5224 356
rect 5258 322 5405 356
rect 5005 282 5405 322
rect 5005 248 5152 282
rect 5186 248 5224 282
rect 5258 248 5405 282
rect 5005 208 5405 248
rect 5005 174 5152 208
rect 5186 174 5224 208
rect 5258 174 5405 208
rect 5005 134 5405 174
rect 5005 100 5152 134
rect 5186 100 5224 134
rect 5258 100 5405 134
rect 5005 47 5405 100
tri 5005 42 5010 47 ne
rect 5010 42 5400 47
tri 5400 42 5405 47 nw
tri 5517 3053 5564 3100 se
rect 5564 3053 5670 3100
tri 5670 3053 5717 3100 sw
rect 5517 3000 5717 3053
rect 5517 2966 5564 3000
rect 5598 2966 5636 3000
rect 5670 2966 5717 3000
rect 5517 2927 5717 2966
rect 5517 2893 5564 2927
rect 5598 2893 5636 2927
rect 5670 2893 5717 2927
rect 5517 2854 5717 2893
rect 5517 2820 5564 2854
rect 5598 2820 5636 2854
rect 5670 2820 5717 2854
rect 5517 2781 5717 2820
rect 5517 2747 5564 2781
rect 5598 2747 5636 2781
rect 5670 2747 5717 2781
rect 5517 2708 5717 2747
rect 5517 2674 5564 2708
rect 5598 2674 5636 2708
rect 5670 2674 5717 2708
rect 5517 2635 5717 2674
rect 5517 2601 5564 2635
rect 5598 2601 5636 2635
rect 5670 2601 5717 2635
rect 5517 2562 5717 2601
rect 5517 2528 5564 2562
rect 5598 2528 5636 2562
rect 5670 2528 5717 2562
rect 5517 2489 5717 2528
rect 5517 2455 5564 2489
rect 5598 2455 5636 2489
rect 5670 2455 5717 2489
rect 5517 2416 5717 2455
rect 5517 2382 5564 2416
rect 5598 2382 5636 2416
rect 5670 2382 5717 2416
rect 5517 2343 5717 2382
rect 5517 2309 5564 2343
rect 5598 2309 5636 2343
rect 5670 2309 5717 2343
rect 5517 2270 5717 2309
rect 5517 2236 5564 2270
rect 5598 2236 5636 2270
rect 5670 2236 5717 2270
rect 5517 2197 5717 2236
rect 5517 2163 5564 2197
rect 5598 2163 5636 2197
rect 5670 2163 5717 2197
rect 5517 2124 5717 2163
rect 5517 2090 5564 2124
rect 5598 2090 5636 2124
rect 5670 2090 5717 2124
rect 5517 2051 5717 2090
rect 5517 2017 5564 2051
rect 5598 2017 5636 2051
rect 5670 2017 5717 2051
rect 5517 1978 5717 2017
rect 5517 1944 5564 1978
rect 5598 1944 5636 1978
rect 5670 1944 5717 1978
rect 5517 1905 5717 1944
rect 5517 1871 5564 1905
rect 5598 1871 5636 1905
rect 5670 1871 5717 1905
rect 5517 1832 5717 1871
rect 5517 1798 5564 1832
rect 5598 1798 5636 1832
rect 5670 1798 5717 1832
rect 5517 1759 5717 1798
rect 5517 1725 5564 1759
rect 5598 1725 5636 1759
rect 5670 1725 5717 1759
rect 5517 1686 5717 1725
rect 5517 1652 5564 1686
rect 5598 1652 5636 1686
rect 5670 1652 5717 1686
rect 5517 1613 5717 1652
rect 5517 1579 5564 1613
rect 5598 1579 5636 1613
rect 5670 1579 5717 1613
rect 5517 1540 5717 1579
rect 5517 1506 5564 1540
rect 5598 1506 5636 1540
rect 5670 1506 5717 1540
rect 5517 1466 5717 1506
rect 5517 1432 5564 1466
rect 5598 1432 5636 1466
rect 5670 1432 5717 1466
rect 5517 1392 5717 1432
rect 5517 1358 5564 1392
rect 5598 1358 5636 1392
rect 5670 1358 5717 1392
rect 5517 1318 5717 1358
rect 5517 1284 5564 1318
rect 5598 1284 5636 1318
rect 5670 1284 5717 1318
rect 5517 1244 5717 1284
rect 5517 1210 5564 1244
rect 5598 1210 5636 1244
rect 5670 1210 5717 1244
rect 5517 1170 5717 1210
rect 5517 1136 5564 1170
rect 5598 1136 5636 1170
rect 5670 1136 5717 1170
rect 5517 1096 5717 1136
rect 5517 1062 5564 1096
rect 5598 1062 5636 1096
rect 5670 1062 5717 1096
rect 5517 1022 5717 1062
rect 5517 988 5564 1022
rect 5598 988 5636 1022
rect 5670 988 5717 1022
rect 5517 948 5717 988
rect 5517 914 5564 948
rect 5598 914 5636 948
rect 5670 914 5717 948
rect 5517 874 5717 914
rect 5517 840 5564 874
rect 5598 840 5636 874
rect 5670 840 5717 874
rect 5517 800 5717 840
rect 5517 766 5564 800
rect 5598 766 5636 800
rect 5670 766 5717 800
rect 5517 726 5717 766
rect 5517 692 5564 726
rect 5598 692 5636 726
rect 5670 692 5717 726
rect 5517 652 5717 692
rect 5517 618 5564 652
rect 5598 618 5636 652
rect 5670 618 5717 652
rect 5517 578 5717 618
rect 5517 544 5564 578
rect 5598 544 5636 578
rect 5670 544 5717 578
rect 5517 504 5717 544
rect 5517 470 5564 504
rect 5598 470 5636 504
rect 5670 470 5717 504
rect 5517 430 5717 470
rect 5517 396 5564 430
rect 5598 396 5636 430
rect 5670 396 5717 430
rect 5517 356 5717 396
rect 5517 322 5564 356
rect 5598 322 5636 356
rect 5670 322 5717 356
rect 5517 282 5717 322
rect 5517 248 5564 282
rect 5598 248 5636 282
rect 5670 248 5717 282
rect 5517 208 5717 248
rect 5517 174 5564 208
rect 5598 174 5636 208
rect 5670 174 5717 208
rect 5517 134 5717 174
rect 5517 100 5564 134
rect 5598 100 5636 134
rect 5670 100 5717 134
rect 5517 47 5717 100
tri 5517 42 5522 47 ne
rect 5522 42 5712 47
tri 5712 42 5717 47 nw
tri 5829 3053 5876 3100 se
rect 5876 3053 6182 3100
tri 6182 3053 6229 3100 sw
rect 5829 3000 6229 3053
rect 5829 2966 5976 3000
rect 6010 2966 6048 3000
rect 6082 2966 6229 3000
rect 5829 2927 6229 2966
rect 5829 2893 5976 2927
rect 6010 2893 6048 2927
rect 6082 2893 6229 2927
rect 5829 2854 6229 2893
rect 5829 2820 5976 2854
rect 6010 2820 6048 2854
rect 6082 2820 6229 2854
rect 5829 2781 6229 2820
rect 5829 2747 5976 2781
rect 6010 2747 6048 2781
rect 6082 2747 6229 2781
rect 5829 2708 6229 2747
rect 5829 2674 5976 2708
rect 6010 2674 6048 2708
rect 6082 2674 6229 2708
rect 5829 2635 6229 2674
rect 5829 2601 5976 2635
rect 6010 2601 6048 2635
rect 6082 2601 6229 2635
rect 5829 2562 6229 2601
rect 5829 2528 5976 2562
rect 6010 2528 6048 2562
rect 6082 2528 6229 2562
rect 5829 2489 6229 2528
rect 5829 2455 5976 2489
rect 6010 2455 6048 2489
rect 6082 2455 6229 2489
rect 5829 2416 6229 2455
rect 5829 2382 5976 2416
rect 6010 2382 6048 2416
rect 6082 2382 6229 2416
rect 5829 2343 6229 2382
rect 5829 2309 5976 2343
rect 6010 2309 6048 2343
rect 6082 2309 6229 2343
rect 5829 2270 6229 2309
rect 5829 2236 5976 2270
rect 6010 2236 6048 2270
rect 6082 2236 6229 2270
rect 5829 2197 6229 2236
rect 5829 2163 5976 2197
rect 6010 2163 6048 2197
rect 6082 2163 6229 2197
rect 5829 2124 6229 2163
rect 5829 2090 5976 2124
rect 6010 2090 6048 2124
rect 6082 2090 6229 2124
rect 5829 2051 6229 2090
rect 5829 2017 5976 2051
rect 6010 2017 6048 2051
rect 6082 2017 6229 2051
rect 5829 1978 6229 2017
rect 5829 1944 5976 1978
rect 6010 1944 6048 1978
rect 6082 1944 6229 1978
rect 5829 1905 6229 1944
rect 5829 1871 5976 1905
rect 6010 1871 6048 1905
rect 6082 1871 6229 1905
rect 5829 1832 6229 1871
rect 5829 1798 5976 1832
rect 6010 1798 6048 1832
rect 6082 1798 6229 1832
rect 5829 1759 6229 1798
rect 5829 1725 5976 1759
rect 6010 1725 6048 1759
rect 6082 1725 6229 1759
rect 5829 1686 6229 1725
rect 5829 1652 5976 1686
rect 6010 1652 6048 1686
rect 6082 1652 6229 1686
rect 5829 1613 6229 1652
rect 5829 1579 5976 1613
rect 6010 1579 6048 1613
rect 6082 1579 6229 1613
rect 5829 1540 6229 1579
rect 5829 1506 5976 1540
rect 6010 1506 6048 1540
rect 6082 1506 6229 1540
rect 5829 1466 6229 1506
rect 5829 1432 5976 1466
rect 6010 1432 6048 1466
rect 6082 1432 6229 1466
rect 5829 1392 6229 1432
rect 5829 1358 5976 1392
rect 6010 1358 6048 1392
rect 6082 1358 6229 1392
rect 5829 1318 6229 1358
rect 5829 1284 5976 1318
rect 6010 1284 6048 1318
rect 6082 1284 6229 1318
rect 5829 1244 6229 1284
rect 5829 1210 5976 1244
rect 6010 1210 6048 1244
rect 6082 1210 6229 1244
rect 5829 1170 6229 1210
rect 5829 1136 5976 1170
rect 6010 1136 6048 1170
rect 6082 1136 6229 1170
rect 5829 1096 6229 1136
rect 5829 1062 5976 1096
rect 6010 1062 6048 1096
rect 6082 1062 6229 1096
rect 5829 1022 6229 1062
rect 5829 988 5976 1022
rect 6010 988 6048 1022
rect 6082 988 6229 1022
rect 5829 948 6229 988
rect 5829 914 5976 948
rect 6010 914 6048 948
rect 6082 914 6229 948
rect 5829 874 6229 914
rect 5829 840 5976 874
rect 6010 840 6048 874
rect 6082 840 6229 874
rect 5829 800 6229 840
rect 5829 766 5976 800
rect 6010 766 6048 800
rect 6082 766 6229 800
rect 5829 726 6229 766
rect 5829 692 5976 726
rect 6010 692 6048 726
rect 6082 692 6229 726
rect 5829 652 6229 692
rect 5829 618 5976 652
rect 6010 618 6048 652
rect 6082 618 6229 652
rect 5829 578 6229 618
rect 5829 544 5976 578
rect 6010 544 6048 578
rect 6082 544 6229 578
rect 5829 504 6229 544
rect 5829 470 5976 504
rect 6010 470 6048 504
rect 6082 470 6229 504
rect 5829 430 6229 470
rect 5829 396 5976 430
rect 6010 396 6048 430
rect 6082 396 6229 430
rect 5829 356 6229 396
rect 5829 322 5976 356
rect 6010 322 6048 356
rect 6082 322 6229 356
rect 5829 282 6229 322
rect 5829 248 5976 282
rect 6010 248 6048 282
rect 6082 248 6229 282
rect 5829 208 6229 248
rect 5829 174 5976 208
rect 6010 174 6048 208
rect 6082 174 6229 208
rect 5829 134 6229 174
rect 5829 100 5976 134
rect 6010 100 6048 134
rect 6082 100 6229 134
rect 5829 47 6229 100
tri 5829 42 5834 47 ne
rect 5834 42 6224 47
tri 6224 42 6229 47 nw
tri 6341 3053 6388 3100 se
rect 6388 3053 6494 3100
tri 6494 3053 6541 3100 sw
rect 6341 3000 6541 3053
rect 6341 2966 6388 3000
rect 6422 2966 6460 3000
rect 6494 2966 6541 3000
rect 6341 2927 6541 2966
rect 6341 2893 6388 2927
rect 6422 2893 6460 2927
rect 6494 2893 6541 2927
rect 6341 2854 6541 2893
rect 6341 2820 6388 2854
rect 6422 2820 6460 2854
rect 6494 2820 6541 2854
rect 6341 2781 6541 2820
rect 6341 2747 6388 2781
rect 6422 2747 6460 2781
rect 6494 2747 6541 2781
rect 6341 2708 6541 2747
rect 6341 2674 6388 2708
rect 6422 2674 6460 2708
rect 6494 2674 6541 2708
rect 6341 2635 6541 2674
rect 6341 2601 6388 2635
rect 6422 2601 6460 2635
rect 6494 2601 6541 2635
rect 6341 2562 6541 2601
rect 6341 2528 6388 2562
rect 6422 2528 6460 2562
rect 6494 2528 6541 2562
rect 6341 2489 6541 2528
rect 6341 2455 6388 2489
rect 6422 2455 6460 2489
rect 6494 2455 6541 2489
rect 6341 2416 6541 2455
rect 6341 2382 6388 2416
rect 6422 2382 6460 2416
rect 6494 2382 6541 2416
rect 6341 2343 6541 2382
rect 6341 2309 6388 2343
rect 6422 2309 6460 2343
rect 6494 2309 6541 2343
rect 6341 2270 6541 2309
rect 6341 2236 6388 2270
rect 6422 2236 6460 2270
rect 6494 2236 6541 2270
rect 6341 2197 6541 2236
rect 6341 2163 6388 2197
rect 6422 2163 6460 2197
rect 6494 2163 6541 2197
rect 6341 2124 6541 2163
rect 6341 2090 6388 2124
rect 6422 2090 6460 2124
rect 6494 2090 6541 2124
rect 6341 2051 6541 2090
rect 6341 2017 6388 2051
rect 6422 2017 6460 2051
rect 6494 2017 6541 2051
rect 6341 1978 6541 2017
rect 6341 1944 6388 1978
rect 6422 1944 6460 1978
rect 6494 1944 6541 1978
rect 6341 1905 6541 1944
rect 6341 1871 6388 1905
rect 6422 1871 6460 1905
rect 6494 1871 6541 1905
rect 6341 1832 6541 1871
rect 6341 1798 6388 1832
rect 6422 1798 6460 1832
rect 6494 1798 6541 1832
rect 6341 1759 6541 1798
rect 6341 1725 6388 1759
rect 6422 1725 6460 1759
rect 6494 1725 6541 1759
rect 6341 1686 6541 1725
rect 6341 1652 6388 1686
rect 6422 1652 6460 1686
rect 6494 1652 6541 1686
rect 6341 1613 6541 1652
rect 6341 1579 6388 1613
rect 6422 1579 6460 1613
rect 6494 1579 6541 1613
rect 6341 1540 6541 1579
rect 6341 1506 6388 1540
rect 6422 1506 6460 1540
rect 6494 1506 6541 1540
rect 6341 1466 6541 1506
rect 6341 1432 6388 1466
rect 6422 1432 6460 1466
rect 6494 1432 6541 1466
rect 6341 1392 6541 1432
rect 6341 1358 6388 1392
rect 6422 1358 6460 1392
rect 6494 1358 6541 1392
rect 6341 1318 6541 1358
rect 6341 1284 6388 1318
rect 6422 1284 6460 1318
rect 6494 1284 6541 1318
rect 6341 1244 6541 1284
rect 6341 1210 6388 1244
rect 6422 1210 6460 1244
rect 6494 1210 6541 1244
rect 6341 1170 6541 1210
rect 6341 1136 6388 1170
rect 6422 1136 6460 1170
rect 6494 1136 6541 1170
rect 6341 1096 6541 1136
rect 6341 1062 6388 1096
rect 6422 1062 6460 1096
rect 6494 1062 6541 1096
rect 6341 1022 6541 1062
rect 6341 988 6388 1022
rect 6422 988 6460 1022
rect 6494 988 6541 1022
rect 6341 948 6541 988
rect 6341 914 6388 948
rect 6422 914 6460 948
rect 6494 914 6541 948
rect 6341 874 6541 914
rect 6341 840 6388 874
rect 6422 840 6460 874
rect 6494 840 6541 874
rect 6341 800 6541 840
rect 6341 766 6388 800
rect 6422 766 6460 800
rect 6494 766 6541 800
rect 6341 726 6541 766
rect 6341 692 6388 726
rect 6422 692 6460 726
rect 6494 692 6541 726
rect 6341 652 6541 692
rect 6341 618 6388 652
rect 6422 618 6460 652
rect 6494 618 6541 652
rect 6341 578 6541 618
rect 6341 544 6388 578
rect 6422 544 6460 578
rect 6494 544 6541 578
rect 6341 504 6541 544
rect 6341 470 6388 504
rect 6422 470 6460 504
rect 6494 470 6541 504
rect 6341 430 6541 470
rect 6341 396 6388 430
rect 6422 396 6460 430
rect 6494 396 6541 430
rect 6341 356 6541 396
rect 6341 322 6388 356
rect 6422 322 6460 356
rect 6494 322 6541 356
rect 6341 282 6541 322
rect 6341 248 6388 282
rect 6422 248 6460 282
rect 6494 248 6541 282
rect 6341 208 6541 248
rect 6341 174 6388 208
rect 6422 174 6460 208
rect 6494 174 6541 208
rect 6341 134 6541 174
rect 6341 100 6388 134
rect 6422 100 6460 134
rect 6494 100 6541 134
rect 6341 47 6541 100
tri 6341 42 6346 47 ne
rect 6346 42 6536 47
tri 6536 42 6541 47 nw
tri 6653 3053 6700 3100 se
rect 6700 3053 7006 3100
tri 7006 3053 7053 3100 sw
rect 6653 3000 7053 3053
rect 6653 2966 6800 3000
rect 6834 2966 6872 3000
rect 6906 2966 7053 3000
rect 6653 2927 7053 2966
rect 6653 2893 6800 2927
rect 6834 2893 6872 2927
rect 6906 2893 7053 2927
rect 6653 2854 7053 2893
rect 6653 2820 6800 2854
rect 6834 2820 6872 2854
rect 6906 2820 7053 2854
rect 6653 2781 7053 2820
rect 6653 2747 6800 2781
rect 6834 2747 6872 2781
rect 6906 2747 7053 2781
rect 6653 2708 7053 2747
rect 6653 2674 6800 2708
rect 6834 2674 6872 2708
rect 6906 2674 7053 2708
rect 6653 2635 7053 2674
rect 6653 2601 6800 2635
rect 6834 2601 6872 2635
rect 6906 2601 7053 2635
rect 6653 2562 7053 2601
rect 6653 2528 6800 2562
rect 6834 2528 6872 2562
rect 6906 2528 7053 2562
rect 6653 2489 7053 2528
rect 6653 2455 6800 2489
rect 6834 2455 6872 2489
rect 6906 2455 7053 2489
rect 6653 2416 7053 2455
rect 6653 2382 6800 2416
rect 6834 2382 6872 2416
rect 6906 2382 7053 2416
rect 6653 2343 7053 2382
rect 6653 2309 6800 2343
rect 6834 2309 6872 2343
rect 6906 2309 7053 2343
rect 6653 2270 7053 2309
rect 6653 2236 6800 2270
rect 6834 2236 6872 2270
rect 6906 2236 7053 2270
rect 6653 2197 7053 2236
rect 6653 2163 6800 2197
rect 6834 2163 6872 2197
rect 6906 2163 7053 2197
rect 6653 2124 7053 2163
rect 6653 2090 6800 2124
rect 6834 2090 6872 2124
rect 6906 2090 7053 2124
rect 6653 2051 7053 2090
rect 6653 2017 6800 2051
rect 6834 2017 6872 2051
rect 6906 2017 7053 2051
rect 6653 1978 7053 2017
rect 6653 1944 6800 1978
rect 6834 1944 6872 1978
rect 6906 1944 7053 1978
rect 6653 1905 7053 1944
rect 6653 1871 6800 1905
rect 6834 1871 6872 1905
rect 6906 1871 7053 1905
rect 6653 1832 7053 1871
rect 6653 1798 6800 1832
rect 6834 1798 6872 1832
rect 6906 1798 7053 1832
rect 6653 1759 7053 1798
rect 6653 1725 6800 1759
rect 6834 1725 6872 1759
rect 6906 1725 7053 1759
rect 6653 1686 7053 1725
rect 6653 1652 6800 1686
rect 6834 1652 6872 1686
rect 6906 1652 7053 1686
rect 6653 1613 7053 1652
rect 6653 1579 6800 1613
rect 6834 1579 6872 1613
rect 6906 1579 7053 1613
rect 6653 1540 7053 1579
rect 6653 1506 6800 1540
rect 6834 1506 6872 1540
rect 6906 1506 7053 1540
rect 6653 1466 7053 1506
rect 6653 1432 6800 1466
rect 6834 1432 6872 1466
rect 6906 1432 7053 1466
rect 6653 1392 7053 1432
rect 6653 1358 6800 1392
rect 6834 1358 6872 1392
rect 6906 1358 7053 1392
rect 6653 1318 7053 1358
rect 6653 1284 6800 1318
rect 6834 1284 6872 1318
rect 6906 1284 7053 1318
rect 6653 1244 7053 1284
rect 6653 1210 6800 1244
rect 6834 1210 6872 1244
rect 6906 1210 7053 1244
rect 6653 1170 7053 1210
rect 6653 1136 6800 1170
rect 6834 1136 6872 1170
rect 6906 1136 7053 1170
rect 6653 1096 7053 1136
rect 6653 1062 6800 1096
rect 6834 1062 6872 1096
rect 6906 1062 7053 1096
rect 6653 1022 7053 1062
rect 6653 988 6800 1022
rect 6834 988 6872 1022
rect 6906 988 7053 1022
rect 6653 948 7053 988
rect 6653 914 6800 948
rect 6834 914 6872 948
rect 6906 914 7053 948
rect 6653 874 7053 914
rect 6653 840 6800 874
rect 6834 840 6872 874
rect 6906 840 7053 874
rect 6653 800 7053 840
rect 6653 766 6800 800
rect 6834 766 6872 800
rect 6906 766 7053 800
rect 6653 726 7053 766
rect 6653 692 6800 726
rect 6834 692 6872 726
rect 6906 692 7053 726
rect 6653 652 7053 692
rect 6653 618 6800 652
rect 6834 618 6872 652
rect 6906 618 7053 652
rect 6653 578 7053 618
rect 6653 544 6800 578
rect 6834 544 6872 578
rect 6906 544 7053 578
rect 6653 504 7053 544
rect 6653 470 6800 504
rect 6834 470 6872 504
rect 6906 470 7053 504
rect 6653 430 7053 470
rect 6653 396 6800 430
rect 6834 396 6872 430
rect 6906 396 7053 430
rect 6653 356 7053 396
rect 6653 322 6800 356
rect 6834 322 6872 356
rect 6906 322 7053 356
rect 6653 282 7053 322
rect 6653 248 6800 282
rect 6834 248 6872 282
rect 6906 248 7053 282
rect 6653 208 7053 248
rect 6653 174 6800 208
rect 6834 174 6872 208
rect 6906 174 7053 208
rect 6653 134 7053 174
rect 6653 100 6800 134
rect 6834 100 6872 134
rect 6906 100 7053 134
rect 6653 47 7053 100
tri 6653 42 6658 47 ne
rect 6658 42 7048 47
tri 7048 42 7053 47 nw
tri 7165 3053 7212 3100 se
rect 7212 3053 7318 3100
tri 7318 3053 7365 3100 sw
rect 7165 3000 7365 3053
rect 7165 2966 7212 3000
rect 7246 2966 7284 3000
rect 7318 2966 7365 3000
rect 7165 2927 7365 2966
rect 7165 2893 7212 2927
rect 7246 2893 7284 2927
rect 7318 2893 7365 2927
rect 7165 2854 7365 2893
rect 7165 2820 7212 2854
rect 7246 2820 7284 2854
rect 7318 2820 7365 2854
rect 7165 2781 7365 2820
rect 7165 2747 7212 2781
rect 7246 2747 7284 2781
rect 7318 2747 7365 2781
rect 7165 2708 7365 2747
rect 7165 2674 7212 2708
rect 7246 2674 7284 2708
rect 7318 2674 7365 2708
rect 7165 2635 7365 2674
rect 7165 2601 7212 2635
rect 7246 2601 7284 2635
rect 7318 2601 7365 2635
rect 7165 2562 7365 2601
rect 7165 2528 7212 2562
rect 7246 2528 7284 2562
rect 7318 2528 7365 2562
rect 7165 2489 7365 2528
rect 7165 2455 7212 2489
rect 7246 2455 7284 2489
rect 7318 2455 7365 2489
rect 7165 2416 7365 2455
rect 7165 2382 7212 2416
rect 7246 2382 7284 2416
rect 7318 2382 7365 2416
rect 7165 2343 7365 2382
rect 7165 2309 7212 2343
rect 7246 2309 7284 2343
rect 7318 2309 7365 2343
rect 7165 2270 7365 2309
rect 7165 2236 7212 2270
rect 7246 2236 7284 2270
rect 7318 2236 7365 2270
rect 7165 2197 7365 2236
rect 7165 2163 7212 2197
rect 7246 2163 7284 2197
rect 7318 2163 7365 2197
rect 7165 2124 7365 2163
rect 7165 2090 7212 2124
rect 7246 2090 7284 2124
rect 7318 2090 7365 2124
rect 7165 2051 7365 2090
rect 7165 2017 7212 2051
rect 7246 2017 7284 2051
rect 7318 2017 7365 2051
rect 7165 1978 7365 2017
rect 7165 1944 7212 1978
rect 7246 1944 7284 1978
rect 7318 1944 7365 1978
rect 7165 1905 7365 1944
rect 7165 1871 7212 1905
rect 7246 1871 7284 1905
rect 7318 1871 7365 1905
rect 7165 1832 7365 1871
rect 7165 1798 7212 1832
rect 7246 1798 7284 1832
rect 7318 1798 7365 1832
rect 7165 1759 7365 1798
rect 7165 1725 7212 1759
rect 7246 1725 7284 1759
rect 7318 1725 7365 1759
rect 7165 1686 7365 1725
rect 7165 1652 7212 1686
rect 7246 1652 7284 1686
rect 7318 1652 7365 1686
rect 7165 1613 7365 1652
rect 7165 1579 7212 1613
rect 7246 1579 7284 1613
rect 7318 1579 7365 1613
rect 7165 1540 7365 1579
rect 7165 1506 7212 1540
rect 7246 1506 7284 1540
rect 7318 1506 7365 1540
rect 7165 1466 7365 1506
rect 7165 1432 7212 1466
rect 7246 1432 7284 1466
rect 7318 1432 7365 1466
rect 7165 1392 7365 1432
rect 7165 1358 7212 1392
rect 7246 1358 7284 1392
rect 7318 1358 7365 1392
rect 7165 1318 7365 1358
rect 7165 1284 7212 1318
rect 7246 1284 7284 1318
rect 7318 1284 7365 1318
rect 7165 1244 7365 1284
rect 7165 1210 7212 1244
rect 7246 1210 7284 1244
rect 7318 1210 7365 1244
rect 7165 1170 7365 1210
rect 7165 1136 7212 1170
rect 7246 1136 7284 1170
rect 7318 1136 7365 1170
rect 7165 1096 7365 1136
rect 7165 1062 7212 1096
rect 7246 1062 7284 1096
rect 7318 1062 7365 1096
rect 7165 1022 7365 1062
rect 7165 988 7212 1022
rect 7246 988 7284 1022
rect 7318 988 7365 1022
rect 7165 948 7365 988
rect 7165 914 7212 948
rect 7246 914 7284 948
rect 7318 914 7365 948
rect 7165 874 7365 914
rect 7165 840 7212 874
rect 7246 840 7284 874
rect 7318 840 7365 874
rect 7165 800 7365 840
rect 7165 766 7212 800
rect 7246 766 7284 800
rect 7318 766 7365 800
rect 7165 726 7365 766
rect 7165 692 7212 726
rect 7246 692 7284 726
rect 7318 692 7365 726
rect 7165 652 7365 692
rect 7165 618 7212 652
rect 7246 618 7284 652
rect 7318 618 7365 652
rect 7165 578 7365 618
rect 7165 544 7212 578
rect 7246 544 7284 578
rect 7318 544 7365 578
rect 7165 504 7365 544
rect 7165 470 7212 504
rect 7246 470 7284 504
rect 7318 470 7365 504
rect 7165 430 7365 470
rect 7165 396 7212 430
rect 7246 396 7284 430
rect 7318 396 7365 430
rect 7165 356 7365 396
rect 7165 322 7212 356
rect 7246 322 7284 356
rect 7318 322 7365 356
rect 7165 282 7365 322
rect 7165 248 7212 282
rect 7246 248 7284 282
rect 7318 248 7365 282
rect 7165 208 7365 248
rect 7165 174 7212 208
rect 7246 174 7284 208
rect 7318 174 7365 208
rect 7165 134 7365 174
rect 7165 100 7212 134
rect 7246 100 7284 134
rect 7318 100 7365 134
rect 7165 47 7365 100
tri 7165 42 7170 47 ne
rect 7170 42 7360 47
tri 7360 42 7365 47 nw
tri 7477 3053 7524 3100 se
rect 7524 3053 7830 3100
tri 7830 3053 7877 3100 sw
rect 7477 3000 7877 3053
rect 7477 2966 7624 3000
rect 7658 2966 7696 3000
rect 7730 2966 7877 3000
rect 7477 2927 7877 2966
rect 7477 2893 7624 2927
rect 7658 2893 7696 2927
rect 7730 2893 7877 2927
rect 7477 2854 7877 2893
rect 7477 2820 7624 2854
rect 7658 2820 7696 2854
rect 7730 2820 7877 2854
rect 7477 2781 7877 2820
rect 7477 2747 7624 2781
rect 7658 2747 7696 2781
rect 7730 2747 7877 2781
rect 7477 2708 7877 2747
rect 7477 2674 7624 2708
rect 7658 2674 7696 2708
rect 7730 2674 7877 2708
rect 7477 2635 7877 2674
rect 7477 2601 7624 2635
rect 7658 2601 7696 2635
rect 7730 2601 7877 2635
rect 7477 2562 7877 2601
rect 7477 2528 7624 2562
rect 7658 2528 7696 2562
rect 7730 2528 7877 2562
rect 7477 2489 7877 2528
rect 7477 2455 7624 2489
rect 7658 2455 7696 2489
rect 7730 2455 7877 2489
rect 7477 2416 7877 2455
rect 7477 2382 7624 2416
rect 7658 2382 7696 2416
rect 7730 2382 7877 2416
rect 7477 2343 7877 2382
rect 7477 2309 7624 2343
rect 7658 2309 7696 2343
rect 7730 2309 7877 2343
rect 7477 2270 7877 2309
rect 7477 2236 7624 2270
rect 7658 2236 7696 2270
rect 7730 2236 7877 2270
rect 7477 2197 7877 2236
rect 7477 2163 7624 2197
rect 7658 2163 7696 2197
rect 7730 2163 7877 2197
rect 7477 2124 7877 2163
rect 7477 2090 7624 2124
rect 7658 2090 7696 2124
rect 7730 2090 7877 2124
rect 7477 2051 7877 2090
rect 7477 2017 7624 2051
rect 7658 2017 7696 2051
rect 7730 2017 7877 2051
rect 7477 1978 7877 2017
rect 7477 1944 7624 1978
rect 7658 1944 7696 1978
rect 7730 1944 7877 1978
rect 7477 1905 7877 1944
rect 7477 1871 7624 1905
rect 7658 1871 7696 1905
rect 7730 1871 7877 1905
rect 7477 1832 7877 1871
rect 7477 1798 7624 1832
rect 7658 1798 7696 1832
rect 7730 1798 7877 1832
rect 7477 1759 7877 1798
rect 7477 1725 7624 1759
rect 7658 1725 7696 1759
rect 7730 1725 7877 1759
rect 7477 1686 7877 1725
rect 7477 1652 7624 1686
rect 7658 1652 7696 1686
rect 7730 1652 7877 1686
rect 7477 1613 7877 1652
rect 7477 1579 7624 1613
rect 7658 1579 7696 1613
rect 7730 1579 7877 1613
rect 7477 1540 7877 1579
rect 7477 1506 7624 1540
rect 7658 1506 7696 1540
rect 7730 1506 7877 1540
rect 7477 1466 7877 1506
rect 7477 1432 7624 1466
rect 7658 1432 7696 1466
rect 7730 1432 7877 1466
rect 7477 1392 7877 1432
rect 7477 1358 7624 1392
rect 7658 1358 7696 1392
rect 7730 1358 7877 1392
rect 7477 1318 7877 1358
rect 7477 1284 7624 1318
rect 7658 1284 7696 1318
rect 7730 1284 7877 1318
rect 7477 1244 7877 1284
rect 7477 1210 7624 1244
rect 7658 1210 7696 1244
rect 7730 1210 7877 1244
rect 7477 1170 7877 1210
rect 7477 1136 7624 1170
rect 7658 1136 7696 1170
rect 7730 1136 7877 1170
rect 7477 1096 7877 1136
rect 7477 1062 7624 1096
rect 7658 1062 7696 1096
rect 7730 1062 7877 1096
rect 7477 1022 7877 1062
rect 7477 988 7624 1022
rect 7658 988 7696 1022
rect 7730 988 7877 1022
rect 7477 948 7877 988
rect 7477 914 7624 948
rect 7658 914 7696 948
rect 7730 914 7877 948
rect 7477 874 7877 914
rect 7477 840 7624 874
rect 7658 840 7696 874
rect 7730 840 7877 874
rect 7477 800 7877 840
rect 7477 766 7624 800
rect 7658 766 7696 800
rect 7730 766 7877 800
rect 7477 726 7877 766
rect 7477 692 7624 726
rect 7658 692 7696 726
rect 7730 692 7877 726
rect 7477 652 7877 692
rect 7477 618 7624 652
rect 7658 618 7696 652
rect 7730 618 7877 652
rect 7477 578 7877 618
rect 7477 544 7624 578
rect 7658 544 7696 578
rect 7730 544 7877 578
rect 7477 504 7877 544
rect 7477 470 7624 504
rect 7658 470 7696 504
rect 7730 470 7877 504
rect 7477 430 7877 470
rect 7477 396 7624 430
rect 7658 396 7696 430
rect 7730 396 7877 430
rect 7477 356 7877 396
rect 7477 322 7624 356
rect 7658 322 7696 356
rect 7730 322 7877 356
rect 7477 282 7877 322
rect 7477 248 7624 282
rect 7658 248 7696 282
rect 7730 248 7877 282
rect 7477 208 7877 248
rect 7477 174 7624 208
rect 7658 174 7696 208
rect 7730 174 7877 208
rect 7477 134 7877 174
rect 7477 100 7624 134
rect 7658 100 7696 134
rect 7730 100 7877 134
rect 7477 47 7877 100
tri 7477 42 7482 47 ne
rect 7482 42 7872 47
tri 7872 42 7877 47 nw
tri 7989 3053 8036 3100 se
rect 8036 3053 8142 3100
tri 8142 3053 8189 3100 sw
rect 7989 3000 8189 3053
rect 7989 2966 8036 3000
rect 8070 2966 8108 3000
rect 8142 2966 8189 3000
rect 7989 2927 8189 2966
rect 7989 2893 8036 2927
rect 8070 2893 8108 2927
rect 8142 2893 8189 2927
rect 7989 2854 8189 2893
rect 7989 2820 8036 2854
rect 8070 2820 8108 2854
rect 8142 2820 8189 2854
rect 7989 2781 8189 2820
rect 7989 2747 8036 2781
rect 8070 2747 8108 2781
rect 8142 2747 8189 2781
rect 7989 2708 8189 2747
rect 7989 2674 8036 2708
rect 8070 2674 8108 2708
rect 8142 2674 8189 2708
rect 7989 2635 8189 2674
rect 7989 2601 8036 2635
rect 8070 2601 8108 2635
rect 8142 2601 8189 2635
rect 7989 2562 8189 2601
rect 7989 2528 8036 2562
rect 8070 2528 8108 2562
rect 8142 2528 8189 2562
rect 7989 2489 8189 2528
rect 7989 2455 8036 2489
rect 8070 2455 8108 2489
rect 8142 2455 8189 2489
rect 7989 2416 8189 2455
rect 7989 2382 8036 2416
rect 8070 2382 8108 2416
rect 8142 2382 8189 2416
rect 7989 2343 8189 2382
rect 7989 2309 8036 2343
rect 8070 2309 8108 2343
rect 8142 2309 8189 2343
rect 7989 2270 8189 2309
rect 7989 2236 8036 2270
rect 8070 2236 8108 2270
rect 8142 2236 8189 2270
rect 7989 2197 8189 2236
rect 7989 2163 8036 2197
rect 8070 2163 8108 2197
rect 8142 2163 8189 2197
rect 7989 2124 8189 2163
rect 7989 2090 8036 2124
rect 8070 2090 8108 2124
rect 8142 2090 8189 2124
rect 7989 2051 8189 2090
rect 7989 2017 8036 2051
rect 8070 2017 8108 2051
rect 8142 2017 8189 2051
rect 7989 1978 8189 2017
rect 7989 1944 8036 1978
rect 8070 1944 8108 1978
rect 8142 1944 8189 1978
rect 7989 1905 8189 1944
rect 7989 1871 8036 1905
rect 8070 1871 8108 1905
rect 8142 1871 8189 1905
rect 7989 1832 8189 1871
rect 7989 1798 8036 1832
rect 8070 1798 8108 1832
rect 8142 1798 8189 1832
rect 7989 1759 8189 1798
rect 7989 1725 8036 1759
rect 8070 1725 8108 1759
rect 8142 1725 8189 1759
rect 7989 1686 8189 1725
rect 7989 1652 8036 1686
rect 8070 1652 8108 1686
rect 8142 1652 8189 1686
rect 7989 1613 8189 1652
rect 7989 1579 8036 1613
rect 8070 1579 8108 1613
rect 8142 1579 8189 1613
rect 7989 1540 8189 1579
rect 7989 1506 8036 1540
rect 8070 1506 8108 1540
rect 8142 1506 8189 1540
rect 7989 1466 8189 1506
rect 7989 1432 8036 1466
rect 8070 1432 8108 1466
rect 8142 1432 8189 1466
rect 7989 1392 8189 1432
rect 7989 1358 8036 1392
rect 8070 1358 8108 1392
rect 8142 1358 8189 1392
rect 7989 1318 8189 1358
rect 7989 1284 8036 1318
rect 8070 1284 8108 1318
rect 8142 1284 8189 1318
rect 7989 1244 8189 1284
rect 7989 1210 8036 1244
rect 8070 1210 8108 1244
rect 8142 1210 8189 1244
rect 7989 1170 8189 1210
rect 7989 1136 8036 1170
rect 8070 1136 8108 1170
rect 8142 1136 8189 1170
rect 7989 1096 8189 1136
rect 7989 1062 8036 1096
rect 8070 1062 8108 1096
rect 8142 1062 8189 1096
rect 7989 1022 8189 1062
rect 7989 988 8036 1022
rect 8070 988 8108 1022
rect 8142 988 8189 1022
rect 7989 948 8189 988
rect 7989 914 8036 948
rect 8070 914 8108 948
rect 8142 914 8189 948
rect 7989 874 8189 914
rect 7989 840 8036 874
rect 8070 840 8108 874
rect 8142 840 8189 874
rect 7989 800 8189 840
rect 7989 766 8036 800
rect 8070 766 8108 800
rect 8142 766 8189 800
rect 7989 726 8189 766
rect 7989 692 8036 726
rect 8070 692 8108 726
rect 8142 692 8189 726
rect 7989 652 8189 692
rect 7989 618 8036 652
rect 8070 618 8108 652
rect 8142 618 8189 652
rect 7989 578 8189 618
rect 7989 544 8036 578
rect 8070 544 8108 578
rect 8142 544 8189 578
rect 7989 504 8189 544
rect 7989 470 8036 504
rect 8070 470 8108 504
rect 8142 470 8189 504
rect 7989 430 8189 470
rect 7989 396 8036 430
rect 8070 396 8108 430
rect 8142 396 8189 430
rect 7989 356 8189 396
rect 7989 322 8036 356
rect 8070 322 8108 356
rect 8142 322 8189 356
rect 7989 282 8189 322
rect 7989 248 8036 282
rect 8070 248 8108 282
rect 8142 248 8189 282
rect 7989 208 8189 248
rect 7989 174 8036 208
rect 8070 174 8108 208
rect 8142 174 8189 208
rect 7989 134 8189 174
rect 7989 100 8036 134
rect 8070 100 8108 134
rect 8142 100 8189 134
rect 7989 47 8189 100
tri 7989 42 7994 47 ne
rect 7994 42 8184 47
tri 8184 42 8189 47 nw
tri 8301 3053 8348 3100 se
rect 8348 3053 8654 3100
tri 8654 3053 8701 3100 sw
rect 8301 3000 8701 3053
rect 8301 2966 8448 3000
rect 8482 2966 8520 3000
rect 8554 2966 8701 3000
rect 8301 2927 8701 2966
rect 8301 2893 8448 2927
rect 8482 2893 8520 2927
rect 8554 2893 8701 2927
rect 8301 2854 8701 2893
rect 8301 2820 8448 2854
rect 8482 2820 8520 2854
rect 8554 2820 8701 2854
rect 8301 2781 8701 2820
rect 8301 2747 8448 2781
rect 8482 2747 8520 2781
rect 8554 2747 8701 2781
rect 8301 2708 8701 2747
rect 8301 2674 8448 2708
rect 8482 2674 8520 2708
rect 8554 2674 8701 2708
rect 8301 2635 8701 2674
rect 8301 2601 8448 2635
rect 8482 2601 8520 2635
rect 8554 2601 8701 2635
rect 8301 2562 8701 2601
rect 8301 2528 8448 2562
rect 8482 2528 8520 2562
rect 8554 2528 8701 2562
rect 8301 2489 8701 2528
rect 8301 2455 8448 2489
rect 8482 2455 8520 2489
rect 8554 2455 8701 2489
rect 8301 2416 8701 2455
rect 8301 2382 8448 2416
rect 8482 2382 8520 2416
rect 8554 2382 8701 2416
rect 8301 2343 8701 2382
rect 8301 2309 8448 2343
rect 8482 2309 8520 2343
rect 8554 2309 8701 2343
rect 8301 2270 8701 2309
rect 8301 2236 8448 2270
rect 8482 2236 8520 2270
rect 8554 2236 8701 2270
rect 8301 2197 8701 2236
rect 8301 2163 8448 2197
rect 8482 2163 8520 2197
rect 8554 2163 8701 2197
rect 8301 2124 8701 2163
rect 8301 2090 8448 2124
rect 8482 2090 8520 2124
rect 8554 2090 8701 2124
rect 8301 2051 8701 2090
rect 8301 2017 8448 2051
rect 8482 2017 8520 2051
rect 8554 2017 8701 2051
rect 8301 1978 8701 2017
rect 8301 1944 8448 1978
rect 8482 1944 8520 1978
rect 8554 1944 8701 1978
rect 8301 1905 8701 1944
rect 8301 1871 8448 1905
rect 8482 1871 8520 1905
rect 8554 1871 8701 1905
rect 8301 1832 8701 1871
rect 8301 1798 8448 1832
rect 8482 1798 8520 1832
rect 8554 1798 8701 1832
rect 8301 1759 8701 1798
rect 8301 1725 8448 1759
rect 8482 1725 8520 1759
rect 8554 1725 8701 1759
rect 8301 1686 8701 1725
rect 8301 1652 8448 1686
rect 8482 1652 8520 1686
rect 8554 1652 8701 1686
rect 8301 1613 8701 1652
rect 8301 1579 8448 1613
rect 8482 1579 8520 1613
rect 8554 1579 8701 1613
rect 8301 1540 8701 1579
rect 8301 1506 8448 1540
rect 8482 1506 8520 1540
rect 8554 1506 8701 1540
rect 8301 1466 8701 1506
rect 8301 1432 8448 1466
rect 8482 1432 8520 1466
rect 8554 1432 8701 1466
rect 8301 1392 8701 1432
rect 8301 1358 8448 1392
rect 8482 1358 8520 1392
rect 8554 1358 8701 1392
rect 8301 1318 8701 1358
rect 8301 1284 8448 1318
rect 8482 1284 8520 1318
rect 8554 1284 8701 1318
rect 8301 1244 8701 1284
rect 8301 1210 8448 1244
rect 8482 1210 8520 1244
rect 8554 1210 8701 1244
rect 8301 1170 8701 1210
rect 8301 1136 8448 1170
rect 8482 1136 8520 1170
rect 8554 1136 8701 1170
rect 8301 1096 8701 1136
rect 8301 1062 8448 1096
rect 8482 1062 8520 1096
rect 8554 1062 8701 1096
rect 8301 1022 8701 1062
rect 8301 988 8448 1022
rect 8482 988 8520 1022
rect 8554 988 8701 1022
rect 8301 948 8701 988
rect 8301 914 8448 948
rect 8482 914 8520 948
rect 8554 914 8701 948
rect 8301 874 8701 914
rect 8301 840 8448 874
rect 8482 840 8520 874
rect 8554 840 8701 874
rect 8301 800 8701 840
rect 8301 766 8448 800
rect 8482 766 8520 800
rect 8554 766 8701 800
rect 8301 726 8701 766
rect 8301 692 8448 726
rect 8482 692 8520 726
rect 8554 692 8701 726
rect 8301 652 8701 692
rect 8301 618 8448 652
rect 8482 618 8520 652
rect 8554 618 8701 652
rect 8301 578 8701 618
rect 8301 544 8448 578
rect 8482 544 8520 578
rect 8554 544 8701 578
rect 8301 504 8701 544
rect 8301 470 8448 504
rect 8482 470 8520 504
rect 8554 470 8701 504
rect 8301 430 8701 470
rect 8301 396 8448 430
rect 8482 396 8520 430
rect 8554 396 8701 430
rect 8301 356 8701 396
rect 8301 322 8448 356
rect 8482 322 8520 356
rect 8554 322 8701 356
rect 8301 282 8701 322
rect 8301 248 8448 282
rect 8482 248 8520 282
rect 8554 248 8701 282
rect 8301 208 8701 248
rect 8301 174 8448 208
rect 8482 174 8520 208
rect 8554 174 8701 208
rect 8301 134 8701 174
rect 8301 100 8448 134
rect 8482 100 8520 134
rect 8554 100 8701 134
rect 8301 47 8701 100
tri 8301 42 8306 47 ne
rect 8306 42 8696 47
tri 8696 42 8701 47 nw
tri 8813 3053 8860 3100 se
rect 8860 3053 8966 3100
tri 8966 3053 9013 3100 sw
rect 8813 3000 9013 3053
rect 8813 2966 8860 3000
rect 8894 2966 8932 3000
rect 8966 2966 9013 3000
rect 8813 2927 9013 2966
rect 8813 2893 8860 2927
rect 8894 2893 8932 2927
rect 8966 2893 9013 2927
rect 8813 2854 9013 2893
rect 8813 2820 8860 2854
rect 8894 2820 8932 2854
rect 8966 2820 9013 2854
rect 8813 2781 9013 2820
rect 8813 2747 8860 2781
rect 8894 2747 8932 2781
rect 8966 2747 9013 2781
rect 8813 2708 9013 2747
rect 8813 2674 8860 2708
rect 8894 2674 8932 2708
rect 8966 2674 9013 2708
rect 8813 2635 9013 2674
rect 8813 2601 8860 2635
rect 8894 2601 8932 2635
rect 8966 2601 9013 2635
rect 8813 2562 9013 2601
rect 8813 2528 8860 2562
rect 8894 2528 8932 2562
rect 8966 2528 9013 2562
rect 8813 2489 9013 2528
rect 8813 2455 8860 2489
rect 8894 2455 8932 2489
rect 8966 2455 9013 2489
rect 8813 2416 9013 2455
rect 8813 2382 8860 2416
rect 8894 2382 8932 2416
rect 8966 2382 9013 2416
rect 8813 2343 9013 2382
rect 8813 2309 8860 2343
rect 8894 2309 8932 2343
rect 8966 2309 9013 2343
rect 8813 2270 9013 2309
rect 8813 2236 8860 2270
rect 8894 2236 8932 2270
rect 8966 2236 9013 2270
rect 8813 2197 9013 2236
rect 8813 2163 8860 2197
rect 8894 2163 8932 2197
rect 8966 2163 9013 2197
rect 8813 2124 9013 2163
rect 8813 2090 8860 2124
rect 8894 2090 8932 2124
rect 8966 2090 9013 2124
rect 8813 2051 9013 2090
rect 8813 2017 8860 2051
rect 8894 2017 8932 2051
rect 8966 2017 9013 2051
rect 8813 1978 9013 2017
rect 8813 1944 8860 1978
rect 8894 1944 8932 1978
rect 8966 1944 9013 1978
rect 8813 1905 9013 1944
rect 8813 1871 8860 1905
rect 8894 1871 8932 1905
rect 8966 1871 9013 1905
rect 8813 1832 9013 1871
rect 8813 1798 8860 1832
rect 8894 1798 8932 1832
rect 8966 1798 9013 1832
rect 8813 1759 9013 1798
rect 8813 1725 8860 1759
rect 8894 1725 8932 1759
rect 8966 1725 9013 1759
rect 8813 1686 9013 1725
rect 8813 1652 8860 1686
rect 8894 1652 8932 1686
rect 8966 1652 9013 1686
rect 8813 1613 9013 1652
rect 8813 1579 8860 1613
rect 8894 1579 8932 1613
rect 8966 1579 9013 1613
rect 8813 1540 9013 1579
rect 8813 1506 8860 1540
rect 8894 1506 8932 1540
rect 8966 1506 9013 1540
rect 8813 1466 9013 1506
rect 8813 1432 8860 1466
rect 8894 1432 8932 1466
rect 8966 1432 9013 1466
rect 8813 1392 9013 1432
rect 8813 1358 8860 1392
rect 8894 1358 8932 1392
rect 8966 1358 9013 1392
rect 8813 1318 9013 1358
rect 8813 1284 8860 1318
rect 8894 1284 8932 1318
rect 8966 1284 9013 1318
rect 8813 1244 9013 1284
rect 8813 1210 8860 1244
rect 8894 1210 8932 1244
rect 8966 1210 9013 1244
rect 8813 1170 9013 1210
rect 8813 1136 8860 1170
rect 8894 1136 8932 1170
rect 8966 1136 9013 1170
rect 8813 1096 9013 1136
rect 8813 1062 8860 1096
rect 8894 1062 8932 1096
rect 8966 1062 9013 1096
rect 8813 1022 9013 1062
rect 8813 988 8860 1022
rect 8894 988 8932 1022
rect 8966 988 9013 1022
rect 8813 948 9013 988
rect 8813 914 8860 948
rect 8894 914 8932 948
rect 8966 914 9013 948
rect 8813 874 9013 914
rect 8813 840 8860 874
rect 8894 840 8932 874
rect 8966 840 9013 874
rect 8813 800 9013 840
rect 8813 766 8860 800
rect 8894 766 8932 800
rect 8966 766 9013 800
rect 8813 726 9013 766
rect 8813 692 8860 726
rect 8894 692 8932 726
rect 8966 692 9013 726
rect 8813 652 9013 692
rect 8813 618 8860 652
rect 8894 618 8932 652
rect 8966 618 9013 652
rect 8813 578 9013 618
rect 8813 544 8860 578
rect 8894 544 8932 578
rect 8966 544 9013 578
rect 8813 504 9013 544
rect 8813 470 8860 504
rect 8894 470 8932 504
rect 8966 470 9013 504
rect 8813 430 9013 470
rect 8813 396 8860 430
rect 8894 396 8932 430
rect 8966 396 9013 430
rect 8813 356 9013 396
rect 8813 322 8860 356
rect 8894 322 8932 356
rect 8966 322 9013 356
rect 8813 282 9013 322
rect 8813 248 8860 282
rect 8894 248 8932 282
rect 8966 248 9013 282
rect 8813 208 9013 248
rect 8813 174 8860 208
rect 8894 174 8932 208
rect 8966 174 9013 208
rect 8813 134 9013 174
rect 8813 100 8860 134
rect 8894 100 8932 134
rect 8966 100 9013 134
rect 8813 47 9013 100
tri 8813 42 8818 47 ne
rect 8818 42 9008 47
tri 9008 42 9013 47 nw
tri 9125 3053 9172 3100 se
rect 9172 3053 9478 3100
tri 9478 3053 9525 3100 sw
rect 9125 3000 9525 3053
rect 9125 2966 9272 3000
rect 9306 2966 9344 3000
rect 9378 2966 9525 3000
rect 9125 2927 9525 2966
rect 9125 2893 9272 2927
rect 9306 2893 9344 2927
rect 9378 2893 9525 2927
rect 9125 2854 9525 2893
rect 9125 2820 9272 2854
rect 9306 2820 9344 2854
rect 9378 2820 9525 2854
rect 9125 2781 9525 2820
rect 9125 2747 9272 2781
rect 9306 2747 9344 2781
rect 9378 2747 9525 2781
rect 9125 2708 9525 2747
rect 9125 2674 9272 2708
rect 9306 2674 9344 2708
rect 9378 2674 9525 2708
rect 9125 2635 9525 2674
rect 9125 2601 9272 2635
rect 9306 2601 9344 2635
rect 9378 2601 9525 2635
rect 9125 2562 9525 2601
rect 9125 2528 9272 2562
rect 9306 2528 9344 2562
rect 9378 2528 9525 2562
rect 9125 2489 9525 2528
rect 9125 2455 9272 2489
rect 9306 2455 9344 2489
rect 9378 2455 9525 2489
rect 9125 2416 9525 2455
rect 9125 2382 9272 2416
rect 9306 2382 9344 2416
rect 9378 2382 9525 2416
rect 9125 2343 9525 2382
rect 9125 2309 9272 2343
rect 9306 2309 9344 2343
rect 9378 2309 9525 2343
rect 9125 2270 9525 2309
rect 9125 2236 9272 2270
rect 9306 2236 9344 2270
rect 9378 2236 9525 2270
rect 9125 2197 9525 2236
rect 9125 2163 9272 2197
rect 9306 2163 9344 2197
rect 9378 2163 9525 2197
rect 9125 2124 9525 2163
rect 9125 2090 9272 2124
rect 9306 2090 9344 2124
rect 9378 2090 9525 2124
rect 9125 2051 9525 2090
rect 9125 2017 9272 2051
rect 9306 2017 9344 2051
rect 9378 2017 9525 2051
rect 9125 1978 9525 2017
rect 9125 1944 9272 1978
rect 9306 1944 9344 1978
rect 9378 1944 9525 1978
rect 9125 1905 9525 1944
rect 9125 1871 9272 1905
rect 9306 1871 9344 1905
rect 9378 1871 9525 1905
rect 9125 1832 9525 1871
rect 9125 1798 9272 1832
rect 9306 1798 9344 1832
rect 9378 1798 9525 1832
rect 9125 1759 9525 1798
rect 9125 1725 9272 1759
rect 9306 1725 9344 1759
rect 9378 1725 9525 1759
rect 9125 1686 9525 1725
rect 9125 1652 9272 1686
rect 9306 1652 9344 1686
rect 9378 1652 9525 1686
rect 9125 1613 9525 1652
rect 9125 1579 9272 1613
rect 9306 1579 9344 1613
rect 9378 1579 9525 1613
rect 9125 1540 9525 1579
rect 9125 1506 9272 1540
rect 9306 1506 9344 1540
rect 9378 1506 9525 1540
rect 9125 1466 9525 1506
rect 9125 1432 9272 1466
rect 9306 1432 9344 1466
rect 9378 1432 9525 1466
rect 9125 1392 9525 1432
rect 9125 1358 9272 1392
rect 9306 1358 9344 1392
rect 9378 1358 9525 1392
rect 9125 1318 9525 1358
rect 9125 1284 9272 1318
rect 9306 1284 9344 1318
rect 9378 1284 9525 1318
rect 9125 1244 9525 1284
rect 9125 1210 9272 1244
rect 9306 1210 9344 1244
rect 9378 1210 9525 1244
rect 9125 1170 9525 1210
rect 9125 1136 9272 1170
rect 9306 1136 9344 1170
rect 9378 1136 9525 1170
rect 9125 1096 9525 1136
rect 9125 1062 9272 1096
rect 9306 1062 9344 1096
rect 9378 1062 9525 1096
rect 9125 1022 9525 1062
rect 9125 988 9272 1022
rect 9306 988 9344 1022
rect 9378 988 9525 1022
rect 9125 948 9525 988
rect 9125 914 9272 948
rect 9306 914 9344 948
rect 9378 914 9525 948
rect 9125 874 9525 914
rect 9125 840 9272 874
rect 9306 840 9344 874
rect 9378 840 9525 874
rect 9125 800 9525 840
rect 9125 766 9272 800
rect 9306 766 9344 800
rect 9378 766 9525 800
rect 9125 726 9525 766
rect 9125 692 9272 726
rect 9306 692 9344 726
rect 9378 692 9525 726
rect 9125 652 9525 692
rect 9125 618 9272 652
rect 9306 618 9344 652
rect 9378 618 9525 652
rect 9125 578 9525 618
rect 9125 544 9272 578
rect 9306 544 9344 578
rect 9378 544 9525 578
rect 9125 504 9525 544
rect 9125 470 9272 504
rect 9306 470 9344 504
rect 9378 470 9525 504
rect 9125 430 9525 470
rect 9125 396 9272 430
rect 9306 396 9344 430
rect 9378 396 9525 430
rect 9125 356 9525 396
rect 9125 322 9272 356
rect 9306 322 9344 356
rect 9378 322 9525 356
rect 9125 282 9525 322
rect 9125 248 9272 282
rect 9306 248 9344 282
rect 9378 248 9525 282
rect 9125 208 9525 248
rect 9125 174 9272 208
rect 9306 174 9344 208
rect 9378 174 9525 208
rect 9125 134 9525 174
rect 9125 100 9272 134
rect 9306 100 9344 134
rect 9378 100 9525 134
rect 9125 47 9525 100
tri 9125 42 9130 47 ne
rect 9130 42 9520 47
tri 9520 42 9525 47 nw
tri 9637 3053 9684 3100 se
rect 9684 3053 9790 3100
tri 9790 3053 9837 3100 sw
rect 9637 3000 9837 3053
rect 9637 2966 9684 3000
rect 9718 2966 9756 3000
rect 9790 2966 9837 3000
rect 9637 2927 9837 2966
rect 9637 2893 9684 2927
rect 9718 2893 9756 2927
rect 9790 2893 9837 2927
rect 9637 2854 9837 2893
rect 9637 2820 9684 2854
rect 9718 2820 9756 2854
rect 9790 2820 9837 2854
rect 9637 2781 9837 2820
rect 9637 2747 9684 2781
rect 9718 2747 9756 2781
rect 9790 2747 9837 2781
rect 9637 2708 9837 2747
rect 9637 2674 9684 2708
rect 9718 2674 9756 2708
rect 9790 2674 9837 2708
rect 9637 2635 9837 2674
rect 9637 2601 9684 2635
rect 9718 2601 9756 2635
rect 9790 2601 9837 2635
rect 9637 2562 9837 2601
rect 9637 2528 9684 2562
rect 9718 2528 9756 2562
rect 9790 2528 9837 2562
rect 9637 2489 9837 2528
rect 9637 2455 9684 2489
rect 9718 2455 9756 2489
rect 9790 2455 9837 2489
rect 9637 2416 9837 2455
rect 9637 2382 9684 2416
rect 9718 2382 9756 2416
rect 9790 2382 9837 2416
rect 9637 2343 9837 2382
rect 9637 2309 9684 2343
rect 9718 2309 9756 2343
rect 9790 2309 9837 2343
rect 9637 2270 9837 2309
rect 9637 2236 9684 2270
rect 9718 2236 9756 2270
rect 9790 2236 9837 2270
rect 9637 2197 9837 2236
rect 9637 2163 9684 2197
rect 9718 2163 9756 2197
rect 9790 2163 9837 2197
rect 9637 2124 9837 2163
rect 9637 2090 9684 2124
rect 9718 2090 9756 2124
rect 9790 2090 9837 2124
rect 9637 2051 9837 2090
rect 9637 2017 9684 2051
rect 9718 2017 9756 2051
rect 9790 2017 9837 2051
rect 9637 1978 9837 2017
rect 9637 1944 9684 1978
rect 9718 1944 9756 1978
rect 9790 1944 9837 1978
rect 9637 1905 9837 1944
rect 9637 1871 9684 1905
rect 9718 1871 9756 1905
rect 9790 1871 9837 1905
rect 9637 1832 9837 1871
rect 9637 1798 9684 1832
rect 9718 1798 9756 1832
rect 9790 1798 9837 1832
rect 9637 1759 9837 1798
rect 9637 1725 9684 1759
rect 9718 1725 9756 1759
rect 9790 1725 9837 1759
rect 9637 1686 9837 1725
rect 9637 1652 9684 1686
rect 9718 1652 9756 1686
rect 9790 1652 9837 1686
rect 9637 1613 9837 1652
rect 9637 1579 9684 1613
rect 9718 1579 9756 1613
rect 9790 1579 9837 1613
rect 9637 1540 9837 1579
rect 9637 1506 9684 1540
rect 9718 1506 9756 1540
rect 9790 1506 9837 1540
rect 9637 1466 9837 1506
rect 9637 1432 9684 1466
rect 9718 1432 9756 1466
rect 9790 1432 9837 1466
rect 9637 1392 9837 1432
rect 9637 1358 9684 1392
rect 9718 1358 9756 1392
rect 9790 1358 9837 1392
rect 9637 1318 9837 1358
rect 9637 1284 9684 1318
rect 9718 1284 9756 1318
rect 9790 1284 9837 1318
rect 9637 1244 9837 1284
rect 9637 1210 9684 1244
rect 9718 1210 9756 1244
rect 9790 1210 9837 1244
rect 9637 1170 9837 1210
rect 9637 1136 9684 1170
rect 9718 1136 9756 1170
rect 9790 1136 9837 1170
rect 9637 1096 9837 1136
rect 9637 1062 9684 1096
rect 9718 1062 9756 1096
rect 9790 1062 9837 1096
rect 9637 1022 9837 1062
rect 9637 988 9684 1022
rect 9718 988 9756 1022
rect 9790 988 9837 1022
rect 9637 948 9837 988
rect 9637 914 9684 948
rect 9718 914 9756 948
rect 9790 914 9837 948
rect 9637 874 9837 914
rect 9637 840 9684 874
rect 9718 840 9756 874
rect 9790 840 9837 874
rect 9637 800 9837 840
rect 9637 766 9684 800
rect 9718 766 9756 800
rect 9790 766 9837 800
rect 9637 726 9837 766
rect 9637 692 9684 726
rect 9718 692 9756 726
rect 9790 692 9837 726
rect 9637 652 9837 692
rect 9637 618 9684 652
rect 9718 618 9756 652
rect 9790 618 9837 652
rect 9637 578 9837 618
rect 9637 544 9684 578
rect 9718 544 9756 578
rect 9790 544 9837 578
rect 9637 504 9837 544
rect 9637 470 9684 504
rect 9718 470 9756 504
rect 9790 470 9837 504
rect 9637 430 9837 470
rect 9637 396 9684 430
rect 9718 396 9756 430
rect 9790 396 9837 430
rect 9637 356 9837 396
rect 9637 322 9684 356
rect 9718 322 9756 356
rect 9790 322 9837 356
rect 9637 282 9837 322
rect 9637 248 9684 282
rect 9718 248 9756 282
rect 9790 248 9837 282
rect 9637 208 9837 248
rect 9637 174 9684 208
rect 9718 174 9756 208
rect 9790 174 9837 208
rect 9637 134 9837 174
rect 9637 100 9684 134
rect 9718 100 9756 134
rect 9790 100 9837 134
rect 9637 47 9837 100
tri 9637 42 9642 47 ne
rect 9642 42 9832 47
tri 9832 42 9837 47 nw
tri 9949 3053 9996 3100 se
rect 9996 3053 10302 3100
tri 10302 3053 10349 3100 sw
rect 9949 3000 10349 3053
rect 9949 2966 10096 3000
rect 10130 2966 10168 3000
rect 10202 2966 10349 3000
rect 9949 2927 10349 2966
rect 9949 2893 10096 2927
rect 10130 2893 10168 2927
rect 10202 2893 10349 2927
rect 9949 2854 10349 2893
rect 9949 2820 10096 2854
rect 10130 2820 10168 2854
rect 10202 2820 10349 2854
rect 9949 2781 10349 2820
rect 9949 2747 10096 2781
rect 10130 2747 10168 2781
rect 10202 2747 10349 2781
rect 9949 2708 10349 2747
rect 9949 2674 10096 2708
rect 10130 2674 10168 2708
rect 10202 2674 10349 2708
rect 9949 2635 10349 2674
rect 9949 2601 10096 2635
rect 10130 2601 10168 2635
rect 10202 2601 10349 2635
rect 9949 2562 10349 2601
rect 9949 2528 10096 2562
rect 10130 2528 10168 2562
rect 10202 2528 10349 2562
rect 9949 2489 10349 2528
rect 9949 2455 10096 2489
rect 10130 2455 10168 2489
rect 10202 2455 10349 2489
rect 9949 2416 10349 2455
rect 9949 2382 10096 2416
rect 10130 2382 10168 2416
rect 10202 2382 10349 2416
rect 9949 2343 10349 2382
rect 9949 2309 10096 2343
rect 10130 2309 10168 2343
rect 10202 2309 10349 2343
rect 9949 2270 10349 2309
rect 9949 2236 10096 2270
rect 10130 2236 10168 2270
rect 10202 2236 10349 2270
rect 9949 2197 10349 2236
rect 9949 2163 10096 2197
rect 10130 2163 10168 2197
rect 10202 2163 10349 2197
rect 9949 2124 10349 2163
rect 9949 2090 10096 2124
rect 10130 2090 10168 2124
rect 10202 2090 10349 2124
rect 9949 2051 10349 2090
rect 9949 2017 10096 2051
rect 10130 2017 10168 2051
rect 10202 2017 10349 2051
rect 9949 1978 10349 2017
rect 9949 1944 10096 1978
rect 10130 1944 10168 1978
rect 10202 1944 10349 1978
rect 9949 1905 10349 1944
rect 9949 1871 10096 1905
rect 10130 1871 10168 1905
rect 10202 1871 10349 1905
rect 9949 1832 10349 1871
rect 9949 1798 10096 1832
rect 10130 1798 10168 1832
rect 10202 1798 10349 1832
rect 9949 1759 10349 1798
rect 9949 1725 10096 1759
rect 10130 1725 10168 1759
rect 10202 1725 10349 1759
rect 9949 1686 10349 1725
rect 9949 1652 10096 1686
rect 10130 1652 10168 1686
rect 10202 1652 10349 1686
rect 9949 1613 10349 1652
rect 9949 1579 10096 1613
rect 10130 1579 10168 1613
rect 10202 1579 10349 1613
rect 9949 1540 10349 1579
rect 9949 1506 10096 1540
rect 10130 1506 10168 1540
rect 10202 1506 10349 1540
rect 9949 1466 10349 1506
rect 9949 1432 10096 1466
rect 10130 1432 10168 1466
rect 10202 1432 10349 1466
rect 9949 1392 10349 1432
rect 9949 1358 10096 1392
rect 10130 1358 10168 1392
rect 10202 1358 10349 1392
rect 9949 1318 10349 1358
rect 9949 1284 10096 1318
rect 10130 1284 10168 1318
rect 10202 1284 10349 1318
rect 9949 1244 10349 1284
rect 9949 1210 10096 1244
rect 10130 1210 10168 1244
rect 10202 1210 10349 1244
rect 9949 1170 10349 1210
rect 9949 1136 10096 1170
rect 10130 1136 10168 1170
rect 10202 1136 10349 1170
rect 9949 1096 10349 1136
rect 9949 1062 10096 1096
rect 10130 1062 10168 1096
rect 10202 1062 10349 1096
rect 9949 1022 10349 1062
rect 9949 988 10096 1022
rect 10130 988 10168 1022
rect 10202 988 10349 1022
rect 9949 948 10349 988
rect 9949 914 10096 948
rect 10130 914 10168 948
rect 10202 914 10349 948
rect 9949 874 10349 914
rect 9949 840 10096 874
rect 10130 840 10168 874
rect 10202 840 10349 874
rect 9949 800 10349 840
rect 9949 766 10096 800
rect 10130 766 10168 800
rect 10202 766 10349 800
rect 9949 726 10349 766
rect 9949 692 10096 726
rect 10130 692 10168 726
rect 10202 692 10349 726
rect 9949 652 10349 692
rect 9949 618 10096 652
rect 10130 618 10168 652
rect 10202 618 10349 652
rect 9949 578 10349 618
rect 9949 544 10096 578
rect 10130 544 10168 578
rect 10202 544 10349 578
rect 9949 504 10349 544
rect 9949 470 10096 504
rect 10130 470 10168 504
rect 10202 470 10349 504
rect 9949 430 10349 470
rect 9949 396 10096 430
rect 10130 396 10168 430
rect 10202 396 10349 430
rect 9949 356 10349 396
rect 9949 322 10096 356
rect 10130 322 10168 356
rect 10202 322 10349 356
rect 9949 282 10349 322
rect 9949 248 10096 282
rect 10130 248 10168 282
rect 10202 248 10349 282
rect 9949 208 10349 248
rect 9949 174 10096 208
rect 10130 174 10168 208
rect 10202 174 10349 208
rect 9949 134 10349 174
rect 9949 100 10096 134
rect 10130 100 10168 134
rect 10202 100 10349 134
rect 9949 47 10349 100
tri 9949 42 9954 47 ne
rect 9954 42 10344 47
tri 10344 42 10349 47 nw
tri 10461 3053 10508 3100 se
rect 10508 3053 10614 3100
tri 10614 3053 10661 3100 sw
rect 10461 3000 10661 3053
rect 10461 2966 10508 3000
rect 10542 2966 10580 3000
rect 10614 2966 10661 3000
rect 10461 2927 10661 2966
rect 10461 2893 10508 2927
rect 10542 2893 10580 2927
rect 10614 2893 10661 2927
rect 10461 2854 10661 2893
rect 10461 2820 10508 2854
rect 10542 2820 10580 2854
rect 10614 2820 10661 2854
rect 10461 2781 10661 2820
rect 10461 2747 10508 2781
rect 10542 2747 10580 2781
rect 10614 2747 10661 2781
rect 10461 2708 10661 2747
rect 10461 2674 10508 2708
rect 10542 2674 10580 2708
rect 10614 2674 10661 2708
rect 10461 2635 10661 2674
rect 10461 2601 10508 2635
rect 10542 2601 10580 2635
rect 10614 2601 10661 2635
rect 10461 2562 10661 2601
rect 10461 2528 10508 2562
rect 10542 2528 10580 2562
rect 10614 2528 10661 2562
rect 10461 2489 10661 2528
rect 10461 2455 10508 2489
rect 10542 2455 10580 2489
rect 10614 2455 10661 2489
rect 10461 2416 10661 2455
rect 10461 2382 10508 2416
rect 10542 2382 10580 2416
rect 10614 2382 10661 2416
rect 10461 2343 10661 2382
rect 10461 2309 10508 2343
rect 10542 2309 10580 2343
rect 10614 2309 10661 2343
rect 10461 2270 10661 2309
rect 10461 2236 10508 2270
rect 10542 2236 10580 2270
rect 10614 2236 10661 2270
rect 10461 2197 10661 2236
rect 10461 2163 10508 2197
rect 10542 2163 10580 2197
rect 10614 2163 10661 2197
rect 10461 2124 10661 2163
rect 10461 2090 10508 2124
rect 10542 2090 10580 2124
rect 10614 2090 10661 2124
rect 10461 2051 10661 2090
rect 10461 2017 10508 2051
rect 10542 2017 10580 2051
rect 10614 2017 10661 2051
rect 10461 1978 10661 2017
rect 10461 1944 10508 1978
rect 10542 1944 10580 1978
rect 10614 1944 10661 1978
rect 10461 1905 10661 1944
rect 10461 1871 10508 1905
rect 10542 1871 10580 1905
rect 10614 1871 10661 1905
rect 10461 1832 10661 1871
rect 10461 1798 10508 1832
rect 10542 1798 10580 1832
rect 10614 1798 10661 1832
rect 10461 1759 10661 1798
rect 10461 1725 10508 1759
rect 10542 1725 10580 1759
rect 10614 1725 10661 1759
rect 10461 1686 10661 1725
rect 10461 1652 10508 1686
rect 10542 1652 10580 1686
rect 10614 1652 10661 1686
rect 10461 1613 10661 1652
rect 10461 1579 10508 1613
rect 10542 1579 10580 1613
rect 10614 1579 10661 1613
rect 10461 1540 10661 1579
rect 10461 1506 10508 1540
rect 10542 1506 10580 1540
rect 10614 1506 10661 1540
rect 10461 1466 10661 1506
rect 10461 1432 10508 1466
rect 10542 1432 10580 1466
rect 10614 1432 10661 1466
rect 10461 1392 10661 1432
rect 10461 1358 10508 1392
rect 10542 1358 10580 1392
rect 10614 1358 10661 1392
rect 10461 1318 10661 1358
rect 10461 1284 10508 1318
rect 10542 1284 10580 1318
rect 10614 1284 10661 1318
rect 10461 1244 10661 1284
rect 10461 1210 10508 1244
rect 10542 1210 10580 1244
rect 10614 1210 10661 1244
rect 10461 1170 10661 1210
rect 10461 1136 10508 1170
rect 10542 1136 10580 1170
rect 10614 1136 10661 1170
rect 10461 1096 10661 1136
rect 10461 1062 10508 1096
rect 10542 1062 10580 1096
rect 10614 1062 10661 1096
rect 10461 1022 10661 1062
rect 10461 988 10508 1022
rect 10542 988 10580 1022
rect 10614 988 10661 1022
rect 10461 948 10661 988
rect 10461 914 10508 948
rect 10542 914 10580 948
rect 10614 914 10661 948
rect 10461 874 10661 914
rect 10461 840 10508 874
rect 10542 840 10580 874
rect 10614 840 10661 874
rect 10461 800 10661 840
rect 10461 766 10508 800
rect 10542 766 10580 800
rect 10614 766 10661 800
rect 10461 726 10661 766
rect 10461 692 10508 726
rect 10542 692 10580 726
rect 10614 692 10661 726
rect 10461 652 10661 692
rect 10461 618 10508 652
rect 10542 618 10580 652
rect 10614 618 10661 652
rect 10461 578 10661 618
rect 10461 544 10508 578
rect 10542 544 10580 578
rect 10614 544 10661 578
rect 10461 504 10661 544
rect 10461 470 10508 504
rect 10542 470 10580 504
rect 10614 470 10661 504
rect 10461 430 10661 470
rect 10461 396 10508 430
rect 10542 396 10580 430
rect 10614 396 10661 430
rect 10461 356 10661 396
rect 10461 322 10508 356
rect 10542 322 10580 356
rect 10614 322 10661 356
rect 10461 282 10661 322
rect 10461 248 10508 282
rect 10542 248 10580 282
rect 10614 248 10661 282
rect 10461 208 10661 248
rect 10461 174 10508 208
rect 10542 174 10580 208
rect 10614 174 10661 208
rect 10461 134 10661 174
rect 10461 100 10508 134
rect 10542 100 10580 134
rect 10614 100 10661 134
rect 10461 47 10661 100
tri 10461 42 10466 47 ne
rect 10466 42 10656 47
tri 10656 42 10661 47 nw
tri 10773 3053 10820 3100 se
rect 10820 3053 11126 3100
tri 11126 3053 11173 3100 sw
rect 10773 3000 11173 3053
rect 10773 2966 10920 3000
rect 10954 2966 10992 3000
rect 11026 2966 11173 3000
rect 10773 2927 11173 2966
rect 10773 2893 10920 2927
rect 10954 2893 10992 2927
rect 11026 2893 11173 2927
rect 10773 2854 11173 2893
rect 10773 2820 10920 2854
rect 10954 2820 10992 2854
rect 11026 2820 11173 2854
rect 10773 2781 11173 2820
rect 10773 2747 10920 2781
rect 10954 2747 10992 2781
rect 11026 2747 11173 2781
rect 10773 2708 11173 2747
rect 10773 2674 10920 2708
rect 10954 2674 10992 2708
rect 11026 2674 11173 2708
rect 10773 2635 11173 2674
rect 10773 2601 10920 2635
rect 10954 2601 10992 2635
rect 11026 2601 11173 2635
rect 10773 2562 11173 2601
rect 10773 2528 10920 2562
rect 10954 2528 10992 2562
rect 11026 2528 11173 2562
rect 10773 2489 11173 2528
rect 10773 2455 10920 2489
rect 10954 2455 10992 2489
rect 11026 2455 11173 2489
rect 10773 2416 11173 2455
rect 10773 2382 10920 2416
rect 10954 2382 10992 2416
rect 11026 2382 11173 2416
rect 10773 2343 11173 2382
rect 10773 2309 10920 2343
rect 10954 2309 10992 2343
rect 11026 2309 11173 2343
rect 10773 2270 11173 2309
rect 10773 2236 10920 2270
rect 10954 2236 10992 2270
rect 11026 2236 11173 2270
rect 10773 2197 11173 2236
rect 10773 2163 10920 2197
rect 10954 2163 10992 2197
rect 11026 2163 11173 2197
rect 10773 2124 11173 2163
rect 10773 2090 10920 2124
rect 10954 2090 10992 2124
rect 11026 2090 11173 2124
rect 10773 2051 11173 2090
rect 10773 2017 10920 2051
rect 10954 2017 10992 2051
rect 11026 2017 11173 2051
rect 10773 1978 11173 2017
rect 10773 1944 10920 1978
rect 10954 1944 10992 1978
rect 11026 1944 11173 1978
rect 10773 1905 11173 1944
rect 10773 1871 10920 1905
rect 10954 1871 10992 1905
rect 11026 1871 11173 1905
rect 10773 1832 11173 1871
rect 10773 1798 10920 1832
rect 10954 1798 10992 1832
rect 11026 1798 11173 1832
rect 10773 1759 11173 1798
rect 10773 1725 10920 1759
rect 10954 1725 10992 1759
rect 11026 1725 11173 1759
rect 10773 1686 11173 1725
rect 10773 1652 10920 1686
rect 10954 1652 10992 1686
rect 11026 1652 11173 1686
rect 10773 1613 11173 1652
rect 10773 1579 10920 1613
rect 10954 1579 10992 1613
rect 11026 1579 11173 1613
rect 10773 1540 11173 1579
rect 10773 1506 10920 1540
rect 10954 1506 10992 1540
rect 11026 1506 11173 1540
rect 10773 1466 11173 1506
rect 10773 1432 10920 1466
rect 10954 1432 10992 1466
rect 11026 1432 11173 1466
rect 10773 1392 11173 1432
rect 10773 1358 10920 1392
rect 10954 1358 10992 1392
rect 11026 1358 11173 1392
rect 10773 1318 11173 1358
rect 10773 1284 10920 1318
rect 10954 1284 10992 1318
rect 11026 1284 11173 1318
rect 10773 1244 11173 1284
rect 10773 1210 10920 1244
rect 10954 1210 10992 1244
rect 11026 1210 11173 1244
rect 10773 1170 11173 1210
rect 10773 1136 10920 1170
rect 10954 1136 10992 1170
rect 11026 1136 11173 1170
rect 10773 1096 11173 1136
rect 10773 1062 10920 1096
rect 10954 1062 10992 1096
rect 11026 1062 11173 1096
rect 10773 1022 11173 1062
rect 10773 988 10920 1022
rect 10954 988 10992 1022
rect 11026 988 11173 1022
rect 10773 948 11173 988
rect 10773 914 10920 948
rect 10954 914 10992 948
rect 11026 914 11173 948
rect 10773 874 11173 914
rect 10773 840 10920 874
rect 10954 840 10992 874
rect 11026 840 11173 874
rect 10773 800 11173 840
rect 10773 766 10920 800
rect 10954 766 10992 800
rect 11026 766 11173 800
rect 10773 726 11173 766
rect 10773 692 10920 726
rect 10954 692 10992 726
rect 11026 692 11173 726
rect 10773 652 11173 692
rect 10773 618 10920 652
rect 10954 618 10992 652
rect 11026 618 11173 652
rect 10773 578 11173 618
rect 10773 544 10920 578
rect 10954 544 10992 578
rect 11026 544 11173 578
rect 10773 504 11173 544
rect 10773 470 10920 504
rect 10954 470 10992 504
rect 11026 470 11173 504
rect 10773 430 11173 470
rect 10773 396 10920 430
rect 10954 396 10992 430
rect 11026 396 11173 430
rect 10773 356 11173 396
rect 10773 322 10920 356
rect 10954 322 10992 356
rect 11026 322 11173 356
rect 10773 282 11173 322
rect 10773 248 10920 282
rect 10954 248 10992 282
rect 11026 248 11173 282
rect 10773 208 11173 248
rect 10773 174 10920 208
rect 10954 174 10992 208
rect 11026 174 11173 208
rect 10773 134 11173 174
rect 10773 100 10920 134
rect 10954 100 10992 134
rect 11026 100 11173 134
rect 10773 47 11173 100
tri 10773 42 10778 47 ne
rect 10778 42 11168 47
tri 11168 42 11173 47 nw
tri 11285 3053 11332 3100 se
rect 11332 3053 11438 3100
tri 11438 3053 11485 3100 sw
rect 11285 3000 11485 3053
rect 11285 2966 11332 3000
rect 11366 2966 11404 3000
rect 11438 2966 11485 3000
rect 11285 2927 11485 2966
rect 11285 2893 11332 2927
rect 11366 2893 11404 2927
rect 11438 2893 11485 2927
rect 11285 2854 11485 2893
rect 11285 2820 11332 2854
rect 11366 2820 11404 2854
rect 11438 2820 11485 2854
rect 11285 2781 11485 2820
rect 11285 2747 11332 2781
rect 11366 2747 11404 2781
rect 11438 2747 11485 2781
rect 11285 2708 11485 2747
rect 11285 2674 11332 2708
rect 11366 2674 11404 2708
rect 11438 2674 11485 2708
rect 11285 2635 11485 2674
rect 11285 2601 11332 2635
rect 11366 2601 11404 2635
rect 11438 2601 11485 2635
rect 11285 2562 11485 2601
rect 11285 2528 11332 2562
rect 11366 2528 11404 2562
rect 11438 2528 11485 2562
rect 11285 2489 11485 2528
rect 11285 2455 11332 2489
rect 11366 2455 11404 2489
rect 11438 2455 11485 2489
rect 11285 2416 11485 2455
rect 11285 2382 11332 2416
rect 11366 2382 11404 2416
rect 11438 2382 11485 2416
rect 11285 2343 11485 2382
rect 11285 2309 11332 2343
rect 11366 2309 11404 2343
rect 11438 2309 11485 2343
rect 11285 2270 11485 2309
rect 11285 2236 11332 2270
rect 11366 2236 11404 2270
rect 11438 2236 11485 2270
rect 11285 2197 11485 2236
rect 11285 2163 11332 2197
rect 11366 2163 11404 2197
rect 11438 2163 11485 2197
rect 11285 2124 11485 2163
rect 11285 2090 11332 2124
rect 11366 2090 11404 2124
rect 11438 2090 11485 2124
rect 11285 2051 11485 2090
rect 11285 2017 11332 2051
rect 11366 2017 11404 2051
rect 11438 2017 11485 2051
rect 11285 1978 11485 2017
rect 11285 1944 11332 1978
rect 11366 1944 11404 1978
rect 11438 1944 11485 1978
rect 11285 1905 11485 1944
rect 11285 1871 11332 1905
rect 11366 1871 11404 1905
rect 11438 1871 11485 1905
rect 11285 1832 11485 1871
rect 11285 1798 11332 1832
rect 11366 1798 11404 1832
rect 11438 1798 11485 1832
rect 11285 1759 11485 1798
rect 11285 1725 11332 1759
rect 11366 1725 11404 1759
rect 11438 1725 11485 1759
rect 11285 1686 11485 1725
rect 11285 1652 11332 1686
rect 11366 1652 11404 1686
rect 11438 1652 11485 1686
rect 11285 1613 11485 1652
rect 11285 1579 11332 1613
rect 11366 1579 11404 1613
rect 11438 1579 11485 1613
rect 11285 1540 11485 1579
rect 11285 1506 11332 1540
rect 11366 1506 11404 1540
rect 11438 1506 11485 1540
rect 11285 1466 11485 1506
rect 11285 1432 11332 1466
rect 11366 1432 11404 1466
rect 11438 1432 11485 1466
rect 11285 1392 11485 1432
rect 11285 1358 11332 1392
rect 11366 1358 11404 1392
rect 11438 1358 11485 1392
rect 11285 1318 11485 1358
rect 11285 1284 11332 1318
rect 11366 1284 11404 1318
rect 11438 1284 11485 1318
rect 11285 1244 11485 1284
rect 11285 1210 11332 1244
rect 11366 1210 11404 1244
rect 11438 1210 11485 1244
rect 11285 1170 11485 1210
rect 11285 1136 11332 1170
rect 11366 1136 11404 1170
rect 11438 1136 11485 1170
rect 11285 1096 11485 1136
rect 11285 1062 11332 1096
rect 11366 1062 11404 1096
rect 11438 1062 11485 1096
rect 11285 1022 11485 1062
rect 11285 988 11332 1022
rect 11366 988 11404 1022
rect 11438 988 11485 1022
rect 11285 948 11485 988
rect 11285 914 11332 948
rect 11366 914 11404 948
rect 11438 914 11485 948
rect 11285 874 11485 914
rect 11285 840 11332 874
rect 11366 840 11404 874
rect 11438 840 11485 874
rect 11285 800 11485 840
rect 11285 766 11332 800
rect 11366 766 11404 800
rect 11438 766 11485 800
rect 11285 726 11485 766
rect 11285 692 11332 726
rect 11366 692 11404 726
rect 11438 692 11485 726
rect 11285 652 11485 692
rect 11285 618 11332 652
rect 11366 618 11404 652
rect 11438 618 11485 652
rect 11285 578 11485 618
rect 11285 544 11332 578
rect 11366 544 11404 578
rect 11438 544 11485 578
rect 11285 504 11485 544
rect 11285 470 11332 504
rect 11366 470 11404 504
rect 11438 470 11485 504
rect 11285 430 11485 470
rect 11285 396 11332 430
rect 11366 396 11404 430
rect 11438 396 11485 430
rect 11285 356 11485 396
rect 11285 322 11332 356
rect 11366 322 11404 356
rect 11438 322 11485 356
rect 11285 282 11485 322
rect 11285 248 11332 282
rect 11366 248 11404 282
rect 11438 248 11485 282
rect 11285 208 11485 248
rect 11285 174 11332 208
rect 11366 174 11404 208
rect 11438 174 11485 208
rect 11285 134 11485 174
rect 11285 100 11332 134
rect 11366 100 11404 134
rect 11438 100 11485 134
rect 11285 47 11485 100
tri 11285 42 11290 47 ne
rect 11290 42 11480 47
tri 11480 42 11485 47 nw
tri 11597 3053 11644 3100 se
rect 11644 3053 11950 3100
tri 11950 3053 11997 3100 sw
rect 11597 3000 11997 3053
rect 11597 2966 11744 3000
rect 11778 2966 11816 3000
rect 11850 2966 11997 3000
rect 11597 2927 11997 2966
rect 11597 2893 11744 2927
rect 11778 2893 11816 2927
rect 11850 2893 11997 2927
rect 11597 2854 11997 2893
rect 11597 2820 11744 2854
rect 11778 2820 11816 2854
rect 11850 2820 11997 2854
rect 11597 2781 11997 2820
rect 11597 2747 11744 2781
rect 11778 2747 11816 2781
rect 11850 2747 11997 2781
rect 11597 2708 11997 2747
rect 11597 2674 11744 2708
rect 11778 2674 11816 2708
rect 11850 2674 11997 2708
rect 11597 2635 11997 2674
rect 11597 2601 11744 2635
rect 11778 2601 11816 2635
rect 11850 2601 11997 2635
rect 11597 2562 11997 2601
rect 11597 2528 11744 2562
rect 11778 2528 11816 2562
rect 11850 2528 11997 2562
rect 11597 2489 11997 2528
rect 11597 2455 11744 2489
rect 11778 2455 11816 2489
rect 11850 2455 11997 2489
rect 11597 2416 11997 2455
rect 11597 2382 11744 2416
rect 11778 2382 11816 2416
rect 11850 2382 11997 2416
rect 11597 2343 11997 2382
rect 11597 2309 11744 2343
rect 11778 2309 11816 2343
rect 11850 2309 11997 2343
rect 11597 2270 11997 2309
rect 11597 2236 11744 2270
rect 11778 2236 11816 2270
rect 11850 2236 11997 2270
rect 11597 2197 11997 2236
rect 11597 2163 11744 2197
rect 11778 2163 11816 2197
rect 11850 2163 11997 2197
rect 11597 2124 11997 2163
rect 11597 2090 11744 2124
rect 11778 2090 11816 2124
rect 11850 2090 11997 2124
rect 11597 2051 11997 2090
rect 11597 2017 11744 2051
rect 11778 2017 11816 2051
rect 11850 2017 11997 2051
rect 11597 1978 11997 2017
rect 11597 1944 11744 1978
rect 11778 1944 11816 1978
rect 11850 1944 11997 1978
rect 11597 1905 11997 1944
rect 11597 1871 11744 1905
rect 11778 1871 11816 1905
rect 11850 1871 11997 1905
rect 11597 1832 11997 1871
rect 11597 1798 11744 1832
rect 11778 1798 11816 1832
rect 11850 1798 11997 1832
rect 11597 1759 11997 1798
rect 11597 1725 11744 1759
rect 11778 1725 11816 1759
rect 11850 1725 11997 1759
rect 11597 1686 11997 1725
rect 11597 1652 11744 1686
rect 11778 1652 11816 1686
rect 11850 1652 11997 1686
rect 11597 1613 11997 1652
rect 11597 1579 11744 1613
rect 11778 1579 11816 1613
rect 11850 1579 11997 1613
rect 11597 1540 11997 1579
rect 11597 1506 11744 1540
rect 11778 1506 11816 1540
rect 11850 1506 11997 1540
rect 11597 1466 11997 1506
rect 11597 1432 11744 1466
rect 11778 1432 11816 1466
rect 11850 1432 11997 1466
rect 11597 1392 11997 1432
rect 11597 1358 11744 1392
rect 11778 1358 11816 1392
rect 11850 1358 11997 1392
rect 11597 1318 11997 1358
rect 11597 1284 11744 1318
rect 11778 1284 11816 1318
rect 11850 1284 11997 1318
rect 11597 1244 11997 1284
rect 11597 1210 11744 1244
rect 11778 1210 11816 1244
rect 11850 1210 11997 1244
rect 11597 1170 11997 1210
rect 11597 1136 11744 1170
rect 11778 1136 11816 1170
rect 11850 1136 11997 1170
rect 11597 1096 11997 1136
rect 11597 1062 11744 1096
rect 11778 1062 11816 1096
rect 11850 1062 11997 1096
rect 11597 1022 11997 1062
rect 11597 988 11744 1022
rect 11778 988 11816 1022
rect 11850 988 11997 1022
rect 11597 948 11997 988
rect 11597 914 11744 948
rect 11778 914 11816 948
rect 11850 914 11997 948
rect 11597 874 11997 914
rect 11597 840 11744 874
rect 11778 840 11816 874
rect 11850 840 11997 874
rect 11597 800 11997 840
rect 11597 766 11744 800
rect 11778 766 11816 800
rect 11850 766 11997 800
rect 11597 726 11997 766
rect 11597 692 11744 726
rect 11778 692 11816 726
rect 11850 692 11997 726
rect 11597 652 11997 692
rect 11597 618 11744 652
rect 11778 618 11816 652
rect 11850 618 11997 652
rect 11597 578 11997 618
rect 11597 544 11744 578
rect 11778 544 11816 578
rect 11850 544 11997 578
rect 11597 504 11997 544
rect 11597 470 11744 504
rect 11778 470 11816 504
rect 11850 470 11997 504
rect 11597 430 11997 470
rect 11597 396 11744 430
rect 11778 396 11816 430
rect 11850 396 11997 430
rect 11597 356 11997 396
rect 11597 322 11744 356
rect 11778 322 11816 356
rect 11850 322 11997 356
rect 11597 282 11997 322
rect 11597 248 11744 282
rect 11778 248 11816 282
rect 11850 248 11997 282
rect 11597 208 11997 248
rect 11597 174 11744 208
rect 11778 174 11816 208
rect 11850 174 11997 208
rect 11597 134 11997 174
rect 11597 100 11744 134
rect 11778 100 11816 134
rect 11850 100 11997 134
rect 11597 47 11997 100
tri 11597 42 11602 47 ne
rect 11602 42 11992 47
tri 11992 42 11997 47 nw
tri 12109 3053 12156 3100 se
rect 12156 3053 12262 3100
tri 12262 3053 12309 3100 sw
rect 12109 3000 12309 3053
rect 12109 2966 12156 3000
rect 12190 2966 12228 3000
rect 12262 2966 12309 3000
rect 12109 2927 12309 2966
rect 12109 2893 12156 2927
rect 12190 2893 12228 2927
rect 12262 2893 12309 2927
rect 12109 2854 12309 2893
rect 12109 2820 12156 2854
rect 12190 2820 12228 2854
rect 12262 2820 12309 2854
rect 12109 2781 12309 2820
rect 12109 2747 12156 2781
rect 12190 2747 12228 2781
rect 12262 2747 12309 2781
rect 12109 2708 12309 2747
rect 12109 2674 12156 2708
rect 12190 2674 12228 2708
rect 12262 2674 12309 2708
rect 12109 2635 12309 2674
rect 12109 2601 12156 2635
rect 12190 2601 12228 2635
rect 12262 2601 12309 2635
rect 12109 2562 12309 2601
rect 12109 2528 12156 2562
rect 12190 2528 12228 2562
rect 12262 2528 12309 2562
rect 12109 2489 12309 2528
rect 12109 2455 12156 2489
rect 12190 2455 12228 2489
rect 12262 2455 12309 2489
rect 12109 2416 12309 2455
rect 12109 2382 12156 2416
rect 12190 2382 12228 2416
rect 12262 2382 12309 2416
rect 12109 2343 12309 2382
rect 12109 2309 12156 2343
rect 12190 2309 12228 2343
rect 12262 2309 12309 2343
rect 12109 2270 12309 2309
rect 12109 2236 12156 2270
rect 12190 2236 12228 2270
rect 12262 2236 12309 2270
rect 12109 2197 12309 2236
rect 12109 2163 12156 2197
rect 12190 2163 12228 2197
rect 12262 2163 12309 2197
rect 12109 2124 12309 2163
rect 12109 2090 12156 2124
rect 12190 2090 12228 2124
rect 12262 2090 12309 2124
rect 12109 2051 12309 2090
rect 12109 2017 12156 2051
rect 12190 2017 12228 2051
rect 12262 2017 12309 2051
rect 12109 1978 12309 2017
rect 12109 1944 12156 1978
rect 12190 1944 12228 1978
rect 12262 1944 12309 1978
rect 12109 1905 12309 1944
rect 12109 1871 12156 1905
rect 12190 1871 12228 1905
rect 12262 1871 12309 1905
rect 12109 1832 12309 1871
rect 12109 1798 12156 1832
rect 12190 1798 12228 1832
rect 12262 1798 12309 1832
rect 12109 1759 12309 1798
rect 12109 1725 12156 1759
rect 12190 1725 12228 1759
rect 12262 1725 12309 1759
rect 12109 1686 12309 1725
rect 12109 1652 12156 1686
rect 12190 1652 12228 1686
rect 12262 1652 12309 1686
rect 12109 1613 12309 1652
rect 12109 1579 12156 1613
rect 12190 1579 12228 1613
rect 12262 1579 12309 1613
rect 12109 1540 12309 1579
rect 12109 1506 12156 1540
rect 12190 1506 12228 1540
rect 12262 1506 12309 1540
rect 12109 1466 12309 1506
rect 12109 1432 12156 1466
rect 12190 1432 12228 1466
rect 12262 1432 12309 1466
rect 12109 1392 12309 1432
rect 12109 1358 12156 1392
rect 12190 1358 12228 1392
rect 12262 1358 12309 1392
rect 12109 1318 12309 1358
rect 12109 1284 12156 1318
rect 12190 1284 12228 1318
rect 12262 1284 12309 1318
rect 12109 1244 12309 1284
rect 12109 1210 12156 1244
rect 12190 1210 12228 1244
rect 12262 1210 12309 1244
rect 12109 1170 12309 1210
rect 12109 1136 12156 1170
rect 12190 1136 12228 1170
rect 12262 1136 12309 1170
rect 12109 1096 12309 1136
rect 12109 1062 12156 1096
rect 12190 1062 12228 1096
rect 12262 1062 12309 1096
rect 12109 1022 12309 1062
rect 12109 988 12156 1022
rect 12190 988 12228 1022
rect 12262 988 12309 1022
rect 12109 948 12309 988
rect 12109 914 12156 948
rect 12190 914 12228 948
rect 12262 914 12309 948
rect 12109 874 12309 914
rect 12109 840 12156 874
rect 12190 840 12228 874
rect 12262 840 12309 874
rect 12109 800 12309 840
rect 12109 766 12156 800
rect 12190 766 12228 800
rect 12262 766 12309 800
rect 12109 726 12309 766
rect 12109 692 12156 726
rect 12190 692 12228 726
rect 12262 692 12309 726
rect 12109 652 12309 692
rect 12109 618 12156 652
rect 12190 618 12228 652
rect 12262 618 12309 652
rect 12109 578 12309 618
rect 12109 544 12156 578
rect 12190 544 12228 578
rect 12262 544 12309 578
rect 12109 504 12309 544
rect 12109 470 12156 504
rect 12190 470 12228 504
rect 12262 470 12309 504
rect 12109 430 12309 470
rect 12109 396 12156 430
rect 12190 396 12228 430
rect 12262 396 12309 430
rect 12109 356 12309 396
rect 12109 322 12156 356
rect 12190 322 12228 356
rect 12262 322 12309 356
rect 12109 282 12309 322
rect 12109 248 12156 282
rect 12190 248 12228 282
rect 12262 248 12309 282
rect 12109 208 12309 248
rect 12109 174 12156 208
rect 12190 174 12228 208
rect 12262 174 12309 208
rect 12109 134 12309 174
rect 12109 100 12156 134
rect 12190 100 12228 134
rect 12262 100 12309 134
rect 12109 47 12309 100
tri 12109 42 12114 47 ne
rect 12114 42 12304 47
tri 12304 42 12309 47 nw
tri 12421 3053 12468 3100 se
rect 12468 3053 12774 3100
tri 12774 3053 12821 3100 sw
rect 12421 3000 12821 3053
rect 12421 2966 12568 3000
rect 12602 2966 12640 3000
rect 12674 2966 12821 3000
rect 12421 2927 12821 2966
rect 12421 2893 12568 2927
rect 12602 2893 12640 2927
rect 12674 2893 12821 2927
rect 12421 2854 12821 2893
rect 12421 2820 12568 2854
rect 12602 2820 12640 2854
rect 12674 2820 12821 2854
rect 12421 2781 12821 2820
rect 12421 2747 12568 2781
rect 12602 2747 12640 2781
rect 12674 2747 12821 2781
rect 12421 2708 12821 2747
rect 12421 2674 12568 2708
rect 12602 2674 12640 2708
rect 12674 2674 12821 2708
rect 12421 2635 12821 2674
rect 12421 2601 12568 2635
rect 12602 2601 12640 2635
rect 12674 2601 12821 2635
rect 12421 2562 12821 2601
rect 12421 2528 12568 2562
rect 12602 2528 12640 2562
rect 12674 2528 12821 2562
rect 12421 2489 12821 2528
rect 12421 2455 12568 2489
rect 12602 2455 12640 2489
rect 12674 2455 12821 2489
rect 12421 2416 12821 2455
rect 12421 2382 12568 2416
rect 12602 2382 12640 2416
rect 12674 2382 12821 2416
rect 12421 2343 12821 2382
rect 12421 2309 12568 2343
rect 12602 2309 12640 2343
rect 12674 2309 12821 2343
rect 12421 2270 12821 2309
rect 12421 2236 12568 2270
rect 12602 2236 12640 2270
rect 12674 2236 12821 2270
rect 12421 2197 12821 2236
rect 12421 2163 12568 2197
rect 12602 2163 12640 2197
rect 12674 2163 12821 2197
rect 12421 2124 12821 2163
rect 12421 2090 12568 2124
rect 12602 2090 12640 2124
rect 12674 2090 12821 2124
rect 12421 2051 12821 2090
rect 12421 2017 12568 2051
rect 12602 2017 12640 2051
rect 12674 2017 12821 2051
rect 12421 1978 12821 2017
rect 12421 1944 12568 1978
rect 12602 1944 12640 1978
rect 12674 1944 12821 1978
rect 12421 1905 12821 1944
rect 12421 1871 12568 1905
rect 12602 1871 12640 1905
rect 12674 1871 12821 1905
rect 12421 1832 12821 1871
rect 12421 1798 12568 1832
rect 12602 1798 12640 1832
rect 12674 1798 12821 1832
rect 12421 1759 12821 1798
rect 12421 1725 12568 1759
rect 12602 1725 12640 1759
rect 12674 1725 12821 1759
rect 12421 1686 12821 1725
rect 12421 1652 12568 1686
rect 12602 1652 12640 1686
rect 12674 1652 12821 1686
rect 12421 1613 12821 1652
rect 12421 1579 12568 1613
rect 12602 1579 12640 1613
rect 12674 1579 12821 1613
rect 12421 1540 12821 1579
rect 12421 1506 12568 1540
rect 12602 1506 12640 1540
rect 12674 1506 12821 1540
rect 12421 1466 12821 1506
rect 12421 1432 12568 1466
rect 12602 1432 12640 1466
rect 12674 1432 12821 1466
rect 12421 1392 12821 1432
rect 12421 1358 12568 1392
rect 12602 1358 12640 1392
rect 12674 1358 12821 1392
rect 12421 1318 12821 1358
rect 12421 1284 12568 1318
rect 12602 1284 12640 1318
rect 12674 1284 12821 1318
rect 12421 1244 12821 1284
rect 12421 1210 12568 1244
rect 12602 1210 12640 1244
rect 12674 1210 12821 1244
rect 12421 1170 12821 1210
rect 12421 1136 12568 1170
rect 12602 1136 12640 1170
rect 12674 1136 12821 1170
rect 12421 1096 12821 1136
rect 12421 1062 12568 1096
rect 12602 1062 12640 1096
rect 12674 1062 12821 1096
rect 12421 1022 12821 1062
rect 12421 988 12568 1022
rect 12602 988 12640 1022
rect 12674 988 12821 1022
rect 12421 948 12821 988
rect 12421 914 12568 948
rect 12602 914 12640 948
rect 12674 914 12821 948
rect 12421 874 12821 914
rect 12421 840 12568 874
rect 12602 840 12640 874
rect 12674 840 12821 874
rect 12421 800 12821 840
rect 12421 766 12568 800
rect 12602 766 12640 800
rect 12674 766 12821 800
rect 12421 726 12821 766
rect 12421 692 12568 726
rect 12602 692 12640 726
rect 12674 692 12821 726
rect 12421 652 12821 692
rect 12421 618 12568 652
rect 12602 618 12640 652
rect 12674 618 12821 652
rect 12421 578 12821 618
rect 12421 544 12568 578
rect 12602 544 12640 578
rect 12674 544 12821 578
rect 12421 504 12821 544
rect 12421 470 12568 504
rect 12602 470 12640 504
rect 12674 470 12821 504
rect 12421 430 12821 470
rect 12421 396 12568 430
rect 12602 396 12640 430
rect 12674 396 12821 430
rect 12421 356 12821 396
rect 12421 322 12568 356
rect 12602 322 12640 356
rect 12674 322 12821 356
rect 12421 282 12821 322
rect 12421 248 12568 282
rect 12602 248 12640 282
rect 12674 248 12821 282
rect 12421 208 12821 248
rect 12421 174 12568 208
rect 12602 174 12640 208
rect 12674 174 12821 208
rect 12421 134 12821 174
rect 12421 100 12568 134
rect 12602 100 12640 134
rect 12674 100 12821 134
rect 12421 47 12821 100
tri 12421 42 12426 47 ne
rect 12426 42 12816 47
tri 12816 42 12821 47 nw
tri 12933 3053 12980 3100 se
rect 12980 3053 13086 3100
tri 13086 3053 13133 3100 sw
rect 12933 3000 13133 3053
rect 12933 2966 12980 3000
rect 13014 2966 13052 3000
rect 13086 2966 13133 3000
rect 12933 2927 13133 2966
rect 12933 2893 12980 2927
rect 13014 2893 13052 2927
rect 13086 2893 13133 2927
rect 12933 2854 13133 2893
rect 12933 2820 12980 2854
rect 13014 2820 13052 2854
rect 13086 2820 13133 2854
rect 12933 2781 13133 2820
rect 12933 2747 12980 2781
rect 13014 2747 13052 2781
rect 13086 2747 13133 2781
rect 12933 2708 13133 2747
rect 12933 2674 12980 2708
rect 13014 2674 13052 2708
rect 13086 2674 13133 2708
rect 12933 2635 13133 2674
rect 12933 2601 12980 2635
rect 13014 2601 13052 2635
rect 13086 2601 13133 2635
rect 12933 2562 13133 2601
rect 12933 2528 12980 2562
rect 13014 2528 13052 2562
rect 13086 2528 13133 2562
rect 12933 2489 13133 2528
rect 12933 2455 12980 2489
rect 13014 2455 13052 2489
rect 13086 2455 13133 2489
rect 12933 2416 13133 2455
rect 12933 2382 12980 2416
rect 13014 2382 13052 2416
rect 13086 2382 13133 2416
rect 12933 2343 13133 2382
rect 12933 2309 12980 2343
rect 13014 2309 13052 2343
rect 13086 2309 13133 2343
rect 12933 2270 13133 2309
rect 12933 2236 12980 2270
rect 13014 2236 13052 2270
rect 13086 2236 13133 2270
rect 12933 2197 13133 2236
rect 12933 2163 12980 2197
rect 13014 2163 13052 2197
rect 13086 2163 13133 2197
rect 12933 2124 13133 2163
rect 12933 2090 12980 2124
rect 13014 2090 13052 2124
rect 13086 2090 13133 2124
rect 12933 2051 13133 2090
rect 12933 2017 12980 2051
rect 13014 2017 13052 2051
rect 13086 2017 13133 2051
rect 12933 1978 13133 2017
rect 12933 1944 12980 1978
rect 13014 1944 13052 1978
rect 13086 1944 13133 1978
rect 12933 1905 13133 1944
rect 12933 1871 12980 1905
rect 13014 1871 13052 1905
rect 13086 1871 13133 1905
rect 12933 1832 13133 1871
rect 12933 1798 12980 1832
rect 13014 1798 13052 1832
rect 13086 1798 13133 1832
rect 12933 1759 13133 1798
rect 12933 1725 12980 1759
rect 13014 1725 13052 1759
rect 13086 1725 13133 1759
rect 12933 1686 13133 1725
rect 12933 1652 12980 1686
rect 13014 1652 13052 1686
rect 13086 1652 13133 1686
rect 12933 1613 13133 1652
rect 12933 1579 12980 1613
rect 13014 1579 13052 1613
rect 13086 1579 13133 1613
rect 12933 1540 13133 1579
rect 12933 1506 12980 1540
rect 13014 1506 13052 1540
rect 13086 1506 13133 1540
rect 12933 1466 13133 1506
rect 12933 1432 12980 1466
rect 13014 1432 13052 1466
rect 13086 1432 13133 1466
rect 12933 1392 13133 1432
rect 12933 1358 12980 1392
rect 13014 1358 13052 1392
rect 13086 1358 13133 1392
rect 12933 1318 13133 1358
rect 12933 1284 12980 1318
rect 13014 1284 13052 1318
rect 13086 1284 13133 1318
rect 12933 1244 13133 1284
rect 12933 1210 12980 1244
rect 13014 1210 13052 1244
rect 13086 1210 13133 1244
rect 12933 1170 13133 1210
rect 12933 1136 12980 1170
rect 13014 1136 13052 1170
rect 13086 1136 13133 1170
rect 12933 1096 13133 1136
rect 12933 1062 12980 1096
rect 13014 1062 13052 1096
rect 13086 1062 13133 1096
rect 12933 1022 13133 1062
rect 12933 988 12980 1022
rect 13014 988 13052 1022
rect 13086 988 13133 1022
rect 12933 948 13133 988
rect 12933 914 12980 948
rect 13014 914 13052 948
rect 13086 914 13133 948
rect 12933 874 13133 914
rect 12933 840 12980 874
rect 13014 840 13052 874
rect 13086 840 13133 874
rect 12933 800 13133 840
rect 12933 766 12980 800
rect 13014 766 13052 800
rect 13086 766 13133 800
rect 12933 726 13133 766
rect 12933 692 12980 726
rect 13014 692 13052 726
rect 13086 692 13133 726
rect 12933 652 13133 692
rect 12933 618 12980 652
rect 13014 618 13052 652
rect 13086 618 13133 652
rect 12933 578 13133 618
rect 12933 544 12980 578
rect 13014 544 13052 578
rect 13086 544 13133 578
rect 12933 504 13133 544
rect 12933 470 12980 504
rect 13014 470 13052 504
rect 13086 470 13133 504
rect 12933 430 13133 470
rect 12933 396 12980 430
rect 13014 396 13052 430
rect 13086 396 13133 430
rect 12933 356 13133 396
rect 12933 322 12980 356
rect 13014 322 13052 356
rect 13086 322 13133 356
rect 12933 282 13133 322
rect 12933 248 12980 282
rect 13014 248 13052 282
rect 13086 248 13133 282
rect 12933 208 13133 248
rect 12933 174 12980 208
rect 13014 174 13052 208
rect 13086 174 13133 208
rect 12933 134 13133 174
rect 12933 100 12980 134
rect 13014 100 13052 134
rect 13086 100 13133 134
rect 12933 47 13133 100
tri 12933 42 12938 47 ne
rect 12938 42 13128 47
tri 13128 42 13133 47 nw
rect 13190 2451 13202 3277
rect 13956 2451 13968 3277
rect 13190 2412 13968 2451
rect 13190 2378 13202 2412
rect 13236 2378 13274 2412
rect 13308 2378 13346 2412
rect 13380 2378 13418 2412
rect 13452 2378 13490 2412
rect 13524 2378 13562 2412
rect 13596 2378 13634 2412
rect 13668 2378 13706 2412
rect 13740 2378 13778 2412
rect 13812 2378 13850 2412
rect 13884 2378 13922 2412
rect 13956 2378 13968 2412
rect 13190 2339 13968 2378
rect 13190 2305 13202 2339
rect 13236 2305 13274 2339
rect 13308 2305 13346 2339
rect 13380 2305 13418 2339
rect 13452 2305 13490 2339
rect 13524 2305 13562 2339
rect 13596 2305 13634 2339
rect 13668 2305 13706 2339
rect 13740 2305 13778 2339
rect 13812 2305 13850 2339
rect 13884 2305 13922 2339
rect 13956 2305 13968 2339
rect 13190 2266 13968 2305
rect 13190 2232 13202 2266
rect 13236 2232 13274 2266
rect 13308 2232 13346 2266
rect 13380 2232 13418 2266
rect 13452 2232 13490 2266
rect 13524 2232 13562 2266
rect 13596 2232 13634 2266
rect 13668 2232 13706 2266
rect 13740 2232 13778 2266
rect 13812 2232 13850 2266
rect 13884 2232 13922 2266
rect 13956 2232 13968 2266
rect 13190 2193 13968 2232
rect 13190 2159 13202 2193
rect 13236 2159 13274 2193
rect 13308 2159 13346 2193
rect 13380 2159 13418 2193
rect 13452 2159 13490 2193
rect 13524 2159 13562 2193
rect 13596 2159 13634 2193
rect 13668 2159 13706 2193
rect 13740 2159 13778 2193
rect 13812 2159 13850 2193
rect 13884 2159 13922 2193
rect 13956 2159 13968 2193
rect 13190 2120 13968 2159
rect 13190 2086 13202 2120
rect 13236 2086 13274 2120
rect 13308 2086 13346 2120
rect 13380 2086 13418 2120
rect 13452 2086 13490 2120
rect 13524 2086 13562 2120
rect 13596 2086 13634 2120
rect 13668 2086 13706 2120
rect 13740 2086 13778 2120
rect 13812 2086 13850 2120
rect 13884 2086 13922 2120
rect 13956 2086 13968 2120
rect 13190 2047 13968 2086
rect 13190 2013 13202 2047
rect 13236 2013 13274 2047
rect 13308 2013 13346 2047
rect 13380 2013 13418 2047
rect 13452 2013 13490 2047
rect 13524 2013 13562 2047
rect 13596 2013 13634 2047
rect 13668 2013 13706 2047
rect 13740 2013 13778 2047
rect 13812 2013 13850 2047
rect 13884 2013 13922 2047
rect 13956 2013 13968 2047
rect 13190 1974 13968 2013
rect 13190 1940 13202 1974
rect 13236 1940 13274 1974
rect 13308 1940 13346 1974
rect 13380 1940 13418 1974
rect 13452 1940 13490 1974
rect 13524 1940 13562 1974
rect 13596 1940 13634 1974
rect 13668 1940 13706 1974
rect 13740 1940 13778 1974
rect 13812 1940 13850 1974
rect 13884 1940 13922 1974
rect 13956 1940 13968 1974
rect 13190 1901 13968 1940
rect 13190 1867 13202 1901
rect 13236 1867 13274 1901
rect 13308 1867 13346 1901
rect 13380 1867 13418 1901
rect 13452 1867 13490 1901
rect 13524 1867 13562 1901
rect 13596 1867 13634 1901
rect 13668 1867 13706 1901
rect 13740 1867 13778 1901
rect 13812 1867 13850 1901
rect 13884 1867 13922 1901
rect 13956 1867 13968 1901
rect 13190 1828 13968 1867
rect 13190 1794 13202 1828
rect 13236 1794 13274 1828
rect 13308 1794 13346 1828
rect 13380 1794 13418 1828
rect 13452 1794 13490 1828
rect 13524 1794 13562 1828
rect 13596 1794 13634 1828
rect 13668 1794 13706 1828
rect 13740 1794 13778 1828
rect 13812 1794 13850 1828
rect 13884 1794 13922 1828
rect 13956 1794 13968 1828
rect 13190 1755 13968 1794
rect 13190 1721 13202 1755
rect 13236 1721 13274 1755
rect 13308 1721 13346 1755
rect 13380 1721 13418 1755
rect 13452 1721 13490 1755
rect 13524 1721 13562 1755
rect 13596 1721 13634 1755
rect 13668 1721 13706 1755
rect 13740 1721 13778 1755
rect 13812 1721 13850 1755
rect 13884 1721 13922 1755
rect 13956 1721 13968 1755
rect 13190 1682 13968 1721
rect 13190 1648 13202 1682
rect 13236 1648 13274 1682
rect 13308 1648 13346 1682
rect 13380 1648 13418 1682
rect 13452 1648 13490 1682
rect 13524 1648 13562 1682
rect 13596 1648 13634 1682
rect 13668 1648 13706 1682
rect 13740 1648 13778 1682
rect 13812 1648 13850 1682
rect 13884 1648 13922 1682
rect 13956 1648 13968 1682
rect 13190 1609 13968 1648
rect 13190 1575 13202 1609
rect 13236 1575 13274 1609
rect 13308 1575 13346 1609
rect 13380 1575 13418 1609
rect 13452 1575 13490 1609
rect 13524 1575 13562 1609
rect 13596 1575 13634 1609
rect 13668 1575 13706 1609
rect 13740 1575 13778 1609
rect 13812 1575 13850 1609
rect 13884 1575 13922 1609
rect 13956 1575 13968 1609
rect 13190 1536 13968 1575
rect 13190 1502 13202 1536
rect 13236 1502 13274 1536
rect 13308 1502 13346 1536
rect 13380 1502 13418 1536
rect 13452 1502 13490 1536
rect 13524 1502 13562 1536
rect 13596 1502 13634 1536
rect 13668 1502 13706 1536
rect 13740 1502 13778 1536
rect 13812 1502 13850 1536
rect 13884 1502 13922 1536
rect 13956 1502 13968 1536
rect 13190 1463 13968 1502
rect 13190 1429 13202 1463
rect 13236 1429 13274 1463
rect 13308 1429 13346 1463
rect 13380 1429 13418 1463
rect 13452 1429 13490 1463
rect 13524 1429 13562 1463
rect 13596 1429 13634 1463
rect 13668 1429 13706 1463
rect 13740 1429 13778 1463
rect 13812 1429 13850 1463
rect 13884 1429 13922 1463
rect 13956 1429 13968 1463
rect 13190 1390 13968 1429
rect 13190 1356 13202 1390
rect 13236 1356 13274 1390
rect 13308 1356 13346 1390
rect 13380 1356 13418 1390
rect 13452 1356 13490 1390
rect 13524 1356 13562 1390
rect 13596 1356 13634 1390
rect 13668 1356 13706 1390
rect 13740 1356 13778 1390
rect 13812 1356 13850 1390
rect 13884 1356 13922 1390
rect 13956 1356 13968 1390
rect 13190 1317 13968 1356
rect 13190 1283 13202 1317
rect 13236 1283 13274 1317
rect 13308 1283 13346 1317
rect 13380 1283 13418 1317
rect 13452 1283 13490 1317
rect 13524 1283 13562 1317
rect 13596 1283 13634 1317
rect 13668 1283 13706 1317
rect 13740 1283 13778 1317
rect 13812 1283 13850 1317
rect 13884 1283 13922 1317
rect 13956 1283 13968 1317
rect 13190 1244 13968 1283
rect 13190 1210 13202 1244
rect 13236 1210 13274 1244
rect 13308 1210 13346 1244
rect 13380 1210 13418 1244
rect 13452 1210 13490 1244
rect 13524 1210 13562 1244
rect 13596 1210 13634 1244
rect 13668 1210 13706 1244
rect 13740 1210 13778 1244
rect 13812 1210 13850 1244
rect 13884 1210 13922 1244
rect 13956 1210 13968 1244
rect 13190 1171 13968 1210
rect 13190 1137 13202 1171
rect 13236 1137 13274 1171
rect 13308 1137 13346 1171
rect 13380 1137 13418 1171
rect 13452 1137 13490 1171
rect 13524 1137 13562 1171
rect 13596 1137 13634 1171
rect 13668 1137 13706 1171
rect 13740 1137 13778 1171
rect 13812 1137 13850 1171
rect 13884 1137 13922 1171
rect 13956 1137 13968 1171
rect 13190 1098 13968 1137
rect 13190 1064 13202 1098
rect 13236 1064 13274 1098
rect 13308 1064 13346 1098
rect 13380 1064 13418 1098
rect 13452 1064 13490 1098
rect 13524 1064 13562 1098
rect 13596 1064 13634 1098
rect 13668 1064 13706 1098
rect 13740 1064 13778 1098
rect 13812 1064 13850 1098
rect 13884 1064 13922 1098
rect 13956 1064 13968 1098
rect 13190 1025 13968 1064
rect 13190 991 13202 1025
rect 13236 991 13274 1025
rect 13308 991 13346 1025
rect 13380 991 13418 1025
rect 13452 991 13490 1025
rect 13524 991 13562 1025
rect 13596 991 13634 1025
rect 13668 991 13706 1025
rect 13740 991 13778 1025
rect 13812 991 13850 1025
rect 13884 991 13922 1025
rect 13956 991 13968 1025
rect 13190 952 13968 991
rect 13190 918 13202 952
rect 13236 918 13274 952
rect 13308 918 13346 952
rect 13380 918 13418 952
rect 13452 918 13490 952
rect 13524 918 13562 952
rect 13596 918 13634 952
rect 13668 918 13706 952
rect 13740 918 13778 952
rect 13812 918 13850 952
rect 13884 918 13922 952
rect 13956 918 13968 952
rect 13190 879 13968 918
rect 13190 845 13202 879
rect 13236 845 13274 879
rect 13308 845 13346 879
rect 13380 845 13418 879
rect 13452 845 13490 879
rect 13524 845 13562 879
rect 13596 845 13634 879
rect 13668 845 13706 879
rect 13740 845 13778 879
rect 13812 845 13850 879
rect 13884 845 13922 879
rect 13956 845 13968 879
rect 13190 806 13968 845
rect 13190 772 13202 806
rect 13236 772 13274 806
rect 13308 772 13346 806
rect 13380 772 13418 806
rect 13452 772 13490 806
rect 13524 772 13562 806
rect 13596 772 13634 806
rect 13668 772 13706 806
rect 13740 772 13778 806
rect 13812 772 13850 806
rect 13884 772 13922 806
rect 13956 772 13968 806
rect 13190 733 13968 772
rect 13190 699 13202 733
rect 13236 699 13274 733
rect 13308 699 13346 733
rect 13380 699 13418 733
rect 13452 699 13490 733
rect 13524 699 13562 733
rect 13596 699 13634 733
rect 13668 699 13706 733
rect 13740 699 13778 733
rect 13812 699 13850 733
rect 13884 699 13922 733
rect 13956 699 13968 733
rect 13190 660 13968 699
rect 13190 626 13202 660
rect 13236 626 13274 660
rect 13308 626 13346 660
rect 13380 626 13418 660
rect 13452 626 13490 660
rect 13524 626 13562 660
rect 13596 626 13634 660
rect 13668 626 13706 660
rect 13740 626 13778 660
rect 13812 626 13850 660
rect 13884 626 13922 660
rect 13956 626 13968 660
rect 13190 587 13968 626
rect 13190 553 13202 587
rect 13236 553 13274 587
rect 13308 553 13346 587
rect 13380 553 13418 587
rect 13452 553 13490 587
rect 13524 553 13562 587
rect 13596 553 13634 587
rect 13668 553 13706 587
rect 13740 553 13778 587
rect 13812 553 13850 587
rect 13884 553 13922 587
rect 13956 553 13968 587
rect 13190 514 13968 553
rect 13190 480 13202 514
rect 13236 480 13274 514
rect 13308 480 13346 514
rect 13380 480 13418 514
rect 13452 480 13490 514
rect 13524 480 13562 514
rect 13596 480 13634 514
rect 13668 480 13706 514
rect 13740 480 13778 514
rect 13812 480 13850 514
rect 13884 480 13922 514
rect 13956 480 13968 514
rect 13190 441 13968 480
rect 13190 407 13202 441
rect 13236 407 13274 441
rect 13308 407 13346 441
rect 13380 407 13418 441
rect 13452 407 13490 441
rect 13524 407 13562 441
rect 13596 407 13634 441
rect 13668 407 13706 441
rect 13740 407 13778 441
rect 13812 407 13850 441
rect 13884 407 13922 441
rect 13956 407 13968 441
rect 13190 368 13968 407
rect 13190 334 13202 368
rect 13236 334 13274 368
rect 13308 334 13346 368
rect 13380 334 13418 368
rect 13452 334 13490 368
rect 13524 334 13562 368
rect 13596 334 13634 368
rect 13668 334 13706 368
rect 13740 334 13778 368
rect 13812 334 13850 368
rect 13884 334 13922 368
rect 13956 334 13968 368
rect 13190 295 13968 334
rect 13190 261 13202 295
rect 13236 261 13274 295
rect 13308 261 13346 295
rect 13380 261 13418 295
rect 13452 261 13490 295
rect 13524 261 13562 295
rect 13596 261 13634 295
rect 13668 261 13706 295
rect 13740 261 13778 295
rect 13812 261 13850 295
rect 13884 261 13922 295
rect 13956 261 13968 295
rect 13190 222 13968 261
rect 13190 188 13202 222
rect 13236 188 13274 222
rect 13308 188 13346 222
rect 13380 188 13418 222
rect 13452 188 13490 222
rect 13524 188 13562 222
rect 13596 188 13634 222
rect 13668 188 13706 222
rect 13740 188 13778 222
rect 13812 188 13850 222
rect 13884 188 13922 222
rect 13956 188 13968 222
rect 13190 149 13968 188
rect 13190 115 13202 149
rect 13236 115 13274 149
rect 13308 115 13346 149
rect 13380 115 13418 149
rect 13452 115 13490 149
rect 13524 115 13562 149
rect 13596 115 13634 149
rect 13668 115 13706 149
rect 13740 115 13778 149
rect 13812 115 13850 149
rect 13884 115 13922 149
rect 13956 115 13968 149
rect 13190 76 13968 115
rect 13190 42 13202 76
rect 13236 42 13274 76
rect 13308 42 13346 76
rect 13380 42 13418 76
rect 13452 42 13490 76
rect 13524 42 13562 76
rect 13596 42 13634 76
rect 13668 42 13706 76
rect 13740 42 13778 76
rect 13812 42 13850 76
rect 13884 42 13922 76
rect 13956 42 13968 76
rect -1086 3 -308 42
tri -246 37 -241 42 ne
rect -241 37 -61 42
tri -61 37 -56 42 nw
tri 66 37 71 42 ne
rect 71 37 451 42
tri 451 37 456 42 nw
tri 578 37 583 42 ne
rect 583 37 763 42
tri 763 37 768 42 nw
tri 890 37 895 42 ne
rect 895 37 1275 42
tri 1275 37 1280 42 nw
tri 1402 37 1407 42 ne
rect 1407 37 1587 42
tri 1587 37 1592 42 nw
tri 1714 37 1719 42 ne
rect 1719 37 2099 42
tri 2099 37 2104 42 nw
tri 2226 37 2231 42 ne
rect 2231 37 2411 42
tri 2411 37 2416 42 nw
tri 2538 37 2543 42 ne
rect 2543 37 2923 42
tri 2923 37 2928 42 nw
tri 3050 37 3055 42 ne
rect 3055 37 3235 42
tri 3235 37 3240 42 nw
tri 3362 37 3367 42 ne
rect 3367 37 3747 42
tri 3747 37 3752 42 nw
tri 3874 37 3879 42 ne
rect 3879 37 4059 42
tri 4059 37 4064 42 nw
tri 4186 37 4191 42 ne
rect 4191 37 4571 42
tri 4571 37 4576 42 nw
tri 4698 37 4703 42 ne
rect 4703 37 4883 42
tri 4883 37 4888 42 nw
tri 5010 37 5015 42 ne
rect 5015 37 5395 42
tri 5395 37 5400 42 nw
tri 5522 37 5527 42 ne
rect 5527 37 5707 42
tri 5707 37 5712 42 nw
tri 5834 37 5839 42 ne
rect 5839 37 6219 42
tri 6219 37 6224 42 nw
tri 6346 37 6351 42 ne
rect 6351 37 6531 42
tri 6531 37 6536 42 nw
tri 6658 37 6663 42 ne
rect 6663 37 7043 42
tri 7043 37 7048 42 nw
tri 7170 37 7175 42 ne
rect 7175 37 7355 42
tri 7355 37 7360 42 nw
tri 7482 37 7487 42 ne
rect 7487 37 7867 42
tri 7867 37 7872 42 nw
tri 7994 37 7999 42 ne
rect 7999 37 8179 42
tri 8179 37 8184 42 nw
tri 8306 37 8311 42 ne
rect 8311 37 8691 42
tri 8691 37 8696 42 nw
tri 8818 37 8823 42 ne
rect 8823 37 9003 42
tri 9003 37 9008 42 nw
tri 9130 37 9135 42 ne
rect 9135 37 9515 42
tri 9515 37 9520 42 nw
tri 9642 37 9647 42 ne
rect 9647 37 9827 42
tri 9827 37 9832 42 nw
tri 9954 37 9959 42 ne
rect 9959 37 10339 42
tri 10339 37 10344 42 nw
tri 10466 37 10471 42 ne
rect 10471 37 10651 42
tri 10651 37 10656 42 nw
tri 10778 37 10783 42 ne
rect 10783 37 11163 42
tri 11163 37 11168 42 nw
tri 11290 37 11295 42 ne
rect 11295 37 11475 42
tri 11475 37 11480 42 nw
tri 11602 37 11607 42 ne
rect 11607 37 11987 42
tri 11987 37 11992 42 nw
tri 12114 37 12119 42 ne
rect 12119 37 12299 42
tri 12299 37 12304 42 nw
tri 12426 37 12431 42 ne
rect 12431 37 12811 42
tri 12811 37 12816 42 nw
tri 12938 37 12943 42 ne
rect 12943 37 13123 42
tri 13123 37 13128 42 nw
tri -241 3 -207 37 ne
rect -207 3 -95 37
tri -95 3 -61 37 nw
tri 71 3 105 37 ne
rect 105 3 417 37
tri 417 3 451 37 nw
tri 583 3 617 37 ne
rect 617 3 729 37
tri 729 3 763 37 nw
tri 895 3 929 37 ne
rect 929 3 1241 37
tri 1241 3 1275 37 nw
tri 1407 3 1441 37 ne
rect 1441 3 1553 37
tri 1553 3 1587 37 nw
tri 1719 3 1753 37 ne
rect 1753 3 2065 37
tri 2065 3 2099 37 nw
tri 2231 3 2265 37 ne
rect 2265 3 2377 37
tri 2377 3 2411 37 nw
tri 2543 3 2577 37 ne
rect 2577 3 2889 37
tri 2889 3 2923 37 nw
tri 3055 3 3089 37 ne
rect 3089 3 3201 37
tri 3201 3 3235 37 nw
tri 3367 3 3401 37 ne
rect 3401 3 3713 37
tri 3713 3 3747 37 nw
tri 3879 3 3913 37 ne
rect 3913 3 4025 37
tri 4025 3 4059 37 nw
tri 4191 3 4225 37 ne
rect 4225 3 4537 37
tri 4537 3 4571 37 nw
tri 4703 3 4737 37 ne
rect 4737 3 4849 37
tri 4849 3 4883 37 nw
tri 5015 3 5049 37 ne
rect 5049 3 5361 37
tri 5361 3 5395 37 nw
tri 5527 3 5561 37 ne
rect 5561 3 5673 37
tri 5673 3 5707 37 nw
tri 5839 3 5873 37 ne
rect 5873 3 6185 37
tri 6185 3 6219 37 nw
tri 6351 3 6385 37 ne
rect 6385 3 6497 37
tri 6497 3 6531 37 nw
tri 6663 3 6697 37 ne
rect 6697 3 7009 37
tri 7009 3 7043 37 nw
tri 7175 3 7209 37 ne
rect 7209 3 7321 37
tri 7321 3 7355 37 nw
tri 7487 3 7521 37 ne
rect 7521 3 7833 37
tri 7833 3 7867 37 nw
tri 7999 3 8033 37 ne
rect 8033 3 8145 37
tri 8145 3 8179 37 nw
tri 8311 3 8345 37 ne
rect 8345 3 8657 37
tri 8657 3 8691 37 nw
tri 8823 3 8857 37 ne
rect 8857 3 8969 37
tri 8969 3 9003 37 nw
tri 9135 3 9169 37 ne
rect 9169 3 9481 37
tri 9481 3 9515 37 nw
tri 9647 3 9681 37 ne
rect 9681 3 9793 37
tri 9793 3 9827 37 nw
tri 9959 3 9993 37 ne
rect 9993 3 10305 37
tri 10305 3 10339 37 nw
tri 10471 3 10505 37 ne
rect 10505 3 10617 37
tri 10617 3 10651 37 nw
tri 10783 3 10817 37 ne
rect 10817 3 11129 37
tri 11129 3 11163 37 nw
tri 11295 3 11329 37 ne
rect 11329 3 11441 37
tri 11441 3 11475 37 nw
tri 11607 3 11641 37 ne
rect 11641 3 11953 37
tri 11953 3 11987 37 nw
tri 12119 3 12153 37 ne
rect 12153 3 12265 37
tri 12265 3 12299 37 nw
tri 12431 3 12465 37 ne
rect 12465 3 12777 37
tri 12777 3 12811 37 nw
tri 12943 3 12977 37 ne
rect 12977 3 13089 37
tri 13089 3 13123 37 nw
rect 13190 3 13968 42
rect -1086 -31 -1074 3
rect -1040 -31 -1002 3
rect -968 -31 -930 3
rect -896 -31 -858 3
rect -824 -31 -786 3
rect -752 -31 -714 3
rect -680 -31 -642 3
rect -608 -31 -570 3
rect -536 -31 -498 3
rect -464 -31 -426 3
rect -392 -31 -354 3
rect -320 -31 -308 3
tri -207 0 -204 3 ne
rect -204 0 -98 3
tri -98 0 -95 3 nw
tri 105 0 108 3 ne
rect 108 0 414 3
tri 414 0 417 3 nw
tri 617 0 620 3 ne
rect 620 0 726 3
tri 726 0 729 3 nw
tri 929 0 932 3 ne
rect 932 0 1238 3
tri 1238 0 1241 3 nw
tri 1441 0 1444 3 ne
rect 1444 0 1550 3
tri 1550 0 1553 3 nw
tri 1753 0 1756 3 ne
rect 1756 0 2062 3
tri 2062 0 2065 3 nw
tri 2265 0 2268 3 ne
rect 2268 0 2374 3
tri 2374 0 2377 3 nw
tri 2577 0 2580 3 ne
rect 2580 0 2886 3
tri 2886 0 2889 3 nw
tri 3089 0 3092 3 ne
rect 3092 0 3198 3
tri 3198 0 3201 3 nw
tri 3401 0 3404 3 ne
rect 3404 0 3710 3
tri 3710 0 3713 3 nw
tri 3913 0 3916 3 ne
rect 3916 0 4022 3
tri 4022 0 4025 3 nw
tri 4225 0 4228 3 ne
rect 4228 0 4534 3
tri 4534 0 4537 3 nw
tri 4737 0 4740 3 ne
rect 4740 0 4846 3
tri 4846 0 4849 3 nw
tri 5049 0 5052 3 ne
rect 5052 0 5358 3
tri 5358 0 5361 3 nw
tri 5561 0 5564 3 ne
rect 5564 0 5670 3
tri 5670 0 5673 3 nw
tri 5873 0 5876 3 ne
rect 5876 0 6182 3
tri 6182 0 6185 3 nw
tri 6385 0 6388 3 ne
rect 6388 0 6494 3
tri 6494 0 6497 3 nw
tri 6697 0 6700 3 ne
rect 6700 0 7006 3
tri 7006 0 7009 3 nw
tri 7209 0 7212 3 ne
rect 7212 0 7318 3
tri 7318 0 7321 3 nw
tri 7521 0 7524 3 ne
rect 7524 0 7830 3
tri 7830 0 7833 3 nw
tri 8033 0 8036 3 ne
rect 8036 0 8142 3
tri 8142 0 8145 3 nw
tri 8345 0 8348 3 ne
rect 8348 0 8654 3
tri 8654 0 8657 3 nw
tri 8857 0 8860 3 ne
rect 8860 0 8966 3
tri 8966 0 8969 3 nw
tri 9169 0 9172 3 ne
rect 9172 0 9478 3
tri 9478 0 9481 3 nw
tri 9681 0 9684 3 ne
rect 9684 0 9790 3
tri 9790 0 9793 3 nw
tri 9993 0 9996 3 ne
rect 9996 0 10302 3
tri 10302 0 10305 3 nw
tri 10505 0 10508 3 ne
rect 10508 0 10614 3
tri 10614 0 10617 3 nw
tri 10817 0 10820 3 ne
rect 10820 0 11126 3
tri 11126 0 11129 3 nw
tri 11329 0 11332 3 ne
rect 11332 0 11438 3
tri 11438 0 11441 3 nw
tri 11641 0 11644 3 ne
rect 11644 0 11950 3
tri 11950 0 11953 3 nw
tri 12153 0 12156 3 ne
rect 12156 0 12262 3
tri 12262 0 12265 3 nw
tri 12465 0 12468 3 ne
rect 12468 0 12774 3
tri 12774 0 12777 3 nw
tri 12977 0 12980 3 ne
rect 12980 0 13086 3
tri 13086 0 13089 3 nw
rect -1086 -70 -308 -31
rect -1086 -104 -1074 -70
rect -1040 -104 -1002 -70
rect -968 -104 -930 -70
rect -896 -104 -858 -70
rect -824 -104 -786 -70
rect -752 -104 -714 -70
rect -680 -104 -642 -70
rect -608 -104 -570 -70
rect -536 -104 -498 -70
rect -464 -104 -426 -70
rect -392 -104 -354 -70
rect -320 -104 -308 -70
rect -1086 -143 -308 -104
rect -1086 -177 -1074 -143
rect -1040 -177 -1002 -143
rect -968 -177 -930 -143
rect -896 -177 -858 -143
rect -824 -177 -786 -143
rect -752 -177 -714 -143
rect -680 -177 -642 -143
rect -608 -177 -570 -143
rect -536 -177 -498 -143
rect -464 -177 -426 -143
rect -392 -177 -354 -143
rect -320 -177 -308 -143
rect -1086 -221 -308 -177
rect 13190 -31 13202 3
rect 13236 -31 13274 3
rect 13308 -31 13346 3
rect 13380 -31 13418 3
rect 13452 -31 13490 3
rect 13524 -31 13562 3
rect 13596 -31 13634 3
rect 13668 -31 13706 3
rect 13740 -31 13778 3
rect 13812 -31 13850 3
rect 13884 -31 13922 3
rect 13956 -31 13968 3
rect 13190 -70 13968 -31
rect 13190 -104 13202 -70
rect 13236 -104 13274 -70
rect 13308 -104 13346 -70
rect 13380 -104 13418 -70
rect 13452 -104 13490 -70
rect 13524 -104 13562 -70
rect 13596 -104 13634 -70
rect 13668 -104 13706 -70
rect 13740 -104 13778 -70
rect 13812 -104 13850 -70
rect 13884 -104 13922 -70
rect 13956 -104 13968 -70
rect 13190 -143 13968 -104
rect 13190 -177 13202 -143
rect 13236 -177 13274 -143
rect 13308 -177 13346 -143
rect 13380 -177 13418 -143
rect 13452 -177 13490 -143
rect 13524 -177 13562 -143
rect 13596 -177 13634 -143
rect 13668 -177 13706 -143
rect 13740 -177 13778 -143
rect 13812 -177 13850 -143
rect 13884 -177 13922 -143
rect 13956 -177 13968 -143
tri -308 -221 -284 -197 sw
tri 13166 -221 13190 -197 se
rect 13190 -221 13968 -177
rect -1086 -249 -284 -221
tri -284 -249 -256 -221 sw
tri 13138 -249 13166 -221 se
rect 13166 -249 13968 -221
rect -1086 -255 -256 -249
tri -256 -255 -250 -249 sw
tri 13132 -255 13138 -249 se
rect 13138 -255 13968 -249
rect -1086 -294 -250 -255
tri -250 -294 -211 -255 sw
tri 13093 -294 13132 -255 se
rect 13132 -294 13968 -255
tri -1086 -306 -1074 -294 ne
rect -1074 -306 13934 -294
rect -1438 -367 -1308 -328
tri -1074 -340 -1040 -306 ne
rect -1040 -340 -886 -306
rect -852 -340 -813 -306
rect -779 -340 -740 -306
rect -706 -340 -667 -306
rect -633 -340 -594 -306
rect -1438 -401 -1426 -367
rect -1392 -401 -1354 -367
rect -1320 -401 -1308 -367
tri -1040 -378 -1002 -340 ne
rect -1002 -378 -594 -340
rect -1438 -440 -1308 -401
tri -1002 -412 -968 -378 ne
rect -968 -412 -886 -378
rect -852 -412 -813 -378
rect -779 -412 -740 -378
rect -706 -412 -667 -378
rect -633 -412 -594 -378
rect 13768 -328 13934 -306
tri 13934 -328 13968 -294 nw
rect 14190 3356 14320 3395
rect 14190 3322 14202 3356
rect 14236 3322 14274 3356
rect 14308 3322 14320 3356
rect 14190 3283 14320 3322
rect 14190 3249 14202 3283
rect 14236 3249 14274 3283
rect 14308 3249 14320 3283
rect 14190 3210 14320 3249
rect 14190 3176 14202 3210
rect 14236 3176 14274 3210
rect 14308 3176 14320 3210
rect 14190 3137 14320 3176
rect 14190 3103 14202 3137
rect 14236 3103 14274 3137
rect 14308 3103 14320 3137
rect 14190 3064 14320 3103
rect 14190 3030 14202 3064
rect 14236 3030 14274 3064
rect 14308 3030 14320 3064
rect 14190 2991 14320 3030
rect 14190 2957 14202 2991
rect 14236 2957 14274 2991
rect 14308 2957 14320 2991
rect 14190 2918 14320 2957
rect 14190 2884 14202 2918
rect 14236 2884 14274 2918
rect 14308 2884 14320 2918
rect 14190 2845 14320 2884
rect 14190 2811 14202 2845
rect 14236 2811 14274 2845
rect 14308 2811 14320 2845
rect 14190 2772 14320 2811
rect 14190 2738 14202 2772
rect 14236 2738 14274 2772
rect 14308 2738 14320 2772
rect 14190 2699 14320 2738
rect 14190 2665 14202 2699
rect 14236 2665 14274 2699
rect 14308 2665 14320 2699
rect 14190 2626 14320 2665
rect 14190 2592 14202 2626
rect 14236 2592 14274 2626
rect 14308 2592 14320 2626
rect 14190 2553 14320 2592
rect 14190 2519 14202 2553
rect 14236 2519 14274 2553
rect 14308 2519 14320 2553
rect 14190 2480 14320 2519
rect 14190 2446 14202 2480
rect 14236 2446 14274 2480
rect 14308 2446 14320 2480
rect 14190 2407 14320 2446
rect 14190 2373 14202 2407
rect 14236 2373 14274 2407
rect 14308 2373 14320 2407
rect 14190 2334 14320 2373
rect 14190 2300 14202 2334
rect 14236 2300 14274 2334
rect 14308 2300 14320 2334
rect 14190 2261 14320 2300
rect 14190 2227 14202 2261
rect 14236 2227 14274 2261
rect 14308 2227 14320 2261
rect 14190 2188 14320 2227
rect 14190 2154 14202 2188
rect 14236 2154 14274 2188
rect 14308 2154 14320 2188
rect 14190 2115 14320 2154
rect 14190 2081 14202 2115
rect 14236 2081 14274 2115
rect 14308 2081 14320 2115
rect 14190 2042 14320 2081
rect 14190 2008 14202 2042
rect 14236 2008 14274 2042
rect 14308 2008 14320 2042
rect 14190 1969 14320 2008
rect 14190 1935 14202 1969
rect 14236 1935 14274 1969
rect 14308 1935 14320 1969
rect 14190 1896 14320 1935
rect 14190 1862 14202 1896
rect 14236 1862 14274 1896
rect 14308 1862 14320 1896
rect 14190 1823 14320 1862
rect 14190 1789 14202 1823
rect 14236 1789 14274 1823
rect 14308 1789 14320 1823
rect 14190 1750 14320 1789
rect 14190 1716 14202 1750
rect 14236 1716 14274 1750
rect 14308 1716 14320 1750
rect 14190 1677 14320 1716
rect 14190 1643 14202 1677
rect 14236 1643 14274 1677
rect 14308 1643 14320 1677
rect 14190 1604 14320 1643
rect 14190 1570 14202 1604
rect 14236 1570 14274 1604
rect 14308 1570 14320 1604
rect 14190 1531 14320 1570
rect 14190 1497 14202 1531
rect 14236 1497 14274 1531
rect 14308 1497 14320 1531
rect 14190 1458 14320 1497
rect 14190 1424 14202 1458
rect 14236 1424 14274 1458
rect 14308 1424 14320 1458
rect 14190 1385 14320 1424
rect 14190 1351 14202 1385
rect 14236 1351 14274 1385
rect 14308 1351 14320 1385
rect 14190 1312 14320 1351
rect 14190 1278 14202 1312
rect 14236 1278 14274 1312
rect 14308 1278 14320 1312
rect 14190 1239 14320 1278
rect 14190 1205 14202 1239
rect 14236 1205 14274 1239
rect 14308 1205 14320 1239
rect 14190 1166 14320 1205
rect 14190 1132 14202 1166
rect 14236 1132 14274 1166
rect 14308 1132 14320 1166
rect 14190 1093 14320 1132
rect 14190 1059 14202 1093
rect 14236 1059 14274 1093
rect 14308 1059 14320 1093
rect 14190 1020 14320 1059
rect 14190 986 14202 1020
rect 14236 986 14274 1020
rect 14308 986 14320 1020
rect 14190 947 14320 986
rect 14190 913 14202 947
rect 14236 913 14274 947
rect 14308 913 14320 947
rect 14190 874 14320 913
rect 14190 840 14202 874
rect 14236 840 14274 874
rect 14308 840 14320 874
rect 14190 801 14320 840
rect 14190 767 14202 801
rect 14236 767 14274 801
rect 14308 767 14320 801
rect 14190 728 14320 767
rect 14190 694 14202 728
rect 14236 694 14274 728
rect 14308 694 14320 728
rect 14190 655 14320 694
rect 14190 621 14202 655
rect 14236 621 14274 655
rect 14308 621 14320 655
rect 14190 582 14320 621
rect 14190 548 14202 582
rect 14236 548 14274 582
rect 14308 548 14320 582
rect 14190 509 14320 548
rect 14190 475 14202 509
rect 14236 475 14274 509
rect 14308 475 14320 509
rect 14190 436 14320 475
rect 14190 402 14202 436
rect 14236 402 14274 436
rect 14308 402 14320 436
rect 14190 363 14320 402
rect 14190 329 14202 363
rect 14236 329 14274 363
rect 14308 329 14320 363
rect 14190 290 14320 329
rect 14190 256 14202 290
rect 14236 256 14274 290
rect 14308 256 14320 290
rect 14190 217 14320 256
rect 14190 183 14202 217
rect 14236 183 14274 217
rect 14308 183 14320 217
rect 14190 144 14320 183
rect 14190 110 14202 144
rect 14236 110 14274 144
rect 14308 110 14320 144
rect 14190 71 14320 110
rect 14190 37 14202 71
rect 14236 37 14274 71
rect 14308 37 14320 71
rect 14190 -2 14320 37
rect 14190 -36 14202 -2
rect 14236 -36 14274 -2
rect 14308 -36 14320 -2
rect 14190 -75 14320 -36
rect 14190 -109 14202 -75
rect 14236 -109 14274 -75
rect 14308 -109 14320 -75
rect 14190 -148 14320 -109
rect 14190 -182 14202 -148
rect 14236 -182 14274 -148
rect 14308 -182 14320 -148
rect 14190 -221 14320 -182
rect 14190 -255 14202 -221
rect 14236 -255 14274 -221
rect 14308 -255 14320 -221
rect 14190 -294 14320 -255
rect 14190 -328 14202 -294
rect 14236 -328 14274 -294
rect 14308 -328 14320 -294
rect 13768 -367 13895 -328
tri 13895 -367 13934 -328 nw
rect 14190 -367 14320 -328
rect 13768 -401 13861 -367
tri 13861 -401 13895 -367 nw
rect 14190 -401 14202 -367
rect 14236 -401 14274 -367
rect 14308 -401 14320 -367
rect 13768 -412 13840 -401
tri -968 -422 -958 -412 ne
rect -958 -424 13840 -412
tri 13840 -422 13861 -401 nw
rect -1438 -474 -1426 -440
rect -1392 -474 -1354 -440
rect -1320 -474 -1308 -440
rect -1438 -513 -1308 -474
rect -1438 -547 -1426 -513
rect -1392 -547 -1354 -513
rect -1320 -547 -1308 -513
rect -1438 -619 -1308 -547
rect 14190 -440 14320 -401
rect 14190 -474 14202 -440
rect 14236 -474 14274 -440
rect 14308 -474 14320 -440
rect 14190 -513 14320 -474
rect 14190 -547 14202 -513
rect 14236 -547 14274 -513
rect 14308 -547 14320 -513
tri -1308 -619 -1245 -556 sw
tri 14127 -619 14190 -556 se
rect 14190 -619 14320 -547
rect -1438 -664 -1245 -619
tri -1245 -664 -1200 -619 sw
tri 14082 -664 14127 -619 se
rect 14127 -664 14320 -619
tri -1438 -676 -1426 -664 ne
rect -1426 -676 14190 -664
tri -1426 -710 -1392 -676 ne
rect -1392 -710 -1191 -676
rect -1157 -710 -1118 -676
rect -1084 -710 -1045 -676
rect -1011 -710 -972 -676
rect -938 -710 -899 -676
rect -865 -710 -826 -676
rect -792 -710 -753 -676
rect -719 -710 -680 -676
rect -646 -710 -607 -676
rect -573 -710 -534 -676
rect -500 -710 -461 -676
rect -427 -710 -388 -676
rect -354 -710 -315 -676
rect -281 -710 -242 -676
rect -208 -710 -169 -676
rect -135 -710 -96 -676
rect -62 -710 -23 -676
rect 11 -710 50 -676
rect 84 -710 123 -676
rect 157 -710 196 -676
rect 230 -710 269 -676
rect 303 -710 342 -676
rect 376 -710 415 -676
rect 449 -710 488 -676
rect 522 -710 561 -676
rect 595 -710 634 -676
rect 668 -710 707 -676
rect 741 -710 780 -676
rect 814 -710 853 -676
rect 887 -710 926 -676
rect 960 -710 999 -676
rect 1033 -710 1072 -676
rect 1106 -710 1145 -676
rect 1179 -710 1218 -676
rect 1252 -710 1291 -676
rect 1325 -710 1364 -676
rect 1398 -710 1437 -676
rect 1471 -710 1510 -676
rect 1544 -710 1583 -676
tri -1392 -748 -1354 -710 ne
rect -1354 -748 1583 -710
tri -1354 -782 -1320 -748 ne
rect -1320 -782 -1191 -748
rect -1157 -782 -1118 -748
rect -1084 -782 -1045 -748
rect -1011 -782 -972 -748
rect -938 -782 -899 -748
rect -865 -782 -826 -748
rect -792 -782 -753 -748
rect -719 -782 -680 -748
rect -646 -782 -607 -748
rect -573 -782 -534 -748
rect -500 -782 -461 -748
rect -427 -782 -388 -748
rect -354 -782 -315 -748
rect -281 -782 -242 -748
rect -208 -782 -169 -748
rect -135 -782 -96 -748
rect -62 -782 -23 -748
rect 11 -782 50 -748
rect 84 -782 123 -748
rect 157 -782 196 -748
rect 230 -782 269 -748
rect 303 -782 342 -748
rect 376 -782 415 -748
rect 449 -782 488 -748
rect 522 -782 561 -748
rect 595 -782 634 -748
rect 668 -782 707 -748
rect 741 -782 780 -748
rect 814 -782 853 -748
rect 887 -782 926 -748
rect 960 -782 999 -748
rect 1033 -782 1072 -748
rect 1106 -782 1145 -748
rect 1179 -782 1218 -748
rect 1252 -782 1291 -748
rect 1325 -782 1364 -748
rect 1398 -782 1437 -748
rect 1471 -782 1510 -748
rect 1544 -782 1583 -748
rect 14073 -782 14190 -676
tri -1320 -794 -1308 -782 ne
rect -1308 -794 14190 -782
tri 14190 -794 14320 -664 nw
<< labels >>
flabel comment s -151 1550 -151 1550 0 FreeSans 1600 0 0 0 S
flabel comment s 673 1550 673 1550 0 FreeSans 1600 0 0 0 S
flabel comment s 1497 1550 1497 1550 0 FreeSans 1600 0 0 0 S
flabel comment s 2321 1550 2321 1550 0 FreeSans 1600 0 0 0 S
flabel comment s 3145 1550 3145 1550 0 FreeSans 1600 0 0 0 S
flabel comment s 3969 1550 3969 1550 0 FreeSans 1600 0 0 0 S
flabel comment s 4793 1550 4793 1550 0 FreeSans 1600 0 0 0 S
flabel comment s 5617 1550 5617 1550 0 FreeSans 1600 0 0 0 S
flabel comment s 6441 1550 6441 1550 0 FreeSans 1600 0 0 0 S
flabel comment s 7265 1550 7265 1550 0 FreeSans 1600 0 0 0 S
flabel comment s 8089 1550 8089 1550 0 FreeSans 1600 0 0 0 S
flabel comment s 8913 1550 8913 1550 0 FreeSans 1600 0 0 0 S
flabel comment s 9737 1550 9737 1550 0 FreeSans 1600 0 0 0 S
flabel comment s 10561 1550 10561 1550 0 FreeSans 1600 0 0 0 S
flabel comment s 11385 1550 11385 1550 0 FreeSans 1600 0 0 0 S
flabel comment s 12209 1550 12209 1550 0 FreeSans 1600 0 0 0 S
flabel comment s 13033 1550 13033 1550 0 FreeSans 1600 0 0 0 S
flabel comment s 261 1550 261 1550 0 FreeSans 1600 0 0 0 D
flabel comment s 1085 1550 1085 1550 0 FreeSans 1600 0 0 0 D
flabel comment s 1909 1550 1909 1550 0 FreeSans 1600 0 0 0 D
flabel comment s 2733 1550 2733 1550 0 FreeSans 1600 0 0 0 D
flabel comment s 3557 1550 3557 1550 0 FreeSans 1600 0 0 0 D
flabel comment s 4381 1550 4381 1550 0 FreeSans 1600 0 0 0 D
flabel comment s 5205 1550 5205 1550 0 FreeSans 1600 0 0 0 D
flabel comment s 6029 1550 6029 1550 0 FreeSans 1600 0 0 0 D
flabel comment s 6853 1550 6853 1550 0 FreeSans 1600 0 0 0 D
flabel comment s 7677 1550 7677 1550 0 FreeSans 1600 0 0 0 D
flabel comment s 8501 1550 8501 1550 0 FreeSans 1600 0 0 0 D
flabel comment s 9325 1550 9325 1550 0 FreeSans 1600 0 0 0 D
flabel comment s 10149 1550 10149 1550 0 FreeSans 1600 0 0 0 D
flabel comment s 10973 1550 10973 1550 0 FreeSans 1600 0 0 0 D
flabel comment s 11797 1550 11797 1550 0 FreeSans 1600 0 0 0 D
flabel comment s 12621 1550 12621 1550 0 FreeSans 1600 0 0 0 D
flabel comment s -697 1900 -697 1900 0 FreeSans 800 0 0 0 CRITICAL TO
flabel comment s -697 1780 -697 1780 0 FreeSans 800 0 0 0 CONNECT WIDE
flabel comment s -697 1660 -697 1660 0 FreeSans 800 0 0 0 SIDES OF
flabel comment s -697 1540 -697 1540 0 FreeSans 800 0 0 0 GUARDRING
flabel comment s 13579 1900 13579 1900 0 FreeSans 800 0 0 0 CRITICAL TO
flabel comment s 13579 1780 13579 1780 0 FreeSans 800 0 0 0 CONNECT WIDE
flabel comment s 13579 1660 13579 1660 0 FreeSans 800 0 0 0 SIDES OF
flabel comment s 13579 1540 13579 1540 0 FreeSans 800 0 0 0 GUARDRING
<< properties >>
string GDS_END 91719338
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 90882822
<< end >>
