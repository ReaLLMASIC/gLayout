magic
tech sky130B
timestamp 1701704242
<< metal1 >>
rect 0 0 3 58
rect 1981 0 1984 58
<< via1 >>
rect 3 0 1981 58
<< metal2 >>
rect 0 0 3 58
rect 1981 0 1984 58
<< properties >>
string GDS_END 78479622
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 78471554
<< end >>
