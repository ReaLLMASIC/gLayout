magic
tech sky130B
timestamp 1701704242
<< poly >>
rect 0 25 271 33
rect 0 8 8 25
rect 25 8 42 25
rect 59 8 76 25
rect 93 8 110 25
rect 127 8 144 25
rect 161 8 178 25
rect 195 8 212 25
rect 229 8 246 25
rect 263 8 271 25
rect 0 0 271 8
<< polycont >>
rect 8 8 25 25
rect 42 8 59 25
rect 76 8 93 25
rect 110 8 127 25
rect 144 8 161 25
rect 178 8 195 25
rect 212 8 229 25
rect 246 8 263 25
<< locali >>
rect 0 8 8 25
rect 25 8 42 25
rect 59 8 76 25
rect 93 8 110 25
rect 127 8 144 25
rect 161 8 178 25
rect 195 8 212 25
rect 229 8 246 25
rect 263 8 271 25
<< properties >>
string GDS_END 90863864
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 90863156
<< end >>
