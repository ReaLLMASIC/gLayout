magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -36 679 2240 1471
<< locali >>
rect 0 1397 2204 1431
rect 64 674 98 740
rect 1047 690 1081 724
rect 0 -17 2204 17
use sky130_sram_2kbyte_1rw1r_32x512_8_pinv_16  sky130_sram_2kbyte_1rw1r_32x512_8_pinv_16_0
timestamp 1701704242
transform 1 0 0 0 1 0
box -36 -17 2240 1471
<< labels >>
rlabel locali s 1064 707 1064 707 4 Z
rlabel locali s 81 707 81 707 4 A
rlabel locali s 1102 0 1102 0 4 gnd
rlabel locali s 1102 1414 1102 1414 4 vdd
<< properties >>
string FIXED_BBOX 0 0 2204 1414
string GDS_END 365692
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_2kbyte_1rw1r_32x512_8.gds
string GDS_START 364860
<< end >>
