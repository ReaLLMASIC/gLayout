magic
tech sky130B
timestamp 1701704242
<< properties >>
string GDS_END 22132186
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 22126204
<< end >>
