magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< pwell >>
rect -79 -26 279 176
<< mvnmos >>
rect 0 0 200 150
<< mvndiff >>
rect -53 114 0 150
rect -53 80 -45 114
rect -11 80 0 114
rect -53 46 0 80
rect -53 12 -45 46
rect -11 12 0 46
rect -53 0 0 12
rect 200 114 253 150
rect 200 80 211 114
rect 245 80 253 114
rect 200 46 253 80
rect 200 12 211 46
rect 245 12 253 46
rect 200 0 253 12
<< mvndiffc >>
rect -45 80 -11 114
rect -45 12 -11 46
rect 211 80 245 114
rect 211 12 245 46
<< poly >>
rect 0 150 200 176
rect 0 -26 200 0
<< locali >>
rect -45 114 -11 130
rect -45 46 -11 68
rect 211 114 245 130
rect 211 46 245 68
<< viali >>
rect -45 80 -11 102
rect -45 68 -11 80
rect -45 12 -11 30
rect -45 -4 -11 12
rect 211 80 245 102
rect 211 68 245 80
rect 211 12 245 30
rect 211 -4 245 12
<< metal1 >>
rect -51 102 -5 114
rect -51 68 -45 102
rect -11 68 -5 102
rect -51 30 -5 68
rect -51 -4 -45 30
rect -11 -4 -5 30
rect -51 -16 -5 -4
rect 205 102 251 114
rect 205 68 211 102
rect 245 68 251 102
rect 205 30 251 68
rect 205 -4 211 30
rect 245 -4 251 30
rect 205 -16 251 -4
use hvDFM1sd_CDNS_52468879185143  hvDFM1sd_CDNS_52468879185143_0
timestamp 1701704242
transform -1 0 0 0 1 0
box 0 0 1 1
use hvDFM1sd_CDNS_52468879185143  hvDFM1sd_CDNS_52468879185143_1
timestamp 1701704242
transform 1 0 200 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s -28 49 -28 49 0 FreeSans 300 0 0 0 S
flabel comment s 228 49 228 49 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 86851742
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86850852
<< end >>
