magic
tech sky130A
magscale 1 2
timestamp 1701704242
use sky130_fd_pr__dfm1sd__example_55959141808173  sky130_fd_pr__dfm1sd__example_55959141808173_0
timestamp 1701704242
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfm1sd__example_55959141808173  sky130_fd_pr__dfm1sd__example_55959141808173_1
timestamp 1701704242
transform 1 0 412 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_5595914180831  sky130_fd_pr__hvdfm1sd2__example_5595914180831_0
timestamp 1701704242
transform 1 0 100 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_5595914180831  sky130_fd_pr__hvdfm1sd2__example_5595914180831_1
timestamp 1701704242
transform 1 0 256 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 70312238
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 70310156
<< end >>
