magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< locali >>
rect 0 1397 1394 1431
rect 330 708 364 1151
rect 330 674 459 708
rect 883 674 917 708
rect 212 485 246 551
rect 112 237 146 303
rect 0 -17 1394 17
use sky130_sram_1kbyte_1rw1r_8x1024_8_pdriver_1  sky130_sram_1kbyte_1rw1r_8x1024_8_pdriver_1_0
timestamp 1701704242
transform 1 0 378 0 1 0
box -36 -17 1052 1471
use sky130_sram_1kbyte_1rw1r_8x1024_8_pnand2_0  sky130_sram_1kbyte_1rw1r_8x1024_8_pnand2_0_0
timestamp 1701704242
transform 1 0 0 0 1 0
box -36 -17 414 1471
<< labels >>
rlabel locali s 900 691 900 691 4 Z
rlabel locali s 129 270 129 270 4 A
rlabel locali s 229 518 229 518 4 B
rlabel locali s 697 0 697 0 4 gnd
rlabel locali s 697 1414 697 1414 4 vdd
<< properties >>
string FIXED_BBOX 0 0 1394 1414
string GDS_END 6093902
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_8x1024_8.gds
string GDS_START 6092760
<< end >>
