magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< dnwell >>
rect 17450 11681 17634 14661
rect 10345 1141 15400 1250
rect 6222 374 15400 1141
<< nwell >>
rect 17530 11761 17553 14581
rect -2860 2277 595 4834
rect 2214 3637 4515 4595
rect 11092 3637 11764 4594
rect 2214 3335 11764 3637
rect 2214 2277 4515 3335
rect -2860 1957 4515 2277
rect -2860 1956 2256 1957
rect 10133 1227 15486 1336
rect 6136 1044 15486 1227
rect 6136 935 10425 1044
rect 6136 371 6428 935
rect 15194 382 15486 1044
<< pwell >>
rect 11923 3266 17241 4387
rect 4589 2150 17241 3266
rect 4589 2149 16758 2150
rect 4589 1896 5742 2149
rect -2885 745 5742 1896
rect -2885 742 5737 745
rect 10502 883 14970 983
rect 10502 865 10602 883
rect 6526 765 10602 865
rect 15912 -2975 16758 2149
rect 15913 -3001 16758 -2975
<< pdiff >>
rect 28689 -1431 28721 -1397
rect 30587 -1431 30615 -1397
rect 28695 -2401 28721 -2367
rect 30587 -2401 30613 -2367
<< psubdiff >>
rect -2859 1846 2 1870
rect -2825 1812 -2790 1846
rect -2756 1812 -2721 1846
rect -2687 1812 -2652 1846
rect -2618 1812 -2583 1846
rect -2549 1812 -2514 1846
rect -2480 1812 -2445 1846
rect -2411 1812 -2376 1846
rect -2342 1812 -2307 1846
rect -2273 1812 -2238 1846
rect -2204 1812 -2169 1846
rect -2135 1812 -2100 1846
rect -2066 1812 -2031 1846
rect -1997 1812 -1962 1846
rect -1928 1812 -1893 1846
rect -1859 1812 -1824 1846
rect -1790 1812 -1755 1846
rect -1721 1812 -1686 1846
rect -1652 1812 -1617 1846
rect -1583 1812 -1548 1846
rect -1514 1812 -1479 1846
rect -1445 1812 -1410 1846
rect -1376 1812 -1341 1846
rect -1307 1812 -1272 1846
rect -1238 1812 -1203 1846
rect -1169 1812 -1134 1846
rect -1100 1812 -1065 1846
rect -1031 1812 -996 1846
rect -962 1812 -927 1846
rect -893 1812 -858 1846
rect -824 1812 -789 1846
rect -755 1812 -720 1846
rect -686 1812 -651 1846
rect -617 1812 -582 1846
rect -548 1812 -513 1846
rect -479 1812 -444 1846
rect -410 1812 -375 1846
rect -2859 1778 -375 1812
rect -2825 1744 -2790 1778
rect -2756 1744 -2721 1778
rect -2687 1744 -2652 1778
rect -2618 1744 -2583 1778
rect -2549 1744 -2514 1778
rect -2480 1744 -2445 1778
rect -2411 1744 -2376 1778
rect -2342 1744 -2307 1778
rect -2273 1744 -2238 1778
rect -2204 1744 -2169 1778
rect -2135 1744 -2100 1778
rect -2066 1744 -2031 1778
rect -1997 1744 -1962 1778
rect -1928 1744 -1893 1778
rect -1859 1744 -1824 1778
rect -1790 1744 -1755 1778
rect -1721 1744 -1686 1778
rect -1652 1744 -1617 1778
rect -1583 1744 -1548 1778
rect -1514 1744 -1479 1778
rect -1445 1744 -1410 1778
rect -1376 1744 -1341 1778
rect -1307 1744 -1272 1778
rect -1238 1744 -1203 1778
rect -1169 1744 -1134 1778
rect -1100 1744 -1065 1778
rect -1031 1744 -996 1778
rect -962 1744 -927 1778
rect -893 1744 -858 1778
rect -824 1744 -789 1778
rect -755 1744 -720 1778
rect -686 1744 -651 1778
rect -617 1744 -582 1778
rect -548 1744 -513 1778
rect -479 1744 -444 1778
rect -410 1744 -375 1778
rect -2859 1710 -375 1744
rect -2825 1676 -2790 1710
rect -2756 1676 -2721 1710
rect -2687 1676 -2652 1710
rect -2618 1676 -2583 1710
rect -2549 1676 -2514 1710
rect -2480 1676 -2445 1710
rect -2411 1676 -2376 1710
rect -2342 1676 -2307 1710
rect -2273 1676 -2238 1710
rect -2204 1676 -2169 1710
rect -2135 1676 -2100 1710
rect -2066 1676 -2031 1710
rect -1997 1676 -1962 1710
rect -1928 1676 -1893 1710
rect -1859 1676 -1824 1710
rect -1790 1676 -1755 1710
rect -1721 1676 -1686 1710
rect -1652 1676 -1617 1710
rect -1583 1676 -1548 1710
rect -1514 1676 -1479 1710
rect -1445 1676 -1410 1710
rect -1376 1676 -1341 1710
rect -1307 1676 -1272 1710
rect -1238 1676 -1203 1710
rect -1169 1676 -1134 1710
rect -1100 1676 -1065 1710
rect -1031 1676 -996 1710
rect -962 1676 -927 1710
rect -893 1676 -858 1710
rect -824 1676 -789 1710
rect -755 1676 -720 1710
rect -686 1676 -651 1710
rect -617 1676 -582 1710
rect -548 1676 -513 1710
rect -479 1676 -444 1710
rect -410 1676 -375 1710
rect -2859 1642 -375 1676
rect -2825 1608 -2790 1642
rect -2756 1608 -2721 1642
rect -2687 1608 -2652 1642
rect -2618 1608 -2583 1642
rect -2549 1608 -2514 1642
rect -2480 1608 -2445 1642
rect -2411 1608 -2376 1642
rect -2342 1608 -2307 1642
rect -2273 1608 -2238 1642
rect -2204 1608 -2169 1642
rect -2135 1608 -2100 1642
rect -2066 1608 -2031 1642
rect -1997 1608 -1962 1642
rect -1928 1608 -1893 1642
rect -1859 1608 -1824 1642
rect -1790 1608 -1755 1642
rect -1721 1608 -1686 1642
rect -1652 1608 -1617 1642
rect -1583 1608 -1548 1642
rect -1514 1608 -1479 1642
rect -1445 1608 -1410 1642
rect -1376 1608 -1341 1642
rect -1307 1608 -1272 1642
rect -1238 1608 -1203 1642
rect -1169 1608 -1134 1642
rect -1100 1608 -1065 1642
rect -1031 1608 -996 1642
rect -962 1608 -927 1642
rect -893 1608 -858 1642
rect -824 1608 -789 1642
rect -755 1608 -720 1642
rect -686 1608 -651 1642
rect -617 1608 -582 1642
rect -548 1608 -513 1642
rect -479 1608 -444 1642
rect -410 1608 -375 1642
rect -2859 1574 -375 1608
rect -2825 1540 -2790 1574
rect -2756 1540 -2721 1574
rect -2687 1540 -2652 1574
rect -2618 1540 -2583 1574
rect -2549 1540 -2514 1574
rect -2480 1540 -2445 1574
rect -2411 1540 -2376 1574
rect -2342 1540 -2307 1574
rect -2273 1540 -2238 1574
rect -2204 1540 -2169 1574
rect -2135 1540 -2100 1574
rect -2066 1540 -2031 1574
rect -1997 1540 -1962 1574
rect -1928 1540 -1893 1574
rect -1859 1540 -1824 1574
rect -1790 1540 -1755 1574
rect -1721 1540 -1686 1574
rect -1652 1540 -1617 1574
rect -1583 1540 -1548 1574
rect -1514 1540 -1479 1574
rect -1445 1540 -1410 1574
rect -1376 1540 -1341 1574
rect -1307 1540 -1272 1574
rect -1238 1540 -1203 1574
rect -1169 1540 -1134 1574
rect -1100 1540 -1065 1574
rect -1031 1540 -996 1574
rect -962 1540 -927 1574
rect -893 1540 -858 1574
rect -824 1540 -789 1574
rect -755 1540 -720 1574
rect -686 1540 -651 1574
rect -617 1540 -582 1574
rect -548 1540 -513 1574
rect -479 1540 -444 1574
rect -410 1540 -375 1574
rect -2859 1506 -375 1540
rect -2825 1472 -2790 1506
rect -2756 1472 -2721 1506
rect -2687 1472 -2652 1506
rect -2618 1472 -2583 1506
rect -2549 1472 -2514 1506
rect -2480 1472 -2445 1506
rect -2411 1472 -2376 1506
rect -2342 1472 -2307 1506
rect -2273 1472 -2238 1506
rect -2204 1472 -2169 1506
rect -2135 1472 -2100 1506
rect -2066 1472 -2031 1506
rect -1997 1472 -1962 1506
rect -1928 1472 -1893 1506
rect -1859 1472 -1824 1506
rect -1790 1472 -1755 1506
rect -1721 1472 -1686 1506
rect -1652 1472 -1617 1506
rect -1583 1472 -1548 1506
rect -1514 1472 -1479 1506
rect -1445 1472 -1410 1506
rect -1376 1472 -1341 1506
rect -1307 1472 -1272 1506
rect -1238 1472 -1203 1506
rect -1169 1472 -1134 1506
rect -1100 1472 -1065 1506
rect -1031 1472 -996 1506
rect -962 1472 -927 1506
rect -893 1472 -858 1506
rect -824 1472 -789 1506
rect -755 1472 -720 1506
rect -686 1472 -651 1506
rect -617 1472 -582 1506
rect -548 1472 -513 1506
rect -479 1472 -444 1506
rect -410 1472 -375 1506
rect -2859 1438 -375 1472
rect -2825 1404 -2790 1438
rect -2756 1404 -2721 1438
rect -2687 1404 -2652 1438
rect -2618 1404 -2583 1438
rect -2549 1404 -2514 1438
rect -2480 1404 -2445 1438
rect -2411 1404 -2376 1438
rect -2342 1404 -2307 1438
rect -2273 1404 -2238 1438
rect -2204 1404 -2169 1438
rect -2135 1404 -2100 1438
rect -2066 1404 -2031 1438
rect -1997 1404 -1962 1438
rect -1928 1404 -1893 1438
rect -1859 1404 -1824 1438
rect -1790 1404 -1755 1438
rect -1721 1404 -1686 1438
rect -1652 1404 -1617 1438
rect -1583 1404 -1548 1438
rect -1514 1404 -1479 1438
rect -1445 1404 -1410 1438
rect -1376 1404 -1341 1438
rect -1307 1404 -1272 1438
rect -1238 1404 -1203 1438
rect -1169 1404 -1134 1438
rect -1100 1404 -1065 1438
rect -1031 1404 -996 1438
rect -962 1404 -927 1438
rect -893 1404 -858 1438
rect -824 1404 -789 1438
rect -755 1404 -720 1438
rect -686 1404 -651 1438
rect -617 1404 -582 1438
rect -548 1404 -513 1438
rect -479 1404 -444 1438
rect -410 1404 -375 1438
rect -2859 1370 -375 1404
rect -2825 1336 -2790 1370
rect -2756 1336 -2721 1370
rect -2687 1336 -2652 1370
rect -2618 1336 -2583 1370
rect -2549 1336 -2514 1370
rect -2480 1336 -2445 1370
rect -2411 1336 -2376 1370
rect -2342 1336 -2307 1370
rect -2273 1336 -2238 1370
rect -2204 1336 -2169 1370
rect -2135 1336 -2100 1370
rect -2066 1336 -2031 1370
rect -1997 1336 -1962 1370
rect -1928 1336 -1893 1370
rect -1859 1336 -1824 1370
rect -1790 1336 -1755 1370
rect -1721 1336 -1686 1370
rect -1652 1336 -1617 1370
rect -1583 1336 -1548 1370
rect -1514 1336 -1479 1370
rect -1445 1336 -1410 1370
rect -1376 1336 -1341 1370
rect -1307 1336 -1272 1370
rect -1238 1336 -1203 1370
rect -1169 1336 -1134 1370
rect -1100 1336 -1065 1370
rect -1031 1336 -996 1370
rect -962 1336 -927 1370
rect -893 1336 -858 1370
rect -824 1336 -789 1370
rect -755 1336 -720 1370
rect -686 1336 -651 1370
rect -617 1336 -582 1370
rect -548 1336 -513 1370
rect -479 1336 -444 1370
rect -410 1336 -375 1370
rect -2859 1302 -375 1336
rect -2825 1268 -2790 1302
rect -2756 1268 -2721 1302
rect -2687 1268 -2652 1302
rect -2618 1268 -2583 1302
rect -2549 1268 -2514 1302
rect -2480 1268 -2445 1302
rect -2411 1268 -2376 1302
rect -2342 1268 -2307 1302
rect -2273 1268 -2238 1302
rect -2204 1268 -2169 1302
rect -2135 1268 -2100 1302
rect -2066 1268 -2031 1302
rect -1997 1268 -1962 1302
rect -1928 1268 -1893 1302
rect -1859 1268 -1824 1302
rect -1790 1268 -1755 1302
rect -1721 1268 -1686 1302
rect -1652 1268 -1617 1302
rect -1583 1268 -1548 1302
rect -1514 1268 -1479 1302
rect -1445 1268 -1410 1302
rect -1376 1268 -1341 1302
rect -1307 1268 -1272 1302
rect -1238 1268 -1203 1302
rect -1169 1268 -1134 1302
rect -1100 1268 -1065 1302
rect -1031 1268 -996 1302
rect -962 1268 -927 1302
rect -893 1268 -858 1302
rect -824 1268 -789 1302
rect -755 1268 -720 1302
rect -686 1268 -651 1302
rect -617 1268 -582 1302
rect -548 1268 -513 1302
rect -479 1268 -444 1302
rect -410 1268 -375 1302
rect -2859 1234 -375 1268
rect -2825 1200 -2790 1234
rect -2756 1200 -2721 1234
rect -2687 1200 -2652 1234
rect -2618 1200 -2583 1234
rect -2549 1200 -2514 1234
rect -2480 1200 -2445 1234
rect -2411 1200 -2376 1234
rect -2342 1200 -2307 1234
rect -2273 1200 -2238 1234
rect -2204 1200 -2169 1234
rect -2135 1200 -2100 1234
rect -2066 1200 -2031 1234
rect -1997 1200 -1962 1234
rect -1928 1200 -1893 1234
rect -1859 1200 -1824 1234
rect -1790 1200 -1755 1234
rect -1721 1200 -1686 1234
rect -1652 1200 -1617 1234
rect -1583 1200 -1548 1234
rect -1514 1200 -1479 1234
rect -1445 1200 -1410 1234
rect -1376 1200 -1341 1234
rect -1307 1200 -1272 1234
rect -1238 1200 -1203 1234
rect -1169 1200 -1134 1234
rect -1100 1200 -1065 1234
rect -1031 1200 -996 1234
rect -962 1200 -927 1234
rect -893 1200 -858 1234
rect -824 1200 -789 1234
rect -755 1200 -720 1234
rect -686 1200 -651 1234
rect -617 1200 -582 1234
rect -548 1200 -513 1234
rect -479 1200 -444 1234
rect -410 1200 -375 1234
rect -2859 1166 -375 1200
rect -2825 1132 -2790 1166
rect -2756 1132 -2721 1166
rect -2687 1132 -2652 1166
rect -2618 1132 -2583 1166
rect -2549 1132 -2514 1166
rect -2480 1132 -2445 1166
rect -2411 1132 -2376 1166
rect -2342 1132 -2307 1166
rect -2273 1132 -2238 1166
rect -2204 1132 -2169 1166
rect -2135 1132 -2100 1166
rect -2066 1132 -2031 1166
rect -1997 1132 -1962 1166
rect -1928 1132 -1893 1166
rect -1859 1132 -1824 1166
rect -1790 1132 -1755 1166
rect -1721 1132 -1686 1166
rect -1652 1132 -1617 1166
rect -1583 1132 -1548 1166
rect -1514 1132 -1479 1166
rect -1445 1132 -1410 1166
rect -1376 1132 -1341 1166
rect -1307 1132 -1272 1166
rect -1238 1132 -1203 1166
rect -1169 1132 -1134 1166
rect -1100 1132 -1065 1166
rect -1031 1132 -996 1166
rect -962 1132 -927 1166
rect -893 1132 -858 1166
rect -824 1132 -789 1166
rect -755 1132 -720 1166
rect -686 1132 -651 1166
rect -617 1132 -582 1166
rect -548 1132 -513 1166
rect -479 1132 -444 1166
rect -410 1132 -375 1166
rect -2859 1098 -375 1132
rect -2825 1064 -2790 1098
rect -2756 1064 -2721 1098
rect -2687 1064 -2652 1098
rect -2618 1064 -2583 1098
rect -2549 1064 -2514 1098
rect -2480 1064 -2445 1098
rect -2411 1064 -2376 1098
rect -2342 1064 -2307 1098
rect -2273 1064 -2238 1098
rect -2204 1064 -2169 1098
rect -2135 1064 -2100 1098
rect -2066 1064 -2031 1098
rect -1997 1064 -1962 1098
rect -1928 1064 -1893 1098
rect -1859 1064 -1824 1098
rect -1790 1064 -1755 1098
rect -1721 1064 -1686 1098
rect -1652 1064 -1617 1098
rect -1583 1064 -1548 1098
rect -1514 1064 -1479 1098
rect -1445 1064 -1410 1098
rect -1376 1064 -1341 1098
rect -1307 1064 -1272 1098
rect -1238 1064 -1203 1098
rect -1169 1064 -1134 1098
rect -1100 1064 -1065 1098
rect -1031 1064 -996 1098
rect -962 1064 -927 1098
rect -893 1064 -858 1098
rect -824 1064 -789 1098
rect -755 1064 -720 1098
rect -686 1064 -651 1098
rect -617 1064 -582 1098
rect -548 1064 -513 1098
rect -479 1064 -444 1098
rect -410 1064 -375 1098
rect -2859 1030 -375 1064
rect -2825 996 -2790 1030
rect -2756 996 -2721 1030
rect -2687 996 -2652 1030
rect -2618 996 -2583 1030
rect -2549 996 -2514 1030
rect -2480 996 -2445 1030
rect -2411 996 -2376 1030
rect -2342 996 -2307 1030
rect -2273 996 -2238 1030
rect -2204 996 -2169 1030
rect -2135 996 -2100 1030
rect -2066 996 -2031 1030
rect -1997 996 -1962 1030
rect -1928 996 -1893 1030
rect -1859 996 -1824 1030
rect -1790 996 -1755 1030
rect -1721 996 -1686 1030
rect -1652 996 -1617 1030
rect -1583 996 -1548 1030
rect -1514 996 -1479 1030
rect -1445 996 -1410 1030
rect -1376 996 -1341 1030
rect -1307 996 -1272 1030
rect -1238 996 -1203 1030
rect -1169 996 -1134 1030
rect -1100 996 -1065 1030
rect -1031 996 -996 1030
rect -962 996 -927 1030
rect -893 996 -858 1030
rect -824 996 -789 1030
rect -755 996 -720 1030
rect -686 996 -651 1030
rect -617 996 -582 1030
rect -548 996 -513 1030
rect -479 996 -444 1030
rect -410 996 -375 1030
rect -2859 962 -375 996
rect -2825 928 -2790 962
rect -2756 928 -2721 962
rect -2687 928 -2652 962
rect -2618 928 -2583 962
rect -2549 928 -2514 962
rect -2480 928 -2445 962
rect -2411 928 -2376 962
rect -2342 928 -2307 962
rect -2273 928 -2238 962
rect -2204 928 -2169 962
rect -2135 928 -2100 962
rect -2066 928 -2031 962
rect -1997 928 -1962 962
rect -1928 928 -1893 962
rect -1859 928 -1824 962
rect -1790 928 -1755 962
rect -1721 928 -1686 962
rect -1652 928 -1617 962
rect -1583 928 -1548 962
rect -1514 928 -1479 962
rect -1445 928 -1410 962
rect -1376 928 -1341 962
rect -1307 928 -1272 962
rect -1238 928 -1203 962
rect -1169 928 -1134 962
rect -1100 928 -1065 962
rect -1031 928 -996 962
rect -962 928 -927 962
rect -893 928 -858 962
rect -824 928 -789 962
rect -755 928 -720 962
rect -686 928 -651 962
rect -617 928 -582 962
rect -548 928 -513 962
rect -479 928 -444 962
rect -410 928 -375 962
rect -2859 894 -375 928
rect -2825 860 -2790 894
rect -2756 860 -2721 894
rect -2687 860 -2652 894
rect -2618 860 -2583 894
rect -2549 860 -2514 894
rect -2480 860 -2445 894
rect -2411 860 -2376 894
rect -2342 860 -2307 894
rect -2273 860 -2238 894
rect -2204 860 -2169 894
rect -2135 860 -2100 894
rect -2066 860 -2031 894
rect -1997 860 -1962 894
rect -1928 860 -1893 894
rect -1859 860 -1824 894
rect -1790 860 -1755 894
rect -1721 860 -1686 894
rect -1652 860 -1617 894
rect -1583 860 -1548 894
rect -1514 860 -1479 894
rect -1445 860 -1410 894
rect -1376 860 -1341 894
rect -1307 860 -1272 894
rect -1238 860 -1203 894
rect -1169 860 -1134 894
rect -1100 860 -1065 894
rect -1031 860 -996 894
rect -962 860 -927 894
rect -893 860 -858 894
rect -824 860 -789 894
rect -755 860 -720 894
rect -686 860 -651 894
rect -617 860 -582 894
rect -548 860 -513 894
rect -479 860 -444 894
rect -410 860 -375 894
rect -2859 826 -375 860
rect -2825 792 -2790 826
rect -2756 792 -2721 826
rect -2687 792 -2652 826
rect -2618 792 -2583 826
rect -2549 792 -2514 826
rect -2480 792 -2445 826
rect -2411 792 -2376 826
rect -2342 792 -2307 826
rect -2273 792 -2238 826
rect -2204 792 -2169 826
rect -2135 792 -2100 826
rect -2066 792 -2031 826
rect -1997 792 -1962 826
rect -1928 792 -1893 826
rect -1859 792 -1824 826
rect -1790 792 -1755 826
rect -1721 792 -1686 826
rect -1652 792 -1617 826
rect -1583 792 -1548 826
rect -1514 792 -1479 826
rect -1445 792 -1410 826
rect -1376 792 -1341 826
rect -1307 792 -1272 826
rect -1238 792 -1203 826
rect -1169 792 -1134 826
rect -1100 792 -1065 826
rect -1031 792 -996 826
rect -962 792 -927 826
rect -893 792 -858 826
rect -824 792 -789 826
rect -755 792 -720 826
rect -686 792 -651 826
rect -617 792 -582 826
rect -548 792 -513 826
rect -479 792 -444 826
rect -410 792 -375 826
rect -1 792 2 1846
rect -2859 768 2 792
<< nsubdiff >>
rect -148 4232 2 4464
rect -148 3230 -101 4232
<< mvpsubdiff >>
rect 11949 4324 17215 4361
rect 11983 4290 12018 4324
rect 12052 4290 12087 4324
rect 12121 4290 12156 4324
rect 12190 4290 12225 4324
rect 12259 4290 12294 4324
rect 12328 4290 12363 4324
rect 12397 4290 12432 4324
rect 12466 4290 12501 4324
rect 12535 4290 12570 4324
rect 12604 4290 12639 4324
rect 12673 4290 12708 4324
rect 12742 4290 12777 4324
rect 12811 4290 12846 4324
rect 12880 4290 12915 4324
rect 12949 4290 12984 4324
rect 13018 4290 13053 4324
rect 13087 4290 13122 4324
rect 13156 4290 13191 4324
rect 13225 4290 13260 4324
rect 13294 4290 13329 4324
rect 13363 4290 13398 4324
rect 13432 4290 13467 4324
rect 13501 4290 13536 4324
rect 13570 4290 13605 4324
rect 13639 4290 13674 4324
rect 13708 4290 13743 4324
rect 13777 4290 13812 4324
rect 13846 4290 13881 4324
rect 13915 4290 13950 4324
rect 13984 4290 14019 4324
rect 14053 4290 14088 4324
rect 14122 4290 14157 4324
rect 14191 4290 14226 4324
rect 14260 4290 14295 4324
rect 14329 4290 14364 4324
rect 14398 4290 14433 4324
rect 14467 4290 14502 4324
rect 14536 4290 14571 4324
rect 14605 4290 14640 4324
rect 14674 4290 14709 4324
rect 14743 4290 14778 4324
rect 14812 4290 14847 4324
rect 14881 4290 14916 4324
rect 14950 4290 14985 4324
rect 15019 4290 15054 4324
rect 15088 4290 15123 4324
rect 15157 4290 15192 4324
rect 15226 4290 15261 4324
rect 15295 4290 15330 4324
rect 15364 4290 15399 4324
rect 15433 4290 15468 4324
rect 15502 4290 15537 4324
rect 15571 4290 15606 4324
rect 15640 4290 15675 4324
rect 15709 4290 15744 4324
rect 15778 4290 15813 4324
rect 15847 4290 15882 4324
rect 15916 4290 15951 4324
rect 15985 4290 16020 4324
rect 16054 4290 16089 4324
rect 16123 4290 16158 4324
rect 16192 4290 16227 4324
rect 16261 4290 16296 4324
rect 16330 4290 16365 4324
rect 11949 4256 16365 4290
rect 11983 4222 12018 4256
rect 12052 4222 12087 4256
rect 12121 4222 12156 4256
rect 12190 4222 12225 4256
rect 12259 4222 12294 4256
rect 12328 4222 12363 4256
rect 12397 4222 12432 4256
rect 12466 4222 12501 4256
rect 12535 4222 12570 4256
rect 12604 4222 12639 4256
rect 12673 4222 12708 4256
rect 12742 4222 12777 4256
rect 12811 4222 12846 4256
rect 12880 4222 12915 4256
rect 12949 4222 12984 4256
rect 13018 4222 13053 4256
rect 13087 4222 13122 4256
rect 13156 4222 13191 4256
rect 13225 4222 13260 4256
rect 13294 4222 13329 4256
rect 13363 4222 13398 4256
rect 13432 4222 13467 4256
rect 13501 4222 13536 4256
rect 13570 4222 13605 4256
rect 13639 4222 13674 4256
rect 13708 4222 13743 4256
rect 13777 4222 13812 4256
rect 13846 4222 13881 4256
rect 13915 4222 13950 4256
rect 13984 4222 14019 4256
rect 14053 4222 14088 4256
rect 14122 4222 14157 4256
rect 14191 4222 14226 4256
rect 14260 4222 14295 4256
rect 14329 4222 14364 4256
rect 14398 4222 14433 4256
rect 14467 4222 14502 4256
rect 14536 4222 14571 4256
rect 14605 4222 14640 4256
rect 14674 4222 14709 4256
rect 14743 4222 14778 4256
rect 14812 4222 14847 4256
rect 14881 4222 14916 4256
rect 14950 4222 14985 4256
rect 15019 4222 15054 4256
rect 15088 4222 15123 4256
rect 15157 4222 15192 4256
rect 15226 4222 15261 4256
rect 15295 4222 15330 4256
rect 15364 4222 15399 4256
rect 15433 4222 15468 4256
rect 15502 4222 15537 4256
rect 15571 4222 15606 4256
rect 15640 4222 15675 4256
rect 15709 4222 15744 4256
rect 15778 4222 15813 4256
rect 15847 4222 15882 4256
rect 15916 4222 15951 4256
rect 15985 4222 16020 4256
rect 16054 4222 16089 4256
rect 16123 4222 16158 4256
rect 16192 4222 16227 4256
rect 16261 4222 16296 4256
rect 16330 4222 16365 4256
rect 11949 4188 16365 4222
rect 11983 4154 12018 4188
rect 12052 4154 12087 4188
rect 12121 4154 12156 4188
rect 12190 4154 12225 4188
rect 12259 4154 12294 4188
rect 12328 4154 12363 4188
rect 12397 4154 12432 4188
rect 12466 4154 12501 4188
rect 12535 4154 12570 4188
rect 12604 4154 12639 4188
rect 12673 4154 12708 4188
rect 12742 4154 12777 4188
rect 12811 4154 12846 4188
rect 12880 4154 12915 4188
rect 12949 4154 12984 4188
rect 13018 4154 13053 4188
rect 13087 4154 13122 4188
rect 13156 4154 13191 4188
rect 13225 4154 13260 4188
rect 13294 4154 13329 4188
rect 13363 4154 13398 4188
rect 13432 4154 13467 4188
rect 13501 4154 13536 4188
rect 13570 4154 13605 4188
rect 13639 4154 13674 4188
rect 13708 4154 13743 4188
rect 13777 4154 13812 4188
rect 13846 4154 13881 4188
rect 13915 4154 13950 4188
rect 13984 4154 14019 4188
rect 14053 4154 14088 4188
rect 14122 4154 14157 4188
rect 14191 4154 14226 4188
rect 14260 4154 14295 4188
rect 14329 4154 14364 4188
rect 14398 4154 14433 4188
rect 14467 4154 14502 4188
rect 14536 4154 14571 4188
rect 14605 4154 14640 4188
rect 14674 4154 14709 4188
rect 14743 4154 14778 4188
rect 14812 4154 14847 4188
rect 14881 4154 14916 4188
rect 14950 4154 14985 4188
rect 15019 4154 15054 4188
rect 15088 4154 15123 4188
rect 15157 4154 15192 4188
rect 15226 4154 15261 4188
rect 15295 4154 15330 4188
rect 15364 4154 15399 4188
rect 15433 4154 15468 4188
rect 15502 4154 15537 4188
rect 15571 4154 15606 4188
rect 15640 4154 15675 4188
rect 15709 4154 15744 4188
rect 15778 4154 15813 4188
rect 15847 4154 15882 4188
rect 15916 4154 15951 4188
rect 15985 4154 16020 4188
rect 16054 4154 16089 4188
rect 16123 4154 16158 4188
rect 16192 4154 16227 4188
rect 16261 4154 16296 4188
rect 16330 4154 16365 4188
rect 11949 4120 16365 4154
rect 11983 4086 12018 4120
rect 12052 4086 12087 4120
rect 12121 4086 12156 4120
rect 12190 4086 12225 4120
rect 12259 4086 12294 4120
rect 12328 4086 12363 4120
rect 12397 4086 12432 4120
rect 12466 4086 12501 4120
rect 12535 4086 12570 4120
rect 12604 4086 12639 4120
rect 12673 4086 12708 4120
rect 12742 4086 12777 4120
rect 12811 4086 12846 4120
rect 12880 4086 12915 4120
rect 12949 4086 12984 4120
rect 13018 4086 13053 4120
rect 13087 4086 13122 4120
rect 13156 4086 13191 4120
rect 13225 4086 13260 4120
rect 13294 4086 13329 4120
rect 13363 4086 13398 4120
rect 13432 4086 13467 4120
rect 13501 4086 13536 4120
rect 13570 4086 13605 4120
rect 13639 4086 13674 4120
rect 13708 4086 13743 4120
rect 13777 4086 13812 4120
rect 13846 4086 13881 4120
rect 13915 4086 13950 4120
rect 13984 4086 14019 4120
rect 14053 4086 14088 4120
rect 14122 4086 14157 4120
rect 14191 4086 14226 4120
rect 14260 4086 14295 4120
rect 14329 4086 14364 4120
rect 14398 4086 14433 4120
rect 14467 4086 14502 4120
rect 14536 4086 14571 4120
rect 14605 4086 14640 4120
rect 14674 4086 14709 4120
rect 14743 4086 14778 4120
rect 14812 4086 14847 4120
rect 14881 4086 14916 4120
rect 14950 4086 14985 4120
rect 15019 4086 15054 4120
rect 15088 4086 15123 4120
rect 15157 4086 15192 4120
rect 15226 4086 15261 4120
rect 15295 4086 15330 4120
rect 15364 4086 15399 4120
rect 15433 4086 15468 4120
rect 15502 4086 15537 4120
rect 15571 4086 15606 4120
rect 15640 4086 15675 4120
rect 15709 4086 15744 4120
rect 15778 4086 15813 4120
rect 15847 4086 15882 4120
rect 15916 4086 15951 4120
rect 15985 4086 16020 4120
rect 16054 4086 16089 4120
rect 16123 4086 16158 4120
rect 16192 4086 16227 4120
rect 16261 4086 16296 4120
rect 16330 4086 16365 4120
rect 11949 4052 16365 4086
rect 11983 4018 12018 4052
rect 12052 4018 12087 4052
rect 12121 4018 12156 4052
rect 12190 4018 12225 4052
rect 12259 4018 12294 4052
rect 12328 4018 12363 4052
rect 12397 4018 12432 4052
rect 12466 4018 12501 4052
rect 12535 4018 12570 4052
rect 12604 4018 12639 4052
rect 12673 4018 12708 4052
rect 12742 4018 12777 4052
rect 12811 4018 12846 4052
rect 12880 4018 12915 4052
rect 12949 4018 12984 4052
rect 13018 4018 13053 4052
rect 13087 4018 13122 4052
rect 13156 4018 13191 4052
rect 13225 4018 13260 4052
rect 13294 4018 13329 4052
rect 13363 4018 13398 4052
rect 13432 4018 13467 4052
rect 13501 4018 13536 4052
rect 13570 4018 13605 4052
rect 13639 4018 13674 4052
rect 13708 4018 13743 4052
rect 13777 4018 13812 4052
rect 13846 4018 13881 4052
rect 13915 4018 13950 4052
rect 13984 4018 14019 4052
rect 14053 4018 14088 4052
rect 14122 4018 14157 4052
rect 14191 4018 14226 4052
rect 14260 4018 14295 4052
rect 14329 4018 14364 4052
rect 14398 4018 14433 4052
rect 14467 4018 14502 4052
rect 14536 4018 14571 4052
rect 14605 4018 14640 4052
rect 14674 4018 14709 4052
rect 14743 4018 14778 4052
rect 14812 4018 14847 4052
rect 14881 4018 14916 4052
rect 14950 4018 14985 4052
rect 15019 4018 15054 4052
rect 15088 4018 15123 4052
rect 15157 4018 15192 4052
rect 15226 4018 15261 4052
rect 15295 4018 15330 4052
rect 15364 4018 15399 4052
rect 15433 4018 15468 4052
rect 15502 4018 15537 4052
rect 15571 4018 15606 4052
rect 15640 4018 15675 4052
rect 15709 4018 15744 4052
rect 15778 4018 15813 4052
rect 15847 4018 15882 4052
rect 15916 4018 15951 4052
rect 15985 4018 16020 4052
rect 16054 4018 16089 4052
rect 16123 4018 16158 4052
rect 16192 4018 16227 4052
rect 16261 4018 16296 4052
rect 16330 4018 16365 4052
rect 11949 3984 16365 4018
rect 11983 3950 12018 3984
rect 12052 3950 12087 3984
rect 12121 3950 12156 3984
rect 12190 3950 12225 3984
rect 12259 3950 12294 3984
rect 12328 3950 12363 3984
rect 12397 3950 12432 3984
rect 12466 3950 12501 3984
rect 12535 3950 12570 3984
rect 12604 3950 12639 3984
rect 12673 3950 12708 3984
rect 12742 3950 12777 3984
rect 12811 3950 12846 3984
rect 12880 3950 12915 3984
rect 12949 3950 12984 3984
rect 13018 3950 13053 3984
rect 13087 3950 13122 3984
rect 13156 3950 13191 3984
rect 13225 3950 13260 3984
rect 13294 3950 13329 3984
rect 13363 3950 13398 3984
rect 13432 3950 13467 3984
rect 13501 3950 13536 3984
rect 13570 3950 13605 3984
rect 13639 3950 13674 3984
rect 13708 3950 13743 3984
rect 13777 3950 13812 3984
rect 13846 3950 13881 3984
rect 13915 3950 13950 3984
rect 13984 3950 14019 3984
rect 14053 3950 14088 3984
rect 14122 3950 14157 3984
rect 14191 3950 14226 3984
rect 14260 3950 14295 3984
rect 14329 3950 14364 3984
rect 14398 3950 14433 3984
rect 14467 3950 14502 3984
rect 14536 3950 14571 3984
rect 14605 3950 14640 3984
rect 14674 3950 14709 3984
rect 14743 3950 14778 3984
rect 14812 3950 14847 3984
rect 14881 3950 14916 3984
rect 14950 3950 14985 3984
rect 15019 3950 15054 3984
rect 15088 3950 15123 3984
rect 15157 3950 15192 3984
rect 15226 3950 15261 3984
rect 15295 3950 15330 3984
rect 15364 3950 15399 3984
rect 15433 3950 15468 3984
rect 15502 3950 15537 3984
rect 15571 3950 15606 3984
rect 15640 3950 15675 3984
rect 15709 3950 15744 3984
rect 15778 3950 15813 3984
rect 15847 3950 15882 3984
rect 15916 3950 15951 3984
rect 15985 3950 16020 3984
rect 16054 3950 16089 3984
rect 16123 3950 16158 3984
rect 16192 3950 16227 3984
rect 16261 3950 16296 3984
rect 16330 3950 16365 3984
rect 11949 3916 16365 3950
rect 11983 3882 12018 3916
rect 12052 3882 12087 3916
rect 12121 3882 12156 3916
rect 12190 3882 12225 3916
rect 12259 3882 12294 3916
rect 12328 3882 12363 3916
rect 12397 3882 12432 3916
rect 12466 3882 12501 3916
rect 12535 3882 12570 3916
rect 12604 3882 12639 3916
rect 12673 3882 12708 3916
rect 12742 3882 12777 3916
rect 12811 3882 12846 3916
rect 12880 3882 12915 3916
rect 12949 3882 12984 3916
rect 13018 3882 13053 3916
rect 13087 3882 13122 3916
rect 13156 3882 13191 3916
rect 13225 3882 13260 3916
rect 13294 3882 13329 3916
rect 13363 3882 13398 3916
rect 13432 3882 13467 3916
rect 13501 3882 13536 3916
rect 13570 3882 13605 3916
rect 13639 3882 13674 3916
rect 13708 3882 13743 3916
rect 13777 3882 13812 3916
rect 13846 3882 13881 3916
rect 13915 3882 13950 3916
rect 13984 3882 14019 3916
rect 14053 3882 14088 3916
rect 14122 3882 14157 3916
rect 14191 3882 14226 3916
rect 14260 3882 14295 3916
rect 14329 3882 14364 3916
rect 14398 3882 14433 3916
rect 14467 3882 14502 3916
rect 14536 3882 14571 3916
rect 14605 3882 14640 3916
rect 14674 3882 14709 3916
rect 14743 3882 14778 3916
rect 14812 3882 14847 3916
rect 14881 3882 14916 3916
rect 14950 3882 14985 3916
rect 15019 3882 15054 3916
rect 15088 3882 15123 3916
rect 15157 3882 15192 3916
rect 15226 3882 15261 3916
rect 15295 3882 15330 3916
rect 15364 3882 15399 3916
rect 15433 3882 15468 3916
rect 15502 3882 15537 3916
rect 15571 3882 15606 3916
rect 15640 3882 15675 3916
rect 15709 3882 15744 3916
rect 15778 3882 15813 3916
rect 15847 3882 15882 3916
rect 15916 3882 15951 3916
rect 15985 3882 16020 3916
rect 16054 3882 16089 3916
rect 16123 3882 16158 3916
rect 16192 3882 16227 3916
rect 16261 3882 16296 3916
rect 16330 3882 16365 3916
rect 11949 3848 16365 3882
rect 11983 3814 12018 3848
rect 12052 3814 12087 3848
rect 12121 3814 12156 3848
rect 12190 3814 12225 3848
rect 12259 3814 12294 3848
rect 12328 3814 12363 3848
rect 12397 3814 12432 3848
rect 12466 3814 12501 3848
rect 12535 3814 12570 3848
rect 12604 3814 12639 3848
rect 12673 3814 12708 3848
rect 12742 3814 12777 3848
rect 12811 3814 12846 3848
rect 12880 3814 12915 3848
rect 12949 3814 12984 3848
rect 13018 3814 13053 3848
rect 13087 3814 13122 3848
rect 13156 3814 13191 3848
rect 13225 3814 13260 3848
rect 13294 3814 13329 3848
rect 13363 3814 13398 3848
rect 13432 3814 13467 3848
rect 13501 3814 13536 3848
rect 13570 3814 13605 3848
rect 13639 3814 13674 3848
rect 13708 3814 13743 3848
rect 13777 3814 13812 3848
rect 13846 3814 13881 3848
rect 13915 3814 13950 3848
rect 13984 3814 14019 3848
rect 14053 3814 14088 3848
rect 14122 3814 14157 3848
rect 14191 3814 14226 3848
rect 14260 3814 14295 3848
rect 14329 3814 14364 3848
rect 14398 3814 14433 3848
rect 14467 3814 14502 3848
rect 14536 3814 14571 3848
rect 14605 3814 14640 3848
rect 14674 3814 14709 3848
rect 14743 3814 14778 3848
rect 14812 3814 14847 3848
rect 14881 3814 14916 3848
rect 14950 3814 14985 3848
rect 15019 3814 15054 3848
rect 15088 3814 15123 3848
rect 15157 3814 15192 3848
rect 15226 3814 15261 3848
rect 15295 3814 15330 3848
rect 15364 3814 15399 3848
rect 15433 3814 15468 3848
rect 15502 3814 15537 3848
rect 15571 3814 15606 3848
rect 15640 3814 15675 3848
rect 15709 3814 15744 3848
rect 15778 3814 15813 3848
rect 15847 3814 15882 3848
rect 15916 3814 15951 3848
rect 15985 3814 16020 3848
rect 16054 3814 16089 3848
rect 16123 3814 16158 3848
rect 16192 3814 16227 3848
rect 16261 3814 16296 3848
rect 16330 3814 16365 3848
rect 11949 3780 16365 3814
rect 11983 3746 12018 3780
rect 12052 3746 12087 3780
rect 12121 3746 12156 3780
rect 12190 3746 12225 3780
rect 12259 3746 12294 3780
rect 12328 3746 12363 3780
rect 12397 3746 12432 3780
rect 12466 3746 12501 3780
rect 12535 3746 12570 3780
rect 12604 3746 12639 3780
rect 12673 3746 12708 3780
rect 12742 3746 12777 3780
rect 12811 3746 12846 3780
rect 12880 3746 12915 3780
rect 12949 3746 12984 3780
rect 13018 3746 13053 3780
rect 13087 3746 13122 3780
rect 13156 3746 13191 3780
rect 13225 3746 13260 3780
rect 13294 3746 13329 3780
rect 13363 3746 13398 3780
rect 13432 3746 13467 3780
rect 13501 3746 13536 3780
rect 13570 3746 13605 3780
rect 13639 3746 13674 3780
rect 13708 3746 13743 3780
rect 13777 3746 13812 3780
rect 13846 3746 13881 3780
rect 13915 3746 13950 3780
rect 13984 3746 14019 3780
rect 14053 3746 14088 3780
rect 14122 3746 14157 3780
rect 14191 3746 14226 3780
rect 14260 3746 14295 3780
rect 14329 3746 14364 3780
rect 14398 3746 14433 3780
rect 14467 3746 14502 3780
rect 14536 3746 14571 3780
rect 14605 3746 14640 3780
rect 14674 3746 14709 3780
rect 14743 3746 14778 3780
rect 14812 3746 14847 3780
rect 14881 3746 14916 3780
rect 14950 3746 14985 3780
rect 15019 3746 15054 3780
rect 15088 3746 15123 3780
rect 15157 3746 15192 3780
rect 15226 3746 15261 3780
rect 15295 3746 15330 3780
rect 15364 3746 15399 3780
rect 15433 3746 15468 3780
rect 15502 3746 15537 3780
rect 15571 3746 15606 3780
rect 15640 3746 15675 3780
rect 15709 3746 15744 3780
rect 15778 3746 15813 3780
rect 15847 3746 15882 3780
rect 15916 3746 15951 3780
rect 15985 3746 16020 3780
rect 16054 3746 16089 3780
rect 16123 3746 16158 3780
rect 16192 3746 16227 3780
rect 16261 3746 16296 3780
rect 16330 3746 16365 3780
rect 11949 3712 16365 3746
rect 11983 3678 12018 3712
rect 12052 3678 12087 3712
rect 12121 3678 12156 3712
rect 12190 3678 12225 3712
rect 12259 3678 12294 3712
rect 12328 3678 12363 3712
rect 12397 3678 12432 3712
rect 12466 3678 12501 3712
rect 12535 3678 12570 3712
rect 12604 3678 12639 3712
rect 12673 3678 12708 3712
rect 12742 3678 12777 3712
rect 12811 3678 12846 3712
rect 12880 3678 12915 3712
rect 12949 3678 12984 3712
rect 13018 3678 13053 3712
rect 13087 3678 13122 3712
rect 13156 3678 13191 3712
rect 13225 3678 13260 3712
rect 13294 3678 13329 3712
rect 13363 3678 13398 3712
rect 13432 3678 13467 3712
rect 13501 3678 13536 3712
rect 13570 3678 13605 3712
rect 13639 3678 13674 3712
rect 13708 3678 13743 3712
rect 13777 3678 13812 3712
rect 13846 3678 13881 3712
rect 13915 3678 13950 3712
rect 13984 3678 14019 3712
rect 14053 3678 14088 3712
rect 14122 3678 14157 3712
rect 14191 3678 14226 3712
rect 14260 3678 14295 3712
rect 14329 3678 14364 3712
rect 14398 3678 14433 3712
rect 14467 3678 14502 3712
rect 14536 3678 14571 3712
rect 14605 3678 14640 3712
rect 14674 3678 14709 3712
rect 14743 3678 14778 3712
rect 14812 3678 14847 3712
rect 14881 3678 14916 3712
rect 14950 3678 14985 3712
rect 15019 3678 15054 3712
rect 15088 3678 15123 3712
rect 15157 3678 15192 3712
rect 15226 3678 15261 3712
rect 15295 3678 15330 3712
rect 15364 3678 15399 3712
rect 15433 3678 15468 3712
rect 15502 3678 15537 3712
rect 15571 3678 15606 3712
rect 15640 3678 15675 3712
rect 15709 3678 15744 3712
rect 15778 3678 15813 3712
rect 15847 3678 15882 3712
rect 15916 3678 15951 3712
rect 15985 3678 16020 3712
rect 16054 3678 16089 3712
rect 16123 3678 16158 3712
rect 16192 3678 16227 3712
rect 16261 3678 16296 3712
rect 16330 3678 16365 3712
rect 11949 3644 16365 3678
rect 11983 3610 12018 3644
rect 12052 3610 12087 3644
rect 12121 3610 12156 3644
rect 12190 3610 12225 3644
rect 12259 3610 12294 3644
rect 12328 3610 12363 3644
rect 12397 3610 12432 3644
rect 12466 3610 12501 3644
rect 12535 3610 12570 3644
rect 12604 3610 12639 3644
rect 12673 3610 12708 3644
rect 12742 3610 12777 3644
rect 12811 3610 12846 3644
rect 12880 3610 12915 3644
rect 12949 3610 12984 3644
rect 13018 3610 13053 3644
rect 13087 3610 13122 3644
rect 13156 3610 13191 3644
rect 13225 3610 13260 3644
rect 13294 3610 13329 3644
rect 13363 3610 13398 3644
rect 13432 3610 13467 3644
rect 13501 3610 13536 3644
rect 13570 3610 13605 3644
rect 13639 3610 13674 3644
rect 13708 3610 13743 3644
rect 13777 3610 13812 3644
rect 13846 3610 13881 3644
rect 13915 3610 13950 3644
rect 13984 3610 14019 3644
rect 14053 3610 14088 3644
rect 14122 3610 14157 3644
rect 14191 3610 14226 3644
rect 14260 3610 14295 3644
rect 14329 3610 14364 3644
rect 14398 3610 14433 3644
rect 14467 3610 14502 3644
rect 14536 3610 14571 3644
rect 14605 3610 14640 3644
rect 14674 3610 14709 3644
rect 14743 3610 14778 3644
rect 14812 3610 14847 3644
rect 14881 3610 14916 3644
rect 14950 3610 14985 3644
rect 15019 3610 15054 3644
rect 15088 3610 15123 3644
rect 15157 3610 15192 3644
rect 15226 3610 15261 3644
rect 15295 3610 15330 3644
rect 15364 3610 15399 3644
rect 15433 3610 15468 3644
rect 15502 3610 15537 3644
rect 15571 3610 15606 3644
rect 15640 3610 15675 3644
rect 15709 3610 15744 3644
rect 15778 3610 15813 3644
rect 15847 3610 15882 3644
rect 15916 3610 15951 3644
rect 15985 3610 16020 3644
rect 16054 3610 16089 3644
rect 16123 3610 16158 3644
rect 16192 3610 16227 3644
rect 16261 3610 16296 3644
rect 16330 3610 16365 3644
rect 11949 3576 16365 3610
rect 11983 3542 12018 3576
rect 12052 3542 12087 3576
rect 12121 3542 12156 3576
rect 12190 3542 12225 3576
rect 12259 3542 12294 3576
rect 12328 3542 12363 3576
rect 12397 3542 12432 3576
rect 12466 3542 12501 3576
rect 12535 3542 12570 3576
rect 12604 3542 12639 3576
rect 12673 3542 12708 3576
rect 12742 3542 12777 3576
rect 12811 3542 12846 3576
rect 12880 3542 12915 3576
rect 12949 3542 12984 3576
rect 13018 3542 13053 3576
rect 13087 3542 13122 3576
rect 13156 3542 13191 3576
rect 13225 3542 13260 3576
rect 13294 3542 13329 3576
rect 13363 3542 13398 3576
rect 13432 3542 13467 3576
rect 13501 3542 13536 3576
rect 13570 3542 13605 3576
rect 13639 3542 13674 3576
rect 13708 3542 13743 3576
rect 13777 3542 13812 3576
rect 13846 3542 13881 3576
rect 13915 3542 13950 3576
rect 13984 3542 14019 3576
rect 14053 3542 14088 3576
rect 14122 3542 14157 3576
rect 14191 3542 14226 3576
rect 14260 3542 14295 3576
rect 14329 3542 14364 3576
rect 14398 3542 14433 3576
rect 14467 3542 14502 3576
rect 14536 3542 14571 3576
rect 14605 3542 14640 3576
rect 14674 3542 14709 3576
rect 14743 3542 14778 3576
rect 14812 3542 14847 3576
rect 14881 3542 14916 3576
rect 14950 3542 14985 3576
rect 15019 3542 15054 3576
rect 15088 3542 15123 3576
rect 15157 3542 15192 3576
rect 15226 3542 15261 3576
rect 15295 3542 15330 3576
rect 15364 3542 15399 3576
rect 15433 3542 15468 3576
rect 15502 3542 15537 3576
rect 15571 3542 15606 3576
rect 15640 3542 15675 3576
rect 15709 3542 15744 3576
rect 15778 3542 15813 3576
rect 15847 3542 15882 3576
rect 15916 3542 15951 3576
rect 15985 3542 16020 3576
rect 16054 3542 16089 3576
rect 16123 3542 16158 3576
rect 16192 3542 16227 3576
rect 16261 3542 16296 3576
rect 16330 3542 16365 3576
rect 11949 3508 16365 3542
rect 11983 3474 12018 3508
rect 12052 3474 12087 3508
rect 12121 3474 12156 3508
rect 12190 3474 12225 3508
rect 12259 3474 12294 3508
rect 12328 3474 12363 3508
rect 12397 3474 12432 3508
rect 12466 3474 12501 3508
rect 12535 3474 12570 3508
rect 12604 3474 12639 3508
rect 12673 3474 12708 3508
rect 12742 3474 12777 3508
rect 12811 3474 12846 3508
rect 12880 3474 12915 3508
rect 12949 3474 12984 3508
rect 13018 3474 13053 3508
rect 13087 3474 13122 3508
rect 13156 3474 13191 3508
rect 13225 3474 13260 3508
rect 13294 3474 13329 3508
rect 13363 3474 13398 3508
rect 13432 3474 13467 3508
rect 13501 3474 13536 3508
rect 13570 3474 13605 3508
rect 13639 3474 13674 3508
rect 13708 3474 13743 3508
rect 13777 3474 13812 3508
rect 13846 3474 13881 3508
rect 13915 3474 13950 3508
rect 13984 3474 14019 3508
rect 14053 3474 14088 3508
rect 14122 3474 14157 3508
rect 14191 3474 14226 3508
rect 14260 3474 14295 3508
rect 14329 3474 14364 3508
rect 14398 3474 14433 3508
rect 14467 3474 14502 3508
rect 14536 3474 14571 3508
rect 14605 3474 14640 3508
rect 14674 3474 14709 3508
rect 14743 3474 14778 3508
rect 14812 3474 14847 3508
rect 14881 3474 14916 3508
rect 14950 3474 14985 3508
rect 15019 3474 15054 3508
rect 15088 3474 15123 3508
rect 15157 3474 15192 3508
rect 15226 3474 15261 3508
rect 15295 3474 15330 3508
rect 15364 3474 15399 3508
rect 15433 3474 15468 3508
rect 15502 3474 15537 3508
rect 15571 3474 15606 3508
rect 15640 3474 15675 3508
rect 15709 3474 15744 3508
rect 15778 3474 15813 3508
rect 15847 3474 15882 3508
rect 15916 3474 15951 3508
rect 15985 3474 16020 3508
rect 16054 3474 16089 3508
rect 16123 3474 16158 3508
rect 16192 3474 16227 3508
rect 16261 3474 16296 3508
rect 16330 3474 16365 3508
rect 11949 3440 16365 3474
rect 11983 3406 12018 3440
rect 12052 3406 12087 3440
rect 12121 3406 12156 3440
rect 12190 3406 12225 3440
rect 12259 3406 12294 3440
rect 12328 3406 12363 3440
rect 12397 3406 12432 3440
rect 12466 3406 12501 3440
rect 12535 3406 12570 3440
rect 12604 3406 12639 3440
rect 12673 3406 12708 3440
rect 12742 3406 12777 3440
rect 12811 3406 12846 3440
rect 12880 3406 12915 3440
rect 12949 3406 12984 3440
rect 13018 3406 13053 3440
rect 13087 3406 13122 3440
rect 13156 3406 13191 3440
rect 13225 3406 13260 3440
rect 13294 3406 13329 3440
rect 13363 3406 13398 3440
rect 13432 3406 13467 3440
rect 13501 3406 13536 3440
rect 13570 3406 13605 3440
rect 13639 3406 13674 3440
rect 13708 3406 13743 3440
rect 13777 3406 13812 3440
rect 13846 3406 13881 3440
rect 13915 3406 13950 3440
rect 13984 3406 14019 3440
rect 14053 3406 14088 3440
rect 14122 3406 14157 3440
rect 14191 3406 14226 3440
rect 14260 3406 14295 3440
rect 14329 3406 14364 3440
rect 14398 3406 14433 3440
rect 14467 3406 14502 3440
rect 14536 3406 14571 3440
rect 14605 3406 14640 3440
rect 14674 3406 14709 3440
rect 14743 3406 14778 3440
rect 14812 3406 14847 3440
rect 14881 3406 14916 3440
rect 14950 3406 14985 3440
rect 15019 3406 15054 3440
rect 15088 3406 15123 3440
rect 15157 3406 15192 3440
rect 15226 3406 15261 3440
rect 15295 3406 15330 3440
rect 15364 3406 15399 3440
rect 15433 3406 15468 3440
rect 15502 3406 15537 3440
rect 15571 3406 15606 3440
rect 15640 3406 15675 3440
rect 15709 3406 15744 3440
rect 15778 3406 15813 3440
rect 15847 3406 15882 3440
rect 15916 3406 15951 3440
rect 15985 3406 16020 3440
rect 16054 3406 16089 3440
rect 16123 3406 16158 3440
rect 16192 3406 16227 3440
rect 16261 3406 16296 3440
rect 16330 3406 16365 3440
rect 11949 3372 16365 3406
rect 11983 3338 12018 3372
rect 12052 3338 12087 3372
rect 12121 3338 12156 3372
rect 12190 3338 12225 3372
rect 12259 3338 12294 3372
rect 12328 3338 12363 3372
rect 12397 3338 12432 3372
rect 12466 3338 12501 3372
rect 12535 3338 12570 3372
rect 12604 3338 12639 3372
rect 12673 3338 12708 3372
rect 12742 3338 12777 3372
rect 12811 3338 12846 3372
rect 12880 3338 12915 3372
rect 12949 3338 12984 3372
rect 13018 3338 13053 3372
rect 13087 3338 13122 3372
rect 13156 3338 13191 3372
rect 13225 3338 13260 3372
rect 13294 3338 13329 3372
rect 13363 3338 13398 3372
rect 13432 3338 13467 3372
rect 13501 3338 13536 3372
rect 13570 3338 13605 3372
rect 13639 3338 13674 3372
rect 13708 3338 13743 3372
rect 13777 3338 13812 3372
rect 13846 3338 13881 3372
rect 13915 3338 13950 3372
rect 13984 3338 14019 3372
rect 14053 3338 14088 3372
rect 14122 3338 14157 3372
rect 14191 3338 14226 3372
rect 14260 3338 14295 3372
rect 14329 3338 14364 3372
rect 14398 3338 14433 3372
rect 14467 3338 14502 3372
rect 14536 3338 14571 3372
rect 14605 3338 14640 3372
rect 14674 3338 14709 3372
rect 14743 3338 14778 3372
rect 14812 3338 14847 3372
rect 14881 3338 14916 3372
rect 14950 3338 14985 3372
rect 15019 3338 15054 3372
rect 15088 3338 15123 3372
rect 15157 3338 15192 3372
rect 15226 3338 15261 3372
rect 15295 3338 15330 3372
rect 15364 3338 15399 3372
rect 15433 3338 15468 3372
rect 15502 3338 15537 3372
rect 15571 3338 15606 3372
rect 15640 3338 15675 3372
rect 15709 3338 15744 3372
rect 15778 3338 15813 3372
rect 15847 3338 15882 3372
rect 15916 3338 15951 3372
rect 15985 3338 16020 3372
rect 16054 3338 16089 3372
rect 16123 3338 16158 3372
rect 16192 3338 16227 3372
rect 16261 3338 16296 3372
rect 16330 3338 16365 3372
rect 11949 3304 16365 3338
rect 11983 3270 12018 3304
rect 12052 3270 12087 3304
rect 12121 3270 12156 3304
rect 12190 3270 12225 3304
rect 12259 3270 12294 3304
rect 12328 3270 12363 3304
rect 12397 3270 12432 3304
rect 12466 3270 12501 3304
rect 12535 3270 12570 3304
rect 12604 3270 12639 3304
rect 12673 3270 12708 3304
rect 12742 3270 12777 3304
rect 12811 3270 12846 3304
rect 12880 3270 12915 3304
rect 12949 3270 12984 3304
rect 13018 3270 13053 3304
rect 13087 3270 13122 3304
rect 13156 3270 13191 3304
rect 13225 3270 13260 3304
rect 13294 3270 13329 3304
rect 13363 3270 13398 3304
rect 13432 3270 13467 3304
rect 13501 3270 13536 3304
rect 13570 3270 13605 3304
rect 13639 3270 13674 3304
rect 13708 3270 13743 3304
rect 13777 3270 13812 3304
rect 13846 3270 13881 3304
rect 13915 3270 13950 3304
rect 13984 3270 14019 3304
rect 14053 3270 14088 3304
rect 14122 3270 14157 3304
rect 14191 3270 14226 3304
rect 14260 3270 14295 3304
rect 14329 3270 14364 3304
rect 14398 3270 14433 3304
rect 14467 3270 14502 3304
rect 14536 3270 14571 3304
rect 14605 3270 14640 3304
rect 14674 3270 14709 3304
rect 14743 3270 14778 3304
rect 14812 3270 14847 3304
rect 14881 3270 14916 3304
rect 14950 3270 14985 3304
rect 15019 3270 15054 3304
rect 15088 3270 15123 3304
rect 15157 3270 15192 3304
rect 15226 3270 15261 3304
rect 15295 3270 15330 3304
rect 15364 3270 15399 3304
rect 15433 3270 15468 3304
rect 15502 3270 15537 3304
rect 15571 3270 15606 3304
rect 15640 3270 15675 3304
rect 15709 3270 15744 3304
rect 15778 3270 15813 3304
rect 15847 3270 15882 3304
rect 15916 3270 15951 3304
rect 15985 3270 16020 3304
rect 16054 3270 16089 3304
rect 16123 3270 16158 3304
rect 16192 3270 16227 3304
rect 16261 3270 16296 3304
rect 16330 3270 16365 3304
rect 11949 3240 17215 3270
rect 4615 3235 17215 3240
rect 4615 3201 4639 3235
rect 4673 3201 4708 3235
rect 4742 3201 4777 3235
rect 4811 3201 4846 3235
rect 4880 3201 4915 3235
rect 4949 3201 4984 3235
rect 5018 3201 5053 3235
rect 4615 3167 5053 3201
rect 4615 3133 4639 3167
rect 4673 3133 4708 3167
rect 4742 3133 4777 3167
rect 4811 3133 4846 3167
rect 4880 3133 4915 3167
rect 4949 3133 4984 3167
rect 5018 3133 5053 3167
rect 4615 3099 5053 3133
rect 4615 3065 4639 3099
rect 4673 3065 4708 3099
rect 4742 3065 4777 3099
rect 4811 3065 4846 3099
rect 4880 3065 4915 3099
rect 4949 3065 4984 3099
rect 5018 3065 5053 3099
rect 4615 3031 5053 3065
rect 4615 2997 4639 3031
rect 4673 2997 4708 3031
rect 4742 2997 4777 3031
rect 4811 2997 4846 3031
rect 4880 2997 4915 3031
rect 4949 2997 4984 3031
rect 5018 2997 5053 3031
rect 4615 2963 5053 2997
rect 4615 2929 4639 2963
rect 4673 2929 4708 2963
rect 4742 2929 4777 2963
rect 4811 2929 4846 2963
rect 4880 2929 4915 2963
rect 4949 2929 4984 2963
rect 5018 2929 5053 2963
rect 4615 2895 5053 2929
rect 4615 2861 4639 2895
rect 4673 2861 4708 2895
rect 4742 2861 4777 2895
rect 4811 2861 4846 2895
rect 4880 2861 4915 2895
rect 4949 2861 4984 2895
rect 5018 2861 5053 2895
rect 4615 2827 5053 2861
rect 4615 2793 4639 2827
rect 4673 2793 4708 2827
rect 4742 2793 4777 2827
rect 4811 2793 4846 2827
rect 4880 2793 4915 2827
rect 4949 2793 4984 2827
rect 5018 2793 5053 2827
rect 4615 2759 5053 2793
rect 4615 2725 4639 2759
rect 4673 2725 4708 2759
rect 4742 2725 4777 2759
rect 4811 2725 4846 2759
rect 4880 2725 4915 2759
rect 4949 2725 4984 2759
rect 5018 2725 5053 2759
rect 4615 2691 5053 2725
rect 4615 2657 4639 2691
rect 4673 2657 4708 2691
rect 4742 2657 4777 2691
rect 4811 2657 4846 2691
rect 4880 2657 4915 2691
rect 4949 2657 4984 2691
rect 5018 2657 5053 2691
rect 4615 2623 5053 2657
rect 4615 2589 4639 2623
rect 4673 2589 4708 2623
rect 4742 2589 4777 2623
rect 4811 2589 4846 2623
rect 4880 2589 4915 2623
rect 4949 2589 4984 2623
rect 5018 2589 5053 2623
rect 4615 2555 5053 2589
rect 4615 2521 4639 2555
rect 4673 2521 4708 2555
rect 4742 2521 4777 2555
rect 4811 2521 4846 2555
rect 4880 2521 4915 2555
rect 4949 2521 4984 2555
rect 5018 2521 5053 2555
rect 4615 2487 5053 2521
rect 4615 2453 4639 2487
rect 4673 2453 4708 2487
rect 4742 2453 4777 2487
rect 4811 2453 4846 2487
rect 4880 2453 4915 2487
rect 4949 2453 4984 2487
rect 5018 2453 5053 2487
rect 4615 2419 5053 2453
rect 4615 2385 4639 2419
rect 4673 2385 4708 2419
rect 4742 2385 4777 2419
rect 4811 2385 4846 2419
rect 4880 2385 4915 2419
rect 4949 2385 4984 2419
rect 5018 2385 5053 2419
rect 4615 2351 5053 2385
rect 4615 2317 4639 2351
rect 4673 2317 4708 2351
rect 4742 2317 4777 2351
rect 4811 2317 4846 2351
rect 4880 2317 4915 2351
rect 4949 2317 4984 2351
rect 5018 2317 5053 2351
rect 4615 2283 5053 2317
rect 4615 2249 4639 2283
rect 4673 2249 4708 2283
rect 4742 2249 4777 2283
rect 4811 2249 4846 2283
rect 4880 2249 4915 2283
rect 4949 2249 4984 2283
rect 5018 2249 5053 2283
rect 4615 2215 5053 2249
rect 4615 2181 4639 2215
rect 4673 2181 4708 2215
rect 4742 2181 4777 2215
rect 4811 2181 4846 2215
rect 4880 2181 4915 2215
rect 4949 2181 4984 2215
rect 5018 2181 5053 2215
rect 17191 2181 17215 3235
rect 4615 2175 15944 2181
rect 4615 2147 5716 2175
rect 4649 2113 4686 2147
rect 4720 2113 4757 2147
rect 4791 2113 4828 2147
rect 4862 2113 4899 2147
rect 4933 2113 4970 2147
rect 5004 2113 5041 2147
rect 5075 2113 5112 2147
rect 5146 2113 5183 2147
rect 5217 2113 5254 2147
rect 5288 2113 5325 2147
rect 5359 2113 5396 2147
rect 5430 2113 5467 2147
rect 5501 2113 5537 2147
rect 5571 2113 5607 2147
rect 5641 2113 5677 2147
rect 5711 2113 5716 2147
rect 4615 2071 5716 2113
rect 4649 2037 4686 2071
rect 4720 2037 4757 2071
rect 4791 2037 4828 2071
rect 4862 2037 4899 2071
rect 4933 2037 4970 2071
rect 5004 2037 5041 2071
rect 5075 2037 5112 2071
rect 5146 2037 5183 2071
rect 5217 2037 5254 2071
rect 5288 2037 5325 2071
rect 5359 2037 5396 2071
rect 5430 2037 5467 2071
rect 5501 2037 5537 2071
rect 5571 2037 5607 2071
rect 5641 2037 5677 2071
rect 5711 2037 5716 2071
rect 4615 1995 5716 2037
rect 4649 1961 4686 1995
rect 4720 1961 4757 1995
rect 4791 1961 4828 1995
rect 4862 1961 4899 1995
rect 4933 1961 4970 1995
rect 5004 1961 5041 1995
rect 5075 1961 5112 1995
rect 5146 1961 5183 1995
rect 5217 1961 5254 1995
rect 5288 1961 5325 1995
rect 5359 1961 5396 1995
rect 5430 1961 5467 1995
rect 5501 1961 5537 1995
rect 5571 1961 5607 1995
rect 5641 1961 5677 1995
rect 5711 1961 5716 1995
rect 4615 1919 5716 1961
rect 4649 1885 4686 1919
rect 4720 1885 4757 1919
rect 4791 1885 4828 1919
rect 4862 1885 4899 1919
rect 4933 1885 4970 1919
rect 5004 1885 5041 1919
rect 5075 1885 5112 1919
rect 5146 1885 5183 1919
rect 5217 1885 5254 1919
rect 5288 1885 5325 1919
rect 5359 1885 5396 1919
rect 5430 1885 5467 1919
rect 5501 1885 5537 1919
rect 5571 1885 5607 1919
rect 5641 1885 5677 1919
rect 5711 1885 5716 1919
rect 4615 1870 5716 1885
rect 2 1846 5716 1870
rect 2 792 33 1846
rect 5711 792 5716 1846
rect 2 771 5716 792
rect 10528 950 14944 957
rect 10528 916 10596 950
rect 10630 916 10665 950
rect 10699 916 10734 950
rect 10768 916 10803 950
rect 10837 916 10872 950
rect 10906 916 10941 950
rect 10975 916 11010 950
rect 11044 916 11078 950
rect 11112 916 11146 950
rect 11180 916 11214 950
rect 11248 916 11282 950
rect 11316 916 11350 950
rect 11384 916 11418 950
rect 11452 916 11486 950
rect 11520 916 11554 950
rect 11588 916 11622 950
rect 11656 916 11690 950
rect 11724 916 11758 950
rect 11792 916 11826 950
rect 11860 916 11894 950
rect 11928 916 11962 950
rect 11996 916 12030 950
rect 12064 916 12098 950
rect 12132 916 12166 950
rect 12200 916 12234 950
rect 12268 916 12302 950
rect 12336 916 12370 950
rect 12404 916 12438 950
rect 12472 916 12506 950
rect 12540 916 12574 950
rect 12608 916 12642 950
rect 12676 916 12710 950
rect 12744 916 12778 950
rect 12812 916 12846 950
rect 12880 916 12914 950
rect 12948 916 12982 950
rect 13016 916 13050 950
rect 13084 916 13118 950
rect 13152 916 13186 950
rect 13220 916 13254 950
rect 13288 916 13322 950
rect 13356 916 13390 950
rect 13424 916 13458 950
rect 13492 916 13526 950
rect 13560 916 13594 950
rect 13628 916 13662 950
rect 13696 916 13730 950
rect 13764 916 13798 950
rect 13832 916 13866 950
rect 13900 916 13934 950
rect 13968 916 14002 950
rect 14036 916 14070 950
rect 14104 916 14138 950
rect 14172 916 14206 950
rect 14240 916 14274 950
rect 14308 916 14342 950
rect 14376 916 14410 950
rect 14444 916 14478 950
rect 14512 916 14546 950
rect 14580 916 14614 950
rect 14648 916 14682 950
rect 14716 916 14750 950
rect 14784 916 14818 950
rect 14852 916 14886 950
rect 14920 916 14944 950
rect 10528 909 14944 916
rect 10528 839 10576 909
rect 2 768 5711 771
rect 6552 832 10576 839
rect 6552 798 6576 832
rect 6610 798 6645 832
rect 6679 798 6714 832
rect 6748 798 6783 832
rect 6817 798 6852 832
rect 6886 798 6921 832
rect 6955 798 6990 832
rect 7024 798 7059 832
rect 7093 798 7128 832
rect 7162 798 7197 832
rect 7231 798 7266 832
rect 7300 798 7335 832
rect 7369 798 7404 832
rect 7438 798 7473 832
rect 7507 798 7542 832
rect 7576 798 7611 832
rect 7645 798 7680 832
rect 7714 798 7749 832
rect 7783 798 7818 832
rect 7852 798 7887 832
rect 7921 798 7956 832
rect 7990 798 8025 832
rect 8059 798 8094 832
rect 8128 798 8162 832
rect 8196 798 8230 832
rect 8264 798 8298 832
rect 8332 798 8366 832
rect 8400 798 8434 832
rect 8468 798 8502 832
rect 8536 798 8570 832
rect 8604 798 8638 832
rect 8672 798 8706 832
rect 8740 798 8774 832
rect 8808 798 8842 832
rect 8876 798 8910 832
rect 8944 798 8978 832
rect 9012 798 9046 832
rect 9080 798 9114 832
rect 9148 798 9182 832
rect 9216 798 9250 832
rect 9284 798 9318 832
rect 9352 798 9386 832
rect 9420 798 9454 832
rect 9488 798 9522 832
rect 9556 798 9590 832
rect 9624 798 9658 832
rect 9692 798 9726 832
rect 9760 798 9794 832
rect 9828 798 9862 832
rect 9896 798 9930 832
rect 9964 798 9998 832
rect 10032 798 10066 832
rect 10100 798 10134 832
rect 10168 798 10202 832
rect 10236 798 10270 832
rect 10304 798 10338 832
rect 10372 798 10406 832
rect 10440 798 10474 832
rect 10508 798 10576 832
rect 6552 791 10576 798
rect 15938 -2511 15944 2175
rect 16726 2176 17215 2181
rect 16726 -2511 16732 2176
rect 15938 -2546 16732 -2511
rect 15938 -2580 15944 -2546
rect 15978 -2580 16012 -2546
rect 16046 -2580 16080 -2546
rect 16114 -2580 16148 -2546
rect 16182 -2580 16216 -2546
rect 16250 -2580 16284 -2546
rect 16318 -2580 16352 -2546
rect 16386 -2580 16420 -2546
rect 16454 -2580 16488 -2546
rect 16522 -2580 16556 -2546
rect 16590 -2580 16624 -2546
rect 16658 -2580 16692 -2546
rect 16726 -2580 16732 -2546
rect 15938 -2615 16732 -2580
rect 15938 -2649 15944 -2615
rect 15978 -2649 16012 -2615
rect 16046 -2649 16080 -2615
rect 16114 -2649 16148 -2615
rect 16182 -2649 16216 -2615
rect 16250 -2649 16284 -2615
rect 16318 -2649 16352 -2615
rect 16386 -2649 16420 -2615
rect 16454 -2649 16488 -2615
rect 16522 -2649 16556 -2615
rect 16590 -2649 16624 -2615
rect 16658 -2649 16692 -2615
rect 16726 -2649 16732 -2615
rect 15938 -2684 16732 -2649
rect 15938 -2718 15944 -2684
rect 15978 -2718 16012 -2684
rect 16046 -2718 16080 -2684
rect 16114 -2718 16148 -2684
rect 16182 -2718 16216 -2684
rect 16250 -2718 16284 -2684
rect 16318 -2718 16352 -2684
rect 16386 -2718 16420 -2684
rect 16454 -2718 16488 -2684
rect 16522 -2718 16556 -2684
rect 16590 -2718 16624 -2684
rect 16658 -2718 16692 -2684
rect 16726 -2718 16732 -2684
rect 15938 -2753 16732 -2718
rect 15938 -2787 15944 -2753
rect 15978 -2787 16012 -2753
rect 16046 -2787 16080 -2753
rect 16114 -2787 16148 -2753
rect 16182 -2787 16216 -2753
rect 16250 -2787 16284 -2753
rect 16318 -2787 16352 -2753
rect 16386 -2787 16420 -2753
rect 16454 -2787 16488 -2753
rect 16522 -2787 16556 -2753
rect 16590 -2787 16624 -2753
rect 16658 -2787 16692 -2753
rect 16726 -2787 16732 -2753
rect 15938 -2822 16732 -2787
rect 15938 -2856 15944 -2822
rect 15978 -2856 16012 -2822
rect 16046 -2856 16080 -2822
rect 16114 -2856 16148 -2822
rect 16182 -2856 16216 -2822
rect 16250 -2856 16284 -2822
rect 16318 -2856 16352 -2822
rect 16386 -2856 16420 -2822
rect 16454 -2856 16488 -2822
rect 16522 -2856 16556 -2822
rect 16590 -2856 16624 -2822
rect 16658 -2856 16692 -2822
rect 16726 -2856 16732 -2822
rect 15938 -2891 16732 -2856
rect 15938 -2925 15944 -2891
rect 15978 -2925 16012 -2891
rect 16046 -2925 16080 -2891
rect 16114 -2925 16148 -2891
rect 16182 -2925 16216 -2891
rect 16250 -2925 16284 -2891
rect 16318 -2925 16352 -2891
rect 16386 -2925 16420 -2891
rect 16454 -2925 16488 -2891
rect 16522 -2925 16556 -2891
rect 16590 -2925 16624 -2891
rect 16658 -2925 16692 -2891
rect 16726 -2925 16732 -2891
rect 15938 -2949 16732 -2925
rect 15939 -2975 16732 -2949
<< mvnsubdiff >>
rect 17430 11598 17677 14647
rect 17430 11498 17464 11598
rect -2750 4638 -88 4682
rect -2750 4498 433 4638
rect -2716 4464 -2680 4498
rect -2646 4464 -2610 4498
rect -2576 4464 -2540 4498
rect -2506 4464 -2470 4498
rect -2436 4464 -2400 4498
rect -2366 4464 -2330 4498
rect -2296 4464 -2260 4498
rect -2226 4464 -2190 4498
rect -2156 4464 -2120 4498
rect -2086 4464 -2050 4498
rect -2016 4464 -1980 4498
rect -1946 4464 -1910 4498
rect -1876 4464 -1840 4498
rect -1806 4464 -1770 4498
rect -1736 4464 -1700 4498
rect -1666 4464 -1630 4498
rect -1596 4464 -1560 4498
rect -1526 4464 -1490 4498
rect -1456 4464 -1421 4498
rect -1387 4464 -1352 4498
rect -1318 4464 -1283 4498
rect -1249 4464 -1214 4498
rect -1180 4464 -1145 4498
rect -1111 4464 -1076 4498
rect -1042 4464 -1007 4498
rect -973 4464 -938 4498
rect -904 4464 -869 4498
rect -835 4464 -800 4498
rect -766 4464 -731 4498
rect -697 4464 -662 4498
rect -628 4464 -593 4498
rect -559 4464 -524 4498
rect -490 4464 -455 4498
rect -421 4464 -386 4498
rect -352 4464 -317 4498
rect -283 4464 -248 4498
rect -214 4464 433 4498
rect -2750 4428 -148 4464
rect -2716 4394 -2680 4428
rect -2646 4394 -2610 4428
rect -2576 4394 -2540 4428
rect -2506 4394 -2470 4428
rect -2436 4394 -2400 4428
rect -2366 4394 -2330 4428
rect -2296 4394 -2260 4428
rect -2226 4394 -2190 4428
rect -2156 4394 -2120 4428
rect -2086 4394 -2050 4428
rect -2016 4394 -1980 4428
rect -1946 4394 -1910 4428
rect -1876 4394 -1840 4428
rect -1806 4394 -1770 4428
rect -1736 4394 -1700 4428
rect -1666 4394 -1630 4428
rect -1596 4394 -1560 4428
rect -1526 4394 -1490 4428
rect -1456 4394 -1421 4428
rect -1387 4394 -1352 4428
rect -1318 4394 -1283 4428
rect -1249 4394 -1214 4428
rect -1180 4394 -1145 4428
rect -1111 4394 -1076 4428
rect -1042 4394 -1007 4428
rect -973 4394 -938 4428
rect -904 4394 -869 4428
rect -835 4394 -800 4428
rect -766 4394 -731 4428
rect -697 4394 -662 4428
rect -628 4394 -593 4428
rect -559 4394 -524 4428
rect -490 4394 -455 4428
rect -421 4394 -386 4428
rect -352 4394 -317 4428
rect -283 4394 -248 4428
rect -214 4394 -148 4428
rect -2750 4358 -148 4394
rect -2716 4324 -2680 4358
rect -2646 4324 -2610 4358
rect -2576 4324 -2540 4358
rect -2506 4324 -2470 4358
rect -2436 4324 -2400 4358
rect -2366 4324 -2330 4358
rect -2296 4324 -2260 4358
rect -2226 4324 -2190 4358
rect -2156 4324 -2120 4358
rect -2086 4324 -2050 4358
rect -2016 4324 -1980 4358
rect -1946 4324 -1910 4358
rect -1876 4324 -1840 4358
rect -1806 4324 -1770 4358
rect -1736 4324 -1700 4358
rect -1666 4324 -1630 4358
rect -1596 4324 -1560 4358
rect -1526 4324 -1490 4358
rect -1456 4324 -1421 4358
rect -1387 4324 -1352 4358
rect -1318 4324 -1283 4358
rect -1249 4324 -1214 4358
rect -1180 4324 -1145 4358
rect -1111 4324 -1076 4358
rect -1042 4324 -1007 4358
rect -973 4324 -938 4358
rect -904 4324 -869 4358
rect -835 4324 -800 4358
rect -766 4324 -731 4358
rect -697 4324 -662 4358
rect -628 4324 -593 4358
rect -559 4324 -524 4358
rect -490 4324 -455 4358
rect -421 4324 -386 4358
rect -352 4324 -317 4358
rect -283 4324 -248 4358
rect -214 4324 -148 4358
rect -2750 4288 -148 4324
rect -2716 4254 -2680 4288
rect -2646 4254 -2610 4288
rect -2576 4254 -2540 4288
rect -2506 4254 -2470 4288
rect -2436 4254 -2400 4288
rect -2366 4254 -2330 4288
rect -2296 4254 -2260 4288
rect -2226 4254 -2190 4288
rect -2156 4254 -2120 4288
rect -2086 4254 -2050 4288
rect -2016 4254 -1980 4288
rect -1946 4254 -1910 4288
rect -1876 4254 -1840 4288
rect -1806 4254 -1770 4288
rect -1736 4254 -1700 4288
rect -1666 4254 -1630 4288
rect -1596 4254 -1560 4288
rect -1526 4254 -1490 4288
rect -1456 4254 -1421 4288
rect -1387 4254 -1352 4288
rect -1318 4254 -1283 4288
rect -1249 4254 -1214 4288
rect -1180 4254 -1145 4288
rect -1111 4254 -1076 4288
rect -1042 4254 -1007 4288
rect -973 4254 -938 4288
rect -904 4254 -869 4288
rect -835 4254 -800 4288
rect -766 4254 -731 4288
rect -697 4254 -662 4288
rect -628 4254 -593 4288
rect -559 4254 -524 4288
rect -490 4254 -455 4288
rect -421 4254 -386 4288
rect -352 4254 -317 4288
rect -283 4254 -248 4288
rect -214 4254 -148 4288
rect -2750 4218 -148 4254
rect 2 4232 433 4464
rect -2716 4184 -2680 4218
rect -2646 4184 -2610 4218
rect -2576 4184 -2540 4218
rect -2506 4184 -2470 4218
rect -2436 4184 -2400 4218
rect -2366 4184 -2330 4218
rect -2296 4184 -2260 4218
rect -2226 4184 -2190 4218
rect -2156 4184 -2120 4218
rect -2086 4184 -2050 4218
rect -2016 4184 -1980 4218
rect -1946 4184 -1910 4218
rect -1876 4184 -1840 4218
rect -1806 4184 -1770 4218
rect -1736 4184 -1700 4218
rect -1666 4184 -1630 4218
rect -1596 4184 -1560 4218
rect -1526 4184 -1490 4218
rect -1456 4184 -1421 4218
rect -1387 4184 -1352 4218
rect -1318 4184 -1283 4218
rect -1249 4184 -1214 4218
rect -1180 4184 -1145 4218
rect -1111 4184 -1076 4218
rect -1042 4184 -1007 4218
rect -973 4184 -938 4218
rect -904 4184 -869 4218
rect -835 4184 -800 4218
rect -766 4184 -731 4218
rect -697 4184 -662 4218
rect -628 4184 -593 4218
rect -559 4184 -524 4218
rect -490 4184 -455 4218
rect -421 4184 -386 4218
rect -352 4184 -317 4218
rect -283 4184 -248 4218
rect -214 4184 -148 4218
rect -2750 4148 -148 4184
rect -2716 4114 -2680 4148
rect -2646 4114 -2610 4148
rect -2576 4114 -2540 4148
rect -2506 4114 -2470 4148
rect -2436 4114 -2400 4148
rect -2366 4114 -2330 4148
rect -2296 4114 -2260 4148
rect -2226 4114 -2190 4148
rect -2156 4114 -2120 4148
rect -2086 4114 -2050 4148
rect -2016 4114 -1980 4148
rect -1946 4114 -1910 4148
rect -1876 4114 -1840 4148
rect -1806 4114 -1770 4148
rect -1736 4114 -1700 4148
rect -1666 4114 -1630 4148
rect -1596 4114 -1560 4148
rect -1526 4114 -1490 4148
rect -1456 4114 -1421 4148
rect -1387 4114 -1352 4148
rect -1318 4114 -1283 4148
rect -1249 4114 -1214 4148
rect -1180 4114 -1145 4148
rect -1111 4114 -1076 4148
rect -1042 4114 -1007 4148
rect -973 4114 -938 4148
rect -904 4114 -869 4148
rect -835 4114 -800 4148
rect -766 4114 -731 4148
rect -697 4114 -662 4148
rect -628 4114 -593 4148
rect -559 4114 -524 4148
rect -490 4114 -455 4148
rect -421 4114 -386 4148
rect -352 4114 -317 4148
rect -283 4114 -248 4148
rect -214 4114 -148 4148
rect -2750 4078 -148 4114
rect -2716 4044 -2680 4078
rect -2646 4044 -2610 4078
rect -2576 4044 -2540 4078
rect -2506 4044 -2470 4078
rect -2436 4044 -2400 4078
rect -2366 4044 -2330 4078
rect -2296 4044 -2260 4078
rect -2226 4044 -2190 4078
rect -2156 4044 -2120 4078
rect -2086 4044 -2050 4078
rect -2016 4044 -1980 4078
rect -1946 4044 -1910 4078
rect -1876 4044 -1840 4078
rect -1806 4044 -1770 4078
rect -1736 4044 -1700 4078
rect -1666 4044 -1630 4078
rect -1596 4044 -1560 4078
rect -1526 4044 -1490 4078
rect -1456 4044 -1421 4078
rect -1387 4044 -1352 4078
rect -1318 4044 -1283 4078
rect -1249 4044 -1214 4078
rect -1180 4044 -1145 4078
rect -1111 4044 -1076 4078
rect -1042 4044 -1007 4078
rect -973 4044 -938 4078
rect -904 4044 -869 4078
rect -835 4044 -800 4078
rect -766 4044 -731 4078
rect -697 4044 -662 4078
rect -628 4044 -593 4078
rect -559 4044 -524 4078
rect -490 4044 -455 4078
rect -421 4044 -386 4078
rect -352 4044 -317 4078
rect -283 4044 -248 4078
rect -214 4044 -148 4078
rect -2750 4008 -148 4044
rect -2716 3974 -2680 4008
rect -2646 3974 -2610 4008
rect -2576 3974 -2540 4008
rect -2506 3974 -2470 4008
rect -2436 3974 -2400 4008
rect -2366 3974 -2330 4008
rect -2296 3974 -2260 4008
rect -2226 3974 -2190 4008
rect -2156 3974 -2120 4008
rect -2086 3974 -2050 4008
rect -2016 3974 -1980 4008
rect -1946 3974 -1910 4008
rect -1876 3974 -1840 4008
rect -1806 3974 -1770 4008
rect -1736 3974 -1700 4008
rect -1666 3974 -1630 4008
rect -1596 3974 -1560 4008
rect -1526 3974 -1490 4008
rect -1456 3974 -1421 4008
rect -1387 3974 -1352 4008
rect -1318 3974 -1283 4008
rect -1249 3974 -1214 4008
rect -1180 3974 -1145 4008
rect -1111 3974 -1076 4008
rect -1042 3974 -1007 4008
rect -973 3974 -938 4008
rect -904 3974 -869 4008
rect -835 3974 -800 4008
rect -766 3974 -731 4008
rect -697 3974 -662 4008
rect -628 3974 -593 4008
rect -559 3974 -524 4008
rect -490 3974 -455 4008
rect -421 3974 -386 4008
rect -352 3974 -317 4008
rect -283 3974 -248 4008
rect -214 3974 -148 4008
rect -2750 3938 -148 3974
rect -2716 3904 -2680 3938
rect -2646 3904 -2610 3938
rect -2576 3904 -2540 3938
rect -2506 3904 -2470 3938
rect -2436 3904 -2400 3938
rect -2366 3904 -2330 3938
rect -2296 3904 -2260 3938
rect -2226 3904 -2190 3938
rect -2156 3904 -2120 3938
rect -2086 3904 -2050 3938
rect -2016 3904 -1980 3938
rect -1946 3904 -1910 3938
rect -1876 3904 -1840 3938
rect -1806 3904 -1770 3938
rect -1736 3904 -1700 3938
rect -1666 3904 -1630 3938
rect -1596 3904 -1560 3938
rect -1526 3904 -1490 3938
rect -1456 3904 -1421 3938
rect -1387 3904 -1352 3938
rect -1318 3904 -1283 3938
rect -1249 3904 -1214 3938
rect -1180 3904 -1145 3938
rect -1111 3904 -1076 3938
rect -1042 3904 -1007 3938
rect -973 3904 -938 3938
rect -904 3904 -869 3938
rect -835 3904 -800 3938
rect -766 3904 -731 3938
rect -697 3904 -662 3938
rect -628 3904 -593 3938
rect -559 3904 -524 3938
rect -490 3904 -455 3938
rect -421 3904 -386 3938
rect -352 3904 -317 3938
rect -283 3904 -248 3938
rect -214 3904 -148 3938
rect -2750 3868 -148 3904
rect -2716 3834 -2680 3868
rect -2646 3834 -2610 3868
rect -2576 3834 -2540 3868
rect -2506 3834 -2470 3868
rect -2436 3834 -2400 3868
rect -2366 3834 -2330 3868
rect -2296 3834 -2260 3868
rect -2226 3834 -2190 3868
rect -2156 3834 -2120 3868
rect -2086 3834 -2050 3868
rect -2016 3834 -1980 3868
rect -1946 3834 -1910 3868
rect -1876 3834 -1840 3868
rect -1806 3834 -1770 3868
rect -1736 3834 -1700 3868
rect -1666 3834 -1630 3868
rect -1596 3834 -1560 3868
rect -1526 3834 -1490 3868
rect -1456 3834 -1421 3868
rect -1387 3834 -1352 3868
rect -1318 3834 -1283 3868
rect -1249 3834 -1214 3868
rect -1180 3834 -1145 3868
rect -1111 3834 -1076 3868
rect -1042 3834 -1007 3868
rect -973 3834 -938 3868
rect -904 3834 -869 3868
rect -835 3834 -800 3868
rect -766 3834 -731 3868
rect -697 3834 -662 3868
rect -628 3834 -593 3868
rect -559 3834 -524 3868
rect -490 3834 -455 3868
rect -421 3834 -386 3868
rect -352 3834 -317 3868
rect -283 3834 -248 3868
rect -214 3834 -148 3868
rect -2750 3798 -148 3834
rect -2716 3764 -2680 3798
rect -2646 3764 -2610 3798
rect -2576 3764 -2540 3798
rect -2506 3764 -2470 3798
rect -2436 3764 -2400 3798
rect -2366 3764 -2330 3798
rect -2296 3764 -2260 3798
rect -2226 3764 -2190 3798
rect -2156 3764 -2120 3798
rect -2086 3764 -2050 3798
rect -2016 3764 -1980 3798
rect -1946 3764 -1910 3798
rect -1876 3764 -1840 3798
rect -1806 3764 -1770 3798
rect -1736 3764 -1700 3798
rect -1666 3764 -1630 3798
rect -1596 3764 -1560 3798
rect -1526 3764 -1490 3798
rect -1456 3764 -1421 3798
rect -1387 3764 -1352 3798
rect -1318 3764 -1283 3798
rect -1249 3764 -1214 3798
rect -1180 3764 -1145 3798
rect -1111 3764 -1076 3798
rect -1042 3764 -1007 3798
rect -973 3764 -938 3798
rect -904 3764 -869 3798
rect -835 3764 -800 3798
rect -766 3764 -731 3798
rect -697 3764 -662 3798
rect -628 3764 -593 3798
rect -559 3764 -524 3798
rect -490 3764 -455 3798
rect -421 3764 -386 3798
rect -352 3764 -317 3798
rect -283 3764 -248 3798
rect -214 3764 -148 3798
rect -2750 3728 -148 3764
rect -2716 3694 -2680 3728
rect -2646 3694 -2610 3728
rect -2576 3694 -2540 3728
rect -2506 3694 -2470 3728
rect -2436 3694 -2400 3728
rect -2366 3694 -2330 3728
rect -2296 3694 -2260 3728
rect -2226 3694 -2190 3728
rect -2156 3694 -2120 3728
rect -2086 3694 -2050 3728
rect -2016 3694 -1980 3728
rect -1946 3694 -1910 3728
rect -1876 3694 -1840 3728
rect -1806 3694 -1770 3728
rect -1736 3694 -1700 3728
rect -1666 3694 -1630 3728
rect -1596 3694 -1560 3728
rect -1526 3694 -1490 3728
rect -1456 3694 -1421 3728
rect -1387 3694 -1352 3728
rect -1318 3694 -1283 3728
rect -1249 3694 -1214 3728
rect -1180 3694 -1145 3728
rect -1111 3694 -1076 3728
rect -1042 3694 -1007 3728
rect -973 3694 -938 3728
rect -904 3694 -869 3728
rect -835 3694 -800 3728
rect -766 3694 -731 3728
rect -697 3694 -662 3728
rect -628 3694 -593 3728
rect -559 3694 -524 3728
rect -490 3694 -455 3728
rect -421 3694 -386 3728
rect -352 3694 -317 3728
rect -283 3694 -248 3728
rect -214 3694 -148 3728
rect -2750 3658 -148 3694
rect -2716 3624 -2680 3658
rect -2646 3624 -2610 3658
rect -2576 3624 -2540 3658
rect -2506 3624 -2470 3658
rect -2436 3624 -2400 3658
rect -2366 3624 -2330 3658
rect -2296 3624 -2260 3658
rect -2226 3624 -2190 3658
rect -2156 3624 -2120 3658
rect -2086 3624 -2050 3658
rect -2016 3624 -1980 3658
rect -1946 3624 -1910 3658
rect -1876 3624 -1840 3658
rect -1806 3624 -1770 3658
rect -1736 3624 -1700 3658
rect -1666 3624 -1630 3658
rect -1596 3624 -1560 3658
rect -1526 3624 -1490 3658
rect -1456 3624 -1421 3658
rect -1387 3624 -1352 3658
rect -1318 3624 -1283 3658
rect -1249 3624 -1214 3658
rect -1180 3624 -1145 3658
rect -1111 3624 -1076 3658
rect -1042 3624 -1007 3658
rect -973 3624 -938 3658
rect -904 3624 -869 3658
rect -835 3624 -800 3658
rect -766 3624 -731 3658
rect -697 3624 -662 3658
rect -628 3624 -593 3658
rect -559 3624 -524 3658
rect -490 3624 -455 3658
rect -421 3624 -386 3658
rect -352 3624 -317 3658
rect -283 3624 -248 3658
rect -214 3624 -148 3658
rect -2750 3588 -148 3624
rect -2716 3554 -2680 3588
rect -2646 3554 -2610 3588
rect -2576 3554 -2540 3588
rect -2506 3554 -2470 3588
rect -2436 3554 -2400 3588
rect -2366 3554 -2330 3588
rect -2296 3554 -2260 3588
rect -2226 3554 -2190 3588
rect -2156 3554 -2120 3588
rect -2086 3554 -2050 3588
rect -2016 3554 -1980 3588
rect -1946 3554 -1910 3588
rect -1876 3554 -1840 3588
rect -1806 3554 -1770 3588
rect -1736 3554 -1700 3588
rect -1666 3554 -1630 3588
rect -1596 3554 -1560 3588
rect -1526 3554 -1490 3588
rect -1456 3554 -1421 3588
rect -1387 3554 -1352 3588
rect -1318 3554 -1283 3588
rect -1249 3554 -1214 3588
rect -1180 3554 -1145 3588
rect -1111 3554 -1076 3588
rect -1042 3554 -1007 3588
rect -973 3554 -938 3588
rect -904 3554 -869 3588
rect -835 3554 -800 3588
rect -766 3554 -731 3588
rect -697 3554 -662 3588
rect -628 3554 -593 3588
rect -559 3554 -524 3588
rect -490 3554 -455 3588
rect -421 3554 -386 3588
rect -352 3554 -317 3588
rect -283 3554 -248 3588
rect -214 3554 -148 3588
rect -2750 3518 -148 3554
rect -2716 3484 -2680 3518
rect -2646 3484 -2610 3518
rect -2576 3484 -2540 3518
rect -2506 3484 -2470 3518
rect -2436 3484 -2400 3518
rect -2366 3484 -2330 3518
rect -2296 3484 -2260 3518
rect -2226 3484 -2190 3518
rect -2156 3484 -2120 3518
rect -2086 3484 -2050 3518
rect -2016 3484 -1980 3518
rect -1946 3484 -1910 3518
rect -1876 3484 -1840 3518
rect -1806 3484 -1770 3518
rect -1736 3484 -1700 3518
rect -1666 3484 -1630 3518
rect -1596 3484 -1560 3518
rect -1526 3484 -1490 3518
rect -1456 3484 -1421 3518
rect -1387 3484 -1352 3518
rect -1318 3484 -1283 3518
rect -1249 3484 -1214 3518
rect -1180 3484 -1145 3518
rect -1111 3484 -1076 3518
rect -1042 3484 -1007 3518
rect -973 3484 -938 3518
rect -904 3484 -869 3518
rect -835 3484 -800 3518
rect -766 3484 -731 3518
rect -697 3484 -662 3518
rect -628 3484 -593 3518
rect -559 3484 -524 3518
rect -490 3484 -455 3518
rect -421 3484 -386 3518
rect -352 3484 -317 3518
rect -283 3484 -248 3518
rect -214 3484 -148 3518
rect -2750 3448 -148 3484
rect -2716 3414 -2680 3448
rect -2646 3414 -2610 3448
rect -2576 3414 -2540 3448
rect -2506 3414 -2470 3448
rect -2436 3414 -2400 3448
rect -2366 3414 -2330 3448
rect -2296 3414 -2260 3448
rect -2226 3414 -2190 3448
rect -2156 3414 -2120 3448
rect -2086 3414 -2050 3448
rect -2016 3414 -1980 3448
rect -1946 3414 -1910 3448
rect -1876 3414 -1840 3448
rect -1806 3414 -1770 3448
rect -1736 3414 -1700 3448
rect -1666 3414 -1630 3448
rect -1596 3414 -1560 3448
rect -1526 3414 -1490 3448
rect -1456 3414 -1421 3448
rect -1387 3414 -1352 3448
rect -1318 3414 -1283 3448
rect -1249 3414 -1214 3448
rect -1180 3414 -1145 3448
rect -1111 3414 -1076 3448
rect -1042 3414 -1007 3448
rect -973 3414 -938 3448
rect -904 3414 -869 3448
rect -835 3414 -800 3448
rect -766 3414 -731 3448
rect -697 3414 -662 3448
rect -628 3414 -593 3448
rect -559 3414 -524 3448
rect -490 3414 -455 3448
rect -421 3414 -386 3448
rect -352 3414 -317 3448
rect -283 3414 -248 3448
rect -214 3414 -148 3448
rect -2750 3378 -148 3414
rect -2716 3344 -2680 3378
rect -2646 3344 -2610 3378
rect -2576 3344 -2540 3378
rect -2506 3344 -2470 3378
rect -2436 3344 -2400 3378
rect -2366 3344 -2330 3378
rect -2296 3344 -2260 3378
rect -2226 3344 -2190 3378
rect -2156 3344 -2120 3378
rect -2086 3344 -2050 3378
rect -2016 3344 -1980 3378
rect -1946 3344 -1910 3378
rect -1876 3344 -1840 3378
rect -1806 3344 -1770 3378
rect -1736 3344 -1700 3378
rect -1666 3344 -1630 3378
rect -1596 3344 -1560 3378
rect -1526 3344 -1490 3378
rect -1456 3344 -1421 3378
rect -1387 3344 -1352 3378
rect -1318 3344 -1283 3378
rect -1249 3344 -1214 3378
rect -1180 3344 -1145 3378
rect -1111 3344 -1076 3378
rect -1042 3344 -1007 3378
rect -973 3344 -938 3378
rect -904 3344 -869 3378
rect -835 3344 -800 3378
rect -766 3344 -731 3378
rect -697 3344 -662 3378
rect -628 3344 -593 3378
rect -559 3344 -524 3378
rect -490 3344 -455 3378
rect -421 3344 -386 3378
rect -352 3344 -317 3378
rect -283 3344 -248 3378
rect -214 3344 -148 3378
rect -2750 3308 -148 3344
rect -2716 3274 -2680 3308
rect -2646 3274 -2610 3308
rect -2576 3274 -2540 3308
rect -2506 3274 -2470 3308
rect -2436 3274 -2400 3308
rect -2366 3274 -2330 3308
rect -2296 3274 -2260 3308
rect -2226 3274 -2190 3308
rect -2156 3274 -2120 3308
rect -2086 3274 -2050 3308
rect -2016 3274 -1980 3308
rect -1946 3274 -1910 3308
rect -1876 3274 -1840 3308
rect -1806 3274 -1770 3308
rect -1736 3274 -1700 3308
rect -1666 3274 -1630 3308
rect -1596 3274 -1560 3308
rect -1526 3274 -1490 3308
rect -1456 3274 -1421 3308
rect -1387 3274 -1352 3308
rect -1318 3274 -1283 3308
rect -1249 3274 -1214 3308
rect -1180 3274 -1145 3308
rect -1111 3274 -1076 3308
rect -1042 3274 -1007 3308
rect -973 3274 -938 3308
rect -904 3274 -869 3308
rect -835 3274 -800 3308
rect -766 3274 -731 3308
rect -697 3274 -662 3308
rect -628 3274 -593 3308
rect -559 3274 -524 3308
rect -490 3274 -455 3308
rect -421 3274 -386 3308
rect -352 3274 -317 3308
rect -283 3274 -248 3308
rect -214 3274 -148 3308
rect -2750 3238 -148 3274
rect -2716 3204 -2680 3238
rect -2646 3204 -2610 3238
rect -2576 3204 -2540 3238
rect -2506 3204 -2470 3238
rect -2436 3204 -2400 3238
rect -2366 3204 -2330 3238
rect -2296 3204 -2260 3238
rect -2226 3204 -2190 3238
rect -2156 3204 -2120 3238
rect -2086 3204 -2050 3238
rect -2016 3204 -1980 3238
rect -1946 3204 -1910 3238
rect -1876 3204 -1840 3238
rect -1806 3204 -1770 3238
rect -1736 3204 -1700 3238
rect -1666 3204 -1630 3238
rect -1596 3204 -1560 3238
rect -1526 3204 -1490 3238
rect -1456 3204 -1421 3238
rect -1387 3204 -1352 3238
rect -1318 3204 -1283 3238
rect -1249 3204 -1214 3238
rect -1180 3204 -1145 3238
rect -1111 3204 -1076 3238
rect -1042 3204 -1007 3238
rect -973 3204 -938 3238
rect -904 3204 -869 3238
rect -835 3204 -800 3238
rect -766 3204 -731 3238
rect -697 3204 -662 3238
rect -628 3204 -593 3238
rect -559 3204 -524 3238
rect -490 3204 -455 3238
rect -421 3204 -386 3238
rect -352 3204 -317 3238
rect -283 3204 -248 3238
rect -214 3230 -148 3238
rect -214 3205 -101 3230
rect 231 3205 433 4232
rect -214 3204 433 3205
rect -2750 3168 433 3204
rect -2716 3134 -2680 3168
rect -2646 3134 -2610 3168
rect -2576 3134 -2540 3168
rect -2506 3134 -2470 3168
rect -2436 3134 -2400 3168
rect -2366 3134 -2330 3168
rect -2296 3134 -2260 3168
rect -2226 3134 -2190 3168
rect -2156 3134 -2120 3168
rect -2086 3134 -2050 3168
rect -2016 3134 -1980 3168
rect -1946 3134 -1910 3168
rect -1876 3134 -1840 3168
rect -1806 3134 -1770 3168
rect -1736 3134 -1700 3168
rect -1666 3134 -1630 3168
rect -1596 3134 -1560 3168
rect -1526 3134 -1490 3168
rect -1456 3134 -1421 3168
rect -1387 3134 -1352 3168
rect -1318 3134 -1283 3168
rect -1249 3134 -1214 3168
rect -1180 3134 -1145 3168
rect -1111 3134 -1076 3168
rect -1042 3134 -1007 3168
rect -973 3134 -938 3168
rect -904 3134 -869 3168
rect -835 3134 -800 3168
rect -766 3134 -731 3168
rect -697 3134 -662 3168
rect -628 3134 -593 3168
rect -559 3134 -524 3168
rect -490 3134 -455 3168
rect -421 3134 -386 3168
rect -352 3134 -317 3168
rect -283 3134 -248 3168
rect -214 3140 433 3168
rect -214 3134 -161 3140
rect -2750 3106 -161 3134
rect -127 3106 -89 3140
rect -55 3106 -17 3140
rect 17 3106 55 3140
rect 89 3106 127 3140
rect 161 3106 199 3140
rect 233 3106 271 3140
rect 305 3106 433 3140
rect -2750 3098 433 3106
rect -2716 3064 -2680 3098
rect -2646 3064 -2610 3098
rect -2576 3064 -2540 3098
rect -2506 3064 -2470 3098
rect -2436 3064 -2400 3098
rect -2366 3064 -2330 3098
rect -2296 3064 -2260 3098
rect -2226 3064 -2190 3098
rect -2156 3064 -2120 3098
rect -2086 3064 -2050 3098
rect -2016 3064 -1980 3098
rect -1946 3064 -1910 3098
rect -1876 3064 -1840 3098
rect -1806 3064 -1770 3098
rect -1736 3064 -1700 3098
rect -1666 3064 -1630 3098
rect -1596 3064 -1560 3098
rect -1526 3064 -1490 3098
rect -1456 3064 -1421 3098
rect -1387 3064 -1352 3098
rect -1318 3064 -1283 3098
rect -1249 3064 -1214 3098
rect -1180 3064 -1145 3098
rect -1111 3064 -1076 3098
rect -1042 3064 -1007 3098
rect -973 3064 -938 3098
rect -904 3064 -869 3098
rect -835 3064 -800 3098
rect -766 3064 -731 3098
rect -697 3064 -662 3098
rect -628 3064 -593 3098
rect -559 3064 -524 3098
rect -490 3064 -455 3098
rect -421 3064 -386 3098
rect -352 3064 -317 3098
rect -283 3064 -248 3098
rect -214 3071 433 3098
rect -214 3064 -161 3071
rect -2750 3037 -161 3064
rect -127 3037 -89 3071
rect -55 3037 -17 3071
rect 17 3037 55 3071
rect 89 3037 127 3071
rect 161 3037 199 3071
rect 233 3037 271 3071
rect 305 3037 433 3071
rect -2750 3028 433 3037
rect -2716 2994 -2680 3028
rect -2646 2994 -2610 3028
rect -2576 2994 -2540 3028
rect -2506 2994 -2470 3028
rect -2436 2994 -2400 3028
rect -2366 2994 -2330 3028
rect -2296 2994 -2260 3028
rect -2226 2994 -2190 3028
rect -2156 2994 -2120 3028
rect -2086 2994 -2050 3028
rect -2016 2994 -1980 3028
rect -1946 2994 -1910 3028
rect -1876 2994 -1840 3028
rect -1806 2994 -1770 3028
rect -1736 2994 -1700 3028
rect -1666 2994 -1630 3028
rect -1596 2994 -1560 3028
rect -1526 2994 -1490 3028
rect -1456 2994 -1421 3028
rect -1387 2994 -1352 3028
rect -1318 2994 -1283 3028
rect -1249 2994 -1214 3028
rect -1180 2994 -1145 3028
rect -1111 2994 -1076 3028
rect -1042 2994 -1007 3028
rect -973 2994 -938 3028
rect -904 2994 -869 3028
rect -835 2994 -800 3028
rect -766 2994 -731 3028
rect -697 2994 -662 3028
rect -628 2994 -593 3028
rect -559 2994 -524 3028
rect -490 2994 -455 3028
rect -421 2994 -386 3028
rect -352 2994 -317 3028
rect -283 2994 -248 3028
rect -214 3002 433 3028
rect -214 2994 -161 3002
rect -2750 2968 -161 2994
rect -127 2968 -89 3002
rect -55 2968 -17 3002
rect 17 2968 55 3002
rect 89 2968 127 3002
rect 161 2968 199 3002
rect 233 2968 271 3002
rect 305 2968 433 3002
rect -2750 2958 433 2968
rect -2716 2924 -2680 2958
rect -2646 2924 -2610 2958
rect -2576 2924 -2540 2958
rect -2506 2924 -2470 2958
rect -2436 2924 -2400 2958
rect -2366 2924 -2330 2958
rect -2296 2924 -2260 2958
rect -2226 2924 -2190 2958
rect -2156 2924 -2120 2958
rect -2086 2924 -2050 2958
rect -2016 2924 -1980 2958
rect -1946 2924 -1910 2958
rect -1876 2924 -1840 2958
rect -1806 2924 -1770 2958
rect -1736 2924 -1700 2958
rect -1666 2924 -1630 2958
rect -1596 2924 -1560 2958
rect -1526 2924 -1490 2958
rect -1456 2924 -1421 2958
rect -1387 2924 -1352 2958
rect -1318 2924 -1283 2958
rect -1249 2924 -1214 2958
rect -1180 2924 -1145 2958
rect -1111 2924 -1076 2958
rect -1042 2924 -1007 2958
rect -973 2924 -938 2958
rect -904 2924 -869 2958
rect -835 2924 -800 2958
rect -766 2924 -731 2958
rect -697 2924 -662 2958
rect -628 2924 -593 2958
rect -559 2924 -524 2958
rect -490 2924 -455 2958
rect -421 2924 -386 2958
rect -352 2924 -317 2958
rect -283 2924 -248 2958
rect -214 2933 433 2958
rect -214 2924 -161 2933
rect -2750 2899 -161 2924
rect -127 2899 -89 2933
rect -55 2899 -17 2933
rect 17 2899 55 2933
rect 89 2899 127 2933
rect 161 2899 199 2933
rect 233 2899 271 2933
rect 305 2899 433 2933
rect -2750 2888 433 2899
rect -2716 2854 -2680 2888
rect -2646 2854 -2610 2888
rect -2576 2854 -2540 2888
rect -2506 2854 -2470 2888
rect -2436 2854 -2400 2888
rect -2366 2854 -2330 2888
rect -2296 2854 -2260 2888
rect -2226 2854 -2190 2888
rect -2156 2854 -2120 2888
rect -2086 2854 -2050 2888
rect -2016 2854 -1980 2888
rect -1946 2854 -1910 2888
rect -1876 2854 -1840 2888
rect -1806 2854 -1770 2888
rect -1736 2854 -1700 2888
rect -1666 2854 -1630 2888
rect -1596 2854 -1560 2888
rect -1526 2854 -1490 2888
rect -1456 2854 -1421 2888
rect -1387 2854 -1352 2888
rect -1318 2854 -1283 2888
rect -1249 2854 -1214 2888
rect -1180 2854 -1145 2888
rect -1111 2854 -1076 2888
rect -1042 2854 -1007 2888
rect -973 2854 -938 2888
rect -904 2854 -869 2888
rect -835 2854 -800 2888
rect -766 2854 -731 2888
rect -697 2854 -662 2888
rect -628 2854 -593 2888
rect -559 2854 -524 2888
rect -490 2854 -455 2888
rect -421 2854 -386 2888
rect -352 2854 -317 2888
rect -283 2854 -248 2888
rect -214 2863 433 2888
rect -214 2854 -161 2863
rect -2750 2829 -161 2854
rect -127 2829 -89 2863
rect -55 2829 -17 2863
rect 17 2829 55 2863
rect 89 2829 127 2863
rect 161 2829 199 2863
rect 233 2829 271 2863
rect 305 2829 433 2863
rect -2750 2818 433 2829
rect -2716 2784 -2680 2818
rect -2646 2784 -2610 2818
rect -2576 2784 -2540 2818
rect -2506 2784 -2470 2818
rect -2436 2784 -2400 2818
rect -2366 2784 -2330 2818
rect -2296 2784 -2260 2818
rect -2226 2784 -2190 2818
rect -2156 2784 -2120 2818
rect -2086 2784 -2050 2818
rect -2016 2784 -1980 2818
rect -1946 2784 -1910 2818
rect -1876 2784 -1840 2818
rect -1806 2784 -1770 2818
rect -1736 2784 -1700 2818
rect -1666 2784 -1630 2818
rect -1596 2784 -1560 2818
rect -1526 2784 -1490 2818
rect -1456 2784 -1421 2818
rect -1387 2784 -1352 2818
rect -1318 2784 -1283 2818
rect -1249 2784 -1214 2818
rect -1180 2784 -1145 2818
rect -1111 2784 -1076 2818
rect -1042 2784 -1007 2818
rect -973 2784 -938 2818
rect -904 2784 -869 2818
rect -835 2784 -800 2818
rect -766 2784 -731 2818
rect -697 2784 -662 2818
rect -628 2784 -593 2818
rect -559 2784 -524 2818
rect -490 2784 -455 2818
rect -421 2784 -386 2818
rect -352 2784 -317 2818
rect -283 2784 -248 2818
rect -214 2793 433 2818
rect -214 2784 -161 2793
rect -2750 2759 -161 2784
rect -127 2759 -89 2793
rect -55 2759 -17 2793
rect 17 2759 55 2793
rect 89 2759 127 2793
rect 161 2759 199 2793
rect 233 2759 271 2793
rect 305 2759 433 2793
rect -2750 2748 433 2759
rect -2716 2714 -2680 2748
rect -2646 2714 -2610 2748
rect -2576 2714 -2540 2748
rect -2506 2714 -2470 2748
rect -2436 2714 -2400 2748
rect -2366 2714 -2330 2748
rect -2296 2714 -2260 2748
rect -2226 2714 -2190 2748
rect -2156 2714 -2120 2748
rect -2086 2714 -2050 2748
rect -2016 2714 -1980 2748
rect -1946 2714 -1910 2748
rect -1876 2714 -1840 2748
rect -1806 2714 -1770 2748
rect -1736 2714 -1700 2748
rect -1666 2714 -1630 2748
rect -1596 2714 -1560 2748
rect -1526 2714 -1490 2748
rect -1456 2714 -1421 2748
rect -1387 2714 -1352 2748
rect -1318 2714 -1283 2748
rect -1249 2714 -1214 2748
rect -1180 2714 -1145 2748
rect -1111 2714 -1076 2748
rect -1042 2714 -1007 2748
rect -973 2714 -938 2748
rect -904 2714 -869 2748
rect -835 2714 -800 2748
rect -766 2714 -731 2748
rect -697 2714 -662 2748
rect -628 2714 -593 2748
rect -559 2714 -524 2748
rect -490 2714 -455 2748
rect -421 2714 -386 2748
rect -352 2714 -317 2748
rect -283 2714 -248 2748
rect -214 2723 433 2748
rect -214 2714 -161 2723
rect -2750 2689 -161 2714
rect -127 2689 -89 2723
rect -55 2689 -17 2723
rect 17 2689 55 2723
rect 89 2689 127 2723
rect 161 2689 199 2723
rect 233 2689 271 2723
rect 305 2689 433 2723
rect -2750 2678 433 2689
rect -2716 2644 -2680 2678
rect -2646 2644 -2610 2678
rect -2576 2644 -2540 2678
rect -2506 2644 -2470 2678
rect -2436 2644 -2400 2678
rect -2366 2644 -2330 2678
rect -2296 2644 -2260 2678
rect -2226 2644 -2190 2678
rect -2156 2644 -2120 2678
rect -2086 2644 -2050 2678
rect -2016 2644 -1980 2678
rect -1946 2644 -1910 2678
rect -1876 2644 -1840 2678
rect -1806 2644 -1770 2678
rect -1736 2644 -1700 2678
rect -1666 2644 -1630 2678
rect -1596 2644 -1560 2678
rect -1526 2644 -1490 2678
rect -1456 2644 -1421 2678
rect -1387 2644 -1352 2678
rect -1318 2644 -1283 2678
rect -1249 2644 -1214 2678
rect -1180 2644 -1145 2678
rect -1111 2644 -1076 2678
rect -1042 2644 -1007 2678
rect -973 2644 -938 2678
rect -904 2644 -869 2678
rect -835 2644 -800 2678
rect -766 2644 -731 2678
rect -697 2644 -662 2678
rect -628 2644 -593 2678
rect -559 2644 -524 2678
rect -490 2644 -455 2678
rect -421 2644 -386 2678
rect -352 2644 -317 2678
rect -283 2644 -248 2678
rect -214 2653 433 2678
rect -214 2644 -161 2653
rect -2750 2619 -161 2644
rect -127 2619 -89 2653
rect -55 2619 -17 2653
rect 17 2619 55 2653
rect 89 2619 127 2653
rect 161 2619 199 2653
rect 233 2619 271 2653
rect 305 2619 433 2653
rect -2750 2608 433 2619
rect -2716 2574 -2680 2608
rect -2646 2574 -2610 2608
rect -2576 2574 -2540 2608
rect -2506 2574 -2470 2608
rect -2436 2574 -2400 2608
rect -2366 2574 -2330 2608
rect -2296 2574 -2260 2608
rect -2226 2574 -2190 2608
rect -2156 2574 -2120 2608
rect -2086 2574 -2050 2608
rect -2016 2574 -1980 2608
rect -1946 2574 -1910 2608
rect -1876 2574 -1840 2608
rect -1806 2574 -1770 2608
rect -1736 2574 -1700 2608
rect -1666 2574 -1630 2608
rect -1596 2574 -1560 2608
rect -1526 2574 -1490 2608
rect -1456 2574 -1421 2608
rect -1387 2574 -1352 2608
rect -1318 2574 -1283 2608
rect -1249 2574 -1214 2608
rect -1180 2574 -1145 2608
rect -1111 2574 -1076 2608
rect -1042 2574 -1007 2608
rect -973 2574 -938 2608
rect -904 2574 -869 2608
rect -835 2574 -800 2608
rect -766 2574 -731 2608
rect -697 2574 -662 2608
rect -628 2574 -593 2608
rect -559 2574 -524 2608
rect -490 2574 -455 2608
rect -421 2574 -386 2608
rect -352 2574 -317 2608
rect -283 2574 -248 2608
rect -214 2583 433 2608
rect -214 2574 -161 2583
rect -2750 2549 -161 2574
rect -127 2549 -89 2583
rect -55 2549 -17 2583
rect 17 2549 55 2583
rect 89 2549 127 2583
rect 161 2549 199 2583
rect 233 2549 271 2583
rect 305 2549 433 2583
rect -2750 2538 433 2549
rect -2716 2504 -2680 2538
rect -2646 2504 -2610 2538
rect -2576 2504 -2540 2538
rect -2506 2504 -2470 2538
rect -2436 2504 -2400 2538
rect -2366 2504 -2330 2538
rect -2296 2504 -2260 2538
rect -2226 2504 -2190 2538
rect -2156 2504 -2120 2538
rect -2086 2504 -2050 2538
rect -2016 2504 -1980 2538
rect -1946 2504 -1910 2538
rect -1876 2504 -1840 2538
rect -1806 2504 -1770 2538
rect -1736 2504 -1700 2538
rect -1666 2504 -1630 2538
rect -1596 2504 -1560 2538
rect -1526 2504 -1490 2538
rect -1456 2504 -1421 2538
rect -1387 2504 -1352 2538
rect -1318 2504 -1283 2538
rect -1249 2504 -1214 2538
rect -1180 2504 -1145 2538
rect -1111 2504 -1076 2538
rect -1042 2504 -1007 2538
rect -973 2504 -938 2538
rect -904 2504 -869 2538
rect -835 2504 -800 2538
rect -766 2504 -731 2538
rect -697 2504 -662 2538
rect -628 2504 -593 2538
rect -559 2504 -524 2538
rect -490 2504 -455 2538
rect -421 2504 -386 2538
rect -352 2504 -317 2538
rect -283 2504 -248 2538
rect -214 2513 433 2538
rect -214 2504 -161 2513
rect -2750 2479 -161 2504
rect -127 2479 -89 2513
rect -55 2479 -17 2513
rect 17 2479 55 2513
rect 89 2479 127 2513
rect 161 2479 199 2513
rect 233 2479 271 2513
rect 305 2479 433 2513
rect -2750 2468 433 2479
rect -2716 2434 -2680 2468
rect -2646 2434 -2610 2468
rect -2576 2434 -2540 2468
rect -2506 2434 -2470 2468
rect -2436 2434 -2400 2468
rect -2366 2434 -2330 2468
rect -2296 2434 -2260 2468
rect -2226 2434 -2190 2468
rect -2156 2434 -2120 2468
rect -2086 2434 -2050 2468
rect -2016 2434 -1980 2468
rect -1946 2434 -1910 2468
rect -1876 2434 -1840 2468
rect -1806 2434 -1770 2468
rect -1736 2434 -1700 2468
rect -1666 2434 -1630 2468
rect -1596 2434 -1560 2468
rect -1526 2434 -1490 2468
rect -1456 2434 -1421 2468
rect -1387 2434 -1352 2468
rect -1318 2434 -1283 2468
rect -1249 2434 -1214 2468
rect -1180 2434 -1145 2468
rect -1111 2434 -1076 2468
rect -1042 2434 -1007 2468
rect -973 2434 -938 2468
rect -904 2434 -869 2468
rect -835 2434 -800 2468
rect -766 2434 -731 2468
rect -697 2434 -662 2468
rect -628 2434 -593 2468
rect -559 2434 -524 2468
rect -490 2434 -455 2468
rect -421 2434 -386 2468
rect -352 2434 -317 2468
rect -283 2434 -248 2468
rect -214 2443 433 2468
rect -214 2434 -161 2443
rect -2750 2409 -161 2434
rect -127 2409 -89 2443
rect -55 2409 -17 2443
rect 17 2409 55 2443
rect 89 2409 127 2443
rect 161 2409 199 2443
rect 233 2409 271 2443
rect 305 2409 433 2443
rect -2750 2398 433 2409
rect -2716 2364 -2680 2398
rect -2646 2364 -2610 2398
rect -2576 2364 -2540 2398
rect -2506 2364 -2470 2398
rect -2436 2364 -2400 2398
rect -2366 2364 -2330 2398
rect -2296 2364 -2260 2398
rect -2226 2364 -2190 2398
rect -2156 2364 -2120 2398
rect -2086 2364 -2050 2398
rect -2016 2364 -1980 2398
rect -1946 2364 -1910 2398
rect -1876 2364 -1840 2398
rect -1806 2364 -1770 2398
rect -1736 2364 -1700 2398
rect -1666 2364 -1630 2398
rect -1596 2364 -1560 2398
rect -1526 2364 -1490 2398
rect -1456 2364 -1421 2398
rect -1387 2364 -1352 2398
rect -1318 2364 -1283 2398
rect -1249 2364 -1214 2398
rect -1180 2364 -1145 2398
rect -1111 2364 -1076 2398
rect -1042 2364 -1007 2398
rect -973 2364 -938 2398
rect -904 2364 -869 2398
rect -835 2364 -800 2398
rect -766 2364 -731 2398
rect -697 2364 -662 2398
rect -628 2364 -593 2398
rect -559 2364 -524 2398
rect -490 2364 -455 2398
rect -421 2364 -386 2398
rect -352 2364 -317 2398
rect -283 2364 -248 2398
rect -214 2373 433 2398
rect -214 2364 -161 2373
rect -2750 2339 -161 2364
rect -127 2339 -89 2373
rect -55 2339 -17 2373
rect 17 2339 55 2373
rect 89 2339 127 2373
rect 161 2339 199 2373
rect 233 2339 271 2373
rect 305 2339 433 2373
rect -2750 2328 433 2339
rect -2716 2294 -2680 2328
rect -2646 2294 -2610 2328
rect -2576 2294 -2540 2328
rect -2506 2294 -2470 2328
rect -2436 2294 -2400 2328
rect -2366 2294 -2330 2328
rect -2296 2294 -2260 2328
rect -2226 2294 -2190 2328
rect -2156 2294 -2120 2328
rect -2086 2294 -2050 2328
rect -2016 2294 -1980 2328
rect -1946 2294 -1910 2328
rect -1876 2294 -1840 2328
rect -1806 2294 -1770 2328
rect -1736 2294 -1700 2328
rect -1666 2294 -1630 2328
rect -1596 2294 -1560 2328
rect -1526 2294 -1490 2328
rect -1456 2294 -1421 2328
rect -1387 2294 -1352 2328
rect -1318 2294 -1283 2328
rect -1249 2294 -1214 2328
rect -1180 2294 -1145 2328
rect -1111 2294 -1076 2328
rect -1042 2294 -1007 2328
rect -973 2294 -938 2328
rect -904 2294 -869 2328
rect -835 2294 -800 2328
rect -766 2294 -731 2328
rect -697 2294 -662 2328
rect -628 2294 -593 2328
rect -559 2294 -524 2328
rect -490 2294 -455 2328
rect -421 2294 -386 2328
rect -352 2294 -317 2328
rect -283 2294 -248 2328
rect -214 2303 433 2328
rect 2154 4564 4549 4655
rect 11032 4564 11698 4654
rect 2154 4528 4449 4564
rect 2154 4494 2304 4528
rect 2338 4494 2374 4528
rect 2408 4494 2444 4528
rect 2478 4494 2514 4528
rect 2548 4494 2584 4528
rect 2618 4494 2654 4528
rect 2688 4494 2724 4528
rect 2758 4494 2794 4528
rect 2828 4494 2864 4528
rect 2898 4494 2934 4528
rect 2968 4494 3004 4528
rect 3038 4494 3074 4528
rect 3108 4494 3144 4528
rect 3178 4494 3214 4528
rect 3248 4494 3284 4528
rect 3318 4494 3354 4528
rect 3388 4494 3424 4528
rect 3458 4494 3494 4528
rect 3528 4494 3563 4528
rect 3597 4494 3632 4528
rect 3666 4494 3701 4528
rect 3735 4494 3770 4528
rect 3804 4494 3839 4528
rect 3873 4494 3908 4528
rect 3942 4494 3977 4528
rect 4011 4494 4046 4528
rect 4080 4494 4115 4528
rect 4149 4494 4184 4528
rect 4218 4494 4253 4528
rect 4287 4494 4322 4528
rect 4356 4494 4391 4528
rect 4425 4494 4449 4528
rect 2154 4460 4449 4494
rect 2154 4426 2304 4460
rect 2338 4426 2374 4460
rect 2408 4426 2444 4460
rect 2478 4426 2514 4460
rect 2548 4426 2584 4460
rect 2618 4426 2654 4460
rect 2688 4426 2724 4460
rect 2758 4426 2794 4460
rect 2828 4426 2864 4460
rect 2898 4426 2934 4460
rect 2968 4426 3004 4460
rect 3038 4426 3074 4460
rect 3108 4426 3144 4460
rect 3178 4426 3214 4460
rect 3248 4426 3284 4460
rect 3318 4426 3354 4460
rect 3388 4426 3424 4460
rect 3458 4426 3494 4460
rect 3528 4426 3563 4460
rect 3597 4426 3632 4460
rect 3666 4426 3701 4460
rect 3735 4426 3770 4460
rect 3804 4426 3839 4460
rect 3873 4426 3908 4460
rect 3942 4426 3977 4460
rect 4011 4426 4046 4460
rect 4080 4426 4115 4460
rect 4149 4426 4184 4460
rect 4218 4426 4253 4460
rect 4287 4426 4322 4460
rect 4356 4426 4391 4460
rect 4425 4426 4449 4460
rect 2154 4392 4449 4426
rect 2154 4358 2304 4392
rect 2338 4358 2374 4392
rect 2408 4358 2444 4392
rect 2478 4358 2514 4392
rect 2548 4358 2584 4392
rect 2618 4358 2654 4392
rect 2688 4358 2724 4392
rect 2758 4358 2794 4392
rect 2828 4358 2864 4392
rect 2898 4358 2934 4392
rect 2968 4358 3004 4392
rect 3038 4358 3074 4392
rect 3108 4358 3144 4392
rect 3178 4358 3214 4392
rect 3248 4358 3284 4392
rect 3318 4358 3354 4392
rect 3388 4358 3424 4392
rect 3458 4358 3494 4392
rect 3528 4358 3563 4392
rect 3597 4358 3632 4392
rect 3666 4358 3701 4392
rect 3735 4358 3770 4392
rect 3804 4358 3839 4392
rect 3873 4358 3908 4392
rect 3942 4358 3977 4392
rect 4011 4358 4046 4392
rect 4080 4358 4115 4392
rect 4149 4358 4184 4392
rect 4218 4358 4253 4392
rect 4287 4358 4322 4392
rect 4356 4358 4391 4392
rect 4425 4358 4449 4392
rect 2154 4324 4449 4358
rect 2154 4290 2304 4324
rect 2338 4290 2374 4324
rect 2408 4290 2444 4324
rect 2478 4290 2514 4324
rect 2548 4290 2584 4324
rect 2618 4290 2654 4324
rect 2688 4290 2724 4324
rect 2758 4290 2794 4324
rect 2828 4290 2864 4324
rect 2898 4290 2934 4324
rect 2968 4290 3004 4324
rect 3038 4290 3074 4324
rect 3108 4290 3144 4324
rect 3178 4290 3214 4324
rect 3248 4290 3284 4324
rect 3318 4290 3354 4324
rect 3388 4290 3424 4324
rect 3458 4290 3494 4324
rect 3528 4290 3563 4324
rect 3597 4290 3632 4324
rect 3666 4290 3701 4324
rect 3735 4290 3770 4324
rect 3804 4290 3839 4324
rect 3873 4290 3908 4324
rect 3942 4290 3977 4324
rect 4011 4290 4046 4324
rect 4080 4290 4115 4324
rect 4149 4290 4184 4324
rect 4218 4290 4253 4324
rect 4287 4290 4322 4324
rect 4356 4290 4391 4324
rect 4425 4290 4449 4324
rect 2154 4256 4449 4290
rect 2154 4222 2304 4256
rect 2338 4222 2374 4256
rect 2408 4222 2444 4256
rect 2478 4222 2514 4256
rect 2548 4222 2584 4256
rect 2618 4222 2654 4256
rect 2688 4222 2724 4256
rect 2758 4222 2794 4256
rect 2828 4222 2864 4256
rect 2898 4222 2934 4256
rect 2968 4222 3004 4256
rect 3038 4222 3074 4256
rect 3108 4222 3144 4256
rect 3178 4222 3214 4256
rect 3248 4222 3284 4256
rect 3318 4222 3354 4256
rect 3388 4222 3424 4256
rect 3458 4222 3494 4256
rect 3528 4222 3563 4256
rect 3597 4222 3632 4256
rect 3666 4222 3701 4256
rect 3735 4222 3770 4256
rect 3804 4222 3839 4256
rect 3873 4222 3908 4256
rect 3942 4222 3977 4256
rect 4011 4222 4046 4256
rect 4080 4222 4115 4256
rect 4149 4222 4184 4256
rect 4218 4222 4253 4256
rect 4287 4222 4322 4256
rect 4356 4222 4391 4256
rect 4425 4222 4449 4256
rect 2154 4188 4449 4222
rect 2154 4154 2304 4188
rect 2338 4154 2374 4188
rect 2408 4154 2444 4188
rect 2478 4154 2514 4188
rect 2548 4154 2584 4188
rect 2618 4154 2654 4188
rect 2688 4154 2724 4188
rect 2758 4154 2794 4188
rect 2828 4154 2864 4188
rect 2898 4154 2934 4188
rect 2968 4154 3004 4188
rect 3038 4154 3074 4188
rect 3108 4154 3144 4188
rect 3178 4154 3214 4188
rect 3248 4154 3284 4188
rect 3318 4154 3354 4188
rect 3388 4154 3424 4188
rect 3458 4154 3494 4188
rect 3528 4154 3563 4188
rect 3597 4154 3632 4188
rect 3666 4154 3701 4188
rect 3735 4154 3770 4188
rect 3804 4154 3839 4188
rect 3873 4154 3908 4188
rect 3942 4154 3977 4188
rect 4011 4154 4046 4188
rect 4080 4154 4115 4188
rect 4149 4154 4184 4188
rect 4218 4154 4253 4188
rect 4287 4154 4322 4188
rect 4356 4154 4391 4188
rect 4425 4154 4449 4188
rect 2154 4120 4449 4154
rect 2154 4086 2304 4120
rect 2338 4086 2374 4120
rect 2408 4086 2444 4120
rect 2478 4086 2514 4120
rect 2548 4086 2584 4120
rect 2618 4086 2654 4120
rect 2688 4086 2724 4120
rect 2758 4086 2794 4120
rect 2828 4086 2864 4120
rect 2898 4086 2934 4120
rect 2968 4086 3004 4120
rect 3038 4086 3074 4120
rect 3108 4086 3144 4120
rect 3178 4086 3214 4120
rect 3248 4086 3284 4120
rect 3318 4086 3354 4120
rect 3388 4086 3424 4120
rect 3458 4086 3494 4120
rect 3528 4086 3563 4120
rect 3597 4086 3632 4120
rect 3666 4086 3701 4120
rect 3735 4086 3770 4120
rect 3804 4086 3839 4120
rect 3873 4086 3908 4120
rect 3942 4086 3977 4120
rect 4011 4086 4046 4120
rect 4080 4086 4115 4120
rect 4149 4086 4184 4120
rect 4218 4086 4253 4120
rect 4287 4086 4322 4120
rect 4356 4086 4391 4120
rect 4425 4086 4449 4120
rect 2154 4052 4449 4086
rect 2154 4018 2304 4052
rect 2338 4018 2374 4052
rect 2408 4018 2444 4052
rect 2478 4018 2514 4052
rect 2548 4018 2584 4052
rect 2618 4018 2654 4052
rect 2688 4018 2724 4052
rect 2758 4018 2794 4052
rect 2828 4018 2864 4052
rect 2898 4018 2934 4052
rect 2968 4018 3004 4052
rect 3038 4018 3074 4052
rect 3108 4018 3144 4052
rect 3178 4018 3214 4052
rect 3248 4018 3284 4052
rect 3318 4018 3354 4052
rect 3388 4018 3424 4052
rect 3458 4018 3494 4052
rect 3528 4018 3563 4052
rect 3597 4018 3632 4052
rect 3666 4018 3701 4052
rect 3735 4018 3770 4052
rect 3804 4018 3839 4052
rect 3873 4018 3908 4052
rect 3942 4018 3977 4052
rect 4011 4018 4046 4052
rect 4080 4018 4115 4052
rect 4149 4018 4184 4052
rect 4218 4018 4253 4052
rect 4287 4018 4322 4052
rect 4356 4018 4391 4052
rect 4425 4018 4449 4052
rect 2154 3984 4449 4018
rect 2154 3950 2304 3984
rect 2338 3950 2374 3984
rect 2408 3950 2444 3984
rect 2478 3950 2514 3984
rect 2548 3950 2584 3984
rect 2618 3950 2654 3984
rect 2688 3950 2724 3984
rect 2758 3950 2794 3984
rect 2828 3950 2864 3984
rect 2898 3950 2934 3984
rect 2968 3950 3004 3984
rect 3038 3950 3074 3984
rect 3108 3950 3144 3984
rect 3178 3950 3214 3984
rect 3248 3950 3284 3984
rect 3318 3950 3354 3984
rect 3388 3950 3424 3984
rect 3458 3950 3494 3984
rect 3528 3950 3563 3984
rect 3597 3950 3632 3984
rect 3666 3950 3701 3984
rect 3735 3950 3770 3984
rect 3804 3950 3839 3984
rect 3873 3950 3908 3984
rect 3942 3950 3977 3984
rect 4011 3950 4046 3984
rect 4080 3950 4115 3984
rect 4149 3950 4184 3984
rect 4218 3950 4253 3984
rect 4287 3950 4322 3984
rect 4356 3950 4391 3984
rect 4425 3950 4449 3984
rect 2154 3916 4449 3950
rect 2154 3882 2304 3916
rect 2338 3882 2374 3916
rect 2408 3882 2444 3916
rect 2478 3882 2514 3916
rect 2548 3882 2584 3916
rect 2618 3882 2654 3916
rect 2688 3882 2724 3916
rect 2758 3882 2794 3916
rect 2828 3882 2864 3916
rect 2898 3882 2934 3916
rect 2968 3882 3004 3916
rect 3038 3882 3074 3916
rect 3108 3882 3144 3916
rect 3178 3882 3214 3916
rect 3248 3882 3284 3916
rect 3318 3882 3354 3916
rect 3388 3882 3424 3916
rect 3458 3882 3494 3916
rect 3528 3882 3563 3916
rect 3597 3882 3632 3916
rect 3666 3882 3701 3916
rect 3735 3882 3770 3916
rect 3804 3882 3839 3916
rect 3873 3882 3908 3916
rect 3942 3882 3977 3916
rect 4011 3882 4046 3916
rect 4080 3882 4115 3916
rect 4149 3882 4184 3916
rect 4218 3882 4253 3916
rect 4287 3882 4322 3916
rect 4356 3882 4391 3916
rect 4425 3882 4449 3916
rect 2154 3848 4449 3882
rect 2154 3814 2304 3848
rect 2338 3814 2374 3848
rect 2408 3814 2444 3848
rect 2478 3814 2514 3848
rect 2548 3814 2584 3848
rect 2618 3814 2654 3848
rect 2688 3814 2724 3848
rect 2758 3814 2794 3848
rect 2828 3814 2864 3848
rect 2898 3814 2934 3848
rect 2968 3814 3004 3848
rect 3038 3814 3074 3848
rect 3108 3814 3144 3848
rect 3178 3814 3214 3848
rect 3248 3814 3284 3848
rect 3318 3814 3354 3848
rect 3388 3814 3424 3848
rect 3458 3814 3494 3848
rect 3528 3814 3563 3848
rect 3597 3814 3632 3848
rect 3666 3814 3701 3848
rect 3735 3814 3770 3848
rect 3804 3814 3839 3848
rect 3873 3814 3908 3848
rect 3942 3814 3977 3848
rect 4011 3814 4046 3848
rect 4080 3814 4115 3848
rect 4149 3814 4184 3848
rect 4218 3814 4253 3848
rect 4287 3814 4322 3848
rect 4356 3814 4391 3848
rect 4425 3814 4449 3848
rect 2154 3780 4449 3814
rect 2154 3746 2304 3780
rect 2338 3746 2374 3780
rect 2408 3746 2444 3780
rect 2478 3746 2514 3780
rect 2548 3746 2584 3780
rect 2618 3746 2654 3780
rect 2688 3746 2724 3780
rect 2758 3746 2794 3780
rect 2828 3746 2864 3780
rect 2898 3746 2934 3780
rect 2968 3746 3004 3780
rect 3038 3746 3074 3780
rect 3108 3746 3144 3780
rect 3178 3746 3214 3780
rect 3248 3746 3284 3780
rect 3318 3746 3354 3780
rect 3388 3746 3424 3780
rect 3458 3746 3494 3780
rect 3528 3746 3563 3780
rect 3597 3746 3632 3780
rect 3666 3746 3701 3780
rect 3735 3746 3770 3780
rect 3804 3746 3839 3780
rect 3873 3746 3908 3780
rect 3942 3746 3977 3780
rect 4011 3746 4046 3780
rect 4080 3746 4115 3780
rect 4149 3746 4184 3780
rect 4218 3746 4253 3780
rect 4287 3746 4322 3780
rect 4356 3746 4391 3780
rect 4425 3746 4449 3780
rect 2154 3712 4449 3746
rect 2154 3678 2304 3712
rect 2338 3678 2374 3712
rect 2408 3678 2444 3712
rect 2478 3678 2514 3712
rect 2548 3678 2584 3712
rect 2618 3678 2654 3712
rect 2688 3678 2724 3712
rect 2758 3678 2794 3712
rect 2828 3678 2864 3712
rect 2898 3678 2934 3712
rect 2968 3678 3004 3712
rect 3038 3678 3074 3712
rect 3108 3678 3144 3712
rect 3178 3678 3214 3712
rect 3248 3678 3284 3712
rect 3318 3678 3354 3712
rect 3388 3678 3424 3712
rect 3458 3678 3494 3712
rect 3528 3678 3563 3712
rect 3597 3678 3632 3712
rect 3666 3678 3701 3712
rect 3735 3678 3770 3712
rect 3804 3678 3839 3712
rect 3873 3678 3908 3712
rect 3942 3678 3977 3712
rect 4011 3678 4046 3712
rect 4080 3678 4115 3712
rect 4149 3678 4184 3712
rect 4218 3678 4253 3712
rect 4287 3678 4322 3712
rect 4356 3678 4391 3712
rect 4425 3678 4449 3712
rect 2154 3644 4449 3678
rect 2154 3610 2304 3644
rect 2338 3610 2374 3644
rect 2408 3610 2444 3644
rect 2478 3610 2514 3644
rect 2548 3610 2584 3644
rect 2618 3610 2654 3644
rect 2688 3610 2724 3644
rect 2758 3610 2794 3644
rect 2828 3610 2864 3644
rect 2898 3610 2934 3644
rect 2968 3610 3004 3644
rect 3038 3610 3074 3644
rect 3108 3610 3144 3644
rect 3178 3610 3214 3644
rect 3248 3610 3284 3644
rect 3318 3610 3354 3644
rect 3388 3610 3424 3644
rect 3458 3610 3494 3644
rect 3528 3610 3563 3644
rect 3597 3610 3632 3644
rect 3666 3610 3701 3644
rect 3735 3610 3770 3644
rect 3804 3610 3839 3644
rect 3873 3610 3908 3644
rect 3942 3610 3977 3644
rect 4011 3610 4046 3644
rect 4080 3610 4115 3644
rect 4149 3610 4184 3644
rect 4218 3610 4253 3644
rect 4287 3610 4322 3644
rect 4356 3610 4391 3644
rect 4425 3610 4449 3644
rect 2154 3576 4449 3610
rect 2154 3542 2304 3576
rect 2338 3542 2374 3576
rect 2408 3542 2444 3576
rect 2478 3542 2514 3576
rect 2548 3542 2584 3576
rect 2618 3542 2654 3576
rect 2688 3542 2724 3576
rect 2758 3542 2794 3576
rect 2828 3542 2864 3576
rect 2898 3542 2934 3576
rect 2968 3542 3004 3576
rect 3038 3542 3074 3576
rect 3108 3542 3144 3576
rect 3178 3542 3214 3576
rect 3248 3542 3284 3576
rect 3318 3542 3354 3576
rect 3388 3542 3424 3576
rect 3458 3542 3494 3576
rect 3528 3542 3563 3576
rect 3597 3542 3632 3576
rect 3666 3542 3701 3576
rect 3735 3542 3770 3576
rect 3804 3542 3839 3576
rect 3873 3542 3908 3576
rect 3942 3542 3977 3576
rect 4011 3542 4046 3576
rect 4080 3542 4115 3576
rect 4149 3542 4184 3576
rect 4218 3542 4253 3576
rect 4287 3542 4322 3576
rect 4356 3542 4391 3576
rect 4425 3542 4449 3576
rect 11076 4504 11698 4564
rect 11076 4470 11159 4504
rect 11193 4470 11231 4504
rect 11265 4470 11303 4504
rect 11337 4470 11375 4504
rect 11409 4470 11447 4504
rect 11481 4470 11519 4504
rect 11553 4470 11591 4504
rect 11625 4470 11663 4504
rect 11697 4470 11698 4504
rect 11076 4434 11698 4470
rect 11076 4400 11159 4434
rect 11193 4400 11231 4434
rect 11265 4400 11303 4434
rect 11337 4400 11375 4434
rect 11409 4400 11447 4434
rect 11481 4400 11519 4434
rect 11553 4400 11591 4434
rect 11625 4400 11663 4434
rect 11697 4400 11698 4434
rect 11076 4364 11698 4400
rect 11076 4330 11159 4364
rect 11193 4330 11231 4364
rect 11265 4330 11303 4364
rect 11337 4330 11375 4364
rect 11409 4330 11447 4364
rect 11481 4330 11519 4364
rect 11553 4330 11591 4364
rect 11625 4330 11663 4364
rect 11697 4330 11698 4364
rect 11076 4294 11698 4330
rect 11076 4260 11159 4294
rect 11193 4260 11231 4294
rect 11265 4260 11303 4294
rect 11337 4260 11375 4294
rect 11409 4260 11447 4294
rect 11481 4260 11519 4294
rect 11553 4260 11591 4294
rect 11625 4260 11663 4294
rect 11697 4260 11698 4294
rect 11076 4223 11698 4260
rect 11076 4189 11159 4223
rect 11193 4189 11231 4223
rect 11265 4189 11303 4223
rect 11337 4189 11375 4223
rect 11409 4189 11447 4223
rect 11481 4189 11519 4223
rect 11553 4189 11591 4223
rect 11625 4189 11663 4223
rect 11697 4189 11698 4223
rect 11076 4152 11698 4189
rect 11076 4118 11159 4152
rect 11193 4118 11231 4152
rect 11265 4118 11303 4152
rect 11337 4118 11375 4152
rect 11409 4118 11447 4152
rect 11481 4118 11519 4152
rect 11553 4118 11591 4152
rect 11625 4118 11663 4152
rect 11697 4118 11698 4152
rect 11076 4081 11698 4118
rect 11076 4047 11159 4081
rect 11193 4047 11231 4081
rect 11265 4047 11303 4081
rect 11337 4047 11375 4081
rect 11409 4047 11447 4081
rect 11481 4047 11519 4081
rect 11553 4047 11591 4081
rect 11625 4047 11663 4081
rect 11697 4047 11698 4081
rect 11076 4010 11698 4047
rect 11076 3976 11159 4010
rect 11193 3976 11231 4010
rect 11265 3976 11303 4010
rect 11337 3976 11375 4010
rect 11409 3976 11447 4010
rect 11481 3976 11519 4010
rect 11553 3976 11591 4010
rect 11625 3976 11663 4010
rect 11697 3976 11698 4010
rect 11076 3939 11698 3976
rect 11076 3905 11159 3939
rect 11193 3905 11231 3939
rect 11265 3905 11303 3939
rect 11337 3905 11375 3939
rect 11409 3905 11447 3939
rect 11481 3905 11519 3939
rect 11553 3905 11591 3939
rect 11625 3905 11663 3939
rect 11697 3905 11698 3939
rect 11076 3868 11698 3905
rect 11076 3834 11159 3868
rect 11193 3834 11231 3868
rect 11265 3834 11303 3868
rect 11337 3834 11375 3868
rect 11409 3834 11447 3868
rect 11481 3834 11519 3868
rect 11553 3834 11591 3868
rect 11625 3834 11663 3868
rect 11697 3834 11698 3868
rect 11076 3797 11698 3834
rect 11076 3763 11159 3797
rect 11193 3763 11231 3797
rect 11265 3763 11303 3797
rect 11337 3763 11375 3797
rect 11409 3763 11447 3797
rect 11481 3763 11519 3797
rect 11553 3763 11591 3797
rect 11625 3763 11663 3797
rect 11697 3763 11698 3797
rect 11076 3726 11698 3763
rect 11076 3692 11159 3726
rect 11193 3692 11231 3726
rect 11265 3692 11303 3726
rect 11337 3692 11375 3726
rect 11409 3692 11447 3726
rect 11481 3692 11519 3726
rect 11553 3692 11591 3726
rect 11625 3692 11663 3726
rect 11697 3692 11698 3726
rect 11076 3655 11698 3692
rect 11076 3621 11159 3655
rect 11193 3621 11231 3655
rect 11265 3621 11303 3655
rect 11337 3621 11375 3655
rect 11409 3621 11447 3655
rect 11481 3621 11519 3655
rect 11553 3621 11591 3655
rect 11625 3621 11663 3655
rect 11697 3621 11698 3655
rect 11076 3571 11698 3621
rect 2154 3508 4449 3542
rect 2154 3474 2304 3508
rect 2338 3474 2374 3508
rect 2408 3474 2444 3508
rect 2478 3474 2514 3508
rect 2548 3474 2584 3508
rect 2618 3474 2654 3508
rect 2688 3474 2724 3508
rect 2758 3474 2794 3508
rect 2828 3474 2864 3508
rect 2898 3474 2934 3508
rect 2968 3474 3004 3508
rect 3038 3474 3074 3508
rect 3108 3474 3144 3508
rect 3178 3474 3214 3508
rect 3248 3474 3284 3508
rect 3318 3474 3354 3508
rect 3388 3474 3424 3508
rect 3458 3474 3494 3508
rect 3528 3474 3563 3508
rect 3597 3474 3632 3508
rect 3666 3474 3701 3508
rect 3735 3474 3770 3508
rect 3804 3474 3839 3508
rect 3873 3474 3908 3508
rect 3942 3474 3977 3508
rect 4011 3474 4046 3508
rect 4080 3474 4115 3508
rect 4149 3474 4184 3508
rect 4218 3474 4253 3508
rect 4287 3474 4322 3508
rect 4356 3474 4391 3508
rect 4425 3474 4449 3508
rect 2154 3440 4449 3474
rect 2154 3406 2304 3440
rect 2338 3406 2374 3440
rect 2408 3406 2444 3440
rect 2478 3406 2514 3440
rect 2548 3406 2584 3440
rect 2618 3406 2654 3440
rect 2688 3406 2724 3440
rect 2758 3406 2794 3440
rect 2828 3406 2864 3440
rect 2898 3406 2934 3440
rect 2968 3406 3004 3440
rect 3038 3406 3074 3440
rect 3108 3406 3144 3440
rect 3178 3406 3214 3440
rect 3248 3406 3284 3440
rect 3318 3406 3354 3440
rect 3388 3406 3424 3440
rect 3458 3406 3494 3440
rect 3528 3406 3563 3440
rect 3597 3406 3632 3440
rect 3666 3406 3701 3440
rect 3735 3406 3770 3440
rect 3804 3406 3839 3440
rect 3873 3406 3908 3440
rect 3942 3406 3977 3440
rect 4011 3406 4046 3440
rect 4080 3406 4115 3440
rect 4149 3406 4184 3440
rect 4218 3406 4253 3440
rect 4287 3406 4322 3440
rect 4356 3406 4391 3440
rect 4425 3406 4449 3440
rect 2154 3372 4449 3406
rect 4505 3537 4529 3571
rect 4563 3537 4598 3571
rect 4632 3537 4667 3571
rect 4701 3537 4736 3571
rect 4770 3537 4805 3571
rect 4839 3537 4874 3571
rect 4908 3537 4943 3571
rect 4977 3537 5012 3571
rect 5046 3537 5081 3571
rect 5115 3537 5150 3571
rect 5184 3537 5219 3571
rect 5253 3537 5288 3571
rect 5322 3537 5357 3571
rect 5391 3537 5426 3571
rect 5460 3537 5495 3571
rect 5529 3537 5564 3571
rect 5598 3537 5633 3571
rect 5667 3537 5702 3571
rect 5736 3537 5771 3571
rect 5805 3537 5840 3571
rect 5874 3537 5909 3571
rect 5943 3537 5978 3571
rect 6012 3537 6047 3571
rect 6081 3537 6116 3571
rect 6150 3537 6185 3571
rect 6219 3537 6254 3571
rect 6288 3537 6323 3571
rect 6357 3537 6392 3571
rect 6426 3537 6461 3571
rect 6495 3537 6530 3571
rect 6564 3537 6599 3571
rect 6633 3537 6668 3571
rect 6702 3537 6737 3571
rect 6771 3537 6806 3571
rect 6840 3537 6875 3571
rect 6909 3537 6944 3571
rect 6978 3537 7013 3571
rect 7047 3537 7082 3571
rect 7116 3537 7151 3571
rect 7185 3537 7220 3571
rect 4505 3503 7220 3537
rect 4505 3469 4529 3503
rect 4563 3469 4598 3503
rect 4632 3469 4667 3503
rect 4701 3469 4736 3503
rect 4770 3469 4805 3503
rect 4839 3469 4874 3503
rect 4908 3469 4943 3503
rect 4977 3469 5012 3503
rect 5046 3469 5081 3503
rect 5115 3469 5150 3503
rect 5184 3469 5219 3503
rect 5253 3469 5288 3503
rect 5322 3469 5357 3503
rect 5391 3469 5426 3503
rect 5460 3469 5495 3503
rect 5529 3469 5564 3503
rect 5598 3469 5633 3503
rect 5667 3469 5702 3503
rect 5736 3469 5771 3503
rect 5805 3469 5840 3503
rect 5874 3469 5909 3503
rect 5943 3469 5978 3503
rect 6012 3469 6047 3503
rect 6081 3469 6116 3503
rect 6150 3469 6185 3503
rect 6219 3469 6254 3503
rect 6288 3469 6323 3503
rect 6357 3469 6392 3503
rect 6426 3469 6461 3503
rect 6495 3469 6530 3503
rect 6564 3469 6599 3503
rect 6633 3469 6668 3503
rect 6702 3469 6737 3503
rect 6771 3469 6806 3503
rect 6840 3469 6875 3503
rect 6909 3469 6944 3503
rect 6978 3469 7013 3503
rect 7047 3469 7082 3503
rect 7116 3469 7151 3503
rect 7185 3469 7220 3503
rect 4505 3435 7220 3469
rect 4505 3401 4529 3435
rect 4563 3401 4598 3435
rect 4632 3401 4667 3435
rect 4701 3401 4736 3435
rect 4770 3401 4805 3435
rect 4839 3401 4874 3435
rect 4908 3401 4943 3435
rect 4977 3401 5012 3435
rect 5046 3401 5081 3435
rect 5115 3401 5150 3435
rect 5184 3401 5219 3435
rect 5253 3401 5288 3435
rect 5322 3401 5357 3435
rect 5391 3401 5426 3435
rect 5460 3401 5495 3435
rect 5529 3401 5564 3435
rect 5598 3401 5633 3435
rect 5667 3401 5702 3435
rect 5736 3401 5771 3435
rect 5805 3401 5840 3435
rect 5874 3401 5909 3435
rect 5943 3401 5978 3435
rect 6012 3401 6047 3435
rect 6081 3401 6116 3435
rect 6150 3401 6185 3435
rect 6219 3401 6254 3435
rect 6288 3401 6323 3435
rect 6357 3401 6392 3435
rect 6426 3401 6461 3435
rect 6495 3401 6530 3435
rect 6564 3401 6599 3435
rect 6633 3401 6668 3435
rect 6702 3401 6737 3435
rect 6771 3401 6806 3435
rect 6840 3401 6875 3435
rect 6909 3401 6944 3435
rect 6978 3401 7013 3435
rect 7047 3401 7082 3435
rect 7116 3401 7151 3435
rect 7185 3401 7220 3435
rect 11674 3401 11698 3571
rect 2154 3338 2304 3372
rect 2338 3338 2374 3372
rect 2408 3338 2444 3372
rect 2478 3338 2514 3372
rect 2548 3338 2584 3372
rect 2618 3338 2654 3372
rect 2688 3338 2724 3372
rect 2758 3338 2794 3372
rect 2828 3338 2864 3372
rect 2898 3338 2934 3372
rect 2968 3338 3004 3372
rect 3038 3338 3074 3372
rect 3108 3338 3144 3372
rect 3178 3338 3214 3372
rect 3248 3338 3284 3372
rect 3318 3338 3354 3372
rect 3388 3338 3424 3372
rect 3458 3338 3494 3372
rect 3528 3338 3563 3372
rect 3597 3338 3632 3372
rect 3666 3338 3701 3372
rect 3735 3338 3770 3372
rect 3804 3338 3839 3372
rect 3873 3338 3908 3372
rect 3942 3338 3977 3372
rect 4011 3338 4046 3372
rect 4080 3338 4115 3372
rect 4149 3338 4184 3372
rect 4218 3338 4253 3372
rect 4287 3338 4322 3372
rect 4356 3338 4391 3372
rect 4425 3338 4449 3372
rect 2154 3304 4449 3338
rect 2154 3270 2304 3304
rect 2338 3270 2374 3304
rect 2408 3270 2444 3304
rect 2478 3270 2514 3304
rect 2548 3270 2584 3304
rect 2618 3270 2654 3304
rect 2688 3270 2724 3304
rect 2758 3270 2794 3304
rect 2828 3270 2864 3304
rect 2898 3270 2934 3304
rect 2968 3270 3004 3304
rect 3038 3270 3074 3304
rect 3108 3270 3144 3304
rect 3178 3270 3214 3304
rect 3248 3270 3284 3304
rect 3318 3270 3354 3304
rect 3388 3270 3424 3304
rect 3458 3270 3494 3304
rect 3528 3270 3563 3304
rect 3597 3270 3632 3304
rect 3666 3270 3701 3304
rect 3735 3270 3770 3304
rect 3804 3270 3839 3304
rect 3873 3270 3908 3304
rect 3942 3270 3977 3304
rect 4011 3270 4046 3304
rect 4080 3270 4115 3304
rect 4149 3270 4184 3304
rect 4218 3270 4253 3304
rect 4287 3270 4322 3304
rect 4356 3270 4391 3304
rect 4425 3270 4449 3304
rect 2154 3236 4449 3270
rect 2154 3202 2304 3236
rect 2338 3202 2374 3236
rect 2408 3202 2444 3236
rect 2478 3202 2514 3236
rect 2548 3202 2584 3236
rect 2618 3202 2654 3236
rect 2688 3202 2724 3236
rect 2758 3202 2794 3236
rect 2828 3202 2864 3236
rect 2898 3202 2934 3236
rect 2968 3202 3004 3236
rect 3038 3202 3074 3236
rect 3108 3202 3144 3236
rect 3178 3202 3214 3236
rect 3248 3202 3284 3236
rect 3318 3202 3354 3236
rect 3388 3202 3424 3236
rect 3458 3202 3494 3236
rect 3528 3202 3563 3236
rect 3597 3202 3632 3236
rect 3666 3202 3701 3236
rect 3735 3202 3770 3236
rect 3804 3202 3839 3236
rect 3873 3202 3908 3236
rect 3942 3202 3977 3236
rect 4011 3202 4046 3236
rect 4080 3202 4115 3236
rect 4149 3202 4184 3236
rect 4218 3202 4253 3236
rect 4287 3202 4322 3236
rect 4356 3202 4391 3236
rect 4425 3202 4449 3236
rect 2154 3168 4449 3202
rect 2154 3134 2304 3168
rect 2338 3134 2374 3168
rect 2408 3134 2444 3168
rect 2478 3134 2514 3168
rect 2548 3134 2584 3168
rect 2618 3134 2654 3168
rect 2688 3134 2724 3168
rect 2758 3134 2794 3168
rect 2828 3134 2864 3168
rect 2898 3134 2934 3168
rect 2968 3134 3004 3168
rect 3038 3134 3074 3168
rect 3108 3134 3144 3168
rect 3178 3134 3214 3168
rect 3248 3134 3284 3168
rect 3318 3134 3354 3168
rect 3388 3134 3424 3168
rect 3458 3134 3494 3168
rect 3528 3134 3563 3168
rect 3597 3134 3632 3168
rect 3666 3134 3701 3168
rect 3735 3134 3770 3168
rect 3804 3134 3839 3168
rect 3873 3134 3908 3168
rect 3942 3134 3977 3168
rect 4011 3134 4046 3168
rect 4080 3134 4115 3168
rect 4149 3134 4184 3168
rect 4218 3134 4253 3168
rect 4287 3134 4322 3168
rect 4356 3134 4391 3168
rect 4425 3134 4449 3168
rect 2154 3100 4449 3134
rect 2154 3066 2304 3100
rect 2338 3066 2374 3100
rect 2408 3066 2444 3100
rect 2478 3066 2514 3100
rect 2548 3066 2584 3100
rect 2618 3066 2654 3100
rect 2688 3066 2724 3100
rect 2758 3066 2794 3100
rect 2828 3066 2864 3100
rect 2898 3066 2934 3100
rect 2968 3066 3004 3100
rect 3038 3066 3074 3100
rect 3108 3066 3144 3100
rect 3178 3066 3214 3100
rect 3248 3066 3284 3100
rect 3318 3066 3354 3100
rect 3388 3066 3424 3100
rect 3458 3066 3494 3100
rect 3528 3066 3563 3100
rect 3597 3066 3632 3100
rect 3666 3066 3701 3100
rect 3735 3066 3770 3100
rect 3804 3066 3839 3100
rect 3873 3066 3908 3100
rect 3942 3066 3977 3100
rect 4011 3066 4046 3100
rect 4080 3066 4115 3100
rect 4149 3066 4184 3100
rect 4218 3066 4253 3100
rect 4287 3066 4322 3100
rect 4356 3066 4391 3100
rect 4425 3066 4449 3100
rect 2154 3032 4449 3066
rect 2154 2998 2304 3032
rect 2338 2998 2374 3032
rect 2408 2998 2444 3032
rect 2478 2998 2514 3032
rect 2548 2998 2584 3032
rect 2618 2998 2654 3032
rect 2688 2998 2724 3032
rect 2758 2998 2794 3032
rect 2828 2998 2864 3032
rect 2898 2998 2934 3032
rect 2968 2998 3004 3032
rect 3038 2998 3074 3032
rect 3108 2998 3144 3032
rect 3178 2998 3214 3032
rect 3248 2998 3284 3032
rect 3318 2998 3354 3032
rect 3388 2998 3424 3032
rect 3458 2998 3494 3032
rect 3528 2998 3563 3032
rect 3597 2998 3632 3032
rect 3666 2998 3701 3032
rect 3735 2998 3770 3032
rect 3804 2998 3839 3032
rect 3873 2998 3908 3032
rect 3942 2998 3977 3032
rect 4011 2998 4046 3032
rect 4080 2998 4115 3032
rect 4149 2998 4184 3032
rect 4218 2998 4253 3032
rect 4287 2998 4322 3032
rect 4356 2998 4391 3032
rect 4425 2998 4449 3032
rect 2154 2964 4449 2998
rect 2154 2930 2304 2964
rect 2338 2930 2374 2964
rect 2408 2930 2444 2964
rect 2478 2930 2514 2964
rect 2548 2930 2584 2964
rect 2618 2930 2654 2964
rect 2688 2930 2724 2964
rect 2758 2930 2794 2964
rect 2828 2930 2864 2964
rect 2898 2930 2934 2964
rect 2968 2930 3004 2964
rect 3038 2930 3074 2964
rect 3108 2930 3144 2964
rect 3178 2930 3214 2964
rect 3248 2930 3284 2964
rect 3318 2930 3354 2964
rect 3388 2930 3424 2964
rect 3458 2930 3494 2964
rect 3528 2930 3563 2964
rect 3597 2930 3632 2964
rect 3666 2930 3701 2964
rect 3735 2930 3770 2964
rect 3804 2930 3839 2964
rect 3873 2930 3908 2964
rect 3942 2930 3977 2964
rect 4011 2930 4046 2964
rect 4080 2930 4115 2964
rect 4149 2930 4184 2964
rect 4218 2930 4253 2964
rect 4287 2930 4322 2964
rect 4356 2930 4391 2964
rect 4425 2930 4449 2964
rect 2154 2896 4449 2930
rect 2154 2862 2304 2896
rect 2338 2862 2374 2896
rect 2408 2862 2444 2896
rect 2478 2862 2514 2896
rect 2548 2862 2584 2896
rect 2618 2862 2654 2896
rect 2688 2862 2724 2896
rect 2758 2862 2794 2896
rect 2828 2862 2864 2896
rect 2898 2862 2934 2896
rect 2968 2862 3004 2896
rect 3038 2862 3074 2896
rect 3108 2862 3144 2896
rect 3178 2862 3214 2896
rect 3248 2862 3284 2896
rect 3318 2862 3354 2896
rect 3388 2862 3424 2896
rect 3458 2862 3494 2896
rect 3528 2862 3563 2896
rect 3597 2862 3632 2896
rect 3666 2862 3701 2896
rect 3735 2862 3770 2896
rect 3804 2862 3839 2896
rect 3873 2862 3908 2896
rect 3942 2862 3977 2896
rect 4011 2862 4046 2896
rect 4080 2862 4115 2896
rect 4149 2862 4184 2896
rect 4218 2862 4253 2896
rect 4287 2862 4322 2896
rect 4356 2862 4391 2896
rect 4425 2862 4449 2896
rect 2154 2828 4449 2862
rect 2154 2794 2304 2828
rect 2338 2794 2374 2828
rect 2408 2794 2444 2828
rect 2478 2794 2514 2828
rect 2548 2794 2584 2828
rect 2618 2794 2654 2828
rect 2688 2794 2724 2828
rect 2758 2794 2794 2828
rect 2828 2794 2864 2828
rect 2898 2794 2934 2828
rect 2968 2794 3004 2828
rect 3038 2794 3074 2828
rect 3108 2794 3144 2828
rect 3178 2794 3214 2828
rect 3248 2794 3284 2828
rect 3318 2794 3354 2828
rect 3388 2794 3424 2828
rect 3458 2794 3494 2828
rect 3528 2794 3563 2828
rect 3597 2794 3632 2828
rect 3666 2794 3701 2828
rect 3735 2794 3770 2828
rect 3804 2794 3839 2828
rect 3873 2794 3908 2828
rect 3942 2794 3977 2828
rect 4011 2794 4046 2828
rect 4080 2794 4115 2828
rect 4149 2794 4184 2828
rect 4218 2794 4253 2828
rect 4287 2794 4322 2828
rect 4356 2794 4391 2828
rect 4425 2794 4449 2828
rect 2154 2760 4449 2794
rect 2154 2726 2304 2760
rect 2338 2726 2374 2760
rect 2408 2726 2444 2760
rect 2478 2726 2514 2760
rect 2548 2726 2584 2760
rect 2618 2726 2654 2760
rect 2688 2726 2724 2760
rect 2758 2726 2794 2760
rect 2828 2726 2864 2760
rect 2898 2726 2934 2760
rect 2968 2726 3004 2760
rect 3038 2726 3074 2760
rect 3108 2726 3144 2760
rect 3178 2726 3214 2760
rect 3248 2726 3284 2760
rect 3318 2726 3354 2760
rect 3388 2726 3424 2760
rect 3458 2726 3494 2760
rect 3528 2726 3563 2760
rect 3597 2726 3632 2760
rect 3666 2726 3701 2760
rect 3735 2726 3770 2760
rect 3804 2726 3839 2760
rect 3873 2726 3908 2760
rect 3942 2726 3977 2760
rect 4011 2726 4046 2760
rect 4080 2726 4115 2760
rect 4149 2726 4184 2760
rect 4218 2726 4253 2760
rect 4287 2726 4322 2760
rect 4356 2726 4391 2760
rect 4425 2726 4449 2760
rect 2154 2692 4449 2726
rect 2154 2658 2304 2692
rect 2338 2658 2374 2692
rect 2408 2658 2444 2692
rect 2478 2658 2514 2692
rect 2548 2658 2584 2692
rect 2618 2658 2654 2692
rect 2688 2658 2724 2692
rect 2758 2658 2794 2692
rect 2828 2658 2864 2692
rect 2898 2658 2934 2692
rect 2968 2658 3004 2692
rect 3038 2658 3074 2692
rect 3108 2658 3144 2692
rect 3178 2658 3214 2692
rect 3248 2658 3284 2692
rect 3318 2658 3354 2692
rect 3388 2658 3424 2692
rect 3458 2658 3494 2692
rect 3528 2658 3563 2692
rect 3597 2658 3632 2692
rect 3666 2658 3701 2692
rect 3735 2658 3770 2692
rect 3804 2658 3839 2692
rect 3873 2658 3908 2692
rect 3942 2658 3977 2692
rect 4011 2658 4046 2692
rect 4080 2658 4115 2692
rect 4149 2658 4184 2692
rect 4218 2658 4253 2692
rect 4287 2658 4322 2692
rect 4356 2658 4391 2692
rect 4425 2658 4449 2692
rect 2154 2624 4449 2658
rect 2154 2590 2304 2624
rect 2338 2590 2374 2624
rect 2408 2590 2444 2624
rect 2478 2590 2514 2624
rect 2548 2590 2584 2624
rect 2618 2590 2654 2624
rect 2688 2590 2724 2624
rect 2758 2590 2794 2624
rect 2828 2590 2864 2624
rect 2898 2590 2934 2624
rect 2968 2590 3004 2624
rect 3038 2590 3074 2624
rect 3108 2590 3144 2624
rect 3178 2590 3214 2624
rect 3248 2590 3284 2624
rect 3318 2590 3354 2624
rect 3388 2590 3424 2624
rect 3458 2590 3494 2624
rect 3528 2590 3563 2624
rect 3597 2590 3632 2624
rect 3666 2590 3701 2624
rect 3735 2590 3770 2624
rect 3804 2590 3839 2624
rect 3873 2590 3908 2624
rect 3942 2590 3977 2624
rect 4011 2590 4046 2624
rect 4080 2590 4115 2624
rect 4149 2590 4184 2624
rect 4218 2590 4253 2624
rect 4287 2590 4322 2624
rect 4356 2590 4391 2624
rect 4425 2590 4449 2624
rect 2154 2556 4449 2590
rect 2154 2522 2304 2556
rect 2338 2522 2374 2556
rect 2408 2522 2444 2556
rect 2478 2522 2514 2556
rect 2548 2522 2584 2556
rect 2618 2522 2654 2556
rect 2688 2522 2724 2556
rect 2758 2522 2794 2556
rect 2828 2522 2864 2556
rect 2898 2522 2934 2556
rect 2968 2522 3004 2556
rect 3038 2522 3074 2556
rect 3108 2522 3144 2556
rect 3178 2522 3214 2556
rect 3248 2522 3284 2556
rect 3318 2522 3354 2556
rect 3388 2522 3424 2556
rect 3458 2522 3494 2556
rect 3528 2522 3563 2556
rect 3597 2522 3632 2556
rect 3666 2522 3701 2556
rect 3735 2522 3770 2556
rect 3804 2522 3839 2556
rect 3873 2522 3908 2556
rect 3942 2522 3977 2556
rect 4011 2522 4046 2556
rect 4080 2522 4115 2556
rect 4149 2522 4184 2556
rect 4218 2522 4253 2556
rect 4287 2522 4322 2556
rect 4356 2522 4391 2556
rect 4425 2522 4449 2556
rect 2154 2488 4449 2522
rect 2154 2454 2304 2488
rect 2338 2454 2374 2488
rect 2408 2454 2444 2488
rect 2478 2454 2514 2488
rect 2548 2454 2584 2488
rect 2618 2454 2654 2488
rect 2688 2454 2724 2488
rect 2758 2454 2794 2488
rect 2828 2454 2864 2488
rect 2898 2454 2934 2488
rect 2968 2454 3004 2488
rect 3038 2454 3074 2488
rect 3108 2454 3144 2488
rect 3178 2454 3214 2488
rect 3248 2454 3284 2488
rect 3318 2454 3354 2488
rect 3388 2454 3424 2488
rect 3458 2454 3494 2488
rect 3528 2454 3563 2488
rect 3597 2454 3632 2488
rect 3666 2454 3701 2488
rect 3735 2454 3770 2488
rect 3804 2454 3839 2488
rect 3873 2454 3908 2488
rect 3942 2454 3977 2488
rect 4011 2454 4046 2488
rect 4080 2454 4115 2488
rect 4149 2454 4184 2488
rect 4218 2454 4253 2488
rect 4287 2454 4322 2488
rect 4356 2454 4391 2488
rect 4425 2454 4449 2488
rect 2154 2420 4449 2454
rect 2154 2386 2304 2420
rect 2338 2386 2374 2420
rect 2408 2386 2444 2420
rect 2478 2386 2514 2420
rect 2548 2386 2584 2420
rect 2618 2386 2654 2420
rect 2688 2386 2724 2420
rect 2758 2386 2794 2420
rect 2828 2386 2864 2420
rect 2898 2386 2934 2420
rect 2968 2386 3004 2420
rect 3038 2386 3074 2420
rect 3108 2386 3144 2420
rect 3178 2386 3214 2420
rect 3248 2386 3284 2420
rect 3318 2386 3354 2420
rect 3388 2386 3424 2420
rect 3458 2386 3494 2420
rect 3528 2386 3563 2420
rect 3597 2386 3632 2420
rect 3666 2386 3701 2420
rect 3735 2386 3770 2420
rect 3804 2386 3839 2420
rect 3873 2386 3908 2420
rect 3942 2386 3977 2420
rect 4011 2386 4046 2420
rect 4080 2386 4115 2420
rect 4149 2386 4184 2420
rect 4218 2386 4253 2420
rect 4287 2386 4322 2420
rect 4356 2386 4391 2420
rect 4425 2386 4449 2420
rect 2154 2352 4449 2386
rect 2154 2319 2304 2352
rect -214 2294 -161 2303
rect -2750 2269 -161 2294
rect -127 2269 -89 2303
rect -55 2269 -17 2303
rect 17 2269 55 2303
rect 89 2269 127 2303
rect 161 2269 199 2303
rect 233 2269 271 2303
rect 305 2269 433 2303
rect -2750 2204 433 2269
rect 2148 2318 2304 2319
rect 2338 2318 2374 2352
rect 2408 2318 2444 2352
rect 2478 2318 2514 2352
rect 2548 2318 2584 2352
rect 2618 2318 2654 2352
rect 2688 2318 2724 2352
rect 2758 2318 2794 2352
rect 2828 2318 2864 2352
rect 2898 2318 2934 2352
rect 2968 2318 3004 2352
rect 3038 2318 3074 2352
rect 3108 2318 3144 2352
rect 3178 2318 3214 2352
rect 3248 2318 3284 2352
rect 3318 2318 3354 2352
rect 3388 2318 3424 2352
rect 3458 2318 3494 2352
rect 3528 2318 3563 2352
rect 3597 2318 3632 2352
rect 3666 2318 3701 2352
rect 3735 2318 3770 2352
rect 3804 2318 3839 2352
rect 3873 2318 3908 2352
rect 3942 2318 3977 2352
rect 4011 2318 4046 2352
rect 4080 2318 4115 2352
rect 4149 2318 4184 2352
rect 4218 2318 4253 2352
rect 4287 2318 4322 2352
rect 4356 2318 4391 2352
rect 4425 2318 4449 2352
rect 2148 2284 4449 2318
rect 2148 2250 2304 2284
rect 2338 2250 2374 2284
rect 2408 2250 2444 2284
rect 2478 2250 2514 2284
rect 2548 2250 2584 2284
rect 2618 2250 2654 2284
rect 2688 2250 2724 2284
rect 2758 2250 2794 2284
rect 2828 2250 2864 2284
rect 2898 2250 2934 2284
rect 2968 2250 3004 2284
rect 3038 2250 3074 2284
rect 3108 2250 3144 2284
rect 3178 2250 3214 2284
rect 3248 2250 3284 2284
rect 3318 2250 3354 2284
rect 3388 2250 3424 2284
rect 3458 2250 3494 2284
rect 3528 2250 3563 2284
rect 3597 2250 3632 2284
rect 3666 2250 3701 2284
rect 3735 2250 3770 2284
rect 3804 2250 3839 2284
rect 3873 2250 3908 2284
rect 3942 2250 3977 2284
rect 4011 2250 4046 2284
rect 4080 2250 4115 2284
rect 4149 2250 4184 2284
rect 4218 2250 4253 2284
rect 4287 2250 4322 2284
rect 4356 2250 4391 2284
rect 4425 2250 4449 2284
rect 2148 2204 4449 2250
rect -2750 2193 529 2204
rect 2094 2193 4449 2204
rect -2750 2159 -2726 2193
rect -2692 2159 -2656 2193
rect -2622 2159 -2586 2193
rect -2552 2159 -2517 2193
rect -2483 2159 -2448 2193
rect -2414 2159 -2379 2193
rect -2345 2159 -2310 2193
rect -2276 2159 -2241 2193
rect -2207 2159 -2172 2193
rect -2138 2159 -2103 2193
rect -2069 2159 -2034 2193
rect -2000 2159 -1965 2193
rect -1931 2159 -1896 2193
rect -1862 2159 -1827 2193
rect -1793 2159 -1758 2193
rect -1724 2159 -1689 2193
rect -1655 2159 -1620 2193
rect -1586 2159 -1551 2193
rect -1517 2159 -1482 2193
rect -1448 2159 -1413 2193
rect -1379 2159 -1344 2193
rect -1310 2159 -1275 2193
rect -1241 2159 -1206 2193
rect -1172 2159 -1137 2193
rect -1103 2159 -1068 2193
rect -1034 2159 -999 2193
rect -965 2159 -930 2193
rect -896 2159 -861 2193
rect -827 2159 -792 2193
rect -758 2159 -723 2193
rect -689 2159 -654 2193
rect -620 2159 -585 2193
rect -551 2159 -516 2193
rect -482 2159 -447 2193
rect -413 2159 -378 2193
rect -344 2159 -309 2193
rect -275 2159 -240 2193
rect -206 2159 -171 2193
rect -137 2159 -102 2193
rect -68 2159 -33 2193
rect 1 2159 36 2193
rect 70 2159 105 2193
rect 139 2159 174 2193
rect 208 2159 243 2193
rect 277 2159 2298 2193
rect 2332 2159 2368 2193
rect 2402 2159 2438 2193
rect 2472 2159 2508 2193
rect 2542 2159 2578 2193
rect 2612 2159 2648 2193
rect 2682 2159 2718 2193
rect 2752 2159 2788 2193
rect 2822 2159 2858 2193
rect 2892 2159 2928 2193
rect 2962 2159 2998 2193
rect 3032 2159 3068 2193
rect 3102 2159 3138 2193
rect 3172 2159 3208 2193
rect 3242 2159 3278 2193
rect 3312 2159 3348 2193
rect 3382 2159 3418 2193
rect 3452 2159 3488 2193
rect 3522 2159 3558 2193
rect 3592 2159 3628 2193
rect 3662 2159 3698 2193
rect 3732 2159 3768 2193
rect 3802 2159 3838 2193
rect 3872 2159 3908 2193
rect 3942 2159 3977 2193
rect 4011 2159 4046 2193
rect 4080 2159 4115 2193
rect 4149 2159 4184 2193
rect 4218 2159 4253 2193
rect 4287 2159 4322 2193
rect 4356 2159 4391 2193
rect 4425 2159 4449 2193
rect -2750 2125 4449 2159
rect -2750 2091 -2726 2125
rect -2692 2091 -2656 2125
rect -2622 2091 -2586 2125
rect -2552 2091 -2517 2125
rect -2483 2091 -2448 2125
rect -2414 2091 -2379 2125
rect -2345 2091 -2310 2125
rect -2276 2091 -2241 2125
rect -2207 2091 -2172 2125
rect -2138 2091 -2103 2125
rect -2069 2091 -2034 2125
rect -2000 2091 -1965 2125
rect -1931 2091 -1896 2125
rect -1862 2091 -1827 2125
rect -1793 2091 -1758 2125
rect -1724 2091 -1689 2125
rect -1655 2091 -1620 2125
rect -1586 2091 -1551 2125
rect -1517 2091 -1482 2125
rect -1448 2091 -1413 2125
rect -1379 2091 -1344 2125
rect -1310 2091 -1275 2125
rect -1241 2091 -1206 2125
rect -1172 2091 -1137 2125
rect -1103 2091 -1068 2125
rect -1034 2091 -999 2125
rect -965 2091 -930 2125
rect -896 2091 -861 2125
rect -827 2091 -792 2125
rect -758 2091 -723 2125
rect -689 2091 -654 2125
rect -620 2091 -585 2125
rect -551 2091 -516 2125
rect -482 2091 -447 2125
rect -413 2091 -378 2125
rect -344 2091 -309 2125
rect -275 2091 -240 2125
rect -206 2091 -171 2125
rect -137 2091 -102 2125
rect -68 2091 -33 2125
rect 1 2091 36 2125
rect 70 2091 105 2125
rect 139 2091 174 2125
rect 208 2091 243 2125
rect 277 2091 2298 2125
rect 2332 2091 2368 2125
rect 2402 2091 2438 2125
rect 2472 2091 2508 2125
rect 2542 2091 2578 2125
rect 2612 2091 2648 2125
rect 2682 2091 2718 2125
rect 2752 2091 2788 2125
rect 2822 2091 2858 2125
rect 2892 2091 2928 2125
rect 2962 2091 2998 2125
rect 3032 2091 3068 2125
rect 3102 2091 3138 2125
rect 3172 2091 3208 2125
rect 3242 2091 3278 2125
rect 3312 2091 3348 2125
rect 3382 2091 3418 2125
rect 3452 2091 3488 2125
rect 3522 2091 3558 2125
rect 3592 2091 3628 2125
rect 3662 2091 3698 2125
rect 3732 2091 3768 2125
rect 3802 2091 3838 2125
rect 3872 2091 3908 2125
rect 3942 2091 3977 2125
rect 4011 2091 4046 2125
rect 4080 2091 4115 2125
rect 4149 2091 4184 2125
rect 4218 2091 4253 2125
rect 4287 2091 4322 2125
rect 4356 2091 4391 2125
rect 4425 2091 4449 2125
rect -2750 2057 4449 2091
rect -2750 2023 -2726 2057
rect -2692 2023 -2656 2057
rect -2622 2023 -2586 2057
rect -2552 2023 -2517 2057
rect -2483 2023 -2448 2057
rect -2414 2023 -2379 2057
rect -2345 2023 -2310 2057
rect -2276 2023 -2241 2057
rect -2207 2023 -2172 2057
rect -2138 2023 -2103 2057
rect -2069 2023 -2034 2057
rect -2000 2023 -1965 2057
rect -1931 2023 -1896 2057
rect -1862 2023 -1827 2057
rect -1793 2023 -1758 2057
rect -1724 2023 -1689 2057
rect -1655 2023 -1620 2057
rect -1586 2023 -1551 2057
rect -1517 2023 -1482 2057
rect -1448 2023 -1413 2057
rect -1379 2023 -1344 2057
rect -1310 2023 -1275 2057
rect -1241 2023 -1206 2057
rect -1172 2023 -1137 2057
rect -1103 2023 -1068 2057
rect -1034 2023 -999 2057
rect -965 2023 -930 2057
rect -896 2023 -861 2057
rect -827 2023 -792 2057
rect -758 2023 -723 2057
rect -689 2023 -654 2057
rect -620 2023 -585 2057
rect -551 2023 -516 2057
rect -482 2023 -447 2057
rect -413 2023 -378 2057
rect -344 2023 -309 2057
rect -275 2023 -240 2057
rect -206 2023 -171 2057
rect -137 2023 -102 2057
rect -68 2023 -33 2057
rect 1 2023 36 2057
rect 70 2023 105 2057
rect 139 2023 174 2057
rect 208 2023 243 2057
rect 277 2023 2298 2057
rect 2332 2023 2368 2057
rect 2402 2023 2438 2057
rect 2472 2023 2508 2057
rect 2542 2023 2578 2057
rect 2612 2023 2648 2057
rect 2682 2023 2718 2057
rect 2752 2023 2788 2057
rect 2822 2023 2858 2057
rect 2892 2023 2928 2057
rect 2962 2023 2998 2057
rect 3032 2023 3068 2057
rect 3102 2023 3138 2057
rect 3172 2023 3208 2057
rect 3242 2023 3278 2057
rect 3312 2023 3348 2057
rect 3382 2023 3418 2057
rect 3452 2023 3488 2057
rect 3522 2023 3558 2057
rect 3592 2023 3628 2057
rect 3662 2023 3698 2057
rect 3732 2023 3768 2057
rect 3802 2023 3838 2057
rect 3872 2023 3908 2057
rect 3942 2023 3977 2057
rect 4011 2023 4046 2057
rect 4080 2023 4115 2057
rect 4149 2023 4184 2057
rect 4218 2023 4253 2057
rect 4287 2023 4322 2057
rect 4356 2023 4391 2057
rect 4425 2023 4449 2057
rect 10199 1236 10267 1270
rect 10301 1236 10335 1270
rect 10369 1236 10403 1270
rect 10437 1236 10471 1270
rect 10505 1236 10539 1270
rect 10573 1236 10607 1270
rect 10641 1236 10675 1270
rect 10709 1236 10743 1270
rect 10777 1236 10811 1270
rect 10845 1236 10879 1270
rect 10913 1236 10947 1270
rect 10981 1236 11015 1270
rect 11049 1236 11083 1270
rect 11117 1236 11151 1270
rect 11185 1236 11219 1270
rect 11253 1236 11287 1270
rect 11321 1236 11355 1270
rect 11389 1236 11423 1270
rect 11457 1236 11491 1270
rect 11525 1236 11559 1270
rect 11593 1236 11627 1270
rect 11661 1236 11695 1270
rect 11729 1236 11763 1270
rect 11797 1236 11831 1270
rect 11865 1236 11899 1270
rect 11933 1236 11967 1270
rect 12001 1236 12035 1270
rect 12069 1236 12103 1270
rect 12137 1236 12171 1270
rect 12205 1236 12239 1270
rect 12273 1236 12307 1270
rect 12341 1236 12375 1270
rect 12409 1236 12443 1270
rect 12477 1236 12511 1270
rect 12545 1236 12579 1270
rect 12613 1236 12647 1270
rect 12681 1236 12715 1270
rect 12749 1236 12783 1270
rect 12817 1236 12851 1270
rect 12885 1236 12919 1270
rect 12953 1236 12987 1270
rect 13021 1236 13055 1270
rect 13089 1236 13123 1270
rect 13157 1236 13191 1270
rect 13225 1236 13259 1270
rect 13293 1236 13327 1270
rect 13361 1236 13395 1270
rect 13429 1236 13463 1270
rect 13497 1236 13531 1270
rect 13565 1236 13599 1270
rect 13633 1236 13667 1270
rect 13701 1236 13735 1270
rect 13769 1236 13803 1270
rect 13837 1236 13871 1270
rect 13905 1236 13939 1270
rect 13973 1236 14007 1270
rect 14041 1236 14076 1270
rect 14110 1236 14145 1270
rect 14179 1236 14214 1270
rect 14248 1236 14283 1270
rect 14317 1236 14352 1270
rect 14386 1236 14421 1270
rect 14455 1236 14490 1270
rect 14524 1236 14559 1270
rect 14593 1236 14628 1270
rect 14662 1236 14697 1270
rect 14731 1236 14766 1270
rect 14800 1236 14835 1270
rect 14869 1236 14904 1270
rect 14938 1236 14973 1270
rect 15007 1236 15042 1270
rect 15076 1236 15111 1270
rect 15145 1236 15180 1270
rect 15214 1236 15249 1270
rect 15283 1236 15318 1270
rect 15352 1236 15420 1270
rect 10199 1201 15420 1236
rect 10199 1167 15386 1201
rect 10199 1161 15420 1167
rect 6202 1127 6270 1161
rect 6304 1127 6338 1161
rect 6372 1127 6406 1161
rect 6440 1127 6474 1161
rect 6508 1127 6542 1161
rect 6576 1127 6611 1161
rect 6645 1127 6680 1161
rect 6714 1127 6749 1161
rect 6783 1127 6818 1161
rect 6852 1127 6887 1161
rect 6921 1127 6956 1161
rect 6990 1127 7025 1161
rect 7059 1127 7094 1161
rect 7128 1127 7163 1161
rect 7197 1127 7232 1161
rect 7266 1127 7301 1161
rect 7335 1127 7370 1161
rect 7404 1127 7439 1161
rect 7473 1127 7508 1161
rect 7542 1127 7577 1161
rect 7611 1127 7646 1161
rect 7680 1127 7715 1161
rect 7749 1127 7784 1161
rect 7818 1127 7853 1161
rect 7887 1127 7922 1161
rect 7956 1127 7991 1161
rect 8025 1127 8060 1161
rect 8094 1127 8129 1161
rect 8163 1127 8198 1161
rect 8232 1127 8267 1161
rect 8301 1127 8336 1161
rect 8370 1127 8405 1161
rect 8439 1127 8474 1161
rect 8508 1127 8543 1161
rect 8577 1127 8612 1161
rect 8646 1127 8681 1161
rect 8715 1127 8750 1161
rect 8784 1127 8819 1161
rect 8853 1127 8888 1161
rect 8922 1127 8957 1161
rect 8991 1127 9026 1161
rect 9060 1127 9095 1161
rect 9129 1127 9164 1161
rect 9198 1127 9233 1161
rect 9267 1127 9302 1161
rect 9336 1127 9371 1161
rect 9405 1127 9440 1161
rect 9474 1127 9509 1161
rect 9543 1127 9578 1161
rect 9612 1127 9647 1161
rect 9681 1127 9716 1161
rect 9750 1127 9785 1161
rect 9819 1127 9854 1161
rect 9888 1127 9923 1161
rect 9957 1127 9992 1161
rect 10026 1127 10061 1161
rect 10095 1127 10130 1161
rect 10164 1127 10199 1161
rect 10233 1144 15420 1161
rect 10233 1127 10393 1144
rect 6202 1124 10393 1127
rect 6202 1093 10325 1124
rect 6236 1090 10325 1093
rect 10359 1110 10393 1124
rect 10427 1110 10461 1144
rect 10495 1110 10529 1144
rect 10563 1110 10597 1144
rect 10631 1110 10665 1144
rect 10699 1110 10733 1144
rect 10767 1110 10801 1144
rect 10835 1110 10869 1144
rect 10903 1110 10937 1144
rect 10971 1110 11005 1144
rect 11039 1110 11073 1144
rect 11107 1110 11141 1144
rect 11175 1110 11209 1144
rect 11243 1110 11277 1144
rect 11311 1110 11345 1144
rect 11379 1110 11413 1144
rect 11447 1110 11481 1144
rect 11515 1110 11549 1144
rect 11583 1110 11617 1144
rect 11651 1110 11685 1144
rect 11719 1110 11753 1144
rect 11787 1110 11821 1144
rect 11855 1110 11889 1144
rect 11923 1110 11957 1144
rect 11991 1110 12025 1144
rect 12059 1110 12093 1144
rect 12127 1110 12161 1144
rect 12195 1110 12229 1144
rect 12263 1110 12297 1144
rect 12331 1110 12365 1144
rect 12399 1110 12433 1144
rect 12467 1110 12501 1144
rect 12535 1110 12569 1144
rect 12603 1110 12638 1144
rect 12672 1110 12707 1144
rect 12741 1110 12776 1144
rect 12810 1110 12845 1144
rect 12879 1110 12914 1144
rect 12948 1110 12983 1144
rect 13017 1110 13052 1144
rect 13086 1110 13121 1144
rect 13155 1110 13190 1144
rect 13224 1110 13259 1144
rect 13293 1110 13328 1144
rect 13362 1110 13397 1144
rect 13431 1110 13466 1144
rect 13500 1110 13535 1144
rect 13569 1110 13604 1144
rect 13638 1110 13673 1144
rect 13707 1110 13742 1144
rect 13776 1110 13811 1144
rect 13845 1110 13880 1144
rect 13914 1110 13949 1144
rect 13983 1110 14018 1144
rect 14052 1110 14087 1144
rect 14121 1110 14156 1144
rect 14190 1110 14225 1144
rect 14259 1110 14294 1144
rect 14328 1110 14363 1144
rect 14397 1110 14432 1144
rect 14466 1110 14501 1144
rect 14535 1110 14570 1144
rect 14604 1110 14639 1144
rect 14673 1110 14708 1144
rect 14742 1110 14777 1144
rect 14811 1110 14846 1144
rect 14880 1110 14915 1144
rect 14949 1110 14984 1144
rect 15018 1110 15053 1144
rect 15087 1110 15122 1144
rect 15156 1110 15191 1144
rect 15225 1110 15260 1144
rect 15294 1132 15420 1144
rect 15294 1110 15386 1132
rect 6236 1059 10359 1090
rect 6202 1035 10359 1059
rect 6202 1018 6328 1035
rect 6236 1001 6328 1018
rect 6362 1001 6396 1035
rect 6430 1001 6464 1035
rect 6498 1001 6532 1035
rect 6566 1001 6600 1035
rect 6634 1001 6669 1035
rect 6703 1001 6738 1035
rect 6772 1001 6807 1035
rect 6841 1001 6876 1035
rect 6910 1001 6945 1035
rect 6979 1001 7014 1035
rect 7048 1001 7083 1035
rect 7117 1001 7152 1035
rect 7186 1001 7221 1035
rect 7255 1001 7290 1035
rect 7324 1001 7359 1035
rect 7393 1001 7428 1035
rect 7462 1001 7497 1035
rect 7531 1001 7566 1035
rect 7600 1001 7635 1035
rect 7669 1001 7704 1035
rect 7738 1001 7773 1035
rect 7807 1001 7842 1035
rect 7876 1001 7911 1035
rect 7945 1001 7980 1035
rect 8014 1001 8049 1035
rect 8083 1001 8118 1035
rect 8152 1001 8187 1035
rect 8221 1001 8256 1035
rect 8290 1001 8325 1035
rect 8359 1001 8394 1035
rect 8428 1001 8463 1035
rect 8497 1001 8532 1035
rect 8566 1001 8601 1035
rect 8635 1001 8670 1035
rect 8704 1001 8739 1035
rect 8773 1001 8808 1035
rect 8842 1001 8877 1035
rect 8911 1001 8946 1035
rect 8980 1001 9015 1035
rect 9049 1001 9084 1035
rect 9118 1001 9153 1035
rect 9187 1001 9222 1035
rect 9256 1001 9291 1035
rect 9325 1001 9360 1035
rect 9394 1001 9429 1035
rect 9463 1001 9498 1035
rect 9532 1001 9567 1035
rect 9601 1001 9636 1035
rect 9670 1001 9705 1035
rect 9739 1001 9774 1035
rect 9808 1001 9843 1035
rect 9877 1001 9912 1035
rect 9946 1001 9981 1035
rect 10015 1001 10050 1035
rect 10084 1001 10119 1035
rect 10153 1001 10188 1035
rect 10222 1001 10257 1035
rect 10291 1001 10359 1035
rect 15260 1098 15386 1110
rect 15260 1074 15420 1098
rect 15294 1063 15420 1074
rect 15294 1040 15386 1063
rect 15260 1029 15386 1040
rect 15260 1003 15420 1029
rect 6236 984 6362 1001
rect 6202 957 6362 984
rect 15294 994 15420 1003
rect 15294 969 15386 994
rect 15260 960 15386 969
rect 6202 943 6328 957
rect 6236 923 6328 943
rect 6236 909 6362 923
rect 6202 880 6362 909
rect 6202 868 6328 880
rect 6236 846 6328 868
rect 6236 834 6362 846
rect 15260 932 15420 960
rect 6202 803 6362 834
rect 6202 793 6328 803
rect 6236 769 6328 793
rect 15294 925 15420 932
rect 15294 898 15386 925
rect 15260 891 15386 898
rect 15260 861 15420 891
rect 15294 856 15420 861
rect 15294 827 15386 856
rect 15260 822 15386 827
rect 6236 759 6362 769
rect 6202 726 6362 759
rect 6202 718 6328 726
rect 6236 692 6328 718
rect 15260 790 15420 822
rect 15294 786 15420 790
rect 15294 756 15386 786
rect 15260 752 15386 756
rect 6236 684 6362 692
rect 6202 649 6362 684
rect 15260 719 15420 752
rect 15294 716 15420 719
rect 15294 685 15386 716
rect 15260 682 15386 685
rect 6202 643 6328 649
rect 6236 615 6328 643
rect 6236 609 6362 615
rect 6202 572 6362 609
rect 6202 569 6328 572
rect 6236 538 6328 569
rect 6236 535 6362 538
rect 6202 495 6362 535
rect 6236 461 6328 495
rect 6202 391 6362 461
rect 15260 648 15420 682
rect 15294 646 15420 648
rect 15294 614 15386 646
rect 15260 612 15386 614
rect 15260 577 15420 612
rect 15294 576 15420 577
rect 15294 543 15386 576
rect 15260 542 15386 543
rect 15260 506 15420 542
rect 15294 472 15386 506
rect 15260 391 15420 472
<< psubdiffcont >>
rect -2859 1812 -2825 1846
rect -2790 1812 -2756 1846
rect -2721 1812 -2687 1846
rect -2652 1812 -2618 1846
rect -2583 1812 -2549 1846
rect -2514 1812 -2480 1846
rect -2445 1812 -2411 1846
rect -2376 1812 -2342 1846
rect -2307 1812 -2273 1846
rect -2238 1812 -2204 1846
rect -2169 1812 -2135 1846
rect -2100 1812 -2066 1846
rect -2031 1812 -1997 1846
rect -1962 1812 -1928 1846
rect -1893 1812 -1859 1846
rect -1824 1812 -1790 1846
rect -1755 1812 -1721 1846
rect -1686 1812 -1652 1846
rect -1617 1812 -1583 1846
rect -1548 1812 -1514 1846
rect -1479 1812 -1445 1846
rect -1410 1812 -1376 1846
rect -1341 1812 -1307 1846
rect -1272 1812 -1238 1846
rect -1203 1812 -1169 1846
rect -1134 1812 -1100 1846
rect -1065 1812 -1031 1846
rect -996 1812 -962 1846
rect -927 1812 -893 1846
rect -858 1812 -824 1846
rect -789 1812 -755 1846
rect -720 1812 -686 1846
rect -651 1812 -617 1846
rect -582 1812 -548 1846
rect -513 1812 -479 1846
rect -444 1812 -410 1846
rect -2859 1744 -2825 1778
rect -2790 1744 -2756 1778
rect -2721 1744 -2687 1778
rect -2652 1744 -2618 1778
rect -2583 1744 -2549 1778
rect -2514 1744 -2480 1778
rect -2445 1744 -2411 1778
rect -2376 1744 -2342 1778
rect -2307 1744 -2273 1778
rect -2238 1744 -2204 1778
rect -2169 1744 -2135 1778
rect -2100 1744 -2066 1778
rect -2031 1744 -1997 1778
rect -1962 1744 -1928 1778
rect -1893 1744 -1859 1778
rect -1824 1744 -1790 1778
rect -1755 1744 -1721 1778
rect -1686 1744 -1652 1778
rect -1617 1744 -1583 1778
rect -1548 1744 -1514 1778
rect -1479 1744 -1445 1778
rect -1410 1744 -1376 1778
rect -1341 1744 -1307 1778
rect -1272 1744 -1238 1778
rect -1203 1744 -1169 1778
rect -1134 1744 -1100 1778
rect -1065 1744 -1031 1778
rect -996 1744 -962 1778
rect -927 1744 -893 1778
rect -858 1744 -824 1778
rect -789 1744 -755 1778
rect -720 1744 -686 1778
rect -651 1744 -617 1778
rect -582 1744 -548 1778
rect -513 1744 -479 1778
rect -444 1744 -410 1778
rect -2859 1676 -2825 1710
rect -2790 1676 -2756 1710
rect -2721 1676 -2687 1710
rect -2652 1676 -2618 1710
rect -2583 1676 -2549 1710
rect -2514 1676 -2480 1710
rect -2445 1676 -2411 1710
rect -2376 1676 -2342 1710
rect -2307 1676 -2273 1710
rect -2238 1676 -2204 1710
rect -2169 1676 -2135 1710
rect -2100 1676 -2066 1710
rect -2031 1676 -1997 1710
rect -1962 1676 -1928 1710
rect -1893 1676 -1859 1710
rect -1824 1676 -1790 1710
rect -1755 1676 -1721 1710
rect -1686 1676 -1652 1710
rect -1617 1676 -1583 1710
rect -1548 1676 -1514 1710
rect -1479 1676 -1445 1710
rect -1410 1676 -1376 1710
rect -1341 1676 -1307 1710
rect -1272 1676 -1238 1710
rect -1203 1676 -1169 1710
rect -1134 1676 -1100 1710
rect -1065 1676 -1031 1710
rect -996 1676 -962 1710
rect -927 1676 -893 1710
rect -858 1676 -824 1710
rect -789 1676 -755 1710
rect -720 1676 -686 1710
rect -651 1676 -617 1710
rect -582 1676 -548 1710
rect -513 1676 -479 1710
rect -444 1676 -410 1710
rect -2859 1608 -2825 1642
rect -2790 1608 -2756 1642
rect -2721 1608 -2687 1642
rect -2652 1608 -2618 1642
rect -2583 1608 -2549 1642
rect -2514 1608 -2480 1642
rect -2445 1608 -2411 1642
rect -2376 1608 -2342 1642
rect -2307 1608 -2273 1642
rect -2238 1608 -2204 1642
rect -2169 1608 -2135 1642
rect -2100 1608 -2066 1642
rect -2031 1608 -1997 1642
rect -1962 1608 -1928 1642
rect -1893 1608 -1859 1642
rect -1824 1608 -1790 1642
rect -1755 1608 -1721 1642
rect -1686 1608 -1652 1642
rect -1617 1608 -1583 1642
rect -1548 1608 -1514 1642
rect -1479 1608 -1445 1642
rect -1410 1608 -1376 1642
rect -1341 1608 -1307 1642
rect -1272 1608 -1238 1642
rect -1203 1608 -1169 1642
rect -1134 1608 -1100 1642
rect -1065 1608 -1031 1642
rect -996 1608 -962 1642
rect -927 1608 -893 1642
rect -858 1608 -824 1642
rect -789 1608 -755 1642
rect -720 1608 -686 1642
rect -651 1608 -617 1642
rect -582 1608 -548 1642
rect -513 1608 -479 1642
rect -444 1608 -410 1642
rect -2859 1540 -2825 1574
rect -2790 1540 -2756 1574
rect -2721 1540 -2687 1574
rect -2652 1540 -2618 1574
rect -2583 1540 -2549 1574
rect -2514 1540 -2480 1574
rect -2445 1540 -2411 1574
rect -2376 1540 -2342 1574
rect -2307 1540 -2273 1574
rect -2238 1540 -2204 1574
rect -2169 1540 -2135 1574
rect -2100 1540 -2066 1574
rect -2031 1540 -1997 1574
rect -1962 1540 -1928 1574
rect -1893 1540 -1859 1574
rect -1824 1540 -1790 1574
rect -1755 1540 -1721 1574
rect -1686 1540 -1652 1574
rect -1617 1540 -1583 1574
rect -1548 1540 -1514 1574
rect -1479 1540 -1445 1574
rect -1410 1540 -1376 1574
rect -1341 1540 -1307 1574
rect -1272 1540 -1238 1574
rect -1203 1540 -1169 1574
rect -1134 1540 -1100 1574
rect -1065 1540 -1031 1574
rect -996 1540 -962 1574
rect -927 1540 -893 1574
rect -858 1540 -824 1574
rect -789 1540 -755 1574
rect -720 1540 -686 1574
rect -651 1540 -617 1574
rect -582 1540 -548 1574
rect -513 1540 -479 1574
rect -444 1540 -410 1574
rect -2859 1472 -2825 1506
rect -2790 1472 -2756 1506
rect -2721 1472 -2687 1506
rect -2652 1472 -2618 1506
rect -2583 1472 -2549 1506
rect -2514 1472 -2480 1506
rect -2445 1472 -2411 1506
rect -2376 1472 -2342 1506
rect -2307 1472 -2273 1506
rect -2238 1472 -2204 1506
rect -2169 1472 -2135 1506
rect -2100 1472 -2066 1506
rect -2031 1472 -1997 1506
rect -1962 1472 -1928 1506
rect -1893 1472 -1859 1506
rect -1824 1472 -1790 1506
rect -1755 1472 -1721 1506
rect -1686 1472 -1652 1506
rect -1617 1472 -1583 1506
rect -1548 1472 -1514 1506
rect -1479 1472 -1445 1506
rect -1410 1472 -1376 1506
rect -1341 1472 -1307 1506
rect -1272 1472 -1238 1506
rect -1203 1472 -1169 1506
rect -1134 1472 -1100 1506
rect -1065 1472 -1031 1506
rect -996 1472 -962 1506
rect -927 1472 -893 1506
rect -858 1472 -824 1506
rect -789 1472 -755 1506
rect -720 1472 -686 1506
rect -651 1472 -617 1506
rect -582 1472 -548 1506
rect -513 1472 -479 1506
rect -444 1472 -410 1506
rect -2859 1404 -2825 1438
rect -2790 1404 -2756 1438
rect -2721 1404 -2687 1438
rect -2652 1404 -2618 1438
rect -2583 1404 -2549 1438
rect -2514 1404 -2480 1438
rect -2445 1404 -2411 1438
rect -2376 1404 -2342 1438
rect -2307 1404 -2273 1438
rect -2238 1404 -2204 1438
rect -2169 1404 -2135 1438
rect -2100 1404 -2066 1438
rect -2031 1404 -1997 1438
rect -1962 1404 -1928 1438
rect -1893 1404 -1859 1438
rect -1824 1404 -1790 1438
rect -1755 1404 -1721 1438
rect -1686 1404 -1652 1438
rect -1617 1404 -1583 1438
rect -1548 1404 -1514 1438
rect -1479 1404 -1445 1438
rect -1410 1404 -1376 1438
rect -1341 1404 -1307 1438
rect -1272 1404 -1238 1438
rect -1203 1404 -1169 1438
rect -1134 1404 -1100 1438
rect -1065 1404 -1031 1438
rect -996 1404 -962 1438
rect -927 1404 -893 1438
rect -858 1404 -824 1438
rect -789 1404 -755 1438
rect -720 1404 -686 1438
rect -651 1404 -617 1438
rect -582 1404 -548 1438
rect -513 1404 -479 1438
rect -444 1404 -410 1438
rect -2859 1336 -2825 1370
rect -2790 1336 -2756 1370
rect -2721 1336 -2687 1370
rect -2652 1336 -2618 1370
rect -2583 1336 -2549 1370
rect -2514 1336 -2480 1370
rect -2445 1336 -2411 1370
rect -2376 1336 -2342 1370
rect -2307 1336 -2273 1370
rect -2238 1336 -2204 1370
rect -2169 1336 -2135 1370
rect -2100 1336 -2066 1370
rect -2031 1336 -1997 1370
rect -1962 1336 -1928 1370
rect -1893 1336 -1859 1370
rect -1824 1336 -1790 1370
rect -1755 1336 -1721 1370
rect -1686 1336 -1652 1370
rect -1617 1336 -1583 1370
rect -1548 1336 -1514 1370
rect -1479 1336 -1445 1370
rect -1410 1336 -1376 1370
rect -1341 1336 -1307 1370
rect -1272 1336 -1238 1370
rect -1203 1336 -1169 1370
rect -1134 1336 -1100 1370
rect -1065 1336 -1031 1370
rect -996 1336 -962 1370
rect -927 1336 -893 1370
rect -858 1336 -824 1370
rect -789 1336 -755 1370
rect -720 1336 -686 1370
rect -651 1336 -617 1370
rect -582 1336 -548 1370
rect -513 1336 -479 1370
rect -444 1336 -410 1370
rect -2859 1268 -2825 1302
rect -2790 1268 -2756 1302
rect -2721 1268 -2687 1302
rect -2652 1268 -2618 1302
rect -2583 1268 -2549 1302
rect -2514 1268 -2480 1302
rect -2445 1268 -2411 1302
rect -2376 1268 -2342 1302
rect -2307 1268 -2273 1302
rect -2238 1268 -2204 1302
rect -2169 1268 -2135 1302
rect -2100 1268 -2066 1302
rect -2031 1268 -1997 1302
rect -1962 1268 -1928 1302
rect -1893 1268 -1859 1302
rect -1824 1268 -1790 1302
rect -1755 1268 -1721 1302
rect -1686 1268 -1652 1302
rect -1617 1268 -1583 1302
rect -1548 1268 -1514 1302
rect -1479 1268 -1445 1302
rect -1410 1268 -1376 1302
rect -1341 1268 -1307 1302
rect -1272 1268 -1238 1302
rect -1203 1268 -1169 1302
rect -1134 1268 -1100 1302
rect -1065 1268 -1031 1302
rect -996 1268 -962 1302
rect -927 1268 -893 1302
rect -858 1268 -824 1302
rect -789 1268 -755 1302
rect -720 1268 -686 1302
rect -651 1268 -617 1302
rect -582 1268 -548 1302
rect -513 1268 -479 1302
rect -444 1268 -410 1302
rect -2859 1200 -2825 1234
rect -2790 1200 -2756 1234
rect -2721 1200 -2687 1234
rect -2652 1200 -2618 1234
rect -2583 1200 -2549 1234
rect -2514 1200 -2480 1234
rect -2445 1200 -2411 1234
rect -2376 1200 -2342 1234
rect -2307 1200 -2273 1234
rect -2238 1200 -2204 1234
rect -2169 1200 -2135 1234
rect -2100 1200 -2066 1234
rect -2031 1200 -1997 1234
rect -1962 1200 -1928 1234
rect -1893 1200 -1859 1234
rect -1824 1200 -1790 1234
rect -1755 1200 -1721 1234
rect -1686 1200 -1652 1234
rect -1617 1200 -1583 1234
rect -1548 1200 -1514 1234
rect -1479 1200 -1445 1234
rect -1410 1200 -1376 1234
rect -1341 1200 -1307 1234
rect -1272 1200 -1238 1234
rect -1203 1200 -1169 1234
rect -1134 1200 -1100 1234
rect -1065 1200 -1031 1234
rect -996 1200 -962 1234
rect -927 1200 -893 1234
rect -858 1200 -824 1234
rect -789 1200 -755 1234
rect -720 1200 -686 1234
rect -651 1200 -617 1234
rect -582 1200 -548 1234
rect -513 1200 -479 1234
rect -444 1200 -410 1234
rect -2859 1132 -2825 1166
rect -2790 1132 -2756 1166
rect -2721 1132 -2687 1166
rect -2652 1132 -2618 1166
rect -2583 1132 -2549 1166
rect -2514 1132 -2480 1166
rect -2445 1132 -2411 1166
rect -2376 1132 -2342 1166
rect -2307 1132 -2273 1166
rect -2238 1132 -2204 1166
rect -2169 1132 -2135 1166
rect -2100 1132 -2066 1166
rect -2031 1132 -1997 1166
rect -1962 1132 -1928 1166
rect -1893 1132 -1859 1166
rect -1824 1132 -1790 1166
rect -1755 1132 -1721 1166
rect -1686 1132 -1652 1166
rect -1617 1132 -1583 1166
rect -1548 1132 -1514 1166
rect -1479 1132 -1445 1166
rect -1410 1132 -1376 1166
rect -1341 1132 -1307 1166
rect -1272 1132 -1238 1166
rect -1203 1132 -1169 1166
rect -1134 1132 -1100 1166
rect -1065 1132 -1031 1166
rect -996 1132 -962 1166
rect -927 1132 -893 1166
rect -858 1132 -824 1166
rect -789 1132 -755 1166
rect -720 1132 -686 1166
rect -651 1132 -617 1166
rect -582 1132 -548 1166
rect -513 1132 -479 1166
rect -444 1132 -410 1166
rect -2859 1064 -2825 1098
rect -2790 1064 -2756 1098
rect -2721 1064 -2687 1098
rect -2652 1064 -2618 1098
rect -2583 1064 -2549 1098
rect -2514 1064 -2480 1098
rect -2445 1064 -2411 1098
rect -2376 1064 -2342 1098
rect -2307 1064 -2273 1098
rect -2238 1064 -2204 1098
rect -2169 1064 -2135 1098
rect -2100 1064 -2066 1098
rect -2031 1064 -1997 1098
rect -1962 1064 -1928 1098
rect -1893 1064 -1859 1098
rect -1824 1064 -1790 1098
rect -1755 1064 -1721 1098
rect -1686 1064 -1652 1098
rect -1617 1064 -1583 1098
rect -1548 1064 -1514 1098
rect -1479 1064 -1445 1098
rect -1410 1064 -1376 1098
rect -1341 1064 -1307 1098
rect -1272 1064 -1238 1098
rect -1203 1064 -1169 1098
rect -1134 1064 -1100 1098
rect -1065 1064 -1031 1098
rect -996 1064 -962 1098
rect -927 1064 -893 1098
rect -858 1064 -824 1098
rect -789 1064 -755 1098
rect -720 1064 -686 1098
rect -651 1064 -617 1098
rect -582 1064 -548 1098
rect -513 1064 -479 1098
rect -444 1064 -410 1098
rect -2859 996 -2825 1030
rect -2790 996 -2756 1030
rect -2721 996 -2687 1030
rect -2652 996 -2618 1030
rect -2583 996 -2549 1030
rect -2514 996 -2480 1030
rect -2445 996 -2411 1030
rect -2376 996 -2342 1030
rect -2307 996 -2273 1030
rect -2238 996 -2204 1030
rect -2169 996 -2135 1030
rect -2100 996 -2066 1030
rect -2031 996 -1997 1030
rect -1962 996 -1928 1030
rect -1893 996 -1859 1030
rect -1824 996 -1790 1030
rect -1755 996 -1721 1030
rect -1686 996 -1652 1030
rect -1617 996 -1583 1030
rect -1548 996 -1514 1030
rect -1479 996 -1445 1030
rect -1410 996 -1376 1030
rect -1341 996 -1307 1030
rect -1272 996 -1238 1030
rect -1203 996 -1169 1030
rect -1134 996 -1100 1030
rect -1065 996 -1031 1030
rect -996 996 -962 1030
rect -927 996 -893 1030
rect -858 996 -824 1030
rect -789 996 -755 1030
rect -720 996 -686 1030
rect -651 996 -617 1030
rect -582 996 -548 1030
rect -513 996 -479 1030
rect -444 996 -410 1030
rect -2859 928 -2825 962
rect -2790 928 -2756 962
rect -2721 928 -2687 962
rect -2652 928 -2618 962
rect -2583 928 -2549 962
rect -2514 928 -2480 962
rect -2445 928 -2411 962
rect -2376 928 -2342 962
rect -2307 928 -2273 962
rect -2238 928 -2204 962
rect -2169 928 -2135 962
rect -2100 928 -2066 962
rect -2031 928 -1997 962
rect -1962 928 -1928 962
rect -1893 928 -1859 962
rect -1824 928 -1790 962
rect -1755 928 -1721 962
rect -1686 928 -1652 962
rect -1617 928 -1583 962
rect -1548 928 -1514 962
rect -1479 928 -1445 962
rect -1410 928 -1376 962
rect -1341 928 -1307 962
rect -1272 928 -1238 962
rect -1203 928 -1169 962
rect -1134 928 -1100 962
rect -1065 928 -1031 962
rect -996 928 -962 962
rect -927 928 -893 962
rect -858 928 -824 962
rect -789 928 -755 962
rect -720 928 -686 962
rect -651 928 -617 962
rect -582 928 -548 962
rect -513 928 -479 962
rect -444 928 -410 962
rect -2859 860 -2825 894
rect -2790 860 -2756 894
rect -2721 860 -2687 894
rect -2652 860 -2618 894
rect -2583 860 -2549 894
rect -2514 860 -2480 894
rect -2445 860 -2411 894
rect -2376 860 -2342 894
rect -2307 860 -2273 894
rect -2238 860 -2204 894
rect -2169 860 -2135 894
rect -2100 860 -2066 894
rect -2031 860 -1997 894
rect -1962 860 -1928 894
rect -1893 860 -1859 894
rect -1824 860 -1790 894
rect -1755 860 -1721 894
rect -1686 860 -1652 894
rect -1617 860 -1583 894
rect -1548 860 -1514 894
rect -1479 860 -1445 894
rect -1410 860 -1376 894
rect -1341 860 -1307 894
rect -1272 860 -1238 894
rect -1203 860 -1169 894
rect -1134 860 -1100 894
rect -1065 860 -1031 894
rect -996 860 -962 894
rect -927 860 -893 894
rect -858 860 -824 894
rect -789 860 -755 894
rect -720 860 -686 894
rect -651 860 -617 894
rect -582 860 -548 894
rect -513 860 -479 894
rect -444 860 -410 894
rect -2859 792 -2825 826
rect -2790 792 -2756 826
rect -2721 792 -2687 826
rect -2652 792 -2618 826
rect -2583 792 -2549 826
rect -2514 792 -2480 826
rect -2445 792 -2411 826
rect -2376 792 -2342 826
rect -2307 792 -2273 826
rect -2238 792 -2204 826
rect -2169 792 -2135 826
rect -2100 792 -2066 826
rect -2031 792 -1997 826
rect -1962 792 -1928 826
rect -1893 792 -1859 826
rect -1824 792 -1790 826
rect -1755 792 -1721 826
rect -1686 792 -1652 826
rect -1617 792 -1583 826
rect -1548 792 -1514 826
rect -1479 792 -1445 826
rect -1410 792 -1376 826
rect -1341 792 -1307 826
rect -1272 792 -1238 826
rect -1203 792 -1169 826
rect -1134 792 -1100 826
rect -1065 792 -1031 826
rect -996 792 -962 826
rect -927 792 -893 826
rect -858 792 -824 826
rect -789 792 -755 826
rect -720 792 -686 826
rect -651 792 -617 826
rect -582 792 -548 826
rect -513 792 -479 826
rect -444 792 -410 826
rect -375 792 -1 1846
<< mvpsubdiffcont >>
rect 11949 4290 11983 4324
rect 12018 4290 12052 4324
rect 12087 4290 12121 4324
rect 12156 4290 12190 4324
rect 12225 4290 12259 4324
rect 12294 4290 12328 4324
rect 12363 4290 12397 4324
rect 12432 4290 12466 4324
rect 12501 4290 12535 4324
rect 12570 4290 12604 4324
rect 12639 4290 12673 4324
rect 12708 4290 12742 4324
rect 12777 4290 12811 4324
rect 12846 4290 12880 4324
rect 12915 4290 12949 4324
rect 12984 4290 13018 4324
rect 13053 4290 13087 4324
rect 13122 4290 13156 4324
rect 13191 4290 13225 4324
rect 13260 4290 13294 4324
rect 13329 4290 13363 4324
rect 13398 4290 13432 4324
rect 13467 4290 13501 4324
rect 13536 4290 13570 4324
rect 13605 4290 13639 4324
rect 13674 4290 13708 4324
rect 13743 4290 13777 4324
rect 13812 4290 13846 4324
rect 13881 4290 13915 4324
rect 13950 4290 13984 4324
rect 14019 4290 14053 4324
rect 14088 4290 14122 4324
rect 14157 4290 14191 4324
rect 14226 4290 14260 4324
rect 14295 4290 14329 4324
rect 14364 4290 14398 4324
rect 14433 4290 14467 4324
rect 14502 4290 14536 4324
rect 14571 4290 14605 4324
rect 14640 4290 14674 4324
rect 14709 4290 14743 4324
rect 14778 4290 14812 4324
rect 14847 4290 14881 4324
rect 14916 4290 14950 4324
rect 14985 4290 15019 4324
rect 15054 4290 15088 4324
rect 15123 4290 15157 4324
rect 15192 4290 15226 4324
rect 15261 4290 15295 4324
rect 15330 4290 15364 4324
rect 15399 4290 15433 4324
rect 15468 4290 15502 4324
rect 15537 4290 15571 4324
rect 15606 4290 15640 4324
rect 15675 4290 15709 4324
rect 15744 4290 15778 4324
rect 15813 4290 15847 4324
rect 15882 4290 15916 4324
rect 15951 4290 15985 4324
rect 16020 4290 16054 4324
rect 16089 4290 16123 4324
rect 16158 4290 16192 4324
rect 16227 4290 16261 4324
rect 16296 4290 16330 4324
rect 11949 4222 11983 4256
rect 12018 4222 12052 4256
rect 12087 4222 12121 4256
rect 12156 4222 12190 4256
rect 12225 4222 12259 4256
rect 12294 4222 12328 4256
rect 12363 4222 12397 4256
rect 12432 4222 12466 4256
rect 12501 4222 12535 4256
rect 12570 4222 12604 4256
rect 12639 4222 12673 4256
rect 12708 4222 12742 4256
rect 12777 4222 12811 4256
rect 12846 4222 12880 4256
rect 12915 4222 12949 4256
rect 12984 4222 13018 4256
rect 13053 4222 13087 4256
rect 13122 4222 13156 4256
rect 13191 4222 13225 4256
rect 13260 4222 13294 4256
rect 13329 4222 13363 4256
rect 13398 4222 13432 4256
rect 13467 4222 13501 4256
rect 13536 4222 13570 4256
rect 13605 4222 13639 4256
rect 13674 4222 13708 4256
rect 13743 4222 13777 4256
rect 13812 4222 13846 4256
rect 13881 4222 13915 4256
rect 13950 4222 13984 4256
rect 14019 4222 14053 4256
rect 14088 4222 14122 4256
rect 14157 4222 14191 4256
rect 14226 4222 14260 4256
rect 14295 4222 14329 4256
rect 14364 4222 14398 4256
rect 14433 4222 14467 4256
rect 14502 4222 14536 4256
rect 14571 4222 14605 4256
rect 14640 4222 14674 4256
rect 14709 4222 14743 4256
rect 14778 4222 14812 4256
rect 14847 4222 14881 4256
rect 14916 4222 14950 4256
rect 14985 4222 15019 4256
rect 15054 4222 15088 4256
rect 15123 4222 15157 4256
rect 15192 4222 15226 4256
rect 15261 4222 15295 4256
rect 15330 4222 15364 4256
rect 15399 4222 15433 4256
rect 15468 4222 15502 4256
rect 15537 4222 15571 4256
rect 15606 4222 15640 4256
rect 15675 4222 15709 4256
rect 15744 4222 15778 4256
rect 15813 4222 15847 4256
rect 15882 4222 15916 4256
rect 15951 4222 15985 4256
rect 16020 4222 16054 4256
rect 16089 4222 16123 4256
rect 16158 4222 16192 4256
rect 16227 4222 16261 4256
rect 16296 4222 16330 4256
rect 11949 4154 11983 4188
rect 12018 4154 12052 4188
rect 12087 4154 12121 4188
rect 12156 4154 12190 4188
rect 12225 4154 12259 4188
rect 12294 4154 12328 4188
rect 12363 4154 12397 4188
rect 12432 4154 12466 4188
rect 12501 4154 12535 4188
rect 12570 4154 12604 4188
rect 12639 4154 12673 4188
rect 12708 4154 12742 4188
rect 12777 4154 12811 4188
rect 12846 4154 12880 4188
rect 12915 4154 12949 4188
rect 12984 4154 13018 4188
rect 13053 4154 13087 4188
rect 13122 4154 13156 4188
rect 13191 4154 13225 4188
rect 13260 4154 13294 4188
rect 13329 4154 13363 4188
rect 13398 4154 13432 4188
rect 13467 4154 13501 4188
rect 13536 4154 13570 4188
rect 13605 4154 13639 4188
rect 13674 4154 13708 4188
rect 13743 4154 13777 4188
rect 13812 4154 13846 4188
rect 13881 4154 13915 4188
rect 13950 4154 13984 4188
rect 14019 4154 14053 4188
rect 14088 4154 14122 4188
rect 14157 4154 14191 4188
rect 14226 4154 14260 4188
rect 14295 4154 14329 4188
rect 14364 4154 14398 4188
rect 14433 4154 14467 4188
rect 14502 4154 14536 4188
rect 14571 4154 14605 4188
rect 14640 4154 14674 4188
rect 14709 4154 14743 4188
rect 14778 4154 14812 4188
rect 14847 4154 14881 4188
rect 14916 4154 14950 4188
rect 14985 4154 15019 4188
rect 15054 4154 15088 4188
rect 15123 4154 15157 4188
rect 15192 4154 15226 4188
rect 15261 4154 15295 4188
rect 15330 4154 15364 4188
rect 15399 4154 15433 4188
rect 15468 4154 15502 4188
rect 15537 4154 15571 4188
rect 15606 4154 15640 4188
rect 15675 4154 15709 4188
rect 15744 4154 15778 4188
rect 15813 4154 15847 4188
rect 15882 4154 15916 4188
rect 15951 4154 15985 4188
rect 16020 4154 16054 4188
rect 16089 4154 16123 4188
rect 16158 4154 16192 4188
rect 16227 4154 16261 4188
rect 16296 4154 16330 4188
rect 11949 4086 11983 4120
rect 12018 4086 12052 4120
rect 12087 4086 12121 4120
rect 12156 4086 12190 4120
rect 12225 4086 12259 4120
rect 12294 4086 12328 4120
rect 12363 4086 12397 4120
rect 12432 4086 12466 4120
rect 12501 4086 12535 4120
rect 12570 4086 12604 4120
rect 12639 4086 12673 4120
rect 12708 4086 12742 4120
rect 12777 4086 12811 4120
rect 12846 4086 12880 4120
rect 12915 4086 12949 4120
rect 12984 4086 13018 4120
rect 13053 4086 13087 4120
rect 13122 4086 13156 4120
rect 13191 4086 13225 4120
rect 13260 4086 13294 4120
rect 13329 4086 13363 4120
rect 13398 4086 13432 4120
rect 13467 4086 13501 4120
rect 13536 4086 13570 4120
rect 13605 4086 13639 4120
rect 13674 4086 13708 4120
rect 13743 4086 13777 4120
rect 13812 4086 13846 4120
rect 13881 4086 13915 4120
rect 13950 4086 13984 4120
rect 14019 4086 14053 4120
rect 14088 4086 14122 4120
rect 14157 4086 14191 4120
rect 14226 4086 14260 4120
rect 14295 4086 14329 4120
rect 14364 4086 14398 4120
rect 14433 4086 14467 4120
rect 14502 4086 14536 4120
rect 14571 4086 14605 4120
rect 14640 4086 14674 4120
rect 14709 4086 14743 4120
rect 14778 4086 14812 4120
rect 14847 4086 14881 4120
rect 14916 4086 14950 4120
rect 14985 4086 15019 4120
rect 15054 4086 15088 4120
rect 15123 4086 15157 4120
rect 15192 4086 15226 4120
rect 15261 4086 15295 4120
rect 15330 4086 15364 4120
rect 15399 4086 15433 4120
rect 15468 4086 15502 4120
rect 15537 4086 15571 4120
rect 15606 4086 15640 4120
rect 15675 4086 15709 4120
rect 15744 4086 15778 4120
rect 15813 4086 15847 4120
rect 15882 4086 15916 4120
rect 15951 4086 15985 4120
rect 16020 4086 16054 4120
rect 16089 4086 16123 4120
rect 16158 4086 16192 4120
rect 16227 4086 16261 4120
rect 16296 4086 16330 4120
rect 11949 4018 11983 4052
rect 12018 4018 12052 4052
rect 12087 4018 12121 4052
rect 12156 4018 12190 4052
rect 12225 4018 12259 4052
rect 12294 4018 12328 4052
rect 12363 4018 12397 4052
rect 12432 4018 12466 4052
rect 12501 4018 12535 4052
rect 12570 4018 12604 4052
rect 12639 4018 12673 4052
rect 12708 4018 12742 4052
rect 12777 4018 12811 4052
rect 12846 4018 12880 4052
rect 12915 4018 12949 4052
rect 12984 4018 13018 4052
rect 13053 4018 13087 4052
rect 13122 4018 13156 4052
rect 13191 4018 13225 4052
rect 13260 4018 13294 4052
rect 13329 4018 13363 4052
rect 13398 4018 13432 4052
rect 13467 4018 13501 4052
rect 13536 4018 13570 4052
rect 13605 4018 13639 4052
rect 13674 4018 13708 4052
rect 13743 4018 13777 4052
rect 13812 4018 13846 4052
rect 13881 4018 13915 4052
rect 13950 4018 13984 4052
rect 14019 4018 14053 4052
rect 14088 4018 14122 4052
rect 14157 4018 14191 4052
rect 14226 4018 14260 4052
rect 14295 4018 14329 4052
rect 14364 4018 14398 4052
rect 14433 4018 14467 4052
rect 14502 4018 14536 4052
rect 14571 4018 14605 4052
rect 14640 4018 14674 4052
rect 14709 4018 14743 4052
rect 14778 4018 14812 4052
rect 14847 4018 14881 4052
rect 14916 4018 14950 4052
rect 14985 4018 15019 4052
rect 15054 4018 15088 4052
rect 15123 4018 15157 4052
rect 15192 4018 15226 4052
rect 15261 4018 15295 4052
rect 15330 4018 15364 4052
rect 15399 4018 15433 4052
rect 15468 4018 15502 4052
rect 15537 4018 15571 4052
rect 15606 4018 15640 4052
rect 15675 4018 15709 4052
rect 15744 4018 15778 4052
rect 15813 4018 15847 4052
rect 15882 4018 15916 4052
rect 15951 4018 15985 4052
rect 16020 4018 16054 4052
rect 16089 4018 16123 4052
rect 16158 4018 16192 4052
rect 16227 4018 16261 4052
rect 16296 4018 16330 4052
rect 11949 3950 11983 3984
rect 12018 3950 12052 3984
rect 12087 3950 12121 3984
rect 12156 3950 12190 3984
rect 12225 3950 12259 3984
rect 12294 3950 12328 3984
rect 12363 3950 12397 3984
rect 12432 3950 12466 3984
rect 12501 3950 12535 3984
rect 12570 3950 12604 3984
rect 12639 3950 12673 3984
rect 12708 3950 12742 3984
rect 12777 3950 12811 3984
rect 12846 3950 12880 3984
rect 12915 3950 12949 3984
rect 12984 3950 13018 3984
rect 13053 3950 13087 3984
rect 13122 3950 13156 3984
rect 13191 3950 13225 3984
rect 13260 3950 13294 3984
rect 13329 3950 13363 3984
rect 13398 3950 13432 3984
rect 13467 3950 13501 3984
rect 13536 3950 13570 3984
rect 13605 3950 13639 3984
rect 13674 3950 13708 3984
rect 13743 3950 13777 3984
rect 13812 3950 13846 3984
rect 13881 3950 13915 3984
rect 13950 3950 13984 3984
rect 14019 3950 14053 3984
rect 14088 3950 14122 3984
rect 14157 3950 14191 3984
rect 14226 3950 14260 3984
rect 14295 3950 14329 3984
rect 14364 3950 14398 3984
rect 14433 3950 14467 3984
rect 14502 3950 14536 3984
rect 14571 3950 14605 3984
rect 14640 3950 14674 3984
rect 14709 3950 14743 3984
rect 14778 3950 14812 3984
rect 14847 3950 14881 3984
rect 14916 3950 14950 3984
rect 14985 3950 15019 3984
rect 15054 3950 15088 3984
rect 15123 3950 15157 3984
rect 15192 3950 15226 3984
rect 15261 3950 15295 3984
rect 15330 3950 15364 3984
rect 15399 3950 15433 3984
rect 15468 3950 15502 3984
rect 15537 3950 15571 3984
rect 15606 3950 15640 3984
rect 15675 3950 15709 3984
rect 15744 3950 15778 3984
rect 15813 3950 15847 3984
rect 15882 3950 15916 3984
rect 15951 3950 15985 3984
rect 16020 3950 16054 3984
rect 16089 3950 16123 3984
rect 16158 3950 16192 3984
rect 16227 3950 16261 3984
rect 16296 3950 16330 3984
rect 11949 3882 11983 3916
rect 12018 3882 12052 3916
rect 12087 3882 12121 3916
rect 12156 3882 12190 3916
rect 12225 3882 12259 3916
rect 12294 3882 12328 3916
rect 12363 3882 12397 3916
rect 12432 3882 12466 3916
rect 12501 3882 12535 3916
rect 12570 3882 12604 3916
rect 12639 3882 12673 3916
rect 12708 3882 12742 3916
rect 12777 3882 12811 3916
rect 12846 3882 12880 3916
rect 12915 3882 12949 3916
rect 12984 3882 13018 3916
rect 13053 3882 13087 3916
rect 13122 3882 13156 3916
rect 13191 3882 13225 3916
rect 13260 3882 13294 3916
rect 13329 3882 13363 3916
rect 13398 3882 13432 3916
rect 13467 3882 13501 3916
rect 13536 3882 13570 3916
rect 13605 3882 13639 3916
rect 13674 3882 13708 3916
rect 13743 3882 13777 3916
rect 13812 3882 13846 3916
rect 13881 3882 13915 3916
rect 13950 3882 13984 3916
rect 14019 3882 14053 3916
rect 14088 3882 14122 3916
rect 14157 3882 14191 3916
rect 14226 3882 14260 3916
rect 14295 3882 14329 3916
rect 14364 3882 14398 3916
rect 14433 3882 14467 3916
rect 14502 3882 14536 3916
rect 14571 3882 14605 3916
rect 14640 3882 14674 3916
rect 14709 3882 14743 3916
rect 14778 3882 14812 3916
rect 14847 3882 14881 3916
rect 14916 3882 14950 3916
rect 14985 3882 15019 3916
rect 15054 3882 15088 3916
rect 15123 3882 15157 3916
rect 15192 3882 15226 3916
rect 15261 3882 15295 3916
rect 15330 3882 15364 3916
rect 15399 3882 15433 3916
rect 15468 3882 15502 3916
rect 15537 3882 15571 3916
rect 15606 3882 15640 3916
rect 15675 3882 15709 3916
rect 15744 3882 15778 3916
rect 15813 3882 15847 3916
rect 15882 3882 15916 3916
rect 15951 3882 15985 3916
rect 16020 3882 16054 3916
rect 16089 3882 16123 3916
rect 16158 3882 16192 3916
rect 16227 3882 16261 3916
rect 16296 3882 16330 3916
rect 11949 3814 11983 3848
rect 12018 3814 12052 3848
rect 12087 3814 12121 3848
rect 12156 3814 12190 3848
rect 12225 3814 12259 3848
rect 12294 3814 12328 3848
rect 12363 3814 12397 3848
rect 12432 3814 12466 3848
rect 12501 3814 12535 3848
rect 12570 3814 12604 3848
rect 12639 3814 12673 3848
rect 12708 3814 12742 3848
rect 12777 3814 12811 3848
rect 12846 3814 12880 3848
rect 12915 3814 12949 3848
rect 12984 3814 13018 3848
rect 13053 3814 13087 3848
rect 13122 3814 13156 3848
rect 13191 3814 13225 3848
rect 13260 3814 13294 3848
rect 13329 3814 13363 3848
rect 13398 3814 13432 3848
rect 13467 3814 13501 3848
rect 13536 3814 13570 3848
rect 13605 3814 13639 3848
rect 13674 3814 13708 3848
rect 13743 3814 13777 3848
rect 13812 3814 13846 3848
rect 13881 3814 13915 3848
rect 13950 3814 13984 3848
rect 14019 3814 14053 3848
rect 14088 3814 14122 3848
rect 14157 3814 14191 3848
rect 14226 3814 14260 3848
rect 14295 3814 14329 3848
rect 14364 3814 14398 3848
rect 14433 3814 14467 3848
rect 14502 3814 14536 3848
rect 14571 3814 14605 3848
rect 14640 3814 14674 3848
rect 14709 3814 14743 3848
rect 14778 3814 14812 3848
rect 14847 3814 14881 3848
rect 14916 3814 14950 3848
rect 14985 3814 15019 3848
rect 15054 3814 15088 3848
rect 15123 3814 15157 3848
rect 15192 3814 15226 3848
rect 15261 3814 15295 3848
rect 15330 3814 15364 3848
rect 15399 3814 15433 3848
rect 15468 3814 15502 3848
rect 15537 3814 15571 3848
rect 15606 3814 15640 3848
rect 15675 3814 15709 3848
rect 15744 3814 15778 3848
rect 15813 3814 15847 3848
rect 15882 3814 15916 3848
rect 15951 3814 15985 3848
rect 16020 3814 16054 3848
rect 16089 3814 16123 3848
rect 16158 3814 16192 3848
rect 16227 3814 16261 3848
rect 16296 3814 16330 3848
rect 11949 3746 11983 3780
rect 12018 3746 12052 3780
rect 12087 3746 12121 3780
rect 12156 3746 12190 3780
rect 12225 3746 12259 3780
rect 12294 3746 12328 3780
rect 12363 3746 12397 3780
rect 12432 3746 12466 3780
rect 12501 3746 12535 3780
rect 12570 3746 12604 3780
rect 12639 3746 12673 3780
rect 12708 3746 12742 3780
rect 12777 3746 12811 3780
rect 12846 3746 12880 3780
rect 12915 3746 12949 3780
rect 12984 3746 13018 3780
rect 13053 3746 13087 3780
rect 13122 3746 13156 3780
rect 13191 3746 13225 3780
rect 13260 3746 13294 3780
rect 13329 3746 13363 3780
rect 13398 3746 13432 3780
rect 13467 3746 13501 3780
rect 13536 3746 13570 3780
rect 13605 3746 13639 3780
rect 13674 3746 13708 3780
rect 13743 3746 13777 3780
rect 13812 3746 13846 3780
rect 13881 3746 13915 3780
rect 13950 3746 13984 3780
rect 14019 3746 14053 3780
rect 14088 3746 14122 3780
rect 14157 3746 14191 3780
rect 14226 3746 14260 3780
rect 14295 3746 14329 3780
rect 14364 3746 14398 3780
rect 14433 3746 14467 3780
rect 14502 3746 14536 3780
rect 14571 3746 14605 3780
rect 14640 3746 14674 3780
rect 14709 3746 14743 3780
rect 14778 3746 14812 3780
rect 14847 3746 14881 3780
rect 14916 3746 14950 3780
rect 14985 3746 15019 3780
rect 15054 3746 15088 3780
rect 15123 3746 15157 3780
rect 15192 3746 15226 3780
rect 15261 3746 15295 3780
rect 15330 3746 15364 3780
rect 15399 3746 15433 3780
rect 15468 3746 15502 3780
rect 15537 3746 15571 3780
rect 15606 3746 15640 3780
rect 15675 3746 15709 3780
rect 15744 3746 15778 3780
rect 15813 3746 15847 3780
rect 15882 3746 15916 3780
rect 15951 3746 15985 3780
rect 16020 3746 16054 3780
rect 16089 3746 16123 3780
rect 16158 3746 16192 3780
rect 16227 3746 16261 3780
rect 16296 3746 16330 3780
rect 11949 3678 11983 3712
rect 12018 3678 12052 3712
rect 12087 3678 12121 3712
rect 12156 3678 12190 3712
rect 12225 3678 12259 3712
rect 12294 3678 12328 3712
rect 12363 3678 12397 3712
rect 12432 3678 12466 3712
rect 12501 3678 12535 3712
rect 12570 3678 12604 3712
rect 12639 3678 12673 3712
rect 12708 3678 12742 3712
rect 12777 3678 12811 3712
rect 12846 3678 12880 3712
rect 12915 3678 12949 3712
rect 12984 3678 13018 3712
rect 13053 3678 13087 3712
rect 13122 3678 13156 3712
rect 13191 3678 13225 3712
rect 13260 3678 13294 3712
rect 13329 3678 13363 3712
rect 13398 3678 13432 3712
rect 13467 3678 13501 3712
rect 13536 3678 13570 3712
rect 13605 3678 13639 3712
rect 13674 3678 13708 3712
rect 13743 3678 13777 3712
rect 13812 3678 13846 3712
rect 13881 3678 13915 3712
rect 13950 3678 13984 3712
rect 14019 3678 14053 3712
rect 14088 3678 14122 3712
rect 14157 3678 14191 3712
rect 14226 3678 14260 3712
rect 14295 3678 14329 3712
rect 14364 3678 14398 3712
rect 14433 3678 14467 3712
rect 14502 3678 14536 3712
rect 14571 3678 14605 3712
rect 14640 3678 14674 3712
rect 14709 3678 14743 3712
rect 14778 3678 14812 3712
rect 14847 3678 14881 3712
rect 14916 3678 14950 3712
rect 14985 3678 15019 3712
rect 15054 3678 15088 3712
rect 15123 3678 15157 3712
rect 15192 3678 15226 3712
rect 15261 3678 15295 3712
rect 15330 3678 15364 3712
rect 15399 3678 15433 3712
rect 15468 3678 15502 3712
rect 15537 3678 15571 3712
rect 15606 3678 15640 3712
rect 15675 3678 15709 3712
rect 15744 3678 15778 3712
rect 15813 3678 15847 3712
rect 15882 3678 15916 3712
rect 15951 3678 15985 3712
rect 16020 3678 16054 3712
rect 16089 3678 16123 3712
rect 16158 3678 16192 3712
rect 16227 3678 16261 3712
rect 16296 3678 16330 3712
rect 11949 3610 11983 3644
rect 12018 3610 12052 3644
rect 12087 3610 12121 3644
rect 12156 3610 12190 3644
rect 12225 3610 12259 3644
rect 12294 3610 12328 3644
rect 12363 3610 12397 3644
rect 12432 3610 12466 3644
rect 12501 3610 12535 3644
rect 12570 3610 12604 3644
rect 12639 3610 12673 3644
rect 12708 3610 12742 3644
rect 12777 3610 12811 3644
rect 12846 3610 12880 3644
rect 12915 3610 12949 3644
rect 12984 3610 13018 3644
rect 13053 3610 13087 3644
rect 13122 3610 13156 3644
rect 13191 3610 13225 3644
rect 13260 3610 13294 3644
rect 13329 3610 13363 3644
rect 13398 3610 13432 3644
rect 13467 3610 13501 3644
rect 13536 3610 13570 3644
rect 13605 3610 13639 3644
rect 13674 3610 13708 3644
rect 13743 3610 13777 3644
rect 13812 3610 13846 3644
rect 13881 3610 13915 3644
rect 13950 3610 13984 3644
rect 14019 3610 14053 3644
rect 14088 3610 14122 3644
rect 14157 3610 14191 3644
rect 14226 3610 14260 3644
rect 14295 3610 14329 3644
rect 14364 3610 14398 3644
rect 14433 3610 14467 3644
rect 14502 3610 14536 3644
rect 14571 3610 14605 3644
rect 14640 3610 14674 3644
rect 14709 3610 14743 3644
rect 14778 3610 14812 3644
rect 14847 3610 14881 3644
rect 14916 3610 14950 3644
rect 14985 3610 15019 3644
rect 15054 3610 15088 3644
rect 15123 3610 15157 3644
rect 15192 3610 15226 3644
rect 15261 3610 15295 3644
rect 15330 3610 15364 3644
rect 15399 3610 15433 3644
rect 15468 3610 15502 3644
rect 15537 3610 15571 3644
rect 15606 3610 15640 3644
rect 15675 3610 15709 3644
rect 15744 3610 15778 3644
rect 15813 3610 15847 3644
rect 15882 3610 15916 3644
rect 15951 3610 15985 3644
rect 16020 3610 16054 3644
rect 16089 3610 16123 3644
rect 16158 3610 16192 3644
rect 16227 3610 16261 3644
rect 16296 3610 16330 3644
rect 11949 3542 11983 3576
rect 12018 3542 12052 3576
rect 12087 3542 12121 3576
rect 12156 3542 12190 3576
rect 12225 3542 12259 3576
rect 12294 3542 12328 3576
rect 12363 3542 12397 3576
rect 12432 3542 12466 3576
rect 12501 3542 12535 3576
rect 12570 3542 12604 3576
rect 12639 3542 12673 3576
rect 12708 3542 12742 3576
rect 12777 3542 12811 3576
rect 12846 3542 12880 3576
rect 12915 3542 12949 3576
rect 12984 3542 13018 3576
rect 13053 3542 13087 3576
rect 13122 3542 13156 3576
rect 13191 3542 13225 3576
rect 13260 3542 13294 3576
rect 13329 3542 13363 3576
rect 13398 3542 13432 3576
rect 13467 3542 13501 3576
rect 13536 3542 13570 3576
rect 13605 3542 13639 3576
rect 13674 3542 13708 3576
rect 13743 3542 13777 3576
rect 13812 3542 13846 3576
rect 13881 3542 13915 3576
rect 13950 3542 13984 3576
rect 14019 3542 14053 3576
rect 14088 3542 14122 3576
rect 14157 3542 14191 3576
rect 14226 3542 14260 3576
rect 14295 3542 14329 3576
rect 14364 3542 14398 3576
rect 14433 3542 14467 3576
rect 14502 3542 14536 3576
rect 14571 3542 14605 3576
rect 14640 3542 14674 3576
rect 14709 3542 14743 3576
rect 14778 3542 14812 3576
rect 14847 3542 14881 3576
rect 14916 3542 14950 3576
rect 14985 3542 15019 3576
rect 15054 3542 15088 3576
rect 15123 3542 15157 3576
rect 15192 3542 15226 3576
rect 15261 3542 15295 3576
rect 15330 3542 15364 3576
rect 15399 3542 15433 3576
rect 15468 3542 15502 3576
rect 15537 3542 15571 3576
rect 15606 3542 15640 3576
rect 15675 3542 15709 3576
rect 15744 3542 15778 3576
rect 15813 3542 15847 3576
rect 15882 3542 15916 3576
rect 15951 3542 15985 3576
rect 16020 3542 16054 3576
rect 16089 3542 16123 3576
rect 16158 3542 16192 3576
rect 16227 3542 16261 3576
rect 16296 3542 16330 3576
rect 11949 3474 11983 3508
rect 12018 3474 12052 3508
rect 12087 3474 12121 3508
rect 12156 3474 12190 3508
rect 12225 3474 12259 3508
rect 12294 3474 12328 3508
rect 12363 3474 12397 3508
rect 12432 3474 12466 3508
rect 12501 3474 12535 3508
rect 12570 3474 12604 3508
rect 12639 3474 12673 3508
rect 12708 3474 12742 3508
rect 12777 3474 12811 3508
rect 12846 3474 12880 3508
rect 12915 3474 12949 3508
rect 12984 3474 13018 3508
rect 13053 3474 13087 3508
rect 13122 3474 13156 3508
rect 13191 3474 13225 3508
rect 13260 3474 13294 3508
rect 13329 3474 13363 3508
rect 13398 3474 13432 3508
rect 13467 3474 13501 3508
rect 13536 3474 13570 3508
rect 13605 3474 13639 3508
rect 13674 3474 13708 3508
rect 13743 3474 13777 3508
rect 13812 3474 13846 3508
rect 13881 3474 13915 3508
rect 13950 3474 13984 3508
rect 14019 3474 14053 3508
rect 14088 3474 14122 3508
rect 14157 3474 14191 3508
rect 14226 3474 14260 3508
rect 14295 3474 14329 3508
rect 14364 3474 14398 3508
rect 14433 3474 14467 3508
rect 14502 3474 14536 3508
rect 14571 3474 14605 3508
rect 14640 3474 14674 3508
rect 14709 3474 14743 3508
rect 14778 3474 14812 3508
rect 14847 3474 14881 3508
rect 14916 3474 14950 3508
rect 14985 3474 15019 3508
rect 15054 3474 15088 3508
rect 15123 3474 15157 3508
rect 15192 3474 15226 3508
rect 15261 3474 15295 3508
rect 15330 3474 15364 3508
rect 15399 3474 15433 3508
rect 15468 3474 15502 3508
rect 15537 3474 15571 3508
rect 15606 3474 15640 3508
rect 15675 3474 15709 3508
rect 15744 3474 15778 3508
rect 15813 3474 15847 3508
rect 15882 3474 15916 3508
rect 15951 3474 15985 3508
rect 16020 3474 16054 3508
rect 16089 3474 16123 3508
rect 16158 3474 16192 3508
rect 16227 3474 16261 3508
rect 16296 3474 16330 3508
rect 11949 3406 11983 3440
rect 12018 3406 12052 3440
rect 12087 3406 12121 3440
rect 12156 3406 12190 3440
rect 12225 3406 12259 3440
rect 12294 3406 12328 3440
rect 12363 3406 12397 3440
rect 12432 3406 12466 3440
rect 12501 3406 12535 3440
rect 12570 3406 12604 3440
rect 12639 3406 12673 3440
rect 12708 3406 12742 3440
rect 12777 3406 12811 3440
rect 12846 3406 12880 3440
rect 12915 3406 12949 3440
rect 12984 3406 13018 3440
rect 13053 3406 13087 3440
rect 13122 3406 13156 3440
rect 13191 3406 13225 3440
rect 13260 3406 13294 3440
rect 13329 3406 13363 3440
rect 13398 3406 13432 3440
rect 13467 3406 13501 3440
rect 13536 3406 13570 3440
rect 13605 3406 13639 3440
rect 13674 3406 13708 3440
rect 13743 3406 13777 3440
rect 13812 3406 13846 3440
rect 13881 3406 13915 3440
rect 13950 3406 13984 3440
rect 14019 3406 14053 3440
rect 14088 3406 14122 3440
rect 14157 3406 14191 3440
rect 14226 3406 14260 3440
rect 14295 3406 14329 3440
rect 14364 3406 14398 3440
rect 14433 3406 14467 3440
rect 14502 3406 14536 3440
rect 14571 3406 14605 3440
rect 14640 3406 14674 3440
rect 14709 3406 14743 3440
rect 14778 3406 14812 3440
rect 14847 3406 14881 3440
rect 14916 3406 14950 3440
rect 14985 3406 15019 3440
rect 15054 3406 15088 3440
rect 15123 3406 15157 3440
rect 15192 3406 15226 3440
rect 15261 3406 15295 3440
rect 15330 3406 15364 3440
rect 15399 3406 15433 3440
rect 15468 3406 15502 3440
rect 15537 3406 15571 3440
rect 15606 3406 15640 3440
rect 15675 3406 15709 3440
rect 15744 3406 15778 3440
rect 15813 3406 15847 3440
rect 15882 3406 15916 3440
rect 15951 3406 15985 3440
rect 16020 3406 16054 3440
rect 16089 3406 16123 3440
rect 16158 3406 16192 3440
rect 16227 3406 16261 3440
rect 16296 3406 16330 3440
rect 11949 3338 11983 3372
rect 12018 3338 12052 3372
rect 12087 3338 12121 3372
rect 12156 3338 12190 3372
rect 12225 3338 12259 3372
rect 12294 3338 12328 3372
rect 12363 3338 12397 3372
rect 12432 3338 12466 3372
rect 12501 3338 12535 3372
rect 12570 3338 12604 3372
rect 12639 3338 12673 3372
rect 12708 3338 12742 3372
rect 12777 3338 12811 3372
rect 12846 3338 12880 3372
rect 12915 3338 12949 3372
rect 12984 3338 13018 3372
rect 13053 3338 13087 3372
rect 13122 3338 13156 3372
rect 13191 3338 13225 3372
rect 13260 3338 13294 3372
rect 13329 3338 13363 3372
rect 13398 3338 13432 3372
rect 13467 3338 13501 3372
rect 13536 3338 13570 3372
rect 13605 3338 13639 3372
rect 13674 3338 13708 3372
rect 13743 3338 13777 3372
rect 13812 3338 13846 3372
rect 13881 3338 13915 3372
rect 13950 3338 13984 3372
rect 14019 3338 14053 3372
rect 14088 3338 14122 3372
rect 14157 3338 14191 3372
rect 14226 3338 14260 3372
rect 14295 3338 14329 3372
rect 14364 3338 14398 3372
rect 14433 3338 14467 3372
rect 14502 3338 14536 3372
rect 14571 3338 14605 3372
rect 14640 3338 14674 3372
rect 14709 3338 14743 3372
rect 14778 3338 14812 3372
rect 14847 3338 14881 3372
rect 14916 3338 14950 3372
rect 14985 3338 15019 3372
rect 15054 3338 15088 3372
rect 15123 3338 15157 3372
rect 15192 3338 15226 3372
rect 15261 3338 15295 3372
rect 15330 3338 15364 3372
rect 15399 3338 15433 3372
rect 15468 3338 15502 3372
rect 15537 3338 15571 3372
rect 15606 3338 15640 3372
rect 15675 3338 15709 3372
rect 15744 3338 15778 3372
rect 15813 3338 15847 3372
rect 15882 3338 15916 3372
rect 15951 3338 15985 3372
rect 16020 3338 16054 3372
rect 16089 3338 16123 3372
rect 16158 3338 16192 3372
rect 16227 3338 16261 3372
rect 16296 3338 16330 3372
rect 11949 3270 11983 3304
rect 12018 3270 12052 3304
rect 12087 3270 12121 3304
rect 12156 3270 12190 3304
rect 12225 3270 12259 3304
rect 12294 3270 12328 3304
rect 12363 3270 12397 3304
rect 12432 3270 12466 3304
rect 12501 3270 12535 3304
rect 12570 3270 12604 3304
rect 12639 3270 12673 3304
rect 12708 3270 12742 3304
rect 12777 3270 12811 3304
rect 12846 3270 12880 3304
rect 12915 3270 12949 3304
rect 12984 3270 13018 3304
rect 13053 3270 13087 3304
rect 13122 3270 13156 3304
rect 13191 3270 13225 3304
rect 13260 3270 13294 3304
rect 13329 3270 13363 3304
rect 13398 3270 13432 3304
rect 13467 3270 13501 3304
rect 13536 3270 13570 3304
rect 13605 3270 13639 3304
rect 13674 3270 13708 3304
rect 13743 3270 13777 3304
rect 13812 3270 13846 3304
rect 13881 3270 13915 3304
rect 13950 3270 13984 3304
rect 14019 3270 14053 3304
rect 14088 3270 14122 3304
rect 14157 3270 14191 3304
rect 14226 3270 14260 3304
rect 14295 3270 14329 3304
rect 14364 3270 14398 3304
rect 14433 3270 14467 3304
rect 14502 3270 14536 3304
rect 14571 3270 14605 3304
rect 14640 3270 14674 3304
rect 14709 3270 14743 3304
rect 14778 3270 14812 3304
rect 14847 3270 14881 3304
rect 14916 3270 14950 3304
rect 14985 3270 15019 3304
rect 15054 3270 15088 3304
rect 15123 3270 15157 3304
rect 15192 3270 15226 3304
rect 15261 3270 15295 3304
rect 15330 3270 15364 3304
rect 15399 3270 15433 3304
rect 15468 3270 15502 3304
rect 15537 3270 15571 3304
rect 15606 3270 15640 3304
rect 15675 3270 15709 3304
rect 15744 3270 15778 3304
rect 15813 3270 15847 3304
rect 15882 3270 15916 3304
rect 15951 3270 15985 3304
rect 16020 3270 16054 3304
rect 16089 3270 16123 3304
rect 16158 3270 16192 3304
rect 16227 3270 16261 3304
rect 16296 3270 16330 3304
rect 16365 3270 17215 4324
rect 4639 3201 4673 3235
rect 4708 3201 4742 3235
rect 4777 3201 4811 3235
rect 4846 3201 4880 3235
rect 4915 3201 4949 3235
rect 4984 3201 5018 3235
rect 4639 3133 4673 3167
rect 4708 3133 4742 3167
rect 4777 3133 4811 3167
rect 4846 3133 4880 3167
rect 4915 3133 4949 3167
rect 4984 3133 5018 3167
rect 4639 3065 4673 3099
rect 4708 3065 4742 3099
rect 4777 3065 4811 3099
rect 4846 3065 4880 3099
rect 4915 3065 4949 3099
rect 4984 3065 5018 3099
rect 4639 2997 4673 3031
rect 4708 2997 4742 3031
rect 4777 2997 4811 3031
rect 4846 2997 4880 3031
rect 4915 2997 4949 3031
rect 4984 2997 5018 3031
rect 4639 2929 4673 2963
rect 4708 2929 4742 2963
rect 4777 2929 4811 2963
rect 4846 2929 4880 2963
rect 4915 2929 4949 2963
rect 4984 2929 5018 2963
rect 4639 2861 4673 2895
rect 4708 2861 4742 2895
rect 4777 2861 4811 2895
rect 4846 2861 4880 2895
rect 4915 2861 4949 2895
rect 4984 2861 5018 2895
rect 4639 2793 4673 2827
rect 4708 2793 4742 2827
rect 4777 2793 4811 2827
rect 4846 2793 4880 2827
rect 4915 2793 4949 2827
rect 4984 2793 5018 2827
rect 4639 2725 4673 2759
rect 4708 2725 4742 2759
rect 4777 2725 4811 2759
rect 4846 2725 4880 2759
rect 4915 2725 4949 2759
rect 4984 2725 5018 2759
rect 4639 2657 4673 2691
rect 4708 2657 4742 2691
rect 4777 2657 4811 2691
rect 4846 2657 4880 2691
rect 4915 2657 4949 2691
rect 4984 2657 5018 2691
rect 4639 2589 4673 2623
rect 4708 2589 4742 2623
rect 4777 2589 4811 2623
rect 4846 2589 4880 2623
rect 4915 2589 4949 2623
rect 4984 2589 5018 2623
rect 4639 2521 4673 2555
rect 4708 2521 4742 2555
rect 4777 2521 4811 2555
rect 4846 2521 4880 2555
rect 4915 2521 4949 2555
rect 4984 2521 5018 2555
rect 4639 2453 4673 2487
rect 4708 2453 4742 2487
rect 4777 2453 4811 2487
rect 4846 2453 4880 2487
rect 4915 2453 4949 2487
rect 4984 2453 5018 2487
rect 4639 2385 4673 2419
rect 4708 2385 4742 2419
rect 4777 2385 4811 2419
rect 4846 2385 4880 2419
rect 4915 2385 4949 2419
rect 4984 2385 5018 2419
rect 4639 2317 4673 2351
rect 4708 2317 4742 2351
rect 4777 2317 4811 2351
rect 4846 2317 4880 2351
rect 4915 2317 4949 2351
rect 4984 2317 5018 2351
rect 4639 2249 4673 2283
rect 4708 2249 4742 2283
rect 4777 2249 4811 2283
rect 4846 2249 4880 2283
rect 4915 2249 4949 2283
rect 4984 2249 5018 2283
rect 4639 2181 4673 2215
rect 4708 2181 4742 2215
rect 4777 2181 4811 2215
rect 4846 2181 4880 2215
rect 4915 2181 4949 2215
rect 4984 2181 5018 2215
rect 5053 2181 17191 3235
rect 4615 2113 4649 2147
rect 4686 2113 4720 2147
rect 4757 2113 4791 2147
rect 4828 2113 4862 2147
rect 4899 2113 4933 2147
rect 4970 2113 5004 2147
rect 5041 2113 5075 2147
rect 5112 2113 5146 2147
rect 5183 2113 5217 2147
rect 5254 2113 5288 2147
rect 5325 2113 5359 2147
rect 5396 2113 5430 2147
rect 5467 2113 5501 2147
rect 5537 2113 5571 2147
rect 5607 2113 5641 2147
rect 5677 2113 5711 2147
rect 4615 2037 4649 2071
rect 4686 2037 4720 2071
rect 4757 2037 4791 2071
rect 4828 2037 4862 2071
rect 4899 2037 4933 2071
rect 4970 2037 5004 2071
rect 5041 2037 5075 2071
rect 5112 2037 5146 2071
rect 5183 2037 5217 2071
rect 5254 2037 5288 2071
rect 5325 2037 5359 2071
rect 5396 2037 5430 2071
rect 5467 2037 5501 2071
rect 5537 2037 5571 2071
rect 5607 2037 5641 2071
rect 5677 2037 5711 2071
rect 4615 1961 4649 1995
rect 4686 1961 4720 1995
rect 4757 1961 4791 1995
rect 4828 1961 4862 1995
rect 4899 1961 4933 1995
rect 4970 1961 5004 1995
rect 5041 1961 5075 1995
rect 5112 1961 5146 1995
rect 5183 1961 5217 1995
rect 5254 1961 5288 1995
rect 5325 1961 5359 1995
rect 5396 1961 5430 1995
rect 5467 1961 5501 1995
rect 5537 1961 5571 1995
rect 5607 1961 5641 1995
rect 5677 1961 5711 1995
rect 4615 1885 4649 1919
rect 4686 1885 4720 1919
rect 4757 1885 4791 1919
rect 4828 1885 4862 1919
rect 4899 1885 4933 1919
rect 4970 1885 5004 1919
rect 5041 1885 5075 1919
rect 5112 1885 5146 1919
rect 5183 1885 5217 1919
rect 5254 1885 5288 1919
rect 5325 1885 5359 1919
rect 5396 1885 5430 1919
rect 5467 1885 5501 1919
rect 5537 1885 5571 1919
rect 5607 1885 5641 1919
rect 5677 1885 5711 1919
rect 33 792 5711 1846
rect 10596 916 10630 950
rect 10665 916 10699 950
rect 10734 916 10768 950
rect 10803 916 10837 950
rect 10872 916 10906 950
rect 10941 916 10975 950
rect 11010 916 11044 950
rect 11078 916 11112 950
rect 11146 916 11180 950
rect 11214 916 11248 950
rect 11282 916 11316 950
rect 11350 916 11384 950
rect 11418 916 11452 950
rect 11486 916 11520 950
rect 11554 916 11588 950
rect 11622 916 11656 950
rect 11690 916 11724 950
rect 11758 916 11792 950
rect 11826 916 11860 950
rect 11894 916 11928 950
rect 11962 916 11996 950
rect 12030 916 12064 950
rect 12098 916 12132 950
rect 12166 916 12200 950
rect 12234 916 12268 950
rect 12302 916 12336 950
rect 12370 916 12404 950
rect 12438 916 12472 950
rect 12506 916 12540 950
rect 12574 916 12608 950
rect 12642 916 12676 950
rect 12710 916 12744 950
rect 12778 916 12812 950
rect 12846 916 12880 950
rect 12914 916 12948 950
rect 12982 916 13016 950
rect 13050 916 13084 950
rect 13118 916 13152 950
rect 13186 916 13220 950
rect 13254 916 13288 950
rect 13322 916 13356 950
rect 13390 916 13424 950
rect 13458 916 13492 950
rect 13526 916 13560 950
rect 13594 916 13628 950
rect 13662 916 13696 950
rect 13730 916 13764 950
rect 13798 916 13832 950
rect 13866 916 13900 950
rect 13934 916 13968 950
rect 14002 916 14036 950
rect 14070 916 14104 950
rect 14138 916 14172 950
rect 14206 916 14240 950
rect 14274 916 14308 950
rect 14342 916 14376 950
rect 14410 916 14444 950
rect 14478 916 14512 950
rect 14546 916 14580 950
rect 14614 916 14648 950
rect 14682 916 14716 950
rect 14750 916 14784 950
rect 14818 916 14852 950
rect 14886 916 14920 950
rect 6576 798 6610 832
rect 6645 798 6679 832
rect 6714 798 6748 832
rect 6783 798 6817 832
rect 6852 798 6886 832
rect 6921 798 6955 832
rect 6990 798 7024 832
rect 7059 798 7093 832
rect 7128 798 7162 832
rect 7197 798 7231 832
rect 7266 798 7300 832
rect 7335 798 7369 832
rect 7404 798 7438 832
rect 7473 798 7507 832
rect 7542 798 7576 832
rect 7611 798 7645 832
rect 7680 798 7714 832
rect 7749 798 7783 832
rect 7818 798 7852 832
rect 7887 798 7921 832
rect 7956 798 7990 832
rect 8025 798 8059 832
rect 8094 798 8128 832
rect 8162 798 8196 832
rect 8230 798 8264 832
rect 8298 798 8332 832
rect 8366 798 8400 832
rect 8434 798 8468 832
rect 8502 798 8536 832
rect 8570 798 8604 832
rect 8638 798 8672 832
rect 8706 798 8740 832
rect 8774 798 8808 832
rect 8842 798 8876 832
rect 8910 798 8944 832
rect 8978 798 9012 832
rect 9046 798 9080 832
rect 9114 798 9148 832
rect 9182 798 9216 832
rect 9250 798 9284 832
rect 9318 798 9352 832
rect 9386 798 9420 832
rect 9454 798 9488 832
rect 9522 798 9556 832
rect 9590 798 9624 832
rect 9658 798 9692 832
rect 9726 798 9760 832
rect 9794 798 9828 832
rect 9862 798 9896 832
rect 9930 798 9964 832
rect 9998 798 10032 832
rect 10066 798 10100 832
rect 10134 798 10168 832
rect 10202 798 10236 832
rect 10270 798 10304 832
rect 10338 798 10372 832
rect 10406 798 10440 832
rect 10474 798 10508 832
rect 15944 -2511 16726 2181
rect 15944 -2580 15978 -2546
rect 16012 -2580 16046 -2546
rect 16080 -2580 16114 -2546
rect 16148 -2580 16182 -2546
rect 16216 -2580 16250 -2546
rect 16284 -2580 16318 -2546
rect 16352 -2580 16386 -2546
rect 16420 -2580 16454 -2546
rect 16488 -2580 16522 -2546
rect 16556 -2580 16590 -2546
rect 16624 -2580 16658 -2546
rect 16692 -2580 16726 -2546
rect 15944 -2649 15978 -2615
rect 16012 -2649 16046 -2615
rect 16080 -2649 16114 -2615
rect 16148 -2649 16182 -2615
rect 16216 -2649 16250 -2615
rect 16284 -2649 16318 -2615
rect 16352 -2649 16386 -2615
rect 16420 -2649 16454 -2615
rect 16488 -2649 16522 -2615
rect 16556 -2649 16590 -2615
rect 16624 -2649 16658 -2615
rect 16692 -2649 16726 -2615
rect 15944 -2718 15978 -2684
rect 16012 -2718 16046 -2684
rect 16080 -2718 16114 -2684
rect 16148 -2718 16182 -2684
rect 16216 -2718 16250 -2684
rect 16284 -2718 16318 -2684
rect 16352 -2718 16386 -2684
rect 16420 -2718 16454 -2684
rect 16488 -2718 16522 -2684
rect 16556 -2718 16590 -2684
rect 16624 -2718 16658 -2684
rect 16692 -2718 16726 -2684
rect 15944 -2787 15978 -2753
rect 16012 -2787 16046 -2753
rect 16080 -2787 16114 -2753
rect 16148 -2787 16182 -2753
rect 16216 -2787 16250 -2753
rect 16284 -2787 16318 -2753
rect 16352 -2787 16386 -2753
rect 16420 -2787 16454 -2753
rect 16488 -2787 16522 -2753
rect 16556 -2787 16590 -2753
rect 16624 -2787 16658 -2753
rect 16692 -2787 16726 -2753
rect 15944 -2856 15978 -2822
rect 16012 -2856 16046 -2822
rect 16080 -2856 16114 -2822
rect 16148 -2856 16182 -2822
rect 16216 -2856 16250 -2822
rect 16284 -2856 16318 -2822
rect 16352 -2856 16386 -2822
rect 16420 -2856 16454 -2822
rect 16488 -2856 16522 -2822
rect 16556 -2856 16590 -2822
rect 16624 -2856 16658 -2822
rect 16692 -2856 16726 -2822
rect 15944 -2925 15978 -2891
rect 16012 -2925 16046 -2891
rect 16080 -2925 16114 -2891
rect 16148 -2925 16182 -2891
rect 16216 -2925 16250 -2891
rect 16284 -2925 16318 -2891
rect 16352 -2925 16386 -2891
rect 16420 -2925 16454 -2891
rect 16488 -2925 16522 -2891
rect 16556 -2925 16590 -2891
rect 16624 -2925 16658 -2891
rect 16692 -2925 16726 -2891
<< mvnsubdiffcont >>
rect -2750 4464 -2716 4498
rect -2680 4464 -2646 4498
rect -2610 4464 -2576 4498
rect -2540 4464 -2506 4498
rect -2470 4464 -2436 4498
rect -2400 4464 -2366 4498
rect -2330 4464 -2296 4498
rect -2260 4464 -2226 4498
rect -2190 4464 -2156 4498
rect -2120 4464 -2086 4498
rect -2050 4464 -2016 4498
rect -1980 4464 -1946 4498
rect -1910 4464 -1876 4498
rect -1840 4464 -1806 4498
rect -1770 4464 -1736 4498
rect -1700 4464 -1666 4498
rect -1630 4464 -1596 4498
rect -1560 4464 -1526 4498
rect -1490 4464 -1456 4498
rect -1421 4464 -1387 4498
rect -1352 4464 -1318 4498
rect -1283 4464 -1249 4498
rect -1214 4464 -1180 4498
rect -1145 4464 -1111 4498
rect -1076 4464 -1042 4498
rect -1007 4464 -973 4498
rect -938 4464 -904 4498
rect -869 4464 -835 4498
rect -800 4464 -766 4498
rect -731 4464 -697 4498
rect -662 4464 -628 4498
rect -593 4464 -559 4498
rect -524 4464 -490 4498
rect -455 4464 -421 4498
rect -386 4464 -352 4498
rect -317 4464 -283 4498
rect -248 4464 -214 4498
rect -2750 4394 -2716 4428
rect -2680 4394 -2646 4428
rect -2610 4394 -2576 4428
rect -2540 4394 -2506 4428
rect -2470 4394 -2436 4428
rect -2400 4394 -2366 4428
rect -2330 4394 -2296 4428
rect -2260 4394 -2226 4428
rect -2190 4394 -2156 4428
rect -2120 4394 -2086 4428
rect -2050 4394 -2016 4428
rect -1980 4394 -1946 4428
rect -1910 4394 -1876 4428
rect -1840 4394 -1806 4428
rect -1770 4394 -1736 4428
rect -1700 4394 -1666 4428
rect -1630 4394 -1596 4428
rect -1560 4394 -1526 4428
rect -1490 4394 -1456 4428
rect -1421 4394 -1387 4428
rect -1352 4394 -1318 4428
rect -1283 4394 -1249 4428
rect -1214 4394 -1180 4428
rect -1145 4394 -1111 4428
rect -1076 4394 -1042 4428
rect -1007 4394 -973 4428
rect -938 4394 -904 4428
rect -869 4394 -835 4428
rect -800 4394 -766 4428
rect -731 4394 -697 4428
rect -662 4394 -628 4428
rect -593 4394 -559 4428
rect -524 4394 -490 4428
rect -455 4394 -421 4428
rect -386 4394 -352 4428
rect -317 4394 -283 4428
rect -248 4394 -214 4428
rect -2750 4324 -2716 4358
rect -2680 4324 -2646 4358
rect -2610 4324 -2576 4358
rect -2540 4324 -2506 4358
rect -2470 4324 -2436 4358
rect -2400 4324 -2366 4358
rect -2330 4324 -2296 4358
rect -2260 4324 -2226 4358
rect -2190 4324 -2156 4358
rect -2120 4324 -2086 4358
rect -2050 4324 -2016 4358
rect -1980 4324 -1946 4358
rect -1910 4324 -1876 4358
rect -1840 4324 -1806 4358
rect -1770 4324 -1736 4358
rect -1700 4324 -1666 4358
rect -1630 4324 -1596 4358
rect -1560 4324 -1526 4358
rect -1490 4324 -1456 4358
rect -1421 4324 -1387 4358
rect -1352 4324 -1318 4358
rect -1283 4324 -1249 4358
rect -1214 4324 -1180 4358
rect -1145 4324 -1111 4358
rect -1076 4324 -1042 4358
rect -1007 4324 -973 4358
rect -938 4324 -904 4358
rect -869 4324 -835 4358
rect -800 4324 -766 4358
rect -731 4324 -697 4358
rect -662 4324 -628 4358
rect -593 4324 -559 4358
rect -524 4324 -490 4358
rect -455 4324 -421 4358
rect -386 4324 -352 4358
rect -317 4324 -283 4358
rect -248 4324 -214 4358
rect -2750 4254 -2716 4288
rect -2680 4254 -2646 4288
rect -2610 4254 -2576 4288
rect -2540 4254 -2506 4288
rect -2470 4254 -2436 4288
rect -2400 4254 -2366 4288
rect -2330 4254 -2296 4288
rect -2260 4254 -2226 4288
rect -2190 4254 -2156 4288
rect -2120 4254 -2086 4288
rect -2050 4254 -2016 4288
rect -1980 4254 -1946 4288
rect -1910 4254 -1876 4288
rect -1840 4254 -1806 4288
rect -1770 4254 -1736 4288
rect -1700 4254 -1666 4288
rect -1630 4254 -1596 4288
rect -1560 4254 -1526 4288
rect -1490 4254 -1456 4288
rect -1421 4254 -1387 4288
rect -1352 4254 -1318 4288
rect -1283 4254 -1249 4288
rect -1214 4254 -1180 4288
rect -1145 4254 -1111 4288
rect -1076 4254 -1042 4288
rect -1007 4254 -973 4288
rect -938 4254 -904 4288
rect -869 4254 -835 4288
rect -800 4254 -766 4288
rect -731 4254 -697 4288
rect -662 4254 -628 4288
rect -593 4254 -559 4288
rect -524 4254 -490 4288
rect -455 4254 -421 4288
rect -386 4254 -352 4288
rect -317 4254 -283 4288
rect -248 4254 -214 4288
rect -2750 4184 -2716 4218
rect -2680 4184 -2646 4218
rect -2610 4184 -2576 4218
rect -2540 4184 -2506 4218
rect -2470 4184 -2436 4218
rect -2400 4184 -2366 4218
rect -2330 4184 -2296 4218
rect -2260 4184 -2226 4218
rect -2190 4184 -2156 4218
rect -2120 4184 -2086 4218
rect -2050 4184 -2016 4218
rect -1980 4184 -1946 4218
rect -1910 4184 -1876 4218
rect -1840 4184 -1806 4218
rect -1770 4184 -1736 4218
rect -1700 4184 -1666 4218
rect -1630 4184 -1596 4218
rect -1560 4184 -1526 4218
rect -1490 4184 -1456 4218
rect -1421 4184 -1387 4218
rect -1352 4184 -1318 4218
rect -1283 4184 -1249 4218
rect -1214 4184 -1180 4218
rect -1145 4184 -1111 4218
rect -1076 4184 -1042 4218
rect -1007 4184 -973 4218
rect -938 4184 -904 4218
rect -869 4184 -835 4218
rect -800 4184 -766 4218
rect -731 4184 -697 4218
rect -662 4184 -628 4218
rect -593 4184 -559 4218
rect -524 4184 -490 4218
rect -455 4184 -421 4218
rect -386 4184 -352 4218
rect -317 4184 -283 4218
rect -248 4184 -214 4218
rect -2750 4114 -2716 4148
rect -2680 4114 -2646 4148
rect -2610 4114 -2576 4148
rect -2540 4114 -2506 4148
rect -2470 4114 -2436 4148
rect -2400 4114 -2366 4148
rect -2330 4114 -2296 4148
rect -2260 4114 -2226 4148
rect -2190 4114 -2156 4148
rect -2120 4114 -2086 4148
rect -2050 4114 -2016 4148
rect -1980 4114 -1946 4148
rect -1910 4114 -1876 4148
rect -1840 4114 -1806 4148
rect -1770 4114 -1736 4148
rect -1700 4114 -1666 4148
rect -1630 4114 -1596 4148
rect -1560 4114 -1526 4148
rect -1490 4114 -1456 4148
rect -1421 4114 -1387 4148
rect -1352 4114 -1318 4148
rect -1283 4114 -1249 4148
rect -1214 4114 -1180 4148
rect -1145 4114 -1111 4148
rect -1076 4114 -1042 4148
rect -1007 4114 -973 4148
rect -938 4114 -904 4148
rect -869 4114 -835 4148
rect -800 4114 -766 4148
rect -731 4114 -697 4148
rect -662 4114 -628 4148
rect -593 4114 -559 4148
rect -524 4114 -490 4148
rect -455 4114 -421 4148
rect -386 4114 -352 4148
rect -317 4114 -283 4148
rect -248 4114 -214 4148
rect -2750 4044 -2716 4078
rect -2680 4044 -2646 4078
rect -2610 4044 -2576 4078
rect -2540 4044 -2506 4078
rect -2470 4044 -2436 4078
rect -2400 4044 -2366 4078
rect -2330 4044 -2296 4078
rect -2260 4044 -2226 4078
rect -2190 4044 -2156 4078
rect -2120 4044 -2086 4078
rect -2050 4044 -2016 4078
rect -1980 4044 -1946 4078
rect -1910 4044 -1876 4078
rect -1840 4044 -1806 4078
rect -1770 4044 -1736 4078
rect -1700 4044 -1666 4078
rect -1630 4044 -1596 4078
rect -1560 4044 -1526 4078
rect -1490 4044 -1456 4078
rect -1421 4044 -1387 4078
rect -1352 4044 -1318 4078
rect -1283 4044 -1249 4078
rect -1214 4044 -1180 4078
rect -1145 4044 -1111 4078
rect -1076 4044 -1042 4078
rect -1007 4044 -973 4078
rect -938 4044 -904 4078
rect -869 4044 -835 4078
rect -800 4044 -766 4078
rect -731 4044 -697 4078
rect -662 4044 -628 4078
rect -593 4044 -559 4078
rect -524 4044 -490 4078
rect -455 4044 -421 4078
rect -386 4044 -352 4078
rect -317 4044 -283 4078
rect -248 4044 -214 4078
rect -2750 3974 -2716 4008
rect -2680 3974 -2646 4008
rect -2610 3974 -2576 4008
rect -2540 3974 -2506 4008
rect -2470 3974 -2436 4008
rect -2400 3974 -2366 4008
rect -2330 3974 -2296 4008
rect -2260 3974 -2226 4008
rect -2190 3974 -2156 4008
rect -2120 3974 -2086 4008
rect -2050 3974 -2016 4008
rect -1980 3974 -1946 4008
rect -1910 3974 -1876 4008
rect -1840 3974 -1806 4008
rect -1770 3974 -1736 4008
rect -1700 3974 -1666 4008
rect -1630 3974 -1596 4008
rect -1560 3974 -1526 4008
rect -1490 3974 -1456 4008
rect -1421 3974 -1387 4008
rect -1352 3974 -1318 4008
rect -1283 3974 -1249 4008
rect -1214 3974 -1180 4008
rect -1145 3974 -1111 4008
rect -1076 3974 -1042 4008
rect -1007 3974 -973 4008
rect -938 3974 -904 4008
rect -869 3974 -835 4008
rect -800 3974 -766 4008
rect -731 3974 -697 4008
rect -662 3974 -628 4008
rect -593 3974 -559 4008
rect -524 3974 -490 4008
rect -455 3974 -421 4008
rect -386 3974 -352 4008
rect -317 3974 -283 4008
rect -248 3974 -214 4008
rect -2750 3904 -2716 3938
rect -2680 3904 -2646 3938
rect -2610 3904 -2576 3938
rect -2540 3904 -2506 3938
rect -2470 3904 -2436 3938
rect -2400 3904 -2366 3938
rect -2330 3904 -2296 3938
rect -2260 3904 -2226 3938
rect -2190 3904 -2156 3938
rect -2120 3904 -2086 3938
rect -2050 3904 -2016 3938
rect -1980 3904 -1946 3938
rect -1910 3904 -1876 3938
rect -1840 3904 -1806 3938
rect -1770 3904 -1736 3938
rect -1700 3904 -1666 3938
rect -1630 3904 -1596 3938
rect -1560 3904 -1526 3938
rect -1490 3904 -1456 3938
rect -1421 3904 -1387 3938
rect -1352 3904 -1318 3938
rect -1283 3904 -1249 3938
rect -1214 3904 -1180 3938
rect -1145 3904 -1111 3938
rect -1076 3904 -1042 3938
rect -1007 3904 -973 3938
rect -938 3904 -904 3938
rect -869 3904 -835 3938
rect -800 3904 -766 3938
rect -731 3904 -697 3938
rect -662 3904 -628 3938
rect -593 3904 -559 3938
rect -524 3904 -490 3938
rect -455 3904 -421 3938
rect -386 3904 -352 3938
rect -317 3904 -283 3938
rect -248 3904 -214 3938
rect -2750 3834 -2716 3868
rect -2680 3834 -2646 3868
rect -2610 3834 -2576 3868
rect -2540 3834 -2506 3868
rect -2470 3834 -2436 3868
rect -2400 3834 -2366 3868
rect -2330 3834 -2296 3868
rect -2260 3834 -2226 3868
rect -2190 3834 -2156 3868
rect -2120 3834 -2086 3868
rect -2050 3834 -2016 3868
rect -1980 3834 -1946 3868
rect -1910 3834 -1876 3868
rect -1840 3834 -1806 3868
rect -1770 3834 -1736 3868
rect -1700 3834 -1666 3868
rect -1630 3834 -1596 3868
rect -1560 3834 -1526 3868
rect -1490 3834 -1456 3868
rect -1421 3834 -1387 3868
rect -1352 3834 -1318 3868
rect -1283 3834 -1249 3868
rect -1214 3834 -1180 3868
rect -1145 3834 -1111 3868
rect -1076 3834 -1042 3868
rect -1007 3834 -973 3868
rect -938 3834 -904 3868
rect -869 3834 -835 3868
rect -800 3834 -766 3868
rect -731 3834 -697 3868
rect -662 3834 -628 3868
rect -593 3834 -559 3868
rect -524 3834 -490 3868
rect -455 3834 -421 3868
rect -386 3834 -352 3868
rect -317 3834 -283 3868
rect -248 3834 -214 3868
rect -2750 3764 -2716 3798
rect -2680 3764 -2646 3798
rect -2610 3764 -2576 3798
rect -2540 3764 -2506 3798
rect -2470 3764 -2436 3798
rect -2400 3764 -2366 3798
rect -2330 3764 -2296 3798
rect -2260 3764 -2226 3798
rect -2190 3764 -2156 3798
rect -2120 3764 -2086 3798
rect -2050 3764 -2016 3798
rect -1980 3764 -1946 3798
rect -1910 3764 -1876 3798
rect -1840 3764 -1806 3798
rect -1770 3764 -1736 3798
rect -1700 3764 -1666 3798
rect -1630 3764 -1596 3798
rect -1560 3764 -1526 3798
rect -1490 3764 -1456 3798
rect -1421 3764 -1387 3798
rect -1352 3764 -1318 3798
rect -1283 3764 -1249 3798
rect -1214 3764 -1180 3798
rect -1145 3764 -1111 3798
rect -1076 3764 -1042 3798
rect -1007 3764 -973 3798
rect -938 3764 -904 3798
rect -869 3764 -835 3798
rect -800 3764 -766 3798
rect -731 3764 -697 3798
rect -662 3764 -628 3798
rect -593 3764 -559 3798
rect -524 3764 -490 3798
rect -455 3764 -421 3798
rect -386 3764 -352 3798
rect -317 3764 -283 3798
rect -248 3764 -214 3798
rect -2750 3694 -2716 3728
rect -2680 3694 -2646 3728
rect -2610 3694 -2576 3728
rect -2540 3694 -2506 3728
rect -2470 3694 -2436 3728
rect -2400 3694 -2366 3728
rect -2330 3694 -2296 3728
rect -2260 3694 -2226 3728
rect -2190 3694 -2156 3728
rect -2120 3694 -2086 3728
rect -2050 3694 -2016 3728
rect -1980 3694 -1946 3728
rect -1910 3694 -1876 3728
rect -1840 3694 -1806 3728
rect -1770 3694 -1736 3728
rect -1700 3694 -1666 3728
rect -1630 3694 -1596 3728
rect -1560 3694 -1526 3728
rect -1490 3694 -1456 3728
rect -1421 3694 -1387 3728
rect -1352 3694 -1318 3728
rect -1283 3694 -1249 3728
rect -1214 3694 -1180 3728
rect -1145 3694 -1111 3728
rect -1076 3694 -1042 3728
rect -1007 3694 -973 3728
rect -938 3694 -904 3728
rect -869 3694 -835 3728
rect -800 3694 -766 3728
rect -731 3694 -697 3728
rect -662 3694 -628 3728
rect -593 3694 -559 3728
rect -524 3694 -490 3728
rect -455 3694 -421 3728
rect -386 3694 -352 3728
rect -317 3694 -283 3728
rect -248 3694 -214 3728
rect -2750 3624 -2716 3658
rect -2680 3624 -2646 3658
rect -2610 3624 -2576 3658
rect -2540 3624 -2506 3658
rect -2470 3624 -2436 3658
rect -2400 3624 -2366 3658
rect -2330 3624 -2296 3658
rect -2260 3624 -2226 3658
rect -2190 3624 -2156 3658
rect -2120 3624 -2086 3658
rect -2050 3624 -2016 3658
rect -1980 3624 -1946 3658
rect -1910 3624 -1876 3658
rect -1840 3624 -1806 3658
rect -1770 3624 -1736 3658
rect -1700 3624 -1666 3658
rect -1630 3624 -1596 3658
rect -1560 3624 -1526 3658
rect -1490 3624 -1456 3658
rect -1421 3624 -1387 3658
rect -1352 3624 -1318 3658
rect -1283 3624 -1249 3658
rect -1214 3624 -1180 3658
rect -1145 3624 -1111 3658
rect -1076 3624 -1042 3658
rect -1007 3624 -973 3658
rect -938 3624 -904 3658
rect -869 3624 -835 3658
rect -800 3624 -766 3658
rect -731 3624 -697 3658
rect -662 3624 -628 3658
rect -593 3624 -559 3658
rect -524 3624 -490 3658
rect -455 3624 -421 3658
rect -386 3624 -352 3658
rect -317 3624 -283 3658
rect -248 3624 -214 3658
rect -2750 3554 -2716 3588
rect -2680 3554 -2646 3588
rect -2610 3554 -2576 3588
rect -2540 3554 -2506 3588
rect -2470 3554 -2436 3588
rect -2400 3554 -2366 3588
rect -2330 3554 -2296 3588
rect -2260 3554 -2226 3588
rect -2190 3554 -2156 3588
rect -2120 3554 -2086 3588
rect -2050 3554 -2016 3588
rect -1980 3554 -1946 3588
rect -1910 3554 -1876 3588
rect -1840 3554 -1806 3588
rect -1770 3554 -1736 3588
rect -1700 3554 -1666 3588
rect -1630 3554 -1596 3588
rect -1560 3554 -1526 3588
rect -1490 3554 -1456 3588
rect -1421 3554 -1387 3588
rect -1352 3554 -1318 3588
rect -1283 3554 -1249 3588
rect -1214 3554 -1180 3588
rect -1145 3554 -1111 3588
rect -1076 3554 -1042 3588
rect -1007 3554 -973 3588
rect -938 3554 -904 3588
rect -869 3554 -835 3588
rect -800 3554 -766 3588
rect -731 3554 -697 3588
rect -662 3554 -628 3588
rect -593 3554 -559 3588
rect -524 3554 -490 3588
rect -455 3554 -421 3588
rect -386 3554 -352 3588
rect -317 3554 -283 3588
rect -248 3554 -214 3588
rect -2750 3484 -2716 3518
rect -2680 3484 -2646 3518
rect -2610 3484 -2576 3518
rect -2540 3484 -2506 3518
rect -2470 3484 -2436 3518
rect -2400 3484 -2366 3518
rect -2330 3484 -2296 3518
rect -2260 3484 -2226 3518
rect -2190 3484 -2156 3518
rect -2120 3484 -2086 3518
rect -2050 3484 -2016 3518
rect -1980 3484 -1946 3518
rect -1910 3484 -1876 3518
rect -1840 3484 -1806 3518
rect -1770 3484 -1736 3518
rect -1700 3484 -1666 3518
rect -1630 3484 -1596 3518
rect -1560 3484 -1526 3518
rect -1490 3484 -1456 3518
rect -1421 3484 -1387 3518
rect -1352 3484 -1318 3518
rect -1283 3484 -1249 3518
rect -1214 3484 -1180 3518
rect -1145 3484 -1111 3518
rect -1076 3484 -1042 3518
rect -1007 3484 -973 3518
rect -938 3484 -904 3518
rect -869 3484 -835 3518
rect -800 3484 -766 3518
rect -731 3484 -697 3518
rect -662 3484 -628 3518
rect -593 3484 -559 3518
rect -524 3484 -490 3518
rect -455 3484 -421 3518
rect -386 3484 -352 3518
rect -317 3484 -283 3518
rect -248 3484 -214 3518
rect -2750 3414 -2716 3448
rect -2680 3414 -2646 3448
rect -2610 3414 -2576 3448
rect -2540 3414 -2506 3448
rect -2470 3414 -2436 3448
rect -2400 3414 -2366 3448
rect -2330 3414 -2296 3448
rect -2260 3414 -2226 3448
rect -2190 3414 -2156 3448
rect -2120 3414 -2086 3448
rect -2050 3414 -2016 3448
rect -1980 3414 -1946 3448
rect -1910 3414 -1876 3448
rect -1840 3414 -1806 3448
rect -1770 3414 -1736 3448
rect -1700 3414 -1666 3448
rect -1630 3414 -1596 3448
rect -1560 3414 -1526 3448
rect -1490 3414 -1456 3448
rect -1421 3414 -1387 3448
rect -1352 3414 -1318 3448
rect -1283 3414 -1249 3448
rect -1214 3414 -1180 3448
rect -1145 3414 -1111 3448
rect -1076 3414 -1042 3448
rect -1007 3414 -973 3448
rect -938 3414 -904 3448
rect -869 3414 -835 3448
rect -800 3414 -766 3448
rect -731 3414 -697 3448
rect -662 3414 -628 3448
rect -593 3414 -559 3448
rect -524 3414 -490 3448
rect -455 3414 -421 3448
rect -386 3414 -352 3448
rect -317 3414 -283 3448
rect -248 3414 -214 3448
rect -2750 3344 -2716 3378
rect -2680 3344 -2646 3378
rect -2610 3344 -2576 3378
rect -2540 3344 -2506 3378
rect -2470 3344 -2436 3378
rect -2400 3344 -2366 3378
rect -2330 3344 -2296 3378
rect -2260 3344 -2226 3378
rect -2190 3344 -2156 3378
rect -2120 3344 -2086 3378
rect -2050 3344 -2016 3378
rect -1980 3344 -1946 3378
rect -1910 3344 -1876 3378
rect -1840 3344 -1806 3378
rect -1770 3344 -1736 3378
rect -1700 3344 -1666 3378
rect -1630 3344 -1596 3378
rect -1560 3344 -1526 3378
rect -1490 3344 -1456 3378
rect -1421 3344 -1387 3378
rect -1352 3344 -1318 3378
rect -1283 3344 -1249 3378
rect -1214 3344 -1180 3378
rect -1145 3344 -1111 3378
rect -1076 3344 -1042 3378
rect -1007 3344 -973 3378
rect -938 3344 -904 3378
rect -869 3344 -835 3378
rect -800 3344 -766 3378
rect -731 3344 -697 3378
rect -662 3344 -628 3378
rect -593 3344 -559 3378
rect -524 3344 -490 3378
rect -455 3344 -421 3378
rect -386 3344 -352 3378
rect -317 3344 -283 3378
rect -248 3344 -214 3378
rect -2750 3274 -2716 3308
rect -2680 3274 -2646 3308
rect -2610 3274 -2576 3308
rect -2540 3274 -2506 3308
rect -2470 3274 -2436 3308
rect -2400 3274 -2366 3308
rect -2330 3274 -2296 3308
rect -2260 3274 -2226 3308
rect -2190 3274 -2156 3308
rect -2120 3274 -2086 3308
rect -2050 3274 -2016 3308
rect -1980 3274 -1946 3308
rect -1910 3274 -1876 3308
rect -1840 3274 -1806 3308
rect -1770 3274 -1736 3308
rect -1700 3274 -1666 3308
rect -1630 3274 -1596 3308
rect -1560 3274 -1526 3308
rect -1490 3274 -1456 3308
rect -1421 3274 -1387 3308
rect -1352 3274 -1318 3308
rect -1283 3274 -1249 3308
rect -1214 3274 -1180 3308
rect -1145 3274 -1111 3308
rect -1076 3274 -1042 3308
rect -1007 3274 -973 3308
rect -938 3274 -904 3308
rect -869 3274 -835 3308
rect -800 3274 -766 3308
rect -731 3274 -697 3308
rect -662 3274 -628 3308
rect -593 3274 -559 3308
rect -524 3274 -490 3308
rect -455 3274 -421 3308
rect -386 3274 -352 3308
rect -317 3274 -283 3308
rect -248 3274 -214 3308
rect -2750 3204 -2716 3238
rect -2680 3204 -2646 3238
rect -2610 3204 -2576 3238
rect -2540 3204 -2506 3238
rect -2470 3204 -2436 3238
rect -2400 3204 -2366 3238
rect -2330 3204 -2296 3238
rect -2260 3204 -2226 3238
rect -2190 3204 -2156 3238
rect -2120 3204 -2086 3238
rect -2050 3204 -2016 3238
rect -1980 3204 -1946 3238
rect -1910 3204 -1876 3238
rect -1840 3204 -1806 3238
rect -1770 3204 -1736 3238
rect -1700 3204 -1666 3238
rect -1630 3204 -1596 3238
rect -1560 3204 -1526 3238
rect -1490 3204 -1456 3238
rect -1421 3204 -1387 3238
rect -1352 3204 -1318 3238
rect -1283 3204 -1249 3238
rect -1214 3204 -1180 3238
rect -1145 3204 -1111 3238
rect -1076 3204 -1042 3238
rect -1007 3204 -973 3238
rect -938 3204 -904 3238
rect -869 3204 -835 3238
rect -800 3204 -766 3238
rect -731 3204 -697 3238
rect -662 3204 -628 3238
rect -593 3204 -559 3238
rect -524 3204 -490 3238
rect -455 3204 -421 3238
rect -386 3204 -352 3238
rect -317 3204 -283 3238
rect -248 3204 -214 3238
rect -2750 3134 -2716 3168
rect -2680 3134 -2646 3168
rect -2610 3134 -2576 3168
rect -2540 3134 -2506 3168
rect -2470 3134 -2436 3168
rect -2400 3134 -2366 3168
rect -2330 3134 -2296 3168
rect -2260 3134 -2226 3168
rect -2190 3134 -2156 3168
rect -2120 3134 -2086 3168
rect -2050 3134 -2016 3168
rect -1980 3134 -1946 3168
rect -1910 3134 -1876 3168
rect -1840 3134 -1806 3168
rect -1770 3134 -1736 3168
rect -1700 3134 -1666 3168
rect -1630 3134 -1596 3168
rect -1560 3134 -1526 3168
rect -1490 3134 -1456 3168
rect -1421 3134 -1387 3168
rect -1352 3134 -1318 3168
rect -1283 3134 -1249 3168
rect -1214 3134 -1180 3168
rect -1145 3134 -1111 3168
rect -1076 3134 -1042 3168
rect -1007 3134 -973 3168
rect -938 3134 -904 3168
rect -869 3134 -835 3168
rect -800 3134 -766 3168
rect -731 3134 -697 3168
rect -662 3134 -628 3168
rect -593 3134 -559 3168
rect -524 3134 -490 3168
rect -455 3134 -421 3168
rect -386 3134 -352 3168
rect -317 3134 -283 3168
rect -248 3134 -214 3168
rect -161 3106 -127 3140
rect -89 3106 -55 3140
rect -17 3106 17 3140
rect 55 3106 89 3140
rect 127 3106 161 3140
rect 199 3106 233 3140
rect 271 3106 305 3140
rect -2750 3064 -2716 3098
rect -2680 3064 -2646 3098
rect -2610 3064 -2576 3098
rect -2540 3064 -2506 3098
rect -2470 3064 -2436 3098
rect -2400 3064 -2366 3098
rect -2330 3064 -2296 3098
rect -2260 3064 -2226 3098
rect -2190 3064 -2156 3098
rect -2120 3064 -2086 3098
rect -2050 3064 -2016 3098
rect -1980 3064 -1946 3098
rect -1910 3064 -1876 3098
rect -1840 3064 -1806 3098
rect -1770 3064 -1736 3098
rect -1700 3064 -1666 3098
rect -1630 3064 -1596 3098
rect -1560 3064 -1526 3098
rect -1490 3064 -1456 3098
rect -1421 3064 -1387 3098
rect -1352 3064 -1318 3098
rect -1283 3064 -1249 3098
rect -1214 3064 -1180 3098
rect -1145 3064 -1111 3098
rect -1076 3064 -1042 3098
rect -1007 3064 -973 3098
rect -938 3064 -904 3098
rect -869 3064 -835 3098
rect -800 3064 -766 3098
rect -731 3064 -697 3098
rect -662 3064 -628 3098
rect -593 3064 -559 3098
rect -524 3064 -490 3098
rect -455 3064 -421 3098
rect -386 3064 -352 3098
rect -317 3064 -283 3098
rect -248 3064 -214 3098
rect -161 3037 -127 3071
rect -89 3037 -55 3071
rect -17 3037 17 3071
rect 55 3037 89 3071
rect 127 3037 161 3071
rect 199 3037 233 3071
rect 271 3037 305 3071
rect -2750 2994 -2716 3028
rect -2680 2994 -2646 3028
rect -2610 2994 -2576 3028
rect -2540 2994 -2506 3028
rect -2470 2994 -2436 3028
rect -2400 2994 -2366 3028
rect -2330 2994 -2296 3028
rect -2260 2994 -2226 3028
rect -2190 2994 -2156 3028
rect -2120 2994 -2086 3028
rect -2050 2994 -2016 3028
rect -1980 2994 -1946 3028
rect -1910 2994 -1876 3028
rect -1840 2994 -1806 3028
rect -1770 2994 -1736 3028
rect -1700 2994 -1666 3028
rect -1630 2994 -1596 3028
rect -1560 2994 -1526 3028
rect -1490 2994 -1456 3028
rect -1421 2994 -1387 3028
rect -1352 2994 -1318 3028
rect -1283 2994 -1249 3028
rect -1214 2994 -1180 3028
rect -1145 2994 -1111 3028
rect -1076 2994 -1042 3028
rect -1007 2994 -973 3028
rect -938 2994 -904 3028
rect -869 2994 -835 3028
rect -800 2994 -766 3028
rect -731 2994 -697 3028
rect -662 2994 -628 3028
rect -593 2994 -559 3028
rect -524 2994 -490 3028
rect -455 2994 -421 3028
rect -386 2994 -352 3028
rect -317 2994 -283 3028
rect -248 2994 -214 3028
rect -161 2968 -127 3002
rect -89 2968 -55 3002
rect -17 2968 17 3002
rect 55 2968 89 3002
rect 127 2968 161 3002
rect 199 2968 233 3002
rect 271 2968 305 3002
rect -2750 2924 -2716 2958
rect -2680 2924 -2646 2958
rect -2610 2924 -2576 2958
rect -2540 2924 -2506 2958
rect -2470 2924 -2436 2958
rect -2400 2924 -2366 2958
rect -2330 2924 -2296 2958
rect -2260 2924 -2226 2958
rect -2190 2924 -2156 2958
rect -2120 2924 -2086 2958
rect -2050 2924 -2016 2958
rect -1980 2924 -1946 2958
rect -1910 2924 -1876 2958
rect -1840 2924 -1806 2958
rect -1770 2924 -1736 2958
rect -1700 2924 -1666 2958
rect -1630 2924 -1596 2958
rect -1560 2924 -1526 2958
rect -1490 2924 -1456 2958
rect -1421 2924 -1387 2958
rect -1352 2924 -1318 2958
rect -1283 2924 -1249 2958
rect -1214 2924 -1180 2958
rect -1145 2924 -1111 2958
rect -1076 2924 -1042 2958
rect -1007 2924 -973 2958
rect -938 2924 -904 2958
rect -869 2924 -835 2958
rect -800 2924 -766 2958
rect -731 2924 -697 2958
rect -662 2924 -628 2958
rect -593 2924 -559 2958
rect -524 2924 -490 2958
rect -455 2924 -421 2958
rect -386 2924 -352 2958
rect -317 2924 -283 2958
rect -248 2924 -214 2958
rect -161 2899 -127 2933
rect -89 2899 -55 2933
rect -17 2899 17 2933
rect 55 2899 89 2933
rect 127 2899 161 2933
rect 199 2899 233 2933
rect 271 2899 305 2933
rect -2750 2854 -2716 2888
rect -2680 2854 -2646 2888
rect -2610 2854 -2576 2888
rect -2540 2854 -2506 2888
rect -2470 2854 -2436 2888
rect -2400 2854 -2366 2888
rect -2330 2854 -2296 2888
rect -2260 2854 -2226 2888
rect -2190 2854 -2156 2888
rect -2120 2854 -2086 2888
rect -2050 2854 -2016 2888
rect -1980 2854 -1946 2888
rect -1910 2854 -1876 2888
rect -1840 2854 -1806 2888
rect -1770 2854 -1736 2888
rect -1700 2854 -1666 2888
rect -1630 2854 -1596 2888
rect -1560 2854 -1526 2888
rect -1490 2854 -1456 2888
rect -1421 2854 -1387 2888
rect -1352 2854 -1318 2888
rect -1283 2854 -1249 2888
rect -1214 2854 -1180 2888
rect -1145 2854 -1111 2888
rect -1076 2854 -1042 2888
rect -1007 2854 -973 2888
rect -938 2854 -904 2888
rect -869 2854 -835 2888
rect -800 2854 -766 2888
rect -731 2854 -697 2888
rect -662 2854 -628 2888
rect -593 2854 -559 2888
rect -524 2854 -490 2888
rect -455 2854 -421 2888
rect -386 2854 -352 2888
rect -317 2854 -283 2888
rect -248 2854 -214 2888
rect -161 2829 -127 2863
rect -89 2829 -55 2863
rect -17 2829 17 2863
rect 55 2829 89 2863
rect 127 2829 161 2863
rect 199 2829 233 2863
rect 271 2829 305 2863
rect -2750 2784 -2716 2818
rect -2680 2784 -2646 2818
rect -2610 2784 -2576 2818
rect -2540 2784 -2506 2818
rect -2470 2784 -2436 2818
rect -2400 2784 -2366 2818
rect -2330 2784 -2296 2818
rect -2260 2784 -2226 2818
rect -2190 2784 -2156 2818
rect -2120 2784 -2086 2818
rect -2050 2784 -2016 2818
rect -1980 2784 -1946 2818
rect -1910 2784 -1876 2818
rect -1840 2784 -1806 2818
rect -1770 2784 -1736 2818
rect -1700 2784 -1666 2818
rect -1630 2784 -1596 2818
rect -1560 2784 -1526 2818
rect -1490 2784 -1456 2818
rect -1421 2784 -1387 2818
rect -1352 2784 -1318 2818
rect -1283 2784 -1249 2818
rect -1214 2784 -1180 2818
rect -1145 2784 -1111 2818
rect -1076 2784 -1042 2818
rect -1007 2784 -973 2818
rect -938 2784 -904 2818
rect -869 2784 -835 2818
rect -800 2784 -766 2818
rect -731 2784 -697 2818
rect -662 2784 -628 2818
rect -593 2784 -559 2818
rect -524 2784 -490 2818
rect -455 2784 -421 2818
rect -386 2784 -352 2818
rect -317 2784 -283 2818
rect -248 2784 -214 2818
rect -161 2759 -127 2793
rect -89 2759 -55 2793
rect -17 2759 17 2793
rect 55 2759 89 2793
rect 127 2759 161 2793
rect 199 2759 233 2793
rect 271 2759 305 2793
rect -2750 2714 -2716 2748
rect -2680 2714 -2646 2748
rect -2610 2714 -2576 2748
rect -2540 2714 -2506 2748
rect -2470 2714 -2436 2748
rect -2400 2714 -2366 2748
rect -2330 2714 -2296 2748
rect -2260 2714 -2226 2748
rect -2190 2714 -2156 2748
rect -2120 2714 -2086 2748
rect -2050 2714 -2016 2748
rect -1980 2714 -1946 2748
rect -1910 2714 -1876 2748
rect -1840 2714 -1806 2748
rect -1770 2714 -1736 2748
rect -1700 2714 -1666 2748
rect -1630 2714 -1596 2748
rect -1560 2714 -1526 2748
rect -1490 2714 -1456 2748
rect -1421 2714 -1387 2748
rect -1352 2714 -1318 2748
rect -1283 2714 -1249 2748
rect -1214 2714 -1180 2748
rect -1145 2714 -1111 2748
rect -1076 2714 -1042 2748
rect -1007 2714 -973 2748
rect -938 2714 -904 2748
rect -869 2714 -835 2748
rect -800 2714 -766 2748
rect -731 2714 -697 2748
rect -662 2714 -628 2748
rect -593 2714 -559 2748
rect -524 2714 -490 2748
rect -455 2714 -421 2748
rect -386 2714 -352 2748
rect -317 2714 -283 2748
rect -248 2714 -214 2748
rect -161 2689 -127 2723
rect -89 2689 -55 2723
rect -17 2689 17 2723
rect 55 2689 89 2723
rect 127 2689 161 2723
rect 199 2689 233 2723
rect 271 2689 305 2723
rect -2750 2644 -2716 2678
rect -2680 2644 -2646 2678
rect -2610 2644 -2576 2678
rect -2540 2644 -2506 2678
rect -2470 2644 -2436 2678
rect -2400 2644 -2366 2678
rect -2330 2644 -2296 2678
rect -2260 2644 -2226 2678
rect -2190 2644 -2156 2678
rect -2120 2644 -2086 2678
rect -2050 2644 -2016 2678
rect -1980 2644 -1946 2678
rect -1910 2644 -1876 2678
rect -1840 2644 -1806 2678
rect -1770 2644 -1736 2678
rect -1700 2644 -1666 2678
rect -1630 2644 -1596 2678
rect -1560 2644 -1526 2678
rect -1490 2644 -1456 2678
rect -1421 2644 -1387 2678
rect -1352 2644 -1318 2678
rect -1283 2644 -1249 2678
rect -1214 2644 -1180 2678
rect -1145 2644 -1111 2678
rect -1076 2644 -1042 2678
rect -1007 2644 -973 2678
rect -938 2644 -904 2678
rect -869 2644 -835 2678
rect -800 2644 -766 2678
rect -731 2644 -697 2678
rect -662 2644 -628 2678
rect -593 2644 -559 2678
rect -524 2644 -490 2678
rect -455 2644 -421 2678
rect -386 2644 -352 2678
rect -317 2644 -283 2678
rect -248 2644 -214 2678
rect -161 2619 -127 2653
rect -89 2619 -55 2653
rect -17 2619 17 2653
rect 55 2619 89 2653
rect 127 2619 161 2653
rect 199 2619 233 2653
rect 271 2619 305 2653
rect -2750 2574 -2716 2608
rect -2680 2574 -2646 2608
rect -2610 2574 -2576 2608
rect -2540 2574 -2506 2608
rect -2470 2574 -2436 2608
rect -2400 2574 -2366 2608
rect -2330 2574 -2296 2608
rect -2260 2574 -2226 2608
rect -2190 2574 -2156 2608
rect -2120 2574 -2086 2608
rect -2050 2574 -2016 2608
rect -1980 2574 -1946 2608
rect -1910 2574 -1876 2608
rect -1840 2574 -1806 2608
rect -1770 2574 -1736 2608
rect -1700 2574 -1666 2608
rect -1630 2574 -1596 2608
rect -1560 2574 -1526 2608
rect -1490 2574 -1456 2608
rect -1421 2574 -1387 2608
rect -1352 2574 -1318 2608
rect -1283 2574 -1249 2608
rect -1214 2574 -1180 2608
rect -1145 2574 -1111 2608
rect -1076 2574 -1042 2608
rect -1007 2574 -973 2608
rect -938 2574 -904 2608
rect -869 2574 -835 2608
rect -800 2574 -766 2608
rect -731 2574 -697 2608
rect -662 2574 -628 2608
rect -593 2574 -559 2608
rect -524 2574 -490 2608
rect -455 2574 -421 2608
rect -386 2574 -352 2608
rect -317 2574 -283 2608
rect -248 2574 -214 2608
rect -161 2549 -127 2583
rect -89 2549 -55 2583
rect -17 2549 17 2583
rect 55 2549 89 2583
rect 127 2549 161 2583
rect 199 2549 233 2583
rect 271 2549 305 2583
rect -2750 2504 -2716 2538
rect -2680 2504 -2646 2538
rect -2610 2504 -2576 2538
rect -2540 2504 -2506 2538
rect -2470 2504 -2436 2538
rect -2400 2504 -2366 2538
rect -2330 2504 -2296 2538
rect -2260 2504 -2226 2538
rect -2190 2504 -2156 2538
rect -2120 2504 -2086 2538
rect -2050 2504 -2016 2538
rect -1980 2504 -1946 2538
rect -1910 2504 -1876 2538
rect -1840 2504 -1806 2538
rect -1770 2504 -1736 2538
rect -1700 2504 -1666 2538
rect -1630 2504 -1596 2538
rect -1560 2504 -1526 2538
rect -1490 2504 -1456 2538
rect -1421 2504 -1387 2538
rect -1352 2504 -1318 2538
rect -1283 2504 -1249 2538
rect -1214 2504 -1180 2538
rect -1145 2504 -1111 2538
rect -1076 2504 -1042 2538
rect -1007 2504 -973 2538
rect -938 2504 -904 2538
rect -869 2504 -835 2538
rect -800 2504 -766 2538
rect -731 2504 -697 2538
rect -662 2504 -628 2538
rect -593 2504 -559 2538
rect -524 2504 -490 2538
rect -455 2504 -421 2538
rect -386 2504 -352 2538
rect -317 2504 -283 2538
rect -248 2504 -214 2538
rect -161 2479 -127 2513
rect -89 2479 -55 2513
rect -17 2479 17 2513
rect 55 2479 89 2513
rect 127 2479 161 2513
rect 199 2479 233 2513
rect 271 2479 305 2513
rect -2750 2434 -2716 2468
rect -2680 2434 -2646 2468
rect -2610 2434 -2576 2468
rect -2540 2434 -2506 2468
rect -2470 2434 -2436 2468
rect -2400 2434 -2366 2468
rect -2330 2434 -2296 2468
rect -2260 2434 -2226 2468
rect -2190 2434 -2156 2468
rect -2120 2434 -2086 2468
rect -2050 2434 -2016 2468
rect -1980 2434 -1946 2468
rect -1910 2434 -1876 2468
rect -1840 2434 -1806 2468
rect -1770 2434 -1736 2468
rect -1700 2434 -1666 2468
rect -1630 2434 -1596 2468
rect -1560 2434 -1526 2468
rect -1490 2434 -1456 2468
rect -1421 2434 -1387 2468
rect -1352 2434 -1318 2468
rect -1283 2434 -1249 2468
rect -1214 2434 -1180 2468
rect -1145 2434 -1111 2468
rect -1076 2434 -1042 2468
rect -1007 2434 -973 2468
rect -938 2434 -904 2468
rect -869 2434 -835 2468
rect -800 2434 -766 2468
rect -731 2434 -697 2468
rect -662 2434 -628 2468
rect -593 2434 -559 2468
rect -524 2434 -490 2468
rect -455 2434 -421 2468
rect -386 2434 -352 2468
rect -317 2434 -283 2468
rect -248 2434 -214 2468
rect -161 2409 -127 2443
rect -89 2409 -55 2443
rect -17 2409 17 2443
rect 55 2409 89 2443
rect 127 2409 161 2443
rect 199 2409 233 2443
rect 271 2409 305 2443
rect -2750 2364 -2716 2398
rect -2680 2364 -2646 2398
rect -2610 2364 -2576 2398
rect -2540 2364 -2506 2398
rect -2470 2364 -2436 2398
rect -2400 2364 -2366 2398
rect -2330 2364 -2296 2398
rect -2260 2364 -2226 2398
rect -2190 2364 -2156 2398
rect -2120 2364 -2086 2398
rect -2050 2364 -2016 2398
rect -1980 2364 -1946 2398
rect -1910 2364 -1876 2398
rect -1840 2364 -1806 2398
rect -1770 2364 -1736 2398
rect -1700 2364 -1666 2398
rect -1630 2364 -1596 2398
rect -1560 2364 -1526 2398
rect -1490 2364 -1456 2398
rect -1421 2364 -1387 2398
rect -1352 2364 -1318 2398
rect -1283 2364 -1249 2398
rect -1214 2364 -1180 2398
rect -1145 2364 -1111 2398
rect -1076 2364 -1042 2398
rect -1007 2364 -973 2398
rect -938 2364 -904 2398
rect -869 2364 -835 2398
rect -800 2364 -766 2398
rect -731 2364 -697 2398
rect -662 2364 -628 2398
rect -593 2364 -559 2398
rect -524 2364 -490 2398
rect -455 2364 -421 2398
rect -386 2364 -352 2398
rect -317 2364 -283 2398
rect -248 2364 -214 2398
rect -161 2339 -127 2373
rect -89 2339 -55 2373
rect -17 2339 17 2373
rect 55 2339 89 2373
rect 127 2339 161 2373
rect 199 2339 233 2373
rect 271 2339 305 2373
rect -2750 2294 -2716 2328
rect -2680 2294 -2646 2328
rect -2610 2294 -2576 2328
rect -2540 2294 -2506 2328
rect -2470 2294 -2436 2328
rect -2400 2294 -2366 2328
rect -2330 2294 -2296 2328
rect -2260 2294 -2226 2328
rect -2190 2294 -2156 2328
rect -2120 2294 -2086 2328
rect -2050 2294 -2016 2328
rect -1980 2294 -1946 2328
rect -1910 2294 -1876 2328
rect -1840 2294 -1806 2328
rect -1770 2294 -1736 2328
rect -1700 2294 -1666 2328
rect -1630 2294 -1596 2328
rect -1560 2294 -1526 2328
rect -1490 2294 -1456 2328
rect -1421 2294 -1387 2328
rect -1352 2294 -1318 2328
rect -1283 2294 -1249 2328
rect -1214 2294 -1180 2328
rect -1145 2294 -1111 2328
rect -1076 2294 -1042 2328
rect -1007 2294 -973 2328
rect -938 2294 -904 2328
rect -869 2294 -835 2328
rect -800 2294 -766 2328
rect -731 2294 -697 2328
rect -662 2294 -628 2328
rect -593 2294 -559 2328
rect -524 2294 -490 2328
rect -455 2294 -421 2328
rect -386 2294 -352 2328
rect -317 2294 -283 2328
rect -248 2294 -214 2328
rect 2304 4494 2338 4528
rect 2374 4494 2408 4528
rect 2444 4494 2478 4528
rect 2514 4494 2548 4528
rect 2584 4494 2618 4528
rect 2654 4494 2688 4528
rect 2724 4494 2758 4528
rect 2794 4494 2828 4528
rect 2864 4494 2898 4528
rect 2934 4494 2968 4528
rect 3004 4494 3038 4528
rect 3074 4494 3108 4528
rect 3144 4494 3178 4528
rect 3214 4494 3248 4528
rect 3284 4494 3318 4528
rect 3354 4494 3388 4528
rect 3424 4494 3458 4528
rect 3494 4494 3528 4528
rect 3563 4494 3597 4528
rect 3632 4494 3666 4528
rect 3701 4494 3735 4528
rect 3770 4494 3804 4528
rect 3839 4494 3873 4528
rect 3908 4494 3942 4528
rect 3977 4494 4011 4528
rect 4046 4494 4080 4528
rect 4115 4494 4149 4528
rect 4184 4494 4218 4528
rect 4253 4494 4287 4528
rect 4322 4494 4356 4528
rect 4391 4494 4425 4528
rect 2304 4426 2338 4460
rect 2374 4426 2408 4460
rect 2444 4426 2478 4460
rect 2514 4426 2548 4460
rect 2584 4426 2618 4460
rect 2654 4426 2688 4460
rect 2724 4426 2758 4460
rect 2794 4426 2828 4460
rect 2864 4426 2898 4460
rect 2934 4426 2968 4460
rect 3004 4426 3038 4460
rect 3074 4426 3108 4460
rect 3144 4426 3178 4460
rect 3214 4426 3248 4460
rect 3284 4426 3318 4460
rect 3354 4426 3388 4460
rect 3424 4426 3458 4460
rect 3494 4426 3528 4460
rect 3563 4426 3597 4460
rect 3632 4426 3666 4460
rect 3701 4426 3735 4460
rect 3770 4426 3804 4460
rect 3839 4426 3873 4460
rect 3908 4426 3942 4460
rect 3977 4426 4011 4460
rect 4046 4426 4080 4460
rect 4115 4426 4149 4460
rect 4184 4426 4218 4460
rect 4253 4426 4287 4460
rect 4322 4426 4356 4460
rect 4391 4426 4425 4460
rect 2304 4358 2338 4392
rect 2374 4358 2408 4392
rect 2444 4358 2478 4392
rect 2514 4358 2548 4392
rect 2584 4358 2618 4392
rect 2654 4358 2688 4392
rect 2724 4358 2758 4392
rect 2794 4358 2828 4392
rect 2864 4358 2898 4392
rect 2934 4358 2968 4392
rect 3004 4358 3038 4392
rect 3074 4358 3108 4392
rect 3144 4358 3178 4392
rect 3214 4358 3248 4392
rect 3284 4358 3318 4392
rect 3354 4358 3388 4392
rect 3424 4358 3458 4392
rect 3494 4358 3528 4392
rect 3563 4358 3597 4392
rect 3632 4358 3666 4392
rect 3701 4358 3735 4392
rect 3770 4358 3804 4392
rect 3839 4358 3873 4392
rect 3908 4358 3942 4392
rect 3977 4358 4011 4392
rect 4046 4358 4080 4392
rect 4115 4358 4149 4392
rect 4184 4358 4218 4392
rect 4253 4358 4287 4392
rect 4322 4358 4356 4392
rect 4391 4358 4425 4392
rect 2304 4290 2338 4324
rect 2374 4290 2408 4324
rect 2444 4290 2478 4324
rect 2514 4290 2548 4324
rect 2584 4290 2618 4324
rect 2654 4290 2688 4324
rect 2724 4290 2758 4324
rect 2794 4290 2828 4324
rect 2864 4290 2898 4324
rect 2934 4290 2968 4324
rect 3004 4290 3038 4324
rect 3074 4290 3108 4324
rect 3144 4290 3178 4324
rect 3214 4290 3248 4324
rect 3284 4290 3318 4324
rect 3354 4290 3388 4324
rect 3424 4290 3458 4324
rect 3494 4290 3528 4324
rect 3563 4290 3597 4324
rect 3632 4290 3666 4324
rect 3701 4290 3735 4324
rect 3770 4290 3804 4324
rect 3839 4290 3873 4324
rect 3908 4290 3942 4324
rect 3977 4290 4011 4324
rect 4046 4290 4080 4324
rect 4115 4290 4149 4324
rect 4184 4290 4218 4324
rect 4253 4290 4287 4324
rect 4322 4290 4356 4324
rect 4391 4290 4425 4324
rect 2304 4222 2338 4256
rect 2374 4222 2408 4256
rect 2444 4222 2478 4256
rect 2514 4222 2548 4256
rect 2584 4222 2618 4256
rect 2654 4222 2688 4256
rect 2724 4222 2758 4256
rect 2794 4222 2828 4256
rect 2864 4222 2898 4256
rect 2934 4222 2968 4256
rect 3004 4222 3038 4256
rect 3074 4222 3108 4256
rect 3144 4222 3178 4256
rect 3214 4222 3248 4256
rect 3284 4222 3318 4256
rect 3354 4222 3388 4256
rect 3424 4222 3458 4256
rect 3494 4222 3528 4256
rect 3563 4222 3597 4256
rect 3632 4222 3666 4256
rect 3701 4222 3735 4256
rect 3770 4222 3804 4256
rect 3839 4222 3873 4256
rect 3908 4222 3942 4256
rect 3977 4222 4011 4256
rect 4046 4222 4080 4256
rect 4115 4222 4149 4256
rect 4184 4222 4218 4256
rect 4253 4222 4287 4256
rect 4322 4222 4356 4256
rect 4391 4222 4425 4256
rect 2304 4154 2338 4188
rect 2374 4154 2408 4188
rect 2444 4154 2478 4188
rect 2514 4154 2548 4188
rect 2584 4154 2618 4188
rect 2654 4154 2688 4188
rect 2724 4154 2758 4188
rect 2794 4154 2828 4188
rect 2864 4154 2898 4188
rect 2934 4154 2968 4188
rect 3004 4154 3038 4188
rect 3074 4154 3108 4188
rect 3144 4154 3178 4188
rect 3214 4154 3248 4188
rect 3284 4154 3318 4188
rect 3354 4154 3388 4188
rect 3424 4154 3458 4188
rect 3494 4154 3528 4188
rect 3563 4154 3597 4188
rect 3632 4154 3666 4188
rect 3701 4154 3735 4188
rect 3770 4154 3804 4188
rect 3839 4154 3873 4188
rect 3908 4154 3942 4188
rect 3977 4154 4011 4188
rect 4046 4154 4080 4188
rect 4115 4154 4149 4188
rect 4184 4154 4218 4188
rect 4253 4154 4287 4188
rect 4322 4154 4356 4188
rect 4391 4154 4425 4188
rect 2304 4086 2338 4120
rect 2374 4086 2408 4120
rect 2444 4086 2478 4120
rect 2514 4086 2548 4120
rect 2584 4086 2618 4120
rect 2654 4086 2688 4120
rect 2724 4086 2758 4120
rect 2794 4086 2828 4120
rect 2864 4086 2898 4120
rect 2934 4086 2968 4120
rect 3004 4086 3038 4120
rect 3074 4086 3108 4120
rect 3144 4086 3178 4120
rect 3214 4086 3248 4120
rect 3284 4086 3318 4120
rect 3354 4086 3388 4120
rect 3424 4086 3458 4120
rect 3494 4086 3528 4120
rect 3563 4086 3597 4120
rect 3632 4086 3666 4120
rect 3701 4086 3735 4120
rect 3770 4086 3804 4120
rect 3839 4086 3873 4120
rect 3908 4086 3942 4120
rect 3977 4086 4011 4120
rect 4046 4086 4080 4120
rect 4115 4086 4149 4120
rect 4184 4086 4218 4120
rect 4253 4086 4287 4120
rect 4322 4086 4356 4120
rect 4391 4086 4425 4120
rect 2304 4018 2338 4052
rect 2374 4018 2408 4052
rect 2444 4018 2478 4052
rect 2514 4018 2548 4052
rect 2584 4018 2618 4052
rect 2654 4018 2688 4052
rect 2724 4018 2758 4052
rect 2794 4018 2828 4052
rect 2864 4018 2898 4052
rect 2934 4018 2968 4052
rect 3004 4018 3038 4052
rect 3074 4018 3108 4052
rect 3144 4018 3178 4052
rect 3214 4018 3248 4052
rect 3284 4018 3318 4052
rect 3354 4018 3388 4052
rect 3424 4018 3458 4052
rect 3494 4018 3528 4052
rect 3563 4018 3597 4052
rect 3632 4018 3666 4052
rect 3701 4018 3735 4052
rect 3770 4018 3804 4052
rect 3839 4018 3873 4052
rect 3908 4018 3942 4052
rect 3977 4018 4011 4052
rect 4046 4018 4080 4052
rect 4115 4018 4149 4052
rect 4184 4018 4218 4052
rect 4253 4018 4287 4052
rect 4322 4018 4356 4052
rect 4391 4018 4425 4052
rect 2304 3950 2338 3984
rect 2374 3950 2408 3984
rect 2444 3950 2478 3984
rect 2514 3950 2548 3984
rect 2584 3950 2618 3984
rect 2654 3950 2688 3984
rect 2724 3950 2758 3984
rect 2794 3950 2828 3984
rect 2864 3950 2898 3984
rect 2934 3950 2968 3984
rect 3004 3950 3038 3984
rect 3074 3950 3108 3984
rect 3144 3950 3178 3984
rect 3214 3950 3248 3984
rect 3284 3950 3318 3984
rect 3354 3950 3388 3984
rect 3424 3950 3458 3984
rect 3494 3950 3528 3984
rect 3563 3950 3597 3984
rect 3632 3950 3666 3984
rect 3701 3950 3735 3984
rect 3770 3950 3804 3984
rect 3839 3950 3873 3984
rect 3908 3950 3942 3984
rect 3977 3950 4011 3984
rect 4046 3950 4080 3984
rect 4115 3950 4149 3984
rect 4184 3950 4218 3984
rect 4253 3950 4287 3984
rect 4322 3950 4356 3984
rect 4391 3950 4425 3984
rect 2304 3882 2338 3916
rect 2374 3882 2408 3916
rect 2444 3882 2478 3916
rect 2514 3882 2548 3916
rect 2584 3882 2618 3916
rect 2654 3882 2688 3916
rect 2724 3882 2758 3916
rect 2794 3882 2828 3916
rect 2864 3882 2898 3916
rect 2934 3882 2968 3916
rect 3004 3882 3038 3916
rect 3074 3882 3108 3916
rect 3144 3882 3178 3916
rect 3214 3882 3248 3916
rect 3284 3882 3318 3916
rect 3354 3882 3388 3916
rect 3424 3882 3458 3916
rect 3494 3882 3528 3916
rect 3563 3882 3597 3916
rect 3632 3882 3666 3916
rect 3701 3882 3735 3916
rect 3770 3882 3804 3916
rect 3839 3882 3873 3916
rect 3908 3882 3942 3916
rect 3977 3882 4011 3916
rect 4046 3882 4080 3916
rect 4115 3882 4149 3916
rect 4184 3882 4218 3916
rect 4253 3882 4287 3916
rect 4322 3882 4356 3916
rect 4391 3882 4425 3916
rect 2304 3814 2338 3848
rect 2374 3814 2408 3848
rect 2444 3814 2478 3848
rect 2514 3814 2548 3848
rect 2584 3814 2618 3848
rect 2654 3814 2688 3848
rect 2724 3814 2758 3848
rect 2794 3814 2828 3848
rect 2864 3814 2898 3848
rect 2934 3814 2968 3848
rect 3004 3814 3038 3848
rect 3074 3814 3108 3848
rect 3144 3814 3178 3848
rect 3214 3814 3248 3848
rect 3284 3814 3318 3848
rect 3354 3814 3388 3848
rect 3424 3814 3458 3848
rect 3494 3814 3528 3848
rect 3563 3814 3597 3848
rect 3632 3814 3666 3848
rect 3701 3814 3735 3848
rect 3770 3814 3804 3848
rect 3839 3814 3873 3848
rect 3908 3814 3942 3848
rect 3977 3814 4011 3848
rect 4046 3814 4080 3848
rect 4115 3814 4149 3848
rect 4184 3814 4218 3848
rect 4253 3814 4287 3848
rect 4322 3814 4356 3848
rect 4391 3814 4425 3848
rect 2304 3746 2338 3780
rect 2374 3746 2408 3780
rect 2444 3746 2478 3780
rect 2514 3746 2548 3780
rect 2584 3746 2618 3780
rect 2654 3746 2688 3780
rect 2724 3746 2758 3780
rect 2794 3746 2828 3780
rect 2864 3746 2898 3780
rect 2934 3746 2968 3780
rect 3004 3746 3038 3780
rect 3074 3746 3108 3780
rect 3144 3746 3178 3780
rect 3214 3746 3248 3780
rect 3284 3746 3318 3780
rect 3354 3746 3388 3780
rect 3424 3746 3458 3780
rect 3494 3746 3528 3780
rect 3563 3746 3597 3780
rect 3632 3746 3666 3780
rect 3701 3746 3735 3780
rect 3770 3746 3804 3780
rect 3839 3746 3873 3780
rect 3908 3746 3942 3780
rect 3977 3746 4011 3780
rect 4046 3746 4080 3780
rect 4115 3746 4149 3780
rect 4184 3746 4218 3780
rect 4253 3746 4287 3780
rect 4322 3746 4356 3780
rect 4391 3746 4425 3780
rect 2304 3678 2338 3712
rect 2374 3678 2408 3712
rect 2444 3678 2478 3712
rect 2514 3678 2548 3712
rect 2584 3678 2618 3712
rect 2654 3678 2688 3712
rect 2724 3678 2758 3712
rect 2794 3678 2828 3712
rect 2864 3678 2898 3712
rect 2934 3678 2968 3712
rect 3004 3678 3038 3712
rect 3074 3678 3108 3712
rect 3144 3678 3178 3712
rect 3214 3678 3248 3712
rect 3284 3678 3318 3712
rect 3354 3678 3388 3712
rect 3424 3678 3458 3712
rect 3494 3678 3528 3712
rect 3563 3678 3597 3712
rect 3632 3678 3666 3712
rect 3701 3678 3735 3712
rect 3770 3678 3804 3712
rect 3839 3678 3873 3712
rect 3908 3678 3942 3712
rect 3977 3678 4011 3712
rect 4046 3678 4080 3712
rect 4115 3678 4149 3712
rect 4184 3678 4218 3712
rect 4253 3678 4287 3712
rect 4322 3678 4356 3712
rect 4391 3678 4425 3712
rect 2304 3610 2338 3644
rect 2374 3610 2408 3644
rect 2444 3610 2478 3644
rect 2514 3610 2548 3644
rect 2584 3610 2618 3644
rect 2654 3610 2688 3644
rect 2724 3610 2758 3644
rect 2794 3610 2828 3644
rect 2864 3610 2898 3644
rect 2934 3610 2968 3644
rect 3004 3610 3038 3644
rect 3074 3610 3108 3644
rect 3144 3610 3178 3644
rect 3214 3610 3248 3644
rect 3284 3610 3318 3644
rect 3354 3610 3388 3644
rect 3424 3610 3458 3644
rect 3494 3610 3528 3644
rect 3563 3610 3597 3644
rect 3632 3610 3666 3644
rect 3701 3610 3735 3644
rect 3770 3610 3804 3644
rect 3839 3610 3873 3644
rect 3908 3610 3942 3644
rect 3977 3610 4011 3644
rect 4046 3610 4080 3644
rect 4115 3610 4149 3644
rect 4184 3610 4218 3644
rect 4253 3610 4287 3644
rect 4322 3610 4356 3644
rect 4391 3610 4425 3644
rect 2304 3542 2338 3576
rect 2374 3542 2408 3576
rect 2444 3542 2478 3576
rect 2514 3542 2548 3576
rect 2584 3542 2618 3576
rect 2654 3542 2688 3576
rect 2724 3542 2758 3576
rect 2794 3542 2828 3576
rect 2864 3542 2898 3576
rect 2934 3542 2968 3576
rect 3004 3542 3038 3576
rect 3074 3542 3108 3576
rect 3144 3542 3178 3576
rect 3214 3542 3248 3576
rect 3284 3542 3318 3576
rect 3354 3542 3388 3576
rect 3424 3542 3458 3576
rect 3494 3542 3528 3576
rect 3563 3542 3597 3576
rect 3632 3542 3666 3576
rect 3701 3542 3735 3576
rect 3770 3542 3804 3576
rect 3839 3542 3873 3576
rect 3908 3542 3942 3576
rect 3977 3542 4011 3576
rect 4046 3542 4080 3576
rect 4115 3542 4149 3576
rect 4184 3542 4218 3576
rect 4253 3542 4287 3576
rect 4322 3542 4356 3576
rect 4391 3542 4425 3576
rect 11159 4470 11193 4504
rect 11231 4470 11265 4504
rect 11303 4470 11337 4504
rect 11375 4470 11409 4504
rect 11447 4470 11481 4504
rect 11519 4470 11553 4504
rect 11591 4470 11625 4504
rect 11663 4470 11697 4504
rect 11159 4400 11193 4434
rect 11231 4400 11265 4434
rect 11303 4400 11337 4434
rect 11375 4400 11409 4434
rect 11447 4400 11481 4434
rect 11519 4400 11553 4434
rect 11591 4400 11625 4434
rect 11663 4400 11697 4434
rect 11159 4330 11193 4364
rect 11231 4330 11265 4364
rect 11303 4330 11337 4364
rect 11375 4330 11409 4364
rect 11447 4330 11481 4364
rect 11519 4330 11553 4364
rect 11591 4330 11625 4364
rect 11663 4330 11697 4364
rect 11159 4260 11193 4294
rect 11231 4260 11265 4294
rect 11303 4260 11337 4294
rect 11375 4260 11409 4294
rect 11447 4260 11481 4294
rect 11519 4260 11553 4294
rect 11591 4260 11625 4294
rect 11663 4260 11697 4294
rect 11159 4189 11193 4223
rect 11231 4189 11265 4223
rect 11303 4189 11337 4223
rect 11375 4189 11409 4223
rect 11447 4189 11481 4223
rect 11519 4189 11553 4223
rect 11591 4189 11625 4223
rect 11663 4189 11697 4223
rect 11159 4118 11193 4152
rect 11231 4118 11265 4152
rect 11303 4118 11337 4152
rect 11375 4118 11409 4152
rect 11447 4118 11481 4152
rect 11519 4118 11553 4152
rect 11591 4118 11625 4152
rect 11663 4118 11697 4152
rect 11159 4047 11193 4081
rect 11231 4047 11265 4081
rect 11303 4047 11337 4081
rect 11375 4047 11409 4081
rect 11447 4047 11481 4081
rect 11519 4047 11553 4081
rect 11591 4047 11625 4081
rect 11663 4047 11697 4081
rect 11159 3976 11193 4010
rect 11231 3976 11265 4010
rect 11303 3976 11337 4010
rect 11375 3976 11409 4010
rect 11447 3976 11481 4010
rect 11519 3976 11553 4010
rect 11591 3976 11625 4010
rect 11663 3976 11697 4010
rect 11159 3905 11193 3939
rect 11231 3905 11265 3939
rect 11303 3905 11337 3939
rect 11375 3905 11409 3939
rect 11447 3905 11481 3939
rect 11519 3905 11553 3939
rect 11591 3905 11625 3939
rect 11663 3905 11697 3939
rect 11159 3834 11193 3868
rect 11231 3834 11265 3868
rect 11303 3834 11337 3868
rect 11375 3834 11409 3868
rect 11447 3834 11481 3868
rect 11519 3834 11553 3868
rect 11591 3834 11625 3868
rect 11663 3834 11697 3868
rect 11159 3763 11193 3797
rect 11231 3763 11265 3797
rect 11303 3763 11337 3797
rect 11375 3763 11409 3797
rect 11447 3763 11481 3797
rect 11519 3763 11553 3797
rect 11591 3763 11625 3797
rect 11663 3763 11697 3797
rect 11159 3692 11193 3726
rect 11231 3692 11265 3726
rect 11303 3692 11337 3726
rect 11375 3692 11409 3726
rect 11447 3692 11481 3726
rect 11519 3692 11553 3726
rect 11591 3692 11625 3726
rect 11663 3692 11697 3726
rect 11159 3621 11193 3655
rect 11231 3621 11265 3655
rect 11303 3621 11337 3655
rect 11375 3621 11409 3655
rect 11447 3621 11481 3655
rect 11519 3621 11553 3655
rect 11591 3621 11625 3655
rect 11663 3621 11697 3655
rect 2304 3474 2338 3508
rect 2374 3474 2408 3508
rect 2444 3474 2478 3508
rect 2514 3474 2548 3508
rect 2584 3474 2618 3508
rect 2654 3474 2688 3508
rect 2724 3474 2758 3508
rect 2794 3474 2828 3508
rect 2864 3474 2898 3508
rect 2934 3474 2968 3508
rect 3004 3474 3038 3508
rect 3074 3474 3108 3508
rect 3144 3474 3178 3508
rect 3214 3474 3248 3508
rect 3284 3474 3318 3508
rect 3354 3474 3388 3508
rect 3424 3474 3458 3508
rect 3494 3474 3528 3508
rect 3563 3474 3597 3508
rect 3632 3474 3666 3508
rect 3701 3474 3735 3508
rect 3770 3474 3804 3508
rect 3839 3474 3873 3508
rect 3908 3474 3942 3508
rect 3977 3474 4011 3508
rect 4046 3474 4080 3508
rect 4115 3474 4149 3508
rect 4184 3474 4218 3508
rect 4253 3474 4287 3508
rect 4322 3474 4356 3508
rect 4391 3474 4425 3508
rect 2304 3406 2338 3440
rect 2374 3406 2408 3440
rect 2444 3406 2478 3440
rect 2514 3406 2548 3440
rect 2584 3406 2618 3440
rect 2654 3406 2688 3440
rect 2724 3406 2758 3440
rect 2794 3406 2828 3440
rect 2864 3406 2898 3440
rect 2934 3406 2968 3440
rect 3004 3406 3038 3440
rect 3074 3406 3108 3440
rect 3144 3406 3178 3440
rect 3214 3406 3248 3440
rect 3284 3406 3318 3440
rect 3354 3406 3388 3440
rect 3424 3406 3458 3440
rect 3494 3406 3528 3440
rect 3563 3406 3597 3440
rect 3632 3406 3666 3440
rect 3701 3406 3735 3440
rect 3770 3406 3804 3440
rect 3839 3406 3873 3440
rect 3908 3406 3942 3440
rect 3977 3406 4011 3440
rect 4046 3406 4080 3440
rect 4115 3406 4149 3440
rect 4184 3406 4218 3440
rect 4253 3406 4287 3440
rect 4322 3406 4356 3440
rect 4391 3406 4425 3440
rect 4529 3537 4563 3571
rect 4598 3537 4632 3571
rect 4667 3537 4701 3571
rect 4736 3537 4770 3571
rect 4805 3537 4839 3571
rect 4874 3537 4908 3571
rect 4943 3537 4977 3571
rect 5012 3537 5046 3571
rect 5081 3537 5115 3571
rect 5150 3537 5184 3571
rect 5219 3537 5253 3571
rect 5288 3537 5322 3571
rect 5357 3537 5391 3571
rect 5426 3537 5460 3571
rect 5495 3537 5529 3571
rect 5564 3537 5598 3571
rect 5633 3537 5667 3571
rect 5702 3537 5736 3571
rect 5771 3537 5805 3571
rect 5840 3537 5874 3571
rect 5909 3537 5943 3571
rect 5978 3537 6012 3571
rect 6047 3537 6081 3571
rect 6116 3537 6150 3571
rect 6185 3537 6219 3571
rect 6254 3537 6288 3571
rect 6323 3537 6357 3571
rect 6392 3537 6426 3571
rect 6461 3537 6495 3571
rect 6530 3537 6564 3571
rect 6599 3537 6633 3571
rect 6668 3537 6702 3571
rect 6737 3537 6771 3571
rect 6806 3537 6840 3571
rect 6875 3537 6909 3571
rect 6944 3537 6978 3571
rect 7013 3537 7047 3571
rect 7082 3537 7116 3571
rect 7151 3537 7185 3571
rect 4529 3469 4563 3503
rect 4598 3469 4632 3503
rect 4667 3469 4701 3503
rect 4736 3469 4770 3503
rect 4805 3469 4839 3503
rect 4874 3469 4908 3503
rect 4943 3469 4977 3503
rect 5012 3469 5046 3503
rect 5081 3469 5115 3503
rect 5150 3469 5184 3503
rect 5219 3469 5253 3503
rect 5288 3469 5322 3503
rect 5357 3469 5391 3503
rect 5426 3469 5460 3503
rect 5495 3469 5529 3503
rect 5564 3469 5598 3503
rect 5633 3469 5667 3503
rect 5702 3469 5736 3503
rect 5771 3469 5805 3503
rect 5840 3469 5874 3503
rect 5909 3469 5943 3503
rect 5978 3469 6012 3503
rect 6047 3469 6081 3503
rect 6116 3469 6150 3503
rect 6185 3469 6219 3503
rect 6254 3469 6288 3503
rect 6323 3469 6357 3503
rect 6392 3469 6426 3503
rect 6461 3469 6495 3503
rect 6530 3469 6564 3503
rect 6599 3469 6633 3503
rect 6668 3469 6702 3503
rect 6737 3469 6771 3503
rect 6806 3469 6840 3503
rect 6875 3469 6909 3503
rect 6944 3469 6978 3503
rect 7013 3469 7047 3503
rect 7082 3469 7116 3503
rect 7151 3469 7185 3503
rect 4529 3401 4563 3435
rect 4598 3401 4632 3435
rect 4667 3401 4701 3435
rect 4736 3401 4770 3435
rect 4805 3401 4839 3435
rect 4874 3401 4908 3435
rect 4943 3401 4977 3435
rect 5012 3401 5046 3435
rect 5081 3401 5115 3435
rect 5150 3401 5184 3435
rect 5219 3401 5253 3435
rect 5288 3401 5322 3435
rect 5357 3401 5391 3435
rect 5426 3401 5460 3435
rect 5495 3401 5529 3435
rect 5564 3401 5598 3435
rect 5633 3401 5667 3435
rect 5702 3401 5736 3435
rect 5771 3401 5805 3435
rect 5840 3401 5874 3435
rect 5909 3401 5943 3435
rect 5978 3401 6012 3435
rect 6047 3401 6081 3435
rect 6116 3401 6150 3435
rect 6185 3401 6219 3435
rect 6254 3401 6288 3435
rect 6323 3401 6357 3435
rect 6392 3401 6426 3435
rect 6461 3401 6495 3435
rect 6530 3401 6564 3435
rect 6599 3401 6633 3435
rect 6668 3401 6702 3435
rect 6737 3401 6771 3435
rect 6806 3401 6840 3435
rect 6875 3401 6909 3435
rect 6944 3401 6978 3435
rect 7013 3401 7047 3435
rect 7082 3401 7116 3435
rect 7151 3401 7185 3435
rect 7220 3401 11674 3571
rect 2304 3338 2338 3372
rect 2374 3338 2408 3372
rect 2444 3338 2478 3372
rect 2514 3338 2548 3372
rect 2584 3338 2618 3372
rect 2654 3338 2688 3372
rect 2724 3338 2758 3372
rect 2794 3338 2828 3372
rect 2864 3338 2898 3372
rect 2934 3338 2968 3372
rect 3004 3338 3038 3372
rect 3074 3338 3108 3372
rect 3144 3338 3178 3372
rect 3214 3338 3248 3372
rect 3284 3338 3318 3372
rect 3354 3338 3388 3372
rect 3424 3338 3458 3372
rect 3494 3338 3528 3372
rect 3563 3338 3597 3372
rect 3632 3338 3666 3372
rect 3701 3338 3735 3372
rect 3770 3338 3804 3372
rect 3839 3338 3873 3372
rect 3908 3338 3942 3372
rect 3977 3338 4011 3372
rect 4046 3338 4080 3372
rect 4115 3338 4149 3372
rect 4184 3338 4218 3372
rect 4253 3338 4287 3372
rect 4322 3338 4356 3372
rect 4391 3338 4425 3372
rect 2304 3270 2338 3304
rect 2374 3270 2408 3304
rect 2444 3270 2478 3304
rect 2514 3270 2548 3304
rect 2584 3270 2618 3304
rect 2654 3270 2688 3304
rect 2724 3270 2758 3304
rect 2794 3270 2828 3304
rect 2864 3270 2898 3304
rect 2934 3270 2968 3304
rect 3004 3270 3038 3304
rect 3074 3270 3108 3304
rect 3144 3270 3178 3304
rect 3214 3270 3248 3304
rect 3284 3270 3318 3304
rect 3354 3270 3388 3304
rect 3424 3270 3458 3304
rect 3494 3270 3528 3304
rect 3563 3270 3597 3304
rect 3632 3270 3666 3304
rect 3701 3270 3735 3304
rect 3770 3270 3804 3304
rect 3839 3270 3873 3304
rect 3908 3270 3942 3304
rect 3977 3270 4011 3304
rect 4046 3270 4080 3304
rect 4115 3270 4149 3304
rect 4184 3270 4218 3304
rect 4253 3270 4287 3304
rect 4322 3270 4356 3304
rect 4391 3270 4425 3304
rect 2304 3202 2338 3236
rect 2374 3202 2408 3236
rect 2444 3202 2478 3236
rect 2514 3202 2548 3236
rect 2584 3202 2618 3236
rect 2654 3202 2688 3236
rect 2724 3202 2758 3236
rect 2794 3202 2828 3236
rect 2864 3202 2898 3236
rect 2934 3202 2968 3236
rect 3004 3202 3038 3236
rect 3074 3202 3108 3236
rect 3144 3202 3178 3236
rect 3214 3202 3248 3236
rect 3284 3202 3318 3236
rect 3354 3202 3388 3236
rect 3424 3202 3458 3236
rect 3494 3202 3528 3236
rect 3563 3202 3597 3236
rect 3632 3202 3666 3236
rect 3701 3202 3735 3236
rect 3770 3202 3804 3236
rect 3839 3202 3873 3236
rect 3908 3202 3942 3236
rect 3977 3202 4011 3236
rect 4046 3202 4080 3236
rect 4115 3202 4149 3236
rect 4184 3202 4218 3236
rect 4253 3202 4287 3236
rect 4322 3202 4356 3236
rect 4391 3202 4425 3236
rect 2304 3134 2338 3168
rect 2374 3134 2408 3168
rect 2444 3134 2478 3168
rect 2514 3134 2548 3168
rect 2584 3134 2618 3168
rect 2654 3134 2688 3168
rect 2724 3134 2758 3168
rect 2794 3134 2828 3168
rect 2864 3134 2898 3168
rect 2934 3134 2968 3168
rect 3004 3134 3038 3168
rect 3074 3134 3108 3168
rect 3144 3134 3178 3168
rect 3214 3134 3248 3168
rect 3284 3134 3318 3168
rect 3354 3134 3388 3168
rect 3424 3134 3458 3168
rect 3494 3134 3528 3168
rect 3563 3134 3597 3168
rect 3632 3134 3666 3168
rect 3701 3134 3735 3168
rect 3770 3134 3804 3168
rect 3839 3134 3873 3168
rect 3908 3134 3942 3168
rect 3977 3134 4011 3168
rect 4046 3134 4080 3168
rect 4115 3134 4149 3168
rect 4184 3134 4218 3168
rect 4253 3134 4287 3168
rect 4322 3134 4356 3168
rect 4391 3134 4425 3168
rect 2304 3066 2338 3100
rect 2374 3066 2408 3100
rect 2444 3066 2478 3100
rect 2514 3066 2548 3100
rect 2584 3066 2618 3100
rect 2654 3066 2688 3100
rect 2724 3066 2758 3100
rect 2794 3066 2828 3100
rect 2864 3066 2898 3100
rect 2934 3066 2968 3100
rect 3004 3066 3038 3100
rect 3074 3066 3108 3100
rect 3144 3066 3178 3100
rect 3214 3066 3248 3100
rect 3284 3066 3318 3100
rect 3354 3066 3388 3100
rect 3424 3066 3458 3100
rect 3494 3066 3528 3100
rect 3563 3066 3597 3100
rect 3632 3066 3666 3100
rect 3701 3066 3735 3100
rect 3770 3066 3804 3100
rect 3839 3066 3873 3100
rect 3908 3066 3942 3100
rect 3977 3066 4011 3100
rect 4046 3066 4080 3100
rect 4115 3066 4149 3100
rect 4184 3066 4218 3100
rect 4253 3066 4287 3100
rect 4322 3066 4356 3100
rect 4391 3066 4425 3100
rect 2304 2998 2338 3032
rect 2374 2998 2408 3032
rect 2444 2998 2478 3032
rect 2514 2998 2548 3032
rect 2584 2998 2618 3032
rect 2654 2998 2688 3032
rect 2724 2998 2758 3032
rect 2794 2998 2828 3032
rect 2864 2998 2898 3032
rect 2934 2998 2968 3032
rect 3004 2998 3038 3032
rect 3074 2998 3108 3032
rect 3144 2998 3178 3032
rect 3214 2998 3248 3032
rect 3284 2998 3318 3032
rect 3354 2998 3388 3032
rect 3424 2998 3458 3032
rect 3494 2998 3528 3032
rect 3563 2998 3597 3032
rect 3632 2998 3666 3032
rect 3701 2998 3735 3032
rect 3770 2998 3804 3032
rect 3839 2998 3873 3032
rect 3908 2998 3942 3032
rect 3977 2998 4011 3032
rect 4046 2998 4080 3032
rect 4115 2998 4149 3032
rect 4184 2998 4218 3032
rect 4253 2998 4287 3032
rect 4322 2998 4356 3032
rect 4391 2998 4425 3032
rect 2304 2930 2338 2964
rect 2374 2930 2408 2964
rect 2444 2930 2478 2964
rect 2514 2930 2548 2964
rect 2584 2930 2618 2964
rect 2654 2930 2688 2964
rect 2724 2930 2758 2964
rect 2794 2930 2828 2964
rect 2864 2930 2898 2964
rect 2934 2930 2968 2964
rect 3004 2930 3038 2964
rect 3074 2930 3108 2964
rect 3144 2930 3178 2964
rect 3214 2930 3248 2964
rect 3284 2930 3318 2964
rect 3354 2930 3388 2964
rect 3424 2930 3458 2964
rect 3494 2930 3528 2964
rect 3563 2930 3597 2964
rect 3632 2930 3666 2964
rect 3701 2930 3735 2964
rect 3770 2930 3804 2964
rect 3839 2930 3873 2964
rect 3908 2930 3942 2964
rect 3977 2930 4011 2964
rect 4046 2930 4080 2964
rect 4115 2930 4149 2964
rect 4184 2930 4218 2964
rect 4253 2930 4287 2964
rect 4322 2930 4356 2964
rect 4391 2930 4425 2964
rect 2304 2862 2338 2896
rect 2374 2862 2408 2896
rect 2444 2862 2478 2896
rect 2514 2862 2548 2896
rect 2584 2862 2618 2896
rect 2654 2862 2688 2896
rect 2724 2862 2758 2896
rect 2794 2862 2828 2896
rect 2864 2862 2898 2896
rect 2934 2862 2968 2896
rect 3004 2862 3038 2896
rect 3074 2862 3108 2896
rect 3144 2862 3178 2896
rect 3214 2862 3248 2896
rect 3284 2862 3318 2896
rect 3354 2862 3388 2896
rect 3424 2862 3458 2896
rect 3494 2862 3528 2896
rect 3563 2862 3597 2896
rect 3632 2862 3666 2896
rect 3701 2862 3735 2896
rect 3770 2862 3804 2896
rect 3839 2862 3873 2896
rect 3908 2862 3942 2896
rect 3977 2862 4011 2896
rect 4046 2862 4080 2896
rect 4115 2862 4149 2896
rect 4184 2862 4218 2896
rect 4253 2862 4287 2896
rect 4322 2862 4356 2896
rect 4391 2862 4425 2896
rect 2304 2794 2338 2828
rect 2374 2794 2408 2828
rect 2444 2794 2478 2828
rect 2514 2794 2548 2828
rect 2584 2794 2618 2828
rect 2654 2794 2688 2828
rect 2724 2794 2758 2828
rect 2794 2794 2828 2828
rect 2864 2794 2898 2828
rect 2934 2794 2968 2828
rect 3004 2794 3038 2828
rect 3074 2794 3108 2828
rect 3144 2794 3178 2828
rect 3214 2794 3248 2828
rect 3284 2794 3318 2828
rect 3354 2794 3388 2828
rect 3424 2794 3458 2828
rect 3494 2794 3528 2828
rect 3563 2794 3597 2828
rect 3632 2794 3666 2828
rect 3701 2794 3735 2828
rect 3770 2794 3804 2828
rect 3839 2794 3873 2828
rect 3908 2794 3942 2828
rect 3977 2794 4011 2828
rect 4046 2794 4080 2828
rect 4115 2794 4149 2828
rect 4184 2794 4218 2828
rect 4253 2794 4287 2828
rect 4322 2794 4356 2828
rect 4391 2794 4425 2828
rect 2304 2726 2338 2760
rect 2374 2726 2408 2760
rect 2444 2726 2478 2760
rect 2514 2726 2548 2760
rect 2584 2726 2618 2760
rect 2654 2726 2688 2760
rect 2724 2726 2758 2760
rect 2794 2726 2828 2760
rect 2864 2726 2898 2760
rect 2934 2726 2968 2760
rect 3004 2726 3038 2760
rect 3074 2726 3108 2760
rect 3144 2726 3178 2760
rect 3214 2726 3248 2760
rect 3284 2726 3318 2760
rect 3354 2726 3388 2760
rect 3424 2726 3458 2760
rect 3494 2726 3528 2760
rect 3563 2726 3597 2760
rect 3632 2726 3666 2760
rect 3701 2726 3735 2760
rect 3770 2726 3804 2760
rect 3839 2726 3873 2760
rect 3908 2726 3942 2760
rect 3977 2726 4011 2760
rect 4046 2726 4080 2760
rect 4115 2726 4149 2760
rect 4184 2726 4218 2760
rect 4253 2726 4287 2760
rect 4322 2726 4356 2760
rect 4391 2726 4425 2760
rect 2304 2658 2338 2692
rect 2374 2658 2408 2692
rect 2444 2658 2478 2692
rect 2514 2658 2548 2692
rect 2584 2658 2618 2692
rect 2654 2658 2688 2692
rect 2724 2658 2758 2692
rect 2794 2658 2828 2692
rect 2864 2658 2898 2692
rect 2934 2658 2968 2692
rect 3004 2658 3038 2692
rect 3074 2658 3108 2692
rect 3144 2658 3178 2692
rect 3214 2658 3248 2692
rect 3284 2658 3318 2692
rect 3354 2658 3388 2692
rect 3424 2658 3458 2692
rect 3494 2658 3528 2692
rect 3563 2658 3597 2692
rect 3632 2658 3666 2692
rect 3701 2658 3735 2692
rect 3770 2658 3804 2692
rect 3839 2658 3873 2692
rect 3908 2658 3942 2692
rect 3977 2658 4011 2692
rect 4046 2658 4080 2692
rect 4115 2658 4149 2692
rect 4184 2658 4218 2692
rect 4253 2658 4287 2692
rect 4322 2658 4356 2692
rect 4391 2658 4425 2692
rect 2304 2590 2338 2624
rect 2374 2590 2408 2624
rect 2444 2590 2478 2624
rect 2514 2590 2548 2624
rect 2584 2590 2618 2624
rect 2654 2590 2688 2624
rect 2724 2590 2758 2624
rect 2794 2590 2828 2624
rect 2864 2590 2898 2624
rect 2934 2590 2968 2624
rect 3004 2590 3038 2624
rect 3074 2590 3108 2624
rect 3144 2590 3178 2624
rect 3214 2590 3248 2624
rect 3284 2590 3318 2624
rect 3354 2590 3388 2624
rect 3424 2590 3458 2624
rect 3494 2590 3528 2624
rect 3563 2590 3597 2624
rect 3632 2590 3666 2624
rect 3701 2590 3735 2624
rect 3770 2590 3804 2624
rect 3839 2590 3873 2624
rect 3908 2590 3942 2624
rect 3977 2590 4011 2624
rect 4046 2590 4080 2624
rect 4115 2590 4149 2624
rect 4184 2590 4218 2624
rect 4253 2590 4287 2624
rect 4322 2590 4356 2624
rect 4391 2590 4425 2624
rect 2304 2522 2338 2556
rect 2374 2522 2408 2556
rect 2444 2522 2478 2556
rect 2514 2522 2548 2556
rect 2584 2522 2618 2556
rect 2654 2522 2688 2556
rect 2724 2522 2758 2556
rect 2794 2522 2828 2556
rect 2864 2522 2898 2556
rect 2934 2522 2968 2556
rect 3004 2522 3038 2556
rect 3074 2522 3108 2556
rect 3144 2522 3178 2556
rect 3214 2522 3248 2556
rect 3284 2522 3318 2556
rect 3354 2522 3388 2556
rect 3424 2522 3458 2556
rect 3494 2522 3528 2556
rect 3563 2522 3597 2556
rect 3632 2522 3666 2556
rect 3701 2522 3735 2556
rect 3770 2522 3804 2556
rect 3839 2522 3873 2556
rect 3908 2522 3942 2556
rect 3977 2522 4011 2556
rect 4046 2522 4080 2556
rect 4115 2522 4149 2556
rect 4184 2522 4218 2556
rect 4253 2522 4287 2556
rect 4322 2522 4356 2556
rect 4391 2522 4425 2556
rect 2304 2454 2338 2488
rect 2374 2454 2408 2488
rect 2444 2454 2478 2488
rect 2514 2454 2548 2488
rect 2584 2454 2618 2488
rect 2654 2454 2688 2488
rect 2724 2454 2758 2488
rect 2794 2454 2828 2488
rect 2864 2454 2898 2488
rect 2934 2454 2968 2488
rect 3004 2454 3038 2488
rect 3074 2454 3108 2488
rect 3144 2454 3178 2488
rect 3214 2454 3248 2488
rect 3284 2454 3318 2488
rect 3354 2454 3388 2488
rect 3424 2454 3458 2488
rect 3494 2454 3528 2488
rect 3563 2454 3597 2488
rect 3632 2454 3666 2488
rect 3701 2454 3735 2488
rect 3770 2454 3804 2488
rect 3839 2454 3873 2488
rect 3908 2454 3942 2488
rect 3977 2454 4011 2488
rect 4046 2454 4080 2488
rect 4115 2454 4149 2488
rect 4184 2454 4218 2488
rect 4253 2454 4287 2488
rect 4322 2454 4356 2488
rect 4391 2454 4425 2488
rect 2304 2386 2338 2420
rect 2374 2386 2408 2420
rect 2444 2386 2478 2420
rect 2514 2386 2548 2420
rect 2584 2386 2618 2420
rect 2654 2386 2688 2420
rect 2724 2386 2758 2420
rect 2794 2386 2828 2420
rect 2864 2386 2898 2420
rect 2934 2386 2968 2420
rect 3004 2386 3038 2420
rect 3074 2386 3108 2420
rect 3144 2386 3178 2420
rect 3214 2386 3248 2420
rect 3284 2386 3318 2420
rect 3354 2386 3388 2420
rect 3424 2386 3458 2420
rect 3494 2386 3528 2420
rect 3563 2386 3597 2420
rect 3632 2386 3666 2420
rect 3701 2386 3735 2420
rect 3770 2386 3804 2420
rect 3839 2386 3873 2420
rect 3908 2386 3942 2420
rect 3977 2386 4011 2420
rect 4046 2386 4080 2420
rect 4115 2386 4149 2420
rect 4184 2386 4218 2420
rect 4253 2386 4287 2420
rect 4322 2386 4356 2420
rect 4391 2386 4425 2420
rect -161 2269 -127 2303
rect -89 2269 -55 2303
rect -17 2269 17 2303
rect 55 2269 89 2303
rect 127 2269 161 2303
rect 199 2269 233 2303
rect 271 2269 305 2303
rect 2304 2318 2338 2352
rect 2374 2318 2408 2352
rect 2444 2318 2478 2352
rect 2514 2318 2548 2352
rect 2584 2318 2618 2352
rect 2654 2318 2688 2352
rect 2724 2318 2758 2352
rect 2794 2318 2828 2352
rect 2864 2318 2898 2352
rect 2934 2318 2968 2352
rect 3004 2318 3038 2352
rect 3074 2318 3108 2352
rect 3144 2318 3178 2352
rect 3214 2318 3248 2352
rect 3284 2318 3318 2352
rect 3354 2318 3388 2352
rect 3424 2318 3458 2352
rect 3494 2318 3528 2352
rect 3563 2318 3597 2352
rect 3632 2318 3666 2352
rect 3701 2318 3735 2352
rect 3770 2318 3804 2352
rect 3839 2318 3873 2352
rect 3908 2318 3942 2352
rect 3977 2318 4011 2352
rect 4046 2318 4080 2352
rect 4115 2318 4149 2352
rect 4184 2318 4218 2352
rect 4253 2318 4287 2352
rect 4322 2318 4356 2352
rect 4391 2318 4425 2352
rect 2304 2250 2338 2284
rect 2374 2250 2408 2284
rect 2444 2250 2478 2284
rect 2514 2250 2548 2284
rect 2584 2250 2618 2284
rect 2654 2250 2688 2284
rect 2724 2250 2758 2284
rect 2794 2250 2828 2284
rect 2864 2250 2898 2284
rect 2934 2250 2968 2284
rect 3004 2250 3038 2284
rect 3074 2250 3108 2284
rect 3144 2250 3178 2284
rect 3214 2250 3248 2284
rect 3284 2250 3318 2284
rect 3354 2250 3388 2284
rect 3424 2250 3458 2284
rect 3494 2250 3528 2284
rect 3563 2250 3597 2284
rect 3632 2250 3666 2284
rect 3701 2250 3735 2284
rect 3770 2250 3804 2284
rect 3839 2250 3873 2284
rect 3908 2250 3942 2284
rect 3977 2250 4011 2284
rect 4046 2250 4080 2284
rect 4115 2250 4149 2284
rect 4184 2250 4218 2284
rect 4253 2250 4287 2284
rect 4322 2250 4356 2284
rect 4391 2250 4425 2284
rect -2726 2159 -2692 2193
rect -2656 2159 -2622 2193
rect -2586 2159 -2552 2193
rect -2517 2159 -2483 2193
rect -2448 2159 -2414 2193
rect -2379 2159 -2345 2193
rect -2310 2159 -2276 2193
rect -2241 2159 -2207 2193
rect -2172 2159 -2138 2193
rect -2103 2159 -2069 2193
rect -2034 2159 -2000 2193
rect -1965 2159 -1931 2193
rect -1896 2159 -1862 2193
rect -1827 2159 -1793 2193
rect -1758 2159 -1724 2193
rect -1689 2159 -1655 2193
rect -1620 2159 -1586 2193
rect -1551 2159 -1517 2193
rect -1482 2159 -1448 2193
rect -1413 2159 -1379 2193
rect -1344 2159 -1310 2193
rect -1275 2159 -1241 2193
rect -1206 2159 -1172 2193
rect -1137 2159 -1103 2193
rect -1068 2159 -1034 2193
rect -999 2159 -965 2193
rect -930 2159 -896 2193
rect -861 2159 -827 2193
rect -792 2159 -758 2193
rect -723 2159 -689 2193
rect -654 2159 -620 2193
rect -585 2159 -551 2193
rect -516 2159 -482 2193
rect -447 2159 -413 2193
rect -378 2159 -344 2193
rect -309 2159 -275 2193
rect -240 2159 -206 2193
rect -171 2159 -137 2193
rect -102 2159 -68 2193
rect -33 2159 1 2193
rect 36 2159 70 2193
rect 105 2159 139 2193
rect 174 2159 208 2193
rect 243 2159 277 2193
rect 2298 2159 2332 2193
rect 2368 2159 2402 2193
rect 2438 2159 2472 2193
rect 2508 2159 2542 2193
rect 2578 2159 2612 2193
rect 2648 2159 2682 2193
rect 2718 2159 2752 2193
rect 2788 2159 2822 2193
rect 2858 2159 2892 2193
rect 2928 2159 2962 2193
rect 2998 2159 3032 2193
rect 3068 2159 3102 2193
rect 3138 2159 3172 2193
rect 3208 2159 3242 2193
rect 3278 2159 3312 2193
rect 3348 2159 3382 2193
rect 3418 2159 3452 2193
rect 3488 2159 3522 2193
rect 3558 2159 3592 2193
rect 3628 2159 3662 2193
rect 3698 2159 3732 2193
rect 3768 2159 3802 2193
rect 3838 2159 3872 2193
rect 3908 2159 3942 2193
rect 3977 2159 4011 2193
rect 4046 2159 4080 2193
rect 4115 2159 4149 2193
rect 4184 2159 4218 2193
rect 4253 2159 4287 2193
rect 4322 2159 4356 2193
rect 4391 2159 4425 2193
rect -2726 2091 -2692 2125
rect -2656 2091 -2622 2125
rect -2586 2091 -2552 2125
rect -2517 2091 -2483 2125
rect -2448 2091 -2414 2125
rect -2379 2091 -2345 2125
rect -2310 2091 -2276 2125
rect -2241 2091 -2207 2125
rect -2172 2091 -2138 2125
rect -2103 2091 -2069 2125
rect -2034 2091 -2000 2125
rect -1965 2091 -1931 2125
rect -1896 2091 -1862 2125
rect -1827 2091 -1793 2125
rect -1758 2091 -1724 2125
rect -1689 2091 -1655 2125
rect -1620 2091 -1586 2125
rect -1551 2091 -1517 2125
rect -1482 2091 -1448 2125
rect -1413 2091 -1379 2125
rect -1344 2091 -1310 2125
rect -1275 2091 -1241 2125
rect -1206 2091 -1172 2125
rect -1137 2091 -1103 2125
rect -1068 2091 -1034 2125
rect -999 2091 -965 2125
rect -930 2091 -896 2125
rect -861 2091 -827 2125
rect -792 2091 -758 2125
rect -723 2091 -689 2125
rect -654 2091 -620 2125
rect -585 2091 -551 2125
rect -516 2091 -482 2125
rect -447 2091 -413 2125
rect -378 2091 -344 2125
rect -309 2091 -275 2125
rect -240 2091 -206 2125
rect -171 2091 -137 2125
rect -102 2091 -68 2125
rect -33 2091 1 2125
rect 36 2091 70 2125
rect 105 2091 139 2125
rect 174 2091 208 2125
rect 243 2091 277 2125
rect 2298 2091 2332 2125
rect 2368 2091 2402 2125
rect 2438 2091 2472 2125
rect 2508 2091 2542 2125
rect 2578 2091 2612 2125
rect 2648 2091 2682 2125
rect 2718 2091 2752 2125
rect 2788 2091 2822 2125
rect 2858 2091 2892 2125
rect 2928 2091 2962 2125
rect 2998 2091 3032 2125
rect 3068 2091 3102 2125
rect 3138 2091 3172 2125
rect 3208 2091 3242 2125
rect 3278 2091 3312 2125
rect 3348 2091 3382 2125
rect 3418 2091 3452 2125
rect 3488 2091 3522 2125
rect 3558 2091 3592 2125
rect 3628 2091 3662 2125
rect 3698 2091 3732 2125
rect 3768 2091 3802 2125
rect 3838 2091 3872 2125
rect 3908 2091 3942 2125
rect 3977 2091 4011 2125
rect 4046 2091 4080 2125
rect 4115 2091 4149 2125
rect 4184 2091 4218 2125
rect 4253 2091 4287 2125
rect 4322 2091 4356 2125
rect 4391 2091 4425 2125
rect -2726 2023 -2692 2057
rect -2656 2023 -2622 2057
rect -2586 2023 -2552 2057
rect -2517 2023 -2483 2057
rect -2448 2023 -2414 2057
rect -2379 2023 -2345 2057
rect -2310 2023 -2276 2057
rect -2241 2023 -2207 2057
rect -2172 2023 -2138 2057
rect -2103 2023 -2069 2057
rect -2034 2023 -2000 2057
rect -1965 2023 -1931 2057
rect -1896 2023 -1862 2057
rect -1827 2023 -1793 2057
rect -1758 2023 -1724 2057
rect -1689 2023 -1655 2057
rect -1620 2023 -1586 2057
rect -1551 2023 -1517 2057
rect -1482 2023 -1448 2057
rect -1413 2023 -1379 2057
rect -1344 2023 -1310 2057
rect -1275 2023 -1241 2057
rect -1206 2023 -1172 2057
rect -1137 2023 -1103 2057
rect -1068 2023 -1034 2057
rect -999 2023 -965 2057
rect -930 2023 -896 2057
rect -861 2023 -827 2057
rect -792 2023 -758 2057
rect -723 2023 -689 2057
rect -654 2023 -620 2057
rect -585 2023 -551 2057
rect -516 2023 -482 2057
rect -447 2023 -413 2057
rect -378 2023 -344 2057
rect -309 2023 -275 2057
rect -240 2023 -206 2057
rect -171 2023 -137 2057
rect -102 2023 -68 2057
rect -33 2023 1 2057
rect 36 2023 70 2057
rect 105 2023 139 2057
rect 174 2023 208 2057
rect 243 2023 277 2057
rect 2298 2023 2332 2057
rect 2368 2023 2402 2057
rect 2438 2023 2472 2057
rect 2508 2023 2542 2057
rect 2578 2023 2612 2057
rect 2648 2023 2682 2057
rect 2718 2023 2752 2057
rect 2788 2023 2822 2057
rect 2858 2023 2892 2057
rect 2928 2023 2962 2057
rect 2998 2023 3032 2057
rect 3068 2023 3102 2057
rect 3138 2023 3172 2057
rect 3208 2023 3242 2057
rect 3278 2023 3312 2057
rect 3348 2023 3382 2057
rect 3418 2023 3452 2057
rect 3488 2023 3522 2057
rect 3558 2023 3592 2057
rect 3628 2023 3662 2057
rect 3698 2023 3732 2057
rect 3768 2023 3802 2057
rect 3838 2023 3872 2057
rect 3908 2023 3942 2057
rect 3977 2023 4011 2057
rect 4046 2023 4080 2057
rect 4115 2023 4149 2057
rect 4184 2023 4218 2057
rect 4253 2023 4287 2057
rect 4322 2023 4356 2057
rect 4391 2023 4425 2057
rect 10267 1236 10301 1270
rect 10335 1236 10369 1270
rect 10403 1236 10437 1270
rect 10471 1236 10505 1270
rect 10539 1236 10573 1270
rect 10607 1236 10641 1270
rect 10675 1236 10709 1270
rect 10743 1236 10777 1270
rect 10811 1236 10845 1270
rect 10879 1236 10913 1270
rect 10947 1236 10981 1270
rect 11015 1236 11049 1270
rect 11083 1236 11117 1270
rect 11151 1236 11185 1270
rect 11219 1236 11253 1270
rect 11287 1236 11321 1270
rect 11355 1236 11389 1270
rect 11423 1236 11457 1270
rect 11491 1236 11525 1270
rect 11559 1236 11593 1270
rect 11627 1236 11661 1270
rect 11695 1236 11729 1270
rect 11763 1236 11797 1270
rect 11831 1236 11865 1270
rect 11899 1236 11933 1270
rect 11967 1236 12001 1270
rect 12035 1236 12069 1270
rect 12103 1236 12137 1270
rect 12171 1236 12205 1270
rect 12239 1236 12273 1270
rect 12307 1236 12341 1270
rect 12375 1236 12409 1270
rect 12443 1236 12477 1270
rect 12511 1236 12545 1270
rect 12579 1236 12613 1270
rect 12647 1236 12681 1270
rect 12715 1236 12749 1270
rect 12783 1236 12817 1270
rect 12851 1236 12885 1270
rect 12919 1236 12953 1270
rect 12987 1236 13021 1270
rect 13055 1236 13089 1270
rect 13123 1236 13157 1270
rect 13191 1236 13225 1270
rect 13259 1236 13293 1270
rect 13327 1236 13361 1270
rect 13395 1236 13429 1270
rect 13463 1236 13497 1270
rect 13531 1236 13565 1270
rect 13599 1236 13633 1270
rect 13667 1236 13701 1270
rect 13735 1236 13769 1270
rect 13803 1236 13837 1270
rect 13871 1236 13905 1270
rect 13939 1236 13973 1270
rect 14007 1236 14041 1270
rect 14076 1236 14110 1270
rect 14145 1236 14179 1270
rect 14214 1236 14248 1270
rect 14283 1236 14317 1270
rect 14352 1236 14386 1270
rect 14421 1236 14455 1270
rect 14490 1236 14524 1270
rect 14559 1236 14593 1270
rect 14628 1236 14662 1270
rect 14697 1236 14731 1270
rect 14766 1236 14800 1270
rect 14835 1236 14869 1270
rect 14904 1236 14938 1270
rect 14973 1236 15007 1270
rect 15042 1236 15076 1270
rect 15111 1236 15145 1270
rect 15180 1236 15214 1270
rect 15249 1236 15283 1270
rect 15318 1236 15352 1270
rect 15386 1167 15420 1201
rect 6270 1127 6304 1161
rect 6338 1127 6372 1161
rect 6406 1127 6440 1161
rect 6474 1127 6508 1161
rect 6542 1127 6576 1161
rect 6611 1127 6645 1161
rect 6680 1127 6714 1161
rect 6749 1127 6783 1161
rect 6818 1127 6852 1161
rect 6887 1127 6921 1161
rect 6956 1127 6990 1161
rect 7025 1127 7059 1161
rect 7094 1127 7128 1161
rect 7163 1127 7197 1161
rect 7232 1127 7266 1161
rect 7301 1127 7335 1161
rect 7370 1127 7404 1161
rect 7439 1127 7473 1161
rect 7508 1127 7542 1161
rect 7577 1127 7611 1161
rect 7646 1127 7680 1161
rect 7715 1127 7749 1161
rect 7784 1127 7818 1161
rect 7853 1127 7887 1161
rect 7922 1127 7956 1161
rect 7991 1127 8025 1161
rect 8060 1127 8094 1161
rect 8129 1127 8163 1161
rect 8198 1127 8232 1161
rect 8267 1127 8301 1161
rect 8336 1127 8370 1161
rect 8405 1127 8439 1161
rect 8474 1127 8508 1161
rect 8543 1127 8577 1161
rect 8612 1127 8646 1161
rect 8681 1127 8715 1161
rect 8750 1127 8784 1161
rect 8819 1127 8853 1161
rect 8888 1127 8922 1161
rect 8957 1127 8991 1161
rect 9026 1127 9060 1161
rect 9095 1127 9129 1161
rect 9164 1127 9198 1161
rect 9233 1127 9267 1161
rect 9302 1127 9336 1161
rect 9371 1127 9405 1161
rect 9440 1127 9474 1161
rect 9509 1127 9543 1161
rect 9578 1127 9612 1161
rect 9647 1127 9681 1161
rect 9716 1127 9750 1161
rect 9785 1127 9819 1161
rect 9854 1127 9888 1161
rect 9923 1127 9957 1161
rect 9992 1127 10026 1161
rect 10061 1127 10095 1161
rect 10130 1127 10164 1161
rect 10199 1127 10233 1161
rect 6202 1059 6236 1093
rect 10325 1090 10359 1124
rect 10393 1110 10427 1144
rect 10461 1110 10495 1144
rect 10529 1110 10563 1144
rect 10597 1110 10631 1144
rect 10665 1110 10699 1144
rect 10733 1110 10767 1144
rect 10801 1110 10835 1144
rect 10869 1110 10903 1144
rect 10937 1110 10971 1144
rect 11005 1110 11039 1144
rect 11073 1110 11107 1144
rect 11141 1110 11175 1144
rect 11209 1110 11243 1144
rect 11277 1110 11311 1144
rect 11345 1110 11379 1144
rect 11413 1110 11447 1144
rect 11481 1110 11515 1144
rect 11549 1110 11583 1144
rect 11617 1110 11651 1144
rect 11685 1110 11719 1144
rect 11753 1110 11787 1144
rect 11821 1110 11855 1144
rect 11889 1110 11923 1144
rect 11957 1110 11991 1144
rect 12025 1110 12059 1144
rect 12093 1110 12127 1144
rect 12161 1110 12195 1144
rect 12229 1110 12263 1144
rect 12297 1110 12331 1144
rect 12365 1110 12399 1144
rect 12433 1110 12467 1144
rect 12501 1110 12535 1144
rect 12569 1110 12603 1144
rect 12638 1110 12672 1144
rect 12707 1110 12741 1144
rect 12776 1110 12810 1144
rect 12845 1110 12879 1144
rect 12914 1110 12948 1144
rect 12983 1110 13017 1144
rect 13052 1110 13086 1144
rect 13121 1110 13155 1144
rect 13190 1110 13224 1144
rect 13259 1110 13293 1144
rect 13328 1110 13362 1144
rect 13397 1110 13431 1144
rect 13466 1110 13500 1144
rect 13535 1110 13569 1144
rect 13604 1110 13638 1144
rect 13673 1110 13707 1144
rect 13742 1110 13776 1144
rect 13811 1110 13845 1144
rect 13880 1110 13914 1144
rect 13949 1110 13983 1144
rect 14018 1110 14052 1144
rect 14087 1110 14121 1144
rect 14156 1110 14190 1144
rect 14225 1110 14259 1144
rect 14294 1110 14328 1144
rect 14363 1110 14397 1144
rect 14432 1110 14466 1144
rect 14501 1110 14535 1144
rect 14570 1110 14604 1144
rect 14639 1110 14673 1144
rect 14708 1110 14742 1144
rect 14777 1110 14811 1144
rect 14846 1110 14880 1144
rect 14915 1110 14949 1144
rect 14984 1110 15018 1144
rect 15053 1110 15087 1144
rect 15122 1110 15156 1144
rect 15191 1110 15225 1144
rect 15260 1110 15294 1144
rect 6202 984 6236 1018
rect 6328 1001 6362 1035
rect 6396 1001 6430 1035
rect 6464 1001 6498 1035
rect 6532 1001 6566 1035
rect 6600 1001 6634 1035
rect 6669 1001 6703 1035
rect 6738 1001 6772 1035
rect 6807 1001 6841 1035
rect 6876 1001 6910 1035
rect 6945 1001 6979 1035
rect 7014 1001 7048 1035
rect 7083 1001 7117 1035
rect 7152 1001 7186 1035
rect 7221 1001 7255 1035
rect 7290 1001 7324 1035
rect 7359 1001 7393 1035
rect 7428 1001 7462 1035
rect 7497 1001 7531 1035
rect 7566 1001 7600 1035
rect 7635 1001 7669 1035
rect 7704 1001 7738 1035
rect 7773 1001 7807 1035
rect 7842 1001 7876 1035
rect 7911 1001 7945 1035
rect 7980 1001 8014 1035
rect 8049 1001 8083 1035
rect 8118 1001 8152 1035
rect 8187 1001 8221 1035
rect 8256 1001 8290 1035
rect 8325 1001 8359 1035
rect 8394 1001 8428 1035
rect 8463 1001 8497 1035
rect 8532 1001 8566 1035
rect 8601 1001 8635 1035
rect 8670 1001 8704 1035
rect 8739 1001 8773 1035
rect 8808 1001 8842 1035
rect 8877 1001 8911 1035
rect 8946 1001 8980 1035
rect 9015 1001 9049 1035
rect 9084 1001 9118 1035
rect 9153 1001 9187 1035
rect 9222 1001 9256 1035
rect 9291 1001 9325 1035
rect 9360 1001 9394 1035
rect 9429 1001 9463 1035
rect 9498 1001 9532 1035
rect 9567 1001 9601 1035
rect 9636 1001 9670 1035
rect 9705 1001 9739 1035
rect 9774 1001 9808 1035
rect 9843 1001 9877 1035
rect 9912 1001 9946 1035
rect 9981 1001 10015 1035
rect 10050 1001 10084 1035
rect 10119 1001 10153 1035
rect 10188 1001 10222 1035
rect 10257 1001 10291 1035
rect 15386 1098 15420 1132
rect 15260 1040 15294 1074
rect 15386 1029 15420 1063
rect 15260 969 15294 1003
rect 15386 960 15420 994
rect 6202 909 6236 943
rect 6328 923 6362 957
rect 6202 834 6236 868
rect 6328 846 6362 880
rect 6202 759 6236 793
rect 6328 769 6362 803
rect 15260 898 15294 932
rect 15386 891 15420 925
rect 15260 827 15294 861
rect 15386 822 15420 856
rect 6202 684 6236 718
rect 6328 692 6362 726
rect 15260 756 15294 790
rect 15386 752 15420 786
rect 15260 685 15294 719
rect 15386 682 15420 716
rect 6202 609 6236 643
rect 6328 615 6362 649
rect 6202 535 6236 569
rect 6328 538 6362 572
rect 6202 461 6236 495
rect 6328 461 6362 495
rect 15260 614 15294 648
rect 15386 612 15420 646
rect 15260 543 15294 577
rect 15386 542 15420 576
rect 15260 472 15294 506
rect 15386 472 15420 506
<< poly >>
rect 12 4110 112 4126
rect 12 4076 45 4110
rect 79 4076 112 4110
rect 12 4058 112 4076
rect 12 3340 112 3358
rect 12 3306 45 3340
rect 79 3306 112 3340
rect 12 3290 112 3306
rect 6567 708 14748 725
rect 6567 674 6583 708
rect 6617 674 6652 708
rect 6686 674 6721 708
rect 6755 674 6790 708
rect 6824 674 6859 708
rect 6893 674 6928 708
rect 6962 674 6997 708
rect 7031 674 7066 708
rect 7100 674 7135 708
rect 7169 674 7204 708
rect 7238 674 7273 708
rect 7307 674 7342 708
rect 7376 674 7411 708
rect 7445 674 7480 708
rect 7514 674 7549 708
rect 7583 674 7618 708
rect 7652 674 7687 708
rect 7721 674 7756 708
rect 7790 674 7824 708
rect 7858 674 7892 708
rect 7926 674 7960 708
rect 7994 674 8028 708
rect 8062 674 8096 708
rect 8130 674 8164 708
rect 8198 674 8232 708
rect 8266 674 8300 708
rect 8334 674 8368 708
rect 8402 674 8436 708
rect 8470 674 8504 708
rect 8538 674 8572 708
rect 8606 674 8640 708
rect 8674 674 8708 708
rect 8742 674 8776 708
rect 8810 674 8844 708
rect 8878 674 8912 708
rect 8946 674 8980 708
rect 9014 674 9048 708
rect 9082 674 9116 708
rect 9150 674 9184 708
rect 9218 674 9252 708
rect 9286 674 9320 708
rect 9354 674 9388 708
rect 9422 674 9456 708
rect 9490 674 9524 708
rect 9558 674 9592 708
rect 9626 674 9660 708
rect 9694 674 9728 708
rect 9762 674 9796 708
rect 9830 674 9864 708
rect 9898 674 9932 708
rect 9966 674 10000 708
rect 10034 674 10068 708
rect 10102 674 10136 708
rect 10170 674 10204 708
rect 10238 674 10272 708
rect 10306 674 10340 708
rect 10374 674 10408 708
rect 10442 674 10476 708
rect 10510 674 10801 708
rect 10835 674 10870 708
rect 10904 674 10939 708
rect 10973 674 11008 708
rect 11042 674 11077 708
rect 11111 674 11146 708
rect 11180 674 11215 708
rect 11249 674 11284 708
rect 11318 674 11353 708
rect 11387 674 11422 708
rect 11456 674 11491 708
rect 11525 674 11560 708
rect 11594 674 11629 708
rect 11663 674 11698 708
rect 11732 674 11767 708
rect 11801 674 11836 708
rect 11870 674 11905 708
rect 11939 674 11974 708
rect 12008 674 12043 708
rect 12077 674 12112 708
rect 12146 674 12181 708
rect 12215 674 12250 708
rect 12284 674 12318 708
rect 12352 674 12386 708
rect 12420 674 12454 708
rect 12488 674 12522 708
rect 12556 674 12590 708
rect 12624 674 12658 708
rect 12692 674 12726 708
rect 12760 674 12794 708
rect 12828 674 12862 708
rect 12896 674 12930 708
rect 12964 674 12998 708
rect 13032 674 13066 708
rect 13100 674 13134 708
rect 13168 674 13202 708
rect 13236 674 13270 708
rect 13304 674 13338 708
rect 13372 674 13406 708
rect 13440 674 13474 708
rect 13508 674 13542 708
rect 13576 674 13610 708
rect 13644 674 13678 708
rect 13712 674 13746 708
rect 13780 674 13814 708
rect 13848 674 13882 708
rect 13916 674 13950 708
rect 13984 674 14018 708
rect 14052 674 14086 708
rect 14120 674 14154 708
rect 14188 674 14222 708
rect 14256 674 14290 708
rect 14324 674 14358 708
rect 14392 674 14426 708
rect 14460 674 14494 708
rect 14528 674 14562 708
rect 14596 674 14630 708
rect 14664 674 14698 708
rect 14732 674 14748 708
rect 6567 653 14748 674
<< polycont >>
rect 45 4076 79 4110
rect 45 3306 79 3340
rect 6583 674 6617 708
rect 6652 674 6686 708
rect 6721 674 6755 708
rect 6790 674 6824 708
rect 6859 674 6893 708
rect 6928 674 6962 708
rect 6997 674 7031 708
rect 7066 674 7100 708
rect 7135 674 7169 708
rect 7204 674 7238 708
rect 7273 674 7307 708
rect 7342 674 7376 708
rect 7411 674 7445 708
rect 7480 674 7514 708
rect 7549 674 7583 708
rect 7618 674 7652 708
rect 7687 674 7721 708
rect 7756 674 7790 708
rect 7824 674 7858 708
rect 7892 674 7926 708
rect 7960 674 7994 708
rect 8028 674 8062 708
rect 8096 674 8130 708
rect 8164 674 8198 708
rect 8232 674 8266 708
rect 8300 674 8334 708
rect 8368 674 8402 708
rect 8436 674 8470 708
rect 8504 674 8538 708
rect 8572 674 8606 708
rect 8640 674 8674 708
rect 8708 674 8742 708
rect 8776 674 8810 708
rect 8844 674 8878 708
rect 8912 674 8946 708
rect 8980 674 9014 708
rect 9048 674 9082 708
rect 9116 674 9150 708
rect 9184 674 9218 708
rect 9252 674 9286 708
rect 9320 674 9354 708
rect 9388 674 9422 708
rect 9456 674 9490 708
rect 9524 674 9558 708
rect 9592 674 9626 708
rect 9660 674 9694 708
rect 9728 674 9762 708
rect 9796 674 9830 708
rect 9864 674 9898 708
rect 9932 674 9966 708
rect 10000 674 10034 708
rect 10068 674 10102 708
rect 10136 674 10170 708
rect 10204 674 10238 708
rect 10272 674 10306 708
rect 10340 674 10374 708
rect 10408 674 10442 708
rect 10476 674 10510 708
rect 10801 674 10835 708
rect 10870 674 10904 708
rect 10939 674 10973 708
rect 11008 674 11042 708
rect 11077 674 11111 708
rect 11146 674 11180 708
rect 11215 674 11249 708
rect 11284 674 11318 708
rect 11353 674 11387 708
rect 11422 674 11456 708
rect 11491 674 11525 708
rect 11560 674 11594 708
rect 11629 674 11663 708
rect 11698 674 11732 708
rect 11767 674 11801 708
rect 11836 674 11870 708
rect 11905 674 11939 708
rect 11974 674 12008 708
rect 12043 674 12077 708
rect 12112 674 12146 708
rect 12181 674 12215 708
rect 12250 674 12284 708
rect 12318 674 12352 708
rect 12386 674 12420 708
rect 12454 674 12488 708
rect 12522 674 12556 708
rect 12590 674 12624 708
rect 12658 674 12692 708
rect 12726 674 12760 708
rect 12794 674 12828 708
rect 12862 674 12896 708
rect 12930 674 12964 708
rect 12998 674 13032 708
rect 13066 674 13100 708
rect 13134 674 13168 708
rect 13202 674 13236 708
rect 13270 674 13304 708
rect 13338 674 13372 708
rect 13406 674 13440 708
rect 13474 674 13508 708
rect 13542 674 13576 708
rect 13610 674 13644 708
rect 13678 674 13712 708
rect 13746 674 13780 708
rect 13814 674 13848 708
rect 13882 674 13916 708
rect 13950 674 13984 708
rect 14018 674 14052 708
rect 14086 674 14120 708
rect 14154 674 14188 708
rect 14222 674 14256 708
rect 14290 674 14324 708
rect 14358 674 14392 708
rect 14426 674 14460 708
rect 14494 674 14528 708
rect 14562 674 14596 708
rect 14630 674 14664 708
rect 14698 674 14732 708
<< locali >>
rect 17430 11598 17677 14647
rect 17430 4564 17464 11598
rect -2750 4498 -214 4564
rect -2716 4464 -2680 4498
rect -2646 4464 -2610 4498
rect -2576 4464 -2540 4498
rect -2506 4464 -2470 4498
rect -2436 4464 -2400 4498
rect -2366 4464 -2330 4498
rect -2296 4464 -2260 4498
rect -2226 4464 -2190 4498
rect -2156 4464 -2120 4498
rect -2086 4464 -2050 4498
rect -2016 4464 -1980 4498
rect -1946 4464 -1910 4498
rect -1876 4464 -1840 4498
rect -1806 4464 -1770 4498
rect -1736 4464 -1700 4498
rect -1666 4464 -1630 4498
rect -1596 4464 -1560 4498
rect -1526 4464 -1490 4498
rect -1456 4464 -1421 4498
rect -1387 4464 -1352 4498
rect -1318 4464 -1283 4498
rect -1249 4464 -1214 4498
rect -1180 4464 -1145 4498
rect -1111 4464 -1076 4498
rect -1042 4464 -1007 4498
rect -973 4464 -938 4498
rect -904 4464 -869 4498
rect -835 4464 -800 4498
rect -766 4464 -731 4498
rect -697 4464 -662 4498
rect -628 4464 -593 4498
rect -559 4464 -524 4498
rect -490 4464 -455 4498
rect -421 4464 -386 4498
rect -352 4464 -317 4498
rect -283 4464 -248 4498
rect 2094 4529 4448 4555
rect 2094 4528 4449 4529
rect 2094 4494 2304 4528
rect 2338 4494 2374 4528
rect 2408 4494 2444 4528
rect 2478 4494 2514 4528
rect 2548 4494 2584 4528
rect 2618 4494 2654 4528
rect 2688 4494 2724 4528
rect 2758 4494 2794 4528
rect 2828 4494 2864 4528
rect 2898 4494 2934 4528
rect 2968 4494 3004 4528
rect 3038 4494 3074 4528
rect 3108 4494 3144 4528
rect 3178 4494 3214 4528
rect 3248 4494 3284 4528
rect 3318 4494 3354 4528
rect 3388 4494 3424 4528
rect 3458 4494 3494 4528
rect 3528 4494 3563 4528
rect 3597 4494 3632 4528
rect 3666 4494 3701 4528
rect 3735 4494 3770 4528
rect 3804 4494 3839 4528
rect 3873 4501 3908 4528
rect 3942 4501 3977 4528
rect 4011 4501 4046 4528
rect 3873 4494 3891 4501
rect 3942 4494 3967 4501
rect 4011 4494 4043 4501
rect 4080 4494 4115 4528
rect 4149 4501 4184 4528
rect 4218 4501 4253 4528
rect 4287 4501 4322 4528
rect 4356 4501 4391 4528
rect 4425 4501 4449 4528
rect 11158 4504 11698 4528
rect 4153 4494 4184 4501
rect 4229 4494 4253 4501
rect 4305 4494 4322 4501
rect 4381 4494 4391 4501
rect 2094 4474 3891 4494
rect -2750 4428 -214 4464
rect -2716 4394 -2680 4428
rect -2646 4394 -2610 4428
rect -2576 4394 -2540 4428
rect -2506 4394 -2470 4428
rect -2436 4394 -2400 4428
rect -2366 4394 -2330 4428
rect -2296 4394 -2260 4428
rect -2226 4394 -2190 4428
rect -2156 4394 -2120 4428
rect -2086 4394 -2050 4428
rect -2016 4394 -1980 4428
rect -1946 4394 -1910 4428
rect -1876 4394 -1840 4428
rect -1806 4394 -1770 4428
rect -1736 4394 -1700 4428
rect -1666 4394 -1630 4428
rect -1596 4394 -1560 4428
rect -1526 4394 -1490 4428
rect -1456 4394 -1421 4428
rect -1387 4394 -1352 4428
rect -1318 4394 -1283 4428
rect -1249 4394 -1214 4428
rect -1180 4394 -1145 4428
rect -1111 4394 -1076 4428
rect -1042 4394 -1007 4428
rect -973 4394 -938 4428
rect -904 4394 -869 4428
rect -835 4394 -800 4428
rect -766 4394 -731 4428
rect -697 4394 -662 4428
rect -628 4394 -593 4428
rect -559 4394 -524 4428
rect -490 4394 -455 4428
rect -421 4394 -386 4428
rect -352 4394 -317 4428
rect -283 4394 -248 4428
rect -2750 4358 -214 4394
rect -2716 4324 -2680 4358
rect -2646 4324 -2610 4358
rect -2576 4324 -2540 4358
rect -2506 4324 -2470 4358
rect -2436 4324 -2400 4358
rect -2366 4324 -2330 4358
rect -2296 4324 -2260 4358
rect -2226 4324 -2190 4358
rect -2156 4324 -2120 4358
rect -2086 4324 -2050 4358
rect -2016 4324 -1980 4358
rect -1946 4324 -1910 4358
rect -1876 4324 -1840 4358
rect -1806 4324 -1770 4358
rect -1736 4324 -1700 4358
rect -1666 4324 -1630 4358
rect -1596 4324 -1560 4358
rect -1526 4324 -1490 4358
rect -1456 4324 -1421 4358
rect -1387 4324 -1352 4358
rect -1318 4324 -1283 4358
rect -1249 4324 -1214 4358
rect -1180 4324 -1145 4358
rect -1111 4324 -1076 4358
rect -1042 4324 -1007 4358
rect -973 4324 -938 4358
rect -904 4324 -869 4358
rect -835 4324 -800 4358
rect -766 4324 -731 4358
rect -697 4324 -662 4358
rect -628 4324 -593 4358
rect -559 4324 -524 4358
rect -490 4324 -455 4358
rect -421 4324 -386 4358
rect -352 4324 -317 4358
rect -283 4324 -248 4358
rect -2750 4288 -214 4324
rect -2716 4254 -2680 4288
rect -2646 4254 -2610 4288
rect -2576 4254 -2540 4288
rect -2506 4254 -2470 4288
rect -2436 4254 -2400 4288
rect -2366 4254 -2330 4288
rect -2296 4254 -2260 4288
rect -2226 4254 -2190 4288
rect -2156 4254 -2120 4288
rect -2086 4254 -2050 4288
rect -2016 4254 -1980 4288
rect -1946 4254 -1910 4288
rect -1876 4254 -1840 4288
rect -1806 4254 -1770 4288
rect -1736 4254 -1700 4288
rect -1666 4254 -1630 4288
rect -1596 4254 -1560 4288
rect -1526 4254 -1490 4288
rect -1456 4254 -1421 4288
rect -1387 4254 -1352 4288
rect -1318 4254 -1283 4288
rect -1249 4254 -1214 4288
rect -1180 4254 -1145 4288
rect -1111 4254 -1076 4288
rect -1042 4254 -1007 4288
rect -973 4254 -938 4288
rect -904 4254 -869 4288
rect -835 4254 -800 4288
rect -766 4254 -731 4288
rect -697 4254 -662 4288
rect -628 4254 -593 4288
rect -559 4254 -524 4288
rect -490 4254 -455 4288
rect -421 4254 -386 4288
rect -352 4254 -317 4288
rect -283 4254 -248 4288
rect -2750 4218 -214 4254
rect -2716 4184 -2680 4218
rect -2646 4184 -2610 4218
rect -2576 4184 -2540 4218
rect -2506 4184 -2470 4218
rect -2436 4184 -2400 4218
rect -2366 4184 -2330 4218
rect -2296 4184 -2260 4218
rect -2226 4184 -2190 4218
rect -2156 4184 -2120 4218
rect -2086 4184 -2050 4218
rect -2016 4184 -1980 4218
rect -1946 4184 -1910 4218
rect -1876 4184 -1840 4218
rect -1806 4184 -1770 4218
rect -1736 4184 -1700 4218
rect -1666 4184 -1630 4218
rect -1596 4184 -1560 4218
rect -1526 4184 -1490 4218
rect -1456 4184 -1421 4218
rect -1387 4184 -1352 4218
rect -1318 4184 -1283 4218
rect -1249 4184 -1214 4218
rect -1180 4184 -1145 4218
rect -1111 4184 -1076 4218
rect -1042 4184 -1007 4218
rect -973 4184 -938 4218
rect -904 4184 -869 4218
rect -835 4184 -800 4218
rect -766 4184 -731 4218
rect -697 4184 -662 4218
rect -628 4184 -593 4218
rect -559 4184 -524 4218
rect -490 4184 -455 4218
rect -421 4184 -386 4218
rect -352 4184 -317 4218
rect -283 4184 -248 4218
rect -2750 4148 -214 4184
rect -2716 4114 -2680 4148
rect -2646 4114 -2610 4148
rect -2576 4114 -2540 4148
rect -2506 4114 -2470 4148
rect -2436 4114 -2400 4148
rect -2366 4114 -2330 4148
rect -2296 4114 -2260 4148
rect -2226 4114 -2190 4148
rect -2156 4114 -2120 4148
rect -2086 4114 -2050 4148
rect -2016 4114 -1980 4148
rect -1946 4114 -1910 4148
rect -1876 4114 -1840 4148
rect -1806 4114 -1770 4148
rect -1736 4114 -1700 4148
rect -1666 4114 -1630 4148
rect -1596 4114 -1560 4148
rect -1526 4114 -1490 4148
rect -1456 4114 -1421 4148
rect -1387 4114 -1352 4148
rect -1318 4114 -1283 4148
rect -1249 4114 -1214 4148
rect -1180 4114 -1145 4148
rect -1111 4114 -1076 4148
rect -1042 4114 -1007 4148
rect -973 4114 -938 4148
rect -904 4114 -869 4148
rect -835 4114 -800 4148
rect -766 4114 -731 4148
rect -697 4114 -662 4148
rect -628 4114 -593 4148
rect -559 4114 -524 4148
rect -490 4114 -455 4148
rect -421 4114 -386 4148
rect -352 4114 -317 4148
rect -283 4114 -248 4148
rect 2262 4467 3891 4474
rect 3925 4467 3967 4494
rect 4001 4467 4043 4494
rect 4077 4467 4119 4494
rect 4153 4467 4195 4494
rect 4229 4467 4271 4494
rect 4305 4467 4347 4494
rect 4381 4467 4423 4494
rect 4457 4467 4499 4501
rect 4533 4467 4534 4501
rect 2262 4460 4534 4467
rect 2262 4426 2304 4460
rect 2338 4426 2374 4460
rect 2408 4426 2444 4460
rect 2478 4426 2514 4460
rect 2548 4426 2584 4460
rect 2618 4426 2654 4460
rect 2688 4426 2724 4460
rect 2758 4426 2794 4460
rect 2828 4426 2864 4460
rect 2898 4426 2934 4460
rect 2968 4426 3004 4460
rect 3038 4426 3074 4460
rect 3108 4426 3144 4460
rect 3178 4426 3214 4460
rect 3248 4426 3284 4460
rect 3318 4426 3354 4460
rect 3388 4426 3424 4460
rect 3458 4426 3494 4460
rect 3528 4426 3563 4460
rect 3597 4426 3632 4460
rect 3666 4426 3701 4460
rect 3735 4426 3770 4460
rect 3804 4426 3839 4460
rect 3873 4426 3908 4460
rect 3942 4426 3977 4460
rect 4011 4426 4046 4460
rect 4080 4426 4115 4460
rect 4149 4426 4184 4460
rect 4218 4426 4253 4460
rect 4287 4426 4322 4460
rect 4356 4426 4391 4460
rect 4425 4426 4534 4460
rect 2262 4425 4534 4426
rect 2262 4392 3891 4425
rect 3925 4392 3967 4425
rect 4001 4392 4043 4425
rect 4077 4392 4119 4425
rect 4153 4392 4195 4425
rect 4229 4392 4271 4425
rect 4305 4392 4347 4425
rect 4381 4392 4423 4425
rect 2262 4358 2304 4392
rect 2338 4358 2374 4392
rect 2408 4358 2444 4392
rect 2478 4358 2514 4392
rect 2548 4358 2584 4392
rect 2618 4358 2654 4392
rect 2688 4358 2724 4392
rect 2758 4358 2794 4392
rect 2828 4358 2864 4392
rect 2898 4358 2934 4392
rect 2968 4358 3004 4392
rect 3038 4358 3074 4392
rect 3108 4358 3144 4392
rect 3178 4358 3214 4392
rect 3248 4358 3284 4392
rect 3318 4358 3354 4392
rect 3388 4358 3424 4392
rect 3458 4358 3494 4392
rect 3528 4358 3563 4392
rect 3597 4358 3632 4392
rect 3666 4358 3701 4392
rect 3735 4358 3770 4392
rect 3804 4358 3839 4392
rect 3873 4391 3891 4392
rect 3942 4391 3967 4392
rect 4011 4391 4043 4392
rect 3873 4358 3908 4391
rect 3942 4358 3977 4391
rect 4011 4358 4046 4391
rect 4080 4358 4115 4392
rect 4153 4391 4184 4392
rect 4229 4391 4253 4392
rect 4305 4391 4322 4392
rect 4381 4391 4391 4392
rect 4457 4391 4499 4425
rect 4533 4391 4534 4425
rect 4149 4358 4184 4391
rect 4218 4358 4253 4391
rect 4287 4358 4322 4391
rect 4356 4358 4391 4391
rect 4425 4358 4534 4391
rect 2262 4349 4534 4358
rect 2262 4324 3891 4349
rect 3925 4324 3967 4349
rect 4001 4324 4043 4349
rect 4077 4324 4119 4349
rect 4153 4324 4195 4349
rect 4229 4324 4271 4349
rect 4305 4324 4347 4349
rect 4381 4324 4423 4349
rect 2262 4290 2304 4324
rect 2338 4290 2374 4324
rect 2408 4290 2444 4324
rect 2478 4290 2514 4324
rect 2548 4290 2584 4324
rect 2618 4290 2654 4324
rect 2688 4290 2724 4324
rect 2758 4290 2794 4324
rect 2828 4290 2864 4324
rect 2898 4290 2934 4324
rect 2968 4290 3004 4324
rect 3038 4290 3074 4324
rect 3108 4290 3144 4324
rect 3178 4290 3214 4324
rect 3248 4290 3284 4324
rect 3318 4290 3354 4324
rect 3388 4290 3424 4324
rect 3458 4290 3494 4324
rect 3528 4290 3563 4324
rect 3597 4290 3632 4324
rect 3666 4290 3701 4324
rect 3735 4290 3770 4324
rect 3804 4290 3839 4324
rect 3873 4315 3891 4324
rect 3942 4315 3967 4324
rect 4011 4315 4043 4324
rect 3873 4290 3908 4315
rect 3942 4290 3977 4315
rect 4011 4290 4046 4315
rect 4080 4290 4115 4324
rect 4153 4315 4184 4324
rect 4229 4315 4253 4324
rect 4305 4315 4322 4324
rect 4381 4315 4391 4324
rect 4457 4315 4499 4349
rect 4533 4315 4534 4349
rect 4149 4290 4184 4315
rect 4218 4290 4253 4315
rect 4287 4290 4322 4315
rect 4356 4290 4391 4315
rect 4425 4290 4534 4315
rect 2262 4273 4534 4290
rect 2262 4256 3891 4273
rect 3925 4256 3967 4273
rect 4001 4256 4043 4273
rect 4077 4256 4119 4273
rect 4153 4256 4195 4273
rect 4229 4256 4271 4273
rect 4305 4256 4347 4273
rect 4381 4256 4423 4273
rect 2262 4222 2304 4256
rect 2338 4222 2374 4256
rect 2408 4222 2444 4256
rect 2478 4222 2514 4256
rect 2548 4222 2584 4256
rect 2618 4222 2654 4256
rect 2688 4222 2724 4256
rect 2758 4222 2794 4256
rect 2828 4222 2864 4256
rect 2898 4222 2934 4256
rect 2968 4222 3004 4256
rect 3038 4222 3074 4256
rect 3108 4222 3144 4256
rect 3178 4222 3214 4256
rect 3248 4222 3284 4256
rect 3318 4222 3354 4256
rect 3388 4222 3424 4256
rect 3458 4222 3494 4256
rect 3528 4222 3563 4256
rect 3597 4222 3632 4256
rect 3666 4222 3701 4256
rect 3735 4222 3770 4256
rect 3804 4222 3839 4256
rect 3873 4239 3891 4256
rect 3942 4239 3967 4256
rect 4011 4239 4043 4256
rect 3873 4222 3908 4239
rect 3942 4222 3977 4239
rect 4011 4222 4046 4239
rect 4080 4222 4115 4256
rect 4153 4239 4184 4256
rect 4229 4239 4253 4256
rect 4305 4239 4322 4256
rect 4381 4239 4391 4256
rect 4457 4239 4499 4273
rect 4533 4239 4534 4273
rect 4149 4222 4184 4239
rect 4218 4222 4253 4239
rect 4287 4222 4322 4239
rect 4356 4222 4391 4239
rect 4425 4222 4534 4239
rect 2262 4197 4534 4222
rect 2262 4188 3891 4197
rect 3925 4188 3967 4197
rect 4001 4188 4043 4197
rect 4077 4188 4119 4197
rect 4153 4188 4195 4197
rect 4229 4188 4271 4197
rect 4305 4188 4347 4197
rect 4381 4188 4423 4197
rect 2262 4154 2304 4188
rect 2338 4154 2374 4188
rect 2408 4154 2444 4188
rect 2478 4154 2514 4188
rect 2548 4154 2584 4188
rect 2618 4154 2654 4188
rect 2688 4154 2724 4188
rect 2758 4154 2794 4188
rect 2828 4154 2864 4188
rect 2898 4154 2934 4188
rect 2968 4154 3004 4188
rect 3038 4154 3074 4188
rect 3108 4154 3144 4188
rect 3178 4154 3214 4188
rect 3248 4154 3284 4188
rect 3318 4154 3354 4188
rect 3388 4154 3424 4188
rect 3458 4154 3494 4188
rect 3528 4154 3563 4188
rect 3597 4154 3632 4188
rect 3666 4154 3701 4188
rect 3735 4154 3770 4188
rect 3804 4154 3839 4188
rect 3873 4163 3891 4188
rect 3942 4163 3967 4188
rect 4011 4163 4043 4188
rect 3873 4154 3908 4163
rect 3942 4154 3977 4163
rect 4011 4154 4046 4163
rect 4080 4154 4115 4188
rect 4153 4163 4184 4188
rect 4229 4163 4253 4188
rect 4305 4163 4322 4188
rect 4381 4163 4391 4188
rect 4457 4163 4499 4197
rect 4533 4163 4534 4197
rect 4149 4154 4184 4163
rect 4218 4154 4253 4163
rect 4287 4154 4322 4163
rect 4356 4154 4391 4163
rect 4425 4154 4534 4163
rect -2750 4078 -214 4114
rect -2716 4044 -2680 4078
rect -2646 4044 -2610 4078
rect -2576 4044 -2540 4078
rect -2506 4044 -2470 4078
rect -2436 4044 -2400 4078
rect -2366 4044 -2330 4078
rect -2296 4044 -2260 4078
rect -2226 4044 -2190 4078
rect -2156 4044 -2120 4078
rect -2086 4044 -2050 4078
rect -2016 4044 -1980 4078
rect -1946 4044 -1910 4078
rect -1876 4044 -1840 4078
rect -1806 4044 -1770 4078
rect -1736 4044 -1700 4078
rect -1666 4044 -1630 4078
rect -1596 4044 -1560 4078
rect -1526 4044 -1490 4078
rect -1456 4044 -1421 4078
rect -1387 4044 -1352 4078
rect -1318 4044 -1283 4078
rect -1249 4044 -1214 4078
rect -1180 4044 -1145 4078
rect -1111 4044 -1076 4078
rect -1042 4044 -1007 4078
rect -973 4044 -938 4078
rect -904 4044 -869 4078
rect -835 4044 -800 4078
rect -766 4044 -731 4078
rect -697 4044 -662 4078
rect -628 4044 -593 4078
rect -559 4044 -524 4078
rect -490 4044 -455 4078
rect -421 4044 -386 4078
rect -352 4044 -317 4078
rect -283 4044 -248 4078
rect -2750 4008 -214 4044
rect 12 4110 106 4126
rect 2262 4121 4534 4154
rect 2262 4120 3891 4121
rect 3925 4120 3967 4121
rect 4001 4120 4043 4121
rect 4077 4120 4119 4121
rect 4153 4120 4195 4121
rect 4229 4120 4271 4121
rect 4305 4120 4347 4121
rect 4381 4120 4423 4121
rect 12 4076 45 4110
rect 79 4076 106 4110
rect 12 4031 106 4076
rect -2716 3974 -2680 4008
rect -2646 3974 -2610 4008
rect -2576 3974 -2540 4008
rect -2506 3974 -2470 4008
rect -2436 3974 -2400 4008
rect -2366 3974 -2330 4008
rect -2296 3974 -2260 4008
rect -2226 3974 -2190 4008
rect -2156 3974 -2120 4008
rect -2086 3974 -2050 4008
rect -2016 3974 -1980 4008
rect -1946 3974 -1910 4008
rect -1876 3974 -1840 4008
rect -1806 3974 -1770 4008
rect -1736 3974 -1700 4008
rect -1666 3974 -1630 4008
rect -1596 3974 -1560 4008
rect -1526 3974 -1490 4008
rect -1456 3974 -1421 4008
rect -1387 3974 -1352 4008
rect -1318 3974 -1283 4008
rect -1249 3974 -1214 4008
rect -1180 3974 -1145 4008
rect -1111 3974 -1076 4008
rect -1042 3974 -1007 4008
rect -973 3974 -938 4008
rect -904 3974 -869 4008
rect -835 3974 -800 4008
rect -766 3974 -731 4008
rect -697 3974 -662 4008
rect -628 3974 -593 4008
rect -559 3974 -524 4008
rect -490 3974 -455 4008
rect -421 3974 -386 4008
rect -352 3974 -317 4008
rect -283 3974 -248 4008
rect 30 3997 68 4031
rect 102 3997 106 4031
rect 443 4003 509 4110
rect 2262 4086 2304 4120
rect 2338 4086 2374 4120
rect 2408 4086 2444 4120
rect 2478 4086 2514 4120
rect 2548 4086 2584 4120
rect 2618 4086 2654 4120
rect 2688 4086 2724 4120
rect 2758 4086 2794 4120
rect 2828 4086 2864 4120
rect 2898 4086 2934 4120
rect 2968 4086 3004 4120
rect 3038 4086 3074 4120
rect 3108 4086 3144 4120
rect 3178 4086 3214 4120
rect 3248 4086 3284 4120
rect 3318 4086 3354 4120
rect 3388 4086 3424 4120
rect 3458 4086 3494 4120
rect 3528 4086 3563 4120
rect 3597 4086 3632 4120
rect 3666 4086 3701 4120
rect 3735 4086 3770 4120
rect 3804 4086 3839 4120
rect 3873 4087 3891 4120
rect 3942 4087 3967 4120
rect 4011 4087 4043 4120
rect 3873 4086 3908 4087
rect 3942 4086 3977 4087
rect 4011 4086 4046 4087
rect 4080 4086 4115 4120
rect 4153 4087 4184 4120
rect 4229 4087 4253 4120
rect 4305 4087 4322 4120
rect 4381 4087 4391 4120
rect 4457 4087 4499 4121
rect 4533 4087 4534 4121
rect 4149 4086 4184 4087
rect 4218 4086 4253 4087
rect 4287 4086 4322 4087
rect 4356 4086 4391 4087
rect 4425 4086 4534 4087
rect 2262 4052 4534 4086
rect 2262 4018 2304 4052
rect 2338 4018 2374 4052
rect 2408 4018 2444 4052
rect 2478 4018 2514 4052
rect 2548 4018 2584 4052
rect 2618 4018 2654 4052
rect 2688 4018 2724 4052
rect 2758 4018 2794 4052
rect 2828 4018 2864 4052
rect 2898 4018 2934 4052
rect 2968 4018 3004 4052
rect 3038 4018 3074 4052
rect 3108 4018 3144 4052
rect 3178 4018 3214 4052
rect 3248 4018 3284 4052
rect 3318 4018 3354 4052
rect 3388 4018 3424 4052
rect 3458 4018 3494 4052
rect 3528 4018 3563 4052
rect 3597 4018 3632 4052
rect 3666 4018 3701 4052
rect 3735 4018 3770 4052
rect 3804 4018 3839 4052
rect 3873 4045 3908 4052
rect 3942 4045 3977 4052
rect 4011 4045 4046 4052
rect 3873 4018 3891 4045
rect 3942 4018 3967 4045
rect 4011 4018 4043 4045
rect 4080 4018 4115 4052
rect 4149 4045 4184 4052
rect 4218 4045 4253 4052
rect 4287 4045 4322 4052
rect 4356 4045 4391 4052
rect 4425 4045 4534 4052
rect 4153 4018 4184 4045
rect 4229 4018 4253 4045
rect 4305 4018 4322 4045
rect 4381 4018 4391 4045
rect 2262 4011 3891 4018
rect 3925 4011 3967 4018
rect 4001 4011 4043 4018
rect 4077 4011 4119 4018
rect 4153 4011 4195 4018
rect 4229 4011 4271 4018
rect 4305 4011 4347 4018
rect 4381 4011 4423 4018
rect 4457 4011 4499 4045
rect 4533 4011 4534 4045
rect 12 3991 106 3997
rect -2750 3938 -214 3974
rect -2716 3904 -2680 3938
rect -2646 3904 -2610 3938
rect -2576 3904 -2540 3938
rect -2506 3904 -2470 3938
rect -2436 3904 -2400 3938
rect -2366 3904 -2330 3938
rect -2296 3904 -2260 3938
rect -2226 3904 -2190 3938
rect -2156 3904 -2120 3938
rect -2086 3904 -2050 3938
rect -2016 3904 -1980 3938
rect -1946 3904 -1910 3938
rect -1876 3904 -1840 3938
rect -1806 3904 -1770 3938
rect -1736 3904 -1700 3938
rect -1666 3904 -1630 3938
rect -1596 3904 -1560 3938
rect -1526 3904 -1490 3938
rect -1456 3904 -1421 3938
rect -1387 3904 -1352 3938
rect -1318 3904 -1283 3938
rect -1249 3904 -1214 3938
rect -1180 3904 -1145 3938
rect -1111 3904 -1076 3938
rect -1042 3904 -1007 3938
rect -973 3904 -938 3938
rect -904 3904 -869 3938
rect -835 3904 -800 3938
rect -766 3904 -731 3938
rect -697 3904 -662 3938
rect -628 3904 -593 3938
rect -559 3904 -524 3938
rect -490 3904 -455 3938
rect -421 3904 -386 3938
rect -352 3904 -317 3938
rect -283 3904 -248 3938
rect -2750 3868 -214 3904
rect -2716 3834 -2680 3868
rect -2646 3834 -2610 3868
rect -2576 3834 -2540 3868
rect -2506 3834 -2470 3868
rect -2436 3834 -2400 3868
rect -2366 3834 -2330 3868
rect -2296 3834 -2260 3868
rect -2226 3834 -2190 3868
rect -2156 3834 -2120 3868
rect -2086 3834 -2050 3868
rect -2016 3834 -1980 3868
rect -1946 3834 -1910 3868
rect -1876 3834 -1840 3868
rect -1806 3834 -1770 3868
rect -1736 3834 -1700 3868
rect -1666 3834 -1630 3868
rect -1596 3834 -1560 3868
rect -1526 3834 -1490 3868
rect -1456 3834 -1421 3868
rect -1387 3834 -1352 3868
rect -1318 3834 -1283 3868
rect -1249 3834 -1214 3868
rect -1180 3834 -1145 3868
rect -1111 3834 -1076 3868
rect -1042 3834 -1007 3868
rect -973 3834 -938 3868
rect -904 3834 -869 3868
rect -835 3834 -800 3868
rect -766 3834 -731 3868
rect -697 3834 -662 3868
rect -628 3834 -593 3868
rect -559 3834 -524 3868
rect -490 3834 -455 3868
rect -421 3834 -386 3868
rect -352 3834 -317 3868
rect -283 3834 -248 3868
rect -2750 3798 -214 3834
rect -2716 3764 -2680 3798
rect -2646 3764 -2610 3798
rect -2576 3764 -2540 3798
rect -2506 3764 -2470 3798
rect -2436 3764 -2400 3798
rect -2366 3764 -2330 3798
rect -2296 3764 -2260 3798
rect -2226 3764 -2190 3798
rect -2156 3764 -2120 3798
rect -2086 3764 -2050 3798
rect -2016 3764 -1980 3798
rect -1946 3764 -1910 3798
rect -1876 3764 -1840 3798
rect -1806 3764 -1770 3798
rect -1736 3764 -1700 3798
rect -1666 3764 -1630 3798
rect -1596 3764 -1560 3798
rect -1526 3764 -1490 3798
rect -1456 3764 -1421 3798
rect -1387 3764 -1352 3798
rect -1318 3764 -1283 3798
rect -1249 3764 -1214 3798
rect -1180 3764 -1145 3798
rect -1111 3764 -1076 3798
rect -1042 3764 -1007 3798
rect -973 3764 -938 3798
rect -904 3764 -869 3798
rect -835 3764 -800 3798
rect -766 3764 -731 3798
rect -697 3764 -662 3798
rect -628 3764 -593 3798
rect -559 3764 -524 3798
rect -490 3764 -455 3798
rect -421 3764 -386 3798
rect -352 3764 -317 3798
rect -283 3764 -248 3798
rect -2750 3728 -214 3764
rect -2716 3694 -2680 3728
rect -2646 3694 -2610 3728
rect -2576 3694 -2540 3728
rect -2506 3694 -2470 3728
rect -2436 3694 -2400 3728
rect -2366 3694 -2330 3728
rect -2296 3694 -2260 3728
rect -2226 3694 -2190 3728
rect -2156 3694 -2120 3728
rect -2086 3694 -2050 3728
rect -2016 3694 -1980 3728
rect -1946 3694 -1910 3728
rect -1876 3694 -1840 3728
rect -1806 3694 -1770 3728
rect -1736 3694 -1700 3728
rect -1666 3694 -1630 3728
rect -1596 3694 -1560 3728
rect -1526 3694 -1490 3728
rect -1456 3694 -1421 3728
rect -1387 3694 -1352 3728
rect -1318 3694 -1283 3728
rect -1249 3694 -1214 3728
rect -1180 3694 -1145 3728
rect -1111 3694 -1076 3728
rect -1042 3694 -1007 3728
rect -973 3694 -938 3728
rect -904 3694 -869 3728
rect -835 3694 -800 3728
rect -766 3694 -731 3728
rect -697 3694 -662 3728
rect -628 3694 -593 3728
rect -559 3694 -524 3728
rect -490 3694 -455 3728
rect -421 3694 -386 3728
rect -352 3694 -317 3728
rect -283 3694 -248 3728
rect -2750 3658 -214 3694
rect -2716 3624 -2680 3658
rect -2646 3624 -2610 3658
rect -2576 3624 -2540 3658
rect -2506 3624 -2470 3658
rect -2436 3624 -2400 3658
rect -2366 3624 -2330 3658
rect -2296 3624 -2260 3658
rect -2226 3624 -2190 3658
rect -2156 3624 -2120 3658
rect -2086 3624 -2050 3658
rect -2016 3624 -1980 3658
rect -1946 3624 -1910 3658
rect -1876 3624 -1840 3658
rect -1806 3624 -1770 3658
rect -1736 3624 -1700 3658
rect -1666 3624 -1630 3658
rect -1596 3624 -1560 3658
rect -1526 3624 -1490 3658
rect -1456 3624 -1421 3658
rect -1387 3624 -1352 3658
rect -1318 3624 -1283 3658
rect -1249 3624 -1214 3658
rect -1180 3624 -1145 3658
rect -1111 3624 -1076 3658
rect -1042 3624 -1007 3658
rect -973 3624 -938 3658
rect -904 3624 -869 3658
rect -835 3624 -800 3658
rect -766 3624 -731 3658
rect -697 3624 -662 3658
rect -628 3624 -593 3658
rect -559 3624 -524 3658
rect -490 3624 -455 3658
rect -421 3624 -386 3658
rect -352 3624 -317 3658
rect -283 3624 -248 3658
rect -2750 3588 -214 3624
rect -2716 3554 -2680 3588
rect -2646 3554 -2610 3588
rect -2576 3554 -2540 3588
rect -2506 3554 -2470 3588
rect -2436 3554 -2400 3588
rect -2366 3554 -2330 3588
rect -2296 3554 -2260 3588
rect -2226 3554 -2190 3588
rect -2156 3554 -2120 3588
rect -2086 3554 -2050 3588
rect -2016 3554 -1980 3588
rect -1946 3554 -1910 3588
rect -1876 3554 -1840 3588
rect -1806 3554 -1770 3588
rect -1736 3554 -1700 3588
rect -1666 3554 -1630 3588
rect -1596 3554 -1560 3588
rect -1526 3554 -1490 3588
rect -1456 3554 -1421 3588
rect -1387 3554 -1352 3588
rect -1318 3554 -1283 3588
rect -1249 3554 -1214 3588
rect -1180 3554 -1145 3588
rect -1111 3554 -1076 3588
rect -1042 3554 -1007 3588
rect -973 3554 -938 3588
rect -904 3554 -869 3588
rect -835 3554 -800 3588
rect -766 3554 -731 3588
rect -697 3554 -662 3588
rect -628 3554 -593 3588
rect -559 3554 -524 3588
rect -490 3554 -455 3588
rect -421 3554 -386 3588
rect -352 3554 -317 3588
rect -283 3554 -248 3588
rect -2750 3518 -214 3554
rect -2716 3484 -2680 3518
rect -2646 3484 -2610 3518
rect -2576 3484 -2540 3518
rect -2506 3484 -2470 3518
rect -2436 3484 -2400 3518
rect -2366 3484 -2330 3518
rect -2296 3484 -2260 3518
rect -2226 3484 -2190 3518
rect -2156 3484 -2120 3518
rect -2086 3484 -2050 3518
rect -2016 3484 -1980 3518
rect -1946 3484 -1910 3518
rect -1876 3484 -1840 3518
rect -1806 3484 -1770 3518
rect -1736 3484 -1700 3518
rect -1666 3484 -1630 3518
rect -1596 3484 -1560 3518
rect -1526 3484 -1490 3518
rect -1456 3484 -1421 3518
rect -1387 3484 -1352 3518
rect -1318 3484 -1283 3518
rect -1249 3484 -1214 3518
rect -1180 3484 -1145 3518
rect -1111 3484 -1076 3518
rect -1042 3484 -1007 3518
rect -973 3484 -938 3518
rect -904 3484 -869 3518
rect -835 3484 -800 3518
rect -766 3484 -731 3518
rect -697 3484 -662 3518
rect -628 3484 -593 3518
rect -559 3484 -524 3518
rect -490 3484 -455 3518
rect -421 3484 -386 3518
rect -352 3484 -317 3518
rect -283 3484 -248 3518
rect -2750 3448 -214 3484
rect -2716 3414 -2680 3448
rect -2646 3414 -2610 3448
rect -2576 3414 -2540 3448
rect -2506 3414 -2470 3448
rect -2436 3414 -2400 3448
rect -2366 3414 -2330 3448
rect -2296 3414 -2260 3448
rect -2226 3414 -2190 3448
rect -2156 3414 -2120 3448
rect -2086 3414 -2050 3448
rect -2016 3414 -1980 3448
rect -1946 3414 -1910 3448
rect -1876 3414 -1840 3448
rect -1806 3414 -1770 3448
rect -1736 3414 -1700 3448
rect -1666 3414 -1630 3448
rect -1596 3414 -1560 3448
rect -1526 3414 -1490 3448
rect -1456 3414 -1421 3448
rect -1387 3414 -1352 3448
rect -1318 3414 -1283 3448
rect -1249 3414 -1214 3448
rect -1180 3414 -1145 3448
rect -1111 3414 -1076 3448
rect -1042 3414 -1007 3448
rect -973 3414 -938 3448
rect -904 3414 -869 3448
rect -835 3414 -800 3448
rect -766 3414 -731 3448
rect -697 3414 -662 3448
rect -628 3414 -593 3448
rect -559 3414 -524 3448
rect -490 3414 -455 3448
rect -421 3414 -386 3448
rect -352 3414 -317 3448
rect -283 3414 -248 3448
rect -2750 3378 -214 3414
rect 2262 3984 4534 4011
rect 2262 3950 2304 3984
rect 2338 3950 2374 3984
rect 2408 3950 2444 3984
rect 2478 3950 2514 3984
rect 2548 3950 2584 3984
rect 2618 3950 2654 3984
rect 2688 3950 2724 3984
rect 2758 3950 2794 3984
rect 2828 3950 2864 3984
rect 2898 3950 2934 3984
rect 2968 3950 3004 3984
rect 3038 3950 3074 3984
rect 3108 3950 3144 3984
rect 3178 3950 3214 3984
rect 3248 3950 3284 3984
rect 3318 3950 3354 3984
rect 3388 3950 3424 3984
rect 3458 3950 3494 3984
rect 3528 3950 3563 3984
rect 3597 3950 3632 3984
rect 3666 3950 3701 3984
rect 3735 3950 3770 3984
rect 3804 3950 3839 3984
rect 3873 3968 3908 3984
rect 3942 3968 3977 3984
rect 4011 3968 4046 3984
rect 3873 3950 3891 3968
rect 3942 3950 3967 3968
rect 4011 3950 4043 3968
rect 4080 3950 4115 3984
rect 4149 3968 4184 3984
rect 4218 3968 4253 3984
rect 4287 3968 4322 3984
rect 4356 3968 4391 3984
rect 4425 3968 4534 3984
rect 4153 3950 4184 3968
rect 4229 3950 4253 3968
rect 4305 3950 4322 3968
rect 4381 3950 4391 3968
rect 2262 3934 3891 3950
rect 3925 3934 3967 3950
rect 4001 3934 4043 3950
rect 4077 3934 4119 3950
rect 4153 3934 4195 3950
rect 4229 3934 4271 3950
rect 4305 3934 4347 3950
rect 4381 3934 4423 3950
rect 4457 3934 4499 3968
rect 4533 3934 4534 3968
rect 2262 3916 4534 3934
rect 2262 3882 2304 3916
rect 2338 3882 2374 3916
rect 2408 3882 2444 3916
rect 2478 3882 2514 3916
rect 2548 3882 2584 3916
rect 2618 3882 2654 3916
rect 2688 3882 2724 3916
rect 2758 3882 2794 3916
rect 2828 3882 2864 3916
rect 2898 3882 2934 3916
rect 2968 3882 3004 3916
rect 3038 3882 3074 3916
rect 3108 3882 3144 3916
rect 3178 3882 3214 3916
rect 3248 3882 3284 3916
rect 3318 3882 3354 3916
rect 3388 3882 3424 3916
rect 3458 3882 3494 3916
rect 3528 3882 3563 3916
rect 3597 3882 3632 3916
rect 3666 3882 3701 3916
rect 3735 3882 3770 3916
rect 3804 3882 3839 3916
rect 3873 3891 3908 3916
rect 3942 3891 3977 3916
rect 4011 3891 4046 3916
rect 3873 3882 3891 3891
rect 3942 3882 3967 3891
rect 4011 3882 4043 3891
rect 4080 3882 4115 3916
rect 4149 3891 4184 3916
rect 4218 3891 4253 3916
rect 4287 3891 4322 3916
rect 4356 3891 4391 3916
rect 4425 3891 4534 3916
rect 4153 3882 4184 3891
rect 4229 3882 4253 3891
rect 4305 3882 4322 3891
rect 4381 3882 4391 3891
rect 2262 3857 3891 3882
rect 3925 3857 3967 3882
rect 4001 3857 4043 3882
rect 4077 3857 4119 3882
rect 4153 3857 4195 3882
rect 4229 3857 4271 3882
rect 4305 3857 4347 3882
rect 4381 3857 4423 3882
rect 4457 3857 4499 3891
rect 4533 3857 4534 3891
rect 11158 4470 11159 4504
rect 11193 4470 11231 4504
rect 11265 4470 11303 4504
rect 11337 4470 11375 4504
rect 11409 4470 11447 4504
rect 11481 4470 11519 4504
rect 11553 4470 11591 4504
rect 11625 4470 11663 4504
rect 11697 4470 11698 4504
rect 11158 4434 11698 4470
rect 11158 4400 11159 4434
rect 11193 4400 11231 4434
rect 11265 4400 11303 4434
rect 11337 4400 11375 4434
rect 11409 4400 11447 4434
rect 11481 4400 11519 4434
rect 11553 4400 11591 4434
rect 11625 4400 11663 4434
rect 11697 4400 11698 4434
rect 11158 4364 11698 4400
rect 11158 4330 11159 4364
rect 11193 4330 11231 4364
rect 11265 4330 11303 4364
rect 11337 4330 11375 4364
rect 11409 4330 11447 4364
rect 11481 4330 11519 4364
rect 11553 4330 11591 4364
rect 11625 4330 11663 4364
rect 11697 4330 11698 4364
rect 11158 4294 11698 4330
rect 11158 4260 11159 4294
rect 11193 4260 11231 4294
rect 11265 4260 11303 4294
rect 11337 4260 11375 4294
rect 11409 4260 11447 4294
rect 11481 4260 11519 4294
rect 11553 4260 11591 4294
rect 11625 4260 11663 4294
rect 11697 4260 11698 4294
rect 11158 4223 11698 4260
rect 11158 4189 11159 4223
rect 11193 4189 11231 4223
rect 11265 4189 11303 4223
rect 11337 4189 11375 4223
rect 11409 4189 11447 4223
rect 11481 4189 11519 4223
rect 11553 4189 11591 4223
rect 11625 4189 11663 4223
rect 11697 4189 11698 4223
rect 11158 4152 11698 4189
rect 11158 4118 11159 4152
rect 11193 4118 11231 4152
rect 11265 4118 11303 4152
rect 11337 4118 11375 4152
rect 11409 4118 11447 4152
rect 11481 4118 11519 4152
rect 11553 4118 11591 4152
rect 11625 4118 11663 4152
rect 11697 4118 11698 4152
rect 11158 4081 11698 4118
rect 11158 4047 11159 4081
rect 11193 4047 11231 4081
rect 11265 4047 11303 4081
rect 11337 4047 11375 4081
rect 11409 4047 11447 4081
rect 11481 4047 11519 4081
rect 11553 4047 11591 4081
rect 11625 4047 11663 4081
rect 11697 4047 11698 4081
rect 11158 4010 11698 4047
rect 11158 3976 11159 4010
rect 11193 3976 11231 4010
rect 11265 3976 11303 4010
rect 11337 3976 11375 4010
rect 11409 3976 11447 4010
rect 11481 3976 11519 4010
rect 11553 3976 11591 4010
rect 11625 3976 11663 4010
rect 11697 3976 11698 4010
rect 11158 3939 11698 3976
rect 11158 3905 11159 3939
rect 11193 3905 11231 3939
rect 11265 3905 11303 3939
rect 11337 3905 11375 3939
rect 11409 3905 11447 3939
rect 11481 3905 11519 3939
rect 11553 3905 11591 3939
rect 11625 3905 11663 3939
rect 11697 3905 11698 3939
rect 11158 3868 11698 3905
rect 2262 3848 4449 3857
rect 2262 3814 2304 3848
rect 2338 3814 2374 3848
rect 2408 3814 2444 3848
rect 2478 3814 2514 3848
rect 2548 3814 2584 3848
rect 2618 3814 2654 3848
rect 2688 3814 2724 3848
rect 2758 3814 2794 3848
rect 2828 3814 2864 3848
rect 2898 3814 2934 3848
rect 2968 3814 3004 3848
rect 3038 3814 3074 3848
rect 3108 3814 3144 3848
rect 3178 3814 3214 3848
rect 3248 3814 3284 3848
rect 3318 3814 3354 3848
rect 3388 3814 3424 3848
rect 3458 3814 3494 3848
rect 3528 3814 3563 3848
rect 3597 3814 3632 3848
rect 3666 3814 3701 3848
rect 3735 3814 3770 3848
rect 3804 3814 3839 3848
rect 3873 3814 3908 3848
rect 3942 3814 3977 3848
rect 4011 3814 4046 3848
rect 4080 3814 4115 3848
rect 4149 3814 4184 3848
rect 4218 3814 4253 3848
rect 4287 3814 4322 3848
rect 4356 3814 4391 3848
rect 4425 3814 4449 3848
rect 2262 3780 4449 3814
rect 2262 3746 2304 3780
rect 2338 3746 2374 3780
rect 2408 3746 2444 3780
rect 2478 3746 2514 3780
rect 2548 3746 2584 3780
rect 2618 3746 2654 3780
rect 2688 3746 2724 3780
rect 2758 3746 2794 3780
rect 2828 3746 2864 3780
rect 2898 3746 2934 3780
rect 2968 3746 3004 3780
rect 3038 3746 3074 3780
rect 3108 3746 3144 3780
rect 3178 3746 3214 3780
rect 3248 3746 3284 3780
rect 3318 3746 3354 3780
rect 3388 3746 3424 3780
rect 3458 3746 3494 3780
rect 3528 3746 3563 3780
rect 3597 3746 3632 3780
rect 3666 3746 3701 3780
rect 3735 3746 3770 3780
rect 3804 3746 3839 3780
rect 3873 3746 3908 3780
rect 3942 3746 3977 3780
rect 4011 3746 4046 3780
rect 4080 3746 4115 3780
rect 4149 3746 4184 3780
rect 4218 3746 4253 3780
rect 4287 3746 4322 3780
rect 4356 3746 4391 3780
rect 4425 3746 4449 3780
rect 2262 3712 4449 3746
rect 2262 3678 2304 3712
rect 2338 3678 2374 3712
rect 2408 3678 2444 3712
rect 2478 3678 2514 3712
rect 2548 3678 2584 3712
rect 2618 3678 2654 3712
rect 2688 3678 2724 3712
rect 2758 3678 2794 3712
rect 2828 3678 2864 3712
rect 2898 3678 2934 3712
rect 2968 3678 3004 3712
rect 3038 3678 3074 3712
rect 3108 3678 3144 3712
rect 3178 3678 3214 3712
rect 3248 3678 3284 3712
rect 3318 3678 3354 3712
rect 3388 3678 3424 3712
rect 3458 3678 3494 3712
rect 3528 3678 3563 3712
rect 3597 3678 3632 3712
rect 3666 3678 3701 3712
rect 3735 3678 3770 3712
rect 3804 3678 3839 3712
rect 3873 3678 3908 3712
rect 3942 3678 3977 3712
rect 4011 3678 4046 3712
rect 4080 3678 4115 3712
rect 4149 3678 4184 3712
rect 4218 3678 4253 3712
rect 4287 3678 4322 3712
rect 4356 3678 4391 3712
rect 4425 3678 4449 3712
rect 2262 3644 4449 3678
rect 2262 3610 2304 3644
rect 2338 3610 2374 3644
rect 2408 3610 2444 3644
rect 2478 3610 2514 3644
rect 2548 3610 2584 3644
rect 2618 3610 2654 3644
rect 2688 3610 2724 3644
rect 2758 3610 2794 3644
rect 2828 3610 2864 3644
rect 2898 3610 2934 3644
rect 2968 3610 3004 3644
rect 3038 3610 3074 3644
rect 3108 3610 3144 3644
rect 3178 3610 3214 3644
rect 3248 3610 3284 3644
rect 3318 3610 3354 3644
rect 3388 3610 3424 3644
rect 3458 3610 3494 3644
rect 3528 3610 3563 3644
rect 3597 3610 3632 3644
rect 3666 3610 3701 3644
rect 3735 3610 3770 3644
rect 3804 3610 3839 3644
rect 3873 3610 3908 3644
rect 3942 3610 3977 3644
rect 4011 3610 4046 3644
rect 4080 3610 4115 3644
rect 4149 3610 4184 3644
rect 4218 3610 4253 3644
rect 4287 3610 4322 3644
rect 4356 3610 4391 3644
rect 4425 3610 4449 3644
rect 2262 3576 4449 3610
rect 11158 3834 11159 3868
rect 11193 3834 11231 3868
rect 11265 3834 11303 3868
rect 11337 3834 11375 3868
rect 11409 3834 11447 3868
rect 11481 3834 11519 3868
rect 11553 3834 11591 3868
rect 11625 3834 11663 3868
rect 11697 3834 11698 3868
rect 11158 3797 11698 3834
rect 11158 3763 11159 3797
rect 11193 3763 11231 3797
rect 11265 3763 11303 3797
rect 11337 3763 11375 3797
rect 11409 3763 11447 3797
rect 11481 3763 11519 3797
rect 11553 3763 11591 3797
rect 11625 3763 11663 3797
rect 11697 3763 11698 3797
rect 11158 3726 11698 3763
rect 11158 3692 11159 3726
rect 11193 3692 11231 3726
rect 11265 3692 11303 3726
rect 11337 3692 11375 3726
rect 11409 3692 11447 3726
rect 11481 3692 11519 3726
rect 11553 3692 11591 3726
rect 11625 3692 11663 3726
rect 11697 3692 11698 3726
rect 11158 3655 11698 3692
rect 11158 3621 11159 3655
rect 11193 3621 11231 3655
rect 11265 3621 11303 3655
rect 11337 3621 11375 3655
rect 11409 3621 11447 3655
rect 11481 3621 11519 3655
rect 11553 3621 11591 3655
rect 11625 3621 11663 3655
rect 11697 3621 11698 3655
rect 11158 3597 11698 3621
rect 11929 4324 17215 4378
rect 11929 4322 11949 4324
rect 11983 4322 12018 4324
rect 12052 4322 12087 4324
rect 11929 4288 11937 4322
rect 11983 4290 12010 4322
rect 12052 4290 12083 4322
rect 12121 4290 12156 4324
rect 12190 4290 12225 4324
rect 12259 4322 12294 4324
rect 12328 4322 12363 4324
rect 12397 4322 12432 4324
rect 12466 4322 12501 4324
rect 12535 4322 12570 4324
rect 12604 4322 12639 4324
rect 12673 4322 12708 4324
rect 12742 4322 12777 4324
rect 12263 4290 12294 4322
rect 12336 4290 12363 4322
rect 12409 4290 12432 4322
rect 12482 4290 12501 4322
rect 12555 4290 12570 4322
rect 12628 4290 12639 4322
rect 12701 4290 12708 4322
rect 12774 4290 12777 4322
rect 12811 4322 12846 4324
rect 12880 4322 12915 4324
rect 12949 4322 12984 4324
rect 13018 4322 13053 4324
rect 13087 4322 13122 4324
rect 13156 4322 13191 4324
rect 13225 4322 13260 4324
rect 13294 4322 13329 4324
rect 13363 4322 13398 4324
rect 12811 4290 12813 4322
rect 12880 4290 12886 4322
rect 12949 4290 12959 4322
rect 13018 4290 13032 4322
rect 13087 4290 13105 4322
rect 13156 4290 13178 4322
rect 13225 4290 13251 4322
rect 13294 4290 13324 4322
rect 13363 4290 13397 4322
rect 13432 4290 13467 4324
rect 13501 4322 13536 4324
rect 13570 4322 13605 4324
rect 13639 4322 13674 4324
rect 13708 4322 13743 4324
rect 13777 4322 13812 4324
rect 13846 4322 13881 4324
rect 13915 4322 13950 4324
rect 13984 4322 14019 4324
rect 13504 4290 13536 4322
rect 13577 4290 13605 4322
rect 13650 4290 13674 4322
rect 13723 4290 13743 4322
rect 13796 4290 13812 4322
rect 13869 4290 13881 4322
rect 13942 4290 13950 4322
rect 14015 4290 14019 4322
rect 14053 4322 14088 4324
rect 14053 4290 14054 4322
rect 11971 4288 12010 4290
rect 12044 4288 12083 4290
rect 12117 4288 12156 4290
rect 12190 4288 12229 4290
rect 12263 4288 12302 4290
rect 12336 4288 12375 4290
rect 12409 4288 12448 4290
rect 12482 4288 12521 4290
rect 12555 4288 12594 4290
rect 12628 4288 12667 4290
rect 12701 4288 12740 4290
rect 12774 4288 12813 4290
rect 12847 4288 12886 4290
rect 12920 4288 12959 4290
rect 12993 4288 13032 4290
rect 13066 4288 13105 4290
rect 13139 4288 13178 4290
rect 13212 4288 13251 4290
rect 13285 4288 13324 4290
rect 13358 4288 13397 4290
rect 13431 4288 13470 4290
rect 13504 4288 13543 4290
rect 13577 4288 13616 4290
rect 13650 4288 13689 4290
rect 13723 4288 13762 4290
rect 13796 4288 13835 4290
rect 13869 4288 13908 4290
rect 13942 4288 13981 4290
rect 14015 4288 14054 4290
rect 14122 4322 14157 4324
rect 14191 4322 14226 4324
rect 14260 4322 14295 4324
rect 14329 4322 14364 4324
rect 14398 4322 14433 4324
rect 14467 4322 14502 4324
rect 14536 4322 14571 4324
rect 14605 4322 14640 4324
rect 14122 4290 14127 4322
rect 14191 4290 14200 4322
rect 14260 4290 14273 4322
rect 14329 4290 14346 4322
rect 14398 4290 14419 4322
rect 14467 4290 14492 4322
rect 14536 4290 14565 4322
rect 14605 4290 14638 4322
rect 14674 4290 14709 4324
rect 14743 4322 14778 4324
rect 14812 4322 14847 4324
rect 14881 4322 14916 4324
rect 14950 4322 14985 4324
rect 15019 4322 15054 4324
rect 15088 4322 15123 4324
rect 15157 4322 15192 4324
rect 15226 4322 15261 4324
rect 14745 4290 14778 4322
rect 14818 4290 14847 4322
rect 14891 4290 14916 4322
rect 14964 4290 14985 4322
rect 15037 4290 15054 4322
rect 15110 4290 15123 4322
rect 15183 4290 15192 4322
rect 15256 4290 15261 4322
rect 15295 4322 15330 4324
rect 14088 4288 14127 4290
rect 14161 4288 14200 4290
rect 14234 4288 14273 4290
rect 14307 4288 14346 4290
rect 14380 4288 14419 4290
rect 14453 4288 14492 4290
rect 14526 4288 14565 4290
rect 14599 4288 14638 4290
rect 14672 4288 14711 4290
rect 14745 4288 14784 4290
rect 14818 4288 14857 4290
rect 14891 4288 14930 4290
rect 14964 4288 15003 4290
rect 15037 4288 15076 4290
rect 15110 4288 15149 4290
rect 15183 4288 15222 4290
rect 15256 4288 15295 4290
rect 15329 4290 15330 4322
rect 15364 4322 15399 4324
rect 15433 4322 15468 4324
rect 15502 4322 15537 4324
rect 15571 4322 15606 4324
rect 15640 4322 15675 4324
rect 15709 4322 15744 4324
rect 15778 4322 15813 4324
rect 15847 4322 15882 4324
rect 15364 4290 15368 4322
rect 15433 4290 15441 4322
rect 15502 4290 15514 4322
rect 15571 4290 15587 4322
rect 15640 4290 15660 4322
rect 15709 4290 15733 4322
rect 15778 4290 15806 4322
rect 15847 4290 15879 4322
rect 15916 4290 15951 4324
rect 15985 4322 16020 4324
rect 16054 4322 16089 4324
rect 16123 4322 16158 4324
rect 16192 4322 16227 4324
rect 16261 4322 16296 4324
rect 16330 4322 16365 4324
rect 15986 4290 16020 4322
rect 16059 4290 16089 4322
rect 16132 4290 16158 4322
rect 16205 4290 16227 4322
rect 16278 4290 16296 4322
rect 15329 4288 15368 4290
rect 15402 4288 15441 4290
rect 15475 4288 15514 4290
rect 15548 4288 15587 4290
rect 15621 4288 15660 4290
rect 15694 4288 15733 4290
rect 15767 4288 15806 4290
rect 15840 4288 15879 4290
rect 15913 4288 15952 4290
rect 15986 4288 16025 4290
rect 16059 4288 16098 4290
rect 16132 4288 16171 4290
rect 16205 4288 16244 4290
rect 16278 4288 16317 4290
rect 16351 4288 16365 4322
rect 11929 4256 16365 4288
rect 11929 4250 11949 4256
rect 11983 4250 12018 4256
rect 12052 4250 12087 4256
rect 11929 4216 11937 4250
rect 11983 4222 12010 4250
rect 12052 4222 12083 4250
rect 12121 4222 12156 4256
rect 12190 4222 12225 4256
rect 12259 4250 12294 4256
rect 12328 4250 12363 4256
rect 12397 4250 12432 4256
rect 12466 4250 12501 4256
rect 12535 4250 12570 4256
rect 12604 4250 12639 4256
rect 12673 4250 12708 4256
rect 12742 4250 12777 4256
rect 12263 4222 12294 4250
rect 12336 4222 12363 4250
rect 12409 4222 12432 4250
rect 12482 4222 12501 4250
rect 12555 4222 12570 4250
rect 12628 4222 12639 4250
rect 12701 4222 12708 4250
rect 12774 4222 12777 4250
rect 12811 4250 12846 4256
rect 12880 4250 12915 4256
rect 12949 4250 12984 4256
rect 13018 4250 13053 4256
rect 13087 4250 13122 4256
rect 13156 4250 13191 4256
rect 13225 4250 13260 4256
rect 13294 4250 13329 4256
rect 13363 4250 13398 4256
rect 12811 4222 12813 4250
rect 12880 4222 12886 4250
rect 12949 4222 12959 4250
rect 13018 4222 13032 4250
rect 13087 4222 13105 4250
rect 13156 4222 13178 4250
rect 13225 4222 13251 4250
rect 13294 4222 13324 4250
rect 13363 4222 13397 4250
rect 13432 4222 13467 4256
rect 13501 4250 13536 4256
rect 13570 4250 13605 4256
rect 13639 4250 13674 4256
rect 13708 4250 13743 4256
rect 13777 4250 13812 4256
rect 13846 4250 13881 4256
rect 13915 4250 13950 4256
rect 13984 4250 14019 4256
rect 13504 4222 13536 4250
rect 13577 4222 13605 4250
rect 13650 4222 13674 4250
rect 13723 4222 13743 4250
rect 13796 4222 13812 4250
rect 13869 4222 13881 4250
rect 13942 4222 13950 4250
rect 14015 4222 14019 4250
rect 14053 4250 14088 4256
rect 14053 4222 14054 4250
rect 11971 4216 12010 4222
rect 12044 4216 12083 4222
rect 12117 4216 12156 4222
rect 12190 4216 12229 4222
rect 12263 4216 12302 4222
rect 12336 4216 12375 4222
rect 12409 4216 12448 4222
rect 12482 4216 12521 4222
rect 12555 4216 12594 4222
rect 12628 4216 12667 4222
rect 12701 4216 12740 4222
rect 12774 4216 12813 4222
rect 12847 4216 12886 4222
rect 12920 4216 12959 4222
rect 12993 4216 13032 4222
rect 13066 4216 13105 4222
rect 13139 4216 13178 4222
rect 13212 4216 13251 4222
rect 13285 4216 13324 4222
rect 13358 4216 13397 4222
rect 13431 4216 13470 4222
rect 13504 4216 13543 4222
rect 13577 4216 13616 4222
rect 13650 4216 13689 4222
rect 13723 4216 13762 4222
rect 13796 4216 13835 4222
rect 13869 4216 13908 4222
rect 13942 4216 13981 4222
rect 14015 4216 14054 4222
rect 14122 4250 14157 4256
rect 14191 4250 14226 4256
rect 14260 4250 14295 4256
rect 14329 4250 14364 4256
rect 14398 4250 14433 4256
rect 14467 4250 14502 4256
rect 14536 4250 14571 4256
rect 14605 4250 14640 4256
rect 14122 4222 14127 4250
rect 14191 4222 14200 4250
rect 14260 4222 14273 4250
rect 14329 4222 14346 4250
rect 14398 4222 14419 4250
rect 14467 4222 14492 4250
rect 14536 4222 14565 4250
rect 14605 4222 14638 4250
rect 14674 4222 14709 4256
rect 14743 4250 14778 4256
rect 14812 4250 14847 4256
rect 14881 4250 14916 4256
rect 14950 4250 14985 4256
rect 15019 4250 15054 4256
rect 15088 4250 15123 4256
rect 15157 4250 15192 4256
rect 15226 4250 15261 4256
rect 14745 4222 14778 4250
rect 14818 4222 14847 4250
rect 14891 4222 14916 4250
rect 14964 4222 14985 4250
rect 15037 4222 15054 4250
rect 15110 4222 15123 4250
rect 15183 4222 15192 4250
rect 15256 4222 15261 4250
rect 15295 4250 15330 4256
rect 14088 4216 14127 4222
rect 14161 4216 14200 4222
rect 14234 4216 14273 4222
rect 14307 4216 14346 4222
rect 14380 4216 14419 4222
rect 14453 4216 14492 4222
rect 14526 4216 14565 4222
rect 14599 4216 14638 4222
rect 14672 4216 14711 4222
rect 14745 4216 14784 4222
rect 14818 4216 14857 4222
rect 14891 4216 14930 4222
rect 14964 4216 15003 4222
rect 15037 4216 15076 4222
rect 15110 4216 15149 4222
rect 15183 4216 15222 4222
rect 15256 4216 15295 4222
rect 15329 4222 15330 4250
rect 15364 4250 15399 4256
rect 15433 4250 15468 4256
rect 15502 4250 15537 4256
rect 15571 4250 15606 4256
rect 15640 4250 15675 4256
rect 15709 4250 15744 4256
rect 15778 4250 15813 4256
rect 15847 4250 15882 4256
rect 15364 4222 15368 4250
rect 15433 4222 15441 4250
rect 15502 4222 15514 4250
rect 15571 4222 15587 4250
rect 15640 4222 15660 4250
rect 15709 4222 15733 4250
rect 15778 4222 15806 4250
rect 15847 4222 15879 4250
rect 15916 4222 15951 4256
rect 15985 4250 16020 4256
rect 16054 4250 16089 4256
rect 16123 4250 16158 4256
rect 16192 4250 16227 4256
rect 16261 4250 16296 4256
rect 16330 4250 16365 4256
rect 15986 4222 16020 4250
rect 16059 4222 16089 4250
rect 16132 4222 16158 4250
rect 16205 4222 16227 4250
rect 16278 4222 16296 4250
rect 15329 4216 15368 4222
rect 15402 4216 15441 4222
rect 15475 4216 15514 4222
rect 15548 4216 15587 4222
rect 15621 4216 15660 4222
rect 15694 4216 15733 4222
rect 15767 4216 15806 4222
rect 15840 4216 15879 4222
rect 15913 4216 15952 4222
rect 15986 4216 16025 4222
rect 16059 4216 16098 4222
rect 16132 4216 16171 4222
rect 16205 4216 16244 4222
rect 16278 4216 16317 4222
rect 16351 4216 16365 4250
rect 11929 4188 16365 4216
rect 11929 4178 11949 4188
rect 11983 4178 12018 4188
rect 12052 4178 12087 4188
rect 11929 4144 11937 4178
rect 11983 4154 12010 4178
rect 12052 4154 12083 4178
rect 12121 4154 12156 4188
rect 12190 4154 12225 4188
rect 12259 4178 12294 4188
rect 12328 4178 12363 4188
rect 12397 4178 12432 4188
rect 12466 4178 12501 4188
rect 12535 4178 12570 4188
rect 12604 4178 12639 4188
rect 12673 4178 12708 4188
rect 12742 4178 12777 4188
rect 12263 4154 12294 4178
rect 12336 4154 12363 4178
rect 12409 4154 12432 4178
rect 12482 4154 12501 4178
rect 12555 4154 12570 4178
rect 12628 4154 12639 4178
rect 12701 4154 12708 4178
rect 12774 4154 12777 4178
rect 12811 4178 12846 4188
rect 12880 4178 12915 4188
rect 12949 4178 12984 4188
rect 13018 4178 13053 4188
rect 13087 4178 13122 4188
rect 13156 4178 13191 4188
rect 13225 4178 13260 4188
rect 13294 4178 13329 4188
rect 13363 4178 13398 4188
rect 12811 4154 12813 4178
rect 12880 4154 12886 4178
rect 12949 4154 12959 4178
rect 13018 4154 13032 4178
rect 13087 4154 13105 4178
rect 13156 4154 13178 4178
rect 13225 4154 13251 4178
rect 13294 4154 13324 4178
rect 13363 4154 13397 4178
rect 13432 4154 13467 4188
rect 13501 4178 13536 4188
rect 13570 4178 13605 4188
rect 13639 4178 13674 4188
rect 13708 4178 13743 4188
rect 13777 4178 13812 4188
rect 13846 4178 13881 4188
rect 13915 4178 13950 4188
rect 13984 4178 14019 4188
rect 13504 4154 13536 4178
rect 13577 4154 13605 4178
rect 13650 4154 13674 4178
rect 13723 4154 13743 4178
rect 13796 4154 13812 4178
rect 13869 4154 13881 4178
rect 13942 4154 13950 4178
rect 14015 4154 14019 4178
rect 14053 4178 14088 4188
rect 14053 4154 14054 4178
rect 11971 4144 12010 4154
rect 12044 4144 12083 4154
rect 12117 4144 12156 4154
rect 12190 4144 12229 4154
rect 12263 4144 12302 4154
rect 12336 4144 12375 4154
rect 12409 4144 12448 4154
rect 12482 4144 12521 4154
rect 12555 4144 12594 4154
rect 12628 4144 12667 4154
rect 12701 4144 12740 4154
rect 12774 4144 12813 4154
rect 12847 4144 12886 4154
rect 12920 4144 12959 4154
rect 12993 4144 13032 4154
rect 13066 4144 13105 4154
rect 13139 4144 13178 4154
rect 13212 4144 13251 4154
rect 13285 4144 13324 4154
rect 13358 4144 13397 4154
rect 13431 4144 13470 4154
rect 13504 4144 13543 4154
rect 13577 4144 13616 4154
rect 13650 4144 13689 4154
rect 13723 4144 13762 4154
rect 13796 4144 13835 4154
rect 13869 4144 13908 4154
rect 13942 4144 13981 4154
rect 14015 4144 14054 4154
rect 14122 4178 14157 4188
rect 14191 4178 14226 4188
rect 14260 4178 14295 4188
rect 14329 4178 14364 4188
rect 14398 4178 14433 4188
rect 14467 4178 14502 4188
rect 14536 4178 14571 4188
rect 14605 4178 14640 4188
rect 14122 4154 14127 4178
rect 14191 4154 14200 4178
rect 14260 4154 14273 4178
rect 14329 4154 14346 4178
rect 14398 4154 14419 4178
rect 14467 4154 14492 4178
rect 14536 4154 14565 4178
rect 14605 4154 14638 4178
rect 14674 4154 14709 4188
rect 14743 4178 14778 4188
rect 14812 4178 14847 4188
rect 14881 4178 14916 4188
rect 14950 4178 14985 4188
rect 15019 4178 15054 4188
rect 15088 4178 15123 4188
rect 15157 4178 15192 4188
rect 15226 4178 15261 4188
rect 14745 4154 14778 4178
rect 14818 4154 14847 4178
rect 14891 4154 14916 4178
rect 14964 4154 14985 4178
rect 15037 4154 15054 4178
rect 15110 4154 15123 4178
rect 15183 4154 15192 4178
rect 15256 4154 15261 4178
rect 15295 4178 15330 4188
rect 14088 4144 14127 4154
rect 14161 4144 14200 4154
rect 14234 4144 14273 4154
rect 14307 4144 14346 4154
rect 14380 4144 14419 4154
rect 14453 4144 14492 4154
rect 14526 4144 14565 4154
rect 14599 4144 14638 4154
rect 14672 4144 14711 4154
rect 14745 4144 14784 4154
rect 14818 4144 14857 4154
rect 14891 4144 14930 4154
rect 14964 4144 15003 4154
rect 15037 4144 15076 4154
rect 15110 4144 15149 4154
rect 15183 4144 15222 4154
rect 15256 4144 15295 4154
rect 15329 4154 15330 4178
rect 15364 4178 15399 4188
rect 15433 4178 15468 4188
rect 15502 4178 15537 4188
rect 15571 4178 15606 4188
rect 15640 4178 15675 4188
rect 15709 4178 15744 4188
rect 15778 4178 15813 4188
rect 15847 4178 15882 4188
rect 15364 4154 15368 4178
rect 15433 4154 15441 4178
rect 15502 4154 15514 4178
rect 15571 4154 15587 4178
rect 15640 4154 15660 4178
rect 15709 4154 15733 4178
rect 15778 4154 15806 4178
rect 15847 4154 15879 4178
rect 15916 4154 15951 4188
rect 15985 4178 16020 4188
rect 16054 4178 16089 4188
rect 16123 4178 16158 4188
rect 16192 4178 16227 4188
rect 16261 4178 16296 4188
rect 16330 4178 16365 4188
rect 15986 4154 16020 4178
rect 16059 4154 16089 4178
rect 16132 4154 16158 4178
rect 16205 4154 16227 4178
rect 16278 4154 16296 4178
rect 15329 4144 15368 4154
rect 15402 4144 15441 4154
rect 15475 4144 15514 4154
rect 15548 4144 15587 4154
rect 15621 4144 15660 4154
rect 15694 4144 15733 4154
rect 15767 4144 15806 4154
rect 15840 4144 15879 4154
rect 15913 4144 15952 4154
rect 15986 4144 16025 4154
rect 16059 4144 16098 4154
rect 16132 4144 16171 4154
rect 16205 4144 16244 4154
rect 16278 4144 16317 4154
rect 16351 4144 16365 4178
rect 11929 4120 16365 4144
rect 11929 4106 11949 4120
rect 11983 4106 12018 4120
rect 12052 4106 12087 4120
rect 11929 4072 11937 4106
rect 11983 4086 12010 4106
rect 12052 4086 12083 4106
rect 12121 4086 12156 4120
rect 12190 4086 12225 4120
rect 12259 4106 12294 4120
rect 12328 4106 12363 4120
rect 12397 4106 12432 4120
rect 12466 4106 12501 4120
rect 12535 4106 12570 4120
rect 12604 4106 12639 4120
rect 12673 4106 12708 4120
rect 12742 4106 12777 4120
rect 12263 4086 12294 4106
rect 12336 4086 12363 4106
rect 12409 4086 12432 4106
rect 12482 4086 12501 4106
rect 12555 4086 12570 4106
rect 12628 4086 12639 4106
rect 12701 4086 12708 4106
rect 12774 4086 12777 4106
rect 12811 4106 12846 4120
rect 12880 4106 12915 4120
rect 12949 4106 12984 4120
rect 13018 4106 13053 4120
rect 13087 4106 13122 4120
rect 13156 4106 13191 4120
rect 13225 4106 13260 4120
rect 13294 4106 13329 4120
rect 13363 4106 13398 4120
rect 12811 4086 12813 4106
rect 12880 4086 12886 4106
rect 12949 4086 12959 4106
rect 13018 4086 13032 4106
rect 13087 4086 13105 4106
rect 13156 4086 13178 4106
rect 13225 4086 13251 4106
rect 13294 4086 13324 4106
rect 13363 4086 13397 4106
rect 13432 4086 13467 4120
rect 13501 4106 13536 4120
rect 13570 4106 13605 4120
rect 13639 4106 13674 4120
rect 13708 4106 13743 4120
rect 13777 4106 13812 4120
rect 13846 4106 13881 4120
rect 13915 4106 13950 4120
rect 13984 4106 14019 4120
rect 13504 4086 13536 4106
rect 13577 4086 13605 4106
rect 13650 4086 13674 4106
rect 13723 4086 13743 4106
rect 13796 4086 13812 4106
rect 13869 4086 13881 4106
rect 13942 4086 13950 4106
rect 14015 4086 14019 4106
rect 14053 4106 14088 4120
rect 14053 4086 14054 4106
rect 11971 4072 12010 4086
rect 12044 4072 12083 4086
rect 12117 4072 12156 4086
rect 12190 4072 12229 4086
rect 12263 4072 12302 4086
rect 12336 4072 12375 4086
rect 12409 4072 12448 4086
rect 12482 4072 12521 4086
rect 12555 4072 12594 4086
rect 12628 4072 12667 4086
rect 12701 4072 12740 4086
rect 12774 4072 12813 4086
rect 12847 4072 12886 4086
rect 12920 4072 12959 4086
rect 12993 4072 13032 4086
rect 13066 4072 13105 4086
rect 13139 4072 13178 4086
rect 13212 4072 13251 4086
rect 13285 4072 13324 4086
rect 13358 4072 13397 4086
rect 13431 4072 13470 4086
rect 13504 4072 13543 4086
rect 13577 4072 13616 4086
rect 13650 4072 13689 4086
rect 13723 4072 13762 4086
rect 13796 4072 13835 4086
rect 13869 4072 13908 4086
rect 13942 4072 13981 4086
rect 14015 4072 14054 4086
rect 14122 4106 14157 4120
rect 14191 4106 14226 4120
rect 14260 4106 14295 4120
rect 14329 4106 14364 4120
rect 14398 4106 14433 4120
rect 14467 4106 14502 4120
rect 14536 4106 14571 4120
rect 14605 4106 14640 4120
rect 14122 4086 14127 4106
rect 14191 4086 14200 4106
rect 14260 4086 14273 4106
rect 14329 4086 14346 4106
rect 14398 4086 14419 4106
rect 14467 4086 14492 4106
rect 14536 4086 14565 4106
rect 14605 4086 14638 4106
rect 14674 4086 14709 4120
rect 14743 4106 14778 4120
rect 14812 4106 14847 4120
rect 14881 4106 14916 4120
rect 14950 4106 14985 4120
rect 15019 4106 15054 4120
rect 15088 4106 15123 4120
rect 15157 4106 15192 4120
rect 15226 4106 15261 4120
rect 14745 4086 14778 4106
rect 14818 4086 14847 4106
rect 14891 4086 14916 4106
rect 14964 4086 14985 4106
rect 15037 4086 15054 4106
rect 15110 4086 15123 4106
rect 15183 4086 15192 4106
rect 15256 4086 15261 4106
rect 15295 4106 15330 4120
rect 14088 4072 14127 4086
rect 14161 4072 14200 4086
rect 14234 4072 14273 4086
rect 14307 4072 14346 4086
rect 14380 4072 14419 4086
rect 14453 4072 14492 4086
rect 14526 4072 14565 4086
rect 14599 4072 14638 4086
rect 14672 4072 14711 4086
rect 14745 4072 14784 4086
rect 14818 4072 14857 4086
rect 14891 4072 14930 4086
rect 14964 4072 15003 4086
rect 15037 4072 15076 4086
rect 15110 4072 15149 4086
rect 15183 4072 15222 4086
rect 15256 4072 15295 4086
rect 15329 4086 15330 4106
rect 15364 4106 15399 4120
rect 15433 4106 15468 4120
rect 15502 4106 15537 4120
rect 15571 4106 15606 4120
rect 15640 4106 15675 4120
rect 15709 4106 15744 4120
rect 15778 4106 15813 4120
rect 15847 4106 15882 4120
rect 15364 4086 15368 4106
rect 15433 4086 15441 4106
rect 15502 4086 15514 4106
rect 15571 4086 15587 4106
rect 15640 4086 15660 4106
rect 15709 4086 15733 4106
rect 15778 4086 15806 4106
rect 15847 4086 15879 4106
rect 15916 4086 15951 4120
rect 15985 4106 16020 4120
rect 16054 4106 16089 4120
rect 16123 4106 16158 4120
rect 16192 4106 16227 4120
rect 16261 4106 16296 4120
rect 16330 4106 16365 4120
rect 15986 4086 16020 4106
rect 16059 4086 16089 4106
rect 16132 4086 16158 4106
rect 16205 4086 16227 4106
rect 16278 4086 16296 4106
rect 15329 4072 15368 4086
rect 15402 4072 15441 4086
rect 15475 4072 15514 4086
rect 15548 4072 15587 4086
rect 15621 4072 15660 4086
rect 15694 4072 15733 4086
rect 15767 4072 15806 4086
rect 15840 4072 15879 4086
rect 15913 4072 15952 4086
rect 15986 4072 16025 4086
rect 16059 4072 16098 4086
rect 16132 4072 16171 4086
rect 16205 4072 16244 4086
rect 16278 4072 16317 4086
rect 16351 4072 16365 4106
rect 11929 4052 16365 4072
rect 11929 4034 11949 4052
rect 11983 4034 12018 4052
rect 12052 4034 12087 4052
rect 11929 4000 11937 4034
rect 11983 4018 12010 4034
rect 12052 4018 12083 4034
rect 12121 4018 12156 4052
rect 12190 4018 12225 4052
rect 12259 4034 12294 4052
rect 12328 4034 12363 4052
rect 12397 4034 12432 4052
rect 12466 4034 12501 4052
rect 12535 4034 12570 4052
rect 12604 4034 12639 4052
rect 12673 4034 12708 4052
rect 12742 4034 12777 4052
rect 12263 4018 12294 4034
rect 12336 4018 12363 4034
rect 12409 4018 12432 4034
rect 12482 4018 12501 4034
rect 12555 4018 12570 4034
rect 12628 4018 12639 4034
rect 12701 4018 12708 4034
rect 12774 4018 12777 4034
rect 12811 4034 12846 4052
rect 12880 4034 12915 4052
rect 12949 4034 12984 4052
rect 13018 4034 13053 4052
rect 13087 4034 13122 4052
rect 13156 4034 13191 4052
rect 13225 4034 13260 4052
rect 13294 4034 13329 4052
rect 13363 4034 13398 4052
rect 12811 4018 12813 4034
rect 12880 4018 12886 4034
rect 12949 4018 12959 4034
rect 13018 4018 13032 4034
rect 13087 4018 13105 4034
rect 13156 4018 13178 4034
rect 13225 4018 13251 4034
rect 13294 4018 13324 4034
rect 13363 4018 13397 4034
rect 13432 4018 13467 4052
rect 13501 4034 13536 4052
rect 13570 4034 13605 4052
rect 13639 4034 13674 4052
rect 13708 4034 13743 4052
rect 13777 4034 13812 4052
rect 13846 4034 13881 4052
rect 13915 4034 13950 4052
rect 13984 4034 14019 4052
rect 13504 4018 13536 4034
rect 13577 4018 13605 4034
rect 13650 4018 13674 4034
rect 13723 4018 13743 4034
rect 13796 4018 13812 4034
rect 13869 4018 13881 4034
rect 13942 4018 13950 4034
rect 14015 4018 14019 4034
rect 14053 4034 14088 4052
rect 14053 4018 14054 4034
rect 11971 4000 12010 4018
rect 12044 4000 12083 4018
rect 12117 4000 12156 4018
rect 12190 4000 12229 4018
rect 12263 4000 12302 4018
rect 12336 4000 12375 4018
rect 12409 4000 12448 4018
rect 12482 4000 12521 4018
rect 12555 4000 12594 4018
rect 12628 4000 12667 4018
rect 12701 4000 12740 4018
rect 12774 4000 12813 4018
rect 12847 4000 12886 4018
rect 12920 4000 12959 4018
rect 12993 4000 13032 4018
rect 13066 4000 13105 4018
rect 13139 4000 13178 4018
rect 13212 4000 13251 4018
rect 13285 4000 13324 4018
rect 13358 4000 13397 4018
rect 13431 4000 13470 4018
rect 13504 4000 13543 4018
rect 13577 4000 13616 4018
rect 13650 4000 13689 4018
rect 13723 4000 13762 4018
rect 13796 4000 13835 4018
rect 13869 4000 13908 4018
rect 13942 4000 13981 4018
rect 14015 4000 14054 4018
rect 14122 4034 14157 4052
rect 14191 4034 14226 4052
rect 14260 4034 14295 4052
rect 14329 4034 14364 4052
rect 14398 4034 14433 4052
rect 14467 4034 14502 4052
rect 14536 4034 14571 4052
rect 14605 4034 14640 4052
rect 14122 4018 14127 4034
rect 14191 4018 14200 4034
rect 14260 4018 14273 4034
rect 14329 4018 14346 4034
rect 14398 4018 14419 4034
rect 14467 4018 14492 4034
rect 14536 4018 14565 4034
rect 14605 4018 14638 4034
rect 14674 4018 14709 4052
rect 14743 4034 14778 4052
rect 14812 4034 14847 4052
rect 14881 4034 14916 4052
rect 14950 4034 14985 4052
rect 15019 4034 15054 4052
rect 15088 4034 15123 4052
rect 15157 4034 15192 4052
rect 15226 4034 15261 4052
rect 14745 4018 14778 4034
rect 14818 4018 14847 4034
rect 14891 4018 14916 4034
rect 14964 4018 14985 4034
rect 15037 4018 15054 4034
rect 15110 4018 15123 4034
rect 15183 4018 15192 4034
rect 15256 4018 15261 4034
rect 15295 4034 15330 4052
rect 14088 4000 14127 4018
rect 14161 4000 14200 4018
rect 14234 4000 14273 4018
rect 14307 4000 14346 4018
rect 14380 4000 14419 4018
rect 14453 4000 14492 4018
rect 14526 4000 14565 4018
rect 14599 4000 14638 4018
rect 14672 4000 14711 4018
rect 14745 4000 14784 4018
rect 14818 4000 14857 4018
rect 14891 4000 14930 4018
rect 14964 4000 15003 4018
rect 15037 4000 15076 4018
rect 15110 4000 15149 4018
rect 15183 4000 15222 4018
rect 15256 4000 15295 4018
rect 15329 4018 15330 4034
rect 15364 4034 15399 4052
rect 15433 4034 15468 4052
rect 15502 4034 15537 4052
rect 15571 4034 15606 4052
rect 15640 4034 15675 4052
rect 15709 4034 15744 4052
rect 15778 4034 15813 4052
rect 15847 4034 15882 4052
rect 15364 4018 15368 4034
rect 15433 4018 15441 4034
rect 15502 4018 15514 4034
rect 15571 4018 15587 4034
rect 15640 4018 15660 4034
rect 15709 4018 15733 4034
rect 15778 4018 15806 4034
rect 15847 4018 15879 4034
rect 15916 4018 15951 4052
rect 15985 4034 16020 4052
rect 16054 4034 16089 4052
rect 16123 4034 16158 4052
rect 16192 4034 16227 4052
rect 16261 4034 16296 4052
rect 16330 4034 16365 4052
rect 15986 4018 16020 4034
rect 16059 4018 16089 4034
rect 16132 4018 16158 4034
rect 16205 4018 16227 4034
rect 16278 4018 16296 4034
rect 15329 4000 15368 4018
rect 15402 4000 15441 4018
rect 15475 4000 15514 4018
rect 15548 4000 15587 4018
rect 15621 4000 15660 4018
rect 15694 4000 15733 4018
rect 15767 4000 15806 4018
rect 15840 4000 15879 4018
rect 15913 4000 15952 4018
rect 15986 4000 16025 4018
rect 16059 4000 16098 4018
rect 16132 4000 16171 4018
rect 16205 4000 16244 4018
rect 16278 4000 16317 4018
rect 16351 4000 16365 4034
rect 11929 3984 16365 4000
rect 11929 3962 11949 3984
rect 11983 3962 12018 3984
rect 12052 3962 12087 3984
rect 11929 3928 11937 3962
rect 11983 3950 12010 3962
rect 12052 3950 12083 3962
rect 12121 3950 12156 3984
rect 12190 3950 12225 3984
rect 12259 3962 12294 3984
rect 12328 3962 12363 3984
rect 12397 3962 12432 3984
rect 12466 3962 12501 3984
rect 12535 3962 12570 3984
rect 12604 3962 12639 3984
rect 12673 3962 12708 3984
rect 12742 3962 12777 3984
rect 12263 3950 12294 3962
rect 12336 3950 12363 3962
rect 12409 3950 12432 3962
rect 12482 3950 12501 3962
rect 12555 3950 12570 3962
rect 12628 3950 12639 3962
rect 12701 3950 12708 3962
rect 12774 3950 12777 3962
rect 12811 3962 12846 3984
rect 12880 3962 12915 3984
rect 12949 3962 12984 3984
rect 13018 3962 13053 3984
rect 13087 3962 13122 3984
rect 13156 3962 13191 3984
rect 13225 3962 13260 3984
rect 13294 3962 13329 3984
rect 13363 3962 13398 3984
rect 12811 3950 12813 3962
rect 12880 3950 12886 3962
rect 12949 3950 12959 3962
rect 13018 3950 13032 3962
rect 13087 3950 13105 3962
rect 13156 3950 13178 3962
rect 13225 3950 13251 3962
rect 13294 3950 13324 3962
rect 13363 3950 13397 3962
rect 13432 3950 13467 3984
rect 13501 3962 13536 3984
rect 13570 3962 13605 3984
rect 13639 3962 13674 3984
rect 13708 3962 13743 3984
rect 13777 3962 13812 3984
rect 13846 3962 13881 3984
rect 13915 3962 13950 3984
rect 13984 3962 14019 3984
rect 13504 3950 13536 3962
rect 13577 3950 13605 3962
rect 13650 3950 13674 3962
rect 13723 3950 13743 3962
rect 13796 3950 13812 3962
rect 13869 3950 13881 3962
rect 13942 3950 13950 3962
rect 14015 3950 14019 3962
rect 14053 3962 14088 3984
rect 14053 3950 14054 3962
rect 11971 3928 12010 3950
rect 12044 3928 12083 3950
rect 12117 3928 12156 3950
rect 12190 3928 12229 3950
rect 12263 3928 12302 3950
rect 12336 3928 12375 3950
rect 12409 3928 12448 3950
rect 12482 3928 12521 3950
rect 12555 3928 12594 3950
rect 12628 3928 12667 3950
rect 12701 3928 12740 3950
rect 12774 3928 12813 3950
rect 12847 3928 12886 3950
rect 12920 3928 12959 3950
rect 12993 3928 13032 3950
rect 13066 3928 13105 3950
rect 13139 3928 13178 3950
rect 13212 3928 13251 3950
rect 13285 3928 13324 3950
rect 13358 3928 13397 3950
rect 13431 3928 13470 3950
rect 13504 3928 13543 3950
rect 13577 3928 13616 3950
rect 13650 3928 13689 3950
rect 13723 3928 13762 3950
rect 13796 3928 13835 3950
rect 13869 3928 13908 3950
rect 13942 3928 13981 3950
rect 14015 3928 14054 3950
rect 14122 3962 14157 3984
rect 14191 3962 14226 3984
rect 14260 3962 14295 3984
rect 14329 3962 14364 3984
rect 14398 3962 14433 3984
rect 14467 3962 14502 3984
rect 14536 3962 14571 3984
rect 14605 3962 14640 3984
rect 14122 3950 14127 3962
rect 14191 3950 14200 3962
rect 14260 3950 14273 3962
rect 14329 3950 14346 3962
rect 14398 3950 14419 3962
rect 14467 3950 14492 3962
rect 14536 3950 14565 3962
rect 14605 3950 14638 3962
rect 14674 3950 14709 3984
rect 14743 3962 14778 3984
rect 14812 3962 14847 3984
rect 14881 3962 14916 3984
rect 14950 3962 14985 3984
rect 15019 3962 15054 3984
rect 15088 3962 15123 3984
rect 15157 3962 15192 3984
rect 15226 3962 15261 3984
rect 14745 3950 14778 3962
rect 14818 3950 14847 3962
rect 14891 3950 14916 3962
rect 14964 3950 14985 3962
rect 15037 3950 15054 3962
rect 15110 3950 15123 3962
rect 15183 3950 15192 3962
rect 15256 3950 15261 3962
rect 15295 3962 15330 3984
rect 14088 3928 14127 3950
rect 14161 3928 14200 3950
rect 14234 3928 14273 3950
rect 14307 3928 14346 3950
rect 14380 3928 14419 3950
rect 14453 3928 14492 3950
rect 14526 3928 14565 3950
rect 14599 3928 14638 3950
rect 14672 3928 14711 3950
rect 14745 3928 14784 3950
rect 14818 3928 14857 3950
rect 14891 3928 14930 3950
rect 14964 3928 15003 3950
rect 15037 3928 15076 3950
rect 15110 3928 15149 3950
rect 15183 3928 15222 3950
rect 15256 3928 15295 3950
rect 15329 3950 15330 3962
rect 15364 3962 15399 3984
rect 15433 3962 15468 3984
rect 15502 3962 15537 3984
rect 15571 3962 15606 3984
rect 15640 3962 15675 3984
rect 15709 3962 15744 3984
rect 15778 3962 15813 3984
rect 15847 3962 15882 3984
rect 15364 3950 15368 3962
rect 15433 3950 15441 3962
rect 15502 3950 15514 3962
rect 15571 3950 15587 3962
rect 15640 3950 15660 3962
rect 15709 3950 15733 3962
rect 15778 3950 15806 3962
rect 15847 3950 15879 3962
rect 15916 3950 15951 3984
rect 15985 3962 16020 3984
rect 16054 3962 16089 3984
rect 16123 3962 16158 3984
rect 16192 3962 16227 3984
rect 16261 3962 16296 3984
rect 16330 3962 16365 3984
rect 15986 3950 16020 3962
rect 16059 3950 16089 3962
rect 16132 3950 16158 3962
rect 16205 3950 16227 3962
rect 16278 3950 16296 3962
rect 15329 3928 15368 3950
rect 15402 3928 15441 3950
rect 15475 3928 15514 3950
rect 15548 3928 15587 3950
rect 15621 3928 15660 3950
rect 15694 3928 15733 3950
rect 15767 3928 15806 3950
rect 15840 3928 15879 3950
rect 15913 3928 15952 3950
rect 15986 3928 16025 3950
rect 16059 3928 16098 3950
rect 16132 3928 16171 3950
rect 16205 3928 16244 3950
rect 16278 3928 16317 3950
rect 16351 3928 16365 3962
rect 11929 3916 16365 3928
rect 11929 3890 11949 3916
rect 11983 3890 12018 3916
rect 12052 3890 12087 3916
rect 11929 3856 11937 3890
rect 11983 3882 12010 3890
rect 12052 3882 12083 3890
rect 12121 3882 12156 3916
rect 12190 3882 12225 3916
rect 12259 3890 12294 3916
rect 12328 3890 12363 3916
rect 12397 3890 12432 3916
rect 12466 3890 12501 3916
rect 12535 3890 12570 3916
rect 12604 3890 12639 3916
rect 12673 3890 12708 3916
rect 12742 3890 12777 3916
rect 12263 3882 12294 3890
rect 12336 3882 12363 3890
rect 12409 3882 12432 3890
rect 12482 3882 12501 3890
rect 12555 3882 12570 3890
rect 12628 3882 12639 3890
rect 12701 3882 12708 3890
rect 12774 3882 12777 3890
rect 12811 3890 12846 3916
rect 12880 3890 12915 3916
rect 12949 3890 12984 3916
rect 13018 3890 13053 3916
rect 13087 3890 13122 3916
rect 13156 3890 13191 3916
rect 13225 3890 13260 3916
rect 13294 3890 13329 3916
rect 13363 3890 13398 3916
rect 12811 3882 12813 3890
rect 12880 3882 12886 3890
rect 12949 3882 12959 3890
rect 13018 3882 13032 3890
rect 13087 3882 13105 3890
rect 13156 3882 13178 3890
rect 13225 3882 13251 3890
rect 13294 3882 13324 3890
rect 13363 3882 13397 3890
rect 13432 3882 13467 3916
rect 13501 3890 13536 3916
rect 13570 3890 13605 3916
rect 13639 3890 13674 3916
rect 13708 3890 13743 3916
rect 13777 3890 13812 3916
rect 13846 3890 13881 3916
rect 13915 3890 13950 3916
rect 13984 3890 14019 3916
rect 13504 3882 13536 3890
rect 13577 3882 13605 3890
rect 13650 3882 13674 3890
rect 13723 3882 13743 3890
rect 13796 3882 13812 3890
rect 13869 3882 13881 3890
rect 13942 3882 13950 3890
rect 14015 3882 14019 3890
rect 14053 3890 14088 3916
rect 14053 3882 14054 3890
rect 11971 3856 12010 3882
rect 12044 3856 12083 3882
rect 12117 3856 12156 3882
rect 12190 3856 12229 3882
rect 12263 3856 12302 3882
rect 12336 3856 12375 3882
rect 12409 3856 12448 3882
rect 12482 3856 12521 3882
rect 12555 3856 12594 3882
rect 12628 3856 12667 3882
rect 12701 3856 12740 3882
rect 12774 3856 12813 3882
rect 12847 3856 12886 3882
rect 12920 3856 12959 3882
rect 12993 3856 13032 3882
rect 13066 3856 13105 3882
rect 13139 3856 13178 3882
rect 13212 3856 13251 3882
rect 13285 3856 13324 3882
rect 13358 3856 13397 3882
rect 13431 3856 13470 3882
rect 13504 3856 13543 3882
rect 13577 3856 13616 3882
rect 13650 3856 13689 3882
rect 13723 3856 13762 3882
rect 13796 3856 13835 3882
rect 13869 3856 13908 3882
rect 13942 3856 13981 3882
rect 14015 3856 14054 3882
rect 14122 3890 14157 3916
rect 14191 3890 14226 3916
rect 14260 3890 14295 3916
rect 14329 3890 14364 3916
rect 14398 3890 14433 3916
rect 14467 3890 14502 3916
rect 14536 3890 14571 3916
rect 14605 3890 14640 3916
rect 14122 3882 14127 3890
rect 14191 3882 14200 3890
rect 14260 3882 14273 3890
rect 14329 3882 14346 3890
rect 14398 3882 14419 3890
rect 14467 3882 14492 3890
rect 14536 3882 14565 3890
rect 14605 3882 14638 3890
rect 14674 3882 14709 3916
rect 14743 3890 14778 3916
rect 14812 3890 14847 3916
rect 14881 3890 14916 3916
rect 14950 3890 14985 3916
rect 15019 3890 15054 3916
rect 15088 3890 15123 3916
rect 15157 3890 15192 3916
rect 15226 3890 15261 3916
rect 14745 3882 14778 3890
rect 14818 3882 14847 3890
rect 14891 3882 14916 3890
rect 14964 3882 14985 3890
rect 15037 3882 15054 3890
rect 15110 3882 15123 3890
rect 15183 3882 15192 3890
rect 15256 3882 15261 3890
rect 15295 3890 15330 3916
rect 14088 3856 14127 3882
rect 14161 3856 14200 3882
rect 14234 3856 14273 3882
rect 14307 3856 14346 3882
rect 14380 3856 14419 3882
rect 14453 3856 14492 3882
rect 14526 3856 14565 3882
rect 14599 3856 14638 3882
rect 14672 3856 14711 3882
rect 14745 3856 14784 3882
rect 14818 3856 14857 3882
rect 14891 3856 14930 3882
rect 14964 3856 15003 3882
rect 15037 3856 15076 3882
rect 15110 3856 15149 3882
rect 15183 3856 15222 3882
rect 15256 3856 15295 3882
rect 15329 3882 15330 3890
rect 15364 3890 15399 3916
rect 15433 3890 15468 3916
rect 15502 3890 15537 3916
rect 15571 3890 15606 3916
rect 15640 3890 15675 3916
rect 15709 3890 15744 3916
rect 15778 3890 15813 3916
rect 15847 3890 15882 3916
rect 15364 3882 15368 3890
rect 15433 3882 15441 3890
rect 15502 3882 15514 3890
rect 15571 3882 15587 3890
rect 15640 3882 15660 3890
rect 15709 3882 15733 3890
rect 15778 3882 15806 3890
rect 15847 3882 15879 3890
rect 15916 3882 15951 3916
rect 15985 3890 16020 3916
rect 16054 3890 16089 3916
rect 16123 3890 16158 3916
rect 16192 3890 16227 3916
rect 16261 3890 16296 3916
rect 16330 3890 16365 3916
rect 15986 3882 16020 3890
rect 16059 3882 16089 3890
rect 16132 3882 16158 3890
rect 16205 3882 16227 3890
rect 16278 3882 16296 3890
rect 15329 3856 15368 3882
rect 15402 3856 15441 3882
rect 15475 3856 15514 3882
rect 15548 3856 15587 3882
rect 15621 3856 15660 3882
rect 15694 3856 15733 3882
rect 15767 3856 15806 3882
rect 15840 3856 15879 3882
rect 15913 3856 15952 3882
rect 15986 3856 16025 3882
rect 16059 3856 16098 3882
rect 16132 3856 16171 3882
rect 16205 3856 16244 3882
rect 16278 3856 16317 3882
rect 16351 3856 16365 3890
rect 11929 3848 16365 3856
rect 11929 3814 11949 3848
rect 11983 3814 12018 3848
rect 12052 3814 12087 3848
rect 12121 3814 12156 3848
rect 12190 3814 12225 3848
rect 12259 3814 12294 3848
rect 12328 3814 12363 3848
rect 12397 3814 12432 3848
rect 12466 3814 12501 3848
rect 12535 3814 12570 3848
rect 12604 3814 12639 3848
rect 12673 3814 12708 3848
rect 12742 3814 12777 3848
rect 12811 3814 12846 3848
rect 12880 3814 12915 3848
rect 12949 3814 12984 3848
rect 13018 3814 13053 3848
rect 13087 3814 13122 3848
rect 13156 3814 13191 3848
rect 13225 3814 13260 3848
rect 13294 3814 13329 3848
rect 13363 3814 13398 3848
rect 13432 3814 13467 3848
rect 13501 3814 13536 3848
rect 13570 3814 13605 3848
rect 13639 3814 13674 3848
rect 13708 3814 13743 3848
rect 13777 3814 13812 3848
rect 13846 3814 13881 3848
rect 13915 3814 13950 3848
rect 13984 3814 14019 3848
rect 14053 3814 14088 3848
rect 14122 3814 14157 3848
rect 14191 3814 14226 3848
rect 14260 3814 14295 3848
rect 14329 3814 14364 3848
rect 14398 3814 14433 3848
rect 14467 3814 14502 3848
rect 14536 3814 14571 3848
rect 14605 3814 14640 3848
rect 14674 3814 14709 3848
rect 14743 3814 14778 3848
rect 14812 3814 14847 3848
rect 14881 3814 14916 3848
rect 14950 3814 14985 3848
rect 15019 3814 15054 3848
rect 15088 3814 15123 3848
rect 15157 3814 15192 3848
rect 15226 3814 15261 3848
rect 15295 3814 15330 3848
rect 15364 3814 15399 3848
rect 15433 3814 15468 3848
rect 15502 3814 15537 3848
rect 15571 3814 15606 3848
rect 15640 3814 15675 3848
rect 15709 3814 15744 3848
rect 15778 3814 15813 3848
rect 15847 3814 15882 3848
rect 15916 3814 15951 3848
rect 15985 3814 16020 3848
rect 16054 3814 16089 3848
rect 16123 3814 16158 3848
rect 16192 3814 16227 3848
rect 16261 3814 16296 3848
rect 16330 3814 16365 3848
rect 11929 3780 16365 3814
rect 11929 3746 11949 3780
rect 11983 3746 12018 3780
rect 12052 3746 12087 3780
rect 12121 3746 12156 3780
rect 12190 3746 12225 3780
rect 12259 3746 12294 3780
rect 12328 3746 12363 3780
rect 12397 3746 12432 3780
rect 12466 3746 12501 3780
rect 12535 3746 12570 3780
rect 12604 3746 12639 3780
rect 12673 3746 12708 3780
rect 12742 3746 12777 3780
rect 12811 3746 12846 3780
rect 12880 3746 12915 3780
rect 12949 3746 12984 3780
rect 13018 3746 13053 3780
rect 13087 3746 13122 3780
rect 13156 3746 13191 3780
rect 13225 3746 13260 3780
rect 13294 3746 13329 3780
rect 13363 3746 13398 3780
rect 13432 3746 13467 3780
rect 13501 3746 13536 3780
rect 13570 3746 13605 3780
rect 13639 3746 13674 3780
rect 13708 3746 13743 3780
rect 13777 3746 13812 3780
rect 13846 3746 13881 3780
rect 13915 3746 13950 3780
rect 13984 3746 14019 3780
rect 14053 3746 14088 3780
rect 14122 3746 14157 3780
rect 14191 3746 14226 3780
rect 14260 3746 14295 3780
rect 14329 3746 14364 3780
rect 14398 3746 14433 3780
rect 14467 3746 14502 3780
rect 14536 3746 14571 3780
rect 14605 3746 14640 3780
rect 14674 3746 14709 3780
rect 14743 3746 14778 3780
rect 14812 3746 14847 3780
rect 14881 3746 14916 3780
rect 14950 3746 14985 3780
rect 15019 3746 15054 3780
rect 15088 3746 15123 3780
rect 15157 3746 15192 3780
rect 15226 3746 15261 3780
rect 15295 3746 15330 3780
rect 15364 3746 15399 3780
rect 15433 3746 15468 3780
rect 15502 3746 15537 3780
rect 15571 3746 15606 3780
rect 15640 3746 15675 3780
rect 15709 3746 15744 3780
rect 15778 3746 15813 3780
rect 15847 3746 15882 3780
rect 15916 3746 15951 3780
rect 15985 3746 16020 3780
rect 16054 3746 16089 3780
rect 16123 3746 16158 3780
rect 16192 3746 16227 3780
rect 16261 3746 16296 3780
rect 16330 3746 16365 3780
rect 11929 3712 16365 3746
rect 11929 3678 11949 3712
rect 11983 3678 12018 3712
rect 12052 3678 12087 3712
rect 12121 3678 12156 3712
rect 12190 3678 12225 3712
rect 12259 3678 12294 3712
rect 12328 3678 12363 3712
rect 12397 3678 12432 3712
rect 12466 3678 12501 3712
rect 12535 3678 12570 3712
rect 12604 3678 12639 3712
rect 12673 3678 12708 3712
rect 12742 3678 12777 3712
rect 12811 3678 12846 3712
rect 12880 3678 12915 3712
rect 12949 3678 12984 3712
rect 13018 3678 13053 3712
rect 13087 3678 13122 3712
rect 13156 3678 13191 3712
rect 13225 3678 13260 3712
rect 13294 3678 13329 3712
rect 13363 3678 13398 3712
rect 13432 3678 13467 3712
rect 13501 3678 13536 3712
rect 13570 3678 13605 3712
rect 13639 3678 13674 3712
rect 13708 3678 13743 3712
rect 13777 3678 13812 3712
rect 13846 3678 13881 3712
rect 13915 3678 13950 3712
rect 13984 3678 14019 3712
rect 14053 3678 14088 3712
rect 14122 3678 14157 3712
rect 14191 3678 14226 3712
rect 14260 3678 14295 3712
rect 14329 3678 14364 3712
rect 14398 3678 14433 3712
rect 14467 3678 14502 3712
rect 14536 3678 14571 3712
rect 14605 3678 14640 3712
rect 14674 3678 14709 3712
rect 14743 3678 14778 3712
rect 14812 3678 14847 3712
rect 14881 3678 14916 3712
rect 14950 3678 14985 3712
rect 15019 3678 15054 3712
rect 15088 3678 15123 3712
rect 15157 3678 15192 3712
rect 15226 3678 15261 3712
rect 15295 3678 15330 3712
rect 15364 3678 15399 3712
rect 15433 3678 15468 3712
rect 15502 3678 15537 3712
rect 15571 3678 15606 3712
rect 15640 3678 15675 3712
rect 15709 3678 15744 3712
rect 15778 3678 15813 3712
rect 15847 3678 15882 3712
rect 15916 3678 15951 3712
rect 15985 3678 16020 3712
rect 16054 3678 16089 3712
rect 16123 3678 16158 3712
rect 16192 3678 16227 3712
rect 16261 3678 16296 3712
rect 16330 3678 16365 3712
rect 11929 3644 16365 3678
rect 11929 3610 11949 3644
rect 11983 3610 12018 3644
rect 12052 3610 12087 3644
rect 12121 3610 12156 3644
rect 12190 3610 12225 3644
rect 12259 3610 12294 3644
rect 12328 3610 12363 3644
rect 12397 3610 12432 3644
rect 12466 3610 12501 3644
rect 12535 3610 12570 3644
rect 12604 3610 12639 3644
rect 12673 3610 12708 3644
rect 12742 3610 12777 3644
rect 12811 3610 12846 3644
rect 12880 3610 12915 3644
rect 12949 3610 12984 3644
rect 13018 3610 13053 3644
rect 13087 3610 13122 3644
rect 13156 3610 13191 3644
rect 13225 3610 13260 3644
rect 13294 3610 13329 3644
rect 13363 3610 13398 3644
rect 13432 3610 13467 3644
rect 13501 3610 13536 3644
rect 13570 3610 13605 3644
rect 13639 3610 13674 3644
rect 13708 3610 13743 3644
rect 13777 3610 13812 3644
rect 13846 3610 13881 3644
rect 13915 3610 13950 3644
rect 13984 3610 14019 3644
rect 14053 3610 14088 3644
rect 14122 3610 14157 3644
rect 14191 3610 14226 3644
rect 14260 3610 14295 3644
rect 14329 3610 14364 3644
rect 14398 3610 14433 3644
rect 14467 3610 14502 3644
rect 14536 3610 14571 3644
rect 14605 3610 14640 3644
rect 14674 3610 14709 3644
rect 14743 3610 14778 3644
rect 14812 3610 14847 3644
rect 14881 3610 14916 3644
rect 14950 3610 14985 3644
rect 15019 3610 15054 3644
rect 15088 3610 15123 3644
rect 15157 3610 15192 3644
rect 15226 3610 15261 3644
rect 15295 3610 15330 3644
rect 15364 3610 15399 3644
rect 15433 3610 15468 3644
rect 15502 3610 15537 3644
rect 15571 3610 15606 3644
rect 15640 3610 15675 3644
rect 15709 3610 15744 3644
rect 15778 3610 15813 3644
rect 15847 3610 15882 3644
rect 15916 3610 15951 3644
rect 15985 3610 16020 3644
rect 16054 3610 16089 3644
rect 16123 3610 16158 3644
rect 16192 3610 16227 3644
rect 16261 3610 16296 3644
rect 16330 3610 16365 3644
rect 11929 3609 16365 3610
rect 2262 3542 2304 3576
rect 2338 3542 2374 3576
rect 2408 3542 2444 3576
rect 2478 3542 2514 3576
rect 2548 3542 2584 3576
rect 2618 3542 2654 3576
rect 2688 3542 2724 3576
rect 2758 3542 2794 3576
rect 2828 3542 2864 3576
rect 2898 3542 2934 3576
rect 2968 3542 3004 3576
rect 3038 3542 3074 3576
rect 3108 3542 3144 3576
rect 3178 3542 3214 3576
rect 3248 3542 3284 3576
rect 3318 3542 3354 3576
rect 3388 3542 3424 3576
rect 3458 3542 3494 3576
rect 3528 3542 3563 3576
rect 3597 3542 3632 3576
rect 3666 3542 3701 3576
rect 3735 3542 3770 3576
rect 3804 3542 3839 3576
rect 3873 3542 3908 3576
rect 3942 3542 3977 3576
rect 4011 3542 4046 3576
rect 4080 3542 4115 3576
rect 4149 3542 4184 3576
rect 4218 3542 4253 3576
rect 4287 3542 4322 3576
rect 4356 3542 4391 3576
rect 4425 3542 4449 3576
rect 11929 3576 11953 3609
rect 11987 3576 12026 3609
rect 12060 3576 12099 3609
rect 12133 3576 12172 3609
rect 12206 3576 12245 3609
rect 12279 3576 12318 3609
rect 12352 3576 12391 3609
rect 12425 3576 12464 3609
rect 12498 3576 12537 3609
rect 12571 3576 12610 3609
rect 12644 3576 12683 3609
rect 12717 3576 12756 3609
rect 12790 3576 12829 3609
rect 12863 3576 12902 3609
rect 12936 3576 12975 3609
rect 13009 3576 13048 3609
rect 13082 3576 13121 3609
rect 13155 3576 13194 3609
rect 13228 3576 13267 3609
rect 13301 3576 13340 3609
rect 13374 3576 13413 3609
rect 13447 3576 13486 3609
rect 13520 3576 13559 3609
rect 13593 3576 13632 3609
rect 13666 3576 13705 3609
rect 13739 3576 13778 3609
rect 2262 3508 4449 3542
rect 2262 3474 2304 3508
rect 2338 3474 2374 3508
rect 2408 3474 2444 3508
rect 2478 3474 2514 3508
rect 2548 3474 2584 3508
rect 2618 3474 2654 3508
rect 2688 3474 2724 3508
rect 2758 3474 2794 3508
rect 2828 3474 2864 3508
rect 2898 3474 2934 3508
rect 2968 3474 3004 3508
rect 3038 3474 3074 3508
rect 3108 3474 3144 3508
rect 3178 3474 3214 3508
rect 3248 3474 3284 3508
rect 3318 3474 3354 3508
rect 3388 3474 3424 3508
rect 3458 3474 3494 3508
rect 3528 3474 3563 3508
rect 3597 3474 3632 3508
rect 3666 3474 3701 3508
rect 3735 3474 3770 3508
rect 3804 3474 3839 3508
rect 3873 3474 3908 3508
rect 3942 3474 3977 3508
rect 4011 3474 4046 3508
rect 4080 3474 4115 3508
rect 4149 3474 4184 3508
rect 4218 3474 4253 3508
rect 4287 3474 4322 3508
rect 4356 3474 4391 3508
rect 4425 3474 4449 3508
rect 2262 3440 4449 3474
rect -2716 3344 -2680 3378
rect -2646 3344 -2610 3378
rect -2576 3344 -2540 3378
rect -2506 3344 -2470 3378
rect -2436 3344 -2400 3378
rect -2366 3344 -2330 3378
rect -2296 3344 -2260 3378
rect -2226 3344 -2190 3378
rect -2156 3344 -2120 3378
rect -2086 3344 -2050 3378
rect -2016 3344 -1980 3378
rect -1946 3344 -1910 3378
rect -1876 3344 -1840 3378
rect -1806 3344 -1770 3378
rect -1736 3344 -1700 3378
rect -1666 3344 -1630 3378
rect -1596 3344 -1560 3378
rect -1526 3344 -1490 3378
rect -1456 3344 -1421 3378
rect -1387 3344 -1352 3378
rect -1318 3344 -1283 3378
rect -1249 3344 -1214 3378
rect -1180 3344 -1145 3378
rect -1111 3344 -1076 3378
rect -1042 3344 -1007 3378
rect -973 3344 -938 3378
rect -904 3344 -869 3378
rect -835 3344 -800 3378
rect -766 3344 -731 3378
rect -697 3344 -662 3378
rect -628 3344 -593 3378
rect -559 3344 -524 3378
rect -490 3344 -455 3378
rect -421 3344 -386 3378
rect -352 3344 -317 3378
rect -283 3344 -248 3378
rect -2750 3308 -214 3344
rect 45 3340 79 3374
rect -2716 3274 -2680 3308
rect -2646 3274 -2610 3308
rect -2576 3274 -2540 3308
rect -2506 3274 -2470 3308
rect -2436 3274 -2400 3308
rect -2366 3274 -2330 3308
rect -2296 3274 -2260 3308
rect -2226 3274 -2190 3308
rect -2156 3274 -2120 3308
rect -2086 3274 -2050 3308
rect -2016 3274 -1980 3308
rect -1946 3274 -1910 3308
rect -1876 3274 -1840 3308
rect -1806 3274 -1770 3308
rect -1736 3274 -1700 3308
rect -1666 3274 -1630 3308
rect -1596 3274 -1560 3308
rect -1526 3274 -1490 3308
rect -1456 3274 -1421 3308
rect -1387 3274 -1352 3308
rect -1318 3274 -1283 3308
rect -1249 3274 -1214 3308
rect -1180 3274 -1145 3308
rect -1111 3274 -1076 3308
rect -1042 3274 -1007 3308
rect -973 3274 -938 3308
rect -904 3274 -869 3308
rect -835 3274 -800 3308
rect -766 3274 -731 3308
rect -697 3274 -662 3308
rect -628 3274 -593 3308
rect -559 3274 -524 3308
rect -490 3274 -455 3308
rect -421 3274 -386 3308
rect -352 3274 -317 3308
rect -283 3274 -248 3308
rect 29 3306 45 3340
rect 79 3306 95 3340
rect 443 3302 509 3408
rect 2262 3406 2304 3440
rect 2338 3406 2374 3440
rect 2408 3406 2444 3440
rect 2478 3406 2514 3440
rect 2548 3406 2584 3440
rect 2618 3406 2654 3440
rect 2688 3406 2724 3440
rect 2758 3406 2794 3440
rect 2828 3406 2864 3440
rect 2898 3406 2934 3440
rect 2968 3406 3004 3440
rect 3038 3406 3074 3440
rect 3108 3406 3144 3440
rect 3178 3406 3214 3440
rect 3248 3406 3284 3440
rect 3318 3406 3354 3440
rect 3388 3406 3424 3440
rect 3458 3406 3494 3440
rect 3528 3406 3563 3440
rect 3597 3406 3632 3440
rect 3666 3406 3701 3440
rect 3735 3406 3770 3440
rect 3804 3406 3839 3440
rect 3873 3406 3908 3440
rect 3942 3406 3977 3440
rect 4011 3406 4046 3440
rect 4080 3406 4115 3440
rect 4149 3406 4184 3440
rect 4218 3406 4253 3440
rect 4287 3406 4322 3440
rect 4356 3406 4391 3440
rect 4425 3406 4449 3440
rect 2262 3372 4449 3406
rect 4505 3537 4529 3571
rect 4563 3537 4598 3571
rect 4632 3537 4667 3571
rect 4701 3537 4736 3571
rect 4770 3537 4805 3571
rect 4839 3537 4874 3571
rect 4908 3537 4943 3571
rect 4977 3537 5012 3571
rect 5046 3537 5081 3571
rect 5115 3537 5150 3571
rect 5184 3537 5219 3571
rect 5253 3537 5288 3571
rect 5322 3537 5357 3571
rect 5391 3537 5426 3571
rect 5460 3537 5495 3571
rect 5529 3537 5564 3571
rect 5598 3537 5633 3571
rect 5667 3537 5702 3571
rect 5736 3537 5771 3571
rect 5805 3537 5840 3571
rect 5874 3537 5909 3571
rect 5943 3537 5978 3571
rect 6012 3537 6047 3571
rect 6081 3537 6116 3571
rect 6150 3537 6185 3571
rect 6219 3537 6254 3571
rect 6288 3537 6323 3571
rect 6357 3537 6392 3571
rect 6426 3537 6461 3571
rect 6495 3537 6530 3571
rect 6564 3537 6599 3571
rect 6633 3537 6668 3571
rect 6702 3537 6737 3571
rect 6771 3537 6806 3571
rect 6840 3537 6875 3571
rect 6909 3537 6944 3571
rect 6978 3537 7013 3571
rect 7047 3537 7082 3571
rect 7116 3537 7151 3571
rect 7185 3537 7220 3571
rect 4505 3503 7220 3537
rect 4505 3469 4529 3503
rect 4563 3469 4598 3503
rect 4632 3469 4667 3503
rect 4701 3469 4736 3503
rect 4770 3469 4805 3503
rect 4839 3469 4874 3503
rect 4908 3469 4943 3503
rect 4977 3469 5012 3503
rect 5046 3469 5081 3503
rect 5115 3469 5150 3503
rect 5184 3469 5219 3503
rect 5253 3469 5288 3503
rect 5322 3469 5357 3503
rect 5391 3469 5426 3503
rect 5460 3469 5495 3503
rect 5529 3469 5564 3503
rect 5598 3469 5633 3503
rect 5667 3469 5702 3503
rect 5736 3469 5771 3503
rect 5805 3469 5840 3503
rect 5874 3469 5909 3503
rect 5943 3469 5978 3503
rect 6012 3469 6047 3503
rect 6081 3469 6116 3503
rect 6150 3469 6185 3503
rect 6219 3469 6254 3503
rect 6288 3469 6323 3503
rect 6357 3469 6392 3503
rect 6426 3469 6461 3503
rect 6495 3469 6530 3503
rect 6564 3469 6599 3503
rect 6633 3469 6668 3503
rect 6702 3469 6737 3503
rect 6771 3469 6806 3503
rect 6840 3469 6875 3503
rect 6909 3469 6944 3503
rect 6978 3469 7013 3503
rect 7047 3469 7082 3503
rect 7116 3469 7151 3503
rect 7185 3469 7220 3503
rect 4505 3435 7220 3469
rect 4505 3401 4529 3435
rect 4563 3401 4598 3435
rect 4632 3401 4667 3435
rect 4701 3401 4736 3435
rect 4770 3401 4805 3435
rect 4839 3401 4874 3435
rect 4908 3401 4943 3435
rect 4977 3401 5012 3435
rect 5046 3401 5081 3435
rect 5115 3401 5150 3435
rect 5184 3401 5219 3435
rect 5253 3401 5288 3435
rect 5322 3401 5357 3435
rect 5391 3401 5426 3435
rect 5460 3401 5495 3435
rect 5529 3401 5564 3435
rect 5598 3401 5633 3435
rect 5667 3401 5702 3435
rect 5736 3401 5771 3435
rect 5805 3401 5840 3435
rect 5874 3401 5909 3435
rect 5943 3401 5978 3435
rect 6012 3401 6047 3435
rect 6081 3401 6116 3435
rect 6150 3401 6185 3435
rect 6219 3401 6254 3435
rect 6288 3401 6323 3435
rect 6357 3401 6392 3435
rect 6426 3401 6461 3435
rect 6495 3401 6530 3435
rect 6564 3401 6599 3435
rect 6633 3401 6668 3435
rect 6702 3401 6737 3435
rect 6771 3401 6806 3435
rect 6840 3401 6875 3435
rect 6909 3401 6944 3435
rect 6978 3401 7013 3435
rect 7047 3401 7082 3435
rect 7116 3401 7151 3435
rect 7185 3401 7220 3435
rect 11674 3401 11698 3571
rect 11929 3542 11949 3576
rect 11987 3575 12018 3576
rect 12060 3575 12087 3576
rect 12133 3575 12156 3576
rect 12206 3575 12225 3576
rect 12279 3575 12294 3576
rect 12352 3575 12363 3576
rect 12425 3575 12432 3576
rect 12498 3575 12501 3576
rect 11983 3542 12018 3575
rect 12052 3542 12087 3575
rect 12121 3542 12156 3575
rect 12190 3542 12225 3575
rect 12259 3542 12294 3575
rect 12328 3542 12363 3575
rect 12397 3542 12432 3575
rect 12466 3542 12501 3575
rect 12535 3575 12537 3576
rect 12604 3575 12610 3576
rect 12673 3575 12683 3576
rect 12742 3575 12756 3576
rect 12811 3575 12829 3576
rect 12880 3575 12902 3576
rect 12949 3575 12975 3576
rect 13018 3575 13048 3576
rect 13087 3575 13121 3576
rect 12535 3542 12570 3575
rect 12604 3542 12639 3575
rect 12673 3542 12708 3575
rect 12742 3542 12777 3575
rect 12811 3542 12846 3575
rect 12880 3542 12915 3575
rect 12949 3542 12984 3575
rect 13018 3542 13053 3575
rect 13087 3542 13122 3575
rect 13156 3542 13191 3576
rect 13228 3575 13260 3576
rect 13301 3575 13329 3576
rect 13374 3575 13398 3576
rect 13447 3575 13467 3576
rect 13520 3575 13536 3576
rect 13593 3575 13605 3576
rect 13666 3575 13674 3576
rect 13739 3575 13743 3576
rect 13225 3542 13260 3575
rect 13294 3542 13329 3575
rect 13363 3542 13398 3575
rect 13432 3542 13467 3575
rect 13501 3542 13536 3575
rect 13570 3542 13605 3575
rect 13639 3542 13674 3575
rect 13708 3542 13743 3575
rect 13777 3575 13778 3576
rect 13812 3576 13851 3609
rect 13885 3576 13924 3609
rect 13958 3576 13997 3609
rect 14031 3576 14070 3609
rect 14104 3576 14143 3609
rect 14177 3576 14216 3609
rect 14250 3576 14289 3609
rect 14323 3576 14362 3609
rect 14396 3576 14435 3609
rect 14469 3576 14508 3609
rect 14542 3576 14581 3609
rect 14615 3576 14654 3609
rect 14688 3576 14727 3609
rect 14761 3576 14800 3609
rect 14834 3576 14873 3609
rect 14907 3576 14946 3609
rect 14980 3576 15019 3609
rect 13777 3542 13812 3575
rect 13846 3575 13851 3576
rect 13915 3575 13924 3576
rect 13984 3575 13997 3576
rect 14053 3575 14070 3576
rect 14122 3575 14143 3576
rect 14191 3575 14216 3576
rect 14260 3575 14289 3576
rect 14329 3575 14362 3576
rect 13846 3542 13881 3575
rect 13915 3542 13950 3575
rect 13984 3542 14019 3575
rect 14053 3542 14088 3575
rect 14122 3542 14157 3575
rect 14191 3542 14226 3575
rect 14260 3542 14295 3575
rect 14329 3542 14364 3575
rect 14398 3542 14433 3576
rect 14469 3575 14502 3576
rect 14542 3575 14571 3576
rect 14615 3575 14640 3576
rect 14688 3575 14709 3576
rect 14761 3575 14778 3576
rect 14834 3575 14847 3576
rect 14907 3575 14916 3576
rect 14980 3575 14985 3576
rect 14467 3542 14502 3575
rect 14536 3542 14571 3575
rect 14605 3542 14640 3575
rect 14674 3542 14709 3575
rect 14743 3542 14778 3575
rect 14812 3542 14847 3575
rect 14881 3542 14916 3575
rect 14950 3542 14985 3575
rect 15053 3576 15092 3609
rect 15126 3576 15165 3609
rect 15199 3576 15238 3609
rect 15272 3576 15311 3609
rect 15345 3576 15384 3609
rect 15418 3576 15457 3609
rect 15491 3576 15530 3609
rect 15564 3576 15603 3609
rect 15637 3576 15676 3609
rect 15710 3576 15749 3609
rect 15783 3576 15822 3609
rect 15856 3576 15895 3609
rect 15929 3576 15968 3609
rect 16002 3576 16041 3609
rect 16075 3576 16114 3609
rect 16148 3576 16187 3609
rect 16221 3576 16260 3609
rect 16294 3576 16333 3609
rect 15053 3575 15054 3576
rect 15019 3542 15054 3575
rect 15088 3575 15092 3576
rect 15157 3575 15165 3576
rect 15226 3575 15238 3576
rect 15295 3575 15311 3576
rect 15364 3575 15384 3576
rect 15433 3575 15457 3576
rect 15502 3575 15530 3576
rect 15571 3575 15603 3576
rect 15088 3542 15123 3575
rect 15157 3542 15192 3575
rect 15226 3542 15261 3575
rect 15295 3542 15330 3575
rect 15364 3542 15399 3575
rect 15433 3542 15468 3575
rect 15502 3542 15537 3575
rect 15571 3542 15606 3575
rect 15640 3542 15675 3576
rect 15710 3575 15744 3576
rect 15783 3575 15813 3576
rect 15856 3575 15882 3576
rect 15929 3575 15951 3576
rect 16002 3575 16020 3576
rect 16075 3575 16089 3576
rect 16148 3575 16158 3576
rect 16221 3575 16227 3576
rect 16294 3575 16296 3576
rect 15709 3542 15744 3575
rect 15778 3542 15813 3575
rect 15847 3542 15882 3575
rect 15916 3542 15951 3575
rect 15985 3542 16020 3575
rect 16054 3542 16089 3575
rect 16123 3542 16158 3575
rect 16192 3542 16227 3575
rect 16261 3542 16296 3575
rect 16330 3575 16333 3576
rect 16330 3542 16365 3575
rect 11929 3537 16365 3542
rect 11929 3508 11953 3537
rect 11987 3508 12026 3537
rect 12060 3508 12099 3537
rect 12133 3508 12172 3537
rect 12206 3508 12245 3537
rect 12279 3508 12318 3537
rect 12352 3508 12391 3537
rect 12425 3508 12464 3537
rect 12498 3508 12537 3537
rect 12571 3508 12610 3537
rect 12644 3508 12683 3537
rect 12717 3508 12756 3537
rect 12790 3508 12829 3537
rect 12863 3508 12902 3537
rect 12936 3508 12975 3537
rect 13009 3508 13048 3537
rect 13082 3508 13121 3537
rect 13155 3508 13194 3537
rect 13228 3508 13267 3537
rect 13301 3508 13340 3537
rect 13374 3508 13413 3537
rect 13447 3508 13486 3537
rect 13520 3508 13559 3537
rect 13593 3508 13632 3537
rect 13666 3508 13705 3537
rect 13739 3508 13778 3537
rect 11929 3474 11949 3508
rect 11987 3503 12018 3508
rect 12060 3503 12087 3508
rect 12133 3503 12156 3508
rect 12206 3503 12225 3508
rect 12279 3503 12294 3508
rect 12352 3503 12363 3508
rect 12425 3503 12432 3508
rect 12498 3503 12501 3508
rect 11983 3474 12018 3503
rect 12052 3474 12087 3503
rect 12121 3474 12156 3503
rect 12190 3474 12225 3503
rect 12259 3474 12294 3503
rect 12328 3474 12363 3503
rect 12397 3474 12432 3503
rect 12466 3474 12501 3503
rect 12535 3503 12537 3508
rect 12604 3503 12610 3508
rect 12673 3503 12683 3508
rect 12742 3503 12756 3508
rect 12811 3503 12829 3508
rect 12880 3503 12902 3508
rect 12949 3503 12975 3508
rect 13018 3503 13048 3508
rect 13087 3503 13121 3508
rect 12535 3474 12570 3503
rect 12604 3474 12639 3503
rect 12673 3474 12708 3503
rect 12742 3474 12777 3503
rect 12811 3474 12846 3503
rect 12880 3474 12915 3503
rect 12949 3474 12984 3503
rect 13018 3474 13053 3503
rect 13087 3474 13122 3503
rect 13156 3474 13191 3508
rect 13228 3503 13260 3508
rect 13301 3503 13329 3508
rect 13374 3503 13398 3508
rect 13447 3503 13467 3508
rect 13520 3503 13536 3508
rect 13593 3503 13605 3508
rect 13666 3503 13674 3508
rect 13739 3503 13743 3508
rect 13225 3474 13260 3503
rect 13294 3474 13329 3503
rect 13363 3474 13398 3503
rect 13432 3474 13467 3503
rect 13501 3474 13536 3503
rect 13570 3474 13605 3503
rect 13639 3474 13674 3503
rect 13708 3474 13743 3503
rect 13777 3503 13778 3508
rect 13812 3508 13851 3537
rect 13885 3508 13924 3537
rect 13958 3508 13997 3537
rect 14031 3508 14070 3537
rect 14104 3508 14143 3537
rect 14177 3508 14216 3537
rect 14250 3508 14289 3537
rect 14323 3508 14362 3537
rect 14396 3508 14435 3537
rect 14469 3508 14508 3537
rect 14542 3508 14581 3537
rect 14615 3508 14654 3537
rect 14688 3508 14727 3537
rect 14761 3508 14800 3537
rect 14834 3508 14873 3537
rect 14907 3508 14946 3537
rect 14980 3508 15019 3537
rect 13777 3474 13812 3503
rect 13846 3503 13851 3508
rect 13915 3503 13924 3508
rect 13984 3503 13997 3508
rect 14053 3503 14070 3508
rect 14122 3503 14143 3508
rect 14191 3503 14216 3508
rect 14260 3503 14289 3508
rect 14329 3503 14362 3508
rect 13846 3474 13881 3503
rect 13915 3474 13950 3503
rect 13984 3474 14019 3503
rect 14053 3474 14088 3503
rect 14122 3474 14157 3503
rect 14191 3474 14226 3503
rect 14260 3474 14295 3503
rect 14329 3474 14364 3503
rect 14398 3474 14433 3508
rect 14469 3503 14502 3508
rect 14542 3503 14571 3508
rect 14615 3503 14640 3508
rect 14688 3503 14709 3508
rect 14761 3503 14778 3508
rect 14834 3503 14847 3508
rect 14907 3503 14916 3508
rect 14980 3503 14985 3508
rect 14467 3474 14502 3503
rect 14536 3474 14571 3503
rect 14605 3474 14640 3503
rect 14674 3474 14709 3503
rect 14743 3474 14778 3503
rect 14812 3474 14847 3503
rect 14881 3474 14916 3503
rect 14950 3474 14985 3503
rect 15053 3508 15092 3537
rect 15126 3508 15165 3537
rect 15199 3508 15238 3537
rect 15272 3508 15311 3537
rect 15345 3508 15384 3537
rect 15418 3508 15457 3537
rect 15491 3508 15530 3537
rect 15564 3508 15603 3537
rect 15637 3508 15676 3537
rect 15710 3508 15749 3537
rect 15783 3508 15822 3537
rect 15856 3508 15895 3537
rect 15929 3508 15968 3537
rect 16002 3508 16041 3537
rect 16075 3508 16114 3537
rect 16148 3508 16187 3537
rect 16221 3508 16260 3537
rect 16294 3508 16333 3537
rect 15053 3503 15054 3508
rect 15019 3474 15054 3503
rect 15088 3503 15092 3508
rect 15157 3503 15165 3508
rect 15226 3503 15238 3508
rect 15295 3503 15311 3508
rect 15364 3503 15384 3508
rect 15433 3503 15457 3508
rect 15502 3503 15530 3508
rect 15571 3503 15603 3508
rect 15088 3474 15123 3503
rect 15157 3474 15192 3503
rect 15226 3474 15261 3503
rect 15295 3474 15330 3503
rect 15364 3474 15399 3503
rect 15433 3474 15468 3503
rect 15502 3474 15537 3503
rect 15571 3474 15606 3503
rect 15640 3474 15675 3508
rect 15710 3503 15744 3508
rect 15783 3503 15813 3508
rect 15856 3503 15882 3508
rect 15929 3503 15951 3508
rect 16002 3503 16020 3508
rect 16075 3503 16089 3508
rect 16148 3503 16158 3508
rect 16221 3503 16227 3508
rect 16294 3503 16296 3508
rect 15709 3474 15744 3503
rect 15778 3474 15813 3503
rect 15847 3474 15882 3503
rect 15916 3474 15951 3503
rect 15985 3474 16020 3503
rect 16054 3474 16089 3503
rect 16123 3474 16158 3503
rect 16192 3474 16227 3503
rect 16261 3474 16296 3503
rect 16330 3503 16333 3508
rect 16330 3474 16365 3503
rect 11929 3465 16365 3474
rect 11929 3440 11953 3465
rect 11987 3440 12026 3465
rect 12060 3440 12099 3465
rect 12133 3440 12172 3465
rect 12206 3440 12245 3465
rect 12279 3440 12318 3465
rect 12352 3440 12391 3465
rect 12425 3440 12464 3465
rect 12498 3440 12537 3465
rect 12571 3440 12610 3465
rect 12644 3440 12683 3465
rect 12717 3440 12756 3465
rect 12790 3440 12829 3465
rect 12863 3440 12902 3465
rect 12936 3440 12975 3465
rect 13009 3440 13048 3465
rect 13082 3440 13121 3465
rect 13155 3440 13194 3465
rect 13228 3440 13267 3465
rect 13301 3440 13340 3465
rect 13374 3440 13413 3465
rect 13447 3440 13486 3465
rect 13520 3440 13559 3465
rect 13593 3440 13632 3465
rect 13666 3440 13705 3465
rect 13739 3440 13778 3465
rect 11929 3406 11949 3440
rect 11987 3431 12018 3440
rect 12060 3431 12087 3440
rect 12133 3431 12156 3440
rect 12206 3431 12225 3440
rect 12279 3431 12294 3440
rect 12352 3431 12363 3440
rect 12425 3431 12432 3440
rect 12498 3431 12501 3440
rect 11983 3406 12018 3431
rect 12052 3406 12087 3431
rect 12121 3406 12156 3431
rect 12190 3406 12225 3431
rect 12259 3406 12294 3431
rect 12328 3406 12363 3431
rect 12397 3406 12432 3431
rect 12466 3406 12501 3431
rect 12535 3431 12537 3440
rect 12604 3431 12610 3440
rect 12673 3431 12683 3440
rect 12742 3431 12756 3440
rect 12811 3431 12829 3440
rect 12880 3431 12902 3440
rect 12949 3431 12975 3440
rect 13018 3431 13048 3440
rect 13087 3431 13121 3440
rect 12535 3406 12570 3431
rect 12604 3406 12639 3431
rect 12673 3406 12708 3431
rect 12742 3406 12777 3431
rect 12811 3406 12846 3431
rect 12880 3406 12915 3431
rect 12949 3406 12984 3431
rect 13018 3406 13053 3431
rect 13087 3406 13122 3431
rect 13156 3406 13191 3440
rect 13228 3431 13260 3440
rect 13301 3431 13329 3440
rect 13374 3431 13398 3440
rect 13447 3431 13467 3440
rect 13520 3431 13536 3440
rect 13593 3431 13605 3440
rect 13666 3431 13674 3440
rect 13739 3431 13743 3440
rect 13225 3406 13260 3431
rect 13294 3406 13329 3431
rect 13363 3406 13398 3431
rect 13432 3406 13467 3431
rect 13501 3406 13536 3431
rect 13570 3406 13605 3431
rect 13639 3406 13674 3431
rect 13708 3406 13743 3431
rect 13777 3431 13778 3440
rect 13812 3440 13851 3465
rect 13885 3440 13924 3465
rect 13958 3440 13997 3465
rect 14031 3440 14070 3465
rect 14104 3440 14143 3465
rect 14177 3440 14216 3465
rect 14250 3440 14289 3465
rect 14323 3440 14362 3465
rect 14396 3440 14435 3465
rect 14469 3440 14508 3465
rect 14542 3440 14581 3465
rect 14615 3440 14654 3465
rect 14688 3440 14727 3465
rect 14761 3440 14800 3465
rect 14834 3440 14873 3465
rect 14907 3440 14946 3465
rect 14980 3440 15019 3465
rect 13777 3406 13812 3431
rect 13846 3431 13851 3440
rect 13915 3431 13924 3440
rect 13984 3431 13997 3440
rect 14053 3431 14070 3440
rect 14122 3431 14143 3440
rect 14191 3431 14216 3440
rect 14260 3431 14289 3440
rect 14329 3431 14362 3440
rect 13846 3406 13881 3431
rect 13915 3406 13950 3431
rect 13984 3406 14019 3431
rect 14053 3406 14088 3431
rect 14122 3406 14157 3431
rect 14191 3406 14226 3431
rect 14260 3406 14295 3431
rect 14329 3406 14364 3431
rect 14398 3406 14433 3440
rect 14469 3431 14502 3440
rect 14542 3431 14571 3440
rect 14615 3431 14640 3440
rect 14688 3431 14709 3440
rect 14761 3431 14778 3440
rect 14834 3431 14847 3440
rect 14907 3431 14916 3440
rect 14980 3431 14985 3440
rect 14467 3406 14502 3431
rect 14536 3406 14571 3431
rect 14605 3406 14640 3431
rect 14674 3406 14709 3431
rect 14743 3406 14778 3431
rect 14812 3406 14847 3431
rect 14881 3406 14916 3431
rect 14950 3406 14985 3431
rect 15053 3440 15092 3465
rect 15126 3440 15165 3465
rect 15199 3440 15238 3465
rect 15272 3440 15311 3465
rect 15345 3440 15384 3465
rect 15418 3440 15457 3465
rect 15491 3440 15530 3465
rect 15564 3440 15603 3465
rect 15637 3440 15676 3465
rect 15710 3440 15749 3465
rect 15783 3440 15822 3465
rect 15856 3440 15895 3465
rect 15929 3440 15968 3465
rect 16002 3440 16041 3465
rect 16075 3440 16114 3465
rect 16148 3440 16187 3465
rect 16221 3440 16260 3465
rect 16294 3440 16333 3465
rect 15053 3431 15054 3440
rect 15019 3406 15054 3431
rect 15088 3431 15092 3440
rect 15157 3431 15165 3440
rect 15226 3431 15238 3440
rect 15295 3431 15311 3440
rect 15364 3431 15384 3440
rect 15433 3431 15457 3440
rect 15502 3431 15530 3440
rect 15571 3431 15603 3440
rect 15088 3406 15123 3431
rect 15157 3406 15192 3431
rect 15226 3406 15261 3431
rect 15295 3406 15330 3431
rect 15364 3406 15399 3431
rect 15433 3406 15468 3431
rect 15502 3406 15537 3431
rect 15571 3406 15606 3431
rect 15640 3406 15675 3440
rect 15710 3431 15744 3440
rect 15783 3431 15813 3440
rect 15856 3431 15882 3440
rect 15929 3431 15951 3440
rect 16002 3431 16020 3440
rect 16075 3431 16089 3440
rect 16148 3431 16158 3440
rect 16221 3431 16227 3440
rect 16294 3431 16296 3440
rect 15709 3406 15744 3431
rect 15778 3406 15813 3431
rect 15847 3406 15882 3431
rect 15916 3406 15951 3431
rect 15985 3406 16020 3431
rect 16054 3406 16089 3431
rect 16123 3406 16158 3431
rect 16192 3406 16227 3431
rect 16261 3406 16296 3431
rect 16330 3431 16333 3440
rect 16330 3406 16365 3431
rect 2262 3338 2304 3372
rect 2338 3338 2374 3372
rect 2408 3338 2444 3372
rect 2478 3338 2514 3372
rect 2548 3338 2584 3372
rect 2618 3338 2654 3372
rect 2688 3338 2724 3372
rect 2758 3338 2794 3372
rect 2828 3338 2864 3372
rect 2898 3338 2934 3372
rect 2968 3338 3004 3372
rect 3038 3338 3074 3372
rect 3108 3338 3144 3372
rect 3178 3338 3214 3372
rect 3248 3338 3284 3372
rect 3318 3338 3354 3372
rect 3388 3338 3424 3372
rect 3458 3338 3494 3372
rect 3528 3338 3563 3372
rect 3597 3338 3632 3372
rect 3666 3338 3701 3372
rect 3735 3338 3770 3372
rect 3804 3338 3839 3372
rect 3873 3338 3908 3372
rect 3942 3338 3977 3372
rect 4011 3338 4046 3372
rect 4080 3338 4115 3372
rect 4149 3338 4184 3372
rect 4218 3338 4253 3372
rect 4287 3338 4322 3372
rect 4356 3338 4391 3372
rect 4425 3338 4449 3372
rect 2262 3304 4449 3338
rect -2750 3238 -214 3274
rect -2716 3204 -2680 3238
rect -2646 3204 -2610 3238
rect -2576 3204 -2540 3238
rect -2506 3204 -2470 3238
rect -2436 3204 -2400 3238
rect -2366 3204 -2330 3238
rect -2296 3204 -2260 3238
rect -2226 3204 -2190 3238
rect -2156 3204 -2120 3238
rect -2086 3204 -2050 3238
rect -2016 3204 -1980 3238
rect -1946 3204 -1910 3238
rect -1876 3204 -1840 3238
rect -1806 3204 -1770 3238
rect -1736 3204 -1700 3238
rect -1666 3204 -1630 3238
rect -1596 3204 -1560 3238
rect -1526 3204 -1490 3238
rect -1456 3204 -1421 3238
rect -1387 3204 -1352 3238
rect -1318 3204 -1283 3238
rect -1249 3204 -1214 3238
rect -1180 3204 -1145 3238
rect -1111 3204 -1076 3238
rect -1042 3204 -1007 3238
rect -973 3204 -938 3238
rect -904 3204 -869 3238
rect -835 3204 -800 3238
rect -766 3204 -731 3238
rect -697 3204 -662 3238
rect -628 3204 -593 3238
rect -559 3204 -524 3238
rect -490 3204 -455 3238
rect -421 3204 -386 3238
rect -352 3204 -317 3238
rect -283 3204 -248 3238
rect -2750 3168 -214 3204
rect -2716 3134 -2680 3168
rect -2646 3134 -2610 3168
rect -2576 3134 -2540 3168
rect -2506 3134 -2470 3168
rect -2436 3134 -2400 3168
rect -2366 3134 -2330 3168
rect -2296 3134 -2260 3168
rect -2226 3134 -2190 3168
rect -2156 3134 -2120 3168
rect -2086 3134 -2050 3168
rect -2016 3134 -1980 3168
rect -1946 3134 -1910 3168
rect -1876 3134 -1840 3168
rect -1806 3134 -1770 3168
rect -1736 3134 -1700 3168
rect -1666 3134 -1630 3168
rect -1596 3134 -1560 3168
rect -1526 3134 -1490 3168
rect -1456 3134 -1421 3168
rect -1387 3134 -1352 3168
rect -1318 3134 -1283 3168
rect -1249 3134 -1214 3168
rect -1180 3134 -1145 3168
rect -1111 3134 -1076 3168
rect -1042 3134 -1007 3168
rect -973 3134 -938 3168
rect -904 3134 -869 3168
rect -835 3134 -800 3168
rect -766 3134 -731 3168
rect -697 3134 -662 3168
rect -628 3134 -593 3168
rect -559 3134 -524 3168
rect -490 3134 -455 3168
rect -421 3134 -386 3168
rect -352 3134 -317 3168
rect -283 3134 -248 3168
rect 2262 3270 2304 3304
rect 2338 3270 2374 3304
rect 2408 3270 2444 3304
rect 2478 3270 2514 3304
rect 2548 3270 2584 3304
rect 2618 3270 2654 3304
rect 2688 3270 2724 3304
rect 2758 3270 2794 3304
rect 2828 3270 2864 3304
rect 2898 3270 2934 3304
rect 2968 3270 3004 3304
rect 3038 3270 3074 3304
rect 3108 3270 3144 3304
rect 3178 3270 3214 3304
rect 3248 3270 3284 3304
rect 3318 3270 3354 3304
rect 3388 3270 3424 3304
rect 3458 3270 3494 3304
rect 3528 3270 3563 3304
rect 3597 3270 3632 3304
rect 3666 3270 3701 3304
rect 3735 3270 3770 3304
rect 3804 3270 3839 3304
rect 3873 3270 3908 3304
rect 3942 3270 3977 3304
rect 4011 3270 4046 3304
rect 4080 3270 4115 3304
rect 4149 3270 4184 3304
rect 4218 3270 4253 3304
rect 4287 3270 4322 3304
rect 4356 3270 4391 3304
rect 4425 3270 4449 3304
rect 2262 3236 4449 3270
rect 11929 3393 16365 3406
rect 11929 3372 11953 3393
rect 11987 3372 12026 3393
rect 12060 3372 12099 3393
rect 12133 3372 12172 3393
rect 12206 3372 12245 3393
rect 12279 3372 12318 3393
rect 12352 3372 12391 3393
rect 12425 3372 12464 3393
rect 12498 3372 12537 3393
rect 12571 3372 12610 3393
rect 12644 3372 12683 3393
rect 12717 3372 12756 3393
rect 12790 3372 12829 3393
rect 12863 3372 12902 3393
rect 12936 3372 12975 3393
rect 13009 3372 13048 3393
rect 13082 3372 13121 3393
rect 13155 3372 13194 3393
rect 13228 3372 13267 3393
rect 13301 3372 13340 3393
rect 13374 3372 13413 3393
rect 13447 3372 13486 3393
rect 13520 3372 13559 3393
rect 13593 3372 13632 3393
rect 13666 3372 13705 3393
rect 13739 3372 13778 3393
rect 11929 3338 11949 3372
rect 11987 3359 12018 3372
rect 12060 3359 12087 3372
rect 12133 3359 12156 3372
rect 12206 3359 12225 3372
rect 12279 3359 12294 3372
rect 12352 3359 12363 3372
rect 12425 3359 12432 3372
rect 12498 3359 12501 3372
rect 11983 3338 12018 3359
rect 12052 3338 12087 3359
rect 12121 3338 12156 3359
rect 12190 3338 12225 3359
rect 12259 3338 12294 3359
rect 12328 3338 12363 3359
rect 12397 3338 12432 3359
rect 12466 3338 12501 3359
rect 12535 3359 12537 3372
rect 12604 3359 12610 3372
rect 12673 3359 12683 3372
rect 12742 3359 12756 3372
rect 12811 3359 12829 3372
rect 12880 3359 12902 3372
rect 12949 3359 12975 3372
rect 13018 3359 13048 3372
rect 13087 3359 13121 3372
rect 12535 3338 12570 3359
rect 12604 3338 12639 3359
rect 12673 3338 12708 3359
rect 12742 3338 12777 3359
rect 12811 3338 12846 3359
rect 12880 3338 12915 3359
rect 12949 3338 12984 3359
rect 13018 3338 13053 3359
rect 13087 3338 13122 3359
rect 13156 3338 13191 3372
rect 13228 3359 13260 3372
rect 13301 3359 13329 3372
rect 13374 3359 13398 3372
rect 13447 3359 13467 3372
rect 13520 3359 13536 3372
rect 13593 3359 13605 3372
rect 13666 3359 13674 3372
rect 13739 3359 13743 3372
rect 13225 3338 13260 3359
rect 13294 3338 13329 3359
rect 13363 3338 13398 3359
rect 13432 3338 13467 3359
rect 13501 3338 13536 3359
rect 13570 3338 13605 3359
rect 13639 3338 13674 3359
rect 13708 3338 13743 3359
rect 13777 3359 13778 3372
rect 13812 3372 13851 3393
rect 13885 3372 13924 3393
rect 13958 3372 13997 3393
rect 14031 3372 14070 3393
rect 14104 3372 14143 3393
rect 14177 3372 14216 3393
rect 14250 3372 14289 3393
rect 14323 3372 14362 3393
rect 14396 3372 14435 3393
rect 14469 3372 14508 3393
rect 14542 3372 14581 3393
rect 14615 3372 14654 3393
rect 14688 3372 14727 3393
rect 14761 3372 14800 3393
rect 14834 3372 14873 3393
rect 14907 3372 14946 3393
rect 14980 3372 15019 3393
rect 13777 3338 13812 3359
rect 13846 3359 13851 3372
rect 13915 3359 13924 3372
rect 13984 3359 13997 3372
rect 14053 3359 14070 3372
rect 14122 3359 14143 3372
rect 14191 3359 14216 3372
rect 14260 3359 14289 3372
rect 14329 3359 14362 3372
rect 13846 3338 13881 3359
rect 13915 3338 13950 3359
rect 13984 3338 14019 3359
rect 14053 3338 14088 3359
rect 14122 3338 14157 3359
rect 14191 3338 14226 3359
rect 14260 3338 14295 3359
rect 14329 3338 14364 3359
rect 14398 3338 14433 3372
rect 14469 3359 14502 3372
rect 14542 3359 14571 3372
rect 14615 3359 14640 3372
rect 14688 3359 14709 3372
rect 14761 3359 14778 3372
rect 14834 3359 14847 3372
rect 14907 3359 14916 3372
rect 14980 3359 14985 3372
rect 14467 3338 14502 3359
rect 14536 3338 14571 3359
rect 14605 3338 14640 3359
rect 14674 3338 14709 3359
rect 14743 3338 14778 3359
rect 14812 3338 14847 3359
rect 14881 3338 14916 3359
rect 14950 3338 14985 3359
rect 15053 3372 15092 3393
rect 15126 3372 15165 3393
rect 15199 3372 15238 3393
rect 15272 3372 15311 3393
rect 15345 3372 15384 3393
rect 15418 3372 15457 3393
rect 15491 3372 15530 3393
rect 15564 3372 15603 3393
rect 15637 3372 15676 3393
rect 15710 3372 15749 3393
rect 15783 3372 15822 3393
rect 15856 3372 15895 3393
rect 15929 3372 15968 3393
rect 16002 3372 16041 3393
rect 16075 3372 16114 3393
rect 16148 3372 16187 3393
rect 16221 3372 16260 3393
rect 16294 3372 16333 3393
rect 15053 3359 15054 3372
rect 15019 3338 15054 3359
rect 15088 3359 15092 3372
rect 15157 3359 15165 3372
rect 15226 3359 15238 3372
rect 15295 3359 15311 3372
rect 15364 3359 15384 3372
rect 15433 3359 15457 3372
rect 15502 3359 15530 3372
rect 15571 3359 15603 3372
rect 15088 3338 15123 3359
rect 15157 3338 15192 3359
rect 15226 3338 15261 3359
rect 15295 3338 15330 3359
rect 15364 3338 15399 3359
rect 15433 3338 15468 3359
rect 15502 3338 15537 3359
rect 15571 3338 15606 3359
rect 15640 3338 15675 3372
rect 15710 3359 15744 3372
rect 15783 3359 15813 3372
rect 15856 3359 15882 3372
rect 15929 3359 15951 3372
rect 16002 3359 16020 3372
rect 16075 3359 16089 3372
rect 16148 3359 16158 3372
rect 16221 3359 16227 3372
rect 16294 3359 16296 3372
rect 15709 3338 15744 3359
rect 15778 3338 15813 3359
rect 15847 3338 15882 3359
rect 15916 3338 15951 3359
rect 15985 3338 16020 3359
rect 16054 3338 16089 3359
rect 16123 3338 16158 3359
rect 16192 3338 16227 3359
rect 16261 3338 16296 3359
rect 16330 3359 16333 3372
rect 16330 3338 16365 3359
rect 11929 3321 16365 3338
rect 11929 3304 11953 3321
rect 11987 3304 12026 3321
rect 12060 3304 12099 3321
rect 12133 3304 12172 3321
rect 12206 3304 12245 3321
rect 12279 3304 12318 3321
rect 12352 3304 12391 3321
rect 12425 3304 12464 3321
rect 12498 3304 12537 3321
rect 12571 3304 12610 3321
rect 12644 3304 12683 3321
rect 12717 3304 12756 3321
rect 12790 3304 12829 3321
rect 12863 3304 12902 3321
rect 12936 3304 12975 3321
rect 13009 3304 13048 3321
rect 13082 3304 13121 3321
rect 13155 3304 13194 3321
rect 13228 3304 13267 3321
rect 13301 3304 13340 3321
rect 13374 3304 13413 3321
rect 13447 3304 13486 3321
rect 13520 3304 13559 3321
rect 13593 3304 13632 3321
rect 13666 3304 13705 3321
rect 13739 3304 13778 3321
rect 11929 3270 11949 3304
rect 11987 3287 12018 3304
rect 12060 3287 12087 3304
rect 12133 3287 12156 3304
rect 12206 3287 12225 3304
rect 12279 3287 12294 3304
rect 12352 3287 12363 3304
rect 12425 3287 12432 3304
rect 12498 3287 12501 3304
rect 11983 3270 12018 3287
rect 12052 3270 12087 3287
rect 12121 3270 12156 3287
rect 12190 3270 12225 3287
rect 12259 3270 12294 3287
rect 12328 3270 12363 3287
rect 12397 3270 12432 3287
rect 12466 3270 12501 3287
rect 12535 3287 12537 3304
rect 12604 3287 12610 3304
rect 12673 3287 12683 3304
rect 12742 3287 12756 3304
rect 12811 3287 12829 3304
rect 12880 3287 12902 3304
rect 12949 3287 12975 3304
rect 13018 3287 13048 3304
rect 13087 3287 13121 3304
rect 12535 3270 12570 3287
rect 12604 3270 12639 3287
rect 12673 3270 12708 3287
rect 12742 3270 12777 3287
rect 12811 3270 12846 3287
rect 12880 3270 12915 3287
rect 12949 3270 12984 3287
rect 13018 3270 13053 3287
rect 13087 3270 13122 3287
rect 13156 3270 13191 3304
rect 13228 3287 13260 3304
rect 13301 3287 13329 3304
rect 13374 3287 13398 3304
rect 13447 3287 13467 3304
rect 13520 3287 13536 3304
rect 13593 3287 13605 3304
rect 13666 3287 13674 3304
rect 13739 3287 13743 3304
rect 13225 3270 13260 3287
rect 13294 3270 13329 3287
rect 13363 3270 13398 3287
rect 13432 3270 13467 3287
rect 13501 3270 13536 3287
rect 13570 3270 13605 3287
rect 13639 3270 13674 3287
rect 13708 3270 13743 3287
rect 13777 3287 13778 3304
rect 13812 3304 13851 3321
rect 13885 3304 13924 3321
rect 13958 3304 13997 3321
rect 14031 3304 14070 3321
rect 14104 3304 14143 3321
rect 14177 3304 14216 3321
rect 14250 3304 14289 3321
rect 14323 3304 14362 3321
rect 14396 3304 14435 3321
rect 14469 3304 14508 3321
rect 14542 3304 14581 3321
rect 14615 3304 14654 3321
rect 14688 3304 14727 3321
rect 14761 3304 14800 3321
rect 14834 3304 14873 3321
rect 14907 3304 14946 3321
rect 14980 3304 15019 3321
rect 13777 3270 13812 3287
rect 13846 3287 13851 3304
rect 13915 3287 13924 3304
rect 13984 3287 13997 3304
rect 14053 3287 14070 3304
rect 14122 3287 14143 3304
rect 14191 3287 14216 3304
rect 14260 3287 14289 3304
rect 14329 3287 14362 3304
rect 13846 3270 13881 3287
rect 13915 3270 13950 3287
rect 13984 3270 14019 3287
rect 14053 3270 14088 3287
rect 14122 3270 14157 3287
rect 14191 3270 14226 3287
rect 14260 3270 14295 3287
rect 14329 3270 14364 3287
rect 14398 3270 14433 3304
rect 14469 3287 14502 3304
rect 14542 3287 14571 3304
rect 14615 3287 14640 3304
rect 14688 3287 14709 3304
rect 14761 3287 14778 3304
rect 14834 3287 14847 3304
rect 14907 3287 14916 3304
rect 14980 3287 14985 3304
rect 14467 3270 14502 3287
rect 14536 3270 14571 3287
rect 14605 3270 14640 3287
rect 14674 3270 14709 3287
rect 14743 3270 14778 3287
rect 14812 3270 14847 3287
rect 14881 3270 14916 3287
rect 14950 3270 14985 3287
rect 15053 3304 15092 3321
rect 15126 3304 15165 3321
rect 15199 3304 15238 3321
rect 15272 3304 15311 3321
rect 15345 3304 15384 3321
rect 15418 3304 15457 3321
rect 15491 3304 15530 3321
rect 15564 3304 15603 3321
rect 15637 3304 15676 3321
rect 15710 3304 15749 3321
rect 15783 3304 15822 3321
rect 15856 3304 15895 3321
rect 15929 3304 15968 3321
rect 16002 3304 16041 3321
rect 16075 3304 16114 3321
rect 16148 3304 16187 3321
rect 16221 3304 16260 3321
rect 16294 3304 16333 3321
rect 15053 3287 15054 3304
rect 15019 3270 15054 3287
rect 15088 3287 15092 3304
rect 15157 3287 15165 3304
rect 15226 3287 15238 3304
rect 15295 3287 15311 3304
rect 15364 3287 15384 3304
rect 15433 3287 15457 3304
rect 15502 3287 15530 3304
rect 15571 3287 15603 3304
rect 15088 3270 15123 3287
rect 15157 3270 15192 3287
rect 15226 3270 15261 3287
rect 15295 3270 15330 3287
rect 15364 3270 15399 3287
rect 15433 3270 15468 3287
rect 15502 3270 15537 3287
rect 15571 3270 15606 3287
rect 15640 3270 15675 3304
rect 15710 3287 15744 3304
rect 15783 3287 15813 3304
rect 15856 3287 15882 3304
rect 15929 3287 15951 3304
rect 16002 3287 16020 3304
rect 16075 3287 16089 3304
rect 16148 3287 16158 3304
rect 16221 3287 16227 3304
rect 16294 3287 16296 3304
rect 15709 3270 15744 3287
rect 15778 3270 15813 3287
rect 15847 3270 15882 3287
rect 15916 3270 15951 3287
rect 15985 3270 16020 3287
rect 16054 3270 16089 3287
rect 16123 3270 16158 3287
rect 16192 3270 16227 3287
rect 16261 3270 16296 3287
rect 16330 3287 16333 3304
rect 16330 3270 16365 3287
rect 11929 3249 16406 3270
rect 11929 3240 11953 3249
rect 2262 3202 2304 3236
rect 2338 3202 2374 3236
rect 2408 3202 2444 3236
rect 2478 3202 2514 3236
rect 2548 3202 2584 3236
rect 2618 3202 2654 3236
rect 2688 3202 2724 3236
rect 2758 3202 2794 3236
rect 2828 3202 2864 3236
rect 2898 3202 2934 3236
rect 2968 3202 3004 3236
rect 3038 3202 3074 3236
rect 3108 3202 3144 3236
rect 3178 3202 3214 3236
rect 3248 3202 3284 3236
rect 3318 3202 3354 3236
rect 3388 3202 3424 3236
rect 3458 3202 3494 3236
rect 3528 3202 3563 3236
rect 3597 3202 3632 3236
rect 3666 3202 3701 3236
rect 3735 3202 3770 3236
rect 3804 3202 3839 3236
rect 3873 3202 3908 3236
rect 3942 3202 3977 3236
rect 4011 3202 4046 3236
rect 4080 3202 4115 3236
rect 4149 3202 4184 3236
rect 4218 3202 4253 3236
rect 4287 3202 4322 3236
rect 4356 3202 4391 3236
rect 4425 3202 4449 3236
rect 2262 3168 4449 3202
rect -2750 3098 -214 3134
rect -2716 3064 -2680 3098
rect -2646 3064 -2610 3098
rect -2576 3064 -2540 3098
rect -2506 3064 -2470 3098
rect -2436 3064 -2400 3098
rect -2366 3064 -2330 3098
rect -2296 3064 -2260 3098
rect -2226 3064 -2190 3098
rect -2156 3064 -2120 3098
rect -2086 3064 -2050 3098
rect -2016 3064 -1980 3098
rect -1946 3064 -1910 3098
rect -1876 3064 -1840 3098
rect -1806 3064 -1770 3098
rect -1736 3064 -1700 3098
rect -1666 3064 -1630 3098
rect -1596 3064 -1560 3098
rect -1526 3064 -1490 3098
rect -1456 3064 -1421 3098
rect -1387 3064 -1352 3098
rect -1318 3064 -1283 3098
rect -1249 3064 -1214 3098
rect -1180 3064 -1145 3098
rect -1111 3064 -1076 3098
rect -1042 3064 -1007 3098
rect -973 3064 -938 3098
rect -904 3064 -869 3098
rect -835 3064 -800 3098
rect -766 3064 -731 3098
rect -697 3064 -662 3098
rect -628 3064 -593 3098
rect -559 3064 -524 3098
rect -490 3064 -455 3098
rect -421 3064 -386 3098
rect -352 3064 -317 3098
rect -283 3064 -248 3098
rect -2750 3028 -214 3064
rect -2716 2994 -2680 3028
rect -2646 2994 -2610 3028
rect -2576 2994 -2540 3028
rect -2506 2994 -2470 3028
rect -2436 2994 -2400 3028
rect -2366 2994 -2330 3028
rect -2296 2994 -2260 3028
rect -2226 2994 -2190 3028
rect -2156 2994 -2120 3028
rect -2086 2994 -2050 3028
rect -2016 2994 -1980 3028
rect -1946 2994 -1910 3028
rect -1876 2994 -1840 3028
rect -1806 2994 -1770 3028
rect -1736 2994 -1700 3028
rect -1666 2994 -1630 3028
rect -1596 2994 -1560 3028
rect -1526 2994 -1490 3028
rect -1456 2994 -1421 3028
rect -1387 2994 -1352 3028
rect -1318 2994 -1283 3028
rect -1249 2994 -1214 3028
rect -1180 2994 -1145 3028
rect -1111 2994 -1076 3028
rect -1042 2994 -1007 3028
rect -973 2994 -938 3028
rect -904 2994 -869 3028
rect -835 2994 -800 3028
rect -766 2994 -731 3028
rect -697 2994 -662 3028
rect -628 2994 -593 3028
rect -559 2994 -524 3028
rect -490 2994 -455 3028
rect -421 2994 -386 3028
rect -352 2994 -317 3028
rect -283 2994 -248 3028
rect -2750 2958 -214 2994
rect -2716 2924 -2680 2958
rect -2646 2924 -2610 2958
rect -2576 2924 -2540 2958
rect -2506 2924 -2470 2958
rect -2436 2924 -2400 2958
rect -2366 2924 -2330 2958
rect -2296 2924 -2260 2958
rect -2226 2924 -2190 2958
rect -2156 2924 -2120 2958
rect -2086 2924 -2050 2958
rect -2016 2924 -1980 2958
rect -1946 2924 -1910 2958
rect -1876 2924 -1840 2958
rect -1806 2924 -1770 2958
rect -1736 2924 -1700 2958
rect -1666 2924 -1630 2958
rect -1596 2924 -1560 2958
rect -1526 2924 -1490 2958
rect -1456 2924 -1421 2958
rect -1387 2924 -1352 2958
rect -1318 2924 -1283 2958
rect -1249 2924 -1214 2958
rect -1180 2924 -1145 2958
rect -1111 2924 -1076 2958
rect -1042 2924 -1007 2958
rect -973 2924 -938 2958
rect -904 2924 -869 2958
rect -835 2924 -800 2958
rect -766 2924 -731 2958
rect -697 2924 -662 2958
rect -628 2924 -593 2958
rect -559 2924 -524 2958
rect -490 2924 -455 2958
rect -421 2924 -386 2958
rect -352 2924 -317 2958
rect -283 2924 -248 2958
rect -2750 2888 -214 2924
rect -2716 2854 -2680 2888
rect -2646 2854 -2610 2888
rect -2576 2854 -2540 2888
rect -2506 2854 -2470 2888
rect -2436 2854 -2400 2888
rect -2366 2854 -2330 2888
rect -2296 2854 -2260 2888
rect -2226 2854 -2190 2888
rect -2156 2854 -2120 2888
rect -2086 2854 -2050 2888
rect -2016 2854 -1980 2888
rect -1946 2854 -1910 2888
rect -1876 2854 -1840 2888
rect -1806 2854 -1770 2888
rect -1736 2854 -1700 2888
rect -1666 2854 -1630 2888
rect -1596 2854 -1560 2888
rect -1526 2854 -1490 2888
rect -1456 2854 -1421 2888
rect -1387 2854 -1352 2888
rect -1318 2854 -1283 2888
rect -1249 2854 -1214 2888
rect -1180 2854 -1145 2888
rect -1111 2854 -1076 2888
rect -1042 2854 -1007 2888
rect -973 2854 -938 2888
rect -904 2854 -869 2888
rect -835 2854 -800 2888
rect -766 2854 -731 2888
rect -697 2854 -662 2888
rect -628 2854 -593 2888
rect -559 2854 -524 2888
rect -490 2854 -455 2888
rect -421 2854 -386 2888
rect -352 2854 -317 2888
rect -283 2854 -248 2888
rect -2750 2818 -214 2854
rect -2716 2784 -2680 2818
rect -2646 2784 -2610 2818
rect -2576 2784 -2540 2818
rect -2506 2784 -2470 2818
rect -2436 2784 -2400 2818
rect -2366 2784 -2330 2818
rect -2296 2784 -2260 2818
rect -2226 2784 -2190 2818
rect -2156 2784 -2120 2818
rect -2086 2784 -2050 2818
rect -2016 2784 -1980 2818
rect -1946 2784 -1910 2818
rect -1876 2784 -1840 2818
rect -1806 2784 -1770 2818
rect -1736 2784 -1700 2818
rect -1666 2784 -1630 2818
rect -1596 2784 -1560 2818
rect -1526 2784 -1490 2818
rect -1456 2784 -1421 2818
rect -1387 2784 -1352 2818
rect -1318 2784 -1283 2818
rect -1249 2784 -1214 2818
rect -1180 2784 -1145 2818
rect -1111 2784 -1076 2818
rect -1042 2784 -1007 2818
rect -973 2784 -938 2818
rect -904 2784 -869 2818
rect -835 2784 -800 2818
rect -766 2784 -731 2818
rect -697 2784 -662 2818
rect -628 2784 -593 2818
rect -559 2784 -524 2818
rect -490 2784 -455 2818
rect -421 2784 -386 2818
rect -352 2784 -317 2818
rect -283 2784 -248 2818
rect -2750 2748 -214 2784
rect -2716 2714 -2680 2748
rect -2646 2714 -2610 2748
rect -2576 2714 -2540 2748
rect -2506 2714 -2470 2748
rect -2436 2714 -2400 2748
rect -2366 2714 -2330 2748
rect -2296 2714 -2260 2748
rect -2226 2714 -2190 2748
rect -2156 2714 -2120 2748
rect -2086 2714 -2050 2748
rect -2016 2714 -1980 2748
rect -1946 2714 -1910 2748
rect -1876 2714 -1840 2748
rect -1806 2714 -1770 2748
rect -1736 2714 -1700 2748
rect -1666 2714 -1630 2748
rect -1596 2714 -1560 2748
rect -1526 2714 -1490 2748
rect -1456 2714 -1421 2748
rect -1387 2714 -1352 2748
rect -1318 2714 -1283 2748
rect -1249 2714 -1214 2748
rect -1180 2714 -1145 2748
rect -1111 2714 -1076 2748
rect -1042 2714 -1007 2748
rect -973 2714 -938 2748
rect -904 2714 -869 2748
rect -835 2714 -800 2748
rect -766 2714 -731 2748
rect -697 2714 -662 2748
rect -628 2714 -593 2748
rect -559 2714 -524 2748
rect -490 2714 -455 2748
rect -421 2714 -386 2748
rect -352 2714 -317 2748
rect -283 2714 -248 2748
rect -2750 2678 -214 2714
rect -2716 2644 -2680 2678
rect -2646 2644 -2610 2678
rect -2576 2644 -2540 2678
rect -2506 2644 -2470 2678
rect -2436 2644 -2400 2678
rect -2366 2644 -2330 2678
rect -2296 2644 -2260 2678
rect -2226 2644 -2190 2678
rect -2156 2644 -2120 2678
rect -2086 2644 -2050 2678
rect -2016 2644 -1980 2678
rect -1946 2644 -1910 2678
rect -1876 2644 -1840 2678
rect -1806 2644 -1770 2678
rect -1736 2644 -1700 2678
rect -1666 2644 -1630 2678
rect -1596 2644 -1560 2678
rect -1526 2644 -1490 2678
rect -1456 2644 -1421 2678
rect -1387 2644 -1352 2678
rect -1318 2644 -1283 2678
rect -1249 2644 -1214 2678
rect -1180 2644 -1145 2678
rect -1111 2644 -1076 2678
rect -1042 2644 -1007 2678
rect -973 2644 -938 2678
rect -904 2644 -869 2678
rect -835 2644 -800 2678
rect -766 2644 -731 2678
rect -697 2644 -662 2678
rect -628 2644 -593 2678
rect -559 2644 -524 2678
rect -490 2644 -455 2678
rect -421 2644 -386 2678
rect -352 2644 -317 2678
rect -283 2644 -248 2678
rect -2750 2608 -214 2644
rect -2716 2574 -2680 2608
rect -2646 2574 -2610 2608
rect -2576 2574 -2540 2608
rect -2506 2574 -2470 2608
rect -2436 2574 -2400 2608
rect -2366 2574 -2330 2608
rect -2296 2574 -2260 2608
rect -2226 2574 -2190 2608
rect -2156 2574 -2120 2608
rect -2086 2574 -2050 2608
rect -2016 2574 -1980 2608
rect -1946 2574 -1910 2608
rect -1876 2574 -1840 2608
rect -1806 2574 -1770 2608
rect -1736 2574 -1700 2608
rect -1666 2574 -1630 2608
rect -1596 2574 -1560 2608
rect -1526 2574 -1490 2608
rect -1456 2574 -1421 2608
rect -1387 2574 -1352 2608
rect -1318 2574 -1283 2608
rect -1249 2574 -1214 2608
rect -1180 2574 -1145 2608
rect -1111 2574 -1076 2608
rect -1042 2574 -1007 2608
rect -973 2574 -938 2608
rect -904 2574 -869 2608
rect -835 2574 -800 2608
rect -766 2574 -731 2608
rect -697 2574 -662 2608
rect -628 2574 -593 2608
rect -559 2574 -524 2608
rect -490 2574 -455 2608
rect -421 2574 -386 2608
rect -352 2574 -317 2608
rect -283 2574 -248 2608
rect -2750 2538 -214 2574
rect -2716 2504 -2680 2538
rect -2646 2504 -2610 2538
rect -2576 2504 -2540 2538
rect -2506 2504 -2470 2538
rect -2436 2504 -2400 2538
rect -2366 2504 -2330 2538
rect -2296 2504 -2260 2538
rect -2226 2504 -2190 2538
rect -2156 2504 -2120 2538
rect -2086 2504 -2050 2538
rect -2016 2504 -1980 2538
rect -1946 2504 -1910 2538
rect -1876 2504 -1840 2538
rect -1806 2504 -1770 2538
rect -1736 2504 -1700 2538
rect -1666 2504 -1630 2538
rect -1596 2504 -1560 2538
rect -1526 2504 -1490 2538
rect -1456 2504 -1421 2538
rect -1387 2504 -1352 2538
rect -1318 2504 -1283 2538
rect -1249 2504 -1214 2538
rect -1180 2504 -1145 2538
rect -1111 2504 -1076 2538
rect -1042 2504 -1007 2538
rect -973 2504 -938 2538
rect -904 2504 -869 2538
rect -835 2504 -800 2538
rect -766 2504 -731 2538
rect -697 2504 -662 2538
rect -628 2504 -593 2538
rect -559 2504 -524 2538
rect -490 2504 -455 2538
rect -421 2504 -386 2538
rect -352 2504 -317 2538
rect -283 2504 -248 2538
rect -2750 2468 -214 2504
rect -2716 2434 -2680 2468
rect -2646 2434 -2610 2468
rect -2576 2434 -2540 2468
rect -2506 2434 -2470 2468
rect -2436 2434 -2400 2468
rect -2366 2434 -2330 2468
rect -2296 2434 -2260 2468
rect -2226 2434 -2190 2468
rect -2156 2434 -2120 2468
rect -2086 2434 -2050 2468
rect -2016 2434 -1980 2468
rect -1946 2434 -1910 2468
rect -1876 2434 -1840 2468
rect -1806 2434 -1770 2468
rect -1736 2434 -1700 2468
rect -1666 2434 -1630 2468
rect -1596 2434 -1560 2468
rect -1526 2434 -1490 2468
rect -1456 2434 -1421 2468
rect -1387 2434 -1352 2468
rect -1318 2434 -1283 2468
rect -1249 2434 -1214 2468
rect -1180 2434 -1145 2468
rect -1111 2434 -1076 2468
rect -1042 2434 -1007 2468
rect -973 2434 -938 2468
rect -904 2434 -869 2468
rect -835 2434 -800 2468
rect -766 2434 -731 2468
rect -697 2434 -662 2468
rect -628 2434 -593 2468
rect -559 2434 -524 2468
rect -490 2434 -455 2468
rect -421 2434 -386 2468
rect -352 2434 -317 2468
rect -283 2434 -248 2468
rect -2750 2398 -214 2434
rect -2716 2364 -2680 2398
rect -2646 2364 -2610 2398
rect -2576 2364 -2540 2398
rect -2506 2364 -2470 2398
rect -2436 2364 -2400 2398
rect -2366 2364 -2330 2398
rect -2296 2364 -2260 2398
rect -2226 2364 -2190 2398
rect -2156 2364 -2120 2398
rect -2086 2364 -2050 2398
rect -2016 2364 -1980 2398
rect -1946 2364 -1910 2398
rect -1876 2364 -1840 2398
rect -1806 2364 -1770 2398
rect -1736 2364 -1700 2398
rect -1666 2364 -1630 2398
rect -1596 2364 -1560 2398
rect -1526 2364 -1490 2398
rect -1456 2364 -1421 2398
rect -1387 2364 -1352 2398
rect -1318 2364 -1283 2398
rect -1249 2364 -1214 2398
rect -1180 2364 -1145 2398
rect -1111 2364 -1076 2398
rect -1042 2364 -1007 2398
rect -973 2364 -938 2398
rect -904 2364 -869 2398
rect -835 2364 -800 2398
rect -766 2364 -731 2398
rect -697 2364 -662 2398
rect -628 2364 -593 2398
rect -559 2364 -524 2398
rect -490 2364 -455 2398
rect -421 2364 -386 2398
rect -352 2364 -317 2398
rect -283 2364 -248 2398
rect -2750 2328 -214 2364
rect -2716 2294 -2680 2328
rect -2646 2294 -2610 2328
rect -2576 2294 -2540 2328
rect -2506 2294 -2470 2328
rect -2436 2294 -2400 2328
rect -2366 2294 -2330 2328
rect -2296 2294 -2260 2328
rect -2226 2294 -2190 2328
rect -2156 2294 -2120 2328
rect -2086 2294 -2050 2328
rect -2016 2294 -1980 2328
rect -1946 2294 -1910 2328
rect -1876 2294 -1840 2328
rect -1806 2294 -1770 2328
rect -1736 2294 -1700 2328
rect -1666 2294 -1630 2328
rect -1596 2294 -1560 2328
rect -1526 2294 -1490 2328
rect -1456 2294 -1421 2328
rect -1387 2294 -1352 2328
rect -1318 2294 -1283 2328
rect -1249 2294 -1214 2328
rect -1180 2294 -1145 2328
rect -1111 2294 -1076 2328
rect -1042 2294 -1007 2328
rect -973 2294 -938 2328
rect -904 2294 -869 2328
rect -835 2294 -800 2328
rect -766 2294 -731 2328
rect -697 2294 -662 2328
rect -628 2294 -593 2328
rect -559 2294 -524 2328
rect -490 2294 -455 2328
rect -421 2294 -386 2328
rect -352 2294 -317 2328
rect -283 2294 -248 2328
rect -2750 2236 -214 2294
rect -163 3140 307 3164
rect -163 3106 -161 3140
rect -127 3106 -89 3140
rect -55 3106 -17 3140
rect 17 3106 55 3140
rect 89 3106 127 3140
rect 161 3106 199 3140
rect 233 3106 271 3140
rect 305 3106 307 3140
rect -163 3071 307 3106
rect -163 3037 -161 3071
rect -127 3037 -89 3071
rect -55 3037 -17 3071
rect 17 3037 55 3071
rect 89 3037 127 3071
rect 161 3037 199 3071
rect 233 3037 271 3071
rect 305 3037 307 3071
rect -163 3002 307 3037
rect -163 2968 -161 3002
rect -127 2968 -89 3002
rect -55 2968 -17 3002
rect 17 2968 55 3002
rect 89 2968 127 3002
rect 161 2968 199 3002
rect 233 2968 271 3002
rect 305 2968 307 3002
rect -163 2933 307 2968
rect -163 2899 -161 2933
rect -127 2899 -89 2933
rect -55 2899 -17 2933
rect 17 2899 55 2933
rect 89 2899 127 2933
rect 161 2899 199 2933
rect 233 2899 271 2933
rect 305 2899 307 2933
rect -163 2863 307 2899
rect -163 2829 -161 2863
rect -127 2829 -89 2863
rect -55 2829 -17 2863
rect 17 2829 55 2863
rect 89 2829 127 2863
rect 161 2829 199 2863
rect 233 2829 271 2863
rect 305 2829 307 2863
rect -163 2793 307 2829
rect -163 2759 -161 2793
rect -127 2759 -89 2793
rect -55 2759 -17 2793
rect 17 2759 55 2793
rect 89 2759 127 2793
rect 161 2759 199 2793
rect 233 2759 271 2793
rect 305 2759 307 2793
rect -163 2723 307 2759
rect -163 2689 -161 2723
rect -127 2689 -89 2723
rect -55 2689 -17 2723
rect 17 2689 55 2723
rect 89 2689 127 2723
rect 161 2689 199 2723
rect 233 2689 271 2723
rect 305 2689 307 2723
rect -163 2653 307 2689
rect -163 2619 -161 2653
rect -127 2619 -89 2653
rect -55 2619 -17 2653
rect 17 2619 55 2653
rect 89 2619 127 2653
rect 161 2619 199 2653
rect 233 2619 271 2653
rect 305 2619 307 2653
rect -163 2583 307 2619
rect -163 2549 -161 2583
rect -127 2549 -89 2583
rect -55 2549 -17 2583
rect 17 2549 55 2583
rect 89 2549 127 2583
rect 161 2549 199 2583
rect 233 2549 271 2583
rect 305 2549 307 2583
rect -163 2513 307 2549
rect -163 2479 -161 2513
rect -127 2479 -89 2513
rect -55 2479 -17 2513
rect 17 2479 55 2513
rect 89 2479 127 2513
rect 161 2479 199 2513
rect 233 2479 271 2513
rect 305 2479 307 2513
rect -163 2443 307 2479
rect -163 2409 -161 2443
rect -127 2409 -89 2443
rect -55 2409 -17 2443
rect 17 2409 55 2443
rect 89 2409 127 2443
rect 161 2409 199 2443
rect 233 2409 271 2443
rect 305 2409 307 2443
rect -163 2373 307 2409
rect -163 2339 -161 2373
rect -127 2339 -89 2373
rect -55 2339 -17 2373
rect 17 2339 55 2373
rect 89 2339 127 2373
rect 161 2339 199 2373
rect 233 2339 271 2373
rect 305 2339 307 2373
rect -163 2303 307 2339
rect -163 2269 -161 2303
rect -127 2269 -89 2303
rect -55 2269 -17 2303
rect 17 2269 55 2303
rect 89 2269 127 2303
rect 161 2269 199 2303
rect 233 2269 271 2303
rect 305 2269 307 2303
rect -163 2245 307 2269
rect 2262 3134 2304 3168
rect 2338 3134 2374 3168
rect 2408 3134 2444 3168
rect 2478 3134 2514 3168
rect 2548 3134 2584 3168
rect 2618 3134 2654 3168
rect 2688 3134 2724 3168
rect 2758 3134 2794 3168
rect 2828 3134 2864 3168
rect 2898 3134 2934 3168
rect 2968 3134 3004 3168
rect 3038 3134 3074 3168
rect 3108 3134 3144 3168
rect 3178 3134 3214 3168
rect 3248 3134 3284 3168
rect 3318 3134 3354 3168
rect 3388 3134 3424 3168
rect 3458 3134 3494 3168
rect 3528 3134 3563 3168
rect 3597 3134 3632 3168
rect 3666 3134 3701 3168
rect 3735 3134 3770 3168
rect 3804 3134 3839 3168
rect 3873 3134 3908 3168
rect 3942 3134 3977 3168
rect 4011 3134 4046 3168
rect 4080 3134 4115 3168
rect 4149 3134 4184 3168
rect 4218 3134 4253 3168
rect 4287 3134 4322 3168
rect 4356 3134 4391 3168
rect 4425 3134 4449 3168
rect 2262 3100 4449 3134
rect 2262 3066 2304 3100
rect 2338 3066 2374 3100
rect 2408 3066 2444 3100
rect 2478 3066 2514 3100
rect 2548 3066 2584 3100
rect 2618 3066 2654 3100
rect 2688 3066 2724 3100
rect 2758 3066 2794 3100
rect 2828 3066 2864 3100
rect 2898 3066 2934 3100
rect 2968 3066 3004 3100
rect 3038 3066 3074 3100
rect 3108 3066 3144 3100
rect 3178 3066 3214 3100
rect 3248 3066 3284 3100
rect 3318 3066 3354 3100
rect 3388 3066 3424 3100
rect 3458 3066 3494 3100
rect 3528 3066 3563 3100
rect 3597 3066 3632 3100
rect 3666 3066 3701 3100
rect 3735 3066 3770 3100
rect 3804 3066 3839 3100
rect 3873 3066 3908 3100
rect 3942 3066 3977 3100
rect 4011 3066 4046 3100
rect 4080 3066 4115 3100
rect 4149 3066 4184 3100
rect 4218 3066 4253 3100
rect 4287 3066 4322 3100
rect 4356 3066 4391 3100
rect 4425 3066 4449 3100
rect 2262 3032 4449 3066
rect 2262 2998 2304 3032
rect 2338 2998 2374 3032
rect 2408 2998 2444 3032
rect 2478 2998 2514 3032
rect 2548 2998 2584 3032
rect 2618 2998 2654 3032
rect 2688 2998 2724 3032
rect 2758 2998 2794 3032
rect 2828 2998 2864 3032
rect 2898 2998 2934 3032
rect 2968 2998 3004 3032
rect 3038 2998 3074 3032
rect 3108 2998 3144 3032
rect 3178 2998 3214 3032
rect 3248 2998 3284 3032
rect 3318 2998 3354 3032
rect 3388 2998 3424 3032
rect 3458 2998 3494 3032
rect 3528 2998 3563 3032
rect 3597 2998 3632 3032
rect 3666 2998 3701 3032
rect 3735 2998 3770 3032
rect 3804 2998 3839 3032
rect 3873 2998 3908 3032
rect 3942 2998 3977 3032
rect 4011 2998 4046 3032
rect 4080 2998 4115 3032
rect 4149 2998 4184 3032
rect 4218 2998 4253 3032
rect 4287 2998 4322 3032
rect 4356 2998 4391 3032
rect 4425 2998 4449 3032
rect 2262 2964 4449 2998
rect 2262 2930 2304 2964
rect 2338 2930 2374 2964
rect 2408 2930 2444 2964
rect 2478 2930 2514 2964
rect 2548 2930 2584 2964
rect 2618 2930 2654 2964
rect 2688 2930 2724 2964
rect 2758 2930 2794 2964
rect 2828 2930 2864 2964
rect 2898 2930 2934 2964
rect 2968 2930 3004 2964
rect 3038 2930 3074 2964
rect 3108 2930 3144 2964
rect 3178 2930 3214 2964
rect 3248 2930 3284 2964
rect 3318 2930 3354 2964
rect 3388 2930 3424 2964
rect 3458 2930 3494 2964
rect 3528 2930 3563 2964
rect 3597 2930 3632 2964
rect 3666 2930 3701 2964
rect 3735 2930 3770 2964
rect 3804 2930 3839 2964
rect 3873 2930 3908 2964
rect 3942 2930 3977 2964
rect 4011 2930 4046 2964
rect 4080 2930 4115 2964
rect 4149 2930 4184 2964
rect 4218 2930 4253 2964
rect 4287 2930 4322 2964
rect 4356 2930 4391 2964
rect 4425 2930 4449 2964
rect 2262 2896 4449 2930
rect 2262 2862 2304 2896
rect 2338 2862 2374 2896
rect 2408 2862 2444 2896
rect 2478 2862 2514 2896
rect 2548 2862 2584 2896
rect 2618 2862 2654 2896
rect 2688 2862 2724 2896
rect 2758 2862 2794 2896
rect 2828 2862 2864 2896
rect 2898 2862 2934 2896
rect 2968 2862 3004 2896
rect 3038 2862 3074 2896
rect 3108 2862 3144 2896
rect 3178 2862 3214 2896
rect 3248 2862 3284 2896
rect 3318 2862 3354 2896
rect 3388 2862 3424 2896
rect 3458 2862 3494 2896
rect 3528 2862 3563 2896
rect 3597 2862 3632 2896
rect 3666 2862 3701 2896
rect 3735 2862 3770 2896
rect 3804 2862 3839 2896
rect 3873 2862 3908 2896
rect 3942 2862 3977 2896
rect 4011 2862 4046 2896
rect 4080 2862 4115 2896
rect 4149 2862 4184 2896
rect 4218 2862 4253 2896
rect 4287 2862 4322 2896
rect 4356 2862 4391 2896
rect 4425 2862 4449 2896
rect 2262 2828 4449 2862
rect 2262 2794 2304 2828
rect 2338 2794 2374 2828
rect 2408 2794 2444 2828
rect 2478 2794 2514 2828
rect 2548 2794 2584 2828
rect 2618 2794 2654 2828
rect 2688 2794 2724 2828
rect 2758 2794 2794 2828
rect 2828 2794 2864 2828
rect 2898 2794 2934 2828
rect 2968 2794 3004 2828
rect 3038 2794 3074 2828
rect 3108 2794 3144 2828
rect 3178 2794 3214 2828
rect 3248 2794 3284 2828
rect 3318 2794 3354 2828
rect 3388 2794 3424 2828
rect 3458 2794 3494 2828
rect 3528 2794 3563 2828
rect 3597 2794 3632 2828
rect 3666 2794 3701 2828
rect 3735 2794 3770 2828
rect 3804 2794 3839 2828
rect 3873 2794 3908 2828
rect 3942 2794 3977 2828
rect 4011 2794 4046 2828
rect 4080 2794 4115 2828
rect 4149 2794 4184 2828
rect 4218 2794 4253 2828
rect 4287 2794 4322 2828
rect 4356 2794 4391 2828
rect 4425 2794 4449 2828
rect 2262 2760 4449 2794
rect 2262 2726 2304 2760
rect 2338 2726 2374 2760
rect 2408 2726 2444 2760
rect 2478 2726 2514 2760
rect 2548 2726 2584 2760
rect 2618 2726 2654 2760
rect 2688 2726 2724 2760
rect 2758 2726 2794 2760
rect 2828 2726 2864 2760
rect 2898 2726 2934 2760
rect 2968 2726 3004 2760
rect 3038 2726 3074 2760
rect 3108 2726 3144 2760
rect 3178 2726 3214 2760
rect 3248 2726 3284 2760
rect 3318 2726 3354 2760
rect 3388 2726 3424 2760
rect 3458 2726 3494 2760
rect 3528 2726 3563 2760
rect 3597 2726 3632 2760
rect 3666 2726 3701 2760
rect 3735 2726 3770 2760
rect 3804 2726 3839 2760
rect 3873 2726 3908 2760
rect 3942 2726 3977 2760
rect 4011 2726 4046 2760
rect 4080 2726 4115 2760
rect 4149 2726 4184 2760
rect 4218 2726 4253 2760
rect 4287 2726 4322 2760
rect 4356 2726 4391 2760
rect 4425 2726 4449 2760
rect 2262 2692 4449 2726
rect 2262 2658 2304 2692
rect 2338 2658 2374 2692
rect 2408 2658 2444 2692
rect 2478 2658 2514 2692
rect 2548 2658 2584 2692
rect 2618 2658 2654 2692
rect 2688 2658 2724 2692
rect 2758 2658 2794 2692
rect 2828 2658 2864 2692
rect 2898 2658 2934 2692
rect 2968 2658 3004 2692
rect 3038 2658 3074 2692
rect 3108 2658 3144 2692
rect 3178 2658 3214 2692
rect 3248 2658 3284 2692
rect 3318 2658 3354 2692
rect 3388 2658 3424 2692
rect 3458 2658 3494 2692
rect 3528 2658 3563 2692
rect 3597 2658 3632 2692
rect 3666 2658 3701 2692
rect 3735 2658 3770 2692
rect 3804 2658 3839 2692
rect 3873 2658 3908 2692
rect 3942 2658 3977 2692
rect 4011 2658 4046 2692
rect 4080 2658 4115 2692
rect 4149 2658 4184 2692
rect 4218 2658 4253 2692
rect 4287 2658 4322 2692
rect 4356 2658 4391 2692
rect 4425 2658 4449 2692
rect 2262 2624 4449 2658
rect 2262 2590 2304 2624
rect 2338 2590 2374 2624
rect 2408 2590 2444 2624
rect 2478 2590 2514 2624
rect 2548 2590 2584 2624
rect 2618 2590 2654 2624
rect 2688 2590 2724 2624
rect 2758 2590 2794 2624
rect 2828 2590 2864 2624
rect 2898 2590 2934 2624
rect 2968 2590 3004 2624
rect 3038 2590 3074 2624
rect 3108 2590 3144 2624
rect 3178 2590 3214 2624
rect 3248 2590 3284 2624
rect 3318 2590 3354 2624
rect 3388 2590 3424 2624
rect 3458 2590 3494 2624
rect 3528 2590 3563 2624
rect 3597 2590 3632 2624
rect 3666 2590 3701 2624
rect 3735 2590 3770 2624
rect 3804 2590 3839 2624
rect 3873 2590 3908 2624
rect 3942 2590 3977 2624
rect 4011 2590 4046 2624
rect 4080 2590 4115 2624
rect 4149 2590 4184 2624
rect 4218 2590 4253 2624
rect 4287 2590 4322 2624
rect 4356 2590 4391 2624
rect 4425 2590 4449 2624
rect 2262 2556 4449 2590
rect 2262 2522 2304 2556
rect 2338 2522 2374 2556
rect 2408 2522 2444 2556
rect 2478 2522 2514 2556
rect 2548 2522 2584 2556
rect 2618 2522 2654 2556
rect 2688 2522 2724 2556
rect 2758 2522 2794 2556
rect 2828 2522 2864 2556
rect 2898 2522 2934 2556
rect 2968 2522 3004 2556
rect 3038 2522 3074 2556
rect 3108 2522 3144 2556
rect 3178 2522 3214 2556
rect 3248 2522 3284 2556
rect 3318 2522 3354 2556
rect 3388 2522 3424 2556
rect 3458 2522 3494 2556
rect 3528 2522 3563 2556
rect 3597 2522 3632 2556
rect 3666 2522 3701 2556
rect 3735 2522 3770 2556
rect 3804 2522 3839 2556
rect 3873 2522 3908 2556
rect 3942 2522 3977 2556
rect 4011 2522 4046 2556
rect 4080 2522 4115 2556
rect 4149 2522 4184 2556
rect 4218 2522 4253 2556
rect 4287 2522 4322 2556
rect 4356 2522 4391 2556
rect 4425 2522 4449 2556
rect 2262 2488 4449 2522
rect 2262 2454 2304 2488
rect 2338 2454 2374 2488
rect 2408 2454 2444 2488
rect 2478 2454 2514 2488
rect 2548 2454 2584 2488
rect 2618 2454 2654 2488
rect 2688 2454 2724 2488
rect 2758 2454 2794 2488
rect 2828 2454 2864 2488
rect 2898 2454 2934 2488
rect 2968 2454 3004 2488
rect 3038 2454 3074 2488
rect 3108 2454 3144 2488
rect 3178 2454 3214 2488
rect 3248 2454 3284 2488
rect 3318 2454 3354 2488
rect 3388 2454 3424 2488
rect 3458 2454 3494 2488
rect 3528 2454 3563 2488
rect 3597 2454 3632 2488
rect 3666 2454 3701 2488
rect 3735 2454 3770 2488
rect 3804 2454 3839 2488
rect 3873 2454 3908 2488
rect 3942 2454 3977 2488
rect 4011 2454 4046 2488
rect 4080 2454 4115 2488
rect 4149 2454 4184 2488
rect 4218 2454 4253 2488
rect 4287 2454 4322 2488
rect 4356 2454 4391 2488
rect 4425 2454 4449 2488
rect 2262 2420 4449 2454
rect 2262 2386 2304 2420
rect 2338 2386 2374 2420
rect 2408 2386 2444 2420
rect 2478 2386 2514 2420
rect 2548 2386 2584 2420
rect 2618 2386 2654 2420
rect 2688 2386 2724 2420
rect 2758 2386 2794 2420
rect 2828 2386 2864 2420
rect 2898 2386 2934 2420
rect 2968 2386 3004 2420
rect 3038 2386 3074 2420
rect 3108 2386 3144 2420
rect 3178 2386 3214 2420
rect 3248 2386 3284 2420
rect 3318 2386 3354 2420
rect 3388 2386 3424 2420
rect 3458 2386 3494 2420
rect 3528 2386 3563 2420
rect 3597 2386 3632 2420
rect 3666 2386 3701 2420
rect 3735 2386 3770 2420
rect 3804 2386 3839 2420
rect 3873 2386 3908 2420
rect 3942 2386 3977 2420
rect 4011 2386 4046 2420
rect 4080 2386 4115 2420
rect 4149 2386 4184 2420
rect 4218 2386 4253 2420
rect 4287 2386 4322 2420
rect 4356 2386 4391 2420
rect 4425 2386 4449 2420
rect 2262 2352 4449 2386
rect 2262 2318 2304 2352
rect 2338 2318 2374 2352
rect 2408 2318 2444 2352
rect 2478 2318 2514 2352
rect 2548 2318 2584 2352
rect 2618 2318 2654 2352
rect 2688 2318 2724 2352
rect 2758 2318 2794 2352
rect 2828 2318 2864 2352
rect 2898 2318 2934 2352
rect 2968 2318 3004 2352
rect 3038 2318 3074 2352
rect 3108 2318 3144 2352
rect 3178 2318 3214 2352
rect 3248 2318 3284 2352
rect 3318 2318 3354 2352
rect 3388 2318 3424 2352
rect 3458 2318 3494 2352
rect 3528 2318 3563 2352
rect 3597 2318 3632 2352
rect 3666 2318 3701 2352
rect 3735 2318 3770 2352
rect 3804 2318 3839 2352
rect 3873 2318 3908 2352
rect 3942 2318 3977 2352
rect 4011 2318 4046 2352
rect 4080 2318 4115 2352
rect 4149 2318 4184 2352
rect 4218 2318 4253 2352
rect 4287 2318 4322 2352
rect 4356 2318 4391 2352
rect 4425 2318 4449 2352
rect 2262 2284 4449 2318
rect 2262 2250 2304 2284
rect 2338 2250 2374 2284
rect 2408 2250 2444 2284
rect 2478 2250 2514 2284
rect 2548 2250 2584 2284
rect 2618 2250 2654 2284
rect 2688 2250 2724 2284
rect 2758 2250 2794 2284
rect 2828 2250 2864 2284
rect 2898 2250 2934 2284
rect 2968 2250 3004 2284
rect 3038 2250 3074 2284
rect 3108 2250 3144 2284
rect 3178 2250 3214 2284
rect 3248 2250 3284 2284
rect 3318 2250 3354 2284
rect 3388 2250 3424 2284
rect 3458 2250 3494 2284
rect 3528 2250 3563 2284
rect 3597 2250 3632 2284
rect 3666 2250 3701 2284
rect 3735 2250 3770 2284
rect 3804 2250 3839 2284
rect 3873 2250 3908 2284
rect 3942 2250 3977 2284
rect 4011 2250 4046 2284
rect 4080 2250 4115 2284
rect 4149 2250 4184 2284
rect 4218 2250 4253 2284
rect 4287 2250 4322 2284
rect 4356 2250 4391 2284
rect 4425 2250 4449 2284
rect 2262 2193 4449 2250
rect -2750 2159 -2726 2193
rect -2692 2159 -2656 2193
rect -2622 2159 -2586 2193
rect -2552 2159 -2517 2193
rect -2483 2159 -2448 2193
rect -2414 2159 -2379 2193
rect -2345 2159 -2310 2193
rect -2276 2159 -2241 2193
rect -2207 2159 -2172 2193
rect -2138 2159 -2103 2193
rect -2069 2159 -2034 2193
rect -2000 2159 -1965 2193
rect -1931 2159 -1896 2193
rect -1862 2159 -1827 2193
rect -1793 2159 -1758 2193
rect -1724 2159 -1689 2193
rect -1655 2159 -1620 2193
rect -1586 2159 -1551 2193
rect -1517 2159 -1482 2193
rect -1448 2159 -1413 2193
rect -1379 2159 -1344 2193
rect -1310 2159 -1275 2193
rect -1241 2159 -1206 2193
rect -1172 2159 -1137 2193
rect -1103 2159 -1068 2193
rect -1034 2159 -999 2193
rect -965 2159 -930 2193
rect -896 2159 -861 2193
rect -827 2159 -792 2193
rect -758 2159 -723 2193
rect -689 2159 -654 2193
rect -620 2159 -585 2193
rect -551 2159 -516 2193
rect -482 2159 -447 2193
rect -413 2159 -378 2193
rect -344 2159 -309 2193
rect -275 2159 -240 2193
rect -206 2159 -171 2193
rect -137 2159 -102 2193
rect -68 2159 -33 2193
rect 1 2159 36 2193
rect 70 2159 105 2193
rect 139 2159 174 2193
rect 208 2159 243 2193
rect 277 2159 301 2193
rect 2262 2177 2298 2193
rect -2750 2125 301 2159
rect -2750 2091 -2726 2125
rect -2692 2091 -2656 2125
rect -2622 2091 -2586 2125
rect -2552 2091 -2517 2125
rect -2483 2091 -2448 2125
rect -2414 2091 -2379 2125
rect -2345 2091 -2310 2125
rect -2276 2091 -2241 2125
rect -2207 2091 -2172 2125
rect -2138 2091 -2103 2125
rect -2069 2091 -2034 2125
rect -2000 2091 -1965 2125
rect -1931 2091 -1896 2125
rect -1862 2091 -1827 2125
rect -1793 2091 -1758 2125
rect -1724 2091 -1689 2125
rect -1655 2091 -1620 2125
rect -1586 2091 -1551 2125
rect -1517 2091 -1482 2125
rect -1448 2091 -1413 2125
rect -1379 2091 -1344 2125
rect -1310 2091 -1275 2125
rect -1241 2091 -1206 2125
rect -1172 2091 -1137 2125
rect -1103 2091 -1068 2125
rect -1034 2091 -999 2125
rect -965 2091 -930 2125
rect -896 2091 -861 2125
rect -827 2091 -792 2125
rect -758 2091 -723 2125
rect -689 2091 -654 2125
rect -620 2091 -585 2125
rect -551 2091 -516 2125
rect -482 2091 -447 2125
rect -413 2091 -378 2125
rect -344 2091 -309 2125
rect -275 2091 -240 2125
rect -206 2091 -171 2125
rect -137 2091 -102 2125
rect -68 2091 -33 2125
rect 1 2091 36 2125
rect 70 2091 105 2125
rect 139 2091 174 2125
rect 208 2091 243 2125
rect 277 2091 301 2125
rect -2750 2057 301 2091
rect -2750 2023 -2726 2057
rect -2692 2023 -2656 2057
rect -2622 2023 -2586 2057
rect -2552 2023 -2517 2057
rect -2483 2023 -2448 2057
rect -2414 2023 -2379 2057
rect -2345 2023 -2310 2057
rect -2276 2023 -2241 2057
rect -2207 2023 -2172 2057
rect -2138 2023 -2103 2057
rect -2069 2023 -2034 2057
rect -2000 2023 -1965 2057
rect -1931 2023 -1896 2057
rect -1862 2023 -1827 2057
rect -1793 2023 -1758 2057
rect -1724 2023 -1689 2057
rect -1655 2023 -1620 2057
rect -1586 2023 -1551 2057
rect -1517 2023 -1482 2057
rect -1448 2023 -1413 2057
rect -1379 2023 -1344 2057
rect -1310 2023 -1275 2057
rect -1241 2023 -1206 2057
rect -1172 2023 -1137 2057
rect -1103 2023 -1068 2057
rect -1034 2023 -999 2057
rect -965 2023 -930 2057
rect -896 2023 -861 2057
rect -827 2023 -792 2057
rect -758 2023 -723 2057
rect -689 2023 -654 2057
rect -620 2023 -585 2057
rect -551 2023 -516 2057
rect -482 2023 -447 2057
rect -413 2023 -378 2057
rect -344 2023 -309 2057
rect -275 2023 -240 2057
rect -206 2023 -171 2057
rect -137 2023 -102 2057
rect -68 2023 -33 2057
rect 1 2023 36 2057
rect 70 2023 105 2057
rect 139 2023 174 2057
rect 208 2023 243 2057
rect 277 2023 301 2057
rect 403 2159 2298 2177
rect 2332 2159 2368 2193
rect 2402 2159 2438 2193
rect 2472 2159 2508 2193
rect 2542 2159 2578 2193
rect 2612 2159 2648 2193
rect 2682 2159 2718 2193
rect 2752 2159 2788 2193
rect 2822 2159 2858 2193
rect 2892 2159 2928 2193
rect 2962 2159 2998 2193
rect 3032 2159 3068 2193
rect 3102 2159 3138 2193
rect 3172 2159 3208 2193
rect 3242 2159 3278 2193
rect 3312 2159 3348 2193
rect 3382 2159 3418 2193
rect 3452 2159 3488 2193
rect 3522 2159 3558 2193
rect 3592 2159 3628 2193
rect 3662 2159 3698 2193
rect 3732 2159 3768 2193
rect 3802 2159 3838 2193
rect 3872 2159 3908 2193
rect 3942 2159 3977 2193
rect 4011 2159 4046 2193
rect 4080 2159 4115 2193
rect 4149 2159 4184 2193
rect 4218 2159 4253 2193
rect 4287 2159 4322 2193
rect 4356 2159 4391 2193
rect 4425 2159 4449 2193
rect 403 2125 4449 2159
rect 403 2091 2298 2125
rect 2332 2091 2368 2125
rect 2402 2091 2438 2125
rect 2472 2091 2508 2125
rect 2542 2091 2578 2125
rect 2612 2091 2648 2125
rect 2682 2091 2718 2125
rect 2752 2091 2788 2125
rect 2822 2091 2858 2125
rect 2892 2091 2928 2125
rect 2962 2091 2998 2125
rect 3032 2091 3068 2125
rect 3102 2091 3138 2125
rect 3172 2091 3208 2125
rect 3242 2091 3278 2125
rect 3312 2091 3348 2125
rect 3382 2091 3418 2125
rect 3452 2091 3488 2125
rect 3522 2091 3558 2125
rect 3592 2091 3628 2125
rect 3662 2091 3698 2125
rect 3732 2091 3768 2125
rect 3802 2091 3838 2125
rect 3872 2091 3908 2125
rect 3942 2091 3977 2125
rect 4011 2091 4046 2125
rect 4080 2091 4115 2125
rect 4149 2091 4184 2125
rect 4218 2091 4253 2125
rect 4287 2091 4322 2125
rect 4356 2091 4391 2125
rect 4425 2091 4449 2125
rect 403 2057 4449 2091
rect 403 2023 2298 2057
rect 2332 2023 2368 2057
rect 2402 2023 2438 2057
rect 2472 2023 2508 2057
rect 2542 2023 2578 2057
rect 2612 2023 2648 2057
rect 2682 2023 2718 2057
rect 2752 2023 2788 2057
rect 2822 2023 2858 2057
rect 2892 2023 2928 2057
rect 2962 2023 2998 2057
rect 3032 2023 3068 2057
rect 3102 2023 3138 2057
rect 3172 2023 3208 2057
rect 3242 2023 3278 2057
rect 3312 2023 3348 2057
rect 3382 2023 3418 2057
rect 3452 2023 3488 2057
rect 3522 2023 3558 2057
rect 3592 2023 3628 2057
rect 3662 2023 3698 2057
rect 3732 2023 3768 2057
rect 3802 2023 3838 2057
rect 3872 2023 3908 2057
rect 3942 2023 3977 2057
rect 4011 2023 4046 2057
rect 4080 2023 4115 2057
rect 4149 2023 4184 2057
rect 4218 2023 4253 2057
rect 4287 2023 4322 2057
rect 4356 2023 4391 2057
rect 4425 2023 4449 2057
rect 4615 3235 11953 3240
rect 11987 3235 12026 3249
rect 12060 3235 12099 3249
rect 12133 3235 12172 3249
rect 12206 3235 12245 3249
rect 12279 3235 12318 3249
rect 12352 3235 12391 3249
rect 12425 3235 12464 3249
rect 12498 3235 12537 3249
rect 12571 3235 12610 3249
rect 12644 3235 12683 3249
rect 12717 3235 12756 3249
rect 12790 3235 12829 3249
rect 12863 3235 12902 3249
rect 12936 3235 12975 3249
rect 13009 3235 13048 3249
rect 13082 3235 13121 3249
rect 13155 3235 13194 3249
rect 13228 3235 13267 3249
rect 13301 3235 13340 3249
rect 13374 3235 13413 3249
rect 13447 3235 13486 3249
rect 13520 3235 13559 3249
rect 13593 3235 13632 3249
rect 13666 3235 13705 3249
rect 13739 3235 13778 3249
rect 13812 3235 13851 3249
rect 13885 3235 13924 3249
rect 13958 3235 13997 3249
rect 14031 3235 14070 3249
rect 14104 3235 14143 3249
rect 14177 3235 14216 3249
rect 14250 3235 14289 3249
rect 14323 3235 14362 3249
rect 14396 3235 14435 3249
rect 14469 3235 14508 3249
rect 14542 3235 14581 3249
rect 14615 3235 14654 3249
rect 14688 3235 14727 3249
rect 14761 3235 14800 3249
rect 14834 3235 14873 3249
rect 14907 3235 14946 3249
rect 14980 3235 15019 3249
rect 15053 3235 15092 3249
rect 15126 3235 15165 3249
rect 15199 3235 15238 3249
rect 15272 3235 15311 3249
rect 15345 3235 15384 3249
rect 15418 3235 15457 3249
rect 15491 3235 15530 3249
rect 15564 3235 15603 3249
rect 15637 3235 15676 3249
rect 15710 3235 15749 3249
rect 15783 3235 15822 3249
rect 15856 3235 15895 3249
rect 15929 3235 15968 3249
rect 16002 3235 16041 3249
rect 16075 3235 16114 3249
rect 16148 3235 16187 3249
rect 16221 3235 16260 3249
rect 16294 3235 16333 3249
rect 16367 3235 16406 3249
rect 16872 3235 17215 3270
rect 4615 3201 4639 3235
rect 4673 3201 4708 3235
rect 4742 3201 4777 3235
rect 4811 3201 4846 3235
rect 4880 3201 4915 3235
rect 4949 3201 4984 3235
rect 5018 3201 5053 3235
rect 4615 3167 5053 3201
rect 4615 3133 4639 3167
rect 4673 3133 4708 3167
rect 4742 3133 4777 3167
rect 4811 3133 4846 3167
rect 4880 3133 4915 3167
rect 4949 3133 4984 3167
rect 5018 3133 5053 3167
rect 4615 3099 5053 3133
rect 4615 3065 4639 3099
rect 4673 3065 4708 3099
rect 4742 3065 4777 3099
rect 4811 3065 4846 3099
rect 4880 3065 4915 3099
rect 4949 3065 4984 3099
rect 5018 3065 5053 3099
rect 4615 3031 5053 3065
rect 4615 2997 4639 3031
rect 4673 2997 4708 3031
rect 4742 2997 4777 3031
rect 4811 2997 4846 3031
rect 4880 2997 4915 3031
rect 4949 2997 4984 3031
rect 5018 2997 5053 3031
rect 4615 2963 5053 2997
rect 4615 2929 4639 2963
rect 4673 2929 4708 2963
rect 4742 2929 4777 2963
rect 4811 2929 4846 2963
rect 4880 2929 4915 2963
rect 4949 2929 4984 2963
rect 5018 2929 5053 2963
rect 4615 2895 5053 2929
rect 4615 2861 4639 2895
rect 4673 2861 4708 2895
rect 4742 2861 4777 2895
rect 4811 2861 4846 2895
rect 4880 2861 4915 2895
rect 4949 2861 4984 2895
rect 5018 2861 5053 2895
rect 4615 2827 5053 2861
rect 4615 2793 4639 2827
rect 4673 2793 4708 2827
rect 4742 2793 4777 2827
rect 4811 2793 4846 2827
rect 4880 2793 4915 2827
rect 4949 2793 4984 2827
rect 5018 2793 5053 2827
rect 4615 2759 5053 2793
rect 4615 2725 4639 2759
rect 4673 2725 4708 2759
rect 4742 2725 4777 2759
rect 4811 2725 4846 2759
rect 4880 2725 4915 2759
rect 4949 2725 4984 2759
rect 5018 2725 5053 2759
rect 4615 2715 5053 2725
rect 4615 2691 4734 2715
rect 4768 2691 4807 2715
rect 4841 2691 4880 2715
rect 4615 2657 4639 2691
rect 4673 2657 4708 2691
rect 4768 2681 4777 2691
rect 4841 2681 4846 2691
rect 4742 2657 4777 2681
rect 4811 2657 4846 2681
rect 4914 2691 4953 2715
rect 4987 2691 5026 2715
rect 4914 2681 4915 2691
rect 4880 2657 4915 2681
rect 4949 2681 4953 2691
rect 5018 2681 5026 2691
rect 4949 2657 4984 2681
rect 5018 2657 5053 2681
rect 4615 2639 5053 2657
rect 4615 2623 4734 2639
rect 4768 2623 4807 2639
rect 4841 2623 4880 2639
rect 4615 2589 4639 2623
rect 4673 2589 4708 2623
rect 4768 2605 4777 2623
rect 4841 2605 4846 2623
rect 4742 2589 4777 2605
rect 4811 2589 4846 2605
rect 4914 2623 4953 2639
rect 4987 2623 5026 2639
rect 4914 2605 4915 2623
rect 4880 2589 4915 2605
rect 4949 2605 4953 2623
rect 5018 2605 5026 2623
rect 4949 2589 4984 2605
rect 5018 2589 5053 2605
rect 4615 2563 5053 2589
rect 4615 2555 4734 2563
rect 4768 2555 4807 2563
rect 4841 2555 4880 2563
rect 4615 2521 4639 2555
rect 4673 2521 4708 2555
rect 4768 2529 4777 2555
rect 4841 2529 4846 2555
rect 4742 2521 4777 2529
rect 4811 2521 4846 2529
rect 4914 2555 4953 2563
rect 4987 2555 5026 2563
rect 4914 2529 4915 2555
rect 4880 2521 4915 2529
rect 4949 2529 4953 2555
rect 5018 2529 5026 2555
rect 4949 2521 4984 2529
rect 5018 2521 5053 2529
rect 4615 2487 5053 2521
rect 4615 2453 4639 2487
rect 4673 2453 4708 2487
rect 4768 2453 4777 2487
rect 4841 2453 4846 2487
rect 4914 2453 4915 2487
rect 4949 2453 4953 2487
rect 5018 2453 5026 2487
rect 4615 2419 5053 2453
rect 4615 2385 4639 2419
rect 4673 2385 4708 2419
rect 4742 2411 4777 2419
rect 4811 2411 4846 2419
rect 4768 2385 4777 2411
rect 4841 2385 4846 2411
rect 4880 2411 4915 2419
rect 4615 2377 4734 2385
rect 4768 2377 4807 2385
rect 4841 2377 4880 2385
rect 4914 2385 4915 2411
rect 4949 2411 4984 2419
rect 5018 2411 5053 2419
rect 4949 2385 4953 2411
rect 5018 2385 5026 2411
rect 4914 2377 4953 2385
rect 4987 2377 5026 2385
rect 4615 2351 5053 2377
rect 4615 2317 4639 2351
rect 4673 2317 4708 2351
rect 4742 2335 4777 2351
rect 4811 2335 4846 2351
rect 4768 2317 4777 2335
rect 4841 2317 4846 2335
rect 4880 2335 4915 2351
rect 4615 2301 4734 2317
rect 4768 2301 4807 2317
rect 4841 2301 4880 2317
rect 4914 2317 4915 2335
rect 4949 2335 4984 2351
rect 5018 2335 5053 2351
rect 4949 2317 4953 2335
rect 5018 2317 5026 2335
rect 4914 2301 4953 2317
rect 4987 2301 5026 2317
rect 4615 2283 5053 2301
rect 4615 2249 4639 2283
rect 4673 2249 4708 2283
rect 4742 2259 4777 2283
rect 4811 2259 4846 2283
rect 4768 2249 4777 2259
rect 4841 2249 4846 2259
rect 4880 2259 4915 2283
rect 4615 2225 4734 2249
rect 4768 2225 4807 2249
rect 4841 2225 4880 2249
rect 4914 2249 4915 2259
rect 4949 2259 4984 2283
rect 5018 2259 5053 2283
rect 4949 2249 4953 2259
rect 5018 2249 5026 2259
rect 4914 2225 4953 2249
rect 4987 2225 5026 2249
rect 4615 2215 5053 2225
rect 4615 2181 4639 2215
rect 4673 2181 4708 2215
rect 4742 2183 4777 2215
rect 4811 2183 4846 2215
rect 4768 2181 4777 2183
rect 4841 2181 4846 2183
rect 4880 2183 4915 2215
rect 4615 2149 4734 2181
rect 4768 2149 4807 2181
rect 4841 2149 4880 2181
rect 4914 2181 4915 2183
rect 4949 2183 4984 2215
rect 5018 2183 5053 2215
rect 4949 2181 4953 2183
rect 5018 2181 5026 2183
rect 17191 2181 17215 3235
rect 4914 2149 4953 2181
rect 4987 2149 5026 2181
rect 5060 2149 5099 2181
rect 5133 2149 5172 2181
rect 5206 2149 5245 2181
rect 5279 2149 5318 2181
rect 5352 2149 5391 2181
rect 5425 2149 5464 2181
rect 5498 2149 5537 2181
rect 5571 2149 5610 2181
rect 5644 2149 5683 2181
rect 5717 2149 5756 2181
rect 5790 2149 5829 2181
rect 5863 2149 5902 2181
rect 5936 2149 5975 2181
rect 6009 2149 6048 2181
rect 6082 2149 6121 2181
rect 6155 2149 6194 2181
rect 6228 2149 6267 2181
rect 6301 2149 6340 2181
rect 6374 2149 6413 2181
rect 6447 2149 6486 2181
rect 6520 2149 6559 2181
rect 6593 2149 6632 2181
rect 6666 2149 6705 2181
rect 6739 2149 6778 2181
rect 6812 2149 6851 2181
rect 6885 2149 6924 2181
rect 6958 2149 6997 2181
rect 7031 2149 7070 2181
rect 7104 2149 7143 2181
rect 7177 2149 7216 2181
rect 7250 2149 7289 2181
rect 7323 2149 7362 2181
rect 7396 2149 7435 2181
rect 7469 2149 7508 2181
rect 7542 2149 7581 2181
rect 7615 2149 7654 2181
rect 7688 2149 7727 2181
rect 7761 2149 7800 2181
rect 7834 2149 7873 2181
rect 7907 2149 7946 2181
rect 7980 2149 8019 2181
rect 8053 2149 8092 2181
rect 8126 2149 8165 2181
rect 8199 2149 8238 2181
rect 8272 2149 8311 2181
rect 8345 2149 8384 2181
rect 8418 2149 8457 2181
rect 8491 2149 8530 2181
rect 8564 2149 8603 2181
rect 8637 2149 8676 2181
rect 8710 2149 8749 2181
rect 8783 2149 8822 2181
rect 8856 2149 8895 2181
rect 8929 2149 8968 2181
rect 9002 2149 9041 2181
rect 9075 2149 9114 2181
rect 9148 2149 9187 2181
rect 9221 2149 9260 2181
rect 9294 2149 9333 2181
rect 9367 2149 9406 2181
rect 9440 2149 9479 2181
rect 9513 2149 9552 2181
rect 9586 2149 9625 2181
rect 9659 2149 9698 2181
rect 9732 2149 9771 2181
rect 9805 2149 9844 2181
rect 9878 2149 9917 2181
rect 9951 2149 9989 2181
rect 10023 2149 10061 2181
rect 10095 2149 10133 2181
rect 10167 2149 10205 2181
rect 10239 2149 10277 2181
rect 10311 2149 10349 2181
rect 10383 2149 10421 2181
rect 10455 2149 10493 2181
rect 10527 2149 10565 2181
rect 10599 2149 10637 2181
rect 10671 2149 10709 2181
rect 10743 2149 10781 2181
rect 10815 2149 10853 2181
rect 10887 2149 10925 2181
rect 10959 2159 11967 2181
rect 12001 2159 12040 2181
rect 12074 2159 12113 2181
rect 12147 2159 12186 2181
rect 12220 2159 12259 2181
rect 12293 2159 12332 2181
rect 12366 2159 12405 2181
rect 12439 2159 12478 2181
rect 12512 2159 12551 2181
rect 12585 2159 12624 2181
rect 12658 2159 12697 2181
rect 12731 2159 12770 2181
rect 12804 2159 12843 2181
rect 12877 2159 12916 2181
rect 12950 2159 12989 2181
rect 13023 2159 13062 2181
rect 13096 2159 13135 2181
rect 13169 2159 13208 2181
rect 13242 2159 13281 2181
rect 13315 2159 13354 2181
rect 13388 2159 13427 2181
rect 13461 2159 13500 2181
rect 13534 2159 13573 2181
rect 13607 2159 13646 2181
rect 13680 2159 13719 2181
rect 13753 2159 13792 2181
rect 13826 2159 13865 2181
rect 13899 2159 13938 2181
rect 13972 2159 14011 2181
rect 14045 2159 14084 2181
rect 14118 2159 14157 2181
rect 16927 2159 17215 2181
rect 10959 2149 15944 2159
rect 4615 2148 15944 2149
rect 4615 2147 5729 2148
rect 4649 2113 4686 2147
rect 4720 2113 4757 2147
rect 4791 2113 4828 2147
rect 4862 2113 4899 2147
rect 4933 2113 4970 2147
rect 5004 2113 5041 2147
rect 5075 2113 5112 2147
rect 5146 2113 5183 2147
rect 5217 2113 5254 2147
rect 5288 2113 5325 2147
rect 5359 2113 5396 2147
rect 5430 2113 5467 2147
rect 5501 2113 5537 2147
rect 5571 2113 5607 2147
rect 5641 2113 5677 2147
rect 5711 2113 5729 2147
rect 4615 2071 5729 2113
rect 4649 2037 4686 2071
rect 4720 2037 4757 2071
rect 4791 2037 4828 2071
rect 4862 2037 4899 2071
rect 4933 2037 4970 2071
rect 5004 2037 5041 2071
rect 5075 2037 5112 2071
rect 5146 2037 5183 2071
rect 5217 2037 5254 2071
rect 5288 2037 5325 2071
rect 5359 2037 5396 2071
rect 5430 2037 5467 2071
rect 5501 2037 5537 2071
rect 5571 2037 5607 2071
rect 5641 2037 5677 2071
rect 5711 2037 5729 2071
rect 4615 1995 5729 2037
rect 4649 1961 4686 1995
rect 4720 1961 4757 1995
rect 4791 1961 4828 1995
rect 4862 1961 4899 1995
rect 4933 1961 4970 1995
rect 5004 1961 5041 1995
rect 5075 1961 5112 1995
rect 5146 1961 5183 1995
rect 5217 1961 5254 1995
rect 5288 1961 5325 1995
rect 5359 1961 5396 1995
rect 5430 1961 5467 1995
rect 5501 1961 5537 1995
rect 5571 1961 5607 1995
rect 5641 1961 5677 1995
rect 5711 1961 5729 1995
rect 4615 1919 5729 1961
rect 4649 1885 4686 1919
rect 4720 1885 4757 1919
rect 4791 1885 4828 1919
rect 4862 1885 4899 1919
rect 4933 1885 4970 1919
rect 5004 1885 5041 1919
rect 5075 1885 5112 1919
rect 5146 1885 5183 1919
rect 5217 1885 5254 1919
rect 5288 1885 5325 1919
rect 5359 1885 5396 1919
rect 5430 1885 5467 1919
rect 5501 1885 5537 1919
rect 5571 1885 5607 1919
rect 5641 1885 5677 1919
rect 5711 1885 5729 1919
rect 6524 1902 15944 2148
rect 4615 1870 5729 1885
rect -2859 1859 5729 1870
rect 15540 1859 15944 1902
rect -2859 1858 15944 1859
rect -2859 1846 4616 1858
rect 4650 1846 4688 1858
rect 4722 1846 4760 1858
rect 4794 1846 4832 1858
rect 4866 1846 4904 1858
rect 4938 1846 4976 1858
rect 5010 1846 5048 1858
rect 5082 1846 5120 1858
rect 5154 1846 5192 1858
rect 5226 1846 5264 1858
rect 5298 1846 5336 1858
rect 5370 1846 5408 1858
rect 5442 1846 5480 1858
rect 5514 1846 5552 1858
rect 5586 1846 5624 1858
rect 5658 1846 5696 1858
rect -2825 1841 -2790 1846
rect -2756 1841 -2721 1846
rect -2798 1812 -2790 1841
rect -2725 1812 -2721 1841
rect -2687 1841 -2652 1846
rect -2687 1812 -2686 1841
rect -2859 1807 -2832 1812
rect -2798 1807 -2759 1812
rect -2725 1807 -2686 1812
rect -2618 1841 -2583 1846
rect -2549 1841 -2514 1846
rect -2480 1841 -2445 1846
rect -2411 1841 -2376 1846
rect -2342 1841 -2307 1846
rect -2273 1841 -2238 1846
rect -2204 1841 -2169 1846
rect -2135 1841 -2100 1846
rect -2618 1812 -2613 1841
rect -2549 1812 -2540 1841
rect -2480 1812 -2467 1841
rect -2411 1812 -2394 1841
rect -2342 1812 -2321 1841
rect -2273 1812 -2248 1841
rect -2204 1812 -2175 1841
rect -2135 1812 -2102 1841
rect -2066 1812 -2031 1846
rect -1997 1841 -1962 1846
rect -1928 1841 -1893 1846
rect -1859 1841 -1824 1846
rect -1790 1841 -1755 1846
rect -1721 1841 -1686 1846
rect -1652 1841 -1617 1846
rect -1583 1841 -1548 1846
rect -1514 1841 -1479 1846
rect -1445 1841 -1410 1846
rect -1376 1841 -1341 1846
rect -1307 1841 -1272 1846
rect -1238 1841 -1203 1846
rect -1169 1841 -1134 1846
rect -1100 1841 -1065 1846
rect -1031 1841 -996 1846
rect -962 1841 -927 1846
rect -893 1841 -858 1846
rect -824 1841 -789 1846
rect -755 1841 -720 1846
rect -686 1841 -651 1846
rect -617 1841 -582 1846
rect -548 1841 -513 1846
rect -479 1841 -444 1846
rect -410 1841 -375 1846
rect -1 1841 33 1846
rect -1995 1812 -1962 1841
rect -1922 1812 -1893 1841
rect -1849 1812 -1824 1841
rect -1776 1812 -1755 1841
rect -2652 1807 -2613 1812
rect -2579 1807 -2540 1812
rect -2506 1807 -2467 1812
rect -2433 1807 -2394 1812
rect -2360 1807 -2321 1812
rect -2287 1807 -2248 1812
rect -2214 1807 -2175 1812
rect -2141 1807 -2102 1812
rect -2068 1807 -2029 1812
rect -1995 1807 -1956 1812
rect -1922 1807 -1883 1812
rect -1849 1807 -1810 1812
rect -1776 1807 -1737 1812
rect -2859 1778 -1737 1807
rect -2825 1769 -2790 1778
rect -2756 1769 -2721 1778
rect -2798 1744 -2790 1769
rect -2725 1744 -2721 1769
rect -2687 1769 -2652 1778
rect -2687 1744 -2686 1769
rect -2859 1735 -2832 1744
rect -2798 1735 -2759 1744
rect -2725 1735 -2686 1744
rect -2618 1769 -2583 1778
rect -2549 1769 -2514 1778
rect -2480 1769 -2445 1778
rect -2411 1769 -2376 1778
rect -2342 1769 -2307 1778
rect -2273 1769 -2238 1778
rect -2204 1769 -2169 1778
rect -2135 1769 -2100 1778
rect -2618 1744 -2613 1769
rect -2549 1744 -2540 1769
rect -2480 1744 -2467 1769
rect -2411 1744 -2394 1769
rect -2342 1744 -2321 1769
rect -2273 1744 -2248 1769
rect -2204 1744 -2175 1769
rect -2135 1744 -2102 1769
rect -2066 1744 -2031 1778
rect -1997 1769 -1962 1778
rect -1928 1769 -1893 1778
rect -1859 1769 -1824 1778
rect -1790 1769 -1755 1778
rect -1995 1744 -1962 1769
rect -1922 1744 -1893 1769
rect -1849 1744 -1824 1769
rect -1776 1744 -1755 1769
rect -2652 1735 -2613 1744
rect -2579 1735 -2540 1744
rect -2506 1735 -2467 1744
rect -2433 1735 -2394 1744
rect -2360 1735 -2321 1744
rect -2287 1735 -2248 1744
rect -2214 1735 -2175 1744
rect -2141 1735 -2102 1744
rect -2068 1735 -2029 1744
rect -1995 1735 -1956 1744
rect -1922 1735 -1883 1744
rect -1849 1735 -1810 1744
rect -1776 1735 -1737 1744
rect -2859 1710 -1737 1735
rect -2825 1697 -2790 1710
rect -2756 1697 -2721 1710
rect -2798 1676 -2790 1697
rect -2725 1676 -2721 1697
rect -2687 1697 -2652 1710
rect -2687 1676 -2686 1697
rect -2859 1663 -2832 1676
rect -2798 1663 -2759 1676
rect -2725 1663 -2686 1676
rect -2618 1697 -2583 1710
rect -2549 1697 -2514 1710
rect -2480 1697 -2445 1710
rect -2411 1697 -2376 1710
rect -2342 1697 -2307 1710
rect -2273 1697 -2238 1710
rect -2204 1697 -2169 1710
rect -2135 1697 -2100 1710
rect -2618 1676 -2613 1697
rect -2549 1676 -2540 1697
rect -2480 1676 -2467 1697
rect -2411 1676 -2394 1697
rect -2342 1676 -2321 1697
rect -2273 1676 -2248 1697
rect -2204 1676 -2175 1697
rect -2135 1676 -2102 1697
rect -2066 1676 -2031 1710
rect -1997 1697 -1962 1710
rect -1928 1697 -1893 1710
rect -1859 1697 -1824 1710
rect -1790 1697 -1755 1710
rect -1995 1676 -1962 1697
rect -1922 1676 -1893 1697
rect -1849 1676 -1824 1697
rect -1776 1676 -1755 1697
rect -2652 1663 -2613 1676
rect -2579 1663 -2540 1676
rect -2506 1663 -2467 1676
rect -2433 1663 -2394 1676
rect -2360 1663 -2321 1676
rect -2287 1663 -2248 1676
rect -2214 1663 -2175 1676
rect -2141 1663 -2102 1676
rect -2068 1663 -2029 1676
rect -1995 1663 -1956 1676
rect -1922 1663 -1883 1676
rect -1849 1663 -1810 1676
rect -1776 1663 -1737 1676
rect -2859 1642 -1737 1663
rect -2825 1625 -2790 1642
rect -2756 1625 -2721 1642
rect -2798 1608 -2790 1625
rect -2725 1608 -2721 1625
rect -2687 1625 -2652 1642
rect -2687 1608 -2686 1625
rect -2859 1591 -2832 1608
rect -2798 1591 -2759 1608
rect -2725 1591 -2686 1608
rect -2618 1625 -2583 1642
rect -2549 1625 -2514 1642
rect -2480 1625 -2445 1642
rect -2411 1625 -2376 1642
rect -2342 1625 -2307 1642
rect -2273 1625 -2238 1642
rect -2204 1625 -2169 1642
rect -2135 1625 -2100 1642
rect -2618 1608 -2613 1625
rect -2549 1608 -2540 1625
rect -2480 1608 -2467 1625
rect -2411 1608 -2394 1625
rect -2342 1608 -2321 1625
rect -2273 1608 -2248 1625
rect -2204 1608 -2175 1625
rect -2135 1608 -2102 1625
rect -2066 1608 -2031 1642
rect -1997 1625 -1962 1642
rect -1928 1625 -1893 1642
rect -1859 1625 -1824 1642
rect -1790 1625 -1755 1642
rect -1995 1608 -1962 1625
rect -1922 1608 -1893 1625
rect -1849 1608 -1824 1625
rect -1776 1608 -1755 1625
rect -2652 1591 -2613 1608
rect -2579 1591 -2540 1608
rect -2506 1591 -2467 1608
rect -2433 1591 -2394 1608
rect -2360 1591 -2321 1608
rect -2287 1591 -2248 1608
rect -2214 1591 -2175 1608
rect -2141 1591 -2102 1608
rect -2068 1591 -2029 1608
rect -1995 1591 -1956 1608
rect -1922 1591 -1883 1608
rect -1849 1591 -1810 1608
rect -1776 1591 -1737 1608
rect -2859 1574 -1737 1591
rect -2825 1553 -2790 1574
rect -2756 1553 -2721 1574
rect -2798 1540 -2790 1553
rect -2725 1540 -2721 1553
rect -2687 1553 -2652 1574
rect -2687 1540 -2686 1553
rect -2859 1519 -2832 1540
rect -2798 1519 -2759 1540
rect -2725 1519 -2686 1540
rect -2618 1553 -2583 1574
rect -2549 1553 -2514 1574
rect -2480 1553 -2445 1574
rect -2411 1553 -2376 1574
rect -2342 1553 -2307 1574
rect -2273 1553 -2238 1574
rect -2204 1553 -2169 1574
rect -2135 1553 -2100 1574
rect -2618 1540 -2613 1553
rect -2549 1540 -2540 1553
rect -2480 1540 -2467 1553
rect -2411 1540 -2394 1553
rect -2342 1540 -2321 1553
rect -2273 1540 -2248 1553
rect -2204 1540 -2175 1553
rect -2135 1540 -2102 1553
rect -2066 1540 -2031 1574
rect -1997 1553 -1962 1574
rect -1928 1553 -1893 1574
rect -1859 1553 -1824 1574
rect -1790 1553 -1755 1574
rect -1995 1540 -1962 1553
rect -1922 1540 -1893 1553
rect -1849 1540 -1824 1553
rect -1776 1540 -1755 1553
rect -2652 1519 -2613 1540
rect -2579 1519 -2540 1540
rect -2506 1519 -2467 1540
rect -2433 1519 -2394 1540
rect -2360 1519 -2321 1540
rect -2287 1519 -2248 1540
rect -2214 1519 -2175 1540
rect -2141 1519 -2102 1540
rect -2068 1519 -2029 1540
rect -1995 1519 -1956 1540
rect -1922 1519 -1883 1540
rect -1849 1519 -1810 1540
rect -1776 1519 -1737 1540
rect -2859 1506 -1737 1519
rect -2825 1481 -2790 1506
rect -2756 1481 -2721 1506
rect -2798 1472 -2790 1481
rect -2725 1472 -2721 1481
rect -2687 1481 -2652 1506
rect -2687 1472 -2686 1481
rect -2859 1447 -2832 1472
rect -2798 1447 -2759 1472
rect -2725 1447 -2686 1472
rect -2618 1481 -2583 1506
rect -2549 1481 -2514 1506
rect -2480 1481 -2445 1506
rect -2411 1481 -2376 1506
rect -2342 1481 -2307 1506
rect -2273 1481 -2238 1506
rect -2204 1481 -2169 1506
rect -2135 1481 -2100 1506
rect -2618 1472 -2613 1481
rect -2549 1472 -2540 1481
rect -2480 1472 -2467 1481
rect -2411 1472 -2394 1481
rect -2342 1472 -2321 1481
rect -2273 1472 -2248 1481
rect -2204 1472 -2175 1481
rect -2135 1472 -2102 1481
rect -2066 1472 -2031 1506
rect -1997 1481 -1962 1506
rect -1928 1481 -1893 1506
rect -1859 1481 -1824 1506
rect -1790 1481 -1755 1506
rect -1995 1472 -1962 1481
rect -1922 1472 -1893 1481
rect -1849 1472 -1824 1481
rect -1776 1472 -1755 1481
rect -2652 1447 -2613 1472
rect -2579 1447 -2540 1472
rect -2506 1447 -2467 1472
rect -2433 1447 -2394 1472
rect -2360 1447 -2321 1472
rect -2287 1447 -2248 1472
rect -2214 1447 -2175 1472
rect -2141 1447 -2102 1472
rect -2068 1447 -2029 1472
rect -1995 1447 -1956 1472
rect -1922 1447 -1883 1472
rect -1849 1447 -1810 1472
rect -1776 1447 -1737 1472
rect -2859 1438 -1737 1447
rect -2825 1409 -2790 1438
rect -2756 1409 -2721 1438
rect -2798 1404 -2790 1409
rect -2725 1404 -2721 1409
rect -2687 1409 -2652 1438
rect -2687 1404 -2686 1409
rect -2859 1375 -2832 1404
rect -2798 1375 -2759 1404
rect -2725 1375 -2686 1404
rect -2618 1409 -2583 1438
rect -2549 1409 -2514 1438
rect -2480 1409 -2445 1438
rect -2411 1409 -2376 1438
rect -2342 1409 -2307 1438
rect -2273 1409 -2238 1438
rect -2204 1409 -2169 1438
rect -2135 1409 -2100 1438
rect -2618 1404 -2613 1409
rect -2549 1404 -2540 1409
rect -2480 1404 -2467 1409
rect -2411 1404 -2394 1409
rect -2342 1404 -2321 1409
rect -2273 1404 -2248 1409
rect -2204 1404 -2175 1409
rect -2135 1404 -2102 1409
rect -2066 1404 -2031 1438
rect -1997 1409 -1962 1438
rect -1928 1409 -1893 1438
rect -1859 1409 -1824 1438
rect -1790 1409 -1755 1438
rect -1995 1404 -1962 1409
rect -1922 1404 -1893 1409
rect -1849 1404 -1824 1409
rect -1776 1404 -1755 1409
rect -2652 1375 -2613 1404
rect -2579 1375 -2540 1404
rect -2506 1375 -2467 1404
rect -2433 1375 -2394 1404
rect -2360 1375 -2321 1404
rect -2287 1375 -2248 1404
rect -2214 1375 -2175 1404
rect -2141 1375 -2102 1404
rect -2068 1375 -2029 1404
rect -1995 1375 -1956 1404
rect -1922 1375 -1883 1404
rect -1849 1375 -1810 1404
rect -1776 1375 -1737 1404
rect -2859 1370 -1737 1375
rect -2825 1337 -2790 1370
rect -2756 1337 -2721 1370
rect -2798 1336 -2790 1337
rect -2725 1336 -2721 1337
rect -2687 1337 -2652 1370
rect -2687 1336 -2686 1337
rect -2859 1303 -2832 1336
rect -2798 1303 -2759 1336
rect -2725 1303 -2686 1336
rect -2618 1337 -2583 1370
rect -2549 1337 -2514 1370
rect -2480 1337 -2445 1370
rect -2411 1337 -2376 1370
rect -2342 1337 -2307 1370
rect -2273 1337 -2238 1370
rect -2204 1337 -2169 1370
rect -2135 1337 -2100 1370
rect -2618 1336 -2613 1337
rect -2549 1336 -2540 1337
rect -2480 1336 -2467 1337
rect -2411 1336 -2394 1337
rect -2342 1336 -2321 1337
rect -2273 1336 -2248 1337
rect -2204 1336 -2175 1337
rect -2135 1336 -2102 1337
rect -2066 1336 -2031 1370
rect -1997 1337 -1962 1370
rect -1928 1337 -1893 1370
rect -1859 1337 -1824 1370
rect -1790 1337 -1755 1370
rect -1995 1336 -1962 1337
rect -1922 1336 -1893 1337
rect -1849 1336 -1824 1337
rect -1776 1336 -1755 1337
rect -2652 1303 -2613 1336
rect -2579 1303 -2540 1336
rect -2506 1303 -2467 1336
rect -2433 1303 -2394 1336
rect -2360 1303 -2321 1336
rect -2287 1303 -2248 1336
rect -2214 1303 -2175 1336
rect -2141 1303 -2102 1336
rect -2068 1303 -2029 1336
rect -1995 1303 -1956 1336
rect -1922 1303 -1883 1336
rect -1849 1303 -1810 1336
rect -1776 1303 -1737 1336
rect -2859 1302 -1737 1303
rect -2825 1268 -2790 1302
rect -2756 1268 -2721 1302
rect -2687 1268 -2652 1302
rect -2618 1268 -2583 1302
rect -2549 1268 -2514 1302
rect -2480 1268 -2445 1302
rect -2411 1268 -2376 1302
rect -2342 1268 -2307 1302
rect -2273 1268 -2238 1302
rect -2204 1268 -2169 1302
rect -2135 1268 -2100 1302
rect -2066 1268 -2031 1302
rect -1997 1268 -1962 1302
rect -1928 1268 -1893 1302
rect -1859 1268 -1824 1302
rect -1790 1268 -1755 1302
rect -2859 1265 -1737 1268
rect -2859 1234 -2832 1265
rect -2798 1234 -2759 1265
rect -2725 1234 -2686 1265
rect -2798 1231 -2790 1234
rect -2725 1231 -2721 1234
rect -2825 1200 -2790 1231
rect -2756 1200 -2721 1231
rect -2687 1231 -2686 1234
rect -2652 1234 -2613 1265
rect -2579 1234 -2540 1265
rect -2506 1234 -2467 1265
rect -2433 1234 -2394 1265
rect -2360 1234 -2321 1265
rect -2287 1234 -2248 1265
rect -2214 1234 -2175 1265
rect -2141 1234 -2102 1265
rect -2068 1234 -2029 1265
rect -1995 1234 -1956 1265
rect -1922 1234 -1883 1265
rect -1849 1234 -1810 1265
rect -1776 1234 -1737 1265
rect -2687 1200 -2652 1231
rect -2618 1231 -2613 1234
rect -2549 1231 -2540 1234
rect -2480 1231 -2467 1234
rect -2411 1231 -2394 1234
rect -2342 1231 -2321 1234
rect -2273 1231 -2248 1234
rect -2204 1231 -2175 1234
rect -2135 1231 -2102 1234
rect -2618 1200 -2583 1231
rect -2549 1200 -2514 1231
rect -2480 1200 -2445 1231
rect -2411 1200 -2376 1231
rect -2342 1200 -2307 1231
rect -2273 1200 -2238 1231
rect -2204 1200 -2169 1231
rect -2135 1200 -2100 1231
rect -2066 1200 -2031 1234
rect -1995 1231 -1962 1234
rect -1922 1231 -1893 1234
rect -1849 1231 -1824 1234
rect -1776 1231 -1755 1234
rect 5730 1824 5768 1858
rect 5802 1824 5840 1858
rect 5874 1824 5912 1858
rect 5946 1824 5984 1858
rect 6018 1824 6056 1858
rect 6090 1824 6128 1858
rect 6162 1824 6200 1858
rect 6234 1824 6272 1858
rect 6306 1824 6344 1858
rect 6378 1824 6416 1858
rect 6450 1824 6488 1858
rect 6522 1824 6560 1858
rect 6594 1824 6632 1858
rect 6666 1824 6704 1858
rect 6738 1824 6776 1858
rect 6810 1824 6848 1858
rect 6882 1824 6920 1858
rect 6954 1824 6992 1858
rect 7026 1824 7064 1858
rect 7098 1824 7136 1858
rect 7170 1824 7208 1858
rect 7242 1824 7280 1858
rect 7314 1824 7352 1858
rect 7386 1824 7424 1858
rect 7458 1824 7496 1858
rect 7530 1824 7568 1858
rect 7602 1824 7640 1858
rect 7674 1824 7712 1858
rect 7746 1824 7784 1858
rect 7818 1824 7856 1858
rect 7890 1824 7928 1858
rect 7962 1824 8000 1858
rect 8034 1824 8072 1858
rect 8106 1824 8144 1858
rect 8178 1824 8216 1858
rect 8250 1824 8288 1858
rect 8322 1824 8360 1858
rect 8394 1824 8432 1858
rect 8466 1824 8504 1858
rect 8538 1824 8576 1858
rect 8610 1824 8648 1858
rect 8682 1824 8720 1858
rect 8754 1824 8792 1858
rect 8826 1824 8864 1858
rect 8898 1824 8936 1858
rect 8970 1824 9008 1858
rect 9042 1824 9080 1858
rect 9114 1824 9152 1858
rect 9186 1824 9224 1858
rect 9258 1824 9296 1858
rect 9330 1824 9368 1858
rect 9402 1824 9440 1858
rect 9474 1824 9512 1858
rect 9546 1824 9584 1858
rect 9618 1824 9656 1858
rect 9690 1824 9728 1858
rect 9762 1824 9800 1858
rect 9834 1824 9872 1858
rect 9906 1824 9944 1858
rect 9978 1824 10016 1858
rect 10050 1824 10088 1858
rect 10122 1824 10160 1858
rect 10194 1824 10232 1858
rect 10266 1824 10304 1858
rect 10338 1824 10376 1858
rect 10410 1824 10448 1858
rect 10482 1824 10520 1858
rect 10554 1824 10592 1858
rect 10626 1824 10664 1858
rect 10698 1824 10736 1858
rect 10770 1824 10808 1858
rect 10842 1824 10880 1858
rect 10914 1824 10952 1858
rect 10986 1824 11024 1858
rect 11058 1824 11096 1858
rect 11130 1824 11168 1858
rect 11202 1824 11240 1858
rect 11274 1824 11312 1858
rect 11346 1824 11384 1858
rect 11418 1824 11456 1858
rect 11490 1824 11528 1858
rect 11562 1824 11600 1858
rect 11634 1824 11672 1858
rect 11706 1824 11744 1858
rect 11778 1824 11816 1858
rect 11850 1824 11888 1858
rect 11922 1824 11960 1858
rect 11994 1824 12032 1858
rect 12066 1824 12104 1858
rect 12138 1824 12176 1858
rect 12210 1824 12248 1858
rect 12282 1824 12320 1858
rect 12354 1824 12392 1858
rect 12426 1824 12464 1858
rect 12498 1824 12536 1858
rect 12570 1824 12608 1858
rect 12642 1824 12680 1858
rect 12714 1824 12752 1858
rect 12786 1824 12824 1858
rect 12858 1824 12896 1858
rect 12930 1824 12968 1858
rect 13002 1824 13040 1858
rect 13074 1824 13112 1858
rect 13146 1824 13184 1858
rect 13218 1824 13256 1858
rect 13290 1824 13328 1858
rect 13362 1824 13400 1858
rect 13434 1824 13472 1858
rect 13506 1824 13544 1858
rect 13578 1824 13616 1858
rect 13650 1824 13688 1858
rect 13722 1824 13760 1858
rect 13794 1824 13832 1858
rect 13866 1824 13904 1858
rect 13938 1824 13976 1858
rect 14010 1824 14048 1858
rect 14082 1824 14120 1858
rect 14154 1824 14192 1858
rect 14226 1824 14264 1858
rect 14298 1824 14336 1858
rect 14370 1824 14408 1858
rect 14442 1824 14480 1858
rect 14514 1824 14552 1858
rect 14586 1824 14624 1858
rect 14658 1824 14696 1858
rect 14730 1824 14768 1858
rect 14802 1824 14840 1858
rect 14874 1824 14912 1858
rect 14946 1824 14984 1858
rect 15018 1824 15056 1858
rect 15090 1824 15128 1858
rect 15162 1824 15200 1858
rect 15234 1824 15272 1858
rect 15306 1824 15344 1858
rect 15378 1824 15416 1858
rect 15450 1824 15488 1858
rect 15522 1824 15561 1858
rect 15595 1824 15634 1858
rect 15668 1824 15707 1858
rect 15741 1824 15780 1858
rect 15814 1824 15853 1858
rect 15887 1824 15926 1858
rect 5711 1780 15944 1824
rect 5730 1746 5768 1780
rect 5802 1746 5840 1780
rect 5874 1746 5912 1780
rect 5946 1746 5984 1780
rect 6018 1746 6056 1780
rect 6090 1746 6128 1780
rect 6162 1746 6200 1780
rect 6234 1746 6272 1780
rect 6306 1746 6344 1780
rect 6378 1746 6416 1780
rect 6450 1746 6488 1780
rect 6522 1746 6560 1780
rect 6594 1746 6632 1780
rect 6666 1746 6704 1780
rect 6738 1746 6776 1780
rect 6810 1746 6848 1780
rect 6882 1746 6920 1780
rect 6954 1746 6992 1780
rect 7026 1746 7064 1780
rect 7098 1746 7136 1780
rect 7170 1746 7208 1780
rect 7242 1746 7280 1780
rect 7314 1746 7352 1780
rect 7386 1746 7424 1780
rect 7458 1746 7496 1780
rect 7530 1746 7568 1780
rect 7602 1746 7640 1780
rect 7674 1746 7712 1780
rect 7746 1746 7784 1780
rect 7818 1746 7856 1780
rect 7890 1746 7928 1780
rect 7962 1746 8000 1780
rect 8034 1746 8072 1780
rect 8106 1746 8144 1780
rect 8178 1746 8216 1780
rect 8250 1746 8288 1780
rect 8322 1746 8360 1780
rect 8394 1746 8432 1780
rect 8466 1746 8504 1780
rect 8538 1746 8576 1780
rect 8610 1746 8648 1780
rect 8682 1746 8720 1780
rect 8754 1746 8792 1780
rect 8826 1746 8864 1780
rect 8898 1746 8936 1780
rect 8970 1746 9008 1780
rect 9042 1746 9080 1780
rect 9114 1746 9152 1780
rect 9186 1746 9224 1780
rect 9258 1746 9296 1780
rect 9330 1746 9368 1780
rect 9402 1746 9440 1780
rect 9474 1746 9512 1780
rect 9546 1746 9584 1780
rect 9618 1746 9656 1780
rect 9690 1746 9728 1780
rect 9762 1746 9800 1780
rect 9834 1746 9872 1780
rect 9906 1746 9944 1780
rect 9978 1746 10016 1780
rect 10050 1746 10088 1780
rect 10122 1746 10160 1780
rect 10194 1746 10232 1780
rect 10266 1746 10304 1780
rect 10338 1746 10376 1780
rect 10410 1746 10448 1780
rect 10482 1746 10520 1780
rect 10554 1746 10592 1780
rect 10626 1746 10664 1780
rect 10698 1746 10736 1780
rect 10770 1746 10808 1780
rect 10842 1746 10880 1780
rect 10914 1746 10952 1780
rect 10986 1746 11024 1780
rect 11058 1746 11096 1780
rect 11130 1746 11168 1780
rect 11202 1746 11240 1780
rect 11274 1746 11312 1780
rect 11346 1746 11384 1780
rect 11418 1746 11456 1780
rect 11490 1746 11528 1780
rect 11562 1746 11600 1780
rect 11634 1746 11672 1780
rect 11706 1746 11744 1780
rect 11778 1746 11816 1780
rect 11850 1746 11888 1780
rect 11922 1746 11960 1780
rect 11994 1746 12032 1780
rect 12066 1746 12104 1780
rect 12138 1746 12176 1780
rect 12210 1746 12248 1780
rect 12282 1746 12320 1780
rect 12354 1746 12392 1780
rect 12426 1746 12464 1780
rect 12498 1746 12536 1780
rect 12570 1746 12608 1780
rect 12642 1746 12680 1780
rect 12714 1746 12752 1780
rect 12786 1746 12824 1780
rect 12858 1746 12896 1780
rect 12930 1746 12968 1780
rect 13002 1746 13040 1780
rect 13074 1746 13112 1780
rect 13146 1746 13184 1780
rect 13218 1746 13256 1780
rect 13290 1746 13328 1780
rect 13362 1746 13400 1780
rect 13434 1746 13472 1780
rect 13506 1746 13544 1780
rect 13578 1746 13616 1780
rect 13650 1746 13688 1780
rect 13722 1746 13760 1780
rect 13794 1746 13832 1780
rect 13866 1746 13904 1780
rect 13938 1746 13976 1780
rect 14010 1746 14048 1780
rect 14082 1746 14120 1780
rect 14154 1746 14192 1780
rect 14226 1746 14264 1780
rect 14298 1746 14336 1780
rect 14370 1746 14408 1780
rect 14442 1746 14480 1780
rect 14514 1746 14552 1780
rect 14586 1746 14624 1780
rect 14658 1746 14696 1780
rect 14730 1746 14768 1780
rect 14802 1746 14840 1780
rect 14874 1746 14912 1780
rect 14946 1746 14984 1780
rect 15018 1746 15056 1780
rect 15090 1746 15128 1780
rect 15162 1746 15200 1780
rect 15234 1746 15272 1780
rect 15306 1746 15344 1780
rect 15378 1746 15416 1780
rect 15450 1746 15488 1780
rect 15522 1746 15561 1780
rect 15595 1746 15634 1780
rect 15668 1746 15707 1780
rect 15741 1746 15780 1780
rect 15814 1746 15853 1780
rect 15887 1746 15926 1780
rect 5711 1702 15944 1746
rect 5730 1668 5768 1702
rect 5802 1668 5840 1702
rect 5874 1668 5912 1702
rect 5946 1668 5984 1702
rect 6018 1668 6056 1702
rect 6090 1668 6128 1702
rect 6162 1668 6200 1702
rect 6234 1668 6272 1702
rect 6306 1668 6344 1702
rect 6378 1668 6416 1702
rect 6450 1668 6488 1702
rect 6522 1668 6560 1702
rect 6594 1668 6632 1702
rect 6666 1668 6704 1702
rect 6738 1668 6776 1702
rect 6810 1668 6848 1702
rect 6882 1668 6920 1702
rect 6954 1668 6992 1702
rect 7026 1668 7064 1702
rect 7098 1668 7136 1702
rect 7170 1668 7208 1702
rect 7242 1668 7280 1702
rect 7314 1668 7352 1702
rect 7386 1668 7424 1702
rect 7458 1668 7496 1702
rect 7530 1668 7568 1702
rect 7602 1668 7640 1702
rect 7674 1668 7712 1702
rect 7746 1668 7784 1702
rect 7818 1668 7856 1702
rect 7890 1668 7928 1702
rect 7962 1668 8000 1702
rect 8034 1668 8072 1702
rect 8106 1668 8144 1702
rect 8178 1668 8216 1702
rect 8250 1668 8288 1702
rect 8322 1668 8360 1702
rect 8394 1668 8432 1702
rect 8466 1668 8504 1702
rect 8538 1668 8576 1702
rect 8610 1668 8648 1702
rect 8682 1668 8720 1702
rect 8754 1668 8792 1702
rect 8826 1668 8864 1702
rect 8898 1668 8936 1702
rect 8970 1668 9008 1702
rect 9042 1668 9080 1702
rect 9114 1668 9152 1702
rect 9186 1668 9224 1702
rect 9258 1668 9296 1702
rect 9330 1668 9368 1702
rect 9402 1668 9440 1702
rect 9474 1668 9512 1702
rect 9546 1668 9584 1702
rect 9618 1668 9656 1702
rect 9690 1668 9728 1702
rect 9762 1668 9800 1702
rect 9834 1668 9872 1702
rect 9906 1668 9944 1702
rect 9978 1668 10016 1702
rect 10050 1668 10088 1702
rect 10122 1668 10160 1702
rect 10194 1668 10232 1702
rect 10266 1668 10304 1702
rect 10338 1668 10376 1702
rect 10410 1668 10448 1702
rect 10482 1668 10520 1702
rect 10554 1668 10592 1702
rect 10626 1668 10664 1702
rect 10698 1668 10736 1702
rect 10770 1668 10808 1702
rect 10842 1668 10880 1702
rect 10914 1668 10952 1702
rect 10986 1668 11024 1702
rect 11058 1668 11096 1702
rect 11130 1668 11168 1702
rect 11202 1668 11240 1702
rect 11274 1668 11312 1702
rect 11346 1668 11384 1702
rect 11418 1668 11456 1702
rect 11490 1668 11528 1702
rect 11562 1668 11600 1702
rect 11634 1668 11672 1702
rect 11706 1668 11744 1702
rect 11778 1668 11816 1702
rect 11850 1668 11888 1702
rect 11922 1668 11960 1702
rect 11994 1668 12032 1702
rect 12066 1668 12104 1702
rect 12138 1668 12176 1702
rect 12210 1668 12248 1702
rect 12282 1668 12320 1702
rect 12354 1668 12392 1702
rect 12426 1668 12464 1702
rect 12498 1668 12536 1702
rect 12570 1668 12608 1702
rect 12642 1668 12680 1702
rect 12714 1668 12752 1702
rect 12786 1668 12824 1702
rect 12858 1668 12896 1702
rect 12930 1668 12968 1702
rect 13002 1668 13040 1702
rect 13074 1668 13112 1702
rect 13146 1668 13184 1702
rect 13218 1668 13256 1702
rect 13290 1668 13328 1702
rect 13362 1668 13400 1702
rect 13434 1668 13472 1702
rect 13506 1668 13544 1702
rect 13578 1668 13616 1702
rect 13650 1668 13688 1702
rect 13722 1668 13760 1702
rect 13794 1668 13832 1702
rect 13866 1668 13904 1702
rect 13938 1668 13976 1702
rect 14010 1668 14048 1702
rect 14082 1668 14120 1702
rect 14154 1668 14192 1702
rect 14226 1668 14264 1702
rect 14298 1668 14336 1702
rect 14370 1668 14408 1702
rect 14442 1668 14480 1702
rect 14514 1668 14552 1702
rect 14586 1668 14624 1702
rect 14658 1668 14696 1702
rect 14730 1668 14768 1702
rect 14802 1668 14840 1702
rect 14874 1668 14912 1702
rect 14946 1668 14984 1702
rect 15018 1668 15056 1702
rect 15090 1668 15128 1702
rect 15162 1668 15200 1702
rect 15234 1668 15272 1702
rect 15306 1668 15344 1702
rect 15378 1668 15416 1702
rect 15450 1668 15488 1702
rect 15522 1668 15561 1702
rect 15595 1668 15634 1702
rect 15668 1668 15707 1702
rect 15741 1668 15780 1702
rect 15814 1668 15853 1702
rect 15887 1668 15926 1702
rect 5711 1624 15944 1668
rect 5730 1590 5768 1624
rect 5802 1590 5840 1624
rect 5874 1590 5912 1624
rect 5946 1590 5984 1624
rect 6018 1590 6056 1624
rect 6090 1590 6128 1624
rect 6162 1590 6200 1624
rect 6234 1590 6272 1624
rect 6306 1590 6344 1624
rect 6378 1590 6416 1624
rect 6450 1590 6488 1624
rect 6522 1590 6560 1624
rect 6594 1590 6632 1624
rect 6666 1590 6704 1624
rect 6738 1590 6776 1624
rect 6810 1590 6848 1624
rect 6882 1590 6920 1624
rect 6954 1590 6992 1624
rect 7026 1590 7064 1624
rect 7098 1590 7136 1624
rect 7170 1590 7208 1624
rect 7242 1590 7280 1624
rect 7314 1590 7352 1624
rect 7386 1590 7424 1624
rect 7458 1590 7496 1624
rect 7530 1590 7568 1624
rect 7602 1590 7640 1624
rect 7674 1590 7712 1624
rect 7746 1590 7784 1624
rect 7818 1590 7856 1624
rect 7890 1590 7928 1624
rect 7962 1590 8000 1624
rect 8034 1590 8072 1624
rect 8106 1590 8144 1624
rect 8178 1590 8216 1624
rect 8250 1590 8288 1624
rect 8322 1590 8360 1624
rect 8394 1590 8432 1624
rect 8466 1590 8504 1624
rect 8538 1590 8576 1624
rect 8610 1590 8648 1624
rect 8682 1590 8720 1624
rect 8754 1590 8792 1624
rect 8826 1590 8864 1624
rect 8898 1590 8936 1624
rect 8970 1590 9008 1624
rect 9042 1590 9080 1624
rect 9114 1590 9152 1624
rect 9186 1590 9224 1624
rect 9258 1590 9296 1624
rect 9330 1590 9368 1624
rect 9402 1590 9440 1624
rect 9474 1590 9512 1624
rect 9546 1590 9584 1624
rect 9618 1590 9656 1624
rect 9690 1590 9728 1624
rect 9762 1590 9800 1624
rect 9834 1590 9872 1624
rect 9906 1590 9944 1624
rect 9978 1590 10016 1624
rect 10050 1590 10088 1624
rect 10122 1590 10160 1624
rect 10194 1590 10232 1624
rect 10266 1590 10304 1624
rect 10338 1590 10376 1624
rect 10410 1590 10448 1624
rect 10482 1590 10520 1624
rect 10554 1590 10592 1624
rect 10626 1590 10664 1624
rect 10698 1590 10736 1624
rect 10770 1590 10808 1624
rect 10842 1590 10880 1624
rect 10914 1590 10952 1624
rect 10986 1590 11024 1624
rect 11058 1590 11096 1624
rect 11130 1590 11168 1624
rect 11202 1590 11240 1624
rect 11274 1590 11312 1624
rect 11346 1590 11384 1624
rect 11418 1590 11456 1624
rect 11490 1590 11528 1624
rect 11562 1590 11600 1624
rect 11634 1590 11672 1624
rect 11706 1590 11744 1624
rect 11778 1590 11816 1624
rect 11850 1590 11888 1624
rect 11922 1590 11960 1624
rect 11994 1590 12032 1624
rect 12066 1590 12104 1624
rect 12138 1590 12176 1624
rect 12210 1590 12248 1624
rect 12282 1590 12320 1624
rect 12354 1590 12392 1624
rect 12426 1590 12464 1624
rect 12498 1590 12536 1624
rect 12570 1590 12608 1624
rect 12642 1590 12680 1624
rect 12714 1590 12752 1624
rect 12786 1590 12824 1624
rect 12858 1590 12896 1624
rect 12930 1590 12968 1624
rect 13002 1590 13040 1624
rect 13074 1590 13112 1624
rect 13146 1590 13184 1624
rect 13218 1590 13256 1624
rect 13290 1590 13328 1624
rect 13362 1590 13400 1624
rect 13434 1590 13472 1624
rect 13506 1590 13544 1624
rect 13578 1590 13616 1624
rect 13650 1590 13688 1624
rect 13722 1590 13760 1624
rect 13794 1590 13832 1624
rect 13866 1590 13904 1624
rect 13938 1590 13976 1624
rect 14010 1590 14048 1624
rect 14082 1590 14120 1624
rect 14154 1590 14192 1624
rect 14226 1590 14264 1624
rect 14298 1590 14336 1624
rect 14370 1590 14408 1624
rect 14442 1590 14480 1624
rect 14514 1590 14552 1624
rect 14586 1590 14624 1624
rect 14658 1590 14696 1624
rect 14730 1590 14768 1624
rect 14802 1590 14840 1624
rect 14874 1590 14912 1624
rect 14946 1590 14984 1624
rect 15018 1590 15056 1624
rect 15090 1590 15128 1624
rect 15162 1590 15200 1624
rect 15234 1590 15272 1624
rect 15306 1590 15344 1624
rect 15378 1590 15416 1624
rect 15450 1590 15488 1624
rect 15522 1590 15561 1624
rect 15595 1590 15634 1624
rect 15668 1590 15707 1624
rect 15741 1590 15780 1624
rect 15814 1590 15853 1624
rect 15887 1590 15926 1624
rect 5711 1546 15944 1590
rect 5730 1512 5768 1546
rect 5802 1512 5840 1546
rect 5874 1512 5912 1546
rect 5946 1512 5984 1546
rect 6018 1512 6056 1546
rect 6090 1512 6128 1546
rect 6162 1512 6200 1546
rect 6234 1512 6272 1546
rect 6306 1512 6344 1546
rect 6378 1512 6416 1546
rect 6450 1512 6488 1546
rect 6522 1512 6560 1546
rect 6594 1512 6632 1546
rect 6666 1512 6704 1546
rect 6738 1512 6776 1546
rect 6810 1512 6848 1546
rect 6882 1512 6920 1546
rect 6954 1512 6992 1546
rect 7026 1512 7064 1546
rect 7098 1512 7136 1546
rect 7170 1512 7208 1546
rect 7242 1512 7280 1546
rect 7314 1512 7352 1546
rect 7386 1512 7424 1546
rect 7458 1512 7496 1546
rect 7530 1512 7568 1546
rect 7602 1512 7640 1546
rect 7674 1512 7712 1546
rect 7746 1512 7784 1546
rect 7818 1512 7856 1546
rect 7890 1512 7928 1546
rect 7962 1512 8000 1546
rect 8034 1512 8072 1546
rect 8106 1512 8144 1546
rect 8178 1512 8216 1546
rect 8250 1512 8288 1546
rect 8322 1512 8360 1546
rect 8394 1512 8432 1546
rect 8466 1512 8504 1546
rect 8538 1512 8576 1546
rect 8610 1512 8648 1546
rect 8682 1512 8720 1546
rect 8754 1512 8792 1546
rect 8826 1512 8864 1546
rect 8898 1512 8936 1546
rect 8970 1512 9008 1546
rect 9042 1512 9080 1546
rect 9114 1512 9152 1546
rect 9186 1512 9224 1546
rect 9258 1512 9296 1546
rect 9330 1512 9368 1546
rect 9402 1512 9440 1546
rect 9474 1512 9512 1546
rect 9546 1512 9584 1546
rect 9618 1512 9656 1546
rect 9690 1512 9728 1546
rect 9762 1512 9800 1546
rect 9834 1512 9872 1546
rect 9906 1512 9944 1546
rect 9978 1512 10016 1546
rect 10050 1512 10088 1546
rect 10122 1512 10160 1546
rect 10194 1512 10232 1546
rect 10266 1512 10304 1546
rect 10338 1512 10376 1546
rect 10410 1512 10448 1546
rect 10482 1512 10520 1546
rect 10554 1512 10592 1546
rect 10626 1512 10664 1546
rect 10698 1512 10736 1546
rect 10770 1512 10808 1546
rect 10842 1512 10880 1546
rect 10914 1512 10952 1546
rect 10986 1512 11024 1546
rect 11058 1512 11096 1546
rect 11130 1512 11168 1546
rect 11202 1512 11240 1546
rect 11274 1512 11312 1546
rect 11346 1512 11384 1546
rect 11418 1512 11456 1546
rect 11490 1512 11528 1546
rect 11562 1512 11600 1546
rect 11634 1512 11672 1546
rect 11706 1512 11744 1546
rect 11778 1512 11816 1546
rect 11850 1512 11888 1546
rect 11922 1512 11960 1546
rect 11994 1512 12032 1546
rect 12066 1512 12104 1546
rect 12138 1512 12176 1546
rect 12210 1512 12248 1546
rect 12282 1512 12320 1546
rect 12354 1512 12392 1546
rect 12426 1512 12464 1546
rect 12498 1512 12536 1546
rect 12570 1512 12608 1546
rect 12642 1512 12680 1546
rect 12714 1512 12752 1546
rect 12786 1512 12824 1546
rect 12858 1512 12896 1546
rect 12930 1512 12968 1546
rect 13002 1512 13040 1546
rect 13074 1512 13112 1546
rect 13146 1512 13184 1546
rect 13218 1512 13256 1546
rect 13290 1512 13328 1546
rect 13362 1512 13400 1546
rect 13434 1512 13472 1546
rect 13506 1512 13544 1546
rect 13578 1512 13616 1546
rect 13650 1512 13688 1546
rect 13722 1512 13760 1546
rect 13794 1512 13832 1546
rect 13866 1512 13904 1546
rect 13938 1512 13976 1546
rect 14010 1512 14048 1546
rect 14082 1512 14120 1546
rect 14154 1512 14192 1546
rect 14226 1512 14264 1546
rect 14298 1512 14336 1546
rect 14370 1512 14408 1546
rect 14442 1512 14480 1546
rect 14514 1512 14552 1546
rect 14586 1512 14624 1546
rect 14658 1512 14696 1546
rect 14730 1512 14768 1546
rect 14802 1512 14840 1546
rect 14874 1512 14912 1546
rect 14946 1512 14984 1546
rect 15018 1512 15056 1546
rect 15090 1512 15128 1546
rect 15162 1512 15200 1546
rect 15234 1512 15272 1546
rect 15306 1512 15344 1546
rect 15378 1512 15416 1546
rect 15450 1512 15488 1546
rect 15522 1512 15561 1546
rect 15595 1512 15634 1546
rect 15668 1512 15707 1546
rect 15741 1512 15780 1546
rect 15814 1512 15853 1546
rect 15887 1512 15926 1546
rect 5711 1468 15944 1512
rect 5730 1434 5768 1468
rect 5802 1434 5840 1468
rect 5874 1434 5912 1468
rect 5946 1434 5984 1468
rect 6018 1434 6056 1468
rect 6090 1434 6128 1468
rect 6162 1434 6200 1468
rect 6234 1434 6272 1468
rect 6306 1434 6344 1468
rect 6378 1434 6416 1468
rect 6450 1434 6488 1468
rect 6522 1434 6560 1468
rect 6594 1434 6632 1468
rect 6666 1434 6704 1468
rect 6738 1434 6776 1468
rect 6810 1434 6848 1468
rect 6882 1434 6920 1468
rect 6954 1434 6992 1468
rect 7026 1434 7064 1468
rect 7098 1434 7136 1468
rect 7170 1434 7208 1468
rect 7242 1434 7280 1468
rect 7314 1434 7352 1468
rect 7386 1434 7424 1468
rect 7458 1434 7496 1468
rect 7530 1434 7568 1468
rect 7602 1434 7640 1468
rect 7674 1434 7712 1468
rect 7746 1434 7784 1468
rect 7818 1434 7856 1468
rect 7890 1434 7928 1468
rect 7962 1434 8000 1468
rect 8034 1434 8072 1468
rect 8106 1434 8144 1468
rect 8178 1434 8216 1468
rect 8250 1434 8288 1468
rect 8322 1434 8360 1468
rect 8394 1434 8432 1468
rect 8466 1434 8504 1468
rect 8538 1434 8576 1468
rect 8610 1434 8648 1468
rect 8682 1434 8720 1468
rect 8754 1434 8792 1468
rect 8826 1434 8864 1468
rect 8898 1434 8936 1468
rect 8970 1434 9008 1468
rect 9042 1434 9080 1468
rect 9114 1434 9152 1468
rect 9186 1434 9224 1468
rect 9258 1434 9296 1468
rect 9330 1434 9368 1468
rect 9402 1434 9440 1468
rect 9474 1434 9512 1468
rect 9546 1434 9584 1468
rect 9618 1434 9656 1468
rect 9690 1434 9728 1468
rect 9762 1434 9800 1468
rect 9834 1434 9872 1468
rect 9906 1434 9944 1468
rect 9978 1434 10016 1468
rect 10050 1434 10088 1468
rect 10122 1434 10160 1468
rect 10194 1434 10232 1468
rect 10266 1434 10304 1468
rect 10338 1434 10376 1468
rect 10410 1434 10448 1468
rect 10482 1434 10520 1468
rect 10554 1434 10592 1468
rect 10626 1434 10664 1468
rect 10698 1434 10736 1468
rect 10770 1434 10808 1468
rect 10842 1434 10880 1468
rect 10914 1434 10952 1468
rect 10986 1434 11024 1468
rect 11058 1434 11096 1468
rect 11130 1434 11168 1468
rect 11202 1434 11240 1468
rect 11274 1434 11312 1468
rect 11346 1434 11384 1468
rect 11418 1434 11456 1468
rect 11490 1434 11528 1468
rect 11562 1434 11600 1468
rect 11634 1434 11672 1468
rect 11706 1434 11744 1468
rect 11778 1434 11816 1468
rect 11850 1434 11888 1468
rect 11922 1434 11960 1468
rect 11994 1434 12032 1468
rect 12066 1434 12104 1468
rect 12138 1434 12176 1468
rect 12210 1434 12248 1468
rect 12282 1434 12320 1468
rect 12354 1434 12392 1468
rect 12426 1434 12464 1468
rect 12498 1434 12536 1468
rect 12570 1434 12608 1468
rect 12642 1434 12680 1468
rect 12714 1434 12752 1468
rect 12786 1434 12824 1468
rect 12858 1434 12896 1468
rect 12930 1434 12968 1468
rect 13002 1434 13040 1468
rect 13074 1434 13112 1468
rect 13146 1434 13184 1468
rect 13218 1434 13256 1468
rect 13290 1434 13328 1468
rect 13362 1434 13400 1468
rect 13434 1434 13472 1468
rect 13506 1434 13544 1468
rect 13578 1434 13616 1468
rect 13650 1434 13688 1468
rect 13722 1434 13760 1468
rect 13794 1434 13832 1468
rect 13866 1434 13904 1468
rect 13938 1434 13976 1468
rect 14010 1434 14048 1468
rect 14082 1434 14120 1468
rect 14154 1434 14192 1468
rect 14226 1434 14264 1468
rect 14298 1434 14336 1468
rect 14370 1434 14408 1468
rect 14442 1434 14480 1468
rect 14514 1434 14552 1468
rect 14586 1434 14624 1468
rect 14658 1434 14696 1468
rect 14730 1434 14768 1468
rect 14802 1434 14840 1468
rect 14874 1434 14912 1468
rect 14946 1434 14984 1468
rect 15018 1434 15056 1468
rect 15090 1434 15128 1468
rect 15162 1434 15200 1468
rect 15234 1434 15272 1468
rect 15306 1434 15344 1468
rect 15378 1434 15416 1468
rect 15450 1434 15488 1468
rect 15522 1434 15561 1468
rect 15595 1434 15634 1468
rect 15668 1434 15707 1468
rect 15741 1434 15780 1468
rect 15814 1434 15853 1468
rect 15887 1434 15926 1468
rect 5711 1433 15944 1434
rect 5711 1392 5947 1433
rect -1997 1200 -1962 1231
rect -1928 1200 -1893 1231
rect -1859 1200 -1824 1231
rect -1790 1200 -1755 1231
rect -1721 1200 -1686 1231
rect -1652 1200 -1617 1231
rect -1583 1200 -1548 1231
rect -1514 1200 -1479 1231
rect -1445 1200 -1410 1231
rect -1376 1200 -1341 1231
rect -1307 1200 -1272 1231
rect -1238 1200 -1203 1231
rect -1169 1200 -1134 1231
rect -1100 1200 -1065 1231
rect -1031 1200 -996 1231
rect -962 1200 -927 1231
rect -893 1200 -858 1231
rect -824 1200 -789 1231
rect -755 1200 -720 1231
rect -686 1200 -651 1231
rect -617 1200 -582 1231
rect -548 1200 -513 1231
rect -479 1200 -444 1231
rect -410 1200 -375 1231
rect -2859 1166 -375 1200
rect -2825 1132 -2790 1166
rect -2756 1132 -2721 1166
rect -2687 1132 -2652 1166
rect -2618 1132 -2583 1166
rect -2549 1132 -2514 1166
rect -2480 1132 -2445 1166
rect -2411 1132 -2376 1166
rect -2342 1132 -2307 1166
rect -2273 1132 -2238 1166
rect -2204 1132 -2169 1166
rect -2135 1132 -2100 1166
rect -2066 1132 -2031 1166
rect -1997 1132 -1962 1166
rect -1928 1132 -1893 1166
rect -1859 1132 -1824 1166
rect -1790 1132 -1755 1166
rect -1721 1132 -1686 1166
rect -1652 1132 -1617 1166
rect -1583 1132 -1548 1166
rect -1514 1132 -1479 1166
rect -1445 1132 -1410 1166
rect -1376 1132 -1341 1166
rect -1307 1132 -1272 1166
rect -1238 1132 -1203 1166
rect -1169 1132 -1134 1166
rect -1100 1132 -1065 1166
rect -1031 1132 -996 1166
rect -962 1132 -927 1166
rect -893 1132 -858 1166
rect -824 1132 -789 1166
rect -755 1132 -720 1166
rect -686 1132 -651 1166
rect -617 1132 -582 1166
rect -548 1132 -513 1166
rect -479 1132 -444 1166
rect -410 1132 -375 1166
rect -2859 1098 -375 1132
rect -2825 1064 -2790 1098
rect -2756 1064 -2721 1098
rect -2687 1064 -2652 1098
rect -2618 1064 -2583 1098
rect -2549 1064 -2514 1098
rect -2480 1064 -2445 1098
rect -2411 1064 -2376 1098
rect -2342 1064 -2307 1098
rect -2273 1064 -2238 1098
rect -2204 1064 -2169 1098
rect -2135 1064 -2100 1098
rect -2066 1064 -2031 1098
rect -1997 1064 -1962 1098
rect -1928 1064 -1893 1098
rect -1859 1064 -1824 1098
rect -1790 1064 -1755 1098
rect -1721 1064 -1686 1098
rect -1652 1064 -1617 1098
rect -1583 1064 -1548 1098
rect -1514 1064 -1479 1098
rect -1445 1064 -1410 1098
rect -1376 1064 -1341 1098
rect -1307 1064 -1272 1098
rect -1238 1064 -1203 1098
rect -1169 1064 -1134 1098
rect -1100 1064 -1065 1098
rect -1031 1064 -996 1098
rect -962 1064 -927 1098
rect -893 1064 -858 1098
rect -824 1064 -789 1098
rect -755 1064 -720 1098
rect -686 1064 -651 1098
rect -617 1064 -582 1098
rect -548 1064 -513 1098
rect -479 1064 -444 1098
rect -410 1064 -375 1098
rect -2859 1030 -375 1064
rect -2825 996 -2790 1030
rect -2756 996 -2721 1030
rect -2687 996 -2652 1030
rect -2618 996 -2583 1030
rect -2549 996 -2514 1030
rect -2480 996 -2445 1030
rect -2411 996 -2376 1030
rect -2342 996 -2307 1030
rect -2273 996 -2238 1030
rect -2204 996 -2169 1030
rect -2135 996 -2100 1030
rect -2066 996 -2031 1030
rect -1997 996 -1962 1030
rect -1928 996 -1893 1030
rect -1859 996 -1824 1030
rect -1790 996 -1755 1030
rect -1721 996 -1686 1030
rect -1652 996 -1617 1030
rect -1583 996 -1548 1030
rect -1514 996 -1479 1030
rect -1445 996 -1410 1030
rect -1376 996 -1341 1030
rect -1307 996 -1272 1030
rect -1238 996 -1203 1030
rect -1169 996 -1134 1030
rect -1100 996 -1065 1030
rect -1031 996 -996 1030
rect -962 996 -927 1030
rect -893 996 -858 1030
rect -824 996 -789 1030
rect -755 996 -720 1030
rect -686 996 -651 1030
rect -617 996 -582 1030
rect -548 996 -513 1030
rect -479 996 -444 1030
rect -410 996 -375 1030
rect -2859 962 -375 996
rect -2825 928 -2790 962
rect -2756 928 -2721 962
rect -2687 928 -2652 962
rect -2618 928 -2583 962
rect -2549 928 -2514 962
rect -2480 928 -2445 962
rect -2411 928 -2376 962
rect -2342 928 -2307 962
rect -2273 928 -2238 962
rect -2204 928 -2169 962
rect -2135 928 -2100 962
rect -2066 928 -2031 962
rect -1997 928 -1962 962
rect -1928 928 -1893 962
rect -1859 928 -1824 962
rect -1790 928 -1755 962
rect -1721 928 -1686 962
rect -1652 928 -1617 962
rect -1583 928 -1548 962
rect -1514 928 -1479 962
rect -1445 928 -1410 962
rect -1376 928 -1341 962
rect -1307 928 -1272 962
rect -1238 928 -1203 962
rect -1169 928 -1134 962
rect -1100 928 -1065 962
rect -1031 928 -996 962
rect -962 928 -927 962
rect -893 928 -858 962
rect -824 928 -789 962
rect -755 928 -720 962
rect -686 928 -651 962
rect -617 928 -582 962
rect -548 928 -513 962
rect -479 928 -444 962
rect -410 928 -375 962
rect -2859 894 -375 928
rect -2825 860 -2790 894
rect -2756 860 -2721 894
rect -2687 860 -2652 894
rect -2618 860 -2583 894
rect -2549 860 -2514 894
rect -2480 860 -2445 894
rect -2411 860 -2376 894
rect -2342 860 -2307 894
rect -2273 860 -2238 894
rect -2204 860 -2169 894
rect -2135 860 -2100 894
rect -2066 860 -2031 894
rect -1997 860 -1962 894
rect -1928 860 -1893 894
rect -1859 860 -1824 894
rect -1790 860 -1755 894
rect -1721 860 -1686 894
rect -1652 860 -1617 894
rect -1583 860 -1548 894
rect -1514 860 -1479 894
rect -1445 860 -1410 894
rect -1376 860 -1341 894
rect -1307 860 -1272 894
rect -1238 860 -1203 894
rect -1169 860 -1134 894
rect -1100 860 -1065 894
rect -1031 860 -996 894
rect -962 860 -927 894
rect -893 860 -858 894
rect -824 860 -789 894
rect -755 860 -720 894
rect -686 860 -651 894
rect -617 860 -582 894
rect -548 860 -513 894
rect -479 860 -444 894
rect -410 860 -375 894
rect -2859 826 -375 860
rect -2825 792 -2790 826
rect -2756 792 -2721 826
rect -2687 792 -2652 826
rect -2618 792 -2583 826
rect -2549 792 -2514 826
rect -2480 792 -2445 826
rect -2411 792 -2376 826
rect -2342 792 -2307 826
rect -2273 792 -2238 826
rect -2204 792 -2169 826
rect -2135 792 -2100 826
rect -2066 792 -2031 826
rect -1997 792 -1962 826
rect -1928 792 -1893 826
rect -1859 792 -1824 826
rect -1790 792 -1755 826
rect -1721 792 -1686 826
rect -1652 792 -1617 826
rect -1583 792 -1548 826
rect -1514 792 -1479 826
rect -1445 792 -1410 826
rect -1376 792 -1341 826
rect -1307 792 -1272 826
rect -1238 792 -1203 826
rect -1169 792 -1134 826
rect -1100 792 -1065 826
rect -1031 792 -996 826
rect -962 792 -927 826
rect -893 792 -858 826
rect -824 792 -789 826
rect -755 792 -720 826
rect -686 792 -651 826
rect -617 792 -582 826
rect -548 792 -513 826
rect -479 792 -444 826
rect -410 792 -375 826
rect -1 792 33 1231
rect 5711 1358 5736 1392
rect 5770 1358 5809 1392
rect 5843 1358 5882 1392
rect 5916 1358 5947 1392
rect 5711 1320 5947 1358
rect 5711 1286 5736 1320
rect 5770 1286 5809 1320
rect 5843 1286 5882 1320
rect 5916 1286 5947 1320
rect 5711 1248 5947 1286
rect 15540 1393 15944 1433
rect 16726 1393 17215 2159
rect 15540 1359 15560 1393
rect 15594 1359 15633 1393
rect 15667 1359 15706 1393
rect 15740 1359 15779 1393
rect 15813 1359 15852 1393
rect 15886 1359 15925 1393
rect 16726 1359 16732 1393
rect 16766 1359 16806 1393
rect 16840 1359 16880 1393
rect 16914 1359 17215 1393
rect 15540 1319 15944 1359
rect 16726 1319 17215 1359
rect 15540 1285 15560 1319
rect 15594 1285 15633 1319
rect 15667 1285 15706 1319
rect 15740 1285 15779 1319
rect 15813 1285 15852 1319
rect 15886 1285 15925 1319
rect 16726 1285 16732 1319
rect 16766 1285 16806 1319
rect 16840 1285 16880 1319
rect 16914 1285 17215 1319
rect 5711 1214 5736 1248
rect 5770 1214 5809 1248
rect 5843 1214 5882 1248
rect 5916 1214 5947 1248
rect 5711 792 5947 1214
rect 10199 1236 10267 1270
rect 10301 1236 10335 1270
rect 10369 1236 10403 1270
rect 10437 1236 10471 1270
rect 10505 1236 10539 1270
rect 10573 1236 10607 1270
rect 10641 1236 10675 1270
rect 10709 1236 10743 1270
rect 10777 1236 10811 1270
rect 10845 1236 10879 1270
rect 10913 1236 10947 1270
rect 10981 1236 11015 1270
rect 11049 1236 11083 1270
rect 11117 1236 11151 1270
rect 11185 1236 11219 1270
rect 11253 1236 11287 1270
rect 11321 1236 11355 1270
rect 11389 1236 11423 1270
rect 11457 1236 11491 1270
rect 11525 1236 11559 1270
rect 11593 1236 11627 1270
rect 11661 1236 11695 1270
rect 11729 1236 11763 1270
rect 11797 1236 11831 1270
rect 11865 1236 11899 1270
rect 11933 1236 11967 1270
rect 12001 1236 12035 1270
rect 12069 1236 12103 1270
rect 12137 1236 12171 1270
rect 12205 1236 12239 1270
rect 12273 1236 12307 1270
rect 12341 1236 12375 1270
rect 12409 1236 12443 1270
rect 12477 1236 12511 1270
rect 12545 1236 12579 1270
rect 12613 1236 12647 1270
rect 12681 1236 12715 1270
rect 12749 1236 12783 1270
rect 12817 1236 12851 1270
rect 12885 1236 12919 1270
rect 12953 1236 12987 1270
rect 13021 1236 13055 1270
rect 13089 1236 13123 1270
rect 13157 1236 13191 1270
rect 13225 1236 13259 1270
rect 13293 1236 13327 1270
rect 13361 1236 13395 1270
rect 13429 1236 13463 1270
rect 13497 1236 13531 1270
rect 13565 1236 13599 1270
rect 13633 1236 13667 1270
rect 13701 1236 13735 1270
rect 13769 1236 13803 1270
rect 13837 1236 13871 1270
rect 13905 1236 13939 1270
rect 13973 1236 14007 1270
rect 14041 1236 14076 1270
rect 14110 1236 14145 1270
rect 14179 1236 14214 1270
rect 14248 1236 14283 1270
rect 14317 1236 14352 1270
rect 14386 1236 14421 1270
rect 14455 1236 14490 1270
rect 14524 1236 14559 1270
rect 14593 1236 14628 1270
rect 14662 1236 14697 1270
rect 14731 1236 14766 1270
rect 14800 1236 14835 1270
rect 14869 1236 14904 1270
rect 14938 1236 14973 1270
rect 15007 1236 15042 1270
rect 15076 1236 15111 1270
rect 15145 1236 15180 1270
rect 15214 1236 15249 1270
rect 15283 1236 15318 1270
rect 15352 1236 15420 1270
rect 10199 1201 15420 1236
rect 10199 1167 15386 1201
rect 10199 1161 15420 1167
rect -2859 768 5947 792
rect 2162 543 5947 768
rect 6202 1127 6270 1161
rect 6304 1127 6338 1161
rect 6372 1127 6406 1161
rect 6440 1127 6474 1161
rect 6508 1127 6542 1161
rect 6576 1127 6611 1161
rect 6645 1127 6680 1161
rect 6714 1127 6749 1161
rect 6783 1127 6818 1161
rect 6852 1127 6887 1161
rect 6921 1127 6956 1161
rect 6990 1127 7025 1161
rect 7059 1127 7094 1161
rect 7128 1127 7163 1161
rect 7197 1127 7232 1161
rect 7266 1127 7301 1161
rect 7335 1127 7370 1161
rect 7404 1127 7439 1161
rect 7473 1127 7508 1161
rect 7542 1127 7577 1161
rect 7611 1127 7646 1161
rect 7680 1127 7715 1161
rect 7749 1127 7784 1161
rect 7818 1127 7853 1161
rect 7887 1127 7922 1161
rect 7956 1127 7991 1161
rect 8025 1127 8060 1161
rect 8094 1127 8129 1161
rect 8163 1127 8198 1161
rect 8232 1127 8267 1161
rect 8301 1127 8336 1161
rect 8370 1127 8405 1161
rect 8439 1127 8474 1161
rect 8508 1127 8543 1161
rect 8577 1127 8612 1161
rect 8646 1127 8681 1161
rect 8715 1127 8750 1161
rect 8784 1127 8819 1161
rect 8853 1127 8888 1161
rect 8922 1127 8957 1161
rect 8991 1127 9026 1161
rect 9060 1127 9095 1161
rect 9129 1127 9164 1161
rect 9198 1127 9233 1161
rect 9267 1127 9302 1161
rect 9336 1127 9371 1161
rect 9405 1127 9440 1161
rect 9474 1127 9509 1161
rect 9543 1127 9578 1161
rect 9612 1127 9647 1161
rect 9681 1127 9716 1161
rect 9750 1127 9785 1161
rect 9819 1127 9854 1161
rect 9888 1127 9923 1161
rect 9957 1127 9992 1161
rect 10026 1127 10061 1161
rect 10095 1127 10130 1161
rect 10164 1127 10199 1161
rect 10233 1144 15420 1161
rect 10233 1127 10393 1144
rect 6202 1124 10393 1127
rect 6202 1093 10325 1124
rect 6236 1090 10325 1093
rect 10359 1110 10393 1124
rect 10427 1110 10461 1144
rect 10495 1110 10529 1144
rect 10563 1110 10597 1144
rect 10631 1110 10665 1144
rect 10699 1110 10733 1144
rect 10767 1110 10801 1144
rect 10835 1110 10869 1144
rect 10903 1110 10937 1144
rect 10971 1110 11005 1144
rect 11039 1110 11073 1144
rect 11107 1110 11141 1144
rect 11175 1110 11209 1144
rect 11243 1110 11277 1144
rect 11311 1110 11345 1144
rect 11379 1110 11413 1144
rect 11447 1110 11481 1144
rect 11515 1110 11549 1144
rect 11583 1110 11617 1144
rect 11651 1110 11685 1144
rect 11719 1110 11753 1144
rect 11787 1110 11821 1144
rect 11855 1110 11889 1144
rect 11923 1110 11957 1144
rect 11991 1110 12025 1144
rect 12059 1110 12093 1144
rect 12127 1110 12161 1144
rect 12195 1110 12229 1144
rect 12263 1110 12297 1144
rect 12331 1110 12365 1144
rect 12399 1110 12433 1144
rect 12467 1110 12501 1144
rect 12535 1110 12569 1144
rect 12603 1110 12638 1144
rect 12672 1110 12707 1144
rect 12741 1110 12776 1144
rect 12810 1110 12845 1144
rect 12879 1110 12914 1144
rect 12948 1110 12983 1144
rect 13017 1110 13052 1144
rect 13086 1110 13121 1144
rect 13155 1110 13190 1144
rect 13224 1110 13259 1144
rect 13293 1110 13328 1144
rect 13362 1110 13397 1144
rect 13431 1110 13466 1144
rect 13500 1110 13535 1144
rect 13569 1110 13604 1144
rect 13638 1110 13673 1144
rect 13707 1110 13742 1144
rect 13776 1110 13811 1144
rect 13845 1110 13880 1144
rect 13914 1110 13949 1144
rect 13983 1110 14018 1144
rect 14052 1110 14087 1144
rect 14121 1110 14156 1144
rect 14190 1110 14225 1144
rect 14259 1110 14294 1144
rect 14328 1110 14363 1144
rect 14397 1110 14432 1144
rect 14466 1110 14501 1144
rect 14535 1110 14570 1144
rect 14604 1110 14639 1144
rect 14673 1110 14708 1144
rect 14742 1110 14777 1144
rect 14811 1110 14846 1144
rect 14880 1110 14915 1144
rect 14949 1110 14984 1144
rect 15018 1110 15053 1144
rect 15087 1110 15122 1144
rect 15156 1110 15191 1144
rect 15225 1110 15260 1144
rect 15294 1132 15420 1144
rect 15294 1110 15386 1132
rect 6236 1059 10359 1090
rect 6202 1035 10359 1059
rect 6202 1018 6328 1035
rect 6236 1001 6328 1018
rect 6362 1001 6396 1035
rect 6430 1001 6464 1035
rect 6498 1001 6532 1035
rect 6566 1001 6600 1035
rect 6634 1001 6669 1035
rect 6703 1001 6738 1035
rect 6772 1001 6807 1035
rect 6841 1001 6876 1035
rect 6910 1001 6945 1035
rect 6979 1001 7014 1035
rect 7048 1001 7083 1035
rect 7117 1001 7152 1035
rect 7186 1001 7221 1035
rect 7255 1001 7290 1035
rect 7324 1001 7359 1035
rect 7393 1001 7428 1035
rect 7462 1001 7497 1035
rect 7531 1001 7566 1035
rect 7600 1001 7635 1035
rect 7669 1001 7704 1035
rect 7738 1001 7773 1035
rect 7807 1001 7842 1035
rect 7876 1001 7911 1035
rect 7945 1001 7980 1035
rect 8014 1001 8049 1035
rect 8083 1001 8118 1035
rect 8152 1001 8187 1035
rect 8221 1001 8256 1035
rect 8290 1001 8325 1035
rect 8359 1001 8394 1035
rect 8428 1001 8463 1035
rect 8497 1001 8532 1035
rect 8566 1001 8601 1035
rect 8635 1001 8670 1035
rect 8704 1001 8739 1035
rect 8773 1001 8808 1035
rect 8842 1001 8877 1035
rect 8911 1001 8946 1035
rect 8980 1001 9015 1035
rect 9049 1001 9084 1035
rect 9118 1001 9153 1035
rect 9187 1001 9222 1035
rect 9256 1001 9291 1035
rect 9325 1001 9360 1035
rect 9394 1001 9429 1035
rect 9463 1001 9498 1035
rect 9532 1001 9567 1035
rect 9601 1001 9636 1035
rect 9670 1001 9705 1035
rect 9739 1001 9774 1035
rect 9808 1001 9843 1035
rect 9877 1001 9912 1035
rect 9946 1001 9981 1035
rect 10015 1001 10050 1035
rect 10084 1001 10119 1035
rect 10153 1001 10188 1035
rect 10222 1001 10257 1035
rect 10291 1001 10359 1035
rect 15260 1098 15386 1110
rect 15260 1074 15420 1098
rect 15294 1063 15420 1074
rect 15294 1040 15386 1063
rect 15260 1029 15386 1040
rect 15260 1003 15420 1029
rect 6236 984 6362 1001
rect 6202 957 6362 984
rect 15294 994 15420 1003
rect 15294 969 15386 994
rect 15260 960 15386 969
rect 6202 943 6328 957
rect 6236 923 6328 943
rect 6236 909 6362 923
rect 6202 880 6362 909
rect 6202 868 6328 880
rect 6236 846 6328 868
rect 6236 834 6362 846
rect 10528 950 14944 957
rect 10528 916 10596 950
rect 10630 916 10665 950
rect 10699 916 10734 950
rect 10768 916 10803 950
rect 10837 916 10872 950
rect 10906 916 10941 950
rect 10975 916 11010 950
rect 11044 916 11078 950
rect 11112 916 11146 950
rect 11180 916 11214 950
rect 11248 916 11282 950
rect 11316 916 11350 950
rect 11384 916 11418 950
rect 11452 916 11486 950
rect 11520 916 11554 950
rect 11588 916 11622 950
rect 11656 916 11690 950
rect 11724 916 11758 950
rect 11792 916 11826 950
rect 11860 916 11894 950
rect 11928 916 11962 950
rect 11996 916 12030 950
rect 12064 916 12098 950
rect 12132 916 12166 950
rect 12200 916 12234 950
rect 12268 916 12302 950
rect 12336 916 12370 950
rect 12404 916 12438 950
rect 12472 916 12506 950
rect 12540 916 12574 950
rect 12608 916 12642 950
rect 12676 916 12710 950
rect 12744 916 12778 950
rect 12812 916 12846 950
rect 12880 916 12914 950
rect 12948 916 12982 950
rect 13016 916 13050 950
rect 13084 916 13118 950
rect 13152 916 13186 950
rect 13220 916 13254 950
rect 13288 916 13322 950
rect 13356 916 13390 950
rect 13424 916 13458 950
rect 13492 916 13526 950
rect 13560 916 13594 950
rect 13628 916 13662 950
rect 13696 916 13730 950
rect 13764 916 13798 950
rect 13832 916 13866 950
rect 13900 916 13934 950
rect 13968 916 14002 950
rect 14036 916 14070 950
rect 14104 916 14138 950
rect 14172 916 14206 950
rect 14240 916 14274 950
rect 14308 916 14342 950
rect 14376 916 14410 950
rect 14444 916 14478 950
rect 14512 916 14546 950
rect 14580 916 14614 950
rect 14648 916 14682 950
rect 14716 916 14750 950
rect 14784 916 14818 950
rect 14852 916 14886 950
rect 14920 916 14944 950
rect 10528 909 14944 916
rect 15260 932 15420 960
rect 10528 839 10737 909
rect 6202 803 6362 834
rect 6202 793 6328 803
rect 6236 769 6328 793
rect 6552 832 10737 839
rect 6552 798 6576 832
rect 6610 798 6645 832
rect 6679 798 6714 832
rect 6748 798 6783 832
rect 6817 798 6852 832
rect 6886 798 6921 832
rect 6955 798 6990 832
rect 7024 798 7059 832
rect 7093 798 7128 832
rect 7162 798 7197 832
rect 7231 798 7266 832
rect 7300 798 7335 832
rect 7369 798 7404 832
rect 7438 798 7473 832
rect 7507 798 7542 832
rect 7576 798 7611 832
rect 7645 798 7680 832
rect 7714 798 7749 832
rect 7783 798 7818 832
rect 7852 798 7887 832
rect 7921 798 7956 832
rect 7990 798 8025 832
rect 8059 798 8094 832
rect 8128 798 8162 832
rect 8196 798 8230 832
rect 8264 798 8298 832
rect 8332 798 8366 832
rect 8400 798 8434 832
rect 8468 798 8502 832
rect 8536 798 8570 832
rect 8604 798 8638 832
rect 8672 813 8706 832
rect 8740 813 8774 832
rect 8808 813 8842 832
rect 8876 813 8910 832
rect 8944 813 8978 832
rect 8678 798 8706 813
rect 8752 798 8774 813
rect 8826 798 8842 813
rect 8900 798 8910 813
rect 8974 798 8978 813
rect 9012 813 9046 832
rect 9080 813 9114 832
rect 9148 813 9182 832
rect 9216 813 9250 832
rect 9284 813 9318 832
rect 9352 813 9386 832
rect 9012 798 9014 813
rect 9080 798 9088 813
rect 9148 798 9162 813
rect 9216 798 9236 813
rect 9284 798 9310 813
rect 9352 798 9384 813
rect 9420 798 9454 832
rect 9488 813 9522 832
rect 9556 813 9590 832
rect 9624 813 9658 832
rect 9692 813 9726 832
rect 9760 813 9794 832
rect 9828 813 9862 832
rect 9492 798 9522 813
rect 9566 798 9590 813
rect 9640 798 9658 813
rect 9714 798 9726 813
rect 9788 798 9794 813
rect 9861 798 9862 813
rect 9896 813 9930 832
rect 9964 813 9998 832
rect 10032 813 10066 832
rect 10100 813 10134 832
rect 10168 813 10202 832
rect 10236 813 10270 832
rect 9896 798 9900 813
rect 9964 798 9973 813
rect 10032 798 10046 813
rect 10100 798 10119 813
rect 10168 798 10192 813
rect 10236 798 10265 813
rect 10304 798 10338 832
rect 10372 798 10406 832
rect 10440 813 10474 832
rect 10508 813 10737 832
rect 10445 798 10474 813
rect 6552 791 8644 798
rect 6236 759 6362 769
rect 6202 726 6362 759
rect 8678 779 8718 798
rect 8752 779 8792 798
rect 8826 779 8866 798
rect 8900 779 8940 798
rect 8974 779 9014 798
rect 9048 779 9088 798
rect 9122 779 9162 798
rect 9196 779 9236 798
rect 9270 779 9310 798
rect 9344 779 9384 798
rect 9418 779 9458 798
rect 9492 779 9532 798
rect 9566 779 9606 798
rect 9640 779 9680 798
rect 9714 779 9754 798
rect 9788 779 9827 798
rect 9861 779 9900 798
rect 9934 779 9973 798
rect 10007 779 10046 798
rect 10080 779 10119 798
rect 10153 779 10192 798
rect 10226 779 10265 798
rect 10299 779 10338 798
rect 10372 779 10411 798
rect 10445 779 10484 798
rect 10518 779 10557 813
rect 10591 779 10630 813
rect 10664 779 10703 813
rect 15294 925 15420 932
rect 15294 898 15386 925
rect 15260 891 15386 898
rect 15260 861 15420 891
rect 15294 856 15420 861
rect 15294 827 15386 856
rect 15260 822 15386 827
rect 8644 755 10737 779
rect 14716 760 14754 794
rect 15260 790 15420 822
rect 6202 718 6328 726
rect 6236 692 6328 718
rect 6236 684 6362 692
rect 6202 649 6362 684
rect 6567 674 6579 708
rect 6617 674 6652 708
rect 6693 674 6721 708
rect 6773 674 6790 708
rect 6852 674 6859 708
rect 6893 674 6928 708
rect 6962 674 6997 708
rect 7031 674 7066 708
rect 7100 674 7135 708
rect 7169 674 7204 708
rect 7238 674 7273 708
rect 7307 674 7342 708
rect 7376 674 7411 708
rect 7445 674 7480 708
rect 7514 674 7549 708
rect 7583 674 7618 708
rect 7652 674 7687 708
rect 7721 674 7756 708
rect 7790 674 7824 708
rect 7858 674 7892 708
rect 7926 674 7960 708
rect 7994 674 8028 708
rect 8062 674 8096 708
rect 8130 674 8164 708
rect 8198 674 8232 708
rect 8266 674 8300 708
rect 8334 674 8368 708
rect 8402 674 8436 708
rect 8470 674 8504 708
rect 8538 674 8572 708
rect 8606 674 8640 708
rect 8674 674 8708 708
rect 8742 674 8776 708
rect 8810 674 8844 708
rect 8878 674 8912 708
rect 8946 674 8980 708
rect 9014 674 9048 708
rect 9082 674 9116 708
rect 9150 674 9184 708
rect 9218 674 9252 708
rect 9286 674 9320 708
rect 9354 674 9388 708
rect 9422 674 9456 708
rect 9490 674 9524 708
rect 9558 674 9592 708
rect 9626 674 9660 708
rect 9694 674 9728 708
rect 9762 674 9796 708
rect 9830 674 9864 708
rect 9898 674 9932 708
rect 9966 674 10000 708
rect 10034 674 10068 708
rect 10102 674 10136 708
rect 10170 674 10204 708
rect 10238 674 10272 708
rect 10306 674 10340 708
rect 10374 674 10408 708
rect 10442 674 10476 708
rect 10510 674 10526 708
rect 6202 643 6328 649
rect 6236 615 6328 643
rect 6236 609 6362 615
rect 6202 572 6362 609
rect 6556 596 6594 630
rect 6202 569 6328 572
rect 6236 538 6328 569
rect 6236 535 6362 538
rect 6202 495 6362 535
rect 6236 461 6328 495
rect 6202 380 6362 461
rect 10345 489 10478 674
rect 10578 539 10737 755
rect 15294 786 15420 790
rect 15294 756 15386 786
rect 15260 752 15386 756
rect 15260 719 15420 752
rect 10785 674 10801 708
rect 10835 674 10870 708
rect 10904 674 10939 708
rect 10973 674 11008 708
rect 11042 674 11077 708
rect 11111 674 11146 708
rect 11180 674 11215 708
rect 11249 674 11284 708
rect 11318 674 11353 708
rect 11387 674 11422 708
rect 11456 674 11491 708
rect 11525 674 11560 708
rect 11594 674 11629 708
rect 11663 674 11698 708
rect 11732 674 11767 708
rect 11801 674 11836 708
rect 11870 674 11905 708
rect 11939 674 11974 708
rect 12008 674 12043 708
rect 12077 674 12112 708
rect 12146 674 12181 708
rect 12215 674 12250 708
rect 12284 674 12318 708
rect 12352 674 12386 708
rect 12420 674 12454 708
rect 12488 674 12522 708
rect 12556 674 12590 708
rect 12624 674 12658 708
rect 12692 674 12726 708
rect 12760 674 12794 708
rect 12828 674 12862 708
rect 12896 674 12930 708
rect 12964 674 12998 708
rect 13032 674 13066 708
rect 13100 674 13134 708
rect 13168 674 13202 708
rect 13236 674 13270 708
rect 13304 674 13338 708
rect 13372 674 13406 708
rect 13440 674 13474 708
rect 13508 674 13542 708
rect 13576 674 13610 708
rect 13644 674 13678 708
rect 13712 674 13746 708
rect 13780 674 13814 708
rect 13848 674 13882 708
rect 13916 674 13950 708
rect 13984 674 14018 708
rect 14052 674 14086 708
rect 14120 674 14154 708
rect 14188 674 14222 708
rect 14256 674 14290 708
rect 14324 674 14358 708
rect 14392 674 14426 708
rect 14460 674 14494 708
rect 14528 674 14562 708
rect 14596 674 14630 708
rect 14664 674 14698 708
rect 14732 674 14748 708
rect 15294 716 15420 719
rect 15294 685 15386 716
rect 15260 682 15386 685
rect 10883 489 11024 674
rect 15260 648 15420 682
rect 15294 646 15420 648
rect 15294 614 15386 646
rect 15260 612 15386 614
rect 14716 562 14754 596
rect 15260 577 15420 612
rect 10345 432 11024 489
rect 15294 576 15420 577
rect 15294 543 15386 576
rect 15260 542 15386 543
rect 15540 1245 15944 1285
rect 16726 1245 17215 1285
rect 15540 1211 15560 1245
rect 15594 1211 15633 1245
rect 15667 1211 15706 1245
rect 15740 1211 15779 1245
rect 15813 1211 15852 1245
rect 15886 1211 15925 1245
rect 16726 1211 16732 1245
rect 16766 1211 16806 1245
rect 16840 1211 16880 1245
rect 16914 1211 17215 1245
rect 15540 808 15944 1211
rect 15540 542 15648 808
rect 15260 506 15420 542
rect 15294 472 15386 506
rect 15260 381 15420 472
rect 15541 -1314 15648 542
rect 16726 -123 17215 1211
rect 15541 -1353 15944 -1314
rect 15541 -1387 15648 -1353
rect 15682 -1387 15720 -1353
rect 15754 -1387 15792 -1353
rect 15826 -1387 15864 -1353
rect 15898 -1387 15936 -1353
rect 15541 -1426 15944 -1387
rect 15541 -1460 15648 -1426
rect 15682 -1460 15720 -1426
rect 15754 -1460 15792 -1426
rect 15826 -1460 15864 -1426
rect 15898 -1460 15936 -1426
rect 15541 -1499 15944 -1460
rect 15541 -1533 15648 -1499
rect 15682 -1533 15720 -1499
rect 15754 -1533 15792 -1499
rect 15826 -1533 15864 -1499
rect 15898 -1533 15936 -1499
rect 15541 -1572 15944 -1533
rect 15541 -1606 15648 -1572
rect 15682 -1606 15720 -1572
rect 15754 -1606 15792 -1572
rect 15826 -1606 15864 -1572
rect 15898 -1606 15936 -1572
rect 15541 -1645 15944 -1606
rect 15541 -1679 15648 -1645
rect 15682 -1679 15720 -1645
rect 15754 -1679 15792 -1645
rect 15826 -1679 15864 -1645
rect 15898 -1679 15936 -1645
rect 15541 -2076 15944 -1679
rect 15332 -2278 15944 -2076
rect 15938 -2511 15944 -2278
rect 16726 -2511 16732 -123
rect 15938 -2546 16732 -2511
rect 15938 -2580 15944 -2546
rect 15978 -2580 16012 -2546
rect 16046 -2580 16080 -2546
rect 16114 -2580 16148 -2546
rect 16182 -2580 16216 -2546
rect 16250 -2580 16284 -2546
rect 16318 -2580 16352 -2546
rect 16386 -2580 16420 -2546
rect 16454 -2580 16488 -2546
rect 16522 -2580 16556 -2546
rect 16590 -2580 16624 -2546
rect 16658 -2580 16692 -2546
rect 16726 -2580 16732 -2546
rect 15938 -2615 16732 -2580
rect 15938 -2649 15944 -2615
rect 15978 -2649 16012 -2615
rect 16046 -2649 16080 -2615
rect 16114 -2649 16148 -2615
rect 16182 -2649 16216 -2615
rect 16250 -2649 16284 -2615
rect 16318 -2649 16352 -2615
rect 16386 -2649 16420 -2615
rect 16454 -2649 16488 -2615
rect 16522 -2649 16556 -2615
rect 16590 -2649 16624 -2615
rect 16658 -2649 16692 -2615
rect 16726 -2649 16732 -2615
rect 15938 -2684 16732 -2649
rect 15938 -2718 15944 -2684
rect 15978 -2718 16012 -2684
rect 16046 -2718 16080 -2684
rect 16114 -2718 16148 -2684
rect 16182 -2718 16216 -2684
rect 16250 -2718 16284 -2684
rect 16318 -2718 16352 -2684
rect 16386 -2718 16420 -2684
rect 16454 -2718 16488 -2684
rect 16522 -2718 16556 -2684
rect 16590 -2718 16624 -2684
rect 16658 -2718 16692 -2684
rect 16726 -2718 16732 -2684
rect 15938 -2753 16732 -2718
rect 15938 -2787 15944 -2753
rect 15978 -2787 16012 -2753
rect 16046 -2787 16080 -2753
rect 16114 -2787 16148 -2753
rect 16182 -2787 16216 -2753
rect 16250 -2787 16284 -2753
rect 16318 -2787 16352 -2753
rect 16386 -2787 16420 -2753
rect 16454 -2787 16488 -2753
rect 16522 -2787 16556 -2753
rect 16590 -2787 16624 -2753
rect 16658 -2787 16692 -2753
rect 16726 -2787 16732 -2753
rect 15938 -2822 16732 -2787
rect 15938 -2856 15944 -2822
rect 15978 -2856 16012 -2822
rect 16046 -2856 16080 -2822
rect 16114 -2856 16148 -2822
rect 16182 -2856 16216 -2822
rect 16250 -2856 16284 -2822
rect 16318 -2856 16352 -2822
rect 16386 -2856 16420 -2822
rect 16454 -2856 16488 -2822
rect 16522 -2856 16556 -2822
rect 16590 -2856 16624 -2822
rect 16658 -2856 16692 -2822
rect 16726 -2856 16732 -2822
rect 15938 -2891 16732 -2856
rect 15938 -2925 15944 -2891
rect 15978 -2925 16012 -2891
rect 16046 -2925 16080 -2891
rect 16114 -2925 16148 -2891
rect 16182 -2925 16216 -2891
rect 16250 -2925 16284 -2891
rect 16318 -2925 16352 -2891
rect 16386 -2925 16420 -2891
rect 16454 -2925 16488 -2891
rect 16522 -2925 16556 -2891
rect 16590 -2925 16624 -2891
rect 16658 -2925 16692 -2891
rect 16726 -2925 16732 -2891
rect 15938 -2949 16732 -2925
rect 15939 -2975 16732 -2949
<< viali >>
rect 3891 4494 3908 4501
rect 3908 4494 3925 4501
rect 3967 4494 3977 4501
rect 3977 4494 4001 4501
rect 4043 4494 4046 4501
rect 4046 4494 4077 4501
rect 4119 4494 4149 4501
rect 4149 4494 4153 4501
rect 4195 4494 4218 4501
rect 4218 4494 4229 4501
rect 4271 4494 4287 4501
rect 4287 4494 4305 4501
rect 4347 4494 4356 4501
rect 4356 4494 4381 4501
rect 4423 4494 4425 4501
rect 4425 4494 4457 4501
rect 3891 4467 3925 4494
rect 3967 4467 4001 4494
rect 4043 4467 4077 4494
rect 4119 4467 4153 4494
rect 4195 4467 4229 4494
rect 4271 4467 4305 4494
rect 4347 4467 4381 4494
rect 4423 4467 4457 4494
rect 4499 4467 4533 4501
rect 3891 4392 3925 4425
rect 3967 4392 4001 4425
rect 4043 4392 4077 4425
rect 4119 4392 4153 4425
rect 4195 4392 4229 4425
rect 4271 4392 4305 4425
rect 4347 4392 4381 4425
rect 4423 4392 4457 4425
rect 3891 4391 3908 4392
rect 3908 4391 3925 4392
rect 3967 4391 3977 4392
rect 3977 4391 4001 4392
rect 4043 4391 4046 4392
rect 4046 4391 4077 4392
rect 4119 4391 4149 4392
rect 4149 4391 4153 4392
rect 4195 4391 4218 4392
rect 4218 4391 4229 4392
rect 4271 4391 4287 4392
rect 4287 4391 4305 4392
rect 4347 4391 4356 4392
rect 4356 4391 4381 4392
rect 4423 4391 4425 4392
rect 4425 4391 4457 4392
rect 4499 4391 4533 4425
rect 3891 4324 3925 4349
rect 3967 4324 4001 4349
rect 4043 4324 4077 4349
rect 4119 4324 4153 4349
rect 4195 4324 4229 4349
rect 4271 4324 4305 4349
rect 4347 4324 4381 4349
rect 4423 4324 4457 4349
rect 3891 4315 3908 4324
rect 3908 4315 3925 4324
rect 3967 4315 3977 4324
rect 3977 4315 4001 4324
rect 4043 4315 4046 4324
rect 4046 4315 4077 4324
rect 4119 4315 4149 4324
rect 4149 4315 4153 4324
rect 4195 4315 4218 4324
rect 4218 4315 4229 4324
rect 4271 4315 4287 4324
rect 4287 4315 4305 4324
rect 4347 4315 4356 4324
rect 4356 4315 4381 4324
rect 4423 4315 4425 4324
rect 4425 4315 4457 4324
rect 4499 4315 4533 4349
rect 3891 4256 3925 4273
rect 3967 4256 4001 4273
rect 4043 4256 4077 4273
rect 4119 4256 4153 4273
rect 4195 4256 4229 4273
rect 4271 4256 4305 4273
rect 4347 4256 4381 4273
rect 4423 4256 4457 4273
rect 3891 4239 3908 4256
rect 3908 4239 3925 4256
rect 3967 4239 3977 4256
rect 3977 4239 4001 4256
rect 4043 4239 4046 4256
rect 4046 4239 4077 4256
rect 4119 4239 4149 4256
rect 4149 4239 4153 4256
rect 4195 4239 4218 4256
rect 4218 4239 4229 4256
rect 4271 4239 4287 4256
rect 4287 4239 4305 4256
rect 4347 4239 4356 4256
rect 4356 4239 4381 4256
rect 4423 4239 4425 4256
rect 4425 4239 4457 4256
rect 4499 4239 4533 4273
rect 3891 4188 3925 4197
rect 3967 4188 4001 4197
rect 4043 4188 4077 4197
rect 4119 4188 4153 4197
rect 4195 4188 4229 4197
rect 4271 4188 4305 4197
rect 4347 4188 4381 4197
rect 4423 4188 4457 4197
rect 3891 4163 3908 4188
rect 3908 4163 3925 4188
rect 3967 4163 3977 4188
rect 3977 4163 4001 4188
rect 4043 4163 4046 4188
rect 4046 4163 4077 4188
rect 4119 4163 4149 4188
rect 4149 4163 4153 4188
rect 4195 4163 4218 4188
rect 4218 4163 4229 4188
rect 4271 4163 4287 4188
rect 4287 4163 4305 4188
rect 4347 4163 4356 4188
rect 4356 4163 4381 4188
rect 4423 4163 4425 4188
rect 4425 4163 4457 4188
rect 4499 4163 4533 4197
rect 3891 4120 3925 4121
rect 3967 4120 4001 4121
rect 4043 4120 4077 4121
rect 4119 4120 4153 4121
rect 4195 4120 4229 4121
rect 4271 4120 4305 4121
rect 4347 4120 4381 4121
rect 4423 4120 4457 4121
rect -4 3997 30 4031
rect 68 3997 102 4031
rect 3891 4087 3908 4120
rect 3908 4087 3925 4120
rect 3967 4087 3977 4120
rect 3977 4087 4001 4120
rect 4043 4087 4046 4120
rect 4046 4087 4077 4120
rect 4119 4087 4149 4120
rect 4149 4087 4153 4120
rect 4195 4087 4218 4120
rect 4218 4087 4229 4120
rect 4271 4087 4287 4120
rect 4287 4087 4305 4120
rect 4347 4087 4356 4120
rect 4356 4087 4381 4120
rect 4423 4087 4425 4120
rect 4425 4087 4457 4120
rect 4499 4087 4533 4121
rect 3891 4018 3908 4045
rect 3908 4018 3925 4045
rect 3967 4018 3977 4045
rect 3977 4018 4001 4045
rect 4043 4018 4046 4045
rect 4046 4018 4077 4045
rect 4119 4018 4149 4045
rect 4149 4018 4153 4045
rect 4195 4018 4218 4045
rect 4218 4018 4229 4045
rect 4271 4018 4287 4045
rect 4287 4018 4305 4045
rect 4347 4018 4356 4045
rect 4356 4018 4381 4045
rect 4423 4018 4425 4045
rect 4425 4018 4457 4045
rect 3891 4011 3925 4018
rect 3967 4011 4001 4018
rect 4043 4011 4077 4018
rect 4119 4011 4153 4018
rect 4195 4011 4229 4018
rect 4271 4011 4305 4018
rect 4347 4011 4381 4018
rect 4423 4011 4457 4018
rect 4499 4011 4533 4045
rect 3891 3950 3908 3968
rect 3908 3950 3925 3968
rect 3967 3950 3977 3968
rect 3977 3950 4001 3968
rect 4043 3950 4046 3968
rect 4046 3950 4077 3968
rect 4119 3950 4149 3968
rect 4149 3950 4153 3968
rect 4195 3950 4218 3968
rect 4218 3950 4229 3968
rect 4271 3950 4287 3968
rect 4287 3950 4305 3968
rect 4347 3950 4356 3968
rect 4356 3950 4381 3968
rect 4423 3950 4425 3968
rect 4425 3950 4457 3968
rect 3891 3934 3925 3950
rect 3967 3934 4001 3950
rect 4043 3934 4077 3950
rect 4119 3934 4153 3950
rect 4195 3934 4229 3950
rect 4271 3934 4305 3950
rect 4347 3934 4381 3950
rect 4423 3934 4457 3950
rect 4499 3934 4533 3968
rect 3891 3882 3908 3891
rect 3908 3882 3925 3891
rect 3967 3882 3977 3891
rect 3977 3882 4001 3891
rect 4043 3882 4046 3891
rect 4046 3882 4077 3891
rect 4119 3882 4149 3891
rect 4149 3882 4153 3891
rect 4195 3882 4218 3891
rect 4218 3882 4229 3891
rect 4271 3882 4287 3891
rect 4287 3882 4305 3891
rect 4347 3882 4356 3891
rect 4356 3882 4381 3891
rect 4423 3882 4425 3891
rect 4425 3882 4457 3891
rect 3891 3857 3925 3882
rect 3967 3857 4001 3882
rect 4043 3857 4077 3882
rect 4119 3857 4153 3882
rect 4195 3857 4229 3882
rect 4271 3857 4305 3882
rect 4347 3857 4381 3882
rect 4423 3857 4457 3882
rect 4499 3857 4533 3891
rect 11937 4290 11949 4322
rect 11949 4290 11971 4322
rect 12010 4290 12018 4322
rect 12018 4290 12044 4322
rect 12083 4290 12087 4322
rect 12087 4290 12117 4322
rect 12156 4290 12190 4322
rect 12229 4290 12259 4322
rect 12259 4290 12263 4322
rect 12302 4290 12328 4322
rect 12328 4290 12336 4322
rect 12375 4290 12397 4322
rect 12397 4290 12409 4322
rect 12448 4290 12466 4322
rect 12466 4290 12482 4322
rect 12521 4290 12535 4322
rect 12535 4290 12555 4322
rect 12594 4290 12604 4322
rect 12604 4290 12628 4322
rect 12667 4290 12673 4322
rect 12673 4290 12701 4322
rect 12740 4290 12742 4322
rect 12742 4290 12774 4322
rect 12813 4290 12846 4322
rect 12846 4290 12847 4322
rect 12886 4290 12915 4322
rect 12915 4290 12920 4322
rect 12959 4290 12984 4322
rect 12984 4290 12993 4322
rect 13032 4290 13053 4322
rect 13053 4290 13066 4322
rect 13105 4290 13122 4322
rect 13122 4290 13139 4322
rect 13178 4290 13191 4322
rect 13191 4290 13212 4322
rect 13251 4290 13260 4322
rect 13260 4290 13285 4322
rect 13324 4290 13329 4322
rect 13329 4290 13358 4322
rect 13397 4290 13398 4322
rect 13398 4290 13431 4322
rect 13470 4290 13501 4322
rect 13501 4290 13504 4322
rect 13543 4290 13570 4322
rect 13570 4290 13577 4322
rect 13616 4290 13639 4322
rect 13639 4290 13650 4322
rect 13689 4290 13708 4322
rect 13708 4290 13723 4322
rect 13762 4290 13777 4322
rect 13777 4290 13796 4322
rect 13835 4290 13846 4322
rect 13846 4290 13869 4322
rect 13908 4290 13915 4322
rect 13915 4290 13942 4322
rect 13981 4290 13984 4322
rect 13984 4290 14015 4322
rect 11937 4288 11971 4290
rect 12010 4288 12044 4290
rect 12083 4288 12117 4290
rect 12156 4288 12190 4290
rect 12229 4288 12263 4290
rect 12302 4288 12336 4290
rect 12375 4288 12409 4290
rect 12448 4288 12482 4290
rect 12521 4288 12555 4290
rect 12594 4288 12628 4290
rect 12667 4288 12701 4290
rect 12740 4288 12774 4290
rect 12813 4288 12847 4290
rect 12886 4288 12920 4290
rect 12959 4288 12993 4290
rect 13032 4288 13066 4290
rect 13105 4288 13139 4290
rect 13178 4288 13212 4290
rect 13251 4288 13285 4290
rect 13324 4288 13358 4290
rect 13397 4288 13431 4290
rect 13470 4288 13504 4290
rect 13543 4288 13577 4290
rect 13616 4288 13650 4290
rect 13689 4288 13723 4290
rect 13762 4288 13796 4290
rect 13835 4288 13869 4290
rect 13908 4288 13942 4290
rect 13981 4288 14015 4290
rect 14054 4288 14088 4322
rect 14127 4290 14157 4322
rect 14157 4290 14161 4322
rect 14200 4290 14226 4322
rect 14226 4290 14234 4322
rect 14273 4290 14295 4322
rect 14295 4290 14307 4322
rect 14346 4290 14364 4322
rect 14364 4290 14380 4322
rect 14419 4290 14433 4322
rect 14433 4290 14453 4322
rect 14492 4290 14502 4322
rect 14502 4290 14526 4322
rect 14565 4290 14571 4322
rect 14571 4290 14599 4322
rect 14638 4290 14640 4322
rect 14640 4290 14672 4322
rect 14711 4290 14743 4322
rect 14743 4290 14745 4322
rect 14784 4290 14812 4322
rect 14812 4290 14818 4322
rect 14857 4290 14881 4322
rect 14881 4290 14891 4322
rect 14930 4290 14950 4322
rect 14950 4290 14964 4322
rect 15003 4290 15019 4322
rect 15019 4290 15037 4322
rect 15076 4290 15088 4322
rect 15088 4290 15110 4322
rect 15149 4290 15157 4322
rect 15157 4290 15183 4322
rect 15222 4290 15226 4322
rect 15226 4290 15256 4322
rect 14127 4288 14161 4290
rect 14200 4288 14234 4290
rect 14273 4288 14307 4290
rect 14346 4288 14380 4290
rect 14419 4288 14453 4290
rect 14492 4288 14526 4290
rect 14565 4288 14599 4290
rect 14638 4288 14672 4290
rect 14711 4288 14745 4290
rect 14784 4288 14818 4290
rect 14857 4288 14891 4290
rect 14930 4288 14964 4290
rect 15003 4288 15037 4290
rect 15076 4288 15110 4290
rect 15149 4288 15183 4290
rect 15222 4288 15256 4290
rect 15295 4288 15329 4322
rect 15368 4290 15399 4322
rect 15399 4290 15402 4322
rect 15441 4290 15468 4322
rect 15468 4290 15475 4322
rect 15514 4290 15537 4322
rect 15537 4290 15548 4322
rect 15587 4290 15606 4322
rect 15606 4290 15621 4322
rect 15660 4290 15675 4322
rect 15675 4290 15694 4322
rect 15733 4290 15744 4322
rect 15744 4290 15767 4322
rect 15806 4290 15813 4322
rect 15813 4290 15840 4322
rect 15879 4290 15882 4322
rect 15882 4290 15913 4322
rect 15952 4290 15985 4322
rect 15985 4290 15986 4322
rect 16025 4290 16054 4322
rect 16054 4290 16059 4322
rect 16098 4290 16123 4322
rect 16123 4290 16132 4322
rect 16171 4290 16192 4322
rect 16192 4290 16205 4322
rect 16244 4290 16261 4322
rect 16261 4290 16278 4322
rect 16317 4290 16330 4322
rect 16330 4290 16351 4322
rect 15368 4288 15402 4290
rect 15441 4288 15475 4290
rect 15514 4288 15548 4290
rect 15587 4288 15621 4290
rect 15660 4288 15694 4290
rect 15733 4288 15767 4290
rect 15806 4288 15840 4290
rect 15879 4288 15913 4290
rect 15952 4288 15986 4290
rect 16025 4288 16059 4290
rect 16098 4288 16132 4290
rect 16171 4288 16205 4290
rect 16244 4288 16278 4290
rect 16317 4288 16351 4290
rect 11937 4222 11949 4250
rect 11949 4222 11971 4250
rect 12010 4222 12018 4250
rect 12018 4222 12044 4250
rect 12083 4222 12087 4250
rect 12087 4222 12117 4250
rect 12156 4222 12190 4250
rect 12229 4222 12259 4250
rect 12259 4222 12263 4250
rect 12302 4222 12328 4250
rect 12328 4222 12336 4250
rect 12375 4222 12397 4250
rect 12397 4222 12409 4250
rect 12448 4222 12466 4250
rect 12466 4222 12482 4250
rect 12521 4222 12535 4250
rect 12535 4222 12555 4250
rect 12594 4222 12604 4250
rect 12604 4222 12628 4250
rect 12667 4222 12673 4250
rect 12673 4222 12701 4250
rect 12740 4222 12742 4250
rect 12742 4222 12774 4250
rect 12813 4222 12846 4250
rect 12846 4222 12847 4250
rect 12886 4222 12915 4250
rect 12915 4222 12920 4250
rect 12959 4222 12984 4250
rect 12984 4222 12993 4250
rect 13032 4222 13053 4250
rect 13053 4222 13066 4250
rect 13105 4222 13122 4250
rect 13122 4222 13139 4250
rect 13178 4222 13191 4250
rect 13191 4222 13212 4250
rect 13251 4222 13260 4250
rect 13260 4222 13285 4250
rect 13324 4222 13329 4250
rect 13329 4222 13358 4250
rect 13397 4222 13398 4250
rect 13398 4222 13431 4250
rect 13470 4222 13501 4250
rect 13501 4222 13504 4250
rect 13543 4222 13570 4250
rect 13570 4222 13577 4250
rect 13616 4222 13639 4250
rect 13639 4222 13650 4250
rect 13689 4222 13708 4250
rect 13708 4222 13723 4250
rect 13762 4222 13777 4250
rect 13777 4222 13796 4250
rect 13835 4222 13846 4250
rect 13846 4222 13869 4250
rect 13908 4222 13915 4250
rect 13915 4222 13942 4250
rect 13981 4222 13984 4250
rect 13984 4222 14015 4250
rect 11937 4216 11971 4222
rect 12010 4216 12044 4222
rect 12083 4216 12117 4222
rect 12156 4216 12190 4222
rect 12229 4216 12263 4222
rect 12302 4216 12336 4222
rect 12375 4216 12409 4222
rect 12448 4216 12482 4222
rect 12521 4216 12555 4222
rect 12594 4216 12628 4222
rect 12667 4216 12701 4222
rect 12740 4216 12774 4222
rect 12813 4216 12847 4222
rect 12886 4216 12920 4222
rect 12959 4216 12993 4222
rect 13032 4216 13066 4222
rect 13105 4216 13139 4222
rect 13178 4216 13212 4222
rect 13251 4216 13285 4222
rect 13324 4216 13358 4222
rect 13397 4216 13431 4222
rect 13470 4216 13504 4222
rect 13543 4216 13577 4222
rect 13616 4216 13650 4222
rect 13689 4216 13723 4222
rect 13762 4216 13796 4222
rect 13835 4216 13869 4222
rect 13908 4216 13942 4222
rect 13981 4216 14015 4222
rect 14054 4216 14088 4250
rect 14127 4222 14157 4250
rect 14157 4222 14161 4250
rect 14200 4222 14226 4250
rect 14226 4222 14234 4250
rect 14273 4222 14295 4250
rect 14295 4222 14307 4250
rect 14346 4222 14364 4250
rect 14364 4222 14380 4250
rect 14419 4222 14433 4250
rect 14433 4222 14453 4250
rect 14492 4222 14502 4250
rect 14502 4222 14526 4250
rect 14565 4222 14571 4250
rect 14571 4222 14599 4250
rect 14638 4222 14640 4250
rect 14640 4222 14672 4250
rect 14711 4222 14743 4250
rect 14743 4222 14745 4250
rect 14784 4222 14812 4250
rect 14812 4222 14818 4250
rect 14857 4222 14881 4250
rect 14881 4222 14891 4250
rect 14930 4222 14950 4250
rect 14950 4222 14964 4250
rect 15003 4222 15019 4250
rect 15019 4222 15037 4250
rect 15076 4222 15088 4250
rect 15088 4222 15110 4250
rect 15149 4222 15157 4250
rect 15157 4222 15183 4250
rect 15222 4222 15226 4250
rect 15226 4222 15256 4250
rect 14127 4216 14161 4222
rect 14200 4216 14234 4222
rect 14273 4216 14307 4222
rect 14346 4216 14380 4222
rect 14419 4216 14453 4222
rect 14492 4216 14526 4222
rect 14565 4216 14599 4222
rect 14638 4216 14672 4222
rect 14711 4216 14745 4222
rect 14784 4216 14818 4222
rect 14857 4216 14891 4222
rect 14930 4216 14964 4222
rect 15003 4216 15037 4222
rect 15076 4216 15110 4222
rect 15149 4216 15183 4222
rect 15222 4216 15256 4222
rect 15295 4216 15329 4250
rect 15368 4222 15399 4250
rect 15399 4222 15402 4250
rect 15441 4222 15468 4250
rect 15468 4222 15475 4250
rect 15514 4222 15537 4250
rect 15537 4222 15548 4250
rect 15587 4222 15606 4250
rect 15606 4222 15621 4250
rect 15660 4222 15675 4250
rect 15675 4222 15694 4250
rect 15733 4222 15744 4250
rect 15744 4222 15767 4250
rect 15806 4222 15813 4250
rect 15813 4222 15840 4250
rect 15879 4222 15882 4250
rect 15882 4222 15913 4250
rect 15952 4222 15985 4250
rect 15985 4222 15986 4250
rect 16025 4222 16054 4250
rect 16054 4222 16059 4250
rect 16098 4222 16123 4250
rect 16123 4222 16132 4250
rect 16171 4222 16192 4250
rect 16192 4222 16205 4250
rect 16244 4222 16261 4250
rect 16261 4222 16278 4250
rect 16317 4222 16330 4250
rect 16330 4222 16351 4250
rect 15368 4216 15402 4222
rect 15441 4216 15475 4222
rect 15514 4216 15548 4222
rect 15587 4216 15621 4222
rect 15660 4216 15694 4222
rect 15733 4216 15767 4222
rect 15806 4216 15840 4222
rect 15879 4216 15913 4222
rect 15952 4216 15986 4222
rect 16025 4216 16059 4222
rect 16098 4216 16132 4222
rect 16171 4216 16205 4222
rect 16244 4216 16278 4222
rect 16317 4216 16351 4222
rect 11937 4154 11949 4178
rect 11949 4154 11971 4178
rect 12010 4154 12018 4178
rect 12018 4154 12044 4178
rect 12083 4154 12087 4178
rect 12087 4154 12117 4178
rect 12156 4154 12190 4178
rect 12229 4154 12259 4178
rect 12259 4154 12263 4178
rect 12302 4154 12328 4178
rect 12328 4154 12336 4178
rect 12375 4154 12397 4178
rect 12397 4154 12409 4178
rect 12448 4154 12466 4178
rect 12466 4154 12482 4178
rect 12521 4154 12535 4178
rect 12535 4154 12555 4178
rect 12594 4154 12604 4178
rect 12604 4154 12628 4178
rect 12667 4154 12673 4178
rect 12673 4154 12701 4178
rect 12740 4154 12742 4178
rect 12742 4154 12774 4178
rect 12813 4154 12846 4178
rect 12846 4154 12847 4178
rect 12886 4154 12915 4178
rect 12915 4154 12920 4178
rect 12959 4154 12984 4178
rect 12984 4154 12993 4178
rect 13032 4154 13053 4178
rect 13053 4154 13066 4178
rect 13105 4154 13122 4178
rect 13122 4154 13139 4178
rect 13178 4154 13191 4178
rect 13191 4154 13212 4178
rect 13251 4154 13260 4178
rect 13260 4154 13285 4178
rect 13324 4154 13329 4178
rect 13329 4154 13358 4178
rect 13397 4154 13398 4178
rect 13398 4154 13431 4178
rect 13470 4154 13501 4178
rect 13501 4154 13504 4178
rect 13543 4154 13570 4178
rect 13570 4154 13577 4178
rect 13616 4154 13639 4178
rect 13639 4154 13650 4178
rect 13689 4154 13708 4178
rect 13708 4154 13723 4178
rect 13762 4154 13777 4178
rect 13777 4154 13796 4178
rect 13835 4154 13846 4178
rect 13846 4154 13869 4178
rect 13908 4154 13915 4178
rect 13915 4154 13942 4178
rect 13981 4154 13984 4178
rect 13984 4154 14015 4178
rect 11937 4144 11971 4154
rect 12010 4144 12044 4154
rect 12083 4144 12117 4154
rect 12156 4144 12190 4154
rect 12229 4144 12263 4154
rect 12302 4144 12336 4154
rect 12375 4144 12409 4154
rect 12448 4144 12482 4154
rect 12521 4144 12555 4154
rect 12594 4144 12628 4154
rect 12667 4144 12701 4154
rect 12740 4144 12774 4154
rect 12813 4144 12847 4154
rect 12886 4144 12920 4154
rect 12959 4144 12993 4154
rect 13032 4144 13066 4154
rect 13105 4144 13139 4154
rect 13178 4144 13212 4154
rect 13251 4144 13285 4154
rect 13324 4144 13358 4154
rect 13397 4144 13431 4154
rect 13470 4144 13504 4154
rect 13543 4144 13577 4154
rect 13616 4144 13650 4154
rect 13689 4144 13723 4154
rect 13762 4144 13796 4154
rect 13835 4144 13869 4154
rect 13908 4144 13942 4154
rect 13981 4144 14015 4154
rect 14054 4144 14088 4178
rect 14127 4154 14157 4178
rect 14157 4154 14161 4178
rect 14200 4154 14226 4178
rect 14226 4154 14234 4178
rect 14273 4154 14295 4178
rect 14295 4154 14307 4178
rect 14346 4154 14364 4178
rect 14364 4154 14380 4178
rect 14419 4154 14433 4178
rect 14433 4154 14453 4178
rect 14492 4154 14502 4178
rect 14502 4154 14526 4178
rect 14565 4154 14571 4178
rect 14571 4154 14599 4178
rect 14638 4154 14640 4178
rect 14640 4154 14672 4178
rect 14711 4154 14743 4178
rect 14743 4154 14745 4178
rect 14784 4154 14812 4178
rect 14812 4154 14818 4178
rect 14857 4154 14881 4178
rect 14881 4154 14891 4178
rect 14930 4154 14950 4178
rect 14950 4154 14964 4178
rect 15003 4154 15019 4178
rect 15019 4154 15037 4178
rect 15076 4154 15088 4178
rect 15088 4154 15110 4178
rect 15149 4154 15157 4178
rect 15157 4154 15183 4178
rect 15222 4154 15226 4178
rect 15226 4154 15256 4178
rect 14127 4144 14161 4154
rect 14200 4144 14234 4154
rect 14273 4144 14307 4154
rect 14346 4144 14380 4154
rect 14419 4144 14453 4154
rect 14492 4144 14526 4154
rect 14565 4144 14599 4154
rect 14638 4144 14672 4154
rect 14711 4144 14745 4154
rect 14784 4144 14818 4154
rect 14857 4144 14891 4154
rect 14930 4144 14964 4154
rect 15003 4144 15037 4154
rect 15076 4144 15110 4154
rect 15149 4144 15183 4154
rect 15222 4144 15256 4154
rect 15295 4144 15329 4178
rect 15368 4154 15399 4178
rect 15399 4154 15402 4178
rect 15441 4154 15468 4178
rect 15468 4154 15475 4178
rect 15514 4154 15537 4178
rect 15537 4154 15548 4178
rect 15587 4154 15606 4178
rect 15606 4154 15621 4178
rect 15660 4154 15675 4178
rect 15675 4154 15694 4178
rect 15733 4154 15744 4178
rect 15744 4154 15767 4178
rect 15806 4154 15813 4178
rect 15813 4154 15840 4178
rect 15879 4154 15882 4178
rect 15882 4154 15913 4178
rect 15952 4154 15985 4178
rect 15985 4154 15986 4178
rect 16025 4154 16054 4178
rect 16054 4154 16059 4178
rect 16098 4154 16123 4178
rect 16123 4154 16132 4178
rect 16171 4154 16192 4178
rect 16192 4154 16205 4178
rect 16244 4154 16261 4178
rect 16261 4154 16278 4178
rect 16317 4154 16330 4178
rect 16330 4154 16351 4178
rect 15368 4144 15402 4154
rect 15441 4144 15475 4154
rect 15514 4144 15548 4154
rect 15587 4144 15621 4154
rect 15660 4144 15694 4154
rect 15733 4144 15767 4154
rect 15806 4144 15840 4154
rect 15879 4144 15913 4154
rect 15952 4144 15986 4154
rect 16025 4144 16059 4154
rect 16098 4144 16132 4154
rect 16171 4144 16205 4154
rect 16244 4144 16278 4154
rect 16317 4144 16351 4154
rect 11937 4086 11949 4106
rect 11949 4086 11971 4106
rect 12010 4086 12018 4106
rect 12018 4086 12044 4106
rect 12083 4086 12087 4106
rect 12087 4086 12117 4106
rect 12156 4086 12190 4106
rect 12229 4086 12259 4106
rect 12259 4086 12263 4106
rect 12302 4086 12328 4106
rect 12328 4086 12336 4106
rect 12375 4086 12397 4106
rect 12397 4086 12409 4106
rect 12448 4086 12466 4106
rect 12466 4086 12482 4106
rect 12521 4086 12535 4106
rect 12535 4086 12555 4106
rect 12594 4086 12604 4106
rect 12604 4086 12628 4106
rect 12667 4086 12673 4106
rect 12673 4086 12701 4106
rect 12740 4086 12742 4106
rect 12742 4086 12774 4106
rect 12813 4086 12846 4106
rect 12846 4086 12847 4106
rect 12886 4086 12915 4106
rect 12915 4086 12920 4106
rect 12959 4086 12984 4106
rect 12984 4086 12993 4106
rect 13032 4086 13053 4106
rect 13053 4086 13066 4106
rect 13105 4086 13122 4106
rect 13122 4086 13139 4106
rect 13178 4086 13191 4106
rect 13191 4086 13212 4106
rect 13251 4086 13260 4106
rect 13260 4086 13285 4106
rect 13324 4086 13329 4106
rect 13329 4086 13358 4106
rect 13397 4086 13398 4106
rect 13398 4086 13431 4106
rect 13470 4086 13501 4106
rect 13501 4086 13504 4106
rect 13543 4086 13570 4106
rect 13570 4086 13577 4106
rect 13616 4086 13639 4106
rect 13639 4086 13650 4106
rect 13689 4086 13708 4106
rect 13708 4086 13723 4106
rect 13762 4086 13777 4106
rect 13777 4086 13796 4106
rect 13835 4086 13846 4106
rect 13846 4086 13869 4106
rect 13908 4086 13915 4106
rect 13915 4086 13942 4106
rect 13981 4086 13984 4106
rect 13984 4086 14015 4106
rect 11937 4072 11971 4086
rect 12010 4072 12044 4086
rect 12083 4072 12117 4086
rect 12156 4072 12190 4086
rect 12229 4072 12263 4086
rect 12302 4072 12336 4086
rect 12375 4072 12409 4086
rect 12448 4072 12482 4086
rect 12521 4072 12555 4086
rect 12594 4072 12628 4086
rect 12667 4072 12701 4086
rect 12740 4072 12774 4086
rect 12813 4072 12847 4086
rect 12886 4072 12920 4086
rect 12959 4072 12993 4086
rect 13032 4072 13066 4086
rect 13105 4072 13139 4086
rect 13178 4072 13212 4086
rect 13251 4072 13285 4086
rect 13324 4072 13358 4086
rect 13397 4072 13431 4086
rect 13470 4072 13504 4086
rect 13543 4072 13577 4086
rect 13616 4072 13650 4086
rect 13689 4072 13723 4086
rect 13762 4072 13796 4086
rect 13835 4072 13869 4086
rect 13908 4072 13942 4086
rect 13981 4072 14015 4086
rect 14054 4072 14088 4106
rect 14127 4086 14157 4106
rect 14157 4086 14161 4106
rect 14200 4086 14226 4106
rect 14226 4086 14234 4106
rect 14273 4086 14295 4106
rect 14295 4086 14307 4106
rect 14346 4086 14364 4106
rect 14364 4086 14380 4106
rect 14419 4086 14433 4106
rect 14433 4086 14453 4106
rect 14492 4086 14502 4106
rect 14502 4086 14526 4106
rect 14565 4086 14571 4106
rect 14571 4086 14599 4106
rect 14638 4086 14640 4106
rect 14640 4086 14672 4106
rect 14711 4086 14743 4106
rect 14743 4086 14745 4106
rect 14784 4086 14812 4106
rect 14812 4086 14818 4106
rect 14857 4086 14881 4106
rect 14881 4086 14891 4106
rect 14930 4086 14950 4106
rect 14950 4086 14964 4106
rect 15003 4086 15019 4106
rect 15019 4086 15037 4106
rect 15076 4086 15088 4106
rect 15088 4086 15110 4106
rect 15149 4086 15157 4106
rect 15157 4086 15183 4106
rect 15222 4086 15226 4106
rect 15226 4086 15256 4106
rect 14127 4072 14161 4086
rect 14200 4072 14234 4086
rect 14273 4072 14307 4086
rect 14346 4072 14380 4086
rect 14419 4072 14453 4086
rect 14492 4072 14526 4086
rect 14565 4072 14599 4086
rect 14638 4072 14672 4086
rect 14711 4072 14745 4086
rect 14784 4072 14818 4086
rect 14857 4072 14891 4086
rect 14930 4072 14964 4086
rect 15003 4072 15037 4086
rect 15076 4072 15110 4086
rect 15149 4072 15183 4086
rect 15222 4072 15256 4086
rect 15295 4072 15329 4106
rect 15368 4086 15399 4106
rect 15399 4086 15402 4106
rect 15441 4086 15468 4106
rect 15468 4086 15475 4106
rect 15514 4086 15537 4106
rect 15537 4086 15548 4106
rect 15587 4086 15606 4106
rect 15606 4086 15621 4106
rect 15660 4086 15675 4106
rect 15675 4086 15694 4106
rect 15733 4086 15744 4106
rect 15744 4086 15767 4106
rect 15806 4086 15813 4106
rect 15813 4086 15840 4106
rect 15879 4086 15882 4106
rect 15882 4086 15913 4106
rect 15952 4086 15985 4106
rect 15985 4086 15986 4106
rect 16025 4086 16054 4106
rect 16054 4086 16059 4106
rect 16098 4086 16123 4106
rect 16123 4086 16132 4106
rect 16171 4086 16192 4106
rect 16192 4086 16205 4106
rect 16244 4086 16261 4106
rect 16261 4086 16278 4106
rect 16317 4086 16330 4106
rect 16330 4086 16351 4106
rect 15368 4072 15402 4086
rect 15441 4072 15475 4086
rect 15514 4072 15548 4086
rect 15587 4072 15621 4086
rect 15660 4072 15694 4086
rect 15733 4072 15767 4086
rect 15806 4072 15840 4086
rect 15879 4072 15913 4086
rect 15952 4072 15986 4086
rect 16025 4072 16059 4086
rect 16098 4072 16132 4086
rect 16171 4072 16205 4086
rect 16244 4072 16278 4086
rect 16317 4072 16351 4086
rect 11937 4018 11949 4034
rect 11949 4018 11971 4034
rect 12010 4018 12018 4034
rect 12018 4018 12044 4034
rect 12083 4018 12087 4034
rect 12087 4018 12117 4034
rect 12156 4018 12190 4034
rect 12229 4018 12259 4034
rect 12259 4018 12263 4034
rect 12302 4018 12328 4034
rect 12328 4018 12336 4034
rect 12375 4018 12397 4034
rect 12397 4018 12409 4034
rect 12448 4018 12466 4034
rect 12466 4018 12482 4034
rect 12521 4018 12535 4034
rect 12535 4018 12555 4034
rect 12594 4018 12604 4034
rect 12604 4018 12628 4034
rect 12667 4018 12673 4034
rect 12673 4018 12701 4034
rect 12740 4018 12742 4034
rect 12742 4018 12774 4034
rect 12813 4018 12846 4034
rect 12846 4018 12847 4034
rect 12886 4018 12915 4034
rect 12915 4018 12920 4034
rect 12959 4018 12984 4034
rect 12984 4018 12993 4034
rect 13032 4018 13053 4034
rect 13053 4018 13066 4034
rect 13105 4018 13122 4034
rect 13122 4018 13139 4034
rect 13178 4018 13191 4034
rect 13191 4018 13212 4034
rect 13251 4018 13260 4034
rect 13260 4018 13285 4034
rect 13324 4018 13329 4034
rect 13329 4018 13358 4034
rect 13397 4018 13398 4034
rect 13398 4018 13431 4034
rect 13470 4018 13501 4034
rect 13501 4018 13504 4034
rect 13543 4018 13570 4034
rect 13570 4018 13577 4034
rect 13616 4018 13639 4034
rect 13639 4018 13650 4034
rect 13689 4018 13708 4034
rect 13708 4018 13723 4034
rect 13762 4018 13777 4034
rect 13777 4018 13796 4034
rect 13835 4018 13846 4034
rect 13846 4018 13869 4034
rect 13908 4018 13915 4034
rect 13915 4018 13942 4034
rect 13981 4018 13984 4034
rect 13984 4018 14015 4034
rect 11937 4000 11971 4018
rect 12010 4000 12044 4018
rect 12083 4000 12117 4018
rect 12156 4000 12190 4018
rect 12229 4000 12263 4018
rect 12302 4000 12336 4018
rect 12375 4000 12409 4018
rect 12448 4000 12482 4018
rect 12521 4000 12555 4018
rect 12594 4000 12628 4018
rect 12667 4000 12701 4018
rect 12740 4000 12774 4018
rect 12813 4000 12847 4018
rect 12886 4000 12920 4018
rect 12959 4000 12993 4018
rect 13032 4000 13066 4018
rect 13105 4000 13139 4018
rect 13178 4000 13212 4018
rect 13251 4000 13285 4018
rect 13324 4000 13358 4018
rect 13397 4000 13431 4018
rect 13470 4000 13504 4018
rect 13543 4000 13577 4018
rect 13616 4000 13650 4018
rect 13689 4000 13723 4018
rect 13762 4000 13796 4018
rect 13835 4000 13869 4018
rect 13908 4000 13942 4018
rect 13981 4000 14015 4018
rect 14054 4000 14088 4034
rect 14127 4018 14157 4034
rect 14157 4018 14161 4034
rect 14200 4018 14226 4034
rect 14226 4018 14234 4034
rect 14273 4018 14295 4034
rect 14295 4018 14307 4034
rect 14346 4018 14364 4034
rect 14364 4018 14380 4034
rect 14419 4018 14433 4034
rect 14433 4018 14453 4034
rect 14492 4018 14502 4034
rect 14502 4018 14526 4034
rect 14565 4018 14571 4034
rect 14571 4018 14599 4034
rect 14638 4018 14640 4034
rect 14640 4018 14672 4034
rect 14711 4018 14743 4034
rect 14743 4018 14745 4034
rect 14784 4018 14812 4034
rect 14812 4018 14818 4034
rect 14857 4018 14881 4034
rect 14881 4018 14891 4034
rect 14930 4018 14950 4034
rect 14950 4018 14964 4034
rect 15003 4018 15019 4034
rect 15019 4018 15037 4034
rect 15076 4018 15088 4034
rect 15088 4018 15110 4034
rect 15149 4018 15157 4034
rect 15157 4018 15183 4034
rect 15222 4018 15226 4034
rect 15226 4018 15256 4034
rect 14127 4000 14161 4018
rect 14200 4000 14234 4018
rect 14273 4000 14307 4018
rect 14346 4000 14380 4018
rect 14419 4000 14453 4018
rect 14492 4000 14526 4018
rect 14565 4000 14599 4018
rect 14638 4000 14672 4018
rect 14711 4000 14745 4018
rect 14784 4000 14818 4018
rect 14857 4000 14891 4018
rect 14930 4000 14964 4018
rect 15003 4000 15037 4018
rect 15076 4000 15110 4018
rect 15149 4000 15183 4018
rect 15222 4000 15256 4018
rect 15295 4000 15329 4034
rect 15368 4018 15399 4034
rect 15399 4018 15402 4034
rect 15441 4018 15468 4034
rect 15468 4018 15475 4034
rect 15514 4018 15537 4034
rect 15537 4018 15548 4034
rect 15587 4018 15606 4034
rect 15606 4018 15621 4034
rect 15660 4018 15675 4034
rect 15675 4018 15694 4034
rect 15733 4018 15744 4034
rect 15744 4018 15767 4034
rect 15806 4018 15813 4034
rect 15813 4018 15840 4034
rect 15879 4018 15882 4034
rect 15882 4018 15913 4034
rect 15952 4018 15985 4034
rect 15985 4018 15986 4034
rect 16025 4018 16054 4034
rect 16054 4018 16059 4034
rect 16098 4018 16123 4034
rect 16123 4018 16132 4034
rect 16171 4018 16192 4034
rect 16192 4018 16205 4034
rect 16244 4018 16261 4034
rect 16261 4018 16278 4034
rect 16317 4018 16330 4034
rect 16330 4018 16351 4034
rect 15368 4000 15402 4018
rect 15441 4000 15475 4018
rect 15514 4000 15548 4018
rect 15587 4000 15621 4018
rect 15660 4000 15694 4018
rect 15733 4000 15767 4018
rect 15806 4000 15840 4018
rect 15879 4000 15913 4018
rect 15952 4000 15986 4018
rect 16025 4000 16059 4018
rect 16098 4000 16132 4018
rect 16171 4000 16205 4018
rect 16244 4000 16278 4018
rect 16317 4000 16351 4018
rect 11937 3950 11949 3962
rect 11949 3950 11971 3962
rect 12010 3950 12018 3962
rect 12018 3950 12044 3962
rect 12083 3950 12087 3962
rect 12087 3950 12117 3962
rect 12156 3950 12190 3962
rect 12229 3950 12259 3962
rect 12259 3950 12263 3962
rect 12302 3950 12328 3962
rect 12328 3950 12336 3962
rect 12375 3950 12397 3962
rect 12397 3950 12409 3962
rect 12448 3950 12466 3962
rect 12466 3950 12482 3962
rect 12521 3950 12535 3962
rect 12535 3950 12555 3962
rect 12594 3950 12604 3962
rect 12604 3950 12628 3962
rect 12667 3950 12673 3962
rect 12673 3950 12701 3962
rect 12740 3950 12742 3962
rect 12742 3950 12774 3962
rect 12813 3950 12846 3962
rect 12846 3950 12847 3962
rect 12886 3950 12915 3962
rect 12915 3950 12920 3962
rect 12959 3950 12984 3962
rect 12984 3950 12993 3962
rect 13032 3950 13053 3962
rect 13053 3950 13066 3962
rect 13105 3950 13122 3962
rect 13122 3950 13139 3962
rect 13178 3950 13191 3962
rect 13191 3950 13212 3962
rect 13251 3950 13260 3962
rect 13260 3950 13285 3962
rect 13324 3950 13329 3962
rect 13329 3950 13358 3962
rect 13397 3950 13398 3962
rect 13398 3950 13431 3962
rect 13470 3950 13501 3962
rect 13501 3950 13504 3962
rect 13543 3950 13570 3962
rect 13570 3950 13577 3962
rect 13616 3950 13639 3962
rect 13639 3950 13650 3962
rect 13689 3950 13708 3962
rect 13708 3950 13723 3962
rect 13762 3950 13777 3962
rect 13777 3950 13796 3962
rect 13835 3950 13846 3962
rect 13846 3950 13869 3962
rect 13908 3950 13915 3962
rect 13915 3950 13942 3962
rect 13981 3950 13984 3962
rect 13984 3950 14015 3962
rect 11937 3928 11971 3950
rect 12010 3928 12044 3950
rect 12083 3928 12117 3950
rect 12156 3928 12190 3950
rect 12229 3928 12263 3950
rect 12302 3928 12336 3950
rect 12375 3928 12409 3950
rect 12448 3928 12482 3950
rect 12521 3928 12555 3950
rect 12594 3928 12628 3950
rect 12667 3928 12701 3950
rect 12740 3928 12774 3950
rect 12813 3928 12847 3950
rect 12886 3928 12920 3950
rect 12959 3928 12993 3950
rect 13032 3928 13066 3950
rect 13105 3928 13139 3950
rect 13178 3928 13212 3950
rect 13251 3928 13285 3950
rect 13324 3928 13358 3950
rect 13397 3928 13431 3950
rect 13470 3928 13504 3950
rect 13543 3928 13577 3950
rect 13616 3928 13650 3950
rect 13689 3928 13723 3950
rect 13762 3928 13796 3950
rect 13835 3928 13869 3950
rect 13908 3928 13942 3950
rect 13981 3928 14015 3950
rect 14054 3928 14088 3962
rect 14127 3950 14157 3962
rect 14157 3950 14161 3962
rect 14200 3950 14226 3962
rect 14226 3950 14234 3962
rect 14273 3950 14295 3962
rect 14295 3950 14307 3962
rect 14346 3950 14364 3962
rect 14364 3950 14380 3962
rect 14419 3950 14433 3962
rect 14433 3950 14453 3962
rect 14492 3950 14502 3962
rect 14502 3950 14526 3962
rect 14565 3950 14571 3962
rect 14571 3950 14599 3962
rect 14638 3950 14640 3962
rect 14640 3950 14672 3962
rect 14711 3950 14743 3962
rect 14743 3950 14745 3962
rect 14784 3950 14812 3962
rect 14812 3950 14818 3962
rect 14857 3950 14881 3962
rect 14881 3950 14891 3962
rect 14930 3950 14950 3962
rect 14950 3950 14964 3962
rect 15003 3950 15019 3962
rect 15019 3950 15037 3962
rect 15076 3950 15088 3962
rect 15088 3950 15110 3962
rect 15149 3950 15157 3962
rect 15157 3950 15183 3962
rect 15222 3950 15226 3962
rect 15226 3950 15256 3962
rect 14127 3928 14161 3950
rect 14200 3928 14234 3950
rect 14273 3928 14307 3950
rect 14346 3928 14380 3950
rect 14419 3928 14453 3950
rect 14492 3928 14526 3950
rect 14565 3928 14599 3950
rect 14638 3928 14672 3950
rect 14711 3928 14745 3950
rect 14784 3928 14818 3950
rect 14857 3928 14891 3950
rect 14930 3928 14964 3950
rect 15003 3928 15037 3950
rect 15076 3928 15110 3950
rect 15149 3928 15183 3950
rect 15222 3928 15256 3950
rect 15295 3928 15329 3962
rect 15368 3950 15399 3962
rect 15399 3950 15402 3962
rect 15441 3950 15468 3962
rect 15468 3950 15475 3962
rect 15514 3950 15537 3962
rect 15537 3950 15548 3962
rect 15587 3950 15606 3962
rect 15606 3950 15621 3962
rect 15660 3950 15675 3962
rect 15675 3950 15694 3962
rect 15733 3950 15744 3962
rect 15744 3950 15767 3962
rect 15806 3950 15813 3962
rect 15813 3950 15840 3962
rect 15879 3950 15882 3962
rect 15882 3950 15913 3962
rect 15952 3950 15985 3962
rect 15985 3950 15986 3962
rect 16025 3950 16054 3962
rect 16054 3950 16059 3962
rect 16098 3950 16123 3962
rect 16123 3950 16132 3962
rect 16171 3950 16192 3962
rect 16192 3950 16205 3962
rect 16244 3950 16261 3962
rect 16261 3950 16278 3962
rect 16317 3950 16330 3962
rect 16330 3950 16351 3962
rect 15368 3928 15402 3950
rect 15441 3928 15475 3950
rect 15514 3928 15548 3950
rect 15587 3928 15621 3950
rect 15660 3928 15694 3950
rect 15733 3928 15767 3950
rect 15806 3928 15840 3950
rect 15879 3928 15913 3950
rect 15952 3928 15986 3950
rect 16025 3928 16059 3950
rect 16098 3928 16132 3950
rect 16171 3928 16205 3950
rect 16244 3928 16278 3950
rect 16317 3928 16351 3950
rect 11937 3882 11949 3890
rect 11949 3882 11971 3890
rect 12010 3882 12018 3890
rect 12018 3882 12044 3890
rect 12083 3882 12087 3890
rect 12087 3882 12117 3890
rect 12156 3882 12190 3890
rect 12229 3882 12259 3890
rect 12259 3882 12263 3890
rect 12302 3882 12328 3890
rect 12328 3882 12336 3890
rect 12375 3882 12397 3890
rect 12397 3882 12409 3890
rect 12448 3882 12466 3890
rect 12466 3882 12482 3890
rect 12521 3882 12535 3890
rect 12535 3882 12555 3890
rect 12594 3882 12604 3890
rect 12604 3882 12628 3890
rect 12667 3882 12673 3890
rect 12673 3882 12701 3890
rect 12740 3882 12742 3890
rect 12742 3882 12774 3890
rect 12813 3882 12846 3890
rect 12846 3882 12847 3890
rect 12886 3882 12915 3890
rect 12915 3882 12920 3890
rect 12959 3882 12984 3890
rect 12984 3882 12993 3890
rect 13032 3882 13053 3890
rect 13053 3882 13066 3890
rect 13105 3882 13122 3890
rect 13122 3882 13139 3890
rect 13178 3882 13191 3890
rect 13191 3882 13212 3890
rect 13251 3882 13260 3890
rect 13260 3882 13285 3890
rect 13324 3882 13329 3890
rect 13329 3882 13358 3890
rect 13397 3882 13398 3890
rect 13398 3882 13431 3890
rect 13470 3882 13501 3890
rect 13501 3882 13504 3890
rect 13543 3882 13570 3890
rect 13570 3882 13577 3890
rect 13616 3882 13639 3890
rect 13639 3882 13650 3890
rect 13689 3882 13708 3890
rect 13708 3882 13723 3890
rect 13762 3882 13777 3890
rect 13777 3882 13796 3890
rect 13835 3882 13846 3890
rect 13846 3882 13869 3890
rect 13908 3882 13915 3890
rect 13915 3882 13942 3890
rect 13981 3882 13984 3890
rect 13984 3882 14015 3890
rect 11937 3856 11971 3882
rect 12010 3856 12044 3882
rect 12083 3856 12117 3882
rect 12156 3856 12190 3882
rect 12229 3856 12263 3882
rect 12302 3856 12336 3882
rect 12375 3856 12409 3882
rect 12448 3856 12482 3882
rect 12521 3856 12555 3882
rect 12594 3856 12628 3882
rect 12667 3856 12701 3882
rect 12740 3856 12774 3882
rect 12813 3856 12847 3882
rect 12886 3856 12920 3882
rect 12959 3856 12993 3882
rect 13032 3856 13066 3882
rect 13105 3856 13139 3882
rect 13178 3856 13212 3882
rect 13251 3856 13285 3882
rect 13324 3856 13358 3882
rect 13397 3856 13431 3882
rect 13470 3856 13504 3882
rect 13543 3856 13577 3882
rect 13616 3856 13650 3882
rect 13689 3856 13723 3882
rect 13762 3856 13796 3882
rect 13835 3856 13869 3882
rect 13908 3856 13942 3882
rect 13981 3856 14015 3882
rect 14054 3856 14088 3890
rect 14127 3882 14157 3890
rect 14157 3882 14161 3890
rect 14200 3882 14226 3890
rect 14226 3882 14234 3890
rect 14273 3882 14295 3890
rect 14295 3882 14307 3890
rect 14346 3882 14364 3890
rect 14364 3882 14380 3890
rect 14419 3882 14433 3890
rect 14433 3882 14453 3890
rect 14492 3882 14502 3890
rect 14502 3882 14526 3890
rect 14565 3882 14571 3890
rect 14571 3882 14599 3890
rect 14638 3882 14640 3890
rect 14640 3882 14672 3890
rect 14711 3882 14743 3890
rect 14743 3882 14745 3890
rect 14784 3882 14812 3890
rect 14812 3882 14818 3890
rect 14857 3882 14881 3890
rect 14881 3882 14891 3890
rect 14930 3882 14950 3890
rect 14950 3882 14964 3890
rect 15003 3882 15019 3890
rect 15019 3882 15037 3890
rect 15076 3882 15088 3890
rect 15088 3882 15110 3890
rect 15149 3882 15157 3890
rect 15157 3882 15183 3890
rect 15222 3882 15226 3890
rect 15226 3882 15256 3890
rect 14127 3856 14161 3882
rect 14200 3856 14234 3882
rect 14273 3856 14307 3882
rect 14346 3856 14380 3882
rect 14419 3856 14453 3882
rect 14492 3856 14526 3882
rect 14565 3856 14599 3882
rect 14638 3856 14672 3882
rect 14711 3856 14745 3882
rect 14784 3856 14818 3882
rect 14857 3856 14891 3882
rect 14930 3856 14964 3882
rect 15003 3856 15037 3882
rect 15076 3856 15110 3882
rect 15149 3856 15183 3882
rect 15222 3856 15256 3882
rect 15295 3856 15329 3890
rect 15368 3882 15399 3890
rect 15399 3882 15402 3890
rect 15441 3882 15468 3890
rect 15468 3882 15475 3890
rect 15514 3882 15537 3890
rect 15537 3882 15548 3890
rect 15587 3882 15606 3890
rect 15606 3882 15621 3890
rect 15660 3882 15675 3890
rect 15675 3882 15694 3890
rect 15733 3882 15744 3890
rect 15744 3882 15767 3890
rect 15806 3882 15813 3890
rect 15813 3882 15840 3890
rect 15879 3882 15882 3890
rect 15882 3882 15913 3890
rect 15952 3882 15985 3890
rect 15985 3882 15986 3890
rect 16025 3882 16054 3890
rect 16054 3882 16059 3890
rect 16098 3882 16123 3890
rect 16123 3882 16132 3890
rect 16171 3882 16192 3890
rect 16192 3882 16205 3890
rect 16244 3882 16261 3890
rect 16261 3882 16278 3890
rect 16317 3882 16330 3890
rect 16330 3882 16351 3890
rect 15368 3856 15402 3882
rect 15441 3856 15475 3882
rect 15514 3856 15548 3882
rect 15587 3856 15621 3882
rect 15660 3856 15694 3882
rect 15733 3856 15767 3882
rect 15806 3856 15840 3882
rect 15879 3856 15913 3882
rect 15952 3856 15986 3882
rect 16025 3856 16059 3882
rect 16098 3856 16132 3882
rect 16171 3856 16205 3882
rect 16244 3856 16278 3882
rect 16317 3856 16351 3882
rect 16390 3856 16928 4322
rect 11953 3576 11987 3609
rect 12026 3576 12060 3609
rect 12099 3576 12133 3609
rect 12172 3576 12206 3609
rect 12245 3576 12279 3609
rect 12318 3576 12352 3609
rect 12391 3576 12425 3609
rect 12464 3576 12498 3609
rect 12537 3576 12571 3609
rect 12610 3576 12644 3609
rect 12683 3576 12717 3609
rect 12756 3576 12790 3609
rect 12829 3576 12863 3609
rect 12902 3576 12936 3609
rect 12975 3576 13009 3609
rect 13048 3576 13082 3609
rect 13121 3576 13155 3609
rect 13194 3576 13228 3609
rect 13267 3576 13301 3609
rect 13340 3576 13374 3609
rect 13413 3576 13447 3609
rect 13486 3576 13520 3609
rect 13559 3576 13593 3609
rect 13632 3576 13666 3609
rect 13705 3576 13739 3609
rect 45 3374 79 3408
rect 45 3306 79 3336
rect 45 3302 79 3306
rect 11953 3575 11983 3576
rect 11983 3575 11987 3576
rect 12026 3575 12052 3576
rect 12052 3575 12060 3576
rect 12099 3575 12121 3576
rect 12121 3575 12133 3576
rect 12172 3575 12190 3576
rect 12190 3575 12206 3576
rect 12245 3575 12259 3576
rect 12259 3575 12279 3576
rect 12318 3575 12328 3576
rect 12328 3575 12352 3576
rect 12391 3575 12397 3576
rect 12397 3575 12425 3576
rect 12464 3575 12466 3576
rect 12466 3575 12498 3576
rect 12537 3575 12570 3576
rect 12570 3575 12571 3576
rect 12610 3575 12639 3576
rect 12639 3575 12644 3576
rect 12683 3575 12708 3576
rect 12708 3575 12717 3576
rect 12756 3575 12777 3576
rect 12777 3575 12790 3576
rect 12829 3575 12846 3576
rect 12846 3575 12863 3576
rect 12902 3575 12915 3576
rect 12915 3575 12936 3576
rect 12975 3575 12984 3576
rect 12984 3575 13009 3576
rect 13048 3575 13053 3576
rect 13053 3575 13082 3576
rect 13121 3575 13122 3576
rect 13122 3575 13155 3576
rect 13194 3575 13225 3576
rect 13225 3575 13228 3576
rect 13267 3575 13294 3576
rect 13294 3575 13301 3576
rect 13340 3575 13363 3576
rect 13363 3575 13374 3576
rect 13413 3575 13432 3576
rect 13432 3575 13447 3576
rect 13486 3575 13501 3576
rect 13501 3575 13520 3576
rect 13559 3575 13570 3576
rect 13570 3575 13593 3576
rect 13632 3575 13639 3576
rect 13639 3575 13666 3576
rect 13705 3575 13708 3576
rect 13708 3575 13739 3576
rect 13778 3575 13812 3609
rect 13851 3576 13885 3609
rect 13924 3576 13958 3609
rect 13997 3576 14031 3609
rect 14070 3576 14104 3609
rect 14143 3576 14177 3609
rect 14216 3576 14250 3609
rect 14289 3576 14323 3609
rect 14362 3576 14396 3609
rect 14435 3576 14469 3609
rect 14508 3576 14542 3609
rect 14581 3576 14615 3609
rect 14654 3576 14688 3609
rect 14727 3576 14761 3609
rect 14800 3576 14834 3609
rect 14873 3576 14907 3609
rect 14946 3576 14980 3609
rect 13851 3575 13881 3576
rect 13881 3575 13885 3576
rect 13924 3575 13950 3576
rect 13950 3575 13958 3576
rect 13997 3575 14019 3576
rect 14019 3575 14031 3576
rect 14070 3575 14088 3576
rect 14088 3575 14104 3576
rect 14143 3575 14157 3576
rect 14157 3575 14177 3576
rect 14216 3575 14226 3576
rect 14226 3575 14250 3576
rect 14289 3575 14295 3576
rect 14295 3575 14323 3576
rect 14362 3575 14364 3576
rect 14364 3575 14396 3576
rect 14435 3575 14467 3576
rect 14467 3575 14469 3576
rect 14508 3575 14536 3576
rect 14536 3575 14542 3576
rect 14581 3575 14605 3576
rect 14605 3575 14615 3576
rect 14654 3575 14674 3576
rect 14674 3575 14688 3576
rect 14727 3575 14743 3576
rect 14743 3575 14761 3576
rect 14800 3575 14812 3576
rect 14812 3575 14834 3576
rect 14873 3575 14881 3576
rect 14881 3575 14907 3576
rect 14946 3575 14950 3576
rect 14950 3575 14980 3576
rect 15019 3575 15053 3609
rect 15092 3576 15126 3609
rect 15165 3576 15199 3609
rect 15238 3576 15272 3609
rect 15311 3576 15345 3609
rect 15384 3576 15418 3609
rect 15457 3576 15491 3609
rect 15530 3576 15564 3609
rect 15603 3576 15637 3609
rect 15676 3576 15710 3609
rect 15749 3576 15783 3609
rect 15822 3576 15856 3609
rect 15895 3576 15929 3609
rect 15968 3576 16002 3609
rect 16041 3576 16075 3609
rect 16114 3576 16148 3609
rect 16187 3576 16221 3609
rect 16260 3576 16294 3609
rect 15092 3575 15123 3576
rect 15123 3575 15126 3576
rect 15165 3575 15192 3576
rect 15192 3575 15199 3576
rect 15238 3575 15261 3576
rect 15261 3575 15272 3576
rect 15311 3575 15330 3576
rect 15330 3575 15345 3576
rect 15384 3575 15399 3576
rect 15399 3575 15418 3576
rect 15457 3575 15468 3576
rect 15468 3575 15491 3576
rect 15530 3575 15537 3576
rect 15537 3575 15564 3576
rect 15603 3575 15606 3576
rect 15606 3575 15637 3576
rect 15676 3575 15709 3576
rect 15709 3575 15710 3576
rect 15749 3575 15778 3576
rect 15778 3575 15783 3576
rect 15822 3575 15847 3576
rect 15847 3575 15856 3576
rect 15895 3575 15916 3576
rect 15916 3575 15929 3576
rect 15968 3575 15985 3576
rect 15985 3575 16002 3576
rect 16041 3575 16054 3576
rect 16054 3575 16075 3576
rect 16114 3575 16123 3576
rect 16123 3575 16148 3576
rect 16187 3575 16192 3576
rect 16192 3575 16221 3576
rect 16260 3575 16261 3576
rect 16261 3575 16294 3576
rect 16333 3575 16365 3609
rect 16365 3575 16367 3609
rect 11953 3508 11987 3537
rect 12026 3508 12060 3537
rect 12099 3508 12133 3537
rect 12172 3508 12206 3537
rect 12245 3508 12279 3537
rect 12318 3508 12352 3537
rect 12391 3508 12425 3537
rect 12464 3508 12498 3537
rect 12537 3508 12571 3537
rect 12610 3508 12644 3537
rect 12683 3508 12717 3537
rect 12756 3508 12790 3537
rect 12829 3508 12863 3537
rect 12902 3508 12936 3537
rect 12975 3508 13009 3537
rect 13048 3508 13082 3537
rect 13121 3508 13155 3537
rect 13194 3508 13228 3537
rect 13267 3508 13301 3537
rect 13340 3508 13374 3537
rect 13413 3508 13447 3537
rect 13486 3508 13520 3537
rect 13559 3508 13593 3537
rect 13632 3508 13666 3537
rect 13705 3508 13739 3537
rect 11953 3503 11983 3508
rect 11983 3503 11987 3508
rect 12026 3503 12052 3508
rect 12052 3503 12060 3508
rect 12099 3503 12121 3508
rect 12121 3503 12133 3508
rect 12172 3503 12190 3508
rect 12190 3503 12206 3508
rect 12245 3503 12259 3508
rect 12259 3503 12279 3508
rect 12318 3503 12328 3508
rect 12328 3503 12352 3508
rect 12391 3503 12397 3508
rect 12397 3503 12425 3508
rect 12464 3503 12466 3508
rect 12466 3503 12498 3508
rect 12537 3503 12570 3508
rect 12570 3503 12571 3508
rect 12610 3503 12639 3508
rect 12639 3503 12644 3508
rect 12683 3503 12708 3508
rect 12708 3503 12717 3508
rect 12756 3503 12777 3508
rect 12777 3503 12790 3508
rect 12829 3503 12846 3508
rect 12846 3503 12863 3508
rect 12902 3503 12915 3508
rect 12915 3503 12936 3508
rect 12975 3503 12984 3508
rect 12984 3503 13009 3508
rect 13048 3503 13053 3508
rect 13053 3503 13082 3508
rect 13121 3503 13122 3508
rect 13122 3503 13155 3508
rect 13194 3503 13225 3508
rect 13225 3503 13228 3508
rect 13267 3503 13294 3508
rect 13294 3503 13301 3508
rect 13340 3503 13363 3508
rect 13363 3503 13374 3508
rect 13413 3503 13432 3508
rect 13432 3503 13447 3508
rect 13486 3503 13501 3508
rect 13501 3503 13520 3508
rect 13559 3503 13570 3508
rect 13570 3503 13593 3508
rect 13632 3503 13639 3508
rect 13639 3503 13666 3508
rect 13705 3503 13708 3508
rect 13708 3503 13739 3508
rect 13778 3503 13812 3537
rect 13851 3508 13885 3537
rect 13924 3508 13958 3537
rect 13997 3508 14031 3537
rect 14070 3508 14104 3537
rect 14143 3508 14177 3537
rect 14216 3508 14250 3537
rect 14289 3508 14323 3537
rect 14362 3508 14396 3537
rect 14435 3508 14469 3537
rect 14508 3508 14542 3537
rect 14581 3508 14615 3537
rect 14654 3508 14688 3537
rect 14727 3508 14761 3537
rect 14800 3508 14834 3537
rect 14873 3508 14907 3537
rect 14946 3508 14980 3537
rect 13851 3503 13881 3508
rect 13881 3503 13885 3508
rect 13924 3503 13950 3508
rect 13950 3503 13958 3508
rect 13997 3503 14019 3508
rect 14019 3503 14031 3508
rect 14070 3503 14088 3508
rect 14088 3503 14104 3508
rect 14143 3503 14157 3508
rect 14157 3503 14177 3508
rect 14216 3503 14226 3508
rect 14226 3503 14250 3508
rect 14289 3503 14295 3508
rect 14295 3503 14323 3508
rect 14362 3503 14364 3508
rect 14364 3503 14396 3508
rect 14435 3503 14467 3508
rect 14467 3503 14469 3508
rect 14508 3503 14536 3508
rect 14536 3503 14542 3508
rect 14581 3503 14605 3508
rect 14605 3503 14615 3508
rect 14654 3503 14674 3508
rect 14674 3503 14688 3508
rect 14727 3503 14743 3508
rect 14743 3503 14761 3508
rect 14800 3503 14812 3508
rect 14812 3503 14834 3508
rect 14873 3503 14881 3508
rect 14881 3503 14907 3508
rect 14946 3503 14950 3508
rect 14950 3503 14980 3508
rect 15019 3503 15053 3537
rect 15092 3508 15126 3537
rect 15165 3508 15199 3537
rect 15238 3508 15272 3537
rect 15311 3508 15345 3537
rect 15384 3508 15418 3537
rect 15457 3508 15491 3537
rect 15530 3508 15564 3537
rect 15603 3508 15637 3537
rect 15676 3508 15710 3537
rect 15749 3508 15783 3537
rect 15822 3508 15856 3537
rect 15895 3508 15929 3537
rect 15968 3508 16002 3537
rect 16041 3508 16075 3537
rect 16114 3508 16148 3537
rect 16187 3508 16221 3537
rect 16260 3508 16294 3537
rect 15092 3503 15123 3508
rect 15123 3503 15126 3508
rect 15165 3503 15192 3508
rect 15192 3503 15199 3508
rect 15238 3503 15261 3508
rect 15261 3503 15272 3508
rect 15311 3503 15330 3508
rect 15330 3503 15345 3508
rect 15384 3503 15399 3508
rect 15399 3503 15418 3508
rect 15457 3503 15468 3508
rect 15468 3503 15491 3508
rect 15530 3503 15537 3508
rect 15537 3503 15564 3508
rect 15603 3503 15606 3508
rect 15606 3503 15637 3508
rect 15676 3503 15709 3508
rect 15709 3503 15710 3508
rect 15749 3503 15778 3508
rect 15778 3503 15783 3508
rect 15822 3503 15847 3508
rect 15847 3503 15856 3508
rect 15895 3503 15916 3508
rect 15916 3503 15929 3508
rect 15968 3503 15985 3508
rect 15985 3503 16002 3508
rect 16041 3503 16054 3508
rect 16054 3503 16075 3508
rect 16114 3503 16123 3508
rect 16123 3503 16148 3508
rect 16187 3503 16192 3508
rect 16192 3503 16221 3508
rect 16260 3503 16261 3508
rect 16261 3503 16294 3508
rect 16333 3503 16365 3537
rect 16365 3503 16367 3537
rect 11953 3440 11987 3465
rect 12026 3440 12060 3465
rect 12099 3440 12133 3465
rect 12172 3440 12206 3465
rect 12245 3440 12279 3465
rect 12318 3440 12352 3465
rect 12391 3440 12425 3465
rect 12464 3440 12498 3465
rect 12537 3440 12571 3465
rect 12610 3440 12644 3465
rect 12683 3440 12717 3465
rect 12756 3440 12790 3465
rect 12829 3440 12863 3465
rect 12902 3440 12936 3465
rect 12975 3440 13009 3465
rect 13048 3440 13082 3465
rect 13121 3440 13155 3465
rect 13194 3440 13228 3465
rect 13267 3440 13301 3465
rect 13340 3440 13374 3465
rect 13413 3440 13447 3465
rect 13486 3440 13520 3465
rect 13559 3440 13593 3465
rect 13632 3440 13666 3465
rect 13705 3440 13739 3465
rect 11953 3431 11983 3440
rect 11983 3431 11987 3440
rect 12026 3431 12052 3440
rect 12052 3431 12060 3440
rect 12099 3431 12121 3440
rect 12121 3431 12133 3440
rect 12172 3431 12190 3440
rect 12190 3431 12206 3440
rect 12245 3431 12259 3440
rect 12259 3431 12279 3440
rect 12318 3431 12328 3440
rect 12328 3431 12352 3440
rect 12391 3431 12397 3440
rect 12397 3431 12425 3440
rect 12464 3431 12466 3440
rect 12466 3431 12498 3440
rect 12537 3431 12570 3440
rect 12570 3431 12571 3440
rect 12610 3431 12639 3440
rect 12639 3431 12644 3440
rect 12683 3431 12708 3440
rect 12708 3431 12717 3440
rect 12756 3431 12777 3440
rect 12777 3431 12790 3440
rect 12829 3431 12846 3440
rect 12846 3431 12863 3440
rect 12902 3431 12915 3440
rect 12915 3431 12936 3440
rect 12975 3431 12984 3440
rect 12984 3431 13009 3440
rect 13048 3431 13053 3440
rect 13053 3431 13082 3440
rect 13121 3431 13122 3440
rect 13122 3431 13155 3440
rect 13194 3431 13225 3440
rect 13225 3431 13228 3440
rect 13267 3431 13294 3440
rect 13294 3431 13301 3440
rect 13340 3431 13363 3440
rect 13363 3431 13374 3440
rect 13413 3431 13432 3440
rect 13432 3431 13447 3440
rect 13486 3431 13501 3440
rect 13501 3431 13520 3440
rect 13559 3431 13570 3440
rect 13570 3431 13593 3440
rect 13632 3431 13639 3440
rect 13639 3431 13666 3440
rect 13705 3431 13708 3440
rect 13708 3431 13739 3440
rect 13778 3431 13812 3465
rect 13851 3440 13885 3465
rect 13924 3440 13958 3465
rect 13997 3440 14031 3465
rect 14070 3440 14104 3465
rect 14143 3440 14177 3465
rect 14216 3440 14250 3465
rect 14289 3440 14323 3465
rect 14362 3440 14396 3465
rect 14435 3440 14469 3465
rect 14508 3440 14542 3465
rect 14581 3440 14615 3465
rect 14654 3440 14688 3465
rect 14727 3440 14761 3465
rect 14800 3440 14834 3465
rect 14873 3440 14907 3465
rect 14946 3440 14980 3465
rect 13851 3431 13881 3440
rect 13881 3431 13885 3440
rect 13924 3431 13950 3440
rect 13950 3431 13958 3440
rect 13997 3431 14019 3440
rect 14019 3431 14031 3440
rect 14070 3431 14088 3440
rect 14088 3431 14104 3440
rect 14143 3431 14157 3440
rect 14157 3431 14177 3440
rect 14216 3431 14226 3440
rect 14226 3431 14250 3440
rect 14289 3431 14295 3440
rect 14295 3431 14323 3440
rect 14362 3431 14364 3440
rect 14364 3431 14396 3440
rect 14435 3431 14467 3440
rect 14467 3431 14469 3440
rect 14508 3431 14536 3440
rect 14536 3431 14542 3440
rect 14581 3431 14605 3440
rect 14605 3431 14615 3440
rect 14654 3431 14674 3440
rect 14674 3431 14688 3440
rect 14727 3431 14743 3440
rect 14743 3431 14761 3440
rect 14800 3431 14812 3440
rect 14812 3431 14834 3440
rect 14873 3431 14881 3440
rect 14881 3431 14907 3440
rect 14946 3431 14950 3440
rect 14950 3431 14980 3440
rect 15019 3431 15053 3465
rect 15092 3440 15126 3465
rect 15165 3440 15199 3465
rect 15238 3440 15272 3465
rect 15311 3440 15345 3465
rect 15384 3440 15418 3465
rect 15457 3440 15491 3465
rect 15530 3440 15564 3465
rect 15603 3440 15637 3465
rect 15676 3440 15710 3465
rect 15749 3440 15783 3465
rect 15822 3440 15856 3465
rect 15895 3440 15929 3465
rect 15968 3440 16002 3465
rect 16041 3440 16075 3465
rect 16114 3440 16148 3465
rect 16187 3440 16221 3465
rect 16260 3440 16294 3465
rect 15092 3431 15123 3440
rect 15123 3431 15126 3440
rect 15165 3431 15192 3440
rect 15192 3431 15199 3440
rect 15238 3431 15261 3440
rect 15261 3431 15272 3440
rect 15311 3431 15330 3440
rect 15330 3431 15345 3440
rect 15384 3431 15399 3440
rect 15399 3431 15418 3440
rect 15457 3431 15468 3440
rect 15468 3431 15491 3440
rect 15530 3431 15537 3440
rect 15537 3431 15564 3440
rect 15603 3431 15606 3440
rect 15606 3431 15637 3440
rect 15676 3431 15709 3440
rect 15709 3431 15710 3440
rect 15749 3431 15778 3440
rect 15778 3431 15783 3440
rect 15822 3431 15847 3440
rect 15847 3431 15856 3440
rect 15895 3431 15916 3440
rect 15916 3431 15929 3440
rect 15968 3431 15985 3440
rect 15985 3431 16002 3440
rect 16041 3431 16054 3440
rect 16054 3431 16075 3440
rect 16114 3431 16123 3440
rect 16123 3431 16148 3440
rect 16187 3431 16192 3440
rect 16192 3431 16221 3440
rect 16260 3431 16261 3440
rect 16261 3431 16294 3440
rect 16333 3431 16365 3465
rect 16365 3431 16367 3465
rect 11953 3372 11987 3393
rect 12026 3372 12060 3393
rect 12099 3372 12133 3393
rect 12172 3372 12206 3393
rect 12245 3372 12279 3393
rect 12318 3372 12352 3393
rect 12391 3372 12425 3393
rect 12464 3372 12498 3393
rect 12537 3372 12571 3393
rect 12610 3372 12644 3393
rect 12683 3372 12717 3393
rect 12756 3372 12790 3393
rect 12829 3372 12863 3393
rect 12902 3372 12936 3393
rect 12975 3372 13009 3393
rect 13048 3372 13082 3393
rect 13121 3372 13155 3393
rect 13194 3372 13228 3393
rect 13267 3372 13301 3393
rect 13340 3372 13374 3393
rect 13413 3372 13447 3393
rect 13486 3372 13520 3393
rect 13559 3372 13593 3393
rect 13632 3372 13666 3393
rect 13705 3372 13739 3393
rect 11953 3359 11983 3372
rect 11983 3359 11987 3372
rect 12026 3359 12052 3372
rect 12052 3359 12060 3372
rect 12099 3359 12121 3372
rect 12121 3359 12133 3372
rect 12172 3359 12190 3372
rect 12190 3359 12206 3372
rect 12245 3359 12259 3372
rect 12259 3359 12279 3372
rect 12318 3359 12328 3372
rect 12328 3359 12352 3372
rect 12391 3359 12397 3372
rect 12397 3359 12425 3372
rect 12464 3359 12466 3372
rect 12466 3359 12498 3372
rect 12537 3359 12570 3372
rect 12570 3359 12571 3372
rect 12610 3359 12639 3372
rect 12639 3359 12644 3372
rect 12683 3359 12708 3372
rect 12708 3359 12717 3372
rect 12756 3359 12777 3372
rect 12777 3359 12790 3372
rect 12829 3359 12846 3372
rect 12846 3359 12863 3372
rect 12902 3359 12915 3372
rect 12915 3359 12936 3372
rect 12975 3359 12984 3372
rect 12984 3359 13009 3372
rect 13048 3359 13053 3372
rect 13053 3359 13082 3372
rect 13121 3359 13122 3372
rect 13122 3359 13155 3372
rect 13194 3359 13225 3372
rect 13225 3359 13228 3372
rect 13267 3359 13294 3372
rect 13294 3359 13301 3372
rect 13340 3359 13363 3372
rect 13363 3359 13374 3372
rect 13413 3359 13432 3372
rect 13432 3359 13447 3372
rect 13486 3359 13501 3372
rect 13501 3359 13520 3372
rect 13559 3359 13570 3372
rect 13570 3359 13593 3372
rect 13632 3359 13639 3372
rect 13639 3359 13666 3372
rect 13705 3359 13708 3372
rect 13708 3359 13739 3372
rect 13778 3359 13812 3393
rect 13851 3372 13885 3393
rect 13924 3372 13958 3393
rect 13997 3372 14031 3393
rect 14070 3372 14104 3393
rect 14143 3372 14177 3393
rect 14216 3372 14250 3393
rect 14289 3372 14323 3393
rect 14362 3372 14396 3393
rect 14435 3372 14469 3393
rect 14508 3372 14542 3393
rect 14581 3372 14615 3393
rect 14654 3372 14688 3393
rect 14727 3372 14761 3393
rect 14800 3372 14834 3393
rect 14873 3372 14907 3393
rect 14946 3372 14980 3393
rect 13851 3359 13881 3372
rect 13881 3359 13885 3372
rect 13924 3359 13950 3372
rect 13950 3359 13958 3372
rect 13997 3359 14019 3372
rect 14019 3359 14031 3372
rect 14070 3359 14088 3372
rect 14088 3359 14104 3372
rect 14143 3359 14157 3372
rect 14157 3359 14177 3372
rect 14216 3359 14226 3372
rect 14226 3359 14250 3372
rect 14289 3359 14295 3372
rect 14295 3359 14323 3372
rect 14362 3359 14364 3372
rect 14364 3359 14396 3372
rect 14435 3359 14467 3372
rect 14467 3359 14469 3372
rect 14508 3359 14536 3372
rect 14536 3359 14542 3372
rect 14581 3359 14605 3372
rect 14605 3359 14615 3372
rect 14654 3359 14674 3372
rect 14674 3359 14688 3372
rect 14727 3359 14743 3372
rect 14743 3359 14761 3372
rect 14800 3359 14812 3372
rect 14812 3359 14834 3372
rect 14873 3359 14881 3372
rect 14881 3359 14907 3372
rect 14946 3359 14950 3372
rect 14950 3359 14980 3372
rect 15019 3359 15053 3393
rect 15092 3372 15126 3393
rect 15165 3372 15199 3393
rect 15238 3372 15272 3393
rect 15311 3372 15345 3393
rect 15384 3372 15418 3393
rect 15457 3372 15491 3393
rect 15530 3372 15564 3393
rect 15603 3372 15637 3393
rect 15676 3372 15710 3393
rect 15749 3372 15783 3393
rect 15822 3372 15856 3393
rect 15895 3372 15929 3393
rect 15968 3372 16002 3393
rect 16041 3372 16075 3393
rect 16114 3372 16148 3393
rect 16187 3372 16221 3393
rect 16260 3372 16294 3393
rect 15092 3359 15123 3372
rect 15123 3359 15126 3372
rect 15165 3359 15192 3372
rect 15192 3359 15199 3372
rect 15238 3359 15261 3372
rect 15261 3359 15272 3372
rect 15311 3359 15330 3372
rect 15330 3359 15345 3372
rect 15384 3359 15399 3372
rect 15399 3359 15418 3372
rect 15457 3359 15468 3372
rect 15468 3359 15491 3372
rect 15530 3359 15537 3372
rect 15537 3359 15564 3372
rect 15603 3359 15606 3372
rect 15606 3359 15637 3372
rect 15676 3359 15709 3372
rect 15709 3359 15710 3372
rect 15749 3359 15778 3372
rect 15778 3359 15783 3372
rect 15822 3359 15847 3372
rect 15847 3359 15856 3372
rect 15895 3359 15916 3372
rect 15916 3359 15929 3372
rect 15968 3359 15985 3372
rect 15985 3359 16002 3372
rect 16041 3359 16054 3372
rect 16054 3359 16075 3372
rect 16114 3359 16123 3372
rect 16123 3359 16148 3372
rect 16187 3359 16192 3372
rect 16192 3359 16221 3372
rect 16260 3359 16261 3372
rect 16261 3359 16294 3372
rect 16333 3359 16365 3393
rect 16365 3359 16367 3393
rect 11953 3304 11987 3321
rect 12026 3304 12060 3321
rect 12099 3304 12133 3321
rect 12172 3304 12206 3321
rect 12245 3304 12279 3321
rect 12318 3304 12352 3321
rect 12391 3304 12425 3321
rect 12464 3304 12498 3321
rect 12537 3304 12571 3321
rect 12610 3304 12644 3321
rect 12683 3304 12717 3321
rect 12756 3304 12790 3321
rect 12829 3304 12863 3321
rect 12902 3304 12936 3321
rect 12975 3304 13009 3321
rect 13048 3304 13082 3321
rect 13121 3304 13155 3321
rect 13194 3304 13228 3321
rect 13267 3304 13301 3321
rect 13340 3304 13374 3321
rect 13413 3304 13447 3321
rect 13486 3304 13520 3321
rect 13559 3304 13593 3321
rect 13632 3304 13666 3321
rect 13705 3304 13739 3321
rect 11953 3287 11983 3304
rect 11983 3287 11987 3304
rect 12026 3287 12052 3304
rect 12052 3287 12060 3304
rect 12099 3287 12121 3304
rect 12121 3287 12133 3304
rect 12172 3287 12190 3304
rect 12190 3287 12206 3304
rect 12245 3287 12259 3304
rect 12259 3287 12279 3304
rect 12318 3287 12328 3304
rect 12328 3287 12352 3304
rect 12391 3287 12397 3304
rect 12397 3287 12425 3304
rect 12464 3287 12466 3304
rect 12466 3287 12498 3304
rect 12537 3287 12570 3304
rect 12570 3287 12571 3304
rect 12610 3287 12639 3304
rect 12639 3287 12644 3304
rect 12683 3287 12708 3304
rect 12708 3287 12717 3304
rect 12756 3287 12777 3304
rect 12777 3287 12790 3304
rect 12829 3287 12846 3304
rect 12846 3287 12863 3304
rect 12902 3287 12915 3304
rect 12915 3287 12936 3304
rect 12975 3287 12984 3304
rect 12984 3287 13009 3304
rect 13048 3287 13053 3304
rect 13053 3287 13082 3304
rect 13121 3287 13122 3304
rect 13122 3287 13155 3304
rect 13194 3287 13225 3304
rect 13225 3287 13228 3304
rect 13267 3287 13294 3304
rect 13294 3287 13301 3304
rect 13340 3287 13363 3304
rect 13363 3287 13374 3304
rect 13413 3287 13432 3304
rect 13432 3287 13447 3304
rect 13486 3287 13501 3304
rect 13501 3287 13520 3304
rect 13559 3287 13570 3304
rect 13570 3287 13593 3304
rect 13632 3287 13639 3304
rect 13639 3287 13666 3304
rect 13705 3287 13708 3304
rect 13708 3287 13739 3304
rect 13778 3287 13812 3321
rect 13851 3304 13885 3321
rect 13924 3304 13958 3321
rect 13997 3304 14031 3321
rect 14070 3304 14104 3321
rect 14143 3304 14177 3321
rect 14216 3304 14250 3321
rect 14289 3304 14323 3321
rect 14362 3304 14396 3321
rect 14435 3304 14469 3321
rect 14508 3304 14542 3321
rect 14581 3304 14615 3321
rect 14654 3304 14688 3321
rect 14727 3304 14761 3321
rect 14800 3304 14834 3321
rect 14873 3304 14907 3321
rect 14946 3304 14980 3321
rect 13851 3287 13881 3304
rect 13881 3287 13885 3304
rect 13924 3287 13950 3304
rect 13950 3287 13958 3304
rect 13997 3287 14019 3304
rect 14019 3287 14031 3304
rect 14070 3287 14088 3304
rect 14088 3287 14104 3304
rect 14143 3287 14157 3304
rect 14157 3287 14177 3304
rect 14216 3287 14226 3304
rect 14226 3287 14250 3304
rect 14289 3287 14295 3304
rect 14295 3287 14323 3304
rect 14362 3287 14364 3304
rect 14364 3287 14396 3304
rect 14435 3287 14467 3304
rect 14467 3287 14469 3304
rect 14508 3287 14536 3304
rect 14536 3287 14542 3304
rect 14581 3287 14605 3304
rect 14605 3287 14615 3304
rect 14654 3287 14674 3304
rect 14674 3287 14688 3304
rect 14727 3287 14743 3304
rect 14743 3287 14761 3304
rect 14800 3287 14812 3304
rect 14812 3287 14834 3304
rect 14873 3287 14881 3304
rect 14881 3287 14907 3304
rect 14946 3287 14950 3304
rect 14950 3287 14980 3304
rect 15019 3287 15053 3321
rect 15092 3304 15126 3321
rect 15165 3304 15199 3321
rect 15238 3304 15272 3321
rect 15311 3304 15345 3321
rect 15384 3304 15418 3321
rect 15457 3304 15491 3321
rect 15530 3304 15564 3321
rect 15603 3304 15637 3321
rect 15676 3304 15710 3321
rect 15749 3304 15783 3321
rect 15822 3304 15856 3321
rect 15895 3304 15929 3321
rect 15968 3304 16002 3321
rect 16041 3304 16075 3321
rect 16114 3304 16148 3321
rect 16187 3304 16221 3321
rect 16260 3304 16294 3321
rect 15092 3287 15123 3304
rect 15123 3287 15126 3304
rect 15165 3287 15192 3304
rect 15192 3287 15199 3304
rect 15238 3287 15261 3304
rect 15261 3287 15272 3304
rect 15311 3287 15330 3304
rect 15330 3287 15345 3304
rect 15384 3287 15399 3304
rect 15399 3287 15418 3304
rect 15457 3287 15468 3304
rect 15468 3287 15491 3304
rect 15530 3287 15537 3304
rect 15537 3287 15564 3304
rect 15603 3287 15606 3304
rect 15606 3287 15637 3304
rect 15676 3287 15709 3304
rect 15709 3287 15710 3304
rect 15749 3287 15778 3304
rect 15778 3287 15783 3304
rect 15822 3287 15847 3304
rect 15847 3287 15856 3304
rect 15895 3287 15916 3304
rect 15916 3287 15929 3304
rect 15968 3287 15985 3304
rect 15985 3287 16002 3304
rect 16041 3287 16054 3304
rect 16054 3287 16075 3304
rect 16114 3287 16123 3304
rect 16123 3287 16148 3304
rect 16187 3287 16192 3304
rect 16192 3287 16221 3304
rect 16260 3287 16261 3304
rect 16261 3287 16294 3304
rect 16333 3287 16365 3321
rect 16365 3287 16367 3321
rect 16406 3270 16872 3609
rect 11953 3235 11987 3249
rect 12026 3235 12060 3249
rect 12099 3235 12133 3249
rect 12172 3235 12206 3249
rect 12245 3235 12279 3249
rect 12318 3235 12352 3249
rect 12391 3235 12425 3249
rect 12464 3235 12498 3249
rect 12537 3235 12571 3249
rect 12610 3235 12644 3249
rect 12683 3235 12717 3249
rect 12756 3235 12790 3249
rect 12829 3235 12863 3249
rect 12902 3235 12936 3249
rect 12975 3235 13009 3249
rect 13048 3235 13082 3249
rect 13121 3235 13155 3249
rect 13194 3235 13228 3249
rect 13267 3235 13301 3249
rect 13340 3235 13374 3249
rect 13413 3235 13447 3249
rect 13486 3235 13520 3249
rect 13559 3235 13593 3249
rect 13632 3235 13666 3249
rect 13705 3235 13739 3249
rect 13778 3235 13812 3249
rect 13851 3235 13885 3249
rect 13924 3235 13958 3249
rect 13997 3235 14031 3249
rect 14070 3235 14104 3249
rect 14143 3235 14177 3249
rect 14216 3235 14250 3249
rect 14289 3235 14323 3249
rect 14362 3235 14396 3249
rect 14435 3235 14469 3249
rect 14508 3235 14542 3249
rect 14581 3235 14615 3249
rect 14654 3235 14688 3249
rect 14727 3235 14761 3249
rect 14800 3235 14834 3249
rect 14873 3235 14907 3249
rect 14946 3235 14980 3249
rect 15019 3235 15053 3249
rect 15092 3235 15126 3249
rect 15165 3235 15199 3249
rect 15238 3235 15272 3249
rect 15311 3235 15345 3249
rect 15384 3235 15418 3249
rect 15457 3235 15491 3249
rect 15530 3235 15564 3249
rect 15603 3235 15637 3249
rect 15676 3235 15710 3249
rect 15749 3235 15783 3249
rect 15822 3235 15856 3249
rect 15895 3235 15929 3249
rect 15968 3235 16002 3249
rect 16041 3235 16075 3249
rect 16114 3235 16148 3249
rect 16187 3235 16221 3249
rect 16260 3235 16294 3249
rect 16333 3235 16367 3249
rect 16406 3235 16872 3270
rect 11953 3215 11987 3235
rect 12026 3215 12060 3235
rect 12099 3215 12133 3235
rect 12172 3215 12206 3235
rect 12245 3215 12279 3235
rect 12318 3215 12352 3235
rect 12391 3215 12425 3235
rect 12464 3215 12498 3235
rect 12537 3215 12571 3235
rect 12610 3215 12644 3235
rect 12683 3215 12717 3235
rect 12756 3215 12790 3235
rect 12829 3215 12863 3235
rect 12902 3215 12936 3235
rect 12975 3215 13009 3235
rect 13048 3215 13082 3235
rect 13121 3215 13155 3235
rect 13194 3215 13228 3235
rect 13267 3215 13301 3235
rect 13340 3215 13374 3235
rect 13413 3215 13447 3235
rect 13486 3215 13520 3235
rect 13559 3215 13593 3235
rect 13632 3215 13666 3235
rect 13705 3215 13739 3235
rect 13778 3215 13812 3235
rect 13851 3215 13885 3235
rect 13924 3215 13958 3235
rect 13997 3215 14031 3235
rect 14070 3215 14104 3235
rect 14143 3215 14177 3235
rect 14216 3215 14250 3235
rect 14289 3215 14323 3235
rect 14362 3215 14396 3235
rect 14435 3215 14469 3235
rect 14508 3215 14542 3235
rect 14581 3215 14615 3235
rect 14654 3215 14688 3235
rect 14727 3215 14761 3235
rect 14800 3215 14834 3235
rect 14873 3215 14907 3235
rect 14946 3215 14980 3235
rect 15019 3215 15053 3235
rect 15092 3215 15126 3235
rect 15165 3215 15199 3235
rect 15238 3215 15272 3235
rect 15311 3215 15345 3235
rect 15384 3215 15418 3235
rect 15457 3215 15491 3235
rect 15530 3215 15564 3235
rect 15603 3215 15637 3235
rect 15676 3215 15710 3235
rect 15749 3215 15783 3235
rect 15822 3215 15856 3235
rect 15895 3215 15929 3235
rect 15968 3215 16002 3235
rect 16041 3215 16075 3235
rect 16114 3215 16148 3235
rect 16187 3215 16221 3235
rect 16260 3215 16294 3235
rect 16333 3215 16367 3235
rect 11953 3143 11987 3177
rect 12026 3143 12060 3177
rect 12099 3143 12133 3177
rect 12172 3143 12206 3177
rect 12245 3143 12279 3177
rect 12318 3143 12352 3177
rect 12391 3143 12425 3177
rect 12464 3143 12498 3177
rect 12537 3143 12571 3177
rect 12610 3143 12644 3177
rect 12683 3143 12717 3177
rect 12756 3143 12790 3177
rect 12829 3143 12863 3177
rect 12902 3143 12936 3177
rect 12975 3143 13009 3177
rect 13048 3143 13082 3177
rect 13121 3143 13155 3177
rect 13194 3143 13228 3177
rect 13267 3143 13301 3177
rect 13340 3143 13374 3177
rect 13413 3143 13447 3177
rect 13486 3143 13520 3177
rect 13559 3143 13593 3177
rect 13632 3143 13666 3177
rect 13705 3143 13739 3177
rect 13778 3143 13812 3177
rect 13851 3143 13885 3177
rect 13924 3143 13958 3177
rect 13997 3143 14031 3177
rect 14070 3143 14104 3177
rect 14143 3143 14177 3177
rect 14216 3143 14250 3177
rect 14289 3143 14323 3177
rect 14362 3143 14396 3177
rect 14435 3143 14469 3177
rect 14508 3143 14542 3177
rect 14581 3143 14615 3177
rect 14654 3143 14688 3177
rect 14727 3143 14761 3177
rect 14800 3143 14834 3177
rect 14873 3143 14907 3177
rect 14946 3143 14980 3177
rect 15019 3143 15053 3177
rect 15092 3143 15126 3177
rect 15165 3143 15199 3177
rect 15238 3143 15272 3177
rect 15311 3143 15345 3177
rect 15384 3143 15418 3177
rect 15457 3143 15491 3177
rect 15530 3143 15564 3177
rect 15603 3143 15637 3177
rect 15676 3143 15710 3177
rect 15749 3143 15783 3177
rect 15822 3143 15856 3177
rect 15895 3143 15929 3177
rect 15968 3143 16002 3177
rect 16041 3143 16075 3177
rect 16114 3143 16148 3177
rect 16187 3143 16221 3177
rect 16260 3143 16294 3177
rect 16333 3143 16367 3177
rect 11953 3071 11987 3105
rect 12026 3071 12060 3105
rect 12099 3071 12133 3105
rect 12172 3071 12206 3105
rect 12245 3071 12279 3105
rect 12318 3071 12352 3105
rect 12391 3071 12425 3105
rect 12464 3071 12498 3105
rect 12537 3071 12571 3105
rect 12610 3071 12644 3105
rect 12683 3071 12717 3105
rect 12756 3071 12790 3105
rect 12829 3071 12863 3105
rect 12902 3071 12936 3105
rect 12975 3071 13009 3105
rect 13048 3071 13082 3105
rect 13121 3071 13155 3105
rect 13194 3071 13228 3105
rect 13267 3071 13301 3105
rect 13340 3071 13374 3105
rect 13413 3071 13447 3105
rect 13486 3071 13520 3105
rect 13559 3071 13593 3105
rect 13632 3071 13666 3105
rect 13705 3071 13739 3105
rect 13778 3071 13812 3105
rect 13851 3071 13885 3105
rect 13924 3071 13958 3105
rect 13997 3071 14031 3105
rect 14070 3071 14104 3105
rect 14143 3071 14177 3105
rect 14216 3071 14250 3105
rect 14289 3071 14323 3105
rect 14362 3071 14396 3105
rect 14435 3071 14469 3105
rect 14508 3071 14542 3105
rect 14581 3071 14615 3105
rect 14654 3071 14688 3105
rect 14727 3071 14761 3105
rect 14800 3071 14834 3105
rect 14873 3071 14907 3105
rect 14946 3071 14980 3105
rect 15019 3071 15053 3105
rect 15092 3071 15126 3105
rect 15165 3071 15199 3105
rect 15238 3071 15272 3105
rect 15311 3071 15345 3105
rect 15384 3071 15418 3105
rect 15457 3071 15491 3105
rect 15530 3071 15564 3105
rect 15603 3071 15637 3105
rect 15676 3071 15710 3105
rect 15749 3071 15783 3105
rect 15822 3071 15856 3105
rect 15895 3071 15929 3105
rect 15968 3071 16002 3105
rect 16041 3071 16075 3105
rect 16114 3071 16148 3105
rect 16187 3071 16221 3105
rect 16260 3071 16294 3105
rect 16333 3071 16367 3105
rect 11953 2999 11987 3033
rect 12026 2999 12060 3033
rect 12099 2999 12133 3033
rect 12172 2999 12206 3033
rect 12245 2999 12279 3033
rect 12318 2999 12352 3033
rect 12391 2999 12425 3033
rect 12464 2999 12498 3033
rect 12537 2999 12571 3033
rect 12610 2999 12644 3033
rect 12683 2999 12717 3033
rect 12756 2999 12790 3033
rect 12829 2999 12863 3033
rect 12902 2999 12936 3033
rect 12975 2999 13009 3033
rect 13048 2999 13082 3033
rect 13121 2999 13155 3033
rect 13194 2999 13228 3033
rect 13267 2999 13301 3033
rect 13340 2999 13374 3033
rect 13413 2999 13447 3033
rect 13486 2999 13520 3033
rect 13559 2999 13593 3033
rect 13632 2999 13666 3033
rect 13705 2999 13739 3033
rect 13778 2999 13812 3033
rect 13851 2999 13885 3033
rect 13924 2999 13958 3033
rect 13997 2999 14031 3033
rect 14070 2999 14104 3033
rect 14143 2999 14177 3033
rect 14216 2999 14250 3033
rect 14289 2999 14323 3033
rect 14362 2999 14396 3033
rect 14435 2999 14469 3033
rect 14508 2999 14542 3033
rect 14581 2999 14615 3033
rect 14654 2999 14688 3033
rect 14727 2999 14761 3033
rect 14800 2999 14834 3033
rect 14873 2999 14907 3033
rect 14946 2999 14980 3033
rect 15019 2999 15053 3033
rect 15092 2999 15126 3033
rect 15165 2999 15199 3033
rect 15238 2999 15272 3033
rect 15311 2999 15345 3033
rect 15384 2999 15418 3033
rect 15457 2999 15491 3033
rect 15530 2999 15564 3033
rect 15603 2999 15637 3033
rect 15676 2999 15710 3033
rect 15749 2999 15783 3033
rect 15822 2999 15856 3033
rect 15895 2999 15929 3033
rect 15968 2999 16002 3033
rect 16041 2999 16075 3033
rect 16114 2999 16148 3033
rect 16187 2999 16221 3033
rect 16260 2999 16294 3033
rect 16333 2999 16367 3033
rect 16406 2999 16872 3235
rect 4734 2691 4768 2715
rect 4807 2691 4841 2715
rect 4734 2681 4742 2691
rect 4742 2681 4768 2691
rect 4807 2681 4811 2691
rect 4811 2681 4841 2691
rect 4880 2681 4914 2715
rect 4953 2691 4987 2715
rect 4953 2681 4984 2691
rect 4984 2681 4987 2691
rect 5026 2681 5053 2715
rect 5053 2681 5060 2715
rect 5099 2681 5133 2715
rect 5172 2681 5206 2715
rect 5245 2681 5279 2715
rect 5318 2681 5352 2715
rect 5391 2681 5425 2715
rect 5464 2681 5498 2715
rect 5537 2681 5571 2715
rect 5610 2681 5644 2715
rect 5683 2681 5717 2715
rect 5756 2681 5790 2715
rect 5829 2681 5863 2715
rect 5902 2681 5936 2715
rect 5975 2681 6009 2715
rect 6048 2681 6082 2715
rect 6121 2681 6155 2715
rect 6194 2681 6228 2715
rect 6267 2681 6301 2715
rect 6340 2681 6374 2715
rect 6413 2681 6447 2715
rect 6486 2681 6520 2715
rect 6559 2681 6593 2715
rect 6632 2681 6666 2715
rect 6705 2681 6739 2715
rect 6778 2681 6812 2715
rect 6851 2681 6885 2715
rect 6924 2681 6958 2715
rect 6997 2681 7031 2715
rect 7070 2681 7104 2715
rect 7143 2681 7177 2715
rect 7216 2681 7250 2715
rect 7289 2681 7323 2715
rect 7362 2681 7396 2715
rect 7435 2681 7469 2715
rect 7508 2681 7542 2715
rect 7581 2681 7615 2715
rect 7654 2681 7688 2715
rect 7727 2681 7761 2715
rect 7800 2681 7834 2715
rect 7873 2681 7907 2715
rect 7946 2681 7980 2715
rect 8019 2681 8053 2715
rect 8092 2681 8126 2715
rect 8165 2681 8199 2715
rect 8238 2681 8272 2715
rect 8311 2681 8345 2715
rect 8384 2681 8418 2715
rect 8457 2681 8491 2715
rect 8530 2681 8564 2715
rect 8603 2681 8637 2715
rect 8676 2681 8710 2715
rect 8749 2681 8783 2715
rect 8822 2681 8856 2715
rect 8895 2681 8929 2715
rect 8968 2681 9002 2715
rect 9041 2681 9075 2715
rect 9114 2681 9148 2715
rect 9187 2681 9221 2715
rect 9260 2681 9294 2715
rect 9333 2681 9367 2715
rect 9406 2681 9440 2715
rect 9479 2681 9513 2715
rect 9552 2681 9586 2715
rect 9625 2681 9659 2715
rect 9698 2681 9732 2715
rect 9771 2681 9805 2715
rect 9844 2681 9878 2715
rect 9917 2681 9951 2715
rect 9989 2681 10023 2715
rect 10061 2681 10095 2715
rect 10133 2681 10167 2715
rect 10205 2681 10239 2715
rect 10277 2681 10311 2715
rect 10349 2681 10383 2715
rect 10421 2681 10455 2715
rect 10493 2681 10527 2715
rect 10565 2681 10599 2715
rect 10637 2681 10671 2715
rect 10709 2681 10743 2715
rect 10781 2681 10815 2715
rect 10853 2681 10887 2715
rect 10925 2681 10959 2715
rect 11967 2663 12001 2697
rect 12040 2663 12074 2697
rect 12113 2663 12147 2697
rect 12186 2663 12220 2697
rect 12259 2663 12293 2697
rect 12332 2663 12366 2697
rect 12405 2663 12439 2697
rect 12478 2663 12512 2697
rect 12551 2663 12585 2697
rect 12624 2663 12658 2697
rect 12697 2663 12731 2697
rect 12770 2663 12804 2697
rect 12843 2663 12877 2697
rect 12916 2663 12950 2697
rect 12989 2663 13023 2697
rect 13062 2663 13096 2697
rect 13135 2663 13169 2697
rect 13208 2663 13242 2697
rect 13281 2663 13315 2697
rect 13354 2663 13388 2697
rect 13427 2663 13461 2697
rect 13500 2663 13534 2697
rect 13573 2663 13607 2697
rect 13646 2663 13680 2697
rect 13719 2663 13753 2697
rect 13792 2663 13826 2697
rect 13865 2663 13899 2697
rect 13938 2663 13972 2697
rect 14011 2663 14045 2697
rect 14084 2663 14118 2697
rect 4734 2623 4768 2639
rect 4807 2623 4841 2639
rect 4734 2605 4742 2623
rect 4742 2605 4768 2623
rect 4807 2605 4811 2623
rect 4811 2605 4841 2623
rect 4880 2605 4914 2639
rect 4953 2623 4987 2639
rect 4953 2605 4984 2623
rect 4984 2605 4987 2623
rect 5026 2605 5053 2639
rect 5053 2605 5060 2639
rect 5099 2605 5133 2639
rect 5172 2605 5206 2639
rect 5245 2605 5279 2639
rect 5318 2605 5352 2639
rect 5391 2605 5425 2639
rect 5464 2605 5498 2639
rect 5537 2605 5571 2639
rect 5610 2605 5644 2639
rect 5683 2605 5717 2639
rect 5756 2605 5790 2639
rect 5829 2605 5863 2639
rect 5902 2605 5936 2639
rect 5975 2605 6009 2639
rect 6048 2605 6082 2639
rect 6121 2605 6155 2639
rect 6194 2605 6228 2639
rect 6267 2605 6301 2639
rect 6340 2605 6374 2639
rect 6413 2605 6447 2639
rect 6486 2605 6520 2639
rect 6559 2605 6593 2639
rect 6632 2605 6666 2639
rect 6705 2605 6739 2639
rect 6778 2605 6812 2639
rect 6851 2605 6885 2639
rect 6924 2605 6958 2639
rect 6997 2605 7031 2639
rect 7070 2605 7104 2639
rect 7143 2605 7177 2639
rect 7216 2605 7250 2639
rect 7289 2605 7323 2639
rect 7362 2605 7396 2639
rect 7435 2605 7469 2639
rect 7508 2605 7542 2639
rect 7581 2605 7615 2639
rect 7654 2605 7688 2639
rect 7727 2605 7761 2639
rect 7800 2605 7834 2639
rect 7873 2605 7907 2639
rect 7946 2605 7980 2639
rect 8019 2605 8053 2639
rect 8092 2605 8126 2639
rect 8165 2605 8199 2639
rect 8238 2605 8272 2639
rect 8311 2605 8345 2639
rect 8384 2605 8418 2639
rect 8457 2605 8491 2639
rect 8530 2605 8564 2639
rect 8603 2605 8637 2639
rect 8676 2605 8710 2639
rect 8749 2605 8783 2639
rect 8822 2605 8856 2639
rect 8895 2605 8929 2639
rect 8968 2605 9002 2639
rect 9041 2605 9075 2639
rect 9114 2605 9148 2639
rect 9187 2605 9221 2639
rect 9260 2605 9294 2639
rect 9333 2605 9367 2639
rect 9406 2605 9440 2639
rect 9479 2605 9513 2639
rect 9552 2605 9586 2639
rect 9625 2605 9659 2639
rect 9698 2605 9732 2639
rect 9771 2605 9805 2639
rect 9844 2605 9878 2639
rect 9917 2605 9951 2639
rect 9989 2605 10023 2639
rect 10061 2605 10095 2639
rect 10133 2605 10167 2639
rect 10205 2605 10239 2639
rect 10277 2605 10311 2639
rect 10349 2605 10383 2639
rect 10421 2605 10455 2639
rect 10493 2605 10527 2639
rect 10565 2605 10599 2639
rect 10637 2605 10671 2639
rect 10709 2605 10743 2639
rect 10781 2605 10815 2639
rect 10853 2605 10887 2639
rect 10925 2605 10959 2639
rect 11967 2591 12001 2625
rect 12040 2591 12074 2625
rect 12113 2591 12147 2625
rect 12186 2591 12220 2625
rect 12259 2591 12293 2625
rect 12332 2591 12366 2625
rect 12405 2591 12439 2625
rect 12478 2591 12512 2625
rect 12551 2591 12585 2625
rect 12624 2591 12658 2625
rect 12697 2591 12731 2625
rect 12770 2591 12804 2625
rect 12843 2591 12877 2625
rect 12916 2591 12950 2625
rect 12989 2591 13023 2625
rect 13062 2591 13096 2625
rect 13135 2591 13169 2625
rect 13208 2591 13242 2625
rect 13281 2591 13315 2625
rect 13354 2591 13388 2625
rect 13427 2591 13461 2625
rect 13500 2591 13534 2625
rect 13573 2591 13607 2625
rect 13646 2591 13680 2625
rect 13719 2591 13753 2625
rect 13792 2591 13826 2625
rect 13865 2591 13899 2625
rect 13938 2591 13972 2625
rect 14011 2591 14045 2625
rect 14084 2591 14118 2625
rect 4734 2555 4768 2563
rect 4807 2555 4841 2563
rect 4734 2529 4742 2555
rect 4742 2529 4768 2555
rect 4807 2529 4811 2555
rect 4811 2529 4841 2555
rect 4880 2529 4914 2563
rect 4953 2555 4987 2563
rect 4953 2529 4984 2555
rect 4984 2529 4987 2555
rect 5026 2529 5053 2563
rect 5053 2529 5060 2563
rect 5099 2529 5133 2563
rect 5172 2529 5206 2563
rect 5245 2529 5279 2563
rect 5318 2529 5352 2563
rect 5391 2529 5425 2563
rect 5464 2529 5498 2563
rect 5537 2529 5571 2563
rect 5610 2529 5644 2563
rect 5683 2529 5717 2563
rect 5756 2529 5790 2563
rect 5829 2529 5863 2563
rect 5902 2529 5936 2563
rect 5975 2529 6009 2563
rect 6048 2529 6082 2563
rect 6121 2529 6155 2563
rect 6194 2529 6228 2563
rect 6267 2529 6301 2563
rect 6340 2529 6374 2563
rect 6413 2529 6447 2563
rect 6486 2529 6520 2563
rect 6559 2529 6593 2563
rect 6632 2529 6666 2563
rect 6705 2529 6739 2563
rect 6778 2529 6812 2563
rect 6851 2529 6885 2563
rect 6924 2529 6958 2563
rect 6997 2529 7031 2563
rect 7070 2529 7104 2563
rect 7143 2529 7177 2563
rect 7216 2529 7250 2563
rect 7289 2529 7323 2563
rect 7362 2529 7396 2563
rect 7435 2529 7469 2563
rect 7508 2529 7542 2563
rect 7581 2529 7615 2563
rect 7654 2529 7688 2563
rect 7727 2529 7761 2563
rect 7800 2529 7834 2563
rect 7873 2529 7907 2563
rect 7946 2529 7980 2563
rect 8019 2529 8053 2563
rect 8092 2529 8126 2563
rect 8165 2529 8199 2563
rect 8238 2529 8272 2563
rect 8311 2529 8345 2563
rect 8384 2529 8418 2563
rect 8457 2529 8491 2563
rect 8530 2529 8564 2563
rect 8603 2529 8637 2563
rect 8676 2529 8710 2563
rect 8749 2529 8783 2563
rect 8822 2529 8856 2563
rect 8895 2529 8929 2563
rect 8968 2529 9002 2563
rect 9041 2529 9075 2563
rect 9114 2529 9148 2563
rect 9187 2529 9221 2563
rect 9260 2529 9294 2563
rect 9333 2529 9367 2563
rect 9406 2529 9440 2563
rect 9479 2529 9513 2563
rect 9552 2529 9586 2563
rect 9625 2529 9659 2563
rect 9698 2529 9732 2563
rect 9771 2529 9805 2563
rect 9844 2529 9878 2563
rect 9917 2529 9951 2563
rect 9989 2529 10023 2563
rect 10061 2529 10095 2563
rect 10133 2529 10167 2563
rect 10205 2529 10239 2563
rect 10277 2529 10311 2563
rect 10349 2529 10383 2563
rect 10421 2529 10455 2563
rect 10493 2529 10527 2563
rect 10565 2529 10599 2563
rect 10637 2529 10671 2563
rect 10709 2529 10743 2563
rect 10781 2529 10815 2563
rect 10853 2529 10887 2563
rect 10925 2529 10959 2563
rect 11967 2519 12001 2553
rect 12040 2519 12074 2553
rect 12113 2519 12147 2553
rect 12186 2519 12220 2553
rect 12259 2519 12293 2553
rect 12332 2519 12366 2553
rect 12405 2519 12439 2553
rect 12478 2519 12512 2553
rect 12551 2519 12585 2553
rect 12624 2519 12658 2553
rect 12697 2519 12731 2553
rect 12770 2519 12804 2553
rect 12843 2519 12877 2553
rect 12916 2519 12950 2553
rect 12989 2519 13023 2553
rect 13062 2519 13096 2553
rect 13135 2519 13169 2553
rect 13208 2519 13242 2553
rect 13281 2519 13315 2553
rect 13354 2519 13388 2553
rect 13427 2519 13461 2553
rect 13500 2519 13534 2553
rect 13573 2519 13607 2553
rect 13646 2519 13680 2553
rect 13719 2519 13753 2553
rect 13792 2519 13826 2553
rect 13865 2519 13899 2553
rect 13938 2519 13972 2553
rect 14011 2519 14045 2553
rect 14084 2519 14118 2553
rect 4734 2453 4742 2487
rect 4742 2453 4768 2487
rect 4807 2453 4811 2487
rect 4811 2453 4841 2487
rect 4880 2453 4914 2487
rect 4953 2453 4984 2487
rect 4984 2453 4987 2487
rect 5026 2453 5053 2487
rect 5053 2453 5060 2487
rect 5099 2453 5133 2487
rect 5172 2453 5206 2487
rect 5245 2453 5279 2487
rect 5318 2453 5352 2487
rect 5391 2453 5425 2487
rect 5464 2453 5498 2487
rect 5537 2453 5571 2487
rect 5610 2453 5644 2487
rect 5683 2453 5717 2487
rect 5756 2453 5790 2487
rect 5829 2453 5863 2487
rect 5902 2453 5936 2487
rect 5975 2453 6009 2487
rect 6048 2453 6082 2487
rect 6121 2453 6155 2487
rect 6194 2453 6228 2487
rect 6267 2453 6301 2487
rect 6340 2453 6374 2487
rect 6413 2453 6447 2487
rect 6486 2453 6520 2487
rect 6559 2453 6593 2487
rect 6632 2453 6666 2487
rect 6705 2453 6739 2487
rect 6778 2453 6812 2487
rect 6851 2453 6885 2487
rect 6924 2453 6958 2487
rect 6997 2453 7031 2487
rect 7070 2453 7104 2487
rect 7143 2453 7177 2487
rect 7216 2453 7250 2487
rect 7289 2453 7323 2487
rect 7362 2453 7396 2487
rect 7435 2453 7469 2487
rect 7508 2453 7542 2487
rect 7581 2453 7615 2487
rect 7654 2453 7688 2487
rect 7727 2453 7761 2487
rect 7800 2453 7834 2487
rect 7873 2453 7907 2487
rect 7946 2453 7980 2487
rect 8019 2453 8053 2487
rect 8092 2453 8126 2487
rect 8165 2453 8199 2487
rect 8238 2453 8272 2487
rect 8311 2453 8345 2487
rect 8384 2453 8418 2487
rect 8457 2453 8491 2487
rect 8530 2453 8564 2487
rect 8603 2453 8637 2487
rect 8676 2453 8710 2487
rect 8749 2453 8783 2487
rect 8822 2453 8856 2487
rect 8895 2453 8929 2487
rect 8968 2453 9002 2487
rect 9041 2453 9075 2487
rect 9114 2453 9148 2487
rect 9187 2453 9221 2487
rect 9260 2453 9294 2487
rect 9333 2453 9367 2487
rect 9406 2453 9440 2487
rect 9479 2453 9513 2487
rect 9552 2453 9586 2487
rect 9625 2453 9659 2487
rect 9698 2453 9732 2487
rect 9771 2453 9805 2487
rect 9844 2453 9878 2487
rect 9917 2453 9951 2487
rect 9989 2453 10023 2487
rect 10061 2453 10095 2487
rect 10133 2453 10167 2487
rect 10205 2453 10239 2487
rect 10277 2453 10311 2487
rect 10349 2453 10383 2487
rect 10421 2453 10455 2487
rect 10493 2453 10527 2487
rect 10565 2453 10599 2487
rect 10637 2453 10671 2487
rect 10709 2453 10743 2487
rect 10781 2453 10815 2487
rect 10853 2453 10887 2487
rect 10925 2453 10959 2487
rect 11967 2447 12001 2481
rect 12040 2447 12074 2481
rect 12113 2447 12147 2481
rect 12186 2447 12220 2481
rect 12259 2447 12293 2481
rect 12332 2447 12366 2481
rect 12405 2447 12439 2481
rect 12478 2447 12512 2481
rect 12551 2447 12585 2481
rect 12624 2447 12658 2481
rect 12697 2447 12731 2481
rect 12770 2447 12804 2481
rect 12843 2447 12877 2481
rect 12916 2447 12950 2481
rect 12989 2447 13023 2481
rect 13062 2447 13096 2481
rect 13135 2447 13169 2481
rect 13208 2447 13242 2481
rect 13281 2447 13315 2481
rect 13354 2447 13388 2481
rect 13427 2447 13461 2481
rect 13500 2447 13534 2481
rect 13573 2447 13607 2481
rect 13646 2447 13680 2481
rect 13719 2447 13753 2481
rect 13792 2447 13826 2481
rect 13865 2447 13899 2481
rect 13938 2447 13972 2481
rect 14011 2447 14045 2481
rect 14084 2447 14118 2481
rect 4734 2385 4742 2411
rect 4742 2385 4768 2411
rect 4807 2385 4811 2411
rect 4811 2385 4841 2411
rect 4734 2377 4768 2385
rect 4807 2377 4841 2385
rect 4880 2377 4914 2411
rect 4953 2385 4984 2411
rect 4984 2385 4987 2411
rect 4953 2377 4987 2385
rect 5026 2377 5053 2411
rect 5053 2377 5060 2411
rect 5099 2377 5133 2411
rect 5172 2377 5206 2411
rect 5245 2377 5279 2411
rect 5318 2377 5352 2411
rect 5391 2377 5425 2411
rect 5464 2377 5498 2411
rect 5537 2377 5571 2411
rect 5610 2377 5644 2411
rect 5683 2377 5717 2411
rect 5756 2377 5790 2411
rect 5829 2377 5863 2411
rect 5902 2377 5936 2411
rect 5975 2377 6009 2411
rect 6048 2377 6082 2411
rect 6121 2377 6155 2411
rect 6194 2377 6228 2411
rect 6267 2377 6301 2411
rect 6340 2377 6374 2411
rect 6413 2377 6447 2411
rect 6486 2377 6520 2411
rect 6559 2377 6593 2411
rect 6632 2377 6666 2411
rect 6705 2377 6739 2411
rect 6778 2377 6812 2411
rect 6851 2377 6885 2411
rect 6924 2377 6958 2411
rect 6997 2377 7031 2411
rect 7070 2377 7104 2411
rect 7143 2377 7177 2411
rect 7216 2377 7250 2411
rect 7289 2377 7323 2411
rect 7362 2377 7396 2411
rect 7435 2377 7469 2411
rect 7508 2377 7542 2411
rect 7581 2377 7615 2411
rect 7654 2377 7688 2411
rect 7727 2377 7761 2411
rect 7800 2377 7834 2411
rect 7873 2377 7907 2411
rect 7946 2377 7980 2411
rect 8019 2377 8053 2411
rect 8092 2377 8126 2411
rect 8165 2377 8199 2411
rect 8238 2377 8272 2411
rect 8311 2377 8345 2411
rect 8384 2377 8418 2411
rect 8457 2377 8491 2411
rect 8530 2377 8564 2411
rect 8603 2377 8637 2411
rect 8676 2377 8710 2411
rect 8749 2377 8783 2411
rect 8822 2377 8856 2411
rect 8895 2377 8929 2411
rect 8968 2377 9002 2411
rect 9041 2377 9075 2411
rect 9114 2377 9148 2411
rect 9187 2377 9221 2411
rect 9260 2377 9294 2411
rect 9333 2377 9367 2411
rect 9406 2377 9440 2411
rect 9479 2377 9513 2411
rect 9552 2377 9586 2411
rect 9625 2377 9659 2411
rect 9698 2377 9732 2411
rect 9771 2377 9805 2411
rect 9844 2377 9878 2411
rect 9917 2377 9951 2411
rect 9989 2377 10023 2411
rect 10061 2377 10095 2411
rect 10133 2377 10167 2411
rect 10205 2377 10239 2411
rect 10277 2377 10311 2411
rect 10349 2377 10383 2411
rect 10421 2377 10455 2411
rect 10493 2377 10527 2411
rect 10565 2377 10599 2411
rect 10637 2377 10671 2411
rect 10709 2377 10743 2411
rect 10781 2377 10815 2411
rect 10853 2377 10887 2411
rect 10925 2377 10959 2411
rect 11967 2375 12001 2409
rect 12040 2375 12074 2409
rect 12113 2375 12147 2409
rect 12186 2375 12220 2409
rect 12259 2375 12293 2409
rect 12332 2375 12366 2409
rect 12405 2375 12439 2409
rect 12478 2375 12512 2409
rect 12551 2375 12585 2409
rect 12624 2375 12658 2409
rect 12697 2375 12731 2409
rect 12770 2375 12804 2409
rect 12843 2375 12877 2409
rect 12916 2375 12950 2409
rect 12989 2375 13023 2409
rect 13062 2375 13096 2409
rect 13135 2375 13169 2409
rect 13208 2375 13242 2409
rect 13281 2375 13315 2409
rect 13354 2375 13388 2409
rect 13427 2375 13461 2409
rect 13500 2375 13534 2409
rect 13573 2375 13607 2409
rect 13646 2375 13680 2409
rect 13719 2375 13753 2409
rect 13792 2375 13826 2409
rect 13865 2375 13899 2409
rect 13938 2375 13972 2409
rect 14011 2375 14045 2409
rect 14084 2375 14118 2409
rect 4734 2317 4742 2335
rect 4742 2317 4768 2335
rect 4807 2317 4811 2335
rect 4811 2317 4841 2335
rect 4734 2301 4768 2317
rect 4807 2301 4841 2317
rect 4880 2301 4914 2335
rect 4953 2317 4984 2335
rect 4984 2317 4987 2335
rect 4953 2301 4987 2317
rect 5026 2301 5053 2335
rect 5053 2301 5060 2335
rect 5099 2301 5133 2335
rect 5172 2301 5206 2335
rect 5245 2301 5279 2335
rect 5318 2301 5352 2335
rect 5391 2301 5425 2335
rect 5464 2301 5498 2335
rect 5537 2301 5571 2335
rect 5610 2301 5644 2335
rect 5683 2301 5717 2335
rect 5756 2301 5790 2335
rect 5829 2301 5863 2335
rect 5902 2301 5936 2335
rect 5975 2301 6009 2335
rect 6048 2301 6082 2335
rect 6121 2301 6155 2335
rect 6194 2301 6228 2335
rect 6267 2301 6301 2335
rect 6340 2301 6374 2335
rect 6413 2301 6447 2335
rect 6486 2301 6520 2335
rect 6559 2301 6593 2335
rect 6632 2301 6666 2335
rect 6705 2301 6739 2335
rect 6778 2301 6812 2335
rect 6851 2301 6885 2335
rect 6924 2301 6958 2335
rect 6997 2301 7031 2335
rect 7070 2301 7104 2335
rect 7143 2301 7177 2335
rect 7216 2301 7250 2335
rect 7289 2301 7323 2335
rect 7362 2301 7396 2335
rect 7435 2301 7469 2335
rect 7508 2301 7542 2335
rect 7581 2301 7615 2335
rect 7654 2301 7688 2335
rect 7727 2301 7761 2335
rect 7800 2301 7834 2335
rect 7873 2301 7907 2335
rect 7946 2301 7980 2335
rect 8019 2301 8053 2335
rect 8092 2301 8126 2335
rect 8165 2301 8199 2335
rect 8238 2301 8272 2335
rect 8311 2301 8345 2335
rect 8384 2301 8418 2335
rect 8457 2301 8491 2335
rect 8530 2301 8564 2335
rect 8603 2301 8637 2335
rect 8676 2301 8710 2335
rect 8749 2301 8783 2335
rect 8822 2301 8856 2335
rect 8895 2301 8929 2335
rect 8968 2301 9002 2335
rect 9041 2301 9075 2335
rect 9114 2301 9148 2335
rect 9187 2301 9221 2335
rect 9260 2301 9294 2335
rect 9333 2301 9367 2335
rect 9406 2301 9440 2335
rect 9479 2301 9513 2335
rect 9552 2301 9586 2335
rect 9625 2301 9659 2335
rect 9698 2301 9732 2335
rect 9771 2301 9805 2335
rect 9844 2301 9878 2335
rect 9917 2301 9951 2335
rect 9989 2301 10023 2335
rect 10061 2301 10095 2335
rect 10133 2301 10167 2335
rect 10205 2301 10239 2335
rect 10277 2301 10311 2335
rect 10349 2301 10383 2335
rect 10421 2301 10455 2335
rect 10493 2301 10527 2335
rect 10565 2301 10599 2335
rect 10637 2301 10671 2335
rect 10709 2301 10743 2335
rect 10781 2301 10815 2335
rect 10853 2301 10887 2335
rect 10925 2301 10959 2335
rect 11967 2303 12001 2337
rect 12040 2303 12074 2337
rect 12113 2303 12147 2337
rect 12186 2303 12220 2337
rect 12259 2303 12293 2337
rect 12332 2303 12366 2337
rect 12405 2303 12439 2337
rect 12478 2303 12512 2337
rect 12551 2303 12585 2337
rect 12624 2303 12658 2337
rect 12697 2303 12731 2337
rect 12770 2303 12804 2337
rect 12843 2303 12877 2337
rect 12916 2303 12950 2337
rect 12989 2303 13023 2337
rect 13062 2303 13096 2337
rect 13135 2303 13169 2337
rect 13208 2303 13242 2337
rect 13281 2303 13315 2337
rect 13354 2303 13388 2337
rect 13427 2303 13461 2337
rect 13500 2303 13534 2337
rect 13573 2303 13607 2337
rect 13646 2303 13680 2337
rect 13719 2303 13753 2337
rect 13792 2303 13826 2337
rect 13865 2303 13899 2337
rect 13938 2303 13972 2337
rect 14011 2303 14045 2337
rect 14084 2303 14118 2337
rect 4734 2249 4742 2259
rect 4742 2249 4768 2259
rect 4807 2249 4811 2259
rect 4811 2249 4841 2259
rect 4734 2225 4768 2249
rect 4807 2225 4841 2249
rect 4880 2225 4914 2259
rect 4953 2249 4984 2259
rect 4984 2249 4987 2259
rect 4953 2225 4987 2249
rect 5026 2225 5053 2259
rect 5053 2225 5060 2259
rect 5099 2225 5133 2259
rect 5172 2225 5206 2259
rect 5245 2225 5279 2259
rect 5318 2225 5352 2259
rect 5391 2225 5425 2259
rect 5464 2225 5498 2259
rect 5537 2225 5571 2259
rect 5610 2225 5644 2259
rect 5683 2225 5717 2259
rect 5756 2225 5790 2259
rect 5829 2225 5863 2259
rect 5902 2225 5936 2259
rect 5975 2225 6009 2259
rect 6048 2225 6082 2259
rect 6121 2225 6155 2259
rect 6194 2225 6228 2259
rect 6267 2225 6301 2259
rect 6340 2225 6374 2259
rect 6413 2225 6447 2259
rect 6486 2225 6520 2259
rect 6559 2225 6593 2259
rect 6632 2225 6666 2259
rect 6705 2225 6739 2259
rect 6778 2225 6812 2259
rect 6851 2225 6885 2259
rect 6924 2225 6958 2259
rect 6997 2225 7031 2259
rect 7070 2225 7104 2259
rect 7143 2225 7177 2259
rect 7216 2225 7250 2259
rect 7289 2225 7323 2259
rect 7362 2225 7396 2259
rect 7435 2225 7469 2259
rect 7508 2225 7542 2259
rect 7581 2225 7615 2259
rect 7654 2225 7688 2259
rect 7727 2225 7761 2259
rect 7800 2225 7834 2259
rect 7873 2225 7907 2259
rect 7946 2225 7980 2259
rect 8019 2225 8053 2259
rect 8092 2225 8126 2259
rect 8165 2225 8199 2259
rect 8238 2225 8272 2259
rect 8311 2225 8345 2259
rect 8384 2225 8418 2259
rect 8457 2225 8491 2259
rect 8530 2225 8564 2259
rect 8603 2225 8637 2259
rect 8676 2225 8710 2259
rect 8749 2225 8783 2259
rect 8822 2225 8856 2259
rect 8895 2225 8929 2259
rect 8968 2225 9002 2259
rect 9041 2225 9075 2259
rect 9114 2225 9148 2259
rect 9187 2225 9221 2259
rect 9260 2225 9294 2259
rect 9333 2225 9367 2259
rect 9406 2225 9440 2259
rect 9479 2225 9513 2259
rect 9552 2225 9586 2259
rect 9625 2225 9659 2259
rect 9698 2225 9732 2259
rect 9771 2225 9805 2259
rect 9844 2225 9878 2259
rect 9917 2225 9951 2259
rect 9989 2225 10023 2259
rect 10061 2225 10095 2259
rect 10133 2225 10167 2259
rect 10205 2225 10239 2259
rect 10277 2225 10311 2259
rect 10349 2225 10383 2259
rect 10421 2225 10455 2259
rect 10493 2225 10527 2259
rect 10565 2225 10599 2259
rect 10637 2225 10671 2259
rect 10709 2225 10743 2259
rect 10781 2225 10815 2259
rect 10853 2225 10887 2259
rect 10925 2225 10959 2259
rect 11967 2231 12001 2265
rect 12040 2231 12074 2265
rect 12113 2231 12147 2265
rect 12186 2231 12220 2265
rect 12259 2231 12293 2265
rect 12332 2231 12366 2265
rect 12405 2231 12439 2265
rect 12478 2231 12512 2265
rect 12551 2231 12585 2265
rect 12624 2231 12658 2265
rect 12697 2231 12731 2265
rect 12770 2231 12804 2265
rect 12843 2231 12877 2265
rect 12916 2231 12950 2265
rect 12989 2231 13023 2265
rect 13062 2231 13096 2265
rect 13135 2231 13169 2265
rect 13208 2231 13242 2265
rect 13281 2231 13315 2265
rect 13354 2231 13388 2265
rect 13427 2231 13461 2265
rect 13500 2231 13534 2265
rect 13573 2231 13607 2265
rect 13646 2231 13680 2265
rect 13719 2231 13753 2265
rect 13792 2231 13826 2265
rect 13865 2231 13899 2265
rect 13938 2231 13972 2265
rect 14011 2231 14045 2265
rect 14084 2231 14118 2265
rect 4734 2181 4742 2183
rect 4742 2181 4768 2183
rect 4807 2181 4811 2183
rect 4811 2181 4841 2183
rect 4734 2149 4768 2181
rect 4807 2149 4841 2181
rect 4880 2149 4914 2183
rect 4953 2181 4984 2183
rect 4984 2181 4987 2183
rect 5026 2181 5053 2183
rect 5053 2181 5060 2183
rect 5099 2181 5133 2183
rect 5172 2181 5206 2183
rect 5245 2181 5279 2183
rect 5318 2181 5352 2183
rect 5391 2181 5425 2183
rect 5464 2181 5498 2183
rect 5537 2181 5571 2183
rect 5610 2181 5644 2183
rect 5683 2181 5717 2183
rect 5756 2181 5790 2183
rect 5829 2181 5863 2183
rect 5902 2181 5936 2183
rect 5975 2181 6009 2183
rect 6048 2181 6082 2183
rect 6121 2181 6155 2183
rect 6194 2181 6228 2183
rect 6267 2181 6301 2183
rect 6340 2181 6374 2183
rect 6413 2181 6447 2183
rect 6486 2181 6520 2183
rect 6559 2181 6593 2183
rect 6632 2181 6666 2183
rect 6705 2181 6739 2183
rect 6778 2181 6812 2183
rect 6851 2181 6885 2183
rect 6924 2181 6958 2183
rect 6997 2181 7031 2183
rect 7070 2181 7104 2183
rect 7143 2181 7177 2183
rect 7216 2181 7250 2183
rect 7289 2181 7323 2183
rect 7362 2181 7396 2183
rect 7435 2181 7469 2183
rect 7508 2181 7542 2183
rect 7581 2181 7615 2183
rect 7654 2181 7688 2183
rect 7727 2181 7761 2183
rect 7800 2181 7834 2183
rect 7873 2181 7907 2183
rect 7946 2181 7980 2183
rect 8019 2181 8053 2183
rect 8092 2181 8126 2183
rect 8165 2181 8199 2183
rect 8238 2181 8272 2183
rect 8311 2181 8345 2183
rect 8384 2181 8418 2183
rect 8457 2181 8491 2183
rect 8530 2181 8564 2183
rect 8603 2181 8637 2183
rect 8676 2181 8710 2183
rect 8749 2181 8783 2183
rect 8822 2181 8856 2183
rect 8895 2181 8929 2183
rect 8968 2181 9002 2183
rect 9041 2181 9075 2183
rect 9114 2181 9148 2183
rect 9187 2181 9221 2183
rect 9260 2181 9294 2183
rect 9333 2181 9367 2183
rect 9406 2181 9440 2183
rect 9479 2181 9513 2183
rect 9552 2181 9586 2183
rect 9625 2181 9659 2183
rect 9698 2181 9732 2183
rect 9771 2181 9805 2183
rect 9844 2181 9878 2183
rect 9917 2181 9951 2183
rect 9989 2181 10023 2183
rect 10061 2181 10095 2183
rect 10133 2181 10167 2183
rect 10205 2181 10239 2183
rect 10277 2181 10311 2183
rect 10349 2181 10383 2183
rect 10421 2181 10455 2183
rect 10493 2181 10527 2183
rect 10565 2181 10599 2183
rect 10637 2181 10671 2183
rect 10709 2181 10743 2183
rect 10781 2181 10815 2183
rect 10853 2181 10887 2183
rect 10925 2181 10959 2183
rect 11967 2181 12001 2193
rect 12040 2181 12074 2193
rect 12113 2181 12147 2193
rect 12186 2181 12220 2193
rect 12259 2181 12293 2193
rect 12332 2181 12366 2193
rect 12405 2181 12439 2193
rect 12478 2181 12512 2193
rect 12551 2181 12585 2193
rect 12624 2181 12658 2193
rect 12697 2181 12731 2193
rect 12770 2181 12804 2193
rect 12843 2181 12877 2193
rect 12916 2181 12950 2193
rect 12989 2181 13023 2193
rect 13062 2181 13096 2193
rect 13135 2181 13169 2193
rect 13208 2181 13242 2193
rect 13281 2181 13315 2193
rect 13354 2181 13388 2193
rect 13427 2181 13461 2193
rect 13500 2181 13534 2193
rect 13573 2181 13607 2193
rect 13646 2181 13680 2193
rect 13719 2181 13753 2193
rect 13792 2181 13826 2193
rect 13865 2181 13899 2193
rect 13938 2181 13972 2193
rect 14011 2181 14045 2193
rect 14084 2181 14118 2193
rect 14157 2181 16927 2697
rect 4953 2149 4987 2181
rect 5026 2149 5060 2181
rect 5099 2149 5133 2181
rect 5172 2149 5206 2181
rect 5245 2149 5279 2181
rect 5318 2149 5352 2181
rect 5391 2149 5425 2181
rect 5464 2149 5498 2181
rect 5537 2149 5571 2181
rect 5610 2149 5644 2181
rect 5683 2149 5717 2181
rect 5756 2149 5790 2181
rect 5829 2149 5863 2181
rect 5902 2149 5936 2181
rect 5975 2149 6009 2181
rect 6048 2149 6082 2181
rect 6121 2149 6155 2181
rect 6194 2149 6228 2181
rect 6267 2149 6301 2181
rect 6340 2149 6374 2181
rect 6413 2149 6447 2181
rect 6486 2149 6520 2181
rect 6559 2149 6593 2181
rect 6632 2149 6666 2181
rect 6705 2149 6739 2181
rect 6778 2149 6812 2181
rect 6851 2149 6885 2181
rect 6924 2149 6958 2181
rect 6997 2149 7031 2181
rect 7070 2149 7104 2181
rect 7143 2149 7177 2181
rect 7216 2149 7250 2181
rect 7289 2149 7323 2181
rect 7362 2149 7396 2181
rect 7435 2149 7469 2181
rect 7508 2149 7542 2181
rect 7581 2149 7615 2181
rect 7654 2149 7688 2181
rect 7727 2149 7761 2181
rect 7800 2149 7834 2181
rect 7873 2149 7907 2181
rect 7946 2149 7980 2181
rect 8019 2149 8053 2181
rect 8092 2149 8126 2181
rect 8165 2149 8199 2181
rect 8238 2149 8272 2181
rect 8311 2149 8345 2181
rect 8384 2149 8418 2181
rect 8457 2149 8491 2181
rect 8530 2149 8564 2181
rect 8603 2149 8637 2181
rect 8676 2149 8710 2181
rect 8749 2149 8783 2181
rect 8822 2149 8856 2181
rect 8895 2149 8929 2181
rect 8968 2149 9002 2181
rect 9041 2149 9075 2181
rect 9114 2149 9148 2181
rect 9187 2149 9221 2181
rect 9260 2149 9294 2181
rect 9333 2149 9367 2181
rect 9406 2149 9440 2181
rect 9479 2149 9513 2181
rect 9552 2149 9586 2181
rect 9625 2149 9659 2181
rect 9698 2149 9732 2181
rect 9771 2149 9805 2181
rect 9844 2149 9878 2181
rect 9917 2149 9951 2181
rect 9989 2149 10023 2181
rect 10061 2149 10095 2181
rect 10133 2149 10167 2181
rect 10205 2149 10239 2181
rect 10277 2149 10311 2181
rect 10349 2149 10383 2181
rect 10421 2149 10455 2181
rect 10493 2149 10527 2181
rect 10565 2149 10599 2181
rect 10637 2149 10671 2181
rect 10709 2149 10743 2181
rect 10781 2149 10815 2181
rect 10853 2149 10887 2181
rect 10925 2149 10959 2181
rect 11967 2159 12001 2181
rect 12040 2159 12074 2181
rect 12113 2159 12147 2181
rect 12186 2159 12220 2181
rect 12259 2159 12293 2181
rect 12332 2159 12366 2181
rect 12405 2159 12439 2181
rect 12478 2159 12512 2181
rect 12551 2159 12585 2181
rect 12624 2159 12658 2181
rect 12697 2159 12731 2181
rect 12770 2159 12804 2181
rect 12843 2159 12877 2181
rect 12916 2159 12950 2181
rect 12989 2159 13023 2181
rect 13062 2159 13096 2181
rect 13135 2159 13169 2181
rect 13208 2159 13242 2181
rect 13281 2159 13315 2181
rect 13354 2159 13388 2181
rect 13427 2159 13461 2181
rect 13500 2159 13534 2181
rect 13573 2159 13607 2181
rect 13646 2159 13680 2181
rect 13719 2159 13753 2181
rect 13792 2159 13826 2181
rect 13865 2159 13899 2181
rect 13938 2159 13972 2181
rect 14011 2159 14045 2181
rect 14084 2159 14118 2181
rect 14157 2159 15944 2181
rect 15944 2159 16726 2181
rect 16726 2159 16927 2181
rect 4616 1846 4650 1858
rect 4688 1846 4722 1858
rect 4760 1846 4794 1858
rect 4832 1846 4866 1858
rect 4904 1846 4938 1858
rect 4976 1846 5010 1858
rect 5048 1846 5082 1858
rect 5120 1846 5154 1858
rect 5192 1846 5226 1858
rect 5264 1846 5298 1858
rect 5336 1846 5370 1858
rect 5408 1846 5442 1858
rect 5480 1846 5514 1858
rect 5552 1846 5586 1858
rect 5624 1846 5658 1858
rect 5696 1846 5730 1858
rect -2832 1812 -2825 1841
rect -2825 1812 -2798 1841
rect -2759 1812 -2756 1841
rect -2756 1812 -2725 1841
rect -2832 1807 -2798 1812
rect -2759 1807 -2725 1812
rect -2686 1807 -2652 1841
rect -2613 1812 -2583 1841
rect -2583 1812 -2579 1841
rect -2540 1812 -2514 1841
rect -2514 1812 -2506 1841
rect -2467 1812 -2445 1841
rect -2445 1812 -2433 1841
rect -2394 1812 -2376 1841
rect -2376 1812 -2360 1841
rect -2321 1812 -2307 1841
rect -2307 1812 -2287 1841
rect -2248 1812 -2238 1841
rect -2238 1812 -2214 1841
rect -2175 1812 -2169 1841
rect -2169 1812 -2141 1841
rect -2102 1812 -2100 1841
rect -2100 1812 -2068 1841
rect -2029 1812 -1997 1841
rect -1997 1812 -1995 1841
rect -1956 1812 -1928 1841
rect -1928 1812 -1922 1841
rect -1883 1812 -1859 1841
rect -1859 1812 -1849 1841
rect -1810 1812 -1790 1841
rect -1790 1812 -1776 1841
rect -1737 1812 -1721 1841
rect -1721 1812 -1686 1841
rect -1686 1812 -1652 1841
rect -1652 1812 -1617 1841
rect -1617 1812 -1583 1841
rect -1583 1812 -1548 1841
rect -1548 1812 -1514 1841
rect -1514 1812 -1479 1841
rect -1479 1812 -1445 1841
rect -1445 1812 -1410 1841
rect -1410 1812 -1376 1841
rect -1376 1812 -1341 1841
rect -1341 1812 -1307 1841
rect -1307 1812 -1272 1841
rect -1272 1812 -1238 1841
rect -1238 1812 -1203 1841
rect -1203 1812 -1169 1841
rect -1169 1812 -1134 1841
rect -1134 1812 -1100 1841
rect -1100 1812 -1065 1841
rect -1065 1812 -1031 1841
rect -1031 1812 -996 1841
rect -996 1812 -962 1841
rect -962 1812 -927 1841
rect -927 1812 -893 1841
rect -893 1812 -858 1841
rect -858 1812 -824 1841
rect -824 1812 -789 1841
rect -789 1812 -755 1841
rect -755 1812 -720 1841
rect -720 1812 -686 1841
rect -686 1812 -651 1841
rect -651 1812 -617 1841
rect -617 1812 -582 1841
rect -582 1812 -548 1841
rect -548 1812 -513 1841
rect -513 1812 -479 1841
rect -479 1812 -444 1841
rect -444 1812 -410 1841
rect -410 1812 -375 1841
rect -2613 1807 -2579 1812
rect -2540 1807 -2506 1812
rect -2467 1807 -2433 1812
rect -2394 1807 -2360 1812
rect -2321 1807 -2287 1812
rect -2248 1807 -2214 1812
rect -2175 1807 -2141 1812
rect -2102 1807 -2068 1812
rect -2029 1807 -1995 1812
rect -1956 1807 -1922 1812
rect -1883 1807 -1849 1812
rect -1810 1807 -1776 1812
rect -1737 1778 -375 1812
rect -2832 1744 -2825 1769
rect -2825 1744 -2798 1769
rect -2759 1744 -2756 1769
rect -2756 1744 -2725 1769
rect -2832 1735 -2798 1744
rect -2759 1735 -2725 1744
rect -2686 1735 -2652 1769
rect -2613 1744 -2583 1769
rect -2583 1744 -2579 1769
rect -2540 1744 -2514 1769
rect -2514 1744 -2506 1769
rect -2467 1744 -2445 1769
rect -2445 1744 -2433 1769
rect -2394 1744 -2376 1769
rect -2376 1744 -2360 1769
rect -2321 1744 -2307 1769
rect -2307 1744 -2287 1769
rect -2248 1744 -2238 1769
rect -2238 1744 -2214 1769
rect -2175 1744 -2169 1769
rect -2169 1744 -2141 1769
rect -2102 1744 -2100 1769
rect -2100 1744 -2068 1769
rect -2029 1744 -1997 1769
rect -1997 1744 -1995 1769
rect -1956 1744 -1928 1769
rect -1928 1744 -1922 1769
rect -1883 1744 -1859 1769
rect -1859 1744 -1849 1769
rect -1810 1744 -1790 1769
rect -1790 1744 -1776 1769
rect -1737 1744 -1721 1778
rect -1721 1744 -1686 1778
rect -1686 1744 -1652 1778
rect -1652 1744 -1617 1778
rect -1617 1744 -1583 1778
rect -1583 1744 -1548 1778
rect -1548 1744 -1514 1778
rect -1514 1744 -1479 1778
rect -1479 1744 -1445 1778
rect -1445 1744 -1410 1778
rect -1410 1744 -1376 1778
rect -1376 1744 -1341 1778
rect -1341 1744 -1307 1778
rect -1307 1744 -1272 1778
rect -1272 1744 -1238 1778
rect -1238 1744 -1203 1778
rect -1203 1744 -1169 1778
rect -1169 1744 -1134 1778
rect -1134 1744 -1100 1778
rect -1100 1744 -1065 1778
rect -1065 1744 -1031 1778
rect -1031 1744 -996 1778
rect -996 1744 -962 1778
rect -962 1744 -927 1778
rect -927 1744 -893 1778
rect -893 1744 -858 1778
rect -858 1744 -824 1778
rect -824 1744 -789 1778
rect -789 1744 -755 1778
rect -755 1744 -720 1778
rect -720 1744 -686 1778
rect -686 1744 -651 1778
rect -651 1744 -617 1778
rect -617 1744 -582 1778
rect -582 1744 -548 1778
rect -548 1744 -513 1778
rect -513 1744 -479 1778
rect -479 1744 -444 1778
rect -444 1744 -410 1778
rect -410 1744 -375 1778
rect -2613 1735 -2579 1744
rect -2540 1735 -2506 1744
rect -2467 1735 -2433 1744
rect -2394 1735 -2360 1744
rect -2321 1735 -2287 1744
rect -2248 1735 -2214 1744
rect -2175 1735 -2141 1744
rect -2102 1735 -2068 1744
rect -2029 1735 -1995 1744
rect -1956 1735 -1922 1744
rect -1883 1735 -1849 1744
rect -1810 1735 -1776 1744
rect -1737 1710 -375 1744
rect -2832 1676 -2825 1697
rect -2825 1676 -2798 1697
rect -2759 1676 -2756 1697
rect -2756 1676 -2725 1697
rect -2832 1663 -2798 1676
rect -2759 1663 -2725 1676
rect -2686 1663 -2652 1697
rect -2613 1676 -2583 1697
rect -2583 1676 -2579 1697
rect -2540 1676 -2514 1697
rect -2514 1676 -2506 1697
rect -2467 1676 -2445 1697
rect -2445 1676 -2433 1697
rect -2394 1676 -2376 1697
rect -2376 1676 -2360 1697
rect -2321 1676 -2307 1697
rect -2307 1676 -2287 1697
rect -2248 1676 -2238 1697
rect -2238 1676 -2214 1697
rect -2175 1676 -2169 1697
rect -2169 1676 -2141 1697
rect -2102 1676 -2100 1697
rect -2100 1676 -2068 1697
rect -2029 1676 -1997 1697
rect -1997 1676 -1995 1697
rect -1956 1676 -1928 1697
rect -1928 1676 -1922 1697
rect -1883 1676 -1859 1697
rect -1859 1676 -1849 1697
rect -1810 1676 -1790 1697
rect -1790 1676 -1776 1697
rect -1737 1676 -1721 1710
rect -1721 1676 -1686 1710
rect -1686 1676 -1652 1710
rect -1652 1676 -1617 1710
rect -1617 1676 -1583 1710
rect -1583 1676 -1548 1710
rect -1548 1676 -1514 1710
rect -1514 1676 -1479 1710
rect -1479 1676 -1445 1710
rect -1445 1676 -1410 1710
rect -1410 1676 -1376 1710
rect -1376 1676 -1341 1710
rect -1341 1676 -1307 1710
rect -1307 1676 -1272 1710
rect -1272 1676 -1238 1710
rect -1238 1676 -1203 1710
rect -1203 1676 -1169 1710
rect -1169 1676 -1134 1710
rect -1134 1676 -1100 1710
rect -1100 1676 -1065 1710
rect -1065 1676 -1031 1710
rect -1031 1676 -996 1710
rect -996 1676 -962 1710
rect -962 1676 -927 1710
rect -927 1676 -893 1710
rect -893 1676 -858 1710
rect -858 1676 -824 1710
rect -824 1676 -789 1710
rect -789 1676 -755 1710
rect -755 1676 -720 1710
rect -720 1676 -686 1710
rect -686 1676 -651 1710
rect -651 1676 -617 1710
rect -617 1676 -582 1710
rect -582 1676 -548 1710
rect -548 1676 -513 1710
rect -513 1676 -479 1710
rect -479 1676 -444 1710
rect -444 1676 -410 1710
rect -410 1676 -375 1710
rect -2613 1663 -2579 1676
rect -2540 1663 -2506 1676
rect -2467 1663 -2433 1676
rect -2394 1663 -2360 1676
rect -2321 1663 -2287 1676
rect -2248 1663 -2214 1676
rect -2175 1663 -2141 1676
rect -2102 1663 -2068 1676
rect -2029 1663 -1995 1676
rect -1956 1663 -1922 1676
rect -1883 1663 -1849 1676
rect -1810 1663 -1776 1676
rect -1737 1642 -375 1676
rect -2832 1608 -2825 1625
rect -2825 1608 -2798 1625
rect -2759 1608 -2756 1625
rect -2756 1608 -2725 1625
rect -2832 1591 -2798 1608
rect -2759 1591 -2725 1608
rect -2686 1591 -2652 1625
rect -2613 1608 -2583 1625
rect -2583 1608 -2579 1625
rect -2540 1608 -2514 1625
rect -2514 1608 -2506 1625
rect -2467 1608 -2445 1625
rect -2445 1608 -2433 1625
rect -2394 1608 -2376 1625
rect -2376 1608 -2360 1625
rect -2321 1608 -2307 1625
rect -2307 1608 -2287 1625
rect -2248 1608 -2238 1625
rect -2238 1608 -2214 1625
rect -2175 1608 -2169 1625
rect -2169 1608 -2141 1625
rect -2102 1608 -2100 1625
rect -2100 1608 -2068 1625
rect -2029 1608 -1997 1625
rect -1997 1608 -1995 1625
rect -1956 1608 -1928 1625
rect -1928 1608 -1922 1625
rect -1883 1608 -1859 1625
rect -1859 1608 -1849 1625
rect -1810 1608 -1790 1625
rect -1790 1608 -1776 1625
rect -1737 1608 -1721 1642
rect -1721 1608 -1686 1642
rect -1686 1608 -1652 1642
rect -1652 1608 -1617 1642
rect -1617 1608 -1583 1642
rect -1583 1608 -1548 1642
rect -1548 1608 -1514 1642
rect -1514 1608 -1479 1642
rect -1479 1608 -1445 1642
rect -1445 1608 -1410 1642
rect -1410 1608 -1376 1642
rect -1376 1608 -1341 1642
rect -1341 1608 -1307 1642
rect -1307 1608 -1272 1642
rect -1272 1608 -1238 1642
rect -1238 1608 -1203 1642
rect -1203 1608 -1169 1642
rect -1169 1608 -1134 1642
rect -1134 1608 -1100 1642
rect -1100 1608 -1065 1642
rect -1065 1608 -1031 1642
rect -1031 1608 -996 1642
rect -996 1608 -962 1642
rect -962 1608 -927 1642
rect -927 1608 -893 1642
rect -893 1608 -858 1642
rect -858 1608 -824 1642
rect -824 1608 -789 1642
rect -789 1608 -755 1642
rect -755 1608 -720 1642
rect -720 1608 -686 1642
rect -686 1608 -651 1642
rect -651 1608 -617 1642
rect -617 1608 -582 1642
rect -582 1608 -548 1642
rect -548 1608 -513 1642
rect -513 1608 -479 1642
rect -479 1608 -444 1642
rect -444 1608 -410 1642
rect -410 1608 -375 1642
rect -2613 1591 -2579 1608
rect -2540 1591 -2506 1608
rect -2467 1591 -2433 1608
rect -2394 1591 -2360 1608
rect -2321 1591 -2287 1608
rect -2248 1591 -2214 1608
rect -2175 1591 -2141 1608
rect -2102 1591 -2068 1608
rect -2029 1591 -1995 1608
rect -1956 1591 -1922 1608
rect -1883 1591 -1849 1608
rect -1810 1591 -1776 1608
rect -1737 1574 -375 1608
rect -2832 1540 -2825 1553
rect -2825 1540 -2798 1553
rect -2759 1540 -2756 1553
rect -2756 1540 -2725 1553
rect -2832 1519 -2798 1540
rect -2759 1519 -2725 1540
rect -2686 1519 -2652 1553
rect -2613 1540 -2583 1553
rect -2583 1540 -2579 1553
rect -2540 1540 -2514 1553
rect -2514 1540 -2506 1553
rect -2467 1540 -2445 1553
rect -2445 1540 -2433 1553
rect -2394 1540 -2376 1553
rect -2376 1540 -2360 1553
rect -2321 1540 -2307 1553
rect -2307 1540 -2287 1553
rect -2248 1540 -2238 1553
rect -2238 1540 -2214 1553
rect -2175 1540 -2169 1553
rect -2169 1540 -2141 1553
rect -2102 1540 -2100 1553
rect -2100 1540 -2068 1553
rect -2029 1540 -1997 1553
rect -1997 1540 -1995 1553
rect -1956 1540 -1928 1553
rect -1928 1540 -1922 1553
rect -1883 1540 -1859 1553
rect -1859 1540 -1849 1553
rect -1810 1540 -1790 1553
rect -1790 1540 -1776 1553
rect -1737 1540 -1721 1574
rect -1721 1540 -1686 1574
rect -1686 1540 -1652 1574
rect -1652 1540 -1617 1574
rect -1617 1540 -1583 1574
rect -1583 1540 -1548 1574
rect -1548 1540 -1514 1574
rect -1514 1540 -1479 1574
rect -1479 1540 -1445 1574
rect -1445 1540 -1410 1574
rect -1410 1540 -1376 1574
rect -1376 1540 -1341 1574
rect -1341 1540 -1307 1574
rect -1307 1540 -1272 1574
rect -1272 1540 -1238 1574
rect -1238 1540 -1203 1574
rect -1203 1540 -1169 1574
rect -1169 1540 -1134 1574
rect -1134 1540 -1100 1574
rect -1100 1540 -1065 1574
rect -1065 1540 -1031 1574
rect -1031 1540 -996 1574
rect -996 1540 -962 1574
rect -962 1540 -927 1574
rect -927 1540 -893 1574
rect -893 1540 -858 1574
rect -858 1540 -824 1574
rect -824 1540 -789 1574
rect -789 1540 -755 1574
rect -755 1540 -720 1574
rect -720 1540 -686 1574
rect -686 1540 -651 1574
rect -651 1540 -617 1574
rect -617 1540 -582 1574
rect -582 1540 -548 1574
rect -548 1540 -513 1574
rect -513 1540 -479 1574
rect -479 1540 -444 1574
rect -444 1540 -410 1574
rect -410 1540 -375 1574
rect -2613 1519 -2579 1540
rect -2540 1519 -2506 1540
rect -2467 1519 -2433 1540
rect -2394 1519 -2360 1540
rect -2321 1519 -2287 1540
rect -2248 1519 -2214 1540
rect -2175 1519 -2141 1540
rect -2102 1519 -2068 1540
rect -2029 1519 -1995 1540
rect -1956 1519 -1922 1540
rect -1883 1519 -1849 1540
rect -1810 1519 -1776 1540
rect -1737 1506 -375 1540
rect -2832 1472 -2825 1481
rect -2825 1472 -2798 1481
rect -2759 1472 -2756 1481
rect -2756 1472 -2725 1481
rect -2832 1447 -2798 1472
rect -2759 1447 -2725 1472
rect -2686 1447 -2652 1481
rect -2613 1472 -2583 1481
rect -2583 1472 -2579 1481
rect -2540 1472 -2514 1481
rect -2514 1472 -2506 1481
rect -2467 1472 -2445 1481
rect -2445 1472 -2433 1481
rect -2394 1472 -2376 1481
rect -2376 1472 -2360 1481
rect -2321 1472 -2307 1481
rect -2307 1472 -2287 1481
rect -2248 1472 -2238 1481
rect -2238 1472 -2214 1481
rect -2175 1472 -2169 1481
rect -2169 1472 -2141 1481
rect -2102 1472 -2100 1481
rect -2100 1472 -2068 1481
rect -2029 1472 -1997 1481
rect -1997 1472 -1995 1481
rect -1956 1472 -1928 1481
rect -1928 1472 -1922 1481
rect -1883 1472 -1859 1481
rect -1859 1472 -1849 1481
rect -1810 1472 -1790 1481
rect -1790 1472 -1776 1481
rect -1737 1472 -1721 1506
rect -1721 1472 -1686 1506
rect -1686 1472 -1652 1506
rect -1652 1472 -1617 1506
rect -1617 1472 -1583 1506
rect -1583 1472 -1548 1506
rect -1548 1472 -1514 1506
rect -1514 1472 -1479 1506
rect -1479 1472 -1445 1506
rect -1445 1472 -1410 1506
rect -1410 1472 -1376 1506
rect -1376 1472 -1341 1506
rect -1341 1472 -1307 1506
rect -1307 1472 -1272 1506
rect -1272 1472 -1238 1506
rect -1238 1472 -1203 1506
rect -1203 1472 -1169 1506
rect -1169 1472 -1134 1506
rect -1134 1472 -1100 1506
rect -1100 1472 -1065 1506
rect -1065 1472 -1031 1506
rect -1031 1472 -996 1506
rect -996 1472 -962 1506
rect -962 1472 -927 1506
rect -927 1472 -893 1506
rect -893 1472 -858 1506
rect -858 1472 -824 1506
rect -824 1472 -789 1506
rect -789 1472 -755 1506
rect -755 1472 -720 1506
rect -720 1472 -686 1506
rect -686 1472 -651 1506
rect -651 1472 -617 1506
rect -617 1472 -582 1506
rect -582 1472 -548 1506
rect -548 1472 -513 1506
rect -513 1472 -479 1506
rect -479 1472 -444 1506
rect -444 1472 -410 1506
rect -410 1472 -375 1506
rect -2613 1447 -2579 1472
rect -2540 1447 -2506 1472
rect -2467 1447 -2433 1472
rect -2394 1447 -2360 1472
rect -2321 1447 -2287 1472
rect -2248 1447 -2214 1472
rect -2175 1447 -2141 1472
rect -2102 1447 -2068 1472
rect -2029 1447 -1995 1472
rect -1956 1447 -1922 1472
rect -1883 1447 -1849 1472
rect -1810 1447 -1776 1472
rect -1737 1438 -375 1472
rect -2832 1404 -2825 1409
rect -2825 1404 -2798 1409
rect -2759 1404 -2756 1409
rect -2756 1404 -2725 1409
rect -2832 1375 -2798 1404
rect -2759 1375 -2725 1404
rect -2686 1375 -2652 1409
rect -2613 1404 -2583 1409
rect -2583 1404 -2579 1409
rect -2540 1404 -2514 1409
rect -2514 1404 -2506 1409
rect -2467 1404 -2445 1409
rect -2445 1404 -2433 1409
rect -2394 1404 -2376 1409
rect -2376 1404 -2360 1409
rect -2321 1404 -2307 1409
rect -2307 1404 -2287 1409
rect -2248 1404 -2238 1409
rect -2238 1404 -2214 1409
rect -2175 1404 -2169 1409
rect -2169 1404 -2141 1409
rect -2102 1404 -2100 1409
rect -2100 1404 -2068 1409
rect -2029 1404 -1997 1409
rect -1997 1404 -1995 1409
rect -1956 1404 -1928 1409
rect -1928 1404 -1922 1409
rect -1883 1404 -1859 1409
rect -1859 1404 -1849 1409
rect -1810 1404 -1790 1409
rect -1790 1404 -1776 1409
rect -1737 1404 -1721 1438
rect -1721 1404 -1686 1438
rect -1686 1404 -1652 1438
rect -1652 1404 -1617 1438
rect -1617 1404 -1583 1438
rect -1583 1404 -1548 1438
rect -1548 1404 -1514 1438
rect -1514 1404 -1479 1438
rect -1479 1404 -1445 1438
rect -1445 1404 -1410 1438
rect -1410 1404 -1376 1438
rect -1376 1404 -1341 1438
rect -1341 1404 -1307 1438
rect -1307 1404 -1272 1438
rect -1272 1404 -1238 1438
rect -1238 1404 -1203 1438
rect -1203 1404 -1169 1438
rect -1169 1404 -1134 1438
rect -1134 1404 -1100 1438
rect -1100 1404 -1065 1438
rect -1065 1404 -1031 1438
rect -1031 1404 -996 1438
rect -996 1404 -962 1438
rect -962 1404 -927 1438
rect -927 1404 -893 1438
rect -893 1404 -858 1438
rect -858 1404 -824 1438
rect -824 1404 -789 1438
rect -789 1404 -755 1438
rect -755 1404 -720 1438
rect -720 1404 -686 1438
rect -686 1404 -651 1438
rect -651 1404 -617 1438
rect -617 1404 -582 1438
rect -582 1404 -548 1438
rect -548 1404 -513 1438
rect -513 1404 -479 1438
rect -479 1404 -444 1438
rect -444 1404 -410 1438
rect -410 1404 -375 1438
rect -2613 1375 -2579 1404
rect -2540 1375 -2506 1404
rect -2467 1375 -2433 1404
rect -2394 1375 -2360 1404
rect -2321 1375 -2287 1404
rect -2248 1375 -2214 1404
rect -2175 1375 -2141 1404
rect -2102 1375 -2068 1404
rect -2029 1375 -1995 1404
rect -1956 1375 -1922 1404
rect -1883 1375 -1849 1404
rect -1810 1375 -1776 1404
rect -1737 1370 -375 1404
rect -2832 1336 -2825 1337
rect -2825 1336 -2798 1337
rect -2759 1336 -2756 1337
rect -2756 1336 -2725 1337
rect -2832 1303 -2798 1336
rect -2759 1303 -2725 1336
rect -2686 1303 -2652 1337
rect -2613 1336 -2583 1337
rect -2583 1336 -2579 1337
rect -2540 1336 -2514 1337
rect -2514 1336 -2506 1337
rect -2467 1336 -2445 1337
rect -2445 1336 -2433 1337
rect -2394 1336 -2376 1337
rect -2376 1336 -2360 1337
rect -2321 1336 -2307 1337
rect -2307 1336 -2287 1337
rect -2248 1336 -2238 1337
rect -2238 1336 -2214 1337
rect -2175 1336 -2169 1337
rect -2169 1336 -2141 1337
rect -2102 1336 -2100 1337
rect -2100 1336 -2068 1337
rect -2029 1336 -1997 1337
rect -1997 1336 -1995 1337
rect -1956 1336 -1928 1337
rect -1928 1336 -1922 1337
rect -1883 1336 -1859 1337
rect -1859 1336 -1849 1337
rect -1810 1336 -1790 1337
rect -1790 1336 -1776 1337
rect -1737 1336 -1721 1370
rect -1721 1336 -1686 1370
rect -1686 1336 -1652 1370
rect -1652 1336 -1617 1370
rect -1617 1336 -1583 1370
rect -1583 1336 -1548 1370
rect -1548 1336 -1514 1370
rect -1514 1336 -1479 1370
rect -1479 1336 -1445 1370
rect -1445 1336 -1410 1370
rect -1410 1336 -1376 1370
rect -1376 1336 -1341 1370
rect -1341 1336 -1307 1370
rect -1307 1336 -1272 1370
rect -1272 1336 -1238 1370
rect -1238 1336 -1203 1370
rect -1203 1336 -1169 1370
rect -1169 1336 -1134 1370
rect -1134 1336 -1100 1370
rect -1100 1336 -1065 1370
rect -1065 1336 -1031 1370
rect -1031 1336 -996 1370
rect -996 1336 -962 1370
rect -962 1336 -927 1370
rect -927 1336 -893 1370
rect -893 1336 -858 1370
rect -858 1336 -824 1370
rect -824 1336 -789 1370
rect -789 1336 -755 1370
rect -755 1336 -720 1370
rect -720 1336 -686 1370
rect -686 1336 -651 1370
rect -651 1336 -617 1370
rect -617 1336 -582 1370
rect -582 1336 -548 1370
rect -548 1336 -513 1370
rect -513 1336 -479 1370
rect -479 1336 -444 1370
rect -444 1336 -410 1370
rect -410 1336 -375 1370
rect -2613 1303 -2579 1336
rect -2540 1303 -2506 1336
rect -2467 1303 -2433 1336
rect -2394 1303 -2360 1336
rect -2321 1303 -2287 1336
rect -2248 1303 -2214 1336
rect -2175 1303 -2141 1336
rect -2102 1303 -2068 1336
rect -2029 1303 -1995 1336
rect -1956 1303 -1922 1336
rect -1883 1303 -1849 1336
rect -1810 1303 -1776 1336
rect -1737 1302 -375 1336
rect -1737 1268 -1721 1302
rect -1721 1268 -1686 1302
rect -1686 1268 -1652 1302
rect -1652 1268 -1617 1302
rect -1617 1268 -1583 1302
rect -1583 1268 -1548 1302
rect -1548 1268 -1514 1302
rect -1514 1268 -1479 1302
rect -1479 1268 -1445 1302
rect -1445 1268 -1410 1302
rect -1410 1268 -1376 1302
rect -1376 1268 -1341 1302
rect -1341 1268 -1307 1302
rect -1307 1268 -1272 1302
rect -1272 1268 -1238 1302
rect -1238 1268 -1203 1302
rect -1203 1268 -1169 1302
rect -1169 1268 -1134 1302
rect -1134 1268 -1100 1302
rect -1100 1268 -1065 1302
rect -1065 1268 -1031 1302
rect -1031 1268 -996 1302
rect -996 1268 -962 1302
rect -962 1268 -927 1302
rect -927 1268 -893 1302
rect -893 1268 -858 1302
rect -858 1268 -824 1302
rect -824 1268 -789 1302
rect -789 1268 -755 1302
rect -755 1268 -720 1302
rect -720 1268 -686 1302
rect -686 1268 -651 1302
rect -651 1268 -617 1302
rect -617 1268 -582 1302
rect -582 1268 -548 1302
rect -548 1268 -513 1302
rect -513 1268 -479 1302
rect -479 1268 -444 1302
rect -444 1268 -410 1302
rect -410 1268 -375 1302
rect -2832 1234 -2798 1265
rect -2759 1234 -2725 1265
rect -2832 1231 -2825 1234
rect -2825 1231 -2798 1234
rect -2759 1231 -2756 1234
rect -2756 1231 -2725 1234
rect -2686 1231 -2652 1265
rect -2613 1234 -2579 1265
rect -2540 1234 -2506 1265
rect -2467 1234 -2433 1265
rect -2394 1234 -2360 1265
rect -2321 1234 -2287 1265
rect -2248 1234 -2214 1265
rect -2175 1234 -2141 1265
rect -2102 1234 -2068 1265
rect -2029 1234 -1995 1265
rect -1956 1234 -1922 1265
rect -1883 1234 -1849 1265
rect -1810 1234 -1776 1265
rect -1737 1234 -375 1268
rect -2613 1231 -2583 1234
rect -2583 1231 -2579 1234
rect -2540 1231 -2514 1234
rect -2514 1231 -2506 1234
rect -2467 1231 -2445 1234
rect -2445 1231 -2433 1234
rect -2394 1231 -2376 1234
rect -2376 1231 -2360 1234
rect -2321 1231 -2307 1234
rect -2307 1231 -2287 1234
rect -2248 1231 -2238 1234
rect -2238 1231 -2214 1234
rect -2175 1231 -2169 1234
rect -2169 1231 -2141 1234
rect -2102 1231 -2100 1234
rect -2100 1231 -2068 1234
rect -2029 1231 -1997 1234
rect -1997 1231 -1995 1234
rect -1956 1231 -1928 1234
rect -1928 1231 -1922 1234
rect -1883 1231 -1859 1234
rect -1859 1231 -1849 1234
rect -1810 1231 -1790 1234
rect -1790 1231 -1776 1234
rect -1737 1231 -1721 1234
rect -1721 1231 -1686 1234
rect -1686 1231 -1652 1234
rect -1652 1231 -1617 1234
rect -1617 1231 -1583 1234
rect -1583 1231 -1548 1234
rect -1548 1231 -1514 1234
rect -1514 1231 -1479 1234
rect -1479 1231 -1445 1234
rect -1445 1231 -1410 1234
rect -1410 1231 -1376 1234
rect -1376 1231 -1341 1234
rect -1341 1231 -1307 1234
rect -1307 1231 -1272 1234
rect -1272 1231 -1238 1234
rect -1238 1231 -1203 1234
rect -1203 1231 -1169 1234
rect -1169 1231 -1134 1234
rect -1134 1231 -1100 1234
rect -1100 1231 -1065 1234
rect -1065 1231 -1031 1234
rect -1031 1231 -996 1234
rect -996 1231 -962 1234
rect -962 1231 -927 1234
rect -927 1231 -893 1234
rect -893 1231 -858 1234
rect -858 1231 -824 1234
rect -824 1231 -789 1234
rect -789 1231 -755 1234
rect -755 1231 -720 1234
rect -720 1231 -686 1234
rect -686 1231 -651 1234
rect -651 1231 -617 1234
rect -617 1231 -582 1234
rect -582 1231 -548 1234
rect -548 1231 -513 1234
rect -513 1231 -479 1234
rect -479 1231 -444 1234
rect -444 1231 -410 1234
rect -410 1231 -375 1234
rect -375 1231 -1 1841
rect -1 1231 33 1841
rect 33 1231 4561 1841
rect 4616 1824 4650 1846
rect 4688 1824 4722 1846
rect 4760 1824 4794 1846
rect 4832 1824 4866 1846
rect 4904 1824 4938 1846
rect 4976 1824 5010 1846
rect 5048 1824 5082 1846
rect 5120 1824 5154 1846
rect 5192 1824 5226 1846
rect 5264 1824 5298 1846
rect 5336 1824 5370 1846
rect 5408 1824 5442 1846
rect 5480 1824 5514 1846
rect 5552 1824 5586 1846
rect 5624 1824 5658 1846
rect 5696 1824 5711 1846
rect 5711 1824 5730 1846
rect 5768 1824 5802 1858
rect 5840 1824 5874 1858
rect 5912 1824 5946 1858
rect 5984 1824 6018 1858
rect 6056 1824 6090 1858
rect 6128 1824 6162 1858
rect 6200 1824 6234 1858
rect 6272 1824 6306 1858
rect 6344 1824 6378 1858
rect 6416 1824 6450 1858
rect 6488 1824 6522 1858
rect 6560 1824 6594 1858
rect 6632 1824 6666 1858
rect 6704 1824 6738 1858
rect 6776 1824 6810 1858
rect 6848 1824 6882 1858
rect 6920 1824 6954 1858
rect 6992 1824 7026 1858
rect 7064 1824 7098 1858
rect 7136 1824 7170 1858
rect 7208 1824 7242 1858
rect 7280 1824 7314 1858
rect 7352 1824 7386 1858
rect 7424 1824 7458 1858
rect 7496 1824 7530 1858
rect 7568 1824 7602 1858
rect 7640 1824 7674 1858
rect 7712 1824 7746 1858
rect 7784 1824 7818 1858
rect 7856 1824 7890 1858
rect 7928 1824 7962 1858
rect 8000 1824 8034 1858
rect 8072 1824 8106 1858
rect 8144 1824 8178 1858
rect 8216 1824 8250 1858
rect 8288 1824 8322 1858
rect 8360 1824 8394 1858
rect 8432 1824 8466 1858
rect 8504 1824 8538 1858
rect 8576 1824 8610 1858
rect 8648 1824 8682 1858
rect 8720 1824 8754 1858
rect 8792 1824 8826 1858
rect 8864 1824 8898 1858
rect 8936 1824 8970 1858
rect 9008 1824 9042 1858
rect 9080 1824 9114 1858
rect 9152 1824 9186 1858
rect 9224 1824 9258 1858
rect 9296 1824 9330 1858
rect 9368 1824 9402 1858
rect 9440 1824 9474 1858
rect 9512 1824 9546 1858
rect 9584 1824 9618 1858
rect 9656 1824 9690 1858
rect 9728 1824 9762 1858
rect 9800 1824 9834 1858
rect 9872 1824 9906 1858
rect 9944 1824 9978 1858
rect 10016 1824 10050 1858
rect 10088 1824 10122 1858
rect 10160 1824 10194 1858
rect 10232 1824 10266 1858
rect 10304 1824 10338 1858
rect 10376 1824 10410 1858
rect 10448 1824 10482 1858
rect 10520 1824 10554 1858
rect 10592 1824 10626 1858
rect 10664 1824 10698 1858
rect 10736 1824 10770 1858
rect 10808 1824 10842 1858
rect 10880 1824 10914 1858
rect 10952 1824 10986 1858
rect 11024 1824 11058 1858
rect 11096 1824 11130 1858
rect 11168 1824 11202 1858
rect 11240 1824 11274 1858
rect 11312 1824 11346 1858
rect 11384 1824 11418 1858
rect 11456 1824 11490 1858
rect 11528 1824 11562 1858
rect 11600 1824 11634 1858
rect 11672 1824 11706 1858
rect 11744 1824 11778 1858
rect 11816 1824 11850 1858
rect 11888 1824 11922 1858
rect 11960 1824 11994 1858
rect 12032 1824 12066 1858
rect 12104 1824 12138 1858
rect 12176 1824 12210 1858
rect 12248 1824 12282 1858
rect 12320 1824 12354 1858
rect 12392 1824 12426 1858
rect 12464 1824 12498 1858
rect 12536 1824 12570 1858
rect 12608 1824 12642 1858
rect 12680 1824 12714 1858
rect 12752 1824 12786 1858
rect 12824 1824 12858 1858
rect 12896 1824 12930 1858
rect 12968 1824 13002 1858
rect 13040 1824 13074 1858
rect 13112 1824 13146 1858
rect 13184 1824 13218 1858
rect 13256 1824 13290 1858
rect 13328 1824 13362 1858
rect 13400 1824 13434 1858
rect 13472 1824 13506 1858
rect 13544 1824 13578 1858
rect 13616 1824 13650 1858
rect 13688 1824 13722 1858
rect 13760 1824 13794 1858
rect 13832 1824 13866 1858
rect 13904 1824 13938 1858
rect 13976 1824 14010 1858
rect 14048 1824 14082 1858
rect 14120 1824 14154 1858
rect 14192 1824 14226 1858
rect 14264 1824 14298 1858
rect 14336 1824 14370 1858
rect 14408 1824 14442 1858
rect 14480 1824 14514 1858
rect 14552 1824 14586 1858
rect 14624 1824 14658 1858
rect 14696 1824 14730 1858
rect 14768 1824 14802 1858
rect 14840 1824 14874 1858
rect 14912 1824 14946 1858
rect 14984 1824 15018 1858
rect 15056 1824 15090 1858
rect 15128 1824 15162 1858
rect 15200 1824 15234 1858
rect 15272 1824 15306 1858
rect 15344 1824 15378 1858
rect 15416 1824 15450 1858
rect 15488 1824 15522 1858
rect 15561 1824 15595 1858
rect 15634 1824 15668 1858
rect 15707 1824 15741 1858
rect 15780 1824 15814 1858
rect 15853 1824 15887 1858
rect 15926 1824 15944 1858
rect 15944 1824 15960 1858
rect 15999 1824 16033 1858
rect 16072 1824 16106 1858
rect 16145 1824 16179 1858
rect 16218 1824 16252 1858
rect 16291 1824 16325 1858
rect 16364 1824 16398 1858
rect 16437 1824 16471 1858
rect 16510 1824 16544 1858
rect 16583 1824 16617 1858
rect 16656 1824 16690 1858
rect 4616 1746 4650 1780
rect 4688 1746 4722 1780
rect 4760 1746 4794 1780
rect 4832 1746 4866 1780
rect 4904 1746 4938 1780
rect 4976 1746 5010 1780
rect 5048 1746 5082 1780
rect 5120 1746 5154 1780
rect 5192 1746 5226 1780
rect 5264 1746 5298 1780
rect 5336 1746 5370 1780
rect 5408 1746 5442 1780
rect 5480 1746 5514 1780
rect 5552 1746 5586 1780
rect 5624 1746 5658 1780
rect 5696 1746 5711 1780
rect 5711 1746 5730 1780
rect 5768 1746 5802 1780
rect 5840 1746 5874 1780
rect 5912 1746 5946 1780
rect 5984 1746 6018 1780
rect 6056 1746 6090 1780
rect 6128 1746 6162 1780
rect 6200 1746 6234 1780
rect 6272 1746 6306 1780
rect 6344 1746 6378 1780
rect 6416 1746 6450 1780
rect 6488 1746 6522 1780
rect 6560 1746 6594 1780
rect 6632 1746 6666 1780
rect 6704 1746 6738 1780
rect 6776 1746 6810 1780
rect 6848 1746 6882 1780
rect 6920 1746 6954 1780
rect 6992 1746 7026 1780
rect 7064 1746 7098 1780
rect 7136 1746 7170 1780
rect 7208 1746 7242 1780
rect 7280 1746 7314 1780
rect 7352 1746 7386 1780
rect 7424 1746 7458 1780
rect 7496 1746 7530 1780
rect 7568 1746 7602 1780
rect 7640 1746 7674 1780
rect 7712 1746 7746 1780
rect 7784 1746 7818 1780
rect 7856 1746 7890 1780
rect 7928 1746 7962 1780
rect 8000 1746 8034 1780
rect 8072 1746 8106 1780
rect 8144 1746 8178 1780
rect 8216 1746 8250 1780
rect 8288 1746 8322 1780
rect 8360 1746 8394 1780
rect 8432 1746 8466 1780
rect 8504 1746 8538 1780
rect 8576 1746 8610 1780
rect 8648 1746 8682 1780
rect 8720 1746 8754 1780
rect 8792 1746 8826 1780
rect 8864 1746 8898 1780
rect 8936 1746 8970 1780
rect 9008 1746 9042 1780
rect 9080 1746 9114 1780
rect 9152 1746 9186 1780
rect 9224 1746 9258 1780
rect 9296 1746 9330 1780
rect 9368 1746 9402 1780
rect 9440 1746 9474 1780
rect 9512 1746 9546 1780
rect 9584 1746 9618 1780
rect 9656 1746 9690 1780
rect 9728 1746 9762 1780
rect 9800 1746 9834 1780
rect 9872 1746 9906 1780
rect 9944 1746 9978 1780
rect 10016 1746 10050 1780
rect 10088 1746 10122 1780
rect 10160 1746 10194 1780
rect 10232 1746 10266 1780
rect 10304 1746 10338 1780
rect 10376 1746 10410 1780
rect 10448 1746 10482 1780
rect 10520 1746 10554 1780
rect 10592 1746 10626 1780
rect 10664 1746 10698 1780
rect 10736 1746 10770 1780
rect 10808 1746 10842 1780
rect 10880 1746 10914 1780
rect 10952 1746 10986 1780
rect 11024 1746 11058 1780
rect 11096 1746 11130 1780
rect 11168 1746 11202 1780
rect 11240 1746 11274 1780
rect 11312 1746 11346 1780
rect 11384 1746 11418 1780
rect 11456 1746 11490 1780
rect 11528 1746 11562 1780
rect 11600 1746 11634 1780
rect 11672 1746 11706 1780
rect 11744 1746 11778 1780
rect 11816 1746 11850 1780
rect 11888 1746 11922 1780
rect 11960 1746 11994 1780
rect 12032 1746 12066 1780
rect 12104 1746 12138 1780
rect 12176 1746 12210 1780
rect 12248 1746 12282 1780
rect 12320 1746 12354 1780
rect 12392 1746 12426 1780
rect 12464 1746 12498 1780
rect 12536 1746 12570 1780
rect 12608 1746 12642 1780
rect 12680 1746 12714 1780
rect 12752 1746 12786 1780
rect 12824 1746 12858 1780
rect 12896 1746 12930 1780
rect 12968 1746 13002 1780
rect 13040 1746 13074 1780
rect 13112 1746 13146 1780
rect 13184 1746 13218 1780
rect 13256 1746 13290 1780
rect 13328 1746 13362 1780
rect 13400 1746 13434 1780
rect 13472 1746 13506 1780
rect 13544 1746 13578 1780
rect 13616 1746 13650 1780
rect 13688 1746 13722 1780
rect 13760 1746 13794 1780
rect 13832 1746 13866 1780
rect 13904 1746 13938 1780
rect 13976 1746 14010 1780
rect 14048 1746 14082 1780
rect 14120 1746 14154 1780
rect 14192 1746 14226 1780
rect 14264 1746 14298 1780
rect 14336 1746 14370 1780
rect 14408 1746 14442 1780
rect 14480 1746 14514 1780
rect 14552 1746 14586 1780
rect 14624 1746 14658 1780
rect 14696 1746 14730 1780
rect 14768 1746 14802 1780
rect 14840 1746 14874 1780
rect 14912 1746 14946 1780
rect 14984 1746 15018 1780
rect 15056 1746 15090 1780
rect 15128 1746 15162 1780
rect 15200 1746 15234 1780
rect 15272 1746 15306 1780
rect 15344 1746 15378 1780
rect 15416 1746 15450 1780
rect 15488 1746 15522 1780
rect 15561 1746 15595 1780
rect 15634 1746 15668 1780
rect 15707 1746 15741 1780
rect 15780 1746 15814 1780
rect 15853 1746 15887 1780
rect 15926 1746 15944 1780
rect 15944 1746 15960 1780
rect 15999 1746 16033 1780
rect 16072 1746 16106 1780
rect 16145 1746 16179 1780
rect 16218 1746 16252 1780
rect 16291 1746 16325 1780
rect 16364 1746 16398 1780
rect 16437 1746 16471 1780
rect 16510 1746 16544 1780
rect 16583 1746 16617 1780
rect 16656 1746 16690 1780
rect 4616 1668 4650 1702
rect 4688 1668 4722 1702
rect 4760 1668 4794 1702
rect 4832 1668 4866 1702
rect 4904 1668 4938 1702
rect 4976 1668 5010 1702
rect 5048 1668 5082 1702
rect 5120 1668 5154 1702
rect 5192 1668 5226 1702
rect 5264 1668 5298 1702
rect 5336 1668 5370 1702
rect 5408 1668 5442 1702
rect 5480 1668 5514 1702
rect 5552 1668 5586 1702
rect 5624 1668 5658 1702
rect 5696 1668 5711 1702
rect 5711 1668 5730 1702
rect 5768 1668 5802 1702
rect 5840 1668 5874 1702
rect 5912 1668 5946 1702
rect 5984 1668 6018 1702
rect 6056 1668 6090 1702
rect 6128 1668 6162 1702
rect 6200 1668 6234 1702
rect 6272 1668 6306 1702
rect 6344 1668 6378 1702
rect 6416 1668 6450 1702
rect 6488 1668 6522 1702
rect 6560 1668 6594 1702
rect 6632 1668 6666 1702
rect 6704 1668 6738 1702
rect 6776 1668 6810 1702
rect 6848 1668 6882 1702
rect 6920 1668 6954 1702
rect 6992 1668 7026 1702
rect 7064 1668 7098 1702
rect 7136 1668 7170 1702
rect 7208 1668 7242 1702
rect 7280 1668 7314 1702
rect 7352 1668 7386 1702
rect 7424 1668 7458 1702
rect 7496 1668 7530 1702
rect 7568 1668 7602 1702
rect 7640 1668 7674 1702
rect 7712 1668 7746 1702
rect 7784 1668 7818 1702
rect 7856 1668 7890 1702
rect 7928 1668 7962 1702
rect 8000 1668 8034 1702
rect 8072 1668 8106 1702
rect 8144 1668 8178 1702
rect 8216 1668 8250 1702
rect 8288 1668 8322 1702
rect 8360 1668 8394 1702
rect 8432 1668 8466 1702
rect 8504 1668 8538 1702
rect 8576 1668 8610 1702
rect 8648 1668 8682 1702
rect 8720 1668 8754 1702
rect 8792 1668 8826 1702
rect 8864 1668 8898 1702
rect 8936 1668 8970 1702
rect 9008 1668 9042 1702
rect 9080 1668 9114 1702
rect 9152 1668 9186 1702
rect 9224 1668 9258 1702
rect 9296 1668 9330 1702
rect 9368 1668 9402 1702
rect 9440 1668 9474 1702
rect 9512 1668 9546 1702
rect 9584 1668 9618 1702
rect 9656 1668 9690 1702
rect 9728 1668 9762 1702
rect 9800 1668 9834 1702
rect 9872 1668 9906 1702
rect 9944 1668 9978 1702
rect 10016 1668 10050 1702
rect 10088 1668 10122 1702
rect 10160 1668 10194 1702
rect 10232 1668 10266 1702
rect 10304 1668 10338 1702
rect 10376 1668 10410 1702
rect 10448 1668 10482 1702
rect 10520 1668 10554 1702
rect 10592 1668 10626 1702
rect 10664 1668 10698 1702
rect 10736 1668 10770 1702
rect 10808 1668 10842 1702
rect 10880 1668 10914 1702
rect 10952 1668 10986 1702
rect 11024 1668 11058 1702
rect 11096 1668 11130 1702
rect 11168 1668 11202 1702
rect 11240 1668 11274 1702
rect 11312 1668 11346 1702
rect 11384 1668 11418 1702
rect 11456 1668 11490 1702
rect 11528 1668 11562 1702
rect 11600 1668 11634 1702
rect 11672 1668 11706 1702
rect 11744 1668 11778 1702
rect 11816 1668 11850 1702
rect 11888 1668 11922 1702
rect 11960 1668 11994 1702
rect 12032 1668 12066 1702
rect 12104 1668 12138 1702
rect 12176 1668 12210 1702
rect 12248 1668 12282 1702
rect 12320 1668 12354 1702
rect 12392 1668 12426 1702
rect 12464 1668 12498 1702
rect 12536 1668 12570 1702
rect 12608 1668 12642 1702
rect 12680 1668 12714 1702
rect 12752 1668 12786 1702
rect 12824 1668 12858 1702
rect 12896 1668 12930 1702
rect 12968 1668 13002 1702
rect 13040 1668 13074 1702
rect 13112 1668 13146 1702
rect 13184 1668 13218 1702
rect 13256 1668 13290 1702
rect 13328 1668 13362 1702
rect 13400 1668 13434 1702
rect 13472 1668 13506 1702
rect 13544 1668 13578 1702
rect 13616 1668 13650 1702
rect 13688 1668 13722 1702
rect 13760 1668 13794 1702
rect 13832 1668 13866 1702
rect 13904 1668 13938 1702
rect 13976 1668 14010 1702
rect 14048 1668 14082 1702
rect 14120 1668 14154 1702
rect 14192 1668 14226 1702
rect 14264 1668 14298 1702
rect 14336 1668 14370 1702
rect 14408 1668 14442 1702
rect 14480 1668 14514 1702
rect 14552 1668 14586 1702
rect 14624 1668 14658 1702
rect 14696 1668 14730 1702
rect 14768 1668 14802 1702
rect 14840 1668 14874 1702
rect 14912 1668 14946 1702
rect 14984 1668 15018 1702
rect 15056 1668 15090 1702
rect 15128 1668 15162 1702
rect 15200 1668 15234 1702
rect 15272 1668 15306 1702
rect 15344 1668 15378 1702
rect 15416 1668 15450 1702
rect 15488 1668 15522 1702
rect 15561 1668 15595 1702
rect 15634 1668 15668 1702
rect 15707 1668 15741 1702
rect 15780 1668 15814 1702
rect 15853 1668 15887 1702
rect 15926 1668 15944 1702
rect 15944 1668 15960 1702
rect 15999 1668 16033 1702
rect 16072 1668 16106 1702
rect 16145 1668 16179 1702
rect 16218 1668 16252 1702
rect 16291 1668 16325 1702
rect 16364 1668 16398 1702
rect 16437 1668 16471 1702
rect 16510 1668 16544 1702
rect 16583 1668 16617 1702
rect 16656 1668 16690 1702
rect 4616 1590 4650 1624
rect 4688 1590 4722 1624
rect 4760 1590 4794 1624
rect 4832 1590 4866 1624
rect 4904 1590 4938 1624
rect 4976 1590 5010 1624
rect 5048 1590 5082 1624
rect 5120 1590 5154 1624
rect 5192 1590 5226 1624
rect 5264 1590 5298 1624
rect 5336 1590 5370 1624
rect 5408 1590 5442 1624
rect 5480 1590 5514 1624
rect 5552 1590 5586 1624
rect 5624 1590 5658 1624
rect 5696 1590 5711 1624
rect 5711 1590 5730 1624
rect 5768 1590 5802 1624
rect 5840 1590 5874 1624
rect 5912 1590 5946 1624
rect 5984 1590 6018 1624
rect 6056 1590 6090 1624
rect 6128 1590 6162 1624
rect 6200 1590 6234 1624
rect 6272 1590 6306 1624
rect 6344 1590 6378 1624
rect 6416 1590 6450 1624
rect 6488 1590 6522 1624
rect 6560 1590 6594 1624
rect 6632 1590 6666 1624
rect 6704 1590 6738 1624
rect 6776 1590 6810 1624
rect 6848 1590 6882 1624
rect 6920 1590 6954 1624
rect 6992 1590 7026 1624
rect 7064 1590 7098 1624
rect 7136 1590 7170 1624
rect 7208 1590 7242 1624
rect 7280 1590 7314 1624
rect 7352 1590 7386 1624
rect 7424 1590 7458 1624
rect 7496 1590 7530 1624
rect 7568 1590 7602 1624
rect 7640 1590 7674 1624
rect 7712 1590 7746 1624
rect 7784 1590 7818 1624
rect 7856 1590 7890 1624
rect 7928 1590 7962 1624
rect 8000 1590 8034 1624
rect 8072 1590 8106 1624
rect 8144 1590 8178 1624
rect 8216 1590 8250 1624
rect 8288 1590 8322 1624
rect 8360 1590 8394 1624
rect 8432 1590 8466 1624
rect 8504 1590 8538 1624
rect 8576 1590 8610 1624
rect 8648 1590 8682 1624
rect 8720 1590 8754 1624
rect 8792 1590 8826 1624
rect 8864 1590 8898 1624
rect 8936 1590 8970 1624
rect 9008 1590 9042 1624
rect 9080 1590 9114 1624
rect 9152 1590 9186 1624
rect 9224 1590 9258 1624
rect 9296 1590 9330 1624
rect 9368 1590 9402 1624
rect 9440 1590 9474 1624
rect 9512 1590 9546 1624
rect 9584 1590 9618 1624
rect 9656 1590 9690 1624
rect 9728 1590 9762 1624
rect 9800 1590 9834 1624
rect 9872 1590 9906 1624
rect 9944 1590 9978 1624
rect 10016 1590 10050 1624
rect 10088 1590 10122 1624
rect 10160 1590 10194 1624
rect 10232 1590 10266 1624
rect 10304 1590 10338 1624
rect 10376 1590 10410 1624
rect 10448 1590 10482 1624
rect 10520 1590 10554 1624
rect 10592 1590 10626 1624
rect 10664 1590 10698 1624
rect 10736 1590 10770 1624
rect 10808 1590 10842 1624
rect 10880 1590 10914 1624
rect 10952 1590 10986 1624
rect 11024 1590 11058 1624
rect 11096 1590 11130 1624
rect 11168 1590 11202 1624
rect 11240 1590 11274 1624
rect 11312 1590 11346 1624
rect 11384 1590 11418 1624
rect 11456 1590 11490 1624
rect 11528 1590 11562 1624
rect 11600 1590 11634 1624
rect 11672 1590 11706 1624
rect 11744 1590 11778 1624
rect 11816 1590 11850 1624
rect 11888 1590 11922 1624
rect 11960 1590 11994 1624
rect 12032 1590 12066 1624
rect 12104 1590 12138 1624
rect 12176 1590 12210 1624
rect 12248 1590 12282 1624
rect 12320 1590 12354 1624
rect 12392 1590 12426 1624
rect 12464 1590 12498 1624
rect 12536 1590 12570 1624
rect 12608 1590 12642 1624
rect 12680 1590 12714 1624
rect 12752 1590 12786 1624
rect 12824 1590 12858 1624
rect 12896 1590 12930 1624
rect 12968 1590 13002 1624
rect 13040 1590 13074 1624
rect 13112 1590 13146 1624
rect 13184 1590 13218 1624
rect 13256 1590 13290 1624
rect 13328 1590 13362 1624
rect 13400 1590 13434 1624
rect 13472 1590 13506 1624
rect 13544 1590 13578 1624
rect 13616 1590 13650 1624
rect 13688 1590 13722 1624
rect 13760 1590 13794 1624
rect 13832 1590 13866 1624
rect 13904 1590 13938 1624
rect 13976 1590 14010 1624
rect 14048 1590 14082 1624
rect 14120 1590 14154 1624
rect 14192 1590 14226 1624
rect 14264 1590 14298 1624
rect 14336 1590 14370 1624
rect 14408 1590 14442 1624
rect 14480 1590 14514 1624
rect 14552 1590 14586 1624
rect 14624 1590 14658 1624
rect 14696 1590 14730 1624
rect 14768 1590 14802 1624
rect 14840 1590 14874 1624
rect 14912 1590 14946 1624
rect 14984 1590 15018 1624
rect 15056 1590 15090 1624
rect 15128 1590 15162 1624
rect 15200 1590 15234 1624
rect 15272 1590 15306 1624
rect 15344 1590 15378 1624
rect 15416 1590 15450 1624
rect 15488 1590 15522 1624
rect 15561 1590 15595 1624
rect 15634 1590 15668 1624
rect 15707 1590 15741 1624
rect 15780 1590 15814 1624
rect 15853 1590 15887 1624
rect 15926 1590 15944 1624
rect 15944 1590 15960 1624
rect 15999 1590 16033 1624
rect 16072 1590 16106 1624
rect 16145 1590 16179 1624
rect 16218 1590 16252 1624
rect 16291 1590 16325 1624
rect 16364 1590 16398 1624
rect 16437 1590 16471 1624
rect 16510 1590 16544 1624
rect 16583 1590 16617 1624
rect 16656 1590 16690 1624
rect 4616 1512 4650 1546
rect 4688 1512 4722 1546
rect 4760 1512 4794 1546
rect 4832 1512 4866 1546
rect 4904 1512 4938 1546
rect 4976 1512 5010 1546
rect 5048 1512 5082 1546
rect 5120 1512 5154 1546
rect 5192 1512 5226 1546
rect 5264 1512 5298 1546
rect 5336 1512 5370 1546
rect 5408 1512 5442 1546
rect 5480 1512 5514 1546
rect 5552 1512 5586 1546
rect 5624 1512 5658 1546
rect 5696 1512 5711 1546
rect 5711 1512 5730 1546
rect 5768 1512 5802 1546
rect 5840 1512 5874 1546
rect 5912 1512 5946 1546
rect 5984 1512 6018 1546
rect 6056 1512 6090 1546
rect 6128 1512 6162 1546
rect 6200 1512 6234 1546
rect 6272 1512 6306 1546
rect 6344 1512 6378 1546
rect 6416 1512 6450 1546
rect 6488 1512 6522 1546
rect 6560 1512 6594 1546
rect 6632 1512 6666 1546
rect 6704 1512 6738 1546
rect 6776 1512 6810 1546
rect 6848 1512 6882 1546
rect 6920 1512 6954 1546
rect 6992 1512 7026 1546
rect 7064 1512 7098 1546
rect 7136 1512 7170 1546
rect 7208 1512 7242 1546
rect 7280 1512 7314 1546
rect 7352 1512 7386 1546
rect 7424 1512 7458 1546
rect 7496 1512 7530 1546
rect 7568 1512 7602 1546
rect 7640 1512 7674 1546
rect 7712 1512 7746 1546
rect 7784 1512 7818 1546
rect 7856 1512 7890 1546
rect 7928 1512 7962 1546
rect 8000 1512 8034 1546
rect 8072 1512 8106 1546
rect 8144 1512 8178 1546
rect 8216 1512 8250 1546
rect 8288 1512 8322 1546
rect 8360 1512 8394 1546
rect 8432 1512 8466 1546
rect 8504 1512 8538 1546
rect 8576 1512 8610 1546
rect 8648 1512 8682 1546
rect 8720 1512 8754 1546
rect 8792 1512 8826 1546
rect 8864 1512 8898 1546
rect 8936 1512 8970 1546
rect 9008 1512 9042 1546
rect 9080 1512 9114 1546
rect 9152 1512 9186 1546
rect 9224 1512 9258 1546
rect 9296 1512 9330 1546
rect 9368 1512 9402 1546
rect 9440 1512 9474 1546
rect 9512 1512 9546 1546
rect 9584 1512 9618 1546
rect 9656 1512 9690 1546
rect 9728 1512 9762 1546
rect 9800 1512 9834 1546
rect 9872 1512 9906 1546
rect 9944 1512 9978 1546
rect 10016 1512 10050 1546
rect 10088 1512 10122 1546
rect 10160 1512 10194 1546
rect 10232 1512 10266 1546
rect 10304 1512 10338 1546
rect 10376 1512 10410 1546
rect 10448 1512 10482 1546
rect 10520 1512 10554 1546
rect 10592 1512 10626 1546
rect 10664 1512 10698 1546
rect 10736 1512 10770 1546
rect 10808 1512 10842 1546
rect 10880 1512 10914 1546
rect 10952 1512 10986 1546
rect 11024 1512 11058 1546
rect 11096 1512 11130 1546
rect 11168 1512 11202 1546
rect 11240 1512 11274 1546
rect 11312 1512 11346 1546
rect 11384 1512 11418 1546
rect 11456 1512 11490 1546
rect 11528 1512 11562 1546
rect 11600 1512 11634 1546
rect 11672 1512 11706 1546
rect 11744 1512 11778 1546
rect 11816 1512 11850 1546
rect 11888 1512 11922 1546
rect 11960 1512 11994 1546
rect 12032 1512 12066 1546
rect 12104 1512 12138 1546
rect 12176 1512 12210 1546
rect 12248 1512 12282 1546
rect 12320 1512 12354 1546
rect 12392 1512 12426 1546
rect 12464 1512 12498 1546
rect 12536 1512 12570 1546
rect 12608 1512 12642 1546
rect 12680 1512 12714 1546
rect 12752 1512 12786 1546
rect 12824 1512 12858 1546
rect 12896 1512 12930 1546
rect 12968 1512 13002 1546
rect 13040 1512 13074 1546
rect 13112 1512 13146 1546
rect 13184 1512 13218 1546
rect 13256 1512 13290 1546
rect 13328 1512 13362 1546
rect 13400 1512 13434 1546
rect 13472 1512 13506 1546
rect 13544 1512 13578 1546
rect 13616 1512 13650 1546
rect 13688 1512 13722 1546
rect 13760 1512 13794 1546
rect 13832 1512 13866 1546
rect 13904 1512 13938 1546
rect 13976 1512 14010 1546
rect 14048 1512 14082 1546
rect 14120 1512 14154 1546
rect 14192 1512 14226 1546
rect 14264 1512 14298 1546
rect 14336 1512 14370 1546
rect 14408 1512 14442 1546
rect 14480 1512 14514 1546
rect 14552 1512 14586 1546
rect 14624 1512 14658 1546
rect 14696 1512 14730 1546
rect 14768 1512 14802 1546
rect 14840 1512 14874 1546
rect 14912 1512 14946 1546
rect 14984 1512 15018 1546
rect 15056 1512 15090 1546
rect 15128 1512 15162 1546
rect 15200 1512 15234 1546
rect 15272 1512 15306 1546
rect 15344 1512 15378 1546
rect 15416 1512 15450 1546
rect 15488 1512 15522 1546
rect 15561 1512 15595 1546
rect 15634 1512 15668 1546
rect 15707 1512 15741 1546
rect 15780 1512 15814 1546
rect 15853 1512 15887 1546
rect 15926 1512 15944 1546
rect 15944 1512 15960 1546
rect 15999 1512 16033 1546
rect 16072 1512 16106 1546
rect 16145 1512 16179 1546
rect 16218 1512 16252 1546
rect 16291 1512 16325 1546
rect 16364 1512 16398 1546
rect 16437 1512 16471 1546
rect 16510 1512 16544 1546
rect 16583 1512 16617 1546
rect 16656 1512 16690 1546
rect 4616 1434 4650 1468
rect 4688 1434 4722 1468
rect 4760 1434 4794 1468
rect 4832 1434 4866 1468
rect 4904 1434 4938 1468
rect 4976 1434 5010 1468
rect 5048 1434 5082 1468
rect 5120 1434 5154 1468
rect 5192 1434 5226 1468
rect 5264 1434 5298 1468
rect 5336 1434 5370 1468
rect 5408 1434 5442 1468
rect 5480 1434 5514 1468
rect 5552 1434 5586 1468
rect 5624 1434 5658 1468
rect 5696 1434 5711 1468
rect 5711 1434 5730 1468
rect 5768 1434 5802 1468
rect 5840 1434 5874 1468
rect 5912 1434 5946 1468
rect 5984 1434 6018 1468
rect 6056 1434 6090 1468
rect 6128 1434 6162 1468
rect 6200 1434 6234 1468
rect 6272 1434 6306 1468
rect 6344 1434 6378 1468
rect 6416 1434 6450 1468
rect 6488 1434 6522 1468
rect 6560 1434 6594 1468
rect 6632 1434 6666 1468
rect 6704 1434 6738 1468
rect 6776 1434 6810 1468
rect 6848 1434 6882 1468
rect 6920 1434 6954 1468
rect 6992 1434 7026 1468
rect 7064 1434 7098 1468
rect 7136 1434 7170 1468
rect 7208 1434 7242 1468
rect 7280 1434 7314 1468
rect 7352 1434 7386 1468
rect 7424 1434 7458 1468
rect 7496 1434 7530 1468
rect 7568 1434 7602 1468
rect 7640 1434 7674 1468
rect 7712 1434 7746 1468
rect 7784 1434 7818 1468
rect 7856 1434 7890 1468
rect 7928 1434 7962 1468
rect 8000 1434 8034 1468
rect 8072 1434 8106 1468
rect 8144 1434 8178 1468
rect 8216 1434 8250 1468
rect 8288 1434 8322 1468
rect 8360 1434 8394 1468
rect 8432 1434 8466 1468
rect 8504 1434 8538 1468
rect 8576 1434 8610 1468
rect 8648 1434 8682 1468
rect 8720 1434 8754 1468
rect 8792 1434 8826 1468
rect 8864 1434 8898 1468
rect 8936 1434 8970 1468
rect 9008 1434 9042 1468
rect 9080 1434 9114 1468
rect 9152 1434 9186 1468
rect 9224 1434 9258 1468
rect 9296 1434 9330 1468
rect 9368 1434 9402 1468
rect 9440 1434 9474 1468
rect 9512 1434 9546 1468
rect 9584 1434 9618 1468
rect 9656 1434 9690 1468
rect 9728 1434 9762 1468
rect 9800 1434 9834 1468
rect 9872 1434 9906 1468
rect 9944 1434 9978 1468
rect 10016 1434 10050 1468
rect 10088 1434 10122 1468
rect 10160 1434 10194 1468
rect 10232 1434 10266 1468
rect 10304 1434 10338 1468
rect 10376 1434 10410 1468
rect 10448 1434 10482 1468
rect 10520 1434 10554 1468
rect 10592 1434 10626 1468
rect 10664 1434 10698 1468
rect 10736 1434 10770 1468
rect 10808 1434 10842 1468
rect 10880 1434 10914 1468
rect 10952 1434 10986 1468
rect 11024 1434 11058 1468
rect 11096 1434 11130 1468
rect 11168 1434 11202 1468
rect 11240 1434 11274 1468
rect 11312 1434 11346 1468
rect 11384 1434 11418 1468
rect 11456 1434 11490 1468
rect 11528 1434 11562 1468
rect 11600 1434 11634 1468
rect 11672 1434 11706 1468
rect 11744 1434 11778 1468
rect 11816 1434 11850 1468
rect 11888 1434 11922 1468
rect 11960 1434 11994 1468
rect 12032 1434 12066 1468
rect 12104 1434 12138 1468
rect 12176 1434 12210 1468
rect 12248 1434 12282 1468
rect 12320 1434 12354 1468
rect 12392 1434 12426 1468
rect 12464 1434 12498 1468
rect 12536 1434 12570 1468
rect 12608 1434 12642 1468
rect 12680 1434 12714 1468
rect 12752 1434 12786 1468
rect 12824 1434 12858 1468
rect 12896 1434 12930 1468
rect 12968 1434 13002 1468
rect 13040 1434 13074 1468
rect 13112 1434 13146 1468
rect 13184 1434 13218 1468
rect 13256 1434 13290 1468
rect 13328 1434 13362 1468
rect 13400 1434 13434 1468
rect 13472 1434 13506 1468
rect 13544 1434 13578 1468
rect 13616 1434 13650 1468
rect 13688 1434 13722 1468
rect 13760 1434 13794 1468
rect 13832 1434 13866 1468
rect 13904 1434 13938 1468
rect 13976 1434 14010 1468
rect 14048 1434 14082 1468
rect 14120 1434 14154 1468
rect 14192 1434 14226 1468
rect 14264 1434 14298 1468
rect 14336 1434 14370 1468
rect 14408 1434 14442 1468
rect 14480 1434 14514 1468
rect 14552 1434 14586 1468
rect 14624 1434 14658 1468
rect 14696 1434 14730 1468
rect 14768 1434 14802 1468
rect 14840 1434 14874 1468
rect 14912 1434 14946 1468
rect 14984 1434 15018 1468
rect 15056 1434 15090 1468
rect 15128 1434 15162 1468
rect 15200 1434 15234 1468
rect 15272 1434 15306 1468
rect 15344 1434 15378 1468
rect 15416 1434 15450 1468
rect 15488 1434 15522 1468
rect 15561 1434 15595 1468
rect 15634 1434 15668 1468
rect 15707 1434 15741 1468
rect 15780 1434 15814 1468
rect 15853 1434 15887 1468
rect 15926 1434 15944 1468
rect 15944 1434 15960 1468
rect 15999 1434 16033 1468
rect 16072 1434 16106 1468
rect 16145 1434 16179 1468
rect 16218 1434 16252 1468
rect 16291 1434 16325 1468
rect 16364 1434 16398 1468
rect 16437 1434 16471 1468
rect 16510 1434 16544 1468
rect 16583 1434 16617 1468
rect 16656 1434 16690 1468
rect 4721 1214 5259 1392
rect 5298 1358 5332 1392
rect 5371 1358 5405 1392
rect 5444 1358 5478 1392
rect 5517 1358 5551 1392
rect 5590 1358 5624 1392
rect 5663 1358 5697 1392
rect 5736 1358 5770 1392
rect 5809 1358 5843 1392
rect 5882 1358 5916 1392
rect 5298 1286 5332 1320
rect 5371 1286 5405 1320
rect 5444 1286 5478 1320
rect 5517 1286 5551 1320
rect 5590 1286 5624 1320
rect 5663 1286 5697 1320
rect 5736 1286 5770 1320
rect 5809 1286 5843 1320
rect 5882 1286 5916 1320
rect 15560 1359 15594 1393
rect 15633 1359 15667 1393
rect 15706 1359 15740 1393
rect 15779 1359 15813 1393
rect 15852 1359 15886 1393
rect 15925 1359 15944 1393
rect 15944 1359 15959 1393
rect 15998 1359 16032 1393
rect 16071 1359 16105 1393
rect 16144 1359 16178 1393
rect 16217 1359 16251 1393
rect 16290 1359 16324 1393
rect 16363 1359 16397 1393
rect 16436 1359 16470 1393
rect 16510 1359 16544 1393
rect 16584 1359 16618 1393
rect 16658 1359 16692 1393
rect 16732 1359 16766 1393
rect 16806 1359 16840 1393
rect 16880 1359 16914 1393
rect 15560 1285 15594 1319
rect 15633 1285 15667 1319
rect 15706 1285 15740 1319
rect 15779 1285 15813 1319
rect 15852 1285 15886 1319
rect 15925 1285 15944 1319
rect 15944 1285 15959 1319
rect 15998 1285 16032 1319
rect 16071 1285 16105 1319
rect 16144 1285 16178 1319
rect 16217 1285 16251 1319
rect 16290 1285 16324 1319
rect 16363 1285 16397 1319
rect 16436 1285 16470 1319
rect 16510 1285 16544 1319
rect 16584 1285 16618 1319
rect 16658 1285 16692 1319
rect 16732 1285 16766 1319
rect 16806 1285 16840 1319
rect 16880 1285 16914 1319
rect 5298 1214 5332 1248
rect 5371 1214 5405 1248
rect 5444 1214 5478 1248
rect 5517 1214 5551 1248
rect 5590 1214 5624 1248
rect 5663 1214 5697 1248
rect 5736 1214 5770 1248
rect 5809 1214 5843 1248
rect 5882 1214 5916 1248
rect 8644 798 8672 813
rect 8672 798 8678 813
rect 8718 798 8740 813
rect 8740 798 8752 813
rect 8792 798 8808 813
rect 8808 798 8826 813
rect 8866 798 8876 813
rect 8876 798 8900 813
rect 8940 798 8944 813
rect 8944 798 8974 813
rect 9014 798 9046 813
rect 9046 798 9048 813
rect 9088 798 9114 813
rect 9114 798 9122 813
rect 9162 798 9182 813
rect 9182 798 9196 813
rect 9236 798 9250 813
rect 9250 798 9270 813
rect 9310 798 9318 813
rect 9318 798 9344 813
rect 9384 798 9386 813
rect 9386 798 9418 813
rect 9458 798 9488 813
rect 9488 798 9492 813
rect 9532 798 9556 813
rect 9556 798 9566 813
rect 9606 798 9624 813
rect 9624 798 9640 813
rect 9680 798 9692 813
rect 9692 798 9714 813
rect 9754 798 9760 813
rect 9760 798 9788 813
rect 9827 798 9828 813
rect 9828 798 9861 813
rect 9900 798 9930 813
rect 9930 798 9934 813
rect 9973 798 9998 813
rect 9998 798 10007 813
rect 10046 798 10066 813
rect 10066 798 10080 813
rect 10119 798 10134 813
rect 10134 798 10153 813
rect 10192 798 10202 813
rect 10202 798 10226 813
rect 10265 798 10270 813
rect 10270 798 10299 813
rect 10338 798 10372 813
rect 10411 798 10440 813
rect 10440 798 10445 813
rect 10484 798 10508 813
rect 10508 798 10518 813
rect 8644 779 8678 798
rect 8718 779 8752 798
rect 8792 779 8826 798
rect 8866 779 8900 798
rect 8940 779 8974 798
rect 9014 779 9048 798
rect 9088 779 9122 798
rect 9162 779 9196 798
rect 9236 779 9270 798
rect 9310 779 9344 798
rect 9384 779 9418 798
rect 9458 779 9492 798
rect 9532 779 9566 798
rect 9606 779 9640 798
rect 9680 779 9714 798
rect 9754 779 9788 798
rect 9827 779 9861 798
rect 9900 779 9934 798
rect 9973 779 10007 798
rect 10046 779 10080 798
rect 10119 779 10153 798
rect 10192 779 10226 798
rect 10265 779 10299 798
rect 10338 779 10372 798
rect 10411 779 10445 798
rect 10484 779 10518 798
rect 10557 779 10591 813
rect 10630 779 10664 813
rect 10703 779 10737 813
rect 14682 760 14716 794
rect 14754 760 14788 794
rect 6579 674 6583 708
rect 6583 674 6613 708
rect 6659 674 6686 708
rect 6686 674 6693 708
rect 6739 674 6755 708
rect 6755 674 6773 708
rect 6818 674 6824 708
rect 6824 674 6852 708
rect 6522 596 6556 630
rect 6594 596 6628 630
rect 14682 562 14716 596
rect 14754 562 14788 596
rect 15560 1211 15594 1245
rect 15633 1211 15667 1245
rect 15706 1211 15740 1245
rect 15779 1211 15813 1245
rect 15852 1211 15886 1245
rect 15925 1211 15944 1245
rect 15944 1211 15959 1245
rect 15998 1211 16032 1245
rect 16071 1211 16105 1245
rect 16144 1211 16178 1245
rect 16217 1211 16251 1245
rect 16290 1211 16324 1245
rect 16363 1211 16397 1245
rect 16436 1211 16470 1245
rect 16510 1211 16544 1245
rect 16584 1211 16618 1245
rect 16658 1211 16692 1245
rect 16732 1211 16766 1245
rect 16806 1211 16840 1245
rect 16880 1211 16914 1245
rect 15648 -1314 15944 808
rect 15944 -1314 16546 808
rect 15648 -1387 15682 -1353
rect 15720 -1387 15754 -1353
rect 15792 -1387 15826 -1353
rect 15864 -1387 15898 -1353
rect 15936 -1387 15944 -1353
rect 15944 -1387 15970 -1353
rect 16008 -1387 16042 -1353
rect 16080 -1387 16114 -1353
rect 16152 -1387 16186 -1353
rect 16224 -1387 16258 -1353
rect 16296 -1387 16330 -1353
rect 16368 -1387 16402 -1353
rect 16440 -1387 16474 -1353
rect 16512 -1387 16546 -1353
rect 15648 -1460 15682 -1426
rect 15720 -1460 15754 -1426
rect 15792 -1460 15826 -1426
rect 15864 -1460 15898 -1426
rect 15936 -1460 15944 -1426
rect 15944 -1460 15970 -1426
rect 16008 -1460 16042 -1426
rect 16080 -1460 16114 -1426
rect 16152 -1460 16186 -1426
rect 16224 -1460 16258 -1426
rect 16296 -1460 16330 -1426
rect 16368 -1460 16402 -1426
rect 16440 -1460 16474 -1426
rect 16512 -1460 16546 -1426
rect 15648 -1533 15682 -1499
rect 15720 -1533 15754 -1499
rect 15792 -1533 15826 -1499
rect 15864 -1533 15898 -1499
rect 15936 -1533 15944 -1499
rect 15944 -1533 15970 -1499
rect 16008 -1533 16042 -1499
rect 16080 -1533 16114 -1499
rect 16152 -1533 16186 -1499
rect 16224 -1533 16258 -1499
rect 16296 -1533 16330 -1499
rect 16368 -1533 16402 -1499
rect 16440 -1533 16474 -1499
rect 16512 -1533 16546 -1499
rect 15648 -1606 15682 -1572
rect 15720 -1606 15754 -1572
rect 15792 -1606 15826 -1572
rect 15864 -1606 15898 -1572
rect 15936 -1606 15944 -1572
rect 15944 -1606 15970 -1572
rect 16008 -1606 16042 -1572
rect 16080 -1606 16114 -1572
rect 16152 -1606 16186 -1572
rect 16224 -1606 16258 -1572
rect 16296 -1606 16330 -1572
rect 16368 -1606 16402 -1572
rect 16440 -1606 16474 -1572
rect 16512 -1606 16546 -1572
rect 15648 -1679 15682 -1645
rect 15720 -1679 15754 -1645
rect 15792 -1679 15826 -1645
rect 15864 -1679 15898 -1645
rect 15936 -1679 15944 -1645
rect 15944 -1679 15970 -1645
rect 16008 -1679 16042 -1645
rect 16080 -1679 16114 -1645
rect 16152 -1679 16186 -1645
rect 16224 -1679 16258 -1645
rect 16296 -1679 16330 -1645
rect 16368 -1679 16402 -1645
rect 16440 -1679 16474 -1645
rect 16512 -1679 16546 -1645
<< metal1 >>
tri 6916 27018 6961 27063 sw
tri 859 26814 960 26915 sw
rect 859 26810 960 26814
tri 960 26810 964 26814 sw
rect 24081 26762 24087 26814
rect 24139 26762 24181 26814
rect 24233 26762 24274 26814
rect 24326 26762 24332 26814
rect 24081 26750 24332 26762
rect 24081 26698 24087 26750
rect 24139 26698 24181 26750
rect 24233 26698 24274 26750
rect 24326 26698 24332 26750
rect 19265 22193 19271 22245
rect 19323 22193 19341 22245
rect 19393 22193 19411 22245
rect 19463 22193 19480 22245
rect 19532 22193 19549 22245
rect 19601 22193 19618 22245
rect 19670 22193 19687 22245
rect 19739 22193 19756 22245
rect 19808 22193 19825 22245
rect 19877 22193 19883 22245
rect 19265 22181 19883 22193
rect 19265 22129 19271 22181
rect 19323 22129 19341 22181
rect 19393 22129 19411 22181
rect 19463 22129 19480 22181
rect 19532 22129 19549 22181
rect 19601 22129 19618 22181
rect 19670 22129 19687 22181
rect 19739 22129 19756 22181
rect 19808 22129 19825 22181
rect 19877 22129 19883 22181
rect 21006 22193 21012 22245
rect 21064 22193 21079 22245
rect 21131 22193 21146 22245
rect 21198 22193 21213 22245
rect 21265 22193 21280 22245
rect 21332 22193 21347 22245
rect 21399 22193 21414 22245
rect 21466 22193 21481 22245
rect 21533 22193 21548 22245
rect 21600 22193 21615 22245
rect 21667 22193 21681 22245
rect 21733 22193 21747 22245
rect 21799 22193 21813 22245
rect 21865 22193 21871 22245
rect 21006 22181 21871 22193
rect 21006 22129 21012 22181
rect 21064 22129 21079 22181
rect 21131 22129 21146 22181
rect 21198 22129 21213 22181
rect 21265 22129 21280 22181
rect 21332 22129 21347 22181
rect 21399 22129 21414 22181
rect 21466 22129 21481 22181
rect 21533 22129 21548 22181
rect 21600 22129 21615 22181
rect 21667 22129 21681 22181
rect 21733 22129 21747 22181
rect 21799 22129 21813 22181
rect 21865 22129 21871 22181
rect 17482 22077 17598 22083
tri 16904 22025 16956 22077 se
rect 16956 22071 17443 22077
rect 16956 22025 17327 22071
rect 16938 22007 17327 22025
rect 16911 21955 17327 22007
rect 17482 21955 17598 21961
rect 17636 22077 19469 22089
rect 17752 21961 19347 22077
rect 19463 21961 19469 22077
rect 16938 21931 17443 21955
rect 17636 21951 19469 21961
rect 20260 21827 20266 21879
rect 20318 21827 20355 21879
rect 20407 21827 20443 21879
rect 20495 21827 20501 21879
rect 5518 21776 5592 21822
rect 5518 21763 5579 21776
tri 5579 21763 5592 21776 nw
rect 20260 21815 20501 21827
rect 20260 21763 20266 21815
rect 20318 21763 20355 21815
rect 20407 21763 20443 21815
rect 20495 21763 20501 21815
rect 5518 21706 5522 21763
tri 5522 21706 5579 21763 nw
rect 23736 19733 23742 19785
rect 23794 19733 23806 19785
rect 23858 19733 23864 19785
rect 20260 19649 20266 19701
rect 20318 19649 20355 19701
rect 20407 19649 20444 19701
rect 20496 19649 20502 19701
rect 20260 19637 20502 19649
rect 20260 19585 20266 19637
rect 20318 19585 20355 19637
rect 20407 19585 20444 19637
rect 20496 19585 20502 19637
tri 30847 19474 30872 19499 sw
tri 30952 19474 30977 19499 se
rect 30847 19424 30977 19474
tri 30952 19399 30977 19424 ne
rect 19221 18782 20558 18801
rect 19221 18730 19227 18782
rect 19279 18730 19294 18782
rect 19346 18730 19361 18782
rect 19413 18730 19428 18782
rect 19480 18730 19495 18782
rect 19547 18730 19562 18782
rect 19614 18730 19629 18782
rect 19681 18730 19696 18782
rect 19748 18730 19763 18782
rect 19815 18730 19830 18782
rect 19882 18730 19897 18782
rect 19949 18730 19964 18782
rect 20016 18730 20031 18782
rect 20083 18730 20098 18782
rect 20150 18730 20165 18782
rect 20217 18730 20232 18782
rect 20284 18730 20299 18782
rect 20351 18730 20366 18782
rect 20418 18730 20433 18782
rect 20485 18730 20500 18782
rect 20552 18730 20558 18782
rect 19221 18718 20558 18730
rect 19221 18666 19227 18718
rect 19279 18666 19294 18718
rect 19346 18666 19361 18718
rect 19413 18666 19428 18718
rect 19480 18666 19495 18718
rect 19547 18666 19562 18718
rect 19614 18666 19629 18718
rect 19681 18666 19696 18718
rect 19748 18666 19763 18718
rect 19815 18666 19830 18718
rect 19882 18666 19897 18718
rect 19949 18666 19964 18718
rect 20016 18666 20031 18718
rect 20083 18666 20098 18718
rect 20150 18666 20165 18718
rect 20217 18666 20232 18718
rect 20284 18666 20299 18718
rect 20351 18666 20366 18718
rect 20418 18666 20433 18718
rect 20485 18666 20500 18718
rect 20552 18666 20558 18718
rect 19221 18654 20558 18666
rect 19221 18602 19227 18654
rect 19279 18602 19294 18654
rect 19346 18602 19361 18654
rect 19413 18602 19428 18654
rect 19480 18602 19495 18654
rect 19547 18602 19562 18654
rect 19614 18602 19629 18654
rect 19681 18602 19696 18654
rect 19748 18602 19763 18654
rect 19815 18602 19830 18654
rect 19882 18602 19897 18654
rect 19949 18602 19964 18654
rect 20016 18602 20031 18654
rect 20083 18602 20098 18654
rect 20150 18602 20165 18654
rect 20217 18602 20232 18654
rect 20284 18602 20299 18654
rect 20351 18602 20366 18654
rect 20418 18602 20433 18654
rect 20485 18602 20500 18654
rect 20552 18602 20558 18654
rect 19221 18590 20558 18602
rect 19221 18538 19227 18590
rect 19279 18538 19294 18590
rect 19346 18538 19361 18590
rect 19413 18538 19428 18590
rect 19480 18538 19495 18590
rect 19547 18538 19562 18590
rect 19614 18538 19629 18590
rect 19681 18538 19696 18590
rect 19748 18538 19763 18590
rect 19815 18538 19830 18590
rect 19882 18538 19897 18590
rect 19949 18538 19964 18590
rect 20016 18538 20031 18590
rect 20083 18538 20098 18590
rect 20150 18538 20165 18590
rect 20217 18538 20232 18590
rect 20284 18538 20299 18590
rect 20351 18538 20366 18590
rect 20418 18538 20433 18590
rect 20485 18538 20500 18590
rect 20552 18538 20558 18590
rect 19221 18519 20558 18538
rect 21042 18781 21720 18805
rect 21042 18729 21048 18781
rect 21100 18729 21117 18781
rect 21169 18729 21186 18781
rect 21238 18729 21254 18781
rect 21306 18729 21322 18781
rect 21374 18729 21390 18781
rect 21442 18729 21458 18781
rect 21510 18729 21526 18781
rect 21578 18729 21594 18781
rect 21646 18729 21662 18781
rect 21714 18729 21720 18781
rect 21042 18717 21720 18729
rect 21042 18665 21048 18717
rect 21100 18665 21117 18717
rect 21169 18665 21186 18717
rect 21238 18665 21254 18717
rect 21306 18665 21322 18717
rect 21374 18665 21390 18717
rect 21442 18665 21458 18717
rect 21510 18665 21526 18717
rect 21578 18665 21594 18717
rect 21646 18665 21662 18717
rect 21714 18665 21720 18717
rect 21042 18653 21720 18665
rect 21042 18601 21048 18653
rect 21100 18601 21117 18653
rect 21169 18601 21186 18653
rect 21238 18601 21254 18653
rect 21306 18601 21322 18653
rect 21374 18601 21390 18653
rect 21442 18601 21458 18653
rect 21510 18601 21526 18653
rect 21578 18601 21594 18653
rect 21646 18601 21662 18653
rect 21714 18601 21720 18653
rect 21042 18589 21720 18601
rect 21042 18537 21048 18589
rect 21100 18537 21117 18589
rect 21169 18537 21186 18589
rect 21238 18537 21254 18589
rect 21306 18537 21322 18589
rect 21374 18537 21390 18589
rect 21442 18537 21458 18589
rect 21510 18537 21526 18589
rect 21578 18537 21594 18589
rect 21646 18537 21662 18589
rect 21714 18537 21720 18589
rect 31004 18791 31426 18797
rect 31004 18739 31029 18791
rect 31081 18739 31093 18791
rect 31145 18739 31157 18791
rect 31209 18739 31221 18791
rect 31273 18739 31285 18791
rect 31337 18739 31349 18791
rect 31401 18739 31426 18791
rect 31004 18724 31426 18739
rect 31004 18672 31029 18724
rect 31081 18672 31093 18724
rect 31145 18672 31157 18724
rect 31209 18672 31221 18724
rect 31273 18672 31285 18724
rect 31337 18672 31349 18724
rect 31401 18672 31426 18724
rect 31004 18657 31426 18672
rect 31004 18605 31029 18657
rect 31081 18605 31093 18657
rect 31145 18605 31157 18657
rect 31209 18605 31221 18657
rect 31273 18605 31285 18657
rect 31337 18605 31349 18657
rect 31401 18605 31426 18657
rect 31004 18590 31426 18605
tri 30952 18544 30977 18569 se
rect 21042 18513 21720 18537
rect 31004 18538 31029 18590
rect 31081 18538 31093 18590
rect 31145 18538 31157 18590
rect 31209 18538 31221 18590
rect 31273 18538 31285 18590
rect 31337 18538 31349 18590
rect 31401 18538 31426 18590
rect 31004 18523 31426 18538
tri 30952 18473 30977 18498 ne
rect 31004 18471 31029 18523
rect 31081 18471 31093 18523
rect 31145 18471 31157 18523
rect 31209 18471 31221 18523
rect 31273 18471 31285 18523
rect 31337 18471 31349 18523
rect 31401 18471 31426 18523
rect 31004 18456 31426 18471
rect 31004 18404 31029 18456
rect 31081 18404 31093 18456
rect 31145 18404 31157 18456
rect 31209 18404 31221 18456
rect 31273 18404 31285 18456
rect 31337 18404 31349 18456
rect 31401 18404 31426 18456
rect 31004 18389 31426 18404
rect 31004 18337 31029 18389
rect 31081 18337 31093 18389
rect 31145 18337 31157 18389
rect 31209 18337 31221 18389
rect 31273 18337 31285 18389
rect 31337 18337 31349 18389
rect 31401 18337 31426 18389
rect 31004 18322 31426 18337
rect 31004 18270 31029 18322
rect 31081 18270 31093 18322
rect 31145 18270 31157 18322
rect 31209 18270 31221 18322
rect 31273 18270 31285 18322
rect 31337 18270 31349 18322
rect 31401 18270 31426 18322
rect 31004 18255 31426 18270
rect 31004 18203 31029 18255
rect 31081 18203 31093 18255
rect 31145 18203 31157 18255
rect 31209 18203 31221 18255
rect 31273 18203 31285 18255
rect 31337 18203 31349 18255
rect 31401 18203 31426 18255
rect 31004 18188 31426 18203
tri 22930 18138 22955 18163 nw
rect 31004 18136 31029 18188
rect 31081 18136 31093 18188
rect 31145 18136 31157 18188
rect 31209 18136 31221 18188
rect 31273 18136 31285 18188
rect 31337 18136 31349 18188
rect 31401 18136 31426 18188
rect 31004 18121 31426 18136
rect 31004 18069 31029 18121
rect 31081 18069 31093 18121
rect 31145 18069 31157 18121
rect 31209 18069 31221 18121
rect 31273 18069 31285 18121
rect 31337 18069 31349 18121
rect 31401 18069 31426 18121
rect 31004 18063 31426 18069
rect 16055 15797 16056 15855
rect 23032 14365 23038 14417
rect 23090 14365 23102 14417
rect 23154 14416 23160 14417
tri 23160 14416 23161 14417 sw
tri 23754 14416 23755 14417 se
rect 23755 14416 23761 14417
rect 23154 14376 23761 14416
rect 23154 14365 23160 14376
tri 23160 14365 23171 14376 nw
tri 23744 14365 23755 14376 ne
rect 23755 14365 23761 14376
rect 23813 14365 23825 14417
rect 23877 14365 23883 14417
tri 17561 8545 17720 8704 sw
tri 17561 8140 17720 8299 nw
rect 19429 8083 22725 8113
rect 19429 8031 19435 8083
rect 19487 8031 19503 8083
rect 19555 8031 19571 8083
rect 19623 8031 19639 8083
rect 19691 8031 19707 8083
rect 19759 8031 19775 8083
rect 19827 8031 19842 8083
rect 19894 8031 20844 8083
rect 20896 8031 20926 8083
rect 20978 8031 21008 8083
rect 21060 8031 21090 8083
rect 21142 8031 21634 8083
rect 21686 8031 21701 8083
rect 21753 8031 21768 8083
rect 21820 8031 21834 8083
rect 21886 8031 21900 8083
rect 21952 8031 21966 8083
rect 22018 8031 22239 8083
rect 22291 8031 22309 8083
rect 22361 8031 22379 8083
rect 22431 8031 22448 8083
rect 22500 8031 22517 8083
rect 22569 8031 22586 8083
rect 22638 8031 22655 8083
rect 22707 8031 22725 8083
rect 19429 8019 22725 8031
rect 19429 7967 19435 8019
rect 19487 7967 19503 8019
rect 19555 7967 19571 8019
rect 19623 7967 19639 8019
rect 19691 7967 19707 8019
rect 19759 7967 19775 8019
rect 19827 7967 19842 8019
rect 19894 7967 20844 8019
rect 20896 7967 20926 8019
rect 20978 7967 21008 8019
rect 21060 7967 21090 8019
rect 21142 7967 21634 8019
rect 21686 7967 21701 8019
rect 21753 7967 21768 8019
rect 21820 7967 21834 8019
rect 21886 7967 21900 8019
rect 21952 7967 21966 8019
rect 22018 7967 22239 8019
rect 22291 7967 22309 8019
rect 22361 7967 22379 8019
rect 22431 7967 22448 8019
rect 22500 7967 22517 8019
rect 22569 7967 22586 8019
rect 22638 7967 22655 8019
rect 22707 7967 22725 8019
rect 19429 7955 22725 7967
rect 19429 7903 19435 7955
rect 19487 7903 19503 7955
rect 19555 7903 19571 7955
rect 19623 7903 19639 7955
rect 19691 7903 19707 7955
rect 19759 7903 19775 7955
rect 19827 7903 19842 7955
rect 19894 7903 20844 7955
rect 20896 7903 20926 7955
rect 20978 7903 21008 7955
rect 21060 7903 21090 7955
rect 21142 7903 21634 7955
rect 21686 7903 21701 7955
rect 21753 7903 21768 7955
rect 21820 7903 21834 7955
rect 21886 7903 21900 7955
rect 21952 7903 21966 7955
rect 22018 7903 22239 7955
rect 22291 7903 22309 7955
rect 22361 7903 22379 7955
rect 22431 7903 22448 7955
rect 22500 7903 22517 7955
rect 22569 7903 22586 7955
rect 22638 7903 22655 7955
rect 22707 7903 22725 7955
rect 19429 7872 22725 7903
rect 22460 6184 22466 6300
rect 22582 6184 22588 6300
rect 15813 5198 15868 5252
tri 5958 4714 5996 4752 se
rect -3209 4560 -3157 4566
rect -3209 4496 -3157 4508
rect -2889 4552 -2837 4558
rect -2889 4488 -2837 4500
rect -3209 4438 -3157 4444
tri -3157 4438 -3134 4461 sw
tri -3208 4425 -3195 4438 ne
rect -3195 4430 -3134 4438
tri -3134 4430 -3126 4438 sw
rect -2889 4430 -2837 4436
rect -2809 4552 -2757 4558
rect -2809 4488 -2757 4500
rect -2809 4430 -2757 4436
rect -2729 4539 -2677 4545
rect -2729 4475 -2677 4487
rect -3195 4425 -3126 4430
tri -3126 4425 -3121 4430 sw
tri -3195 4397 -3167 4425 ne
rect -3167 4417 -3121 4425
tri -3121 4417 -3113 4425 sw
rect -2569 4539 -2517 4545
rect -2569 4475 -2517 4487
tri -2677 4425 -2667 4435 sw
rect -2677 4423 -2667 4425
rect -2729 4417 -2667 4423
tri -2667 4417 -2659 4425 sw
rect 3884 4501 4540 4513
rect -2517 4467 3117 4469
tri 3117 4467 3119 4469 sw
rect 3884 4467 3891 4501
rect 3925 4467 3967 4501
rect 4001 4467 4043 4501
rect 4077 4467 4119 4501
rect 4153 4497 4195 4501
rect 4229 4497 4271 4501
rect 4305 4497 4347 4501
rect 4381 4497 4423 4501
rect 4457 4497 4499 4501
rect 4178 4467 4195 4497
rect -2517 4463 3119 4467
tri 3119 4463 3123 4467 sw
rect -2517 4425 3123 4463
tri 3123 4425 3161 4463 sw
rect 3884 4445 4126 4467
rect 4178 4445 4196 4467
rect 4248 4445 4266 4497
rect 4318 4445 4336 4497
rect 4388 4445 4406 4497
rect 4458 4445 4476 4497
rect 4533 4467 4540 4501
rect 4528 4445 4540 4467
rect 3884 4432 4540 4445
rect 3884 4425 4126 4432
rect 4178 4425 4196 4432
rect -2517 4423 3161 4425
rect -2569 4417 3161 4423
tri 3161 4417 3169 4425 sw
rect -3167 4397 -3113 4417
tri -3113 4397 -3093 4417 sw
rect -2729 4413 -2659 4417
tri -2729 4397 -2713 4413 ne
rect -2713 4397 -2659 4413
tri -2659 4397 -2639 4417 sw
tri 3095 4397 3115 4417 ne
rect 3115 4397 3169 4417
tri -3167 4391 -3161 4397 ne
rect -3161 4391 -2803 4397
tri -2803 4391 -2797 4397 sw
tri -2713 4391 -2707 4397 ne
rect -2707 4391 -2639 4397
tri -2639 4391 -2633 4397 sw
tri 3115 4391 3121 4397 ne
rect 3121 4391 3169 4397
tri 3169 4391 3195 4417 sw
rect 3884 4391 3891 4425
rect 3925 4391 3967 4425
rect 4001 4391 4043 4425
rect 4077 4391 4119 4425
rect 4178 4391 4195 4425
tri -3161 4387 -3157 4391 ne
rect -3157 4389 -2797 4391
tri -2797 4389 -2795 4391 sw
tri -2707 4389 -2705 4391 ne
rect -2705 4389 -2633 4391
tri -2633 4389 -2631 4391 sw
tri 3121 4389 3123 4391 ne
rect 3123 4389 3195 4391
tri 3195 4389 3197 4391 sw
rect -3157 4387 -2795 4389
tri -3157 4374 -3144 4387 ne
rect -3144 4374 -2795 4387
tri -2795 4374 -2780 4389 sw
tri -2705 4384 -2700 4389 ne
rect -2700 4384 -2631 4389
tri -2631 4384 -2626 4389 sw
tri 3123 4384 3128 4389 ne
rect 3128 4384 3197 4389
tri -2700 4378 -2694 4384 ne
rect -2694 4378 3069 4384
tri 3069 4378 3075 4384 sw
tri 3128 4378 3134 4384 ne
rect 3134 4378 3197 4384
tri -2694 4374 -2690 4378 ne
rect -2690 4374 3075 4378
tri 3075 4374 3079 4378 sw
tri 3134 4374 3138 4378 ne
rect 3138 4374 3197 4378
tri -3144 4349 -3119 4374 ne
rect -3119 4361 -2780 4374
tri -2780 4361 -2767 4374 sw
tri -2690 4361 -2677 4374 ne
rect -2677 4363 3079 4374
tri 3079 4363 3090 4374 sw
tri 3138 4363 3149 4374 ne
rect 3149 4363 3197 4374
rect -2677 4361 3090 4363
rect -3119 4349 -2767 4361
tri -2767 4349 -2755 4361 sw
tri -2677 4349 -2665 4361 ne
rect -2665 4349 3090 4361
tri 3090 4349 3104 4363 sw
tri 3149 4349 3163 4363 ne
rect 3163 4349 3197 4363
tri 3197 4349 3237 4389 sw
rect 3884 4380 4126 4391
rect 4178 4380 4196 4391
rect 4248 4380 4266 4432
rect 4318 4380 4336 4432
rect 4388 4380 4406 4432
rect 4458 4380 4476 4432
rect 4528 4425 4540 4432
rect 4533 4391 4540 4425
tri 11275 4417 11334 4476 se
rect 11334 4417 16940 4476
rect 4528 4380 4540 4391
rect 3884 4367 4540 4380
rect 3884 4349 4126 4367
rect 4178 4349 4196 4367
tri -3119 4345 -3115 4349 ne
rect -3115 4345 -2755 4349
tri -2821 4315 -2791 4345 ne
rect -2791 4315 -2755 4345
tri -2755 4315 -2721 4349 sw
tri -2665 4332 -2648 4349 ne
rect -2648 4332 3104 4349
tri 3047 4315 3064 4332 ne
rect 3064 4315 3104 4332
tri 3104 4315 3138 4349 sw
tri 3163 4315 3197 4349 ne
rect 3197 4315 3237 4349
tri 3237 4315 3271 4349 sw
rect 3884 4315 3891 4349
rect 3925 4315 3967 4349
rect 4001 4315 4043 4349
rect 4077 4315 4119 4349
rect 4178 4315 4195 4349
rect 4248 4315 4266 4367
rect 4318 4315 4336 4367
rect 4388 4315 4406 4367
rect 4458 4315 4476 4367
rect 4528 4349 4540 4367
rect 4533 4315 4540 4349
tri -2791 4304 -2780 4315 ne
rect -2780 4304 -2721 4315
tri -2721 4304 -2710 4315 sw
tri 3064 4304 3075 4315 ne
rect 3075 4304 3138 4315
tri 3138 4304 3149 4315 sw
tri 3197 4304 3208 4315 ne
rect 3208 4304 3271 4315
tri 3271 4304 3282 4315 sw
tri -2780 4288 -2764 4304 ne
rect -2764 4298 3007 4304
tri 3007 4298 3013 4304 sw
tri 3075 4298 3081 4304 ne
rect 3081 4298 3149 4304
tri 3149 4298 3155 4304 sw
tri 3208 4298 3214 4304 ne
rect 3214 4298 3282 4304
tri 3282 4298 3288 4304 sw
rect 3884 4302 4540 4315
rect -2764 4288 3013 4298
tri 3013 4288 3023 4298 sw
tri 3081 4288 3091 4298 ne
rect 3091 4289 3155 4298
tri 3155 4289 3164 4298 sw
tri 3214 4289 3223 4298 ne
rect 3223 4289 3288 4298
rect 3091 4288 3164 4289
tri 3164 4288 3165 4289 sw
tri 3223 4288 3224 4289 ne
rect 3224 4288 3288 4289
tri 3288 4288 3298 4298 sw
tri -2764 4273 -2749 4288 ne
rect -2749 4273 3023 4288
tri 3023 4273 3038 4288 sw
tri 3091 4273 3106 4288 ne
rect 3106 4273 3165 4288
tri 3165 4273 3180 4288 sw
tri 3224 4273 3239 4288 ne
rect 3239 4273 3298 4288
tri 3298 4273 3313 4288 sw
rect 3884 4273 4126 4302
rect 4178 4273 4196 4302
tri -2749 4252 -2728 4273 ne
rect -2728 4252 3038 4273
tri 2985 4239 2998 4252 ne
rect 2998 4239 3038 4252
tri 3038 4239 3072 4273 sw
tri 3106 4239 3140 4273 ne
rect 3140 4241 3180 4273
tri 3180 4241 3212 4273 sw
tri 3239 4241 3271 4273 ne
rect 3271 4241 3313 4273
tri 3313 4241 3345 4273 sw
rect 3140 4239 3212 4241
tri 3212 4239 3214 4241 sw
tri 3271 4239 3273 4241 ne
rect 3273 4239 3345 4241
tri 3345 4239 3347 4241 sw
rect 3884 4239 3891 4273
rect 3925 4239 3967 4273
rect 4001 4239 4043 4273
rect 4077 4239 4119 4273
rect 4178 4250 4195 4273
rect 4248 4250 4266 4302
rect 4318 4250 4336 4302
rect 4388 4250 4406 4302
rect 4458 4250 4476 4302
rect 4528 4273 4540 4302
rect 4153 4239 4195 4250
rect 4229 4239 4271 4250
rect 4305 4239 4347 4250
rect 4381 4239 4423 4250
rect 4457 4239 4499 4250
rect 4533 4239 4540 4273
tri 2998 4224 3013 4239 ne
rect 3013 4236 3072 4239
tri 3072 4236 3075 4239 sw
tri 3140 4236 3143 4239 ne
rect 3143 4236 3214 4239
rect 3013 4230 3075 4236
tri 3075 4230 3081 4236 sw
tri 3143 4230 3149 4236 ne
rect 3149 4230 3214 4236
tri 3214 4230 3223 4239 sw
tri 3273 4230 3282 4239 ne
rect 3282 4230 3347 4239
rect 3013 4224 3081 4230
tri 3081 4224 3087 4230 sw
tri 3149 4224 3155 4230 ne
rect 3155 4224 3223 4230
tri 3223 4224 3229 4230 sw
tri 3282 4224 3288 4230 ne
rect 3288 4224 3347 4230
tri 3347 4224 3362 4239 sw
rect 3884 4237 4540 4239
tri 3013 4216 3021 4224 ne
rect 3021 4216 3087 4224
tri 3087 4216 3095 4224 sw
tri 3155 4216 3163 4224 ne
rect 3163 4216 3229 4224
tri 3229 4216 3237 4224 sw
tri 3288 4216 3296 4224 ne
rect 3296 4216 3362 4224
tri 3362 4216 3370 4224 sw
tri 3021 4197 3040 4216 ne
rect 3040 4197 3095 4216
tri 3095 4197 3114 4216 sw
tri 3163 4197 3182 4216 ne
rect 3182 4215 3237 4216
tri 3237 4215 3238 4216 sw
tri 3296 4215 3297 4216 ne
rect 3297 4215 3370 4216
rect 3182 4197 3238 4215
tri 3238 4197 3256 4215 sw
tri 3297 4197 3315 4215 ne
rect 3315 4197 3370 4215
tri 3370 4197 3389 4216 sw
rect 3884 4197 4126 4237
rect 4178 4197 4196 4237
tri 3040 4163 3074 4197 ne
rect 3074 4163 3114 4197
tri 3114 4163 3148 4197 sw
tri 3182 4163 3216 4197 ne
rect 3216 4167 3256 4197
tri 3256 4167 3286 4197 sw
tri 3315 4167 3345 4197 ne
rect 3345 4167 3389 4197
tri 3389 4167 3419 4197 sw
rect 3216 4163 3286 4167
tri 3286 4163 3290 4167 sw
tri 3345 4163 3349 4167 ne
rect 3349 4163 3419 4167
tri 3419 4163 3423 4167 sw
rect 3884 4163 3891 4197
rect 3925 4163 3967 4197
rect 4001 4163 4043 4197
rect 4077 4163 4119 4197
rect 4178 4185 4195 4197
rect 4248 4185 4266 4237
rect 4318 4185 4336 4237
rect 4388 4185 4406 4237
rect 4458 4185 4476 4237
rect 4528 4197 4540 4237
rect 4153 4171 4195 4185
rect 4229 4171 4271 4185
rect 4305 4171 4347 4185
rect 4381 4171 4423 4185
rect 4457 4171 4499 4185
rect 4178 4163 4195 4171
tri 3074 4150 3087 4163 ne
rect 3087 4162 3148 4163
tri 3148 4162 3149 4163 sw
tri 3216 4162 3217 4163 ne
rect 3217 4162 3290 4163
rect 3087 4156 3149 4162
tri 3149 4156 3155 4162 sw
tri 3217 4156 3223 4162 ne
rect 3223 4156 3290 4162
tri 3290 4156 3297 4163 sw
tri 3349 4156 3356 4163 ne
rect 3356 4156 3423 4163
rect 3087 4150 3155 4156
tri 3155 4150 3161 4156 sw
tri 3223 4150 3229 4156 ne
rect 3229 4150 3297 4156
tri 3297 4150 3303 4156 sw
tri 3356 4150 3362 4156 ne
rect 3362 4150 3423 4156
tri 3423 4150 3436 4163 sw
tri 3087 4144 3093 4150 ne
rect 3093 4144 3161 4150
tri 3161 4144 3167 4150 sw
tri 3229 4144 3235 4150 ne
rect 3235 4144 3303 4150
tri 3303 4144 3309 4150 sw
tri 3362 4144 3368 4150 ne
rect 3368 4144 3436 4150
tri 3436 4144 3442 4150 sw
tri 3093 4121 3116 4144 ne
rect 3116 4135 3167 4144
tri 3167 4135 3176 4144 sw
tri 3235 4135 3244 4144 ne
rect 3244 4141 3309 4144
tri 3309 4141 3312 4144 sw
tri 3368 4141 3371 4144 ne
rect 3371 4141 3442 4144
rect 3244 4135 3312 4141
tri 3312 4135 3318 4141 sw
tri 3371 4135 3377 4141 ne
rect 3377 4135 3442 4141
tri 3442 4135 3451 4144 sw
rect 3116 4121 3176 4135
tri 3176 4121 3190 4135 sw
tri 3244 4121 3258 4135 ne
rect 3258 4121 3318 4135
tri 3318 4121 3332 4135 sw
tri 3377 4121 3391 4135 ne
rect 3391 4121 3451 4135
tri 3451 4121 3465 4135 sw
rect 3884 4121 4126 4163
rect 4178 4121 4196 4163
tri 3116 4087 3150 4121 ne
rect 3150 4088 3190 4121
tri 3190 4088 3223 4121 sw
tri 3258 4088 3291 4121 ne
rect 3291 4093 3332 4121
tri 3332 4093 3360 4121 sw
tri 3391 4093 3419 4121 ne
rect 3419 4093 3465 4121
tri 3465 4093 3493 4121 sw
rect 3291 4088 3360 4093
rect 3150 4087 3223 4088
tri 3223 4087 3224 4088 sw
tri 3291 4087 3292 4088 ne
rect 3292 4087 3360 4088
tri 3360 4087 3366 4093 sw
tri 3419 4087 3425 4093 ne
rect 3425 4087 3493 4093
tri 3493 4087 3499 4093 sw
rect 3884 4087 3891 4121
rect 3925 4087 3967 4121
rect 4001 4087 4043 4121
rect 4077 4087 4119 4121
rect 4178 4119 4195 4121
rect 4248 4119 4266 4171
rect 4318 4119 4336 4171
rect 4388 4119 4406 4171
rect 4458 4119 4476 4171
rect 4533 4163 4540 4197
rect 4528 4121 4540 4163
tri 11227 4369 11275 4417 se
rect 11275 4369 16940 4417
rect 11227 4322 16940 4369
rect 11227 4288 11937 4322
rect 11971 4288 12010 4322
rect 12044 4288 12083 4322
rect 12117 4288 12156 4322
rect 12190 4288 12229 4322
rect 12263 4288 12302 4322
rect 12336 4288 12375 4322
rect 12409 4288 12448 4322
rect 12482 4288 12521 4322
rect 12555 4288 12594 4322
rect 12628 4288 12667 4322
rect 12701 4288 12740 4322
rect 12774 4288 12813 4322
rect 12847 4288 12886 4322
rect 12920 4288 12959 4322
rect 12993 4288 13032 4322
rect 13066 4288 13105 4322
rect 13139 4288 13178 4322
rect 13212 4288 13251 4322
rect 13285 4288 13324 4322
rect 13358 4288 13397 4322
rect 13431 4288 13470 4322
rect 13504 4288 13543 4322
rect 13577 4288 13616 4322
rect 13650 4288 13689 4322
rect 13723 4288 13762 4322
rect 13796 4288 13835 4322
rect 13869 4288 13908 4322
rect 13942 4288 13981 4322
rect 14015 4288 14054 4322
rect 14088 4288 14127 4322
rect 14161 4288 14200 4322
rect 14234 4288 14273 4322
rect 14307 4288 14346 4322
rect 14380 4288 14419 4322
rect 14453 4288 14492 4322
rect 14526 4288 14565 4322
rect 14599 4288 14638 4322
rect 14672 4288 14711 4322
rect 14745 4288 14784 4322
rect 14818 4288 14857 4322
rect 14891 4288 14930 4322
rect 14964 4288 15003 4322
rect 15037 4288 15076 4322
rect 15110 4288 15149 4322
rect 15183 4288 15222 4322
rect 15256 4288 15295 4322
rect 15329 4288 15368 4322
rect 15402 4288 15441 4322
rect 15475 4288 15514 4322
rect 15548 4288 15587 4322
rect 15621 4288 15660 4322
rect 15694 4288 15733 4322
rect 15767 4288 15806 4322
rect 15840 4288 15879 4322
rect 15913 4288 15952 4322
rect 15986 4288 16025 4322
rect 16059 4288 16098 4322
rect 16132 4288 16171 4322
rect 16205 4288 16244 4322
rect 16278 4288 16317 4322
rect 16351 4288 16390 4322
rect 11227 4250 16390 4288
rect 11227 4216 11937 4250
rect 11971 4216 12010 4250
rect 12044 4216 12083 4250
rect 12117 4216 12156 4250
rect 12190 4216 12229 4250
rect 12263 4216 12302 4250
rect 12336 4216 12375 4250
rect 12409 4216 12448 4250
rect 12482 4216 12521 4250
rect 12555 4216 12594 4250
rect 12628 4216 12667 4250
rect 12701 4216 12740 4250
rect 12774 4216 12813 4250
rect 12847 4216 12886 4250
rect 12920 4216 12959 4250
rect 12993 4216 13032 4250
rect 13066 4216 13105 4250
rect 13139 4216 13178 4250
rect 13212 4216 13251 4250
rect 13285 4216 13324 4250
rect 13358 4216 13397 4250
rect 13431 4216 13470 4250
rect 13504 4216 13543 4250
rect 13577 4216 13616 4250
rect 13650 4216 13689 4250
rect 13723 4216 13762 4250
rect 13796 4216 13835 4250
rect 13869 4216 13908 4250
rect 13942 4216 13981 4250
rect 14015 4216 14054 4250
rect 14088 4216 14127 4250
rect 14161 4216 14200 4250
rect 14234 4216 14273 4250
rect 14307 4216 14346 4250
rect 14380 4216 14419 4250
rect 14453 4216 14492 4250
rect 14526 4216 14565 4250
rect 14599 4216 14638 4250
rect 14672 4216 14711 4250
rect 14745 4216 14784 4250
rect 14818 4216 14857 4250
rect 14891 4216 14930 4250
rect 14964 4216 15003 4250
rect 15037 4216 15076 4250
rect 15110 4216 15149 4250
rect 15183 4216 15222 4250
rect 15256 4216 15295 4250
rect 15329 4216 15368 4250
rect 15402 4216 15441 4250
rect 15475 4216 15514 4250
rect 15548 4216 15587 4250
rect 15621 4216 15660 4250
rect 15694 4216 15733 4250
rect 15767 4216 15806 4250
rect 15840 4216 15879 4250
rect 15913 4216 15952 4250
rect 15986 4216 16025 4250
rect 16059 4216 16098 4250
rect 16132 4216 16171 4250
rect 16205 4216 16244 4250
rect 16278 4216 16317 4250
rect 16351 4216 16390 4250
rect 11227 4178 16390 4216
rect 11227 4144 11937 4178
rect 11971 4144 12010 4178
rect 12044 4144 12083 4178
rect 12117 4144 12156 4178
rect 12190 4144 12229 4178
rect 12263 4144 12302 4178
rect 12336 4144 12375 4178
rect 12409 4144 12448 4178
rect 12482 4144 12521 4178
rect 12555 4144 12594 4178
rect 12628 4144 12667 4178
rect 12701 4144 12740 4178
rect 12774 4144 12813 4178
rect 12847 4144 12886 4178
rect 12920 4144 12959 4178
rect 12993 4144 13032 4178
rect 13066 4144 13105 4178
rect 13139 4144 13178 4178
rect 13212 4144 13251 4178
rect 13285 4144 13324 4178
rect 13358 4144 13397 4178
rect 13431 4144 13470 4178
rect 13504 4144 13543 4178
rect 13577 4144 13616 4178
rect 13650 4144 13689 4178
rect 13723 4144 13762 4178
rect 13796 4144 13835 4178
rect 13869 4144 13908 4178
rect 13942 4144 13981 4178
rect 14015 4144 14054 4178
rect 14088 4144 14127 4178
rect 14161 4144 14200 4178
rect 14234 4144 14273 4178
rect 14307 4144 14346 4178
rect 14380 4144 14419 4178
rect 14453 4144 14492 4178
rect 14526 4144 14565 4178
rect 14599 4144 14638 4178
rect 14672 4144 14711 4178
rect 14745 4144 14784 4178
rect 14818 4144 14857 4178
rect 14891 4144 14930 4178
rect 14964 4144 15003 4178
rect 15037 4144 15076 4178
rect 15110 4144 15149 4178
rect 15183 4144 15222 4178
rect 15256 4144 15295 4178
rect 15329 4144 15368 4178
rect 15402 4144 15441 4178
rect 15475 4144 15514 4178
rect 15548 4144 15587 4178
rect 15621 4144 15660 4178
rect 15694 4144 15733 4178
rect 15767 4144 15806 4178
rect 15840 4144 15879 4178
rect 15913 4144 15952 4178
rect 15986 4144 16025 4178
rect 16059 4144 16098 4178
rect 16132 4144 16171 4178
rect 16205 4144 16244 4178
rect 16278 4144 16317 4178
rect 16351 4144 16390 4178
rect 4153 4105 4195 4119
rect 4229 4105 4271 4119
rect 4305 4105 4347 4119
rect 4381 4105 4423 4119
rect 4457 4105 4499 4119
rect 4178 4087 4195 4105
tri 3150 4076 3161 4087 ne
rect 3161 4083 3224 4087
tri 3224 4083 3228 4087 sw
tri 3292 4083 3296 4087 ne
rect 3296 4083 3366 4087
tri 3366 4083 3370 4087 sw
tri 3425 4083 3429 4087 ne
rect 3429 4083 3499 4087
tri 3499 4083 3503 4087 sw
rect 3161 4082 3228 4083
tri 3228 4082 3229 4083 sw
tri 3296 4082 3297 4083 ne
rect 3297 4082 3370 4083
tri 3370 4082 3371 4083 sw
tri 3429 4082 3430 4083 ne
rect 3430 4082 3503 4083
rect 3161 4076 3229 4082
tri 3229 4076 3235 4082 sw
tri 3297 4076 3303 4082 ne
rect 3303 4076 3371 4082
tri 3371 4076 3377 4082 sw
tri 3430 4076 3436 4082 ne
rect 3436 4076 3503 4082
tri 3503 4076 3510 4083 sw
tri 3161 4072 3165 4076 ne
rect 3165 4072 3235 4076
tri 3235 4072 3239 4076 sw
tri 3303 4072 3307 4076 ne
rect 3307 4072 3377 4076
tri 3377 4072 3381 4076 sw
tri 3436 4072 3440 4076 ne
rect 3440 4072 3510 4076
tri 3510 4072 3514 4076 sw
tri 3165 4067 3170 4072 ne
rect 3170 4067 3239 4072
rect -16 3991 -8 4043
rect 44 3991 56 4043
rect 108 3991 114 4043
rect 1621 4015 1627 4067
rect 1679 4015 1708 4067
rect 1760 4061 2884 4067
tri 2884 4061 2890 4067 sw
tri 3170 4061 3176 4067 ne
rect 3176 4061 3239 4067
rect 1760 4045 2890 4061
tri 2890 4045 2906 4061 sw
tri 3176 4045 3192 4061 ne
rect 3192 4045 3239 4061
tri 3239 4045 3266 4072 sw
tri 3307 4045 3334 4072 ne
rect 3334 4067 3381 4072
tri 3381 4067 3386 4072 sw
tri 3440 4067 3445 4072 ne
rect 3445 4067 3514 4072
rect 3334 4045 3386 4067
tri 3386 4045 3408 4067 sw
tri 3445 4045 3467 4067 ne
rect 3467 4045 3514 4067
tri 3514 4045 3541 4072 sw
rect 3884 4053 4126 4087
rect 4178 4053 4196 4087
rect 4248 4053 4266 4105
rect 4318 4053 4336 4105
rect 4388 4053 4406 4105
rect 4458 4053 4476 4105
rect 4533 4087 4540 4121
rect 4528 4053 4540 4087
rect 4762 4083 6268 4135
rect 6320 4083 6344 4135
rect 6396 4083 6966 4135
rect 8402 4083 8408 4135
rect 8460 4083 8472 4135
rect 8524 4083 8530 4135
rect 11227 4106 16390 4144
rect 3884 4045 4540 4053
rect 1760 4043 2906 4045
tri 2906 4043 2908 4045 sw
tri 3192 4043 3194 4045 ne
rect 3194 4043 3266 4045
tri 3266 4043 3268 4045 sw
tri 3334 4043 3336 4045 ne
rect 3336 4043 3408 4045
tri 3408 4043 3410 4045 sw
tri 3467 4043 3469 4045 ne
rect 3469 4043 3541 4045
tri 3541 4043 3543 4045 sw
rect 1760 4015 2908 4043
tri 2908 4015 2936 4043 sw
tri 3194 4015 3222 4043 ne
rect 3222 4015 3268 4043
tri 2862 4011 2866 4015 ne
rect 2866 4011 2936 4015
tri 2936 4011 2940 4015 sw
tri 3222 4011 3226 4015 ne
rect 3226 4014 3268 4015
tri 3268 4014 3297 4043 sw
tri 3336 4014 3365 4043 ne
rect 3365 4019 3410 4043
tri 3410 4019 3434 4043 sw
tri 3469 4019 3493 4043 ne
rect 3493 4019 3543 4043
tri 3543 4019 3567 4043 sw
rect 3365 4014 3434 4019
rect 3226 4011 3297 4014
tri 3297 4011 3300 4014 sw
tri 3365 4011 3368 4014 ne
rect 3368 4011 3434 4014
tri 3434 4011 3442 4019 sw
tri 3493 4011 3501 4019 ne
rect 3501 4011 3567 4019
tri 3567 4011 3575 4019 sw
rect 3884 4011 3891 4045
rect 3925 4011 3967 4045
rect 4001 4011 4043 4045
rect 4077 4011 4119 4045
rect 4153 4039 4195 4045
rect 4229 4039 4271 4045
rect 4305 4039 4347 4045
rect 4381 4039 4423 4045
rect 4457 4039 4499 4045
rect 4178 4011 4195 4039
tri 2866 4000 2877 4011 ne
rect 2877 4002 2940 4011
tri 2940 4002 2949 4011 sw
tri 3226 4002 3235 4011 ne
rect 3235 4008 3300 4011
tri 3300 4008 3303 4011 sw
tri 3368 4008 3371 4011 ne
rect 3371 4008 3442 4011
tri 3442 4008 3445 4011 sw
tri 3501 4008 3504 4011 ne
rect 3504 4008 3575 4011
rect 3235 4002 3303 4008
tri 3303 4002 3309 4008 sw
tri 3371 4002 3377 4008 ne
rect 3377 4002 3445 4008
tri 3445 4002 3451 4008 sw
tri 3504 4002 3510 4008 ne
rect 3510 4002 3575 4008
tri 3575 4002 3584 4011 sw
rect 2877 4000 2949 4002
tri 2949 4000 2951 4002 sw
tri 3235 4000 3237 4002 ne
rect 3237 4000 3309 4002
tri 3309 4000 3311 4002 sw
tri 3377 4000 3379 4002 ne
rect 3379 4000 3451 4002
tri 3451 4000 3453 4002 sw
tri 3510 4000 3512 4002 ne
rect 3512 4000 3584 4002
tri 3584 4000 3586 4002 sw
tri 2877 3991 2886 4000 ne
rect 2886 3991 2951 4000
tri 2951 3991 2960 4000 sw
tri 3237 3991 3246 4000 ne
rect 3246 3991 3311 4000
tri 3311 3991 3320 4000 sw
tri 3379 3991 3388 4000 ne
rect 3388 3993 3453 4000
tri 3453 3993 3460 4000 sw
tri 3512 3993 3519 4000 ne
rect 3519 3993 3586 4000
rect 3388 3991 3460 3993
tri 3460 3991 3462 3993 sw
tri 3519 3991 3521 3993 ne
rect 3521 3991 3586 3993
tri 3586 3991 3595 4000 sw
tri 2886 3987 2890 3991 ne
rect 2890 3987 2960 3991
tri 2960 3987 2964 3991 sw
tri 3246 3987 3250 3991 ne
rect 3250 3987 3320 3991
tri 2890 3968 2909 3987 ne
rect 2909 3968 2964 3987
tri 2964 3968 2983 3987 sw
tri 3250 3968 3269 3987 ne
rect 3269 3968 3320 3987
tri 3320 3968 3343 3991 sw
tri 3388 3968 3411 3991 ne
rect 3411 3968 3462 3991
tri 3462 3968 3485 3991 sw
tri 3521 3968 3544 3991 ne
rect 3544 3968 3595 3991
tri 3595 3968 3618 3991 sw
rect 3884 3987 4126 4011
rect 4178 3987 4196 4011
rect 4248 3987 4266 4039
rect 4318 3987 4336 4039
rect 4388 3987 4406 4039
rect 4458 3987 4476 4039
rect 4533 4011 4540 4045
rect 4528 3987 4540 4011
rect 3884 3973 4540 3987
rect 3884 3968 4126 3973
rect 4178 3968 4196 3973
tri 2909 3934 2943 3968 ne
rect 2943 3934 2983 3968
tri 2983 3934 3017 3968 sw
tri 3269 3934 3303 3968 ne
rect 3303 3940 3343 3968
tri 3343 3940 3371 3968 sw
tri 3411 3940 3439 3968 ne
rect 3439 3945 3485 3968
tri 3485 3945 3508 3968 sw
tri 3544 3945 3567 3968 ne
rect 3567 3945 3618 3968
tri 3618 3945 3641 3968 sw
rect 3439 3940 3508 3945
rect 3303 3934 3371 3940
tri 3371 3934 3377 3940 sw
tri 3439 3934 3445 3940 ne
rect 3445 3934 3508 3940
tri 3508 3934 3519 3945 sw
tri 3567 3934 3578 3945 ne
rect 3578 3934 3641 3945
tri 3641 3934 3652 3945 sw
rect 3884 3934 3891 3968
rect 3925 3934 3967 3968
rect 4001 3934 4043 3968
rect 4077 3934 4119 3968
rect 4178 3934 4195 3968
tri 2943 3928 2949 3934 ne
rect 2949 3928 3017 3934
tri 3017 3928 3023 3934 sw
tri 3303 3928 3309 3934 ne
rect 3309 3928 3377 3934
tri 3377 3928 3383 3934 sw
tri 3445 3928 3451 3934 ne
rect 3451 3928 3519 3934
tri 3519 3928 3525 3934 sw
tri 3578 3928 3584 3934 ne
rect 3584 3928 3652 3934
tri 3652 3928 3658 3934 sw
tri 2949 3913 2964 3928 ne
rect 2964 3913 3023 3928
tri 3023 3913 3038 3928 sw
tri 3309 3913 3324 3928 ne
rect 3324 3913 3383 3928
tri 2964 3891 2986 3913 ne
rect 2986 3891 3038 3913
tri 3038 3891 3060 3913 sw
tri 3324 3891 3346 3913 ne
rect 3346 3891 3383 3913
tri 3383 3891 3420 3928 sw
tri 3451 3891 3488 3928 ne
rect 3488 3919 3525 3928
tri 3525 3919 3534 3928 sw
tri 3584 3919 3593 3928 ne
rect 3593 3919 3658 3928
rect 3488 3891 3534 3919
tri 3534 3891 3562 3919 sw
tri 3593 3891 3621 3919 ne
rect 3621 3891 3658 3919
tri 3658 3891 3695 3928 sw
rect 3884 3921 4126 3934
rect 4178 3921 4196 3934
rect 4248 3921 4266 3973
rect 4318 3921 4336 3973
rect 4388 3921 4406 3973
rect 4458 3921 4476 3973
rect 4528 3968 4540 3973
rect 4533 3934 4540 3968
rect 4528 3921 4540 3934
rect 3884 3907 4540 3921
rect 3884 3891 4126 3907
rect 4178 3891 4196 3907
tri 2986 3857 3020 3891 ne
rect 3020 3857 3060 3891
tri 3060 3857 3094 3891 sw
tri 3346 3857 3380 3891 ne
rect 3380 3866 3420 3891
tri 3420 3866 3445 3891 sw
tri 3488 3866 3513 3891 ne
rect 3513 3871 3562 3891
tri 3562 3871 3582 3891 sw
tri 3621 3871 3641 3891 ne
rect 3641 3871 3695 3891
tri 3695 3871 3715 3891 sw
rect 3513 3866 3582 3871
rect 3380 3860 3445 3866
tri 3445 3860 3451 3866 sw
tri 3513 3860 3519 3866 ne
rect 3519 3860 3582 3866
tri 3582 3860 3593 3871 sw
tri 3641 3860 3652 3871 ne
rect 3652 3860 3715 3871
rect 3380 3857 3451 3860
tri 3451 3857 3454 3860 sw
tri 3519 3857 3522 3860 ne
rect 3522 3857 3593 3860
tri 3593 3857 3596 3860 sw
tri 3652 3857 3655 3860 ne
rect 3655 3857 3715 3860
tri 3715 3857 3729 3871 sw
rect 3884 3857 3891 3891
rect 3925 3857 3967 3891
rect 4001 3857 4043 3891
rect 4077 3857 4119 3891
rect 4178 3857 4195 3891
tri 3020 3856 3021 3857 ne
rect 3021 3856 3094 3857
tri 3094 3856 3095 3857 sw
tri 3380 3856 3381 3857 ne
rect 3381 3856 3454 3857
tri 3454 3856 3455 3857 sw
tri 3522 3856 3523 3857 ne
rect 3523 3856 3596 3857
tri 3596 3856 3597 3857 sw
tri 3655 3856 3656 3857 ne
rect 3656 3856 3729 3857
tri 3729 3856 3730 3857 sw
tri 3021 3839 3038 3856 ne
rect 3038 3854 3095 3856
tri 3095 3854 3097 3856 sw
tri 3381 3854 3383 3856 ne
rect 3383 3854 3455 3856
tri 3455 3854 3457 3856 sw
tri 3523 3854 3525 3856 ne
rect 3525 3854 3597 3856
tri 3597 3854 3599 3856 sw
tri 3656 3854 3658 3856 ne
rect 3658 3854 3730 3856
tri 3730 3854 3732 3856 sw
rect 3884 3855 4126 3857
rect 4178 3855 4196 3857
rect 4248 3855 4266 3907
rect 4318 3855 4336 3907
rect 4388 3855 4406 3907
rect 4458 3855 4476 3907
rect 4528 3891 4540 3907
rect 4533 3857 4540 3891
rect 4528 3855 4540 3857
rect 3038 3839 3097 3854
tri 3097 3839 3112 3854 sw
tri 3383 3839 3398 3854 ne
rect 3398 3839 3457 3854
tri 3038 3765 3112 3839 ne
tri 3112 3780 3171 3839 sw
tri 3398 3780 3457 3839 ne
tri 3457 3792 3519 3854 sw
tri 3525 3792 3587 3854 ne
rect 3587 3845 3599 3854
tri 3599 3845 3608 3854 sw
tri 3658 3845 3667 3854 ne
rect 3667 3845 3732 3854
rect 3587 3797 3608 3845
tri 3608 3797 3656 3845 sw
tri 3667 3797 3715 3845 ne
rect 3715 3797 3732 3845
tri 3732 3797 3789 3854 sw
rect 3884 3845 4540 3855
rect 11227 4072 11937 4106
rect 11971 4072 12010 4106
rect 12044 4072 12083 4106
rect 12117 4072 12156 4106
rect 12190 4072 12229 4106
rect 12263 4072 12302 4106
rect 12336 4072 12375 4106
rect 12409 4072 12448 4106
rect 12482 4072 12521 4106
rect 12555 4072 12594 4106
rect 12628 4072 12667 4106
rect 12701 4072 12740 4106
rect 12774 4072 12813 4106
rect 12847 4072 12886 4106
rect 12920 4072 12959 4106
rect 12993 4072 13032 4106
rect 13066 4072 13105 4106
rect 13139 4072 13178 4106
rect 13212 4072 13251 4106
rect 13285 4072 13324 4106
rect 13358 4072 13397 4106
rect 13431 4072 13470 4106
rect 13504 4072 13543 4106
rect 13577 4072 13616 4106
rect 13650 4072 13689 4106
rect 13723 4072 13762 4106
rect 13796 4072 13835 4106
rect 13869 4072 13908 4106
rect 13942 4072 13981 4106
rect 14015 4072 14054 4106
rect 14088 4072 14127 4106
rect 14161 4072 14200 4106
rect 14234 4072 14273 4106
rect 14307 4072 14346 4106
rect 14380 4072 14419 4106
rect 14453 4072 14492 4106
rect 14526 4072 14565 4106
rect 14599 4072 14638 4106
rect 14672 4072 14711 4106
rect 14745 4072 14784 4106
rect 14818 4072 14857 4106
rect 14891 4072 14930 4106
rect 14964 4072 15003 4106
rect 15037 4072 15076 4106
rect 15110 4072 15149 4106
rect 15183 4072 15222 4106
rect 15256 4072 15295 4106
rect 15329 4072 15368 4106
rect 15402 4072 15441 4106
rect 15475 4072 15514 4106
rect 15548 4072 15587 4106
rect 15621 4072 15660 4106
rect 15694 4072 15733 4106
rect 15767 4072 15806 4106
rect 15840 4072 15879 4106
rect 15913 4072 15952 4106
rect 15986 4072 16025 4106
rect 16059 4072 16098 4106
rect 16132 4072 16171 4106
rect 16205 4072 16244 4106
rect 16278 4072 16317 4106
rect 16351 4072 16390 4106
rect 11227 4034 16390 4072
rect 11227 4000 11937 4034
rect 11971 4000 12010 4034
rect 12044 4000 12083 4034
rect 12117 4000 12156 4034
rect 12190 4000 12229 4034
rect 12263 4000 12302 4034
rect 12336 4000 12375 4034
rect 12409 4000 12448 4034
rect 12482 4000 12521 4034
rect 12555 4000 12594 4034
rect 12628 4000 12667 4034
rect 12701 4000 12740 4034
rect 12774 4000 12813 4034
rect 12847 4000 12886 4034
rect 12920 4000 12959 4034
rect 12993 4000 13032 4034
rect 13066 4000 13105 4034
rect 13139 4000 13178 4034
rect 13212 4000 13251 4034
rect 13285 4000 13324 4034
rect 13358 4000 13397 4034
rect 13431 4000 13470 4034
rect 13504 4000 13543 4034
rect 13577 4000 13616 4034
rect 13650 4000 13689 4034
rect 13723 4000 13762 4034
rect 13796 4000 13835 4034
rect 13869 4000 13908 4034
rect 13942 4000 13981 4034
rect 14015 4000 14054 4034
rect 14088 4000 14127 4034
rect 14161 4000 14200 4034
rect 14234 4000 14273 4034
rect 14307 4000 14346 4034
rect 14380 4000 14419 4034
rect 14453 4000 14492 4034
rect 14526 4000 14565 4034
rect 14599 4000 14638 4034
rect 14672 4000 14711 4034
rect 14745 4000 14784 4034
rect 14818 4000 14857 4034
rect 14891 4000 14930 4034
rect 14964 4000 15003 4034
rect 15037 4000 15076 4034
rect 15110 4000 15149 4034
rect 15183 4000 15222 4034
rect 15256 4000 15295 4034
rect 15329 4000 15368 4034
rect 15402 4000 15441 4034
rect 15475 4000 15514 4034
rect 15548 4000 15587 4034
rect 15621 4000 15660 4034
rect 15694 4000 15733 4034
rect 15767 4000 15806 4034
rect 15840 4000 15879 4034
rect 15913 4000 15952 4034
rect 15986 4000 16025 4034
rect 16059 4000 16098 4034
rect 16132 4000 16171 4034
rect 16205 4000 16244 4034
rect 16278 4000 16317 4034
rect 16351 4000 16390 4034
rect 11227 3962 16390 4000
rect 11227 3928 11937 3962
rect 11971 3928 12010 3962
rect 12044 3928 12083 3962
rect 12117 3928 12156 3962
rect 12190 3928 12229 3962
rect 12263 3928 12302 3962
rect 12336 3928 12375 3962
rect 12409 3928 12448 3962
rect 12482 3928 12521 3962
rect 12555 3928 12594 3962
rect 12628 3928 12667 3962
rect 12701 3928 12740 3962
rect 12774 3928 12813 3962
rect 12847 3928 12886 3962
rect 12920 3928 12959 3962
rect 12993 3928 13032 3962
rect 13066 3928 13105 3962
rect 13139 3928 13178 3962
rect 13212 3928 13251 3962
rect 13285 3928 13324 3962
rect 13358 3928 13397 3962
rect 13431 3928 13470 3962
rect 13504 3928 13543 3962
rect 13577 3928 13616 3962
rect 13650 3928 13689 3962
rect 13723 3928 13762 3962
rect 13796 3928 13835 3962
rect 13869 3928 13908 3962
rect 13942 3928 13981 3962
rect 14015 3928 14054 3962
rect 14088 3928 14127 3962
rect 14161 3928 14200 3962
rect 14234 3928 14273 3962
rect 14307 3928 14346 3962
rect 14380 3928 14419 3962
rect 14453 3928 14492 3962
rect 14526 3928 14565 3962
rect 14599 3928 14638 3962
rect 14672 3928 14711 3962
rect 14745 3928 14784 3962
rect 14818 3928 14857 3962
rect 14891 3928 14930 3962
rect 14964 3928 15003 3962
rect 15037 3928 15076 3962
rect 15110 3928 15149 3962
rect 15183 3928 15222 3962
rect 15256 3928 15295 3962
rect 15329 3928 15368 3962
rect 15402 3928 15441 3962
rect 15475 3928 15514 3962
rect 15548 3928 15587 3962
rect 15621 3928 15660 3962
rect 15694 3928 15733 3962
rect 15767 3928 15806 3962
rect 15840 3928 15879 3962
rect 15913 3928 15952 3962
rect 15986 3928 16025 3962
rect 16059 3928 16098 3962
rect 16132 3928 16171 3962
rect 16205 3928 16244 3962
rect 16278 3928 16317 3962
rect 16351 3928 16390 3962
rect 11227 3890 16390 3928
rect 11227 3856 11937 3890
rect 11971 3856 12010 3890
rect 12044 3856 12083 3890
rect 12117 3856 12156 3890
rect 12190 3856 12229 3890
rect 12263 3856 12302 3890
rect 12336 3856 12375 3890
rect 12409 3856 12448 3890
rect 12482 3856 12521 3890
rect 12555 3856 12594 3890
rect 12628 3856 12667 3890
rect 12701 3856 12740 3890
rect 12774 3856 12813 3890
rect 12847 3856 12886 3890
rect 12920 3856 12959 3890
rect 12993 3856 13032 3890
rect 13066 3856 13105 3890
rect 13139 3856 13178 3890
rect 13212 3856 13251 3890
rect 13285 3856 13324 3890
rect 13358 3856 13397 3890
rect 13431 3856 13470 3890
rect 13504 3856 13543 3890
rect 13577 3856 13616 3890
rect 13650 3856 13689 3890
rect 13723 3856 13762 3890
rect 13796 3856 13835 3890
rect 13869 3856 13908 3890
rect 13942 3856 13981 3890
rect 14015 3856 14054 3890
rect 14088 3856 14127 3890
rect 14161 3856 14200 3890
rect 14234 3856 14273 3890
rect 14307 3856 14346 3890
rect 14380 3856 14419 3890
rect 14453 3856 14492 3890
rect 14526 3856 14565 3890
rect 14599 3856 14638 3890
rect 14672 3856 14711 3890
rect 14745 3856 14784 3890
rect 14818 3856 14857 3890
rect 14891 3856 14930 3890
rect 14964 3856 15003 3890
rect 15037 3856 15076 3890
rect 15110 3856 15149 3890
rect 15183 3856 15222 3890
rect 15256 3856 15295 3890
rect 15329 3856 15368 3890
rect 15402 3856 15441 3890
rect 15475 3856 15514 3890
rect 15548 3856 15587 3890
rect 15621 3856 15660 3890
rect 15694 3856 15733 3890
rect 15767 3856 15806 3890
rect 15840 3856 15879 3890
rect 15913 3856 15952 3890
rect 15986 3856 16025 3890
rect 16059 3856 16098 3890
rect 16132 3856 16171 3890
rect 16205 3856 16244 3890
rect 16278 3856 16317 3890
rect 16351 3856 16390 3890
rect 16928 3856 16940 4322
rect 3587 3792 3656 3797
rect 3457 3786 3519 3792
tri 3519 3786 3525 3792 sw
tri 3587 3786 3593 3792 ne
rect 3593 3786 3656 3792
tri 3656 3786 3667 3797 sw
tri 3715 3786 3726 3797 ne
rect 3726 3786 3789 3797
rect 3457 3780 3525 3786
tri 3525 3780 3531 3786 sw
tri 3593 3780 3599 3786 ne
rect 3599 3780 3667 3786
tri 3667 3780 3673 3786 sw
tri 3726 3780 3732 3786 ne
rect 3732 3780 3789 3786
tri 3789 3780 3806 3797 sw
rect 3112 3765 3171 3780
tri 3171 3765 3186 3780 sw
tri 3457 3765 3472 3780 ne
rect 3472 3765 3531 3780
tri 3112 3691 3186 3765 ne
tri 3186 3706 3245 3765 sw
tri 3472 3706 3531 3765 ne
tri 3531 3718 3593 3780 sw
tri 3599 3718 3661 3780 ne
rect 3661 3771 3673 3780
tri 3673 3771 3682 3780 sw
tri 3732 3771 3741 3780 ne
rect 3741 3771 3806 3780
rect 3661 3723 3682 3771
tri 3682 3723 3730 3771 sw
tri 3741 3723 3789 3771 ne
rect 3789 3723 3806 3771
tri 3806 3723 3863 3780 sw
rect 3661 3718 3730 3723
rect 3531 3712 3593 3718
tri 3593 3712 3599 3718 sw
tri 3661 3712 3667 3718 ne
rect 3667 3712 3730 3718
tri 3730 3712 3741 3723 sw
tri 3789 3712 3800 3723 ne
rect 3800 3712 3863 3723
rect 3531 3706 3599 3712
tri 3599 3706 3605 3712 sw
tri 3667 3706 3673 3712 ne
rect 3673 3706 3741 3712
tri 3741 3706 3747 3712 sw
tri 3800 3706 3806 3712 ne
rect 3806 3706 3863 3712
tri 3863 3706 3880 3723 sw
rect 3186 3691 3245 3706
tri 3245 3691 3260 3706 sw
tri 3531 3691 3546 3706 ne
rect 3546 3691 3605 3706
tri 3186 3617 3260 3691 ne
tri 3260 3632 3319 3691 sw
tri 3546 3632 3605 3691 ne
tri 3605 3661 3650 3706 sw
tri 3673 3661 3718 3706 ne
rect 3718 3697 3747 3706
tri 3747 3697 3756 3706 sw
tri 3806 3697 3815 3706 ne
rect 3815 3697 3880 3706
rect 3718 3661 3756 3697
tri 3756 3661 3792 3697 sw
tri 3815 3661 3851 3697 ne
rect 3851 3661 3880 3697
tri 3880 3661 3925 3706 sw
rect 3605 3644 3650 3661
tri 3650 3644 3667 3661 sw
tri 3718 3644 3735 3661 ne
rect 3735 3649 3792 3661
tri 3792 3649 3804 3661 sw
tri 3851 3649 3863 3661 ne
rect 3863 3649 3925 3661
tri 3925 3649 3937 3661 sw
rect 3735 3644 3804 3649
rect 3605 3638 3667 3644
tri 3667 3638 3673 3644 sw
tri 3735 3638 3741 3644 ne
rect 3741 3638 3804 3644
tri 3804 3638 3815 3649 sw
tri 3863 3638 3874 3649 ne
rect 3874 3638 3937 3649
rect 3605 3632 3673 3638
tri 3673 3632 3679 3638 sw
tri 3741 3632 3747 3638 ne
rect 3747 3632 3815 3638
tri 3815 3632 3821 3638 sw
tri 3874 3632 3880 3638 ne
rect 3880 3632 3937 3638
tri 3937 3632 3954 3649 sw
rect 3260 3617 3319 3632
tri 3319 3617 3334 3632 sw
tri 3605 3617 3620 3632 ne
rect 3620 3617 3679 3632
tri 3260 3609 3268 3617 ne
rect 3268 3609 3334 3617
tri 3334 3609 3342 3617 sw
tri 3620 3609 3628 3617 ne
rect 3628 3609 3679 3617
tri 3679 3609 3702 3632 sw
tri 3747 3609 3770 3632 ne
rect 3770 3623 3821 3632
tri 3821 3623 3830 3632 sw
tri 3880 3623 3889 3632 ne
rect 3889 3623 3954 3632
rect 3770 3609 3830 3623
tri 3830 3609 3844 3623 sw
tri 3889 3609 3903 3623 ne
rect 3903 3609 3954 3623
tri 3954 3609 3977 3632 sw
rect 6313 3609 6319 3661
rect 6371 3609 6383 3661
rect 6435 3609 9392 3661
rect 9444 3609 9456 3661
rect 9508 3609 9514 3661
rect 11227 3609 16940 3856
tri 3268 3575 3302 3609 ne
rect 3302 3575 3342 3609
tri 3342 3575 3376 3609 sw
tri 3628 3575 3662 3609 ne
rect 3662 3575 3702 3609
tri 3702 3575 3736 3609 sw
tri 3770 3575 3804 3609 ne
rect 3804 3575 3844 3609
tri 3844 3575 3878 3609 sw
tri 3903 3575 3937 3609 ne
rect 3937 3575 3977 3609
tri 3977 3575 4011 3609 sw
rect 11227 3575 11953 3609
rect 11987 3575 12026 3609
rect 12060 3575 12099 3609
rect 12133 3575 12172 3609
rect 12206 3575 12245 3609
rect 12279 3575 12318 3609
rect 12352 3575 12391 3609
rect 12425 3575 12464 3609
rect 12498 3575 12537 3609
rect 12571 3575 12610 3609
rect 12644 3575 12683 3609
rect 12717 3575 12756 3609
rect 12790 3575 12829 3609
rect 12863 3575 12902 3609
rect 12936 3575 12975 3609
rect 13009 3575 13048 3609
rect 13082 3575 13121 3609
rect 13155 3575 13194 3609
rect 13228 3575 13267 3609
rect 13301 3575 13340 3609
rect 13374 3575 13413 3609
rect 13447 3575 13486 3609
rect 13520 3575 13559 3609
rect 13593 3575 13632 3609
rect 13666 3575 13705 3609
rect 13739 3575 13778 3609
rect 13812 3575 13851 3609
rect 13885 3575 13924 3609
rect 13958 3575 13997 3609
rect 14031 3575 14070 3609
rect 14104 3575 14143 3609
rect 14177 3575 14216 3609
rect 14250 3575 14289 3609
rect 14323 3575 14362 3609
rect 14396 3575 14435 3609
rect 14469 3575 14508 3609
rect 14542 3575 14581 3609
rect 14615 3575 14654 3609
rect 14688 3575 14727 3609
rect 14761 3575 14800 3609
rect 14834 3575 14873 3609
rect 14907 3575 14946 3609
rect 14980 3575 15019 3609
rect 15053 3575 15092 3609
rect 15126 3575 15165 3609
rect 15199 3575 15238 3609
rect 15272 3575 15311 3609
rect 15345 3575 15384 3609
rect 15418 3575 15457 3609
rect 15491 3575 15530 3609
rect 15564 3575 15603 3609
rect 15637 3575 15676 3609
rect 15710 3575 15749 3609
rect 15783 3575 15822 3609
rect 15856 3575 15895 3609
rect 15929 3575 15968 3609
rect 16002 3575 16041 3609
rect 16075 3575 16114 3609
rect 16148 3575 16187 3609
rect 16221 3575 16260 3609
rect 16294 3575 16333 3609
rect 16367 3575 16406 3609
tri 3302 3543 3334 3575 ne
rect 3334 3558 3376 3575
tri 3376 3558 3393 3575 sw
tri 3662 3558 3679 3575 ne
rect 3679 3570 3736 3575
tri 3736 3570 3741 3575 sw
tri 3804 3570 3809 3575 ne
rect 3809 3570 3878 3575
rect 3679 3564 3741 3570
tri 3741 3564 3747 3570 sw
tri 3809 3564 3815 3570 ne
rect 3815 3564 3878 3570
tri 3878 3564 3889 3575 sw
tri 3937 3564 3948 3575 ne
rect 3948 3564 8240 3575
rect 3679 3558 3747 3564
tri 3747 3558 3753 3564 sw
tri 3815 3558 3821 3564 ne
rect 3821 3558 3889 3564
tri 3889 3558 3895 3564 sw
tri 3948 3558 3954 3564 ne
rect 3954 3558 8240 3564
rect 3334 3543 3393 3558
tri 3393 3543 3408 3558 sw
tri 3679 3543 3694 3558 ne
rect 3694 3543 3753 3558
tri 3334 3537 3340 3543 ne
rect 3340 3537 3408 3543
tri 3408 3537 3414 3543 sw
tri 3694 3537 3700 3543 ne
rect 3700 3537 3753 3543
tri 3753 3537 3774 3558 sw
tri 3821 3537 3842 3558 ne
rect 3842 3549 3895 3558
tri 3895 3549 3904 3558 sw
tri 3954 3549 3963 3558 ne
rect 3963 3549 8240 3558
rect 3842 3537 3904 3549
tri 3904 3537 3916 3549 sw
tri 3963 3537 3975 3549 ne
rect 3975 3537 8240 3549
tri 3340 3503 3374 3537 ne
rect 3374 3503 3414 3537
tri 3414 3503 3448 3537 sw
tri 3700 3503 3734 3537 ne
rect 3734 3523 3774 3537
tri 3774 3523 3788 3537 sw
tri 3842 3523 3856 3537 ne
rect 3856 3523 3916 3537
tri 3916 3523 3930 3537 sw
tri 3975 3523 3989 3537 ne
rect 3989 3523 8240 3537
rect 8292 3523 8304 3575
rect 8356 3523 8362 3575
rect 11227 3537 16406 3575
rect 3734 3503 3788 3523
tri 3788 3503 3808 3523 sw
tri 3856 3503 3876 3523 ne
rect 3876 3503 3930 3523
tri 3930 3503 3950 3523 sw
rect 11227 3503 11953 3537
rect 11987 3503 12026 3537
rect 12060 3503 12099 3537
rect 12133 3503 12172 3537
rect 12206 3503 12245 3537
rect 12279 3503 12318 3537
rect 12352 3503 12391 3537
rect 12425 3503 12464 3537
rect 12498 3503 12537 3537
rect 12571 3503 12610 3537
rect 12644 3503 12683 3537
rect 12717 3503 12756 3537
rect 12790 3503 12829 3537
rect 12863 3503 12902 3537
rect 12936 3503 12975 3537
rect 13009 3503 13048 3537
rect 13082 3503 13121 3537
rect 13155 3503 13194 3537
rect 13228 3503 13267 3537
rect 13301 3503 13340 3537
rect 13374 3503 13413 3537
rect 13447 3503 13486 3537
rect 13520 3503 13559 3537
rect 13593 3503 13632 3537
rect 13666 3503 13705 3537
rect 13739 3503 13778 3537
rect 13812 3503 13851 3537
rect 13885 3503 13924 3537
rect 13958 3503 13997 3537
rect 14031 3503 14070 3537
rect 14104 3503 14143 3537
rect 14177 3503 14216 3537
rect 14250 3503 14289 3537
rect 14323 3503 14362 3537
rect 14396 3503 14435 3537
rect 14469 3503 14508 3537
rect 14542 3503 14581 3537
rect 14615 3503 14654 3537
rect 14688 3503 14727 3537
rect 14761 3503 14800 3537
rect 14834 3503 14873 3537
rect 14907 3503 14946 3537
rect 14980 3503 15019 3537
rect 15053 3503 15092 3537
rect 15126 3503 15165 3537
rect 15199 3503 15238 3537
rect 15272 3503 15311 3537
rect 15345 3503 15384 3537
rect 15418 3503 15457 3537
rect 15491 3503 15530 3537
rect 15564 3503 15603 3537
rect 15637 3503 15676 3537
rect 15710 3503 15749 3537
rect 15783 3503 15822 3537
rect 15856 3503 15895 3537
rect 15929 3503 15968 3537
rect 16002 3503 16041 3537
rect 16075 3503 16114 3537
rect 16148 3503 16187 3537
rect 16221 3503 16260 3537
rect 16294 3503 16333 3537
rect 16367 3503 16406 3537
tri 3374 3469 3408 3503 ne
rect 3408 3484 3448 3503
tri 3448 3484 3467 3503 sw
tri 3734 3484 3753 3503 ne
rect 3753 3496 3808 3503
tri 3808 3496 3815 3503 sw
tri 3876 3496 3883 3503 ne
rect 3883 3496 3950 3503
rect 3753 3490 3815 3496
tri 3815 3490 3821 3496 sw
tri 3883 3490 3889 3496 ne
rect 3889 3490 3950 3496
tri 3950 3490 3963 3503 sw
rect 3753 3484 3821 3490
tri 3821 3484 3827 3490 sw
tri 3889 3484 3895 3490 ne
rect 3895 3484 10440 3490
rect 3408 3469 3467 3484
tri 3467 3469 3482 3484 sw
tri 3753 3469 3768 3484 ne
rect 3768 3469 3827 3484
tri 3408 3465 3412 3469 ne
rect 3412 3465 3482 3469
tri 3482 3465 3486 3469 sw
tri 3768 3465 3772 3469 ne
rect 3772 3465 3827 3469
tri 3827 3465 3846 3484 sw
tri 3895 3465 3914 3484 ne
rect 3914 3465 10440 3484
tri 3412 3431 3446 3465 ne
rect 3446 3431 3486 3465
tri 3486 3431 3520 3465 sw
tri 3772 3431 3806 3465 ne
rect 3806 3438 3846 3465
tri 3846 3438 3873 3465 sw
tri 3914 3438 3941 3465 ne
rect 3941 3438 10440 3465
rect 10492 3438 10504 3490
rect 10556 3438 10562 3490
rect 11227 3465 16406 3503
rect 3806 3431 3873 3438
tri 3873 3431 3880 3438 sw
rect 11227 3431 11953 3465
rect 11987 3431 12026 3465
rect 12060 3431 12099 3465
rect 12133 3431 12172 3465
rect 12206 3431 12245 3465
rect 12279 3431 12318 3465
rect 12352 3431 12391 3465
rect 12425 3431 12464 3465
rect 12498 3431 12537 3465
rect 12571 3431 12610 3465
rect 12644 3431 12683 3465
rect 12717 3431 12756 3465
rect 12790 3431 12829 3465
rect 12863 3431 12902 3465
rect 12936 3431 12975 3465
rect 13009 3431 13048 3465
rect 13082 3431 13121 3465
rect 13155 3431 13194 3465
rect 13228 3431 13267 3465
rect 13301 3431 13340 3465
rect 13374 3431 13413 3465
rect 13447 3431 13486 3465
rect 13520 3431 13559 3465
rect 13593 3431 13632 3465
rect 13666 3431 13705 3465
rect 13739 3431 13778 3465
rect 13812 3431 13851 3465
rect 13885 3431 13924 3465
rect 13958 3431 13997 3465
rect 14031 3431 14070 3465
rect 14104 3431 14143 3465
rect 14177 3431 14216 3465
rect 14250 3431 14289 3465
rect 14323 3431 14362 3465
rect 14396 3431 14435 3465
rect 14469 3431 14508 3465
rect 14542 3431 14581 3465
rect 14615 3431 14654 3465
rect 14688 3431 14727 3465
rect 14761 3431 14800 3465
rect 14834 3431 14873 3465
rect 14907 3431 14946 3465
rect 14980 3431 15019 3465
rect 15053 3431 15092 3465
rect 15126 3431 15165 3465
rect 15199 3431 15238 3465
rect 15272 3431 15311 3465
rect 15345 3431 15384 3465
rect 15418 3431 15457 3465
rect 15491 3431 15530 3465
rect 15564 3431 15603 3465
rect 15637 3431 15676 3465
rect 15710 3431 15749 3465
rect 15783 3431 15822 3465
rect 15856 3431 15895 3465
rect 15929 3431 15968 3465
rect 16002 3431 16041 3465
rect 16075 3431 16114 3465
rect 16148 3431 16187 3465
rect 16221 3431 16260 3465
rect 16294 3431 16333 3465
rect 16367 3431 16406 3465
tri 3446 3425 3452 3431 ne
rect 3452 3425 3520 3431
tri 3520 3425 3526 3431 sw
tri 3806 3425 3812 3431 ne
rect 3812 3425 3880 3431
tri 3880 3425 3886 3431 sw
rect -3049 3419 -203 3425
rect -2997 3397 -203 3419
rect -2997 3374 -2971 3397
tri -2971 3374 -2948 3397 nw
tri -233 3374 -210 3397 ne
rect -210 3374 -203 3397
rect -2997 3373 -2972 3374
tri -2972 3373 -2971 3374 nw
tri -210 3373 -209 3374 ne
rect -209 3373 -203 3374
rect -151 3373 -139 3425
rect -87 3373 -81 3425
tri 3452 3420 3457 3425 ne
rect 3457 3420 3526 3425
tri 3526 3420 3531 3425 sw
tri 3812 3420 3817 3425 ne
rect 3817 3420 3886 3425
tri 3886 3420 3891 3425 sw
rect 39 3410 91 3420
tri 3457 3416 3461 3420 ne
rect 3461 3416 3531 3420
tri 3531 3416 3535 3420 sw
tri 3817 3416 3821 3420 ne
rect 3821 3416 3891 3420
tri 3891 3416 3895 3420 sw
tri 3461 3395 3482 3416 ne
rect 3482 3410 3535 3416
tri 3535 3410 3541 3416 sw
tri 3821 3410 3827 3416 ne
rect 3827 3410 3895 3416
tri 3895 3410 3901 3416 sw
rect 3482 3395 3541 3410
tri 3541 3395 3556 3410 sw
tri 3827 3395 3842 3410 ne
rect 3842 3395 6330 3410
tri 3482 3393 3484 3395 ne
rect 3484 3393 3556 3395
tri 3556 3393 3558 3395 sw
tri 3842 3393 3844 3395 ne
rect 3844 3393 6330 3395
rect -2997 3367 -2986 3373
rect -3049 3359 -2986 3367
tri -2986 3359 -2972 3373 nw
rect -3049 3355 -2997 3359
tri -2997 3348 -2986 3359 nw
tri 3484 3359 3518 3393 ne
rect 3518 3359 3558 3393
tri 3558 3359 3592 3393 sw
tri 3844 3359 3878 3393 ne
rect 3878 3359 6330 3393
rect -3049 3297 -2997 3303
rect 39 3346 91 3358
tri 3518 3321 3556 3359 ne
rect 3556 3358 3592 3359
tri 3592 3358 3593 3359 sw
tri 3878 3358 3879 3359 ne
rect 3879 3358 6330 3359
rect 6382 3358 6394 3410
rect 6446 3358 6452 3410
rect 11227 3393 16406 3431
rect 11227 3359 11953 3393
rect 11987 3359 12026 3393
rect 12060 3359 12099 3393
rect 12133 3359 12172 3393
rect 12206 3359 12245 3393
rect 12279 3359 12318 3393
rect 12352 3359 12391 3393
rect 12425 3359 12464 3393
rect 12498 3359 12537 3393
rect 12571 3359 12610 3393
rect 12644 3359 12683 3393
rect 12717 3359 12756 3393
rect 12790 3359 12829 3393
rect 12863 3359 12902 3393
rect 12936 3359 12975 3393
rect 13009 3359 13048 3393
rect 13082 3359 13121 3393
rect 13155 3359 13194 3393
rect 13228 3359 13267 3393
rect 13301 3359 13340 3393
rect 13374 3359 13413 3393
rect 13447 3359 13486 3393
rect 13520 3359 13559 3393
rect 13593 3359 13632 3393
rect 13666 3359 13705 3393
rect 13739 3359 13778 3393
rect 13812 3359 13851 3393
rect 13885 3359 13924 3393
rect 13958 3359 13997 3393
rect 14031 3359 14070 3393
rect 14104 3359 14143 3393
rect 14177 3359 14216 3393
rect 14250 3359 14289 3393
rect 14323 3359 14362 3393
rect 14396 3359 14435 3393
rect 14469 3359 14508 3393
rect 14542 3359 14581 3393
rect 14615 3359 14654 3393
rect 14688 3359 14727 3393
rect 14761 3359 14800 3393
rect 14834 3359 14873 3393
rect 14907 3359 14946 3393
rect 14980 3359 15019 3393
rect 15053 3359 15092 3393
rect 15126 3359 15165 3393
rect 15199 3359 15238 3393
rect 15272 3359 15311 3393
rect 15345 3359 15384 3393
rect 15418 3359 15457 3393
rect 15491 3359 15530 3393
rect 15564 3359 15603 3393
rect 15637 3359 15676 3393
rect 15710 3359 15749 3393
rect 15783 3359 15822 3393
rect 15856 3359 15895 3393
rect 15929 3359 15968 3393
rect 16002 3359 16041 3393
rect 16075 3359 16114 3393
rect 16148 3359 16187 3393
rect 16221 3359 16260 3393
rect 16294 3359 16333 3393
rect 16367 3359 16406 3393
rect 3556 3321 3593 3358
tri 3593 3321 3630 3358 sw
rect 11227 3321 16406 3359
rect 39 3288 91 3294
tri 3556 3288 3589 3321 ne
rect 3589 3288 3630 3321
tri 3630 3288 3663 3321 sw
tri 3589 3287 3590 3288 ne
rect 3590 3287 3663 3288
tri 3663 3287 3664 3288 sw
rect 11227 3287 11953 3321
rect 11987 3287 12026 3321
rect 12060 3287 12099 3321
rect 12133 3287 12172 3321
rect 12206 3287 12245 3321
rect 12279 3287 12318 3321
rect 12352 3287 12391 3321
rect 12425 3287 12464 3321
rect 12498 3287 12537 3321
rect 12571 3287 12610 3321
rect 12644 3287 12683 3321
rect 12717 3287 12756 3321
rect 12790 3287 12829 3321
rect 12863 3287 12902 3321
rect 12936 3287 12975 3321
rect 13009 3287 13048 3321
rect 13082 3287 13121 3321
rect 13155 3287 13194 3321
rect 13228 3287 13267 3321
rect 13301 3287 13340 3321
rect 13374 3287 13413 3321
rect 13447 3287 13486 3321
rect 13520 3287 13559 3321
rect 13593 3287 13632 3321
rect 13666 3287 13705 3321
rect 13739 3287 13778 3321
rect 13812 3287 13851 3321
rect 13885 3287 13924 3321
rect 13958 3287 13997 3321
rect 14031 3287 14070 3321
rect 14104 3287 14143 3321
rect 14177 3287 14216 3321
rect 14250 3287 14289 3321
rect 14323 3287 14362 3321
rect 14396 3287 14435 3321
rect 14469 3287 14508 3321
rect 14542 3287 14581 3321
rect 14615 3287 14654 3321
rect 14688 3287 14727 3321
rect 14761 3287 14800 3321
rect 14834 3287 14873 3321
rect 14907 3287 14946 3321
rect 14980 3287 15019 3321
rect 15053 3287 15092 3321
rect 15126 3287 15165 3321
rect 15199 3287 15238 3321
rect 15272 3287 15311 3321
rect 15345 3287 15384 3321
rect 15418 3287 15457 3321
rect 15491 3287 15530 3321
rect 15564 3287 15603 3321
rect 15637 3287 15676 3321
rect 15710 3287 15749 3321
rect 15783 3287 15822 3321
rect 15856 3287 15895 3321
rect 15929 3287 15968 3321
rect 16002 3287 16041 3321
rect 16075 3287 16114 3321
rect 16148 3287 16187 3321
rect 16221 3287 16260 3321
rect 16294 3287 16333 3321
rect 16367 3287 16406 3321
tri 3590 3249 3628 3287 ne
rect 3628 3249 3664 3287
tri 3664 3249 3702 3287 sw
rect 11227 3249 16406 3287
tri 3628 3247 3630 3249 ne
rect 3630 3247 3702 3249
tri 3702 3247 3704 3249 sw
tri 3630 3215 3662 3247 ne
rect 3662 3215 3704 3247
tri 3704 3215 3736 3247 sw
rect 11227 3215 11953 3249
rect 11987 3215 12026 3249
rect 12060 3215 12099 3249
rect 12133 3215 12172 3249
rect 12206 3215 12245 3249
rect 12279 3215 12318 3249
rect 12352 3215 12391 3249
rect 12425 3215 12464 3249
rect 12498 3215 12537 3249
rect 12571 3215 12610 3249
rect 12644 3215 12683 3249
rect 12717 3215 12756 3249
rect 12790 3215 12829 3249
rect 12863 3215 12902 3249
rect 12936 3215 12975 3249
rect 13009 3215 13048 3249
rect 13082 3215 13121 3249
rect 13155 3215 13194 3249
rect 13228 3215 13267 3249
rect 13301 3215 13340 3249
rect 13374 3215 13413 3249
rect 13447 3215 13486 3249
rect 13520 3215 13559 3249
rect 13593 3215 13632 3249
rect 13666 3215 13705 3249
rect 13739 3215 13778 3249
rect 13812 3215 13851 3249
rect 13885 3215 13924 3249
rect 13958 3215 13997 3249
rect 14031 3215 14070 3249
rect 14104 3215 14143 3249
rect 14177 3215 14216 3249
rect 14250 3215 14289 3249
rect 14323 3215 14362 3249
rect 14396 3215 14435 3249
rect 14469 3215 14508 3249
rect 14542 3215 14581 3249
rect 14615 3215 14654 3249
rect 14688 3215 14727 3249
rect 14761 3215 14800 3249
rect 14834 3215 14873 3249
rect 14907 3215 14946 3249
rect 14980 3215 15019 3249
rect 15053 3215 15092 3249
rect 15126 3215 15165 3249
rect 15199 3215 15238 3249
rect 15272 3215 15311 3249
rect 15345 3215 15384 3249
rect 15418 3215 15457 3249
rect 15491 3215 15530 3249
rect 15564 3215 15603 3249
rect 15637 3215 15676 3249
rect 15710 3215 15749 3249
rect 15783 3215 15822 3249
rect 15856 3215 15895 3249
rect 15929 3215 15968 3249
rect 16002 3215 16041 3249
rect 16075 3215 16114 3249
rect 16148 3215 16187 3249
rect 16221 3215 16260 3249
rect 16294 3215 16333 3249
rect 16367 3215 16406 3249
tri 3662 3177 3700 3215 ne
rect 3700 3177 3736 3215
tri 3736 3177 3774 3215 sw
rect 11227 3177 16406 3215
tri 3700 3173 3704 3177 ne
rect 3704 3173 3774 3177
tri 3774 3173 3778 3177 sw
tri 3704 3143 3734 3173 ne
rect 3734 3143 9195 3173
tri 3734 3121 3756 3143 ne
rect 3756 3121 9195 3143
rect 9247 3121 9259 3173
rect 9311 3121 9317 3173
rect 11227 3143 11953 3177
rect 11987 3143 12026 3177
rect 12060 3143 12099 3177
rect 12133 3143 12172 3177
rect 12206 3143 12245 3177
rect 12279 3143 12318 3177
rect 12352 3143 12391 3177
rect 12425 3143 12464 3177
rect 12498 3143 12537 3177
rect 12571 3143 12610 3177
rect 12644 3143 12683 3177
rect 12717 3143 12756 3177
rect 12790 3143 12829 3177
rect 12863 3143 12902 3177
rect 12936 3143 12975 3177
rect 13009 3143 13048 3177
rect 13082 3143 13121 3177
rect 13155 3143 13194 3177
rect 13228 3143 13267 3177
rect 13301 3143 13340 3177
rect 13374 3143 13413 3177
rect 13447 3143 13486 3177
rect 13520 3143 13559 3177
rect 13593 3143 13632 3177
rect 13666 3143 13705 3177
rect 13739 3143 13778 3177
rect 13812 3143 13851 3177
rect 13885 3143 13924 3177
rect 13958 3143 13997 3177
rect 14031 3143 14070 3177
rect 14104 3143 14143 3177
rect 14177 3143 14216 3177
rect 14250 3143 14289 3177
rect 14323 3143 14362 3177
rect 14396 3143 14435 3177
rect 14469 3143 14508 3177
rect 14542 3143 14581 3177
rect 14615 3143 14654 3177
rect 14688 3143 14727 3177
rect 14761 3143 14800 3177
rect 14834 3143 14873 3177
rect 14907 3143 14946 3177
rect 14980 3143 15019 3177
rect 15053 3143 15092 3177
rect 15126 3143 15165 3177
rect 15199 3143 15238 3177
rect 15272 3143 15311 3177
rect 15345 3143 15384 3177
rect 15418 3143 15457 3177
rect 15491 3143 15530 3177
rect 15564 3143 15603 3177
rect 15637 3143 15676 3177
rect 15710 3143 15749 3177
rect 15783 3143 15822 3177
rect 15856 3143 15895 3177
rect 15929 3143 15968 3177
rect 16002 3143 16041 3177
rect 16075 3143 16114 3177
rect 16148 3143 16187 3177
rect 16221 3143 16260 3177
rect 16294 3143 16333 3177
rect 16367 3143 16406 3177
rect 11227 3105 16406 3143
rect 11227 3071 11953 3105
rect 11987 3071 12026 3105
rect 12060 3071 12099 3105
rect 12133 3071 12172 3105
rect 12206 3071 12245 3105
rect 12279 3071 12318 3105
rect 12352 3071 12391 3105
rect 12425 3071 12464 3105
rect 12498 3071 12537 3105
rect 12571 3071 12610 3105
rect 12644 3071 12683 3105
rect 12717 3071 12756 3105
rect 12790 3071 12829 3105
rect 12863 3071 12902 3105
rect 12936 3071 12975 3105
rect 13009 3071 13048 3105
rect 13082 3071 13121 3105
rect 13155 3071 13194 3105
rect 13228 3071 13267 3105
rect 13301 3071 13340 3105
rect 13374 3071 13413 3105
rect 13447 3071 13486 3105
rect 13520 3071 13559 3105
rect 13593 3071 13632 3105
rect 13666 3071 13705 3105
rect 13739 3071 13778 3105
rect 13812 3071 13851 3105
rect 13885 3071 13924 3105
rect 13958 3071 13997 3105
rect 14031 3071 14070 3105
rect 14104 3071 14143 3105
rect 14177 3071 14216 3105
rect 14250 3071 14289 3105
rect 14323 3071 14362 3105
rect 14396 3071 14435 3105
rect 14469 3071 14508 3105
rect 14542 3071 14581 3105
rect 14615 3071 14654 3105
rect 14688 3071 14727 3105
rect 14761 3071 14800 3105
rect 14834 3071 14873 3105
rect 14907 3071 14946 3105
rect 14980 3071 15019 3105
rect 15053 3071 15092 3105
rect 15126 3071 15165 3105
rect 15199 3071 15238 3105
rect 15272 3071 15311 3105
rect 15345 3071 15384 3105
rect 15418 3071 15457 3105
rect 15491 3071 15530 3105
rect 15564 3071 15603 3105
rect 15637 3071 15676 3105
rect 15710 3071 15749 3105
rect 15783 3071 15822 3105
rect 15856 3071 15895 3105
rect 15929 3071 15968 3105
rect 16002 3071 16041 3105
rect 16075 3071 16114 3105
rect 16148 3071 16187 3105
rect 16221 3071 16260 3105
rect 16294 3071 16333 3105
rect 16367 3071 16406 3105
rect 11227 3033 16406 3071
rect 11227 2999 11953 3033
rect 11987 2999 12026 3033
rect 12060 2999 12099 3033
rect 12133 2999 12172 3033
rect 12206 2999 12245 3033
rect 12279 2999 12318 3033
rect 12352 2999 12391 3033
rect 12425 2999 12464 3033
rect 12498 2999 12537 3033
rect 12571 2999 12610 3033
rect 12644 2999 12683 3033
rect 12717 2999 12756 3033
rect 12790 2999 12829 3033
rect 12863 2999 12902 3033
rect 12936 2999 12975 3033
rect 13009 2999 13048 3033
rect 13082 2999 13121 3033
rect 13155 2999 13194 3033
rect 13228 2999 13267 3033
rect 13301 2999 13340 3033
rect 13374 2999 13413 3033
rect 13447 2999 13486 3033
rect 13520 2999 13559 3033
rect 13593 2999 13632 3033
rect 13666 2999 13705 3033
rect 13739 2999 13778 3033
rect 13812 2999 13851 3033
rect 13885 2999 13924 3033
rect 13958 2999 13997 3033
rect 14031 2999 14070 3033
rect 14104 2999 14143 3033
rect 14177 2999 14216 3033
rect 14250 2999 14289 3033
rect 14323 2999 14362 3033
rect 14396 2999 14435 3033
rect 14469 2999 14508 3033
rect 14542 2999 14581 3033
rect 14615 2999 14654 3033
rect 14688 2999 14727 3033
rect 14761 2999 14800 3033
rect 14834 2999 14873 3033
rect 14907 2999 14946 3033
rect 14980 2999 15019 3033
rect 15053 2999 15092 3033
rect 15126 2999 15165 3033
rect 15199 2999 15238 3033
rect 15272 2999 15311 3033
rect 15345 2999 15384 3033
rect 15418 2999 15457 3033
rect 15491 2999 15530 3033
rect 15564 2999 15603 3033
rect 15637 2999 15676 3033
rect 15710 2999 15749 3033
rect 15783 2999 15822 3033
rect 15856 2999 15895 3033
rect 15929 2999 15968 3033
rect 16002 2999 16041 3033
rect 16075 2999 16114 3033
rect 16148 2999 16187 3033
rect 16221 2999 16260 3033
rect 16294 2999 16333 3033
rect 16367 2999 16406 3033
rect 16872 2999 16940 3609
rect 11227 2959 16940 2999
tri 11229 2903 11285 2959 ne
tri 11224 2722 11285 2783 se
rect 11285 2722 11470 2959
tri 11470 2903 11526 2959 nw
tri 11829 2903 11885 2959 ne
tri 11470 2722 11531 2783 sw
tri 11824 2722 11885 2783 se
rect 11885 2722 12070 2959
tri 12070 2903 12126 2959 nw
tri 12429 2903 12485 2959 ne
tri 12070 2722 12131 2783 sw
tri 12424 2722 12485 2783 se
rect 12485 2722 12670 2959
tri 12670 2903 12726 2959 nw
tri 13029 2903 13085 2959 ne
tri 12670 2722 12731 2783 sw
tri 13024 2722 13085 2783 se
rect 13085 2722 13270 2959
tri 13270 2903 13326 2959 nw
tri 13629 2903 13685 2959 ne
tri 13270 2722 13331 2783 sw
tri 13624 2722 13685 2783 se
rect 13685 2722 13870 2959
tri 13870 2903 13926 2959 nw
tri 14229 2903 14285 2959 ne
tri 13870 2722 13931 2783 sw
tri 14224 2722 14285 2783 se
rect 14285 2722 14470 2959
tri 14470 2903 14526 2959 nw
tri 14829 2903 14885 2959 ne
tri 14470 2722 14531 2783 sw
tri 14824 2722 14885 2783 se
rect 14885 2722 15070 2959
tri 15070 2903 15126 2959 nw
tri 15429 2903 15485 2959 ne
tri 15070 2722 15131 2783 sw
tri 15424 2722 15485 2783 se
rect 15485 2722 15670 2959
tri 15670 2903 15726 2959 nw
tri 16029 2903 16085 2959 ne
tri 15670 2722 15731 2783 sw
tri 16024 2722 16085 2783 se
rect 16085 2722 16270 2959
tri 16270 2903 16326 2959 nw
tri 16270 2722 16331 2783 sw
rect 4722 2715 16940 2722
rect 4722 2681 4734 2715
rect 4768 2681 4807 2715
rect 4841 2681 4880 2715
rect 4914 2681 4953 2715
rect 4987 2681 5026 2715
rect 5060 2681 5099 2715
rect 5133 2681 5172 2715
rect 5206 2681 5245 2715
rect 5279 2681 5318 2715
rect 5352 2681 5391 2715
rect 5425 2681 5464 2715
rect 5498 2681 5537 2715
rect 5571 2681 5610 2715
rect 5644 2681 5683 2715
rect 5717 2681 5756 2715
rect 5790 2681 5829 2715
rect 5863 2681 5902 2715
rect 5936 2681 5975 2715
rect 6009 2681 6048 2715
rect 6082 2681 6121 2715
rect 6155 2681 6194 2715
rect 6228 2681 6267 2715
rect 6301 2681 6340 2715
rect 6374 2681 6413 2715
rect 6447 2681 6486 2715
rect 6520 2681 6559 2715
rect 6593 2681 6632 2715
rect 6666 2681 6705 2715
rect 6739 2681 6778 2715
rect 6812 2681 6851 2715
rect 6885 2681 6924 2715
rect 6958 2681 6997 2715
rect 7031 2681 7070 2715
rect 7104 2681 7143 2715
rect 7177 2681 7216 2715
rect 7250 2681 7289 2715
rect 7323 2681 7362 2715
rect 7396 2681 7435 2715
rect 7469 2681 7508 2715
rect 7542 2681 7581 2715
rect 7615 2681 7654 2715
rect 7688 2681 7727 2715
rect 7761 2681 7800 2715
rect 7834 2681 7873 2715
rect 7907 2681 7946 2715
rect 7980 2681 8019 2715
rect 8053 2681 8092 2715
rect 8126 2681 8165 2715
rect 8199 2681 8238 2715
rect 8272 2681 8311 2715
rect 8345 2681 8384 2715
rect 8418 2681 8457 2715
rect 8491 2681 8530 2715
rect 8564 2681 8603 2715
rect 8637 2681 8676 2715
rect 8710 2681 8749 2715
rect 8783 2681 8822 2715
rect 8856 2681 8895 2715
rect 8929 2681 8968 2715
rect 9002 2681 9041 2715
rect 9075 2681 9114 2715
rect 9148 2681 9187 2715
rect 9221 2681 9260 2715
rect 9294 2681 9333 2715
rect 9367 2681 9406 2715
rect 9440 2681 9479 2715
rect 9513 2681 9552 2715
rect 9586 2681 9625 2715
rect 9659 2681 9698 2715
rect 9732 2681 9771 2715
rect 9805 2681 9844 2715
rect 9878 2681 9917 2715
rect 9951 2681 9989 2715
rect 10023 2681 10061 2715
rect 10095 2681 10133 2715
rect 10167 2681 10205 2715
rect 10239 2681 10277 2715
rect 10311 2681 10349 2715
rect 10383 2681 10421 2715
rect 10455 2681 10493 2715
rect 10527 2681 10565 2715
rect 10599 2681 10637 2715
rect 10671 2681 10709 2715
rect 10743 2681 10781 2715
rect 10815 2681 10853 2715
rect 10887 2681 10925 2715
rect 10959 2697 16940 2715
rect 10959 2681 11967 2697
rect 4722 2663 11967 2681
rect 12001 2663 12040 2697
rect 12074 2663 12113 2697
rect 12147 2663 12186 2697
rect 12220 2663 12259 2697
rect 12293 2663 12332 2697
rect 12366 2663 12405 2697
rect 12439 2663 12478 2697
rect 12512 2663 12551 2697
rect 12585 2663 12624 2697
rect 12658 2663 12697 2697
rect 12731 2663 12770 2697
rect 12804 2663 12843 2697
rect 12877 2663 12916 2697
rect 12950 2663 12989 2697
rect 13023 2663 13062 2697
rect 13096 2663 13135 2697
rect 13169 2663 13208 2697
rect 13242 2663 13281 2697
rect 13315 2663 13354 2697
rect 13388 2663 13427 2697
rect 13461 2663 13500 2697
rect 13534 2663 13573 2697
rect 13607 2663 13646 2697
rect 13680 2663 13719 2697
rect 13753 2663 13792 2697
rect 13826 2663 13865 2697
rect 13899 2663 13938 2697
rect 13972 2663 14011 2697
rect 14045 2663 14084 2697
rect 14118 2663 14157 2697
rect 4722 2639 14157 2663
rect 4722 2605 4734 2639
rect 4768 2605 4807 2639
rect 4841 2605 4880 2639
rect 4914 2605 4953 2639
rect 4987 2605 5026 2639
rect 5060 2605 5099 2639
rect 5133 2605 5172 2639
rect 5206 2605 5245 2639
rect 5279 2605 5318 2639
rect 5352 2605 5391 2639
rect 5425 2605 5464 2639
rect 5498 2605 5537 2639
rect 5571 2605 5610 2639
rect 5644 2605 5683 2639
rect 5717 2605 5756 2639
rect 5790 2605 5829 2639
rect 5863 2605 5902 2639
rect 5936 2605 5975 2639
rect 6009 2605 6048 2639
rect 6082 2605 6121 2639
rect 6155 2605 6194 2639
rect 6228 2605 6267 2639
rect 6301 2605 6340 2639
rect 6374 2605 6413 2639
rect 6447 2605 6486 2639
rect 6520 2605 6559 2639
rect 6593 2605 6632 2639
rect 6666 2605 6705 2639
rect 6739 2605 6778 2639
rect 6812 2605 6851 2639
rect 6885 2605 6924 2639
rect 6958 2605 6997 2639
rect 7031 2605 7070 2639
rect 7104 2605 7143 2639
rect 7177 2605 7216 2639
rect 7250 2605 7289 2639
rect 7323 2605 7362 2639
rect 7396 2605 7435 2639
rect 7469 2605 7508 2639
rect 7542 2605 7581 2639
rect 7615 2605 7654 2639
rect 7688 2605 7727 2639
rect 7761 2605 7800 2639
rect 7834 2605 7873 2639
rect 7907 2605 7946 2639
rect 7980 2605 8019 2639
rect 8053 2605 8092 2639
rect 8126 2605 8165 2639
rect 8199 2605 8238 2639
rect 8272 2605 8311 2639
rect 8345 2605 8384 2639
rect 8418 2605 8457 2639
rect 8491 2605 8530 2639
rect 8564 2605 8603 2639
rect 8637 2605 8676 2639
rect 8710 2605 8749 2639
rect 8783 2605 8822 2639
rect 8856 2605 8895 2639
rect 8929 2605 8968 2639
rect 9002 2605 9041 2639
rect 9075 2605 9114 2639
rect 9148 2605 9187 2639
rect 9221 2605 9260 2639
rect 9294 2605 9333 2639
rect 9367 2605 9406 2639
rect 9440 2605 9479 2639
rect 9513 2605 9552 2639
rect 9586 2605 9625 2639
rect 9659 2605 9698 2639
rect 9732 2605 9771 2639
rect 9805 2605 9844 2639
rect 9878 2605 9917 2639
rect 9951 2605 9989 2639
rect 10023 2605 10061 2639
rect 10095 2605 10133 2639
rect 10167 2605 10205 2639
rect 10239 2605 10277 2639
rect 10311 2605 10349 2639
rect 10383 2605 10421 2639
rect 10455 2605 10493 2639
rect 10527 2605 10565 2639
rect 10599 2605 10637 2639
rect 10671 2605 10709 2639
rect 10743 2605 10781 2639
rect 10815 2605 10853 2639
rect 10887 2605 10925 2639
rect 10959 2625 14157 2639
rect 10959 2605 11967 2625
rect 4722 2591 11967 2605
rect 12001 2591 12040 2625
rect 12074 2591 12113 2625
rect 12147 2591 12186 2625
rect 12220 2591 12259 2625
rect 12293 2591 12332 2625
rect 12366 2591 12405 2625
rect 12439 2591 12478 2625
rect 12512 2591 12551 2625
rect 12585 2591 12624 2625
rect 12658 2591 12697 2625
rect 12731 2591 12770 2625
rect 12804 2591 12843 2625
rect 12877 2591 12916 2625
rect 12950 2591 12989 2625
rect 13023 2591 13062 2625
rect 13096 2591 13135 2625
rect 13169 2591 13208 2625
rect 13242 2591 13281 2625
rect 13315 2591 13354 2625
rect 13388 2591 13427 2625
rect 13461 2591 13500 2625
rect 13534 2591 13573 2625
rect 13607 2591 13646 2625
rect 13680 2591 13719 2625
rect 13753 2591 13792 2625
rect 13826 2591 13865 2625
rect 13899 2591 13938 2625
rect 13972 2591 14011 2625
rect 14045 2591 14084 2625
rect 14118 2591 14157 2625
rect 4722 2563 14157 2591
rect 4722 2529 4734 2563
rect 4768 2529 4807 2563
rect 4841 2529 4880 2563
rect 4914 2529 4953 2563
rect 4987 2529 5026 2563
rect 5060 2529 5099 2563
rect 5133 2529 5172 2563
rect 5206 2529 5245 2563
rect 5279 2529 5318 2563
rect 5352 2529 5391 2563
rect 5425 2529 5464 2563
rect 5498 2529 5537 2563
rect 5571 2529 5610 2563
rect 5644 2529 5683 2563
rect 5717 2529 5756 2563
rect 5790 2529 5829 2563
rect 5863 2529 5902 2563
rect 5936 2529 5975 2563
rect 6009 2529 6048 2563
rect 6082 2529 6121 2563
rect 6155 2529 6194 2563
rect 6228 2529 6267 2563
rect 6301 2529 6340 2563
rect 6374 2529 6413 2563
rect 6447 2529 6486 2563
rect 6520 2529 6559 2563
rect 6593 2529 6632 2563
rect 6666 2529 6705 2563
rect 6739 2529 6778 2563
rect 6812 2529 6851 2563
rect 6885 2529 6924 2563
rect 6958 2529 6997 2563
rect 7031 2529 7070 2563
rect 7104 2529 7143 2563
rect 7177 2529 7216 2563
rect 7250 2529 7289 2563
rect 7323 2529 7362 2563
rect 7396 2529 7435 2563
rect 7469 2529 7508 2563
rect 7542 2529 7581 2563
rect 7615 2529 7654 2563
rect 7688 2529 7727 2563
rect 7761 2529 7800 2563
rect 7834 2529 7873 2563
rect 7907 2529 7946 2563
rect 7980 2529 8019 2563
rect 8053 2529 8092 2563
rect 8126 2529 8165 2563
rect 8199 2529 8238 2563
rect 8272 2529 8311 2563
rect 8345 2529 8384 2563
rect 8418 2529 8457 2563
rect 8491 2529 8530 2563
rect 8564 2529 8603 2563
rect 8637 2529 8676 2563
rect 8710 2529 8749 2563
rect 8783 2529 8822 2563
rect 8856 2529 8895 2563
rect 8929 2529 8968 2563
rect 9002 2529 9041 2563
rect 9075 2529 9114 2563
rect 9148 2529 9187 2563
rect 9221 2529 9260 2563
rect 9294 2529 9333 2563
rect 9367 2529 9406 2563
rect 9440 2529 9479 2563
rect 9513 2529 9552 2563
rect 9586 2529 9625 2563
rect 9659 2529 9698 2563
rect 9732 2529 9771 2563
rect 9805 2529 9844 2563
rect 9878 2529 9917 2563
rect 9951 2529 9989 2563
rect 10023 2529 10061 2563
rect 10095 2529 10133 2563
rect 10167 2529 10205 2563
rect 10239 2529 10277 2563
rect 10311 2529 10349 2563
rect 10383 2529 10421 2563
rect 10455 2529 10493 2563
rect 10527 2529 10565 2563
rect 10599 2529 10637 2563
rect 10671 2529 10709 2563
rect 10743 2529 10781 2563
rect 10815 2529 10853 2563
rect 10887 2529 10925 2563
rect 10959 2553 14157 2563
rect 10959 2529 11967 2553
rect 4722 2519 11967 2529
rect 12001 2519 12040 2553
rect 12074 2519 12113 2553
rect 12147 2519 12186 2553
rect 12220 2519 12259 2553
rect 12293 2519 12332 2553
rect 12366 2519 12405 2553
rect 12439 2519 12478 2553
rect 12512 2519 12551 2553
rect 12585 2519 12624 2553
rect 12658 2519 12697 2553
rect 12731 2519 12770 2553
rect 12804 2519 12843 2553
rect 12877 2519 12916 2553
rect 12950 2519 12989 2553
rect 13023 2519 13062 2553
rect 13096 2519 13135 2553
rect 13169 2519 13208 2553
rect 13242 2519 13281 2553
rect 13315 2519 13354 2553
rect 13388 2519 13427 2553
rect 13461 2519 13500 2553
rect 13534 2519 13573 2553
rect 13607 2519 13646 2553
rect 13680 2519 13719 2553
rect 13753 2519 13792 2553
rect 13826 2519 13865 2553
rect 13899 2519 13938 2553
rect 13972 2519 14011 2553
rect 14045 2519 14084 2553
rect 14118 2519 14157 2553
rect 4722 2487 14157 2519
rect 4722 2453 4734 2487
rect 4768 2453 4807 2487
rect 4841 2453 4880 2487
rect 4914 2453 4953 2487
rect 4987 2453 5026 2487
rect 5060 2453 5099 2487
rect 5133 2453 5172 2487
rect 5206 2453 5245 2487
rect 5279 2453 5318 2487
rect 5352 2453 5391 2487
rect 5425 2453 5464 2487
rect 5498 2453 5537 2487
rect 5571 2453 5610 2487
rect 5644 2453 5683 2487
rect 5717 2453 5756 2487
rect 5790 2453 5829 2487
rect 5863 2453 5902 2487
rect 5936 2453 5975 2487
rect 6009 2453 6048 2487
rect 6082 2453 6121 2487
rect 6155 2453 6194 2487
rect 6228 2453 6267 2487
rect 6301 2453 6340 2487
rect 6374 2453 6413 2487
rect 6447 2453 6486 2487
rect 6520 2453 6559 2487
rect 6593 2453 6632 2487
rect 6666 2453 6705 2487
rect 6739 2453 6778 2487
rect 6812 2453 6851 2487
rect 6885 2453 6924 2487
rect 6958 2453 6997 2487
rect 7031 2453 7070 2487
rect 7104 2453 7143 2487
rect 7177 2453 7216 2487
rect 7250 2453 7289 2487
rect 7323 2453 7362 2487
rect 7396 2453 7435 2487
rect 7469 2453 7508 2487
rect 7542 2453 7581 2487
rect 7615 2453 7654 2487
rect 7688 2453 7727 2487
rect 7761 2453 7800 2487
rect 7834 2453 7873 2487
rect 7907 2453 7946 2487
rect 7980 2453 8019 2487
rect 8053 2453 8092 2487
rect 8126 2453 8165 2487
rect 8199 2453 8238 2487
rect 8272 2453 8311 2487
rect 8345 2453 8384 2487
rect 8418 2453 8457 2487
rect 8491 2453 8530 2487
rect 8564 2453 8603 2487
rect 8637 2453 8676 2487
rect 8710 2453 8749 2487
rect 8783 2453 8822 2487
rect 8856 2453 8895 2487
rect 8929 2453 8968 2487
rect 9002 2453 9041 2487
rect 9075 2453 9114 2487
rect 9148 2453 9187 2487
rect 9221 2453 9260 2487
rect 9294 2453 9333 2487
rect 9367 2453 9406 2487
rect 9440 2453 9479 2487
rect 9513 2453 9552 2487
rect 9586 2453 9625 2487
rect 9659 2453 9698 2487
rect 9732 2453 9771 2487
rect 9805 2453 9844 2487
rect 9878 2453 9917 2487
rect 9951 2453 9989 2487
rect 10023 2453 10061 2487
rect 10095 2453 10133 2487
rect 10167 2453 10205 2487
rect 10239 2453 10277 2487
rect 10311 2453 10349 2487
rect 10383 2453 10421 2487
rect 10455 2453 10493 2487
rect 10527 2453 10565 2487
rect 10599 2453 10637 2487
rect 10671 2453 10709 2487
rect 10743 2453 10781 2487
rect 10815 2453 10853 2487
rect 10887 2453 10925 2487
rect 10959 2481 14157 2487
rect 10959 2453 11967 2481
rect 4722 2447 11967 2453
rect 12001 2447 12040 2481
rect 12074 2447 12113 2481
rect 12147 2447 12186 2481
rect 12220 2447 12259 2481
rect 12293 2447 12332 2481
rect 12366 2447 12405 2481
rect 12439 2447 12478 2481
rect 12512 2447 12551 2481
rect 12585 2447 12624 2481
rect 12658 2447 12697 2481
rect 12731 2447 12770 2481
rect 12804 2447 12843 2481
rect 12877 2447 12916 2481
rect 12950 2447 12989 2481
rect 13023 2447 13062 2481
rect 13096 2447 13135 2481
rect 13169 2447 13208 2481
rect 13242 2447 13281 2481
rect 13315 2447 13354 2481
rect 13388 2447 13427 2481
rect 13461 2447 13500 2481
rect 13534 2447 13573 2481
rect 13607 2447 13646 2481
rect 13680 2447 13719 2481
rect 13753 2447 13792 2481
rect 13826 2447 13865 2481
rect 13899 2447 13938 2481
rect 13972 2447 14011 2481
rect 14045 2447 14084 2481
rect 14118 2447 14157 2481
rect 4722 2411 14157 2447
rect 4722 2377 4734 2411
rect 4768 2377 4807 2411
rect 4841 2377 4880 2411
rect 4914 2377 4953 2411
rect 4987 2377 5026 2411
rect 5060 2377 5099 2411
rect 5133 2377 5172 2411
rect 5206 2377 5245 2411
rect 5279 2377 5318 2411
rect 5352 2377 5391 2411
rect 5425 2377 5464 2411
rect 5498 2377 5537 2411
rect 5571 2377 5610 2411
rect 5644 2377 5683 2411
rect 5717 2377 5756 2411
rect 5790 2377 5829 2411
rect 5863 2377 5902 2411
rect 5936 2377 5975 2411
rect 6009 2377 6048 2411
rect 6082 2377 6121 2411
rect 6155 2377 6194 2411
rect 6228 2377 6267 2411
rect 6301 2377 6340 2411
rect 6374 2377 6413 2411
rect 6447 2377 6486 2411
rect 6520 2377 6559 2411
rect 6593 2377 6632 2411
rect 6666 2377 6705 2411
rect 6739 2377 6778 2411
rect 6812 2377 6851 2411
rect 6885 2377 6924 2411
rect 6958 2377 6997 2411
rect 7031 2377 7070 2411
rect 7104 2377 7143 2411
rect 7177 2377 7216 2411
rect 7250 2377 7289 2411
rect 7323 2377 7362 2411
rect 7396 2377 7435 2411
rect 7469 2377 7508 2411
rect 7542 2377 7581 2411
rect 7615 2377 7654 2411
rect 7688 2377 7727 2411
rect 7761 2377 7800 2411
rect 7834 2377 7873 2411
rect 7907 2377 7946 2411
rect 7980 2377 8019 2411
rect 8053 2377 8092 2411
rect 8126 2377 8165 2411
rect 8199 2377 8238 2411
rect 8272 2377 8311 2411
rect 8345 2377 8384 2411
rect 8418 2377 8457 2411
rect 8491 2377 8530 2411
rect 8564 2377 8603 2411
rect 8637 2377 8676 2411
rect 8710 2377 8749 2411
rect 8783 2377 8822 2411
rect 8856 2377 8895 2411
rect 8929 2377 8968 2411
rect 9002 2377 9041 2411
rect 9075 2377 9114 2411
rect 9148 2377 9187 2411
rect 9221 2377 9260 2411
rect 9294 2377 9333 2411
rect 9367 2377 9406 2411
rect 9440 2377 9479 2411
rect 9513 2377 9552 2411
rect 9586 2377 9625 2411
rect 9659 2377 9698 2411
rect 9732 2377 9771 2411
rect 9805 2377 9844 2411
rect 9878 2377 9917 2411
rect 9951 2377 9989 2411
rect 10023 2377 10061 2411
rect 10095 2377 10133 2411
rect 10167 2377 10205 2411
rect 10239 2377 10277 2411
rect 10311 2377 10349 2411
rect 10383 2377 10421 2411
rect 10455 2377 10493 2411
rect 10527 2377 10565 2411
rect 10599 2377 10637 2411
rect 10671 2377 10709 2411
rect 10743 2377 10781 2411
rect 10815 2377 10853 2411
rect 10887 2377 10925 2411
rect 10959 2409 14157 2411
rect 10959 2377 11967 2409
rect 4722 2375 11967 2377
rect 12001 2375 12040 2409
rect 12074 2375 12113 2409
rect 12147 2375 12186 2409
rect 12220 2375 12259 2409
rect 12293 2375 12332 2409
rect 12366 2375 12405 2409
rect 12439 2375 12478 2409
rect 12512 2375 12551 2409
rect 12585 2375 12624 2409
rect 12658 2375 12697 2409
rect 12731 2375 12770 2409
rect 12804 2375 12843 2409
rect 12877 2375 12916 2409
rect 12950 2375 12989 2409
rect 13023 2375 13062 2409
rect 13096 2375 13135 2409
rect 13169 2375 13208 2409
rect 13242 2375 13281 2409
rect 13315 2375 13354 2409
rect 13388 2375 13427 2409
rect 13461 2375 13500 2409
rect 13534 2375 13573 2409
rect 13607 2375 13646 2409
rect 13680 2375 13719 2409
rect 13753 2375 13792 2409
rect 13826 2375 13865 2409
rect 13899 2375 13938 2409
rect 13972 2375 14011 2409
rect 14045 2375 14084 2409
rect 14118 2375 14157 2409
rect 4722 2337 14157 2375
rect 4722 2335 11967 2337
rect 4722 2301 4734 2335
rect 4768 2301 4807 2335
rect 4841 2301 4880 2335
rect 4914 2301 4953 2335
rect 4987 2301 5026 2335
rect 5060 2301 5099 2335
rect 5133 2301 5172 2335
rect 5206 2301 5245 2335
rect 5279 2301 5318 2335
rect 5352 2301 5391 2335
rect 5425 2301 5464 2335
rect 5498 2301 5537 2335
rect 5571 2301 5610 2335
rect 5644 2301 5683 2335
rect 5717 2301 5756 2335
rect 5790 2301 5829 2335
rect 5863 2301 5902 2335
rect 5936 2301 5975 2335
rect 6009 2301 6048 2335
rect 6082 2301 6121 2335
rect 6155 2301 6194 2335
rect 6228 2301 6267 2335
rect 6301 2301 6340 2335
rect 6374 2301 6413 2335
rect 6447 2301 6486 2335
rect 6520 2301 6559 2335
rect 6593 2301 6632 2335
rect 6666 2301 6705 2335
rect 6739 2301 6778 2335
rect 6812 2301 6851 2335
rect 6885 2301 6924 2335
rect 6958 2301 6997 2335
rect 7031 2301 7070 2335
rect 7104 2301 7143 2335
rect 7177 2301 7216 2335
rect 7250 2301 7289 2335
rect 7323 2301 7362 2335
rect 7396 2301 7435 2335
rect 7469 2301 7508 2335
rect 7542 2301 7581 2335
rect 7615 2301 7654 2335
rect 7688 2301 7727 2335
rect 7761 2301 7800 2335
rect 7834 2301 7873 2335
rect 7907 2301 7946 2335
rect 7980 2301 8019 2335
rect 8053 2301 8092 2335
rect 8126 2301 8165 2335
rect 8199 2301 8238 2335
rect 8272 2301 8311 2335
rect 8345 2301 8384 2335
rect 8418 2301 8457 2335
rect 8491 2301 8530 2335
rect 8564 2301 8603 2335
rect 8637 2301 8676 2335
rect 8710 2301 8749 2335
rect 8783 2301 8822 2335
rect 8856 2301 8895 2335
rect 8929 2301 8968 2335
rect 9002 2301 9041 2335
rect 9075 2301 9114 2335
rect 9148 2301 9187 2335
rect 9221 2301 9260 2335
rect 9294 2301 9333 2335
rect 9367 2301 9406 2335
rect 9440 2301 9479 2335
rect 9513 2301 9552 2335
rect 9586 2301 9625 2335
rect 9659 2301 9698 2335
rect 9732 2301 9771 2335
rect 9805 2301 9844 2335
rect 9878 2301 9917 2335
rect 9951 2301 9989 2335
rect 10023 2301 10061 2335
rect 10095 2301 10133 2335
rect 10167 2301 10205 2335
rect 10239 2301 10277 2335
rect 10311 2301 10349 2335
rect 10383 2301 10421 2335
rect 10455 2301 10493 2335
rect 10527 2301 10565 2335
rect 10599 2301 10637 2335
rect 10671 2301 10709 2335
rect 10743 2301 10781 2335
rect 10815 2301 10853 2335
rect 10887 2301 10925 2335
rect 10959 2303 11967 2335
rect 12001 2303 12040 2337
rect 12074 2303 12113 2337
rect 12147 2303 12186 2337
rect 12220 2303 12259 2337
rect 12293 2303 12332 2337
rect 12366 2303 12405 2337
rect 12439 2303 12478 2337
rect 12512 2303 12551 2337
rect 12585 2303 12624 2337
rect 12658 2303 12697 2337
rect 12731 2303 12770 2337
rect 12804 2303 12843 2337
rect 12877 2303 12916 2337
rect 12950 2303 12989 2337
rect 13023 2303 13062 2337
rect 13096 2303 13135 2337
rect 13169 2303 13208 2337
rect 13242 2303 13281 2337
rect 13315 2303 13354 2337
rect 13388 2303 13427 2337
rect 13461 2303 13500 2337
rect 13534 2303 13573 2337
rect 13607 2303 13646 2337
rect 13680 2303 13719 2337
rect 13753 2303 13792 2337
rect 13826 2303 13865 2337
rect 13899 2303 13938 2337
rect 13972 2303 14011 2337
rect 14045 2303 14084 2337
rect 14118 2303 14157 2337
rect 10959 2301 14157 2303
rect 4722 2265 14157 2301
rect 4722 2259 11967 2265
rect 4722 2225 4734 2259
rect 4768 2225 4807 2259
rect 4841 2225 4880 2259
rect 4914 2225 4953 2259
rect 4987 2225 5026 2259
rect 5060 2225 5099 2259
rect 5133 2225 5172 2259
rect 5206 2225 5245 2259
rect 5279 2225 5318 2259
rect 5352 2225 5391 2259
rect 5425 2225 5464 2259
rect 5498 2225 5537 2259
rect 5571 2225 5610 2259
rect 5644 2225 5683 2259
rect 5717 2225 5756 2259
rect 5790 2225 5829 2259
rect 5863 2225 5902 2259
rect 5936 2225 5975 2259
rect 6009 2225 6048 2259
rect 6082 2225 6121 2259
rect 6155 2225 6194 2259
rect 6228 2225 6267 2259
rect 6301 2225 6340 2259
rect 6374 2225 6413 2259
rect 6447 2225 6486 2259
rect 6520 2225 6559 2259
rect 6593 2225 6632 2259
rect 6666 2225 6705 2259
rect 6739 2225 6778 2259
rect 6812 2225 6851 2259
rect 6885 2225 6924 2259
rect 6958 2225 6997 2259
rect 7031 2225 7070 2259
rect 7104 2225 7143 2259
rect 7177 2225 7216 2259
rect 7250 2225 7289 2259
rect 7323 2225 7362 2259
rect 7396 2225 7435 2259
rect 7469 2225 7508 2259
rect 7542 2225 7581 2259
rect 7615 2225 7654 2259
rect 7688 2225 7727 2259
rect 7761 2225 7800 2259
rect 7834 2225 7873 2259
rect 7907 2225 7946 2259
rect 7980 2225 8019 2259
rect 8053 2225 8092 2259
rect 8126 2225 8165 2259
rect 8199 2225 8238 2259
rect 8272 2225 8311 2259
rect 8345 2225 8384 2259
rect 8418 2225 8457 2259
rect 8491 2225 8530 2259
rect 8564 2225 8603 2259
rect 8637 2225 8676 2259
rect 8710 2225 8749 2259
rect 8783 2225 8822 2259
rect 8856 2225 8895 2259
rect 8929 2225 8968 2259
rect 9002 2225 9041 2259
rect 9075 2225 9114 2259
rect 9148 2225 9187 2259
rect 9221 2225 9260 2259
rect 9294 2225 9333 2259
rect 9367 2225 9406 2259
rect 9440 2225 9479 2259
rect 9513 2225 9552 2259
rect 9586 2225 9625 2259
rect 9659 2225 9698 2259
rect 9732 2225 9771 2259
rect 9805 2225 9844 2259
rect 9878 2225 9917 2259
rect 9951 2225 9989 2259
rect 10023 2225 10061 2259
rect 10095 2225 10133 2259
rect 10167 2225 10205 2259
rect 10239 2225 10277 2259
rect 10311 2225 10349 2259
rect 10383 2225 10421 2259
rect 10455 2225 10493 2259
rect 10527 2225 10565 2259
rect 10599 2225 10637 2259
rect 10671 2225 10709 2259
rect 10743 2225 10781 2259
rect 10815 2225 10853 2259
rect 10887 2225 10925 2259
rect 10959 2231 11967 2259
rect 12001 2231 12040 2265
rect 12074 2231 12113 2265
rect 12147 2231 12186 2265
rect 12220 2231 12259 2265
rect 12293 2231 12332 2265
rect 12366 2231 12405 2265
rect 12439 2231 12478 2265
rect 12512 2231 12551 2265
rect 12585 2231 12624 2265
rect 12658 2231 12697 2265
rect 12731 2231 12770 2265
rect 12804 2231 12843 2265
rect 12877 2231 12916 2265
rect 12950 2231 12989 2265
rect 13023 2231 13062 2265
rect 13096 2231 13135 2265
rect 13169 2231 13208 2265
rect 13242 2231 13281 2265
rect 13315 2231 13354 2265
rect 13388 2231 13427 2265
rect 13461 2231 13500 2265
rect 13534 2231 13573 2265
rect 13607 2231 13646 2265
rect 13680 2231 13719 2265
rect 13753 2231 13792 2265
rect 13826 2231 13865 2265
rect 13899 2231 13938 2265
rect 13972 2231 14011 2265
rect 14045 2231 14084 2265
rect 14118 2231 14157 2265
rect 10959 2225 14157 2231
rect 4722 2193 14157 2225
rect 4722 2183 11967 2193
rect 4722 2149 4734 2183
rect 4768 2149 4807 2183
rect 4841 2149 4880 2183
rect 4914 2149 4953 2183
rect 4987 2149 5026 2183
rect 5060 2149 5099 2183
rect 5133 2149 5172 2183
rect 5206 2149 5245 2183
rect 5279 2149 5318 2183
rect 5352 2149 5391 2183
rect 5425 2149 5464 2183
rect 5498 2149 5537 2183
rect 5571 2149 5610 2183
rect 5644 2149 5683 2183
rect 5717 2149 5756 2183
rect 5790 2149 5829 2183
rect 5863 2149 5902 2183
rect 5936 2149 5975 2183
rect 6009 2149 6048 2183
rect 6082 2149 6121 2183
rect 6155 2149 6194 2183
rect 6228 2149 6267 2183
rect 6301 2149 6340 2183
rect 6374 2149 6413 2183
rect 6447 2149 6486 2183
rect 6520 2149 6559 2183
rect 6593 2149 6632 2183
rect 6666 2149 6705 2183
rect 6739 2149 6778 2183
rect 6812 2149 6851 2183
rect 6885 2149 6924 2183
rect 6958 2149 6997 2183
rect 7031 2149 7070 2183
rect 7104 2149 7143 2183
rect 7177 2149 7216 2183
rect 7250 2149 7289 2183
rect 7323 2149 7362 2183
rect 7396 2149 7435 2183
rect 7469 2149 7508 2183
rect 7542 2149 7581 2183
rect 7615 2149 7654 2183
rect 7688 2149 7727 2183
rect 7761 2149 7800 2183
rect 7834 2149 7873 2183
rect 7907 2149 7946 2183
rect 7980 2149 8019 2183
rect 8053 2149 8092 2183
rect 8126 2149 8165 2183
rect 8199 2149 8238 2183
rect 8272 2149 8311 2183
rect 8345 2149 8384 2183
rect 8418 2149 8457 2183
rect 8491 2149 8530 2183
rect 8564 2149 8603 2183
rect 8637 2149 8676 2183
rect 8710 2149 8749 2183
rect 8783 2149 8822 2183
rect 8856 2149 8895 2183
rect 8929 2149 8968 2183
rect 9002 2149 9041 2183
rect 9075 2149 9114 2183
rect 9148 2149 9187 2183
rect 9221 2149 9260 2183
rect 9294 2149 9333 2183
rect 9367 2149 9406 2183
rect 9440 2149 9479 2183
rect 9513 2149 9552 2183
rect 9586 2149 9625 2183
rect 9659 2149 9698 2183
rect 9732 2149 9771 2183
rect 9805 2149 9844 2183
rect 9878 2149 9917 2183
rect 9951 2149 9989 2183
rect 10023 2149 10061 2183
rect 10095 2149 10133 2183
rect 10167 2149 10205 2183
rect 10239 2149 10277 2183
rect 10311 2149 10349 2183
rect 10383 2149 10421 2183
rect 10455 2149 10493 2183
rect 10527 2149 10565 2183
rect 10599 2149 10637 2183
rect 10671 2149 10709 2183
rect 10743 2149 10781 2183
rect 10815 2149 10853 2183
rect 10887 2149 10925 2183
rect 10959 2159 11967 2183
rect 12001 2159 12040 2193
rect 12074 2159 12113 2193
rect 12147 2159 12186 2193
rect 12220 2159 12259 2193
rect 12293 2159 12332 2193
rect 12366 2159 12405 2193
rect 12439 2159 12478 2193
rect 12512 2159 12551 2193
rect 12585 2159 12624 2193
rect 12658 2159 12697 2193
rect 12731 2159 12770 2193
rect 12804 2159 12843 2193
rect 12877 2159 12916 2193
rect 12950 2159 12989 2193
rect 13023 2159 13062 2193
rect 13096 2159 13135 2193
rect 13169 2159 13208 2193
rect 13242 2159 13281 2193
rect 13315 2159 13354 2193
rect 13388 2159 13427 2193
rect 13461 2159 13500 2193
rect 13534 2159 13573 2193
rect 13607 2159 13646 2193
rect 13680 2159 13719 2193
rect 13753 2159 13792 2193
rect 13826 2159 13865 2193
rect 13899 2159 13938 2193
rect 13972 2159 14011 2193
rect 14045 2159 14084 2193
rect 14118 2159 14157 2193
rect 16927 2159 16940 2697
rect 10959 2149 16940 2159
rect 4722 2142 16940 2149
tri 10970 2141 10971 2142 ne
rect 10971 2141 16940 2142
rect 1999 1921 17332 2086
tri 424 1865 450 1891 se
rect 450 1865 705 1891
tri 705 1865 731 1891 sw
tri 1024 1865 1050 1891 se
rect 1050 1865 1305 1891
tri 1305 1865 1331 1891 sw
tri 113 1864 114 1865 se
rect 114 1864 17064 1865
rect -2844 1858 17064 1864
rect -2844 1841 4616 1858
rect -2844 1807 -2832 1841
rect -2798 1807 -2759 1841
rect -2725 1807 -2686 1841
rect -2652 1807 -2613 1841
rect -2579 1807 -2540 1841
rect -2506 1807 -2467 1841
rect -2433 1807 -2394 1841
rect -2360 1807 -2321 1841
rect -2287 1807 -2248 1841
rect -2214 1807 -2175 1841
rect -2141 1807 -2102 1841
rect -2068 1807 -2029 1841
rect -1995 1807 -1956 1841
rect -1922 1807 -1883 1841
rect -1849 1807 -1810 1841
rect -1776 1807 -1737 1841
rect -2844 1769 -1737 1807
rect 4561 1824 4616 1841
rect 4650 1824 4688 1858
rect 4722 1824 4760 1858
rect 4794 1824 4832 1858
rect 4866 1824 4904 1858
rect 4938 1824 4976 1858
rect 5010 1824 5048 1858
rect 5082 1824 5120 1858
rect 5154 1824 5192 1858
rect 5226 1824 5264 1858
rect 5298 1824 5336 1858
rect 5370 1824 5408 1858
rect 5442 1824 5480 1858
rect 5514 1824 5552 1858
rect 5586 1824 5624 1858
rect 5658 1824 5696 1858
rect 5730 1824 5768 1858
rect 5802 1824 5840 1858
rect 5874 1824 5912 1858
rect 5946 1824 5984 1858
rect 6018 1824 6056 1858
rect 6090 1824 6128 1858
rect 6162 1824 6200 1858
rect 6234 1824 6272 1858
rect 6306 1824 6344 1858
rect 6378 1824 6416 1858
rect 6450 1824 6488 1858
rect 6522 1824 6560 1858
rect 6594 1824 6632 1858
rect 6666 1824 6704 1858
rect 6738 1824 6776 1858
rect 6810 1824 6848 1858
rect 6882 1824 6920 1858
rect 6954 1824 6992 1858
rect 7026 1824 7064 1858
rect 7098 1824 7136 1858
rect 7170 1824 7208 1858
rect 7242 1824 7280 1858
rect 7314 1824 7352 1858
rect 7386 1824 7424 1858
rect 7458 1824 7496 1858
rect 7530 1824 7568 1858
rect 7602 1824 7640 1858
rect 7674 1824 7712 1858
rect 7746 1824 7784 1858
rect 7818 1824 7856 1858
rect 7890 1824 7928 1858
rect 7962 1824 8000 1858
rect 8034 1824 8072 1858
rect 8106 1824 8144 1858
rect 8178 1824 8216 1858
rect 8250 1824 8288 1858
rect 8322 1824 8360 1858
rect 8394 1824 8432 1858
rect 8466 1824 8504 1858
rect 8538 1824 8576 1858
rect 8610 1824 8648 1858
rect 8682 1824 8720 1858
rect 8754 1824 8792 1858
rect 8826 1824 8864 1858
rect 8898 1824 8936 1858
rect 8970 1824 9008 1858
rect 9042 1824 9080 1858
rect 9114 1824 9152 1858
rect 9186 1824 9224 1858
rect 9258 1824 9296 1858
rect 9330 1824 9368 1858
rect 9402 1824 9440 1858
rect 9474 1824 9512 1858
rect 9546 1824 9584 1858
rect 9618 1824 9656 1858
rect 9690 1824 9728 1858
rect 9762 1824 9800 1858
rect 9834 1824 9872 1858
rect 9906 1824 9944 1858
rect 9978 1824 10016 1858
rect 10050 1824 10088 1858
rect 10122 1824 10160 1858
rect 10194 1824 10232 1858
rect 10266 1824 10304 1858
rect 10338 1824 10376 1858
rect 10410 1824 10448 1858
rect 10482 1824 10520 1858
rect 10554 1824 10592 1858
rect 10626 1824 10664 1858
rect 10698 1824 10736 1858
rect 10770 1824 10808 1858
rect 10842 1824 10880 1858
rect 10914 1824 10952 1858
rect 10986 1824 11024 1858
rect 11058 1824 11096 1858
rect 11130 1824 11168 1858
rect 11202 1824 11240 1858
rect 11274 1824 11312 1858
rect 11346 1824 11384 1858
rect 11418 1824 11456 1858
rect 11490 1824 11528 1858
rect 11562 1824 11600 1858
rect 11634 1824 11672 1858
rect 11706 1824 11744 1858
rect 11778 1824 11816 1858
rect 11850 1824 11888 1858
rect 11922 1824 11960 1858
rect 11994 1824 12032 1858
rect 12066 1824 12104 1858
rect 12138 1824 12176 1858
rect 12210 1824 12248 1858
rect 12282 1824 12320 1858
rect 12354 1824 12392 1858
rect 12426 1824 12464 1858
rect 12498 1824 12536 1858
rect 12570 1824 12608 1858
rect 12642 1824 12680 1858
rect 12714 1824 12752 1858
rect 12786 1824 12824 1858
rect 12858 1824 12896 1858
rect 12930 1824 12968 1858
rect 13002 1824 13040 1858
rect 13074 1824 13112 1858
rect 13146 1824 13184 1858
rect 13218 1824 13256 1858
rect 13290 1824 13328 1858
rect 13362 1824 13400 1858
rect 13434 1824 13472 1858
rect 13506 1824 13544 1858
rect 13578 1824 13616 1858
rect 13650 1824 13688 1858
rect 13722 1824 13760 1858
rect 13794 1824 13832 1858
rect 13866 1824 13904 1858
rect 13938 1824 13976 1858
rect 14010 1824 14048 1858
rect 14082 1824 14120 1858
rect 14154 1824 14192 1858
rect 14226 1824 14264 1858
rect 14298 1824 14336 1858
rect 14370 1824 14408 1858
rect 14442 1824 14480 1858
rect 14514 1824 14552 1858
rect 14586 1824 14624 1858
rect 14658 1824 14696 1858
rect 14730 1824 14768 1858
rect 14802 1824 14840 1858
rect 14874 1824 14912 1858
rect 14946 1824 14984 1858
rect 15018 1824 15056 1858
rect 15090 1824 15128 1858
rect 15162 1824 15200 1858
rect 15234 1824 15272 1858
rect 15306 1824 15344 1858
rect 15378 1824 15416 1858
rect 15450 1824 15488 1858
rect 15522 1824 15561 1858
rect 15595 1824 15634 1858
rect 15668 1824 15707 1858
rect 15741 1824 15780 1858
rect 15814 1824 15853 1858
rect 15887 1824 15926 1858
rect 15960 1824 15999 1858
rect 16033 1824 16072 1858
rect 16106 1824 16145 1858
rect 16179 1824 16218 1858
rect 16252 1824 16291 1858
rect 16325 1824 16364 1858
rect 16398 1824 16437 1858
rect 16471 1824 16510 1858
rect 16544 1824 16583 1858
rect 16617 1824 16656 1858
rect 16690 1824 17064 1858
rect 4561 1801 17064 1824
tri 17064 1801 17128 1865 sw
rect 4561 1780 17128 1801
rect -2844 1735 -2832 1769
rect -2798 1735 -2759 1769
rect -2725 1735 -2686 1769
rect -2652 1735 -2613 1769
rect -2579 1735 -2540 1769
rect -2506 1735 -2467 1769
rect -2433 1735 -2394 1769
rect -2360 1735 -2321 1769
rect -2287 1735 -2248 1769
rect -2214 1735 -2175 1769
rect -2141 1735 -2102 1769
rect -2068 1735 -2029 1769
rect -1995 1735 -1956 1769
rect -1922 1735 -1883 1769
rect -1849 1735 -1810 1769
rect -1776 1735 -1737 1769
rect -2844 1697 -1737 1735
rect 4561 1750 4616 1780
rect 4650 1750 4688 1780
rect 4722 1750 4760 1780
rect 4561 1698 4563 1750
rect 4615 1746 4616 1750
rect 4679 1746 4688 1750
rect 4743 1746 4760 1750
rect 4794 1746 4832 1780
rect 4866 1746 4904 1780
rect 4938 1746 4976 1780
rect 5010 1746 5048 1780
rect 5082 1746 5120 1780
rect 5154 1746 5192 1780
rect 5226 1746 5264 1780
rect 5298 1746 5336 1780
rect 5370 1746 5408 1780
rect 5442 1746 5480 1780
rect 5514 1746 5552 1780
rect 5586 1746 5624 1780
rect 5658 1746 5696 1780
rect 5730 1746 5768 1780
rect 5802 1746 5840 1780
rect 5874 1746 5912 1780
rect 5946 1746 5984 1780
rect 6018 1746 6056 1780
rect 6090 1746 6128 1780
rect 6162 1746 6200 1780
rect 6234 1746 6272 1780
rect 6306 1746 6344 1780
rect 6378 1746 6416 1780
rect 6450 1746 6488 1780
rect 6522 1746 6560 1780
rect 6594 1746 6632 1780
rect 6666 1746 6704 1780
rect 6738 1746 6776 1780
rect 6810 1746 6848 1780
rect 6882 1746 6920 1780
rect 6954 1746 6992 1780
rect 7026 1746 7064 1780
rect 7098 1746 7136 1780
rect 7170 1746 7208 1780
rect 7242 1746 7280 1780
rect 7314 1746 7352 1780
rect 7386 1746 7424 1780
rect 7458 1746 7496 1780
rect 7530 1746 7568 1780
rect 7602 1746 7640 1780
rect 7674 1746 7712 1780
rect 7746 1746 7784 1780
rect 7818 1746 7856 1780
rect 7890 1746 7928 1780
rect 7962 1746 8000 1780
rect 8034 1746 8072 1780
rect 8106 1746 8144 1780
rect 8178 1746 8216 1780
rect 8250 1746 8288 1780
rect 8322 1746 8360 1780
rect 8394 1746 8432 1780
rect 8466 1746 8504 1780
rect 8538 1746 8576 1780
rect 8610 1746 8648 1780
rect 8682 1746 8720 1780
rect 8754 1746 8792 1780
rect 8826 1746 8864 1780
rect 8898 1746 8936 1780
rect 8970 1746 9008 1780
rect 9042 1746 9080 1780
rect 9114 1746 9152 1780
rect 9186 1746 9224 1780
rect 9258 1746 9296 1780
rect 9330 1746 9368 1780
rect 9402 1746 9440 1780
rect 9474 1746 9512 1780
rect 9546 1746 9584 1780
rect 9618 1746 9656 1780
rect 9690 1746 9728 1780
rect 9762 1746 9800 1780
rect 9834 1746 9872 1780
rect 9906 1746 9944 1780
rect 9978 1746 10016 1780
rect 10050 1746 10088 1780
rect 10122 1746 10160 1780
rect 10194 1746 10232 1780
rect 10266 1746 10304 1780
rect 10338 1746 10376 1780
rect 10410 1746 10448 1780
rect 10482 1746 10520 1780
rect 10554 1746 10592 1780
rect 10626 1746 10664 1780
rect 10698 1746 10736 1780
rect 10770 1746 10808 1780
rect 10842 1746 10880 1780
rect 10914 1746 10952 1780
rect 10986 1746 11024 1780
rect 11058 1746 11096 1780
rect 11130 1746 11168 1780
rect 11202 1746 11240 1780
rect 11274 1746 11312 1780
rect 11346 1746 11384 1780
rect 11418 1746 11456 1780
rect 11490 1746 11528 1780
rect 11562 1746 11600 1780
rect 11634 1746 11672 1780
rect 11706 1746 11744 1780
rect 11778 1746 11816 1780
rect 11850 1746 11888 1780
rect 11922 1746 11960 1780
rect 11994 1746 12032 1780
rect 12066 1746 12104 1780
rect 12138 1746 12176 1780
rect 12210 1746 12248 1780
rect 12282 1746 12320 1780
rect 12354 1746 12392 1780
rect 12426 1746 12464 1780
rect 12498 1746 12536 1780
rect 12570 1746 12608 1780
rect 12642 1746 12680 1780
rect 12714 1746 12752 1780
rect 12786 1746 12824 1780
rect 12858 1746 12896 1780
rect 12930 1746 12968 1780
rect 13002 1746 13040 1780
rect 13074 1746 13112 1780
rect 13146 1746 13184 1780
rect 13218 1746 13256 1780
rect 13290 1746 13328 1780
rect 13362 1746 13400 1780
rect 13434 1746 13472 1780
rect 13506 1746 13544 1780
rect 13578 1746 13616 1780
rect 13650 1746 13688 1780
rect 13722 1746 13760 1780
rect 13794 1746 13832 1780
rect 13866 1746 13904 1780
rect 13938 1746 13976 1780
rect 14010 1746 14048 1780
rect 14082 1746 14120 1780
rect 14154 1746 14192 1780
rect 14226 1746 14264 1780
rect 14298 1746 14336 1780
rect 14370 1746 14408 1780
rect 14442 1746 14480 1780
rect 14514 1746 14552 1780
rect 14586 1746 14624 1780
rect 14658 1746 14696 1780
rect 14730 1746 14768 1780
rect 14802 1746 14840 1780
rect 14874 1746 14912 1780
rect 14946 1746 14984 1780
rect 15018 1746 15056 1780
rect 15090 1746 15128 1780
rect 15162 1746 15200 1780
rect 15234 1746 15272 1780
rect 15306 1746 15344 1780
rect 15378 1746 15416 1780
rect 15450 1746 15488 1780
rect 15522 1746 15561 1780
rect 15595 1746 15634 1780
rect 15668 1746 15707 1780
rect 15741 1746 15780 1780
rect 15814 1746 15853 1780
rect 15887 1746 15926 1780
rect 15960 1746 15999 1780
rect 16033 1746 16072 1780
rect 16106 1746 16145 1780
rect 16179 1746 16218 1780
rect 16252 1746 16291 1780
rect 16325 1746 16364 1780
rect 16398 1746 16437 1780
rect 16471 1746 16510 1780
rect 16544 1746 16583 1780
rect 16617 1746 16656 1780
rect 16690 1746 17128 1780
rect 4615 1702 4627 1746
rect 4679 1702 4691 1746
rect 4743 1702 17128 1746
rect 4615 1698 4616 1702
rect 4679 1698 4688 1702
rect 4743 1698 4760 1702
rect -2844 1663 -2832 1697
rect -2798 1663 -2759 1697
rect -2725 1663 -2686 1697
rect -2652 1663 -2613 1697
rect -2579 1663 -2540 1697
rect -2506 1663 -2467 1697
rect -2433 1663 -2394 1697
rect -2360 1663 -2321 1697
rect -2287 1663 -2248 1697
rect -2214 1663 -2175 1697
rect -2141 1663 -2102 1697
rect -2068 1663 -2029 1697
rect -1995 1663 -1956 1697
rect -1922 1663 -1883 1697
rect -1849 1663 -1810 1697
rect -1776 1663 -1737 1697
rect -2844 1625 -1737 1663
rect 4561 1682 4616 1698
rect 4650 1682 4688 1698
rect 4722 1682 4760 1698
rect 4561 1630 4563 1682
rect 4615 1668 4616 1682
rect 4679 1668 4688 1682
rect 4743 1668 4760 1682
rect 4794 1668 4832 1702
rect 4866 1668 4904 1702
rect 4938 1668 4976 1702
rect 5010 1668 5048 1702
rect 5082 1668 5120 1702
rect 5154 1668 5192 1702
rect 5226 1668 5264 1702
rect 5298 1668 5336 1702
rect 5370 1668 5408 1702
rect 5442 1668 5480 1702
rect 5514 1668 5552 1702
rect 5586 1668 5624 1702
rect 5658 1668 5696 1702
rect 5730 1668 5768 1702
rect 5802 1668 5840 1702
rect 5874 1668 5912 1702
rect 5946 1668 5984 1702
rect 6018 1668 6056 1702
rect 6090 1668 6128 1702
rect 6162 1668 6200 1702
rect 6234 1668 6272 1702
rect 6306 1668 6344 1702
rect 6378 1668 6416 1702
rect 6450 1668 6488 1702
rect 6522 1668 6560 1702
rect 6594 1668 6632 1702
rect 6666 1668 6704 1702
rect 6738 1668 6776 1702
rect 6810 1668 6848 1702
rect 6882 1668 6920 1702
rect 6954 1668 6992 1702
rect 7026 1668 7064 1702
rect 7098 1668 7136 1702
rect 7170 1668 7208 1702
rect 7242 1668 7280 1702
rect 7314 1668 7352 1702
rect 7386 1668 7424 1702
rect 7458 1668 7496 1702
rect 7530 1668 7568 1702
rect 7602 1668 7640 1702
rect 7674 1668 7712 1702
rect 7746 1668 7784 1702
rect 7818 1668 7856 1702
rect 7890 1668 7928 1702
rect 7962 1668 8000 1702
rect 8034 1668 8072 1702
rect 8106 1668 8144 1702
rect 8178 1668 8216 1702
rect 8250 1668 8288 1702
rect 8322 1668 8360 1702
rect 8394 1668 8432 1702
rect 8466 1668 8504 1702
rect 8538 1668 8576 1702
rect 8610 1668 8648 1702
rect 8682 1668 8720 1702
rect 8754 1668 8792 1702
rect 8826 1668 8864 1702
rect 8898 1668 8936 1702
rect 8970 1668 9008 1702
rect 9042 1668 9080 1702
rect 9114 1668 9152 1702
rect 9186 1668 9224 1702
rect 9258 1668 9296 1702
rect 9330 1668 9368 1702
rect 9402 1668 9440 1702
rect 9474 1668 9512 1702
rect 9546 1668 9584 1702
rect 9618 1668 9656 1702
rect 9690 1668 9728 1702
rect 9762 1668 9800 1702
rect 9834 1668 9872 1702
rect 9906 1668 9944 1702
rect 9978 1668 10016 1702
rect 10050 1668 10088 1702
rect 10122 1668 10160 1702
rect 10194 1668 10232 1702
rect 10266 1668 10304 1702
rect 10338 1668 10376 1702
rect 10410 1668 10448 1702
rect 10482 1668 10520 1702
rect 10554 1668 10592 1702
rect 10626 1668 10664 1702
rect 10698 1668 10736 1702
rect 10770 1668 10808 1702
rect 10842 1668 10880 1702
rect 10914 1668 10952 1702
rect 10986 1668 11024 1702
rect 11058 1668 11096 1702
rect 11130 1668 11168 1702
rect 11202 1668 11240 1702
rect 11274 1668 11312 1702
rect 11346 1668 11384 1702
rect 11418 1668 11456 1702
rect 11490 1668 11528 1702
rect 11562 1668 11600 1702
rect 11634 1668 11672 1702
rect 11706 1668 11744 1702
rect 11778 1668 11816 1702
rect 11850 1668 11888 1702
rect 11922 1668 11960 1702
rect 11994 1668 12032 1702
rect 12066 1668 12104 1702
rect 12138 1668 12176 1702
rect 12210 1668 12248 1702
rect 12282 1668 12320 1702
rect 12354 1668 12392 1702
rect 12426 1668 12464 1702
rect 12498 1668 12536 1702
rect 12570 1668 12608 1702
rect 12642 1668 12680 1702
rect 12714 1668 12752 1702
rect 12786 1668 12824 1702
rect 12858 1668 12896 1702
rect 12930 1668 12968 1702
rect 13002 1668 13040 1702
rect 13074 1668 13112 1702
rect 13146 1668 13184 1702
rect 13218 1668 13256 1702
rect 13290 1668 13328 1702
rect 13362 1668 13400 1702
rect 13434 1668 13472 1702
rect 13506 1668 13544 1702
rect 13578 1668 13616 1702
rect 13650 1668 13688 1702
rect 13722 1668 13760 1702
rect 13794 1668 13832 1702
rect 13866 1668 13904 1702
rect 13938 1668 13976 1702
rect 14010 1668 14048 1702
rect 14082 1668 14120 1702
rect 14154 1668 14192 1702
rect 14226 1668 14264 1702
rect 14298 1668 14336 1702
rect 14370 1668 14408 1702
rect 14442 1668 14480 1702
rect 14514 1668 14552 1702
rect 14586 1668 14624 1702
rect 14658 1668 14696 1702
rect 14730 1668 14768 1702
rect 14802 1668 14840 1702
rect 14874 1668 14912 1702
rect 14946 1668 14984 1702
rect 15018 1668 15056 1702
rect 15090 1668 15128 1702
rect 15162 1668 15200 1702
rect 15234 1668 15272 1702
rect 15306 1668 15344 1702
rect 15378 1668 15416 1702
rect 15450 1668 15488 1702
rect 15522 1668 15561 1702
rect 15595 1668 15634 1702
rect 15668 1668 15707 1702
rect 15741 1668 15780 1702
rect 15814 1668 15853 1702
rect 15887 1668 15926 1702
rect 15960 1668 15999 1702
rect 16033 1668 16072 1702
rect 16106 1668 16145 1702
rect 16179 1668 16218 1702
rect 16252 1668 16291 1702
rect 16325 1668 16364 1702
rect 16398 1668 16437 1702
rect 16471 1668 16510 1702
rect 16544 1668 16583 1702
rect 16617 1668 16656 1702
rect 16690 1668 17128 1702
rect 4615 1630 4627 1668
rect 4679 1630 4691 1668
rect 4743 1630 17128 1668
rect -2844 1591 -2832 1625
rect -2798 1591 -2759 1625
rect -2725 1591 -2686 1625
rect -2652 1591 -2613 1625
rect -2579 1591 -2540 1625
rect -2506 1591 -2467 1625
rect -2433 1591 -2394 1625
rect -2360 1591 -2321 1625
rect -2287 1591 -2248 1625
rect -2214 1591 -2175 1625
rect -2141 1591 -2102 1625
rect -2068 1591 -2029 1625
rect -1995 1591 -1956 1625
rect -1922 1591 -1883 1625
rect -1849 1591 -1810 1625
rect -1776 1591 -1737 1625
rect -2844 1553 -1737 1591
rect 4561 1624 17128 1630
rect 4561 1614 4616 1624
rect 4650 1614 4688 1624
rect 4722 1614 4760 1624
rect 4561 1562 4563 1614
rect 4615 1590 4616 1614
rect 4679 1590 4688 1614
rect 4743 1590 4760 1614
rect 4794 1590 4832 1624
rect 4866 1590 4904 1624
rect 4938 1590 4976 1624
rect 5010 1590 5048 1624
rect 5082 1590 5120 1624
rect 5154 1590 5192 1624
rect 5226 1590 5264 1624
rect 5298 1590 5336 1624
rect 5370 1590 5408 1624
rect 5442 1590 5480 1624
rect 5514 1590 5552 1624
rect 5586 1590 5624 1624
rect 5658 1590 5696 1624
rect 5730 1590 5768 1624
rect 5802 1590 5840 1624
rect 5874 1590 5912 1624
rect 5946 1590 5984 1624
rect 6018 1590 6056 1624
rect 6090 1590 6128 1624
rect 6162 1590 6200 1624
rect 6234 1590 6272 1624
rect 6306 1590 6344 1624
rect 6378 1590 6416 1624
rect 6450 1590 6488 1624
rect 6522 1590 6560 1624
rect 6594 1590 6632 1624
rect 6666 1590 6704 1624
rect 6738 1590 6776 1624
rect 6810 1590 6848 1624
rect 6882 1590 6920 1624
rect 6954 1590 6992 1624
rect 7026 1590 7064 1624
rect 7098 1590 7136 1624
rect 7170 1590 7208 1624
rect 7242 1590 7280 1624
rect 7314 1590 7352 1624
rect 7386 1590 7424 1624
rect 7458 1590 7496 1624
rect 7530 1590 7568 1624
rect 7602 1590 7640 1624
rect 7674 1590 7712 1624
rect 7746 1590 7784 1624
rect 7818 1590 7856 1624
rect 7890 1590 7928 1624
rect 7962 1590 8000 1624
rect 8034 1590 8072 1624
rect 8106 1590 8144 1624
rect 8178 1590 8216 1624
rect 8250 1590 8288 1624
rect 8322 1590 8360 1624
rect 8394 1590 8432 1624
rect 8466 1590 8504 1624
rect 8538 1590 8576 1624
rect 8610 1590 8648 1624
rect 8682 1590 8720 1624
rect 8754 1590 8792 1624
rect 8826 1590 8864 1624
rect 8898 1590 8936 1624
rect 8970 1590 9008 1624
rect 9042 1590 9080 1624
rect 9114 1590 9152 1624
rect 9186 1590 9224 1624
rect 9258 1590 9296 1624
rect 9330 1590 9368 1624
rect 9402 1590 9440 1624
rect 9474 1590 9512 1624
rect 9546 1590 9584 1624
rect 9618 1590 9656 1624
rect 9690 1590 9728 1624
rect 9762 1590 9800 1624
rect 9834 1590 9872 1624
rect 9906 1590 9944 1624
rect 9978 1590 10016 1624
rect 10050 1590 10088 1624
rect 10122 1590 10160 1624
rect 10194 1590 10232 1624
rect 10266 1590 10304 1624
rect 10338 1590 10376 1624
rect 10410 1590 10448 1624
rect 10482 1590 10520 1624
rect 10554 1590 10592 1624
rect 10626 1590 10664 1624
rect 10698 1590 10736 1624
rect 10770 1590 10808 1624
rect 10842 1590 10880 1624
rect 10914 1590 10952 1624
rect 10986 1590 11024 1624
rect 11058 1590 11096 1624
rect 11130 1590 11168 1624
rect 11202 1590 11240 1624
rect 11274 1590 11312 1624
rect 11346 1590 11384 1624
rect 11418 1590 11456 1624
rect 11490 1590 11528 1624
rect 11562 1590 11600 1624
rect 11634 1590 11672 1624
rect 11706 1590 11744 1624
rect 11778 1590 11816 1624
rect 11850 1590 11888 1624
rect 11922 1590 11960 1624
rect 11994 1590 12032 1624
rect 12066 1590 12104 1624
rect 12138 1590 12176 1624
rect 12210 1590 12248 1624
rect 12282 1590 12320 1624
rect 12354 1590 12392 1624
rect 12426 1590 12464 1624
rect 12498 1590 12536 1624
rect 12570 1590 12608 1624
rect 12642 1590 12680 1624
rect 12714 1590 12752 1624
rect 12786 1590 12824 1624
rect 12858 1590 12896 1624
rect 12930 1590 12968 1624
rect 13002 1590 13040 1624
rect 13074 1590 13112 1624
rect 13146 1590 13184 1624
rect 13218 1590 13256 1624
rect 13290 1590 13328 1624
rect 13362 1590 13400 1624
rect 13434 1590 13472 1624
rect 13506 1590 13544 1624
rect 13578 1590 13616 1624
rect 13650 1590 13688 1624
rect 13722 1590 13760 1624
rect 13794 1590 13832 1624
rect 13866 1590 13904 1624
rect 13938 1590 13976 1624
rect 14010 1590 14048 1624
rect 14082 1590 14120 1624
rect 14154 1590 14192 1624
rect 14226 1590 14264 1624
rect 14298 1590 14336 1624
rect 14370 1590 14408 1624
rect 14442 1590 14480 1624
rect 14514 1590 14552 1624
rect 14586 1590 14624 1624
rect 14658 1590 14696 1624
rect 14730 1590 14768 1624
rect 14802 1590 14840 1624
rect 14874 1590 14912 1624
rect 14946 1590 14984 1624
rect 15018 1590 15056 1624
rect 15090 1590 15128 1624
rect 15162 1590 15200 1624
rect 15234 1590 15272 1624
rect 15306 1590 15344 1624
rect 15378 1590 15416 1624
rect 15450 1590 15488 1624
rect 15522 1590 15561 1624
rect 15595 1590 15634 1624
rect 15668 1590 15707 1624
rect 15741 1590 15780 1624
rect 15814 1590 15853 1624
rect 15887 1590 15926 1624
rect 15960 1590 15999 1624
rect 16033 1590 16072 1624
rect 16106 1590 16145 1624
rect 16179 1590 16218 1624
rect 16252 1590 16291 1624
rect 16325 1590 16364 1624
rect 16398 1590 16437 1624
rect 16471 1590 16510 1624
rect 16544 1590 16583 1624
rect 16617 1590 16656 1624
rect 16690 1599 17128 1624
tri 17128 1599 17330 1801 sw
rect 16690 1590 17330 1599
rect 4615 1562 4627 1590
rect 4679 1562 4691 1590
rect 4743 1562 17330 1590
rect -2844 1519 -2832 1553
rect -2798 1519 -2759 1553
rect -2725 1519 -2686 1553
rect -2652 1519 -2613 1553
rect -2579 1519 -2540 1553
rect -2506 1519 -2467 1553
rect -2433 1519 -2394 1553
rect -2360 1519 -2321 1553
rect -2287 1519 -2248 1553
rect -2214 1519 -2175 1553
rect -2141 1519 -2102 1553
rect -2068 1519 -2029 1553
rect -1995 1519 -1956 1553
rect -1922 1519 -1883 1553
rect -1849 1519 -1810 1553
rect -1776 1519 -1737 1553
rect -2844 1481 -1737 1519
rect 4561 1546 17330 1562
rect 19429 1771 22725 1801
rect 19429 1719 19435 1771
rect 19487 1719 19504 1771
rect 19556 1719 19572 1771
rect 19624 1719 19640 1771
rect 19692 1719 19708 1771
rect 19760 1719 19776 1771
rect 19828 1719 19844 1771
rect 19896 1719 19912 1771
rect 19964 1719 19980 1771
rect 20032 1719 20048 1771
rect 20100 1719 20116 1771
rect 20168 1719 20184 1771
rect 20236 1719 20252 1771
rect 20304 1719 20844 1771
rect 20896 1719 20926 1771
rect 20978 1719 21008 1771
rect 21060 1719 21090 1771
rect 21142 1719 21550 1771
rect 21602 1719 21620 1771
rect 21672 1719 21690 1771
rect 21742 1719 21759 1771
rect 21811 1719 21828 1771
rect 21880 1719 21897 1771
rect 21949 1719 21966 1771
rect 22018 1719 22239 1771
rect 22291 1719 22309 1771
rect 22361 1719 22379 1771
rect 22431 1719 22448 1771
rect 22500 1719 22517 1771
rect 22569 1719 22586 1771
rect 22638 1719 22655 1771
rect 22707 1719 22725 1771
rect 19429 1707 22725 1719
rect 19429 1655 19435 1707
rect 19487 1655 19504 1707
rect 19556 1655 19572 1707
rect 19624 1655 19640 1707
rect 19692 1655 19708 1707
rect 19760 1655 19776 1707
rect 19828 1655 19844 1707
rect 19896 1655 19912 1707
rect 19964 1655 19980 1707
rect 20032 1655 20048 1707
rect 20100 1655 20116 1707
rect 20168 1655 20184 1707
rect 20236 1655 20252 1707
rect 20304 1655 20844 1707
rect 20896 1655 20926 1707
rect 20978 1655 21008 1707
rect 21060 1655 21090 1707
rect 21142 1655 21550 1707
rect 21602 1655 21620 1707
rect 21672 1655 21690 1707
rect 21742 1655 21759 1707
rect 21811 1655 21828 1707
rect 21880 1655 21897 1707
rect 21949 1655 21966 1707
rect 22018 1655 22239 1707
rect 22291 1655 22309 1707
rect 22361 1655 22379 1707
rect 22431 1655 22448 1707
rect 22500 1655 22517 1707
rect 22569 1655 22586 1707
rect 22638 1655 22655 1707
rect 22707 1655 22725 1707
rect 19429 1643 22725 1655
rect 19429 1591 19435 1643
rect 19487 1591 19504 1643
rect 19556 1591 19572 1643
rect 19624 1591 19640 1643
rect 19692 1591 19708 1643
rect 19760 1591 19776 1643
rect 19828 1591 19844 1643
rect 19896 1591 19912 1643
rect 19964 1591 19980 1643
rect 20032 1591 20048 1643
rect 20100 1591 20116 1643
rect 20168 1591 20184 1643
rect 20236 1591 20252 1643
rect 20304 1591 20844 1643
rect 20896 1591 20926 1643
rect 20978 1591 21008 1643
rect 21060 1591 21090 1643
rect 21142 1591 21550 1643
rect 21602 1591 21620 1643
rect 21672 1591 21690 1643
rect 21742 1591 21759 1643
rect 21811 1591 21828 1643
rect 21880 1591 21897 1643
rect 21949 1591 21966 1643
rect 22018 1591 22239 1643
rect 22291 1591 22309 1643
rect 22361 1591 22379 1643
rect 22431 1591 22448 1643
rect 22500 1591 22517 1643
rect 22569 1591 22586 1643
rect 22638 1591 22655 1643
rect 22707 1591 22725 1643
rect 19429 1560 22725 1591
rect 4561 1545 4616 1546
rect 4650 1545 4688 1546
rect 4722 1545 4760 1546
rect 4561 1493 4563 1545
rect 4615 1512 4616 1545
rect 4679 1512 4688 1545
rect 4743 1512 4760 1545
rect 4794 1512 4832 1546
rect 4866 1512 4904 1546
rect 4938 1512 4976 1546
rect 5010 1512 5048 1546
rect 5082 1512 5120 1546
rect 5154 1512 5192 1546
rect 5226 1512 5264 1546
rect 5298 1512 5336 1546
rect 5370 1512 5408 1546
rect 5442 1512 5480 1546
rect 5514 1512 5552 1546
rect 5586 1512 5624 1546
rect 5658 1512 5696 1546
rect 5730 1512 5768 1546
rect 5802 1512 5840 1546
rect 5874 1512 5912 1546
rect 5946 1512 5984 1546
rect 6018 1512 6056 1546
rect 6090 1512 6128 1546
rect 6162 1512 6200 1546
rect 6234 1512 6272 1546
rect 6306 1512 6344 1546
rect 6378 1512 6416 1546
rect 6450 1512 6488 1546
rect 6522 1512 6560 1546
rect 6594 1512 6632 1546
rect 6666 1512 6704 1546
rect 6738 1512 6776 1546
rect 6810 1512 6848 1546
rect 6882 1512 6920 1546
rect 6954 1512 6992 1546
rect 7026 1512 7064 1546
rect 7098 1512 7136 1546
rect 7170 1512 7208 1546
rect 7242 1512 7280 1546
rect 7314 1512 7352 1546
rect 7386 1512 7424 1546
rect 7458 1512 7496 1546
rect 7530 1512 7568 1546
rect 7602 1512 7640 1546
rect 7674 1512 7712 1546
rect 7746 1512 7784 1546
rect 7818 1512 7856 1546
rect 7890 1512 7928 1546
rect 7962 1512 8000 1546
rect 8034 1512 8072 1546
rect 8106 1512 8144 1546
rect 8178 1512 8216 1546
rect 8250 1512 8288 1546
rect 8322 1512 8360 1546
rect 8394 1512 8432 1546
rect 8466 1512 8504 1546
rect 8538 1512 8576 1546
rect 8610 1512 8648 1546
rect 8682 1512 8720 1546
rect 8754 1512 8792 1546
rect 8826 1512 8864 1546
rect 8898 1512 8936 1546
rect 8970 1512 9008 1546
rect 9042 1512 9080 1546
rect 9114 1512 9152 1546
rect 9186 1512 9224 1546
rect 9258 1512 9296 1546
rect 9330 1512 9368 1546
rect 9402 1512 9440 1546
rect 9474 1512 9512 1546
rect 9546 1512 9584 1546
rect 9618 1512 9656 1546
rect 9690 1512 9728 1546
rect 9762 1512 9800 1546
rect 9834 1512 9872 1546
rect 9906 1512 9944 1546
rect 9978 1512 10016 1546
rect 10050 1512 10088 1546
rect 10122 1512 10160 1546
rect 10194 1512 10232 1546
rect 10266 1512 10304 1546
rect 10338 1512 10376 1546
rect 10410 1512 10448 1546
rect 10482 1512 10520 1546
rect 10554 1512 10592 1546
rect 10626 1512 10664 1546
rect 10698 1512 10736 1546
rect 10770 1512 10808 1546
rect 10842 1512 10880 1546
rect 10914 1512 10952 1546
rect 10986 1512 11024 1546
rect 11058 1512 11096 1546
rect 11130 1512 11168 1546
rect 11202 1512 11240 1546
rect 11274 1512 11312 1546
rect 11346 1512 11384 1546
rect 11418 1512 11456 1546
rect 11490 1512 11528 1546
rect 11562 1512 11600 1546
rect 11634 1512 11672 1546
rect 11706 1512 11744 1546
rect 11778 1512 11816 1546
rect 11850 1512 11888 1546
rect 11922 1512 11960 1546
rect 11994 1512 12032 1546
rect 12066 1512 12104 1546
rect 12138 1512 12176 1546
rect 12210 1512 12248 1546
rect 12282 1512 12320 1546
rect 12354 1512 12392 1546
rect 12426 1512 12464 1546
rect 12498 1512 12536 1546
rect 12570 1512 12608 1546
rect 12642 1512 12680 1546
rect 12714 1512 12752 1546
rect 12786 1512 12824 1546
rect 12858 1512 12896 1546
rect 12930 1512 12968 1546
rect 13002 1512 13040 1546
rect 13074 1512 13112 1546
rect 13146 1512 13184 1546
rect 13218 1512 13256 1546
rect 13290 1512 13328 1546
rect 13362 1512 13400 1546
rect 13434 1512 13472 1546
rect 13506 1512 13544 1546
rect 13578 1512 13616 1546
rect 13650 1512 13688 1546
rect 13722 1512 13760 1546
rect 13794 1512 13832 1546
rect 13866 1512 13904 1546
rect 13938 1512 13976 1546
rect 14010 1512 14048 1546
rect 14082 1512 14120 1546
rect 14154 1512 14192 1546
rect 14226 1512 14264 1546
rect 14298 1512 14336 1546
rect 14370 1512 14408 1546
rect 14442 1512 14480 1546
rect 14514 1512 14552 1546
rect 14586 1512 14624 1546
rect 14658 1512 14696 1546
rect 14730 1512 14768 1546
rect 14802 1512 14840 1546
rect 14874 1512 14912 1546
rect 14946 1512 14984 1546
rect 15018 1512 15056 1546
rect 15090 1512 15128 1546
rect 15162 1512 15200 1546
rect 15234 1512 15272 1546
rect 15306 1512 15344 1546
rect 15378 1512 15416 1546
rect 15450 1512 15488 1546
rect 15522 1512 15561 1546
rect 15595 1512 15634 1546
rect 15668 1512 15707 1546
rect 15741 1512 15780 1546
rect 15814 1512 15853 1546
rect 15887 1512 15926 1546
rect 15960 1512 15999 1546
rect 16033 1512 16072 1546
rect 16106 1512 16145 1546
rect 16179 1512 16218 1546
rect 16252 1512 16291 1546
rect 16325 1512 16364 1546
rect 16398 1512 16437 1546
rect 16471 1512 16510 1546
rect 16544 1512 16583 1546
rect 16617 1512 16656 1546
rect 16690 1512 17330 1546
rect 4615 1493 4627 1512
rect 4679 1493 4691 1512
rect 4743 1493 17330 1512
rect -2844 1447 -2832 1481
rect -2798 1447 -2759 1481
rect -2725 1447 -2686 1481
rect -2652 1447 -2613 1481
rect -2579 1447 -2540 1481
rect -2506 1447 -2467 1481
rect -2433 1447 -2394 1481
rect -2360 1447 -2321 1481
rect -2287 1447 -2248 1481
rect -2214 1447 -2175 1481
rect -2141 1447 -2102 1481
rect -2068 1447 -2029 1481
rect -1995 1447 -1956 1481
rect -1922 1447 -1883 1481
rect -1849 1447 -1810 1481
rect -1776 1447 -1737 1481
rect -2844 1409 -1737 1447
rect 4561 1476 17330 1493
rect 4561 1424 4563 1476
rect 4615 1468 4627 1476
rect 4679 1468 4691 1476
rect 4743 1468 17330 1476
rect 4615 1434 4616 1468
rect 4679 1434 4688 1468
rect 4743 1434 4760 1468
rect 4794 1434 4832 1468
rect 4866 1434 4904 1468
rect 4938 1434 4976 1468
rect 5010 1434 5048 1468
rect 5082 1434 5120 1468
rect 5154 1434 5192 1468
rect 5226 1434 5264 1468
rect 5298 1434 5336 1468
rect 5370 1434 5408 1468
rect 5442 1434 5480 1468
rect 5514 1434 5552 1468
rect 5586 1434 5624 1468
rect 5658 1434 5696 1468
rect 5730 1434 5768 1468
rect 5802 1434 5840 1468
rect 5874 1434 5912 1468
rect 5946 1434 5984 1468
rect 6018 1434 6056 1468
rect 6090 1434 6128 1468
rect 6162 1434 6200 1468
rect 6234 1434 6272 1468
rect 6306 1434 6344 1468
rect 6378 1434 6416 1468
rect 6450 1434 6488 1468
rect 6522 1434 6560 1468
rect 6594 1434 6632 1468
rect 6666 1434 6704 1468
rect 6738 1434 6776 1468
rect 6810 1434 6848 1468
rect 6882 1434 6920 1468
rect 6954 1434 6992 1468
rect 7026 1434 7064 1468
rect 7098 1434 7136 1468
rect 7170 1434 7208 1468
rect 7242 1434 7280 1468
rect 7314 1434 7352 1468
rect 7386 1434 7424 1468
rect 7458 1434 7496 1468
rect 7530 1434 7568 1468
rect 7602 1434 7640 1468
rect 7674 1434 7712 1468
rect 7746 1434 7784 1468
rect 7818 1434 7856 1468
rect 7890 1434 7928 1468
rect 7962 1434 8000 1468
rect 8034 1434 8072 1468
rect 8106 1434 8144 1468
rect 8178 1434 8216 1468
rect 8250 1434 8288 1468
rect 8322 1434 8360 1468
rect 8394 1434 8432 1468
rect 8466 1434 8504 1468
rect 8538 1434 8576 1468
rect 8610 1434 8648 1468
rect 8682 1434 8720 1468
rect 8754 1434 8792 1468
rect 8826 1434 8864 1468
rect 8898 1434 8936 1468
rect 8970 1434 9008 1468
rect 9042 1434 9080 1468
rect 9114 1434 9152 1468
rect 9186 1434 9224 1468
rect 9258 1434 9296 1468
rect 9330 1434 9368 1468
rect 9402 1434 9440 1468
rect 9474 1434 9512 1468
rect 9546 1434 9584 1468
rect 9618 1434 9656 1468
rect 9690 1434 9728 1468
rect 9762 1434 9800 1468
rect 9834 1434 9872 1468
rect 9906 1434 9944 1468
rect 9978 1434 10016 1468
rect 10050 1434 10088 1468
rect 10122 1434 10160 1468
rect 10194 1434 10232 1468
rect 10266 1434 10304 1468
rect 10338 1434 10376 1468
rect 10410 1434 10448 1468
rect 10482 1434 10520 1468
rect 10554 1434 10592 1468
rect 10626 1434 10664 1468
rect 10698 1434 10736 1468
rect 10770 1434 10808 1468
rect 10842 1434 10880 1468
rect 10914 1434 10952 1468
rect 10986 1434 11024 1468
rect 11058 1434 11096 1468
rect 11130 1434 11168 1468
rect 11202 1434 11240 1468
rect 11274 1434 11312 1468
rect 11346 1434 11384 1468
rect 11418 1434 11456 1468
rect 11490 1434 11528 1468
rect 11562 1434 11600 1468
rect 11634 1434 11672 1468
rect 11706 1434 11744 1468
rect 11778 1434 11816 1468
rect 11850 1434 11888 1468
rect 11922 1434 11960 1468
rect 11994 1434 12032 1468
rect 12066 1434 12104 1468
rect 12138 1434 12176 1468
rect 12210 1434 12248 1468
rect 12282 1434 12320 1468
rect 12354 1434 12392 1468
rect 12426 1434 12464 1468
rect 12498 1434 12536 1468
rect 12570 1434 12608 1468
rect 12642 1434 12680 1468
rect 12714 1434 12752 1468
rect 12786 1434 12824 1468
rect 12858 1434 12896 1468
rect 12930 1434 12968 1468
rect 13002 1434 13040 1468
rect 13074 1434 13112 1468
rect 13146 1434 13184 1468
rect 13218 1434 13256 1468
rect 13290 1434 13328 1468
rect 13362 1434 13400 1468
rect 13434 1434 13472 1468
rect 13506 1434 13544 1468
rect 13578 1434 13616 1468
rect 13650 1434 13688 1468
rect 13722 1434 13760 1468
rect 13794 1434 13832 1468
rect 13866 1434 13904 1468
rect 13938 1434 13976 1468
rect 14010 1434 14048 1468
rect 14082 1434 14120 1468
rect 14154 1434 14192 1468
rect 14226 1434 14264 1468
rect 14298 1434 14336 1468
rect 14370 1434 14408 1468
rect 14442 1434 14480 1468
rect 14514 1434 14552 1468
rect 14586 1434 14624 1468
rect 14658 1434 14696 1468
rect 14730 1434 14768 1468
rect 14802 1434 14840 1468
rect 14874 1434 14912 1468
rect 14946 1434 14984 1468
rect 15018 1434 15056 1468
rect 15090 1434 15128 1468
rect 15162 1434 15200 1468
rect 15234 1434 15272 1468
rect 15306 1434 15344 1468
rect 15378 1434 15416 1468
rect 15450 1434 15488 1468
rect 15522 1434 15561 1468
rect 15595 1434 15634 1468
rect 15668 1434 15707 1468
rect 15741 1434 15780 1468
rect 15814 1434 15853 1468
rect 15887 1434 15926 1468
rect 15960 1434 15999 1468
rect 16033 1434 16072 1468
rect 16106 1434 16145 1468
rect 16179 1434 16218 1468
rect 16252 1434 16291 1468
rect 16325 1434 16364 1468
rect 16398 1434 16437 1468
rect 16471 1434 16510 1468
rect 16544 1434 16583 1468
rect 16617 1434 16656 1468
rect 16690 1434 17330 1468
rect 4615 1424 4627 1434
rect 4679 1424 4691 1434
rect 4743 1424 17330 1434
rect -2844 1375 -2832 1409
rect -2798 1375 -2759 1409
rect -2725 1375 -2686 1409
rect -2652 1375 -2613 1409
rect -2579 1375 -2540 1409
rect -2506 1375 -2467 1409
rect -2433 1375 -2394 1409
rect -2360 1375 -2321 1409
rect -2287 1375 -2248 1409
rect -2214 1375 -2175 1409
rect -2141 1375 -2102 1409
rect -2068 1375 -2029 1409
rect -1995 1375 -1956 1409
rect -1922 1375 -1883 1409
rect -1849 1375 -1810 1409
rect -1776 1375 -1737 1409
rect -2844 1337 -1737 1375
rect 4561 1407 17330 1424
rect 4561 1355 4563 1407
rect 4615 1355 4627 1407
rect 4679 1355 4691 1407
rect 4743 1393 17330 1407
rect 4743 1392 15560 1393
rect 5259 1358 5298 1392
rect 5332 1358 5371 1392
rect 5405 1358 5444 1392
rect 5478 1358 5517 1392
rect 5551 1358 5590 1392
rect 5624 1358 5663 1392
rect 5697 1358 5736 1392
rect 5770 1358 5809 1392
rect 5843 1358 5882 1392
rect 5916 1359 15560 1392
rect 15594 1359 15633 1393
rect 15667 1359 15706 1393
rect 15740 1359 15779 1393
rect 15813 1359 15852 1393
rect 15886 1359 15925 1393
rect 15959 1359 15998 1393
rect 16032 1359 16071 1393
rect 16105 1359 16144 1393
rect 16178 1359 16217 1393
rect 16251 1359 16290 1393
rect 16324 1359 16363 1393
rect 16397 1359 16436 1393
rect 16470 1359 16510 1393
rect 16544 1359 16584 1393
rect 16618 1359 16658 1393
rect 16692 1359 16732 1393
rect 16766 1359 16806 1393
rect 16840 1359 16880 1393
rect 16914 1359 17330 1393
rect 5916 1358 17330 1359
rect -2844 1303 -2832 1337
rect -2798 1303 -2759 1337
rect -2725 1303 -2686 1337
rect -2652 1303 -2613 1337
rect -2579 1303 -2540 1337
rect -2506 1303 -2467 1337
rect -2433 1303 -2394 1337
rect -2360 1303 -2321 1337
rect -2287 1303 -2248 1337
rect -2214 1303 -2175 1337
rect -2141 1303 -2102 1337
rect -2068 1303 -2029 1337
rect -1995 1303 -1956 1337
rect -1922 1303 -1883 1337
rect -1849 1303 -1810 1337
rect -1776 1303 -1737 1337
rect -2844 1265 -1737 1303
rect 4561 1338 4721 1355
rect 4561 1286 4563 1338
rect 4615 1286 4627 1338
rect 4679 1286 4691 1338
rect 5259 1320 17330 1358
rect 5259 1286 5298 1320
rect 5332 1286 5371 1320
rect 5405 1286 5444 1320
rect 5478 1286 5517 1320
rect 5551 1286 5590 1320
rect 5624 1286 5663 1320
rect 5697 1286 5736 1320
rect 5770 1286 5809 1320
rect 5843 1286 5882 1320
rect 5916 1319 17330 1320
rect 5916 1286 15560 1319
rect -2844 1231 -2832 1265
rect -2798 1231 -2759 1265
rect -2725 1231 -2686 1265
rect -2652 1231 -2613 1265
rect -2579 1231 -2540 1265
rect -2506 1231 -2467 1265
rect -2433 1231 -2394 1265
rect -2360 1231 -2321 1265
rect -2287 1231 -2248 1265
rect -2214 1231 -2175 1265
rect -2141 1231 -2102 1265
rect -2068 1231 -2029 1265
rect -1995 1231 -1956 1265
rect -1922 1231 -1883 1265
rect -1849 1231 -1810 1265
rect -1776 1231 -1737 1265
rect 4561 1269 4721 1286
rect 5259 1285 15560 1286
rect 15594 1285 15633 1319
rect 15667 1285 15706 1319
rect 15740 1285 15779 1319
rect 15813 1285 15852 1319
rect 15886 1285 15925 1319
rect 15959 1285 15998 1319
rect 16032 1285 16071 1319
rect 16105 1285 16144 1319
rect 16178 1285 16217 1319
rect 16251 1285 16290 1319
rect 16324 1285 16363 1319
rect 16397 1285 16436 1319
rect 16470 1285 16510 1319
rect 16544 1285 16584 1319
rect 16618 1285 16658 1319
rect 16692 1285 16732 1319
rect 16766 1285 16806 1319
rect 16840 1285 16880 1319
rect 16914 1285 17330 1319
rect 4561 1231 4563 1269
rect -2844 1230 1128 1231
rect 1180 1230 1192 1231
rect 1244 1230 1256 1231
rect 1308 1230 1320 1231
rect 1372 1230 4243 1231
rect -2844 1217 4243 1230
rect 4295 1217 4307 1231
rect 4359 1217 4371 1231
rect 4423 1217 4435 1231
rect 4487 1217 4499 1231
rect 4551 1217 4563 1231
rect 4615 1217 4627 1269
rect 4679 1217 4691 1269
rect 5259 1260 17330 1285
rect 5259 1248 13839 1260
rect -2844 1214 4721 1217
rect 5259 1214 5298 1248
rect 5332 1214 5371 1248
rect 5405 1214 5444 1248
rect 5478 1214 5517 1248
rect 5551 1214 5590 1248
rect 5624 1214 5663 1248
rect 5697 1214 5736 1248
rect 5770 1214 5809 1248
rect 5843 1214 5882 1248
rect 5916 1245 13839 1248
tri 13839 1245 13854 1260 nw
tri 15112 1245 15127 1260 ne
rect 15127 1245 17330 1260
rect 5916 1214 13805 1245
rect -2844 1211 13805 1214
tri 13805 1211 13839 1245 nw
tri 15127 1211 15161 1245 ne
rect 15161 1211 15560 1245
rect 15594 1211 15633 1245
rect 15667 1211 15706 1245
rect 15740 1211 15779 1245
rect 15813 1211 15852 1245
rect 15886 1211 15925 1245
rect 15959 1211 15998 1245
rect 16032 1211 16071 1245
rect 16105 1211 16144 1245
rect 16178 1211 16217 1245
rect 16251 1211 16290 1245
rect 16324 1211 16363 1245
rect 16397 1211 16436 1245
rect 16470 1211 16510 1245
rect 16544 1211 16584 1245
rect 16618 1211 16658 1245
rect 16692 1211 16732 1245
rect 16766 1211 16806 1245
rect 16840 1211 16880 1245
rect 16914 1211 17330 1245
rect -2844 1208 13801 1211
tri 109 1203 114 1208 ne
rect 114 1207 13801 1208
tri 13801 1207 13805 1211 nw
tri 15161 1207 15165 1211 ne
rect 15165 1207 17330 1211
rect 114 1204 13798 1207
tri 13798 1204 13801 1207 nw
tri 15165 1204 15168 1207 ne
rect 15168 1204 17330 1207
rect 114 1203 13797 1204
tri 13797 1203 13798 1204 nw
tri 15168 1203 15169 1204 ne
rect 15169 1203 17330 1204
rect 13919 1191 13971 1197
rect 13919 1127 13971 1139
rect 6924 1068 6930 1120
rect 6982 1068 6996 1120
rect 7048 1075 13919 1120
rect 7048 1069 13971 1075
rect 14004 1191 14726 1203
rect 14056 1151 14726 1191
rect 14778 1151 14790 1203
rect 14842 1151 14848 1203
rect 14004 1127 14056 1139
rect 14004 1069 14056 1075
rect 7048 1068 13967 1069
rect 14172 1068 14178 1120
rect 14230 1068 14242 1120
rect 14294 1068 14602 1120
rect 14654 1068 14666 1120
rect 14718 1068 14767 1120
rect -209 815 -203 867
rect -151 815 -139 867
rect -87 843 -81 867
tri -81 843 -57 867 sw
rect -87 815 6256 843
tri 6218 813 6220 815 ne
rect 6220 813 6256 815
tri 6256 813 6286 843 sw
rect 8632 822 10749 843
tri 6220 780 6253 813 ne
rect 6253 780 6286 813
tri 6286 780 6319 813 sw
tri 6253 779 6254 780 ne
rect 6254 779 6319 780
tri 6319 779 6320 780 sw
tri 6254 777 6256 779 ne
rect 6256 777 6320 779
tri 6256 760 6273 777 ne
rect 6273 760 6320 777
tri 6320 760 6339 779 sw
rect 8632 770 8639 822
rect 8691 813 8722 822
rect 8774 813 8805 822
rect 8857 813 8888 822
rect 8940 813 8971 822
rect 9023 813 9053 822
rect 9105 813 10749 822
rect 8691 779 8718 813
rect 8774 779 8792 813
rect 8857 779 8866 813
rect 9048 779 9053 813
rect 9122 779 9162 813
rect 9196 779 9236 813
rect 9270 779 9310 813
rect 9344 779 9384 813
rect 9418 779 9458 813
rect 9492 779 9532 813
rect 9566 779 9606 813
rect 9640 779 9680 813
rect 9714 779 9754 813
rect 9788 779 9827 813
rect 9861 779 9900 813
rect 9934 779 9973 813
rect 10007 779 10046 813
rect 10080 779 10119 813
rect 10153 779 10192 813
rect 10226 779 10265 813
rect 10299 779 10338 813
rect 10372 779 10411 813
rect 10445 779 10484 813
rect 10518 779 10557 813
rect 10591 779 10630 813
rect 10664 779 10703 813
rect 10737 779 10749 813
rect 15619 808 17330 820
rect 14672 800 14678 803
rect 8691 770 8722 779
rect 8774 770 8805 779
rect 8857 770 8888 779
rect 8940 770 8971 779
rect 9023 770 9053 779
rect 9105 770 10749 779
tri 6273 714 6319 760 ne
rect 6319 714 6339 760
tri 6339 714 6385 760 sw
rect 8632 749 10749 770
rect 14670 754 14678 800
rect 14672 751 14678 754
rect 14730 751 14742 803
rect 14794 751 14800 803
tri 6319 708 6325 714 ne
rect 6325 708 6864 714
tri 6325 674 6359 708 ne
rect 6359 674 6579 708
rect 6613 674 6659 708
rect 6693 674 6739 708
rect 6773 674 6818 708
rect 6852 674 6864 708
tri 6359 668 6365 674 ne
rect 6365 668 6864 674
tri 6918 636 6924 642 se
rect 6924 636 6930 642
rect 6510 630 6930 636
rect 6510 596 6522 630
rect 6556 596 6594 630
rect 6628 596 6930 630
rect 6510 590 6930 596
rect 6982 590 6996 642
rect 7048 590 7054 642
rect 14672 602 14678 605
rect 7423 508 7429 560
rect 7481 508 7493 560
rect 7545 508 7551 560
rect 14670 556 14678 602
rect 14672 553 14678 556
rect 14730 553 14742 605
rect 14794 553 14800 605
rect 9399 480 9412 508
tri 9412 480 9440 508 nw
rect 9169 428 9175 480
rect 9227 428 9239 480
rect 9291 428 9297 480
tri 9399 467 9412 480 nw
rect 13783 -200 13835 -194
rect 13783 -281 13835 -252
rect 13783 -339 13835 -333
rect 2758 -1094 3040 -1087
rect 2758 -1146 2764 -1094
rect 2816 -1146 2837 -1094
rect 2889 -1146 2910 -1094
rect 2962 -1146 2982 -1094
rect 3034 -1146 3040 -1094
rect 2758 -1158 3040 -1146
rect 2758 -1210 2764 -1158
rect 2816 -1210 2837 -1158
rect 2889 -1210 2910 -1158
rect 2962 -1210 2982 -1158
rect 3034 -1210 3040 -1158
rect 2758 -1222 3040 -1210
rect 2758 -1274 2764 -1222
rect 2816 -1274 2837 -1222
rect 2889 -1274 2910 -1222
rect 2962 -1274 2982 -1222
rect 3034 -1274 3040 -1222
rect 2758 -1281 3040 -1274
rect 15619 -1314 15648 808
rect 16546 425 17330 808
rect 16546 181 17086 425
tri 17086 181 17330 425 nw
rect 19429 436 22725 449
rect 19429 384 19443 436
rect 19495 384 19510 436
rect 19562 384 19577 436
rect 19629 384 19644 436
rect 19696 384 19711 436
rect 19763 384 19778 436
rect 19830 384 19845 436
rect 19897 384 19912 436
rect 19964 384 19979 436
rect 20031 384 20046 436
rect 20098 384 20113 436
rect 20165 384 20179 436
rect 20231 384 20245 436
rect 20297 384 20931 436
rect 20983 384 21011 436
rect 21063 384 21091 436
rect 21143 384 21171 436
rect 21223 384 21550 436
rect 21602 384 21619 436
rect 21671 384 21688 436
rect 21740 384 21757 436
rect 21809 384 21826 436
rect 21878 384 21895 436
rect 21947 384 21964 436
rect 22016 384 22235 436
rect 22287 384 22304 436
rect 22356 384 22373 436
rect 22425 384 22442 436
rect 22494 384 22511 436
rect 22563 384 22580 436
rect 22632 384 22649 436
rect 22701 384 22725 436
rect 19429 372 22725 384
rect 19429 320 19443 372
rect 19495 320 19510 372
rect 19562 320 19577 372
rect 19629 320 19644 372
rect 19696 320 19711 372
rect 19763 320 19778 372
rect 19830 320 19845 372
rect 19897 320 19912 372
rect 19964 320 19979 372
rect 20031 320 20046 372
rect 20098 320 20113 372
rect 20165 320 20179 372
rect 20231 320 20245 372
rect 20297 320 20931 372
rect 20983 320 21011 372
rect 21063 320 21091 372
rect 21143 320 21171 372
rect 21223 320 21550 372
rect 21602 320 21619 372
rect 21671 320 21688 372
rect 21740 320 21757 372
rect 21809 320 21826 372
rect 21878 320 21895 372
rect 21947 320 21964 372
rect 22016 320 22235 372
rect 22287 320 22304 372
rect 22356 320 22373 372
rect 22425 320 22442 372
rect 22494 320 22511 372
rect 22563 320 22580 372
rect 22632 320 22649 372
rect 22701 320 22725 372
rect 19429 308 22725 320
rect 19429 256 19443 308
rect 19495 256 19510 308
rect 19562 256 19577 308
rect 19629 256 19644 308
rect 19696 256 19711 308
rect 19763 256 19778 308
rect 19830 256 19845 308
rect 19897 256 19912 308
rect 19964 256 19979 308
rect 20031 256 20046 308
rect 20098 256 20113 308
rect 20165 256 20179 308
rect 20231 256 20245 308
rect 20297 256 20931 308
rect 20983 256 21011 308
rect 21063 256 21091 308
rect 21143 256 21171 308
rect 21223 256 21550 308
rect 21602 256 21619 308
rect 21671 256 21688 308
rect 21740 256 21757 308
rect 21809 256 21826 308
rect 21878 256 21895 308
rect 21947 256 21964 308
rect 22016 256 22235 308
rect 22287 256 22304 308
rect 22356 256 22373 308
rect 22425 256 22442 308
rect 22494 256 22511 308
rect 22563 256 22580 308
rect 22632 256 22649 308
rect 22701 256 22725 308
rect 19429 244 22725 256
rect 19429 192 19443 244
rect 19495 192 19510 244
rect 19562 192 19577 244
rect 19629 192 19644 244
rect 19696 192 19711 244
rect 19763 192 19778 244
rect 19830 192 19845 244
rect 19897 192 19912 244
rect 19964 192 19979 244
rect 20031 192 20046 244
rect 20098 192 20113 244
rect 20165 192 20179 244
rect 20231 192 20245 244
rect 20297 192 20931 244
rect 20983 192 21011 244
rect 21063 192 21091 244
rect 21143 192 21171 244
rect 21223 192 21550 244
rect 21602 192 21619 244
rect 21671 192 21688 244
rect 21740 192 21757 244
rect 21809 192 21826 244
rect 21878 192 21895 244
rect 21947 192 21964 244
rect 22016 192 22235 244
rect 22287 192 22304 244
rect 22356 192 22373 244
rect 22425 192 22442 244
rect 22494 192 22511 244
rect 22563 192 22580 244
rect 22632 192 22649 244
rect 22701 192 22725 244
rect 19429 181 22725 192
rect 23822 229 23874 235
rect 16546 -1314 16575 181
tri 16575 -330 17086 181 nw
rect 23822 165 23874 177
rect 23822 107 23874 113
rect 17162 -1070 17248 -1018
rect 17162 -1184 17248 -1132
rect 15619 -1353 16575 -1314
rect 15619 -1387 15648 -1353
rect 15682 -1387 15720 -1353
rect 15754 -1387 15792 -1353
rect 15826 -1387 15864 -1353
rect 15898 -1387 15936 -1353
rect 15970 -1387 16008 -1353
rect 16042 -1387 16080 -1353
rect 16114 -1387 16152 -1353
rect 16186 -1387 16224 -1353
rect 16258 -1387 16296 -1353
rect 16330 -1387 16368 -1353
rect 16402 -1387 16440 -1353
rect 16474 -1387 16512 -1353
rect 16546 -1387 16575 -1353
rect 15619 -1426 16575 -1387
rect 15619 -1460 15648 -1426
rect 15682 -1460 15720 -1426
rect 15754 -1460 15792 -1426
rect 15826 -1460 15864 -1426
rect 15898 -1460 15936 -1426
rect 15970 -1460 16008 -1426
rect 16042 -1460 16080 -1426
rect 16114 -1460 16152 -1426
rect 16186 -1460 16224 -1426
rect 16258 -1460 16296 -1426
rect 16330 -1460 16368 -1426
rect 16402 -1460 16440 -1426
rect 16474 -1460 16512 -1426
rect 16546 -1460 16575 -1426
rect 15619 -1499 16575 -1460
rect 15619 -1533 15648 -1499
rect 15682 -1533 15720 -1499
rect 15754 -1533 15792 -1499
rect 15826 -1533 15864 -1499
rect 15898 -1533 15936 -1499
rect 15970 -1533 16008 -1499
rect 16042 -1533 16080 -1499
rect 16114 -1533 16152 -1499
rect 16186 -1533 16224 -1499
rect 16258 -1533 16296 -1499
rect 16330 -1533 16368 -1499
rect 16402 -1533 16440 -1499
rect 16474 -1533 16512 -1499
rect 16546 -1533 16575 -1499
rect 2755 -1575 3041 -1571
rect 2755 -1627 2761 -1575
rect 2813 -1627 2835 -1575
rect 2887 -1627 2909 -1575
rect 2961 -1627 2983 -1575
rect 3035 -1627 3041 -1575
rect 2755 -1639 3041 -1627
rect 2755 -1691 2761 -1639
rect 2813 -1691 2835 -1639
rect 2887 -1691 2909 -1639
rect 2961 -1691 2983 -1639
rect 3035 -1691 3041 -1639
rect 15619 -1572 16575 -1533
rect 15619 -1606 15648 -1572
rect 15682 -1606 15720 -1572
rect 15754 -1606 15792 -1572
rect 15826 -1606 15864 -1572
rect 15898 -1606 15936 -1572
rect 15970 -1606 16008 -1572
rect 16042 -1606 16080 -1572
rect 16114 -1606 16152 -1572
rect 16186 -1606 16224 -1572
rect 16258 -1606 16296 -1572
rect 16330 -1606 16368 -1572
rect 16402 -1606 16440 -1572
rect 16474 -1606 16512 -1572
rect 16546 -1606 16575 -1572
rect 15619 -1645 16575 -1606
rect 15619 -1679 15648 -1645
rect 15682 -1679 15720 -1645
rect 15754 -1679 15792 -1645
rect 15826 -1679 15864 -1645
rect 15898 -1679 15936 -1645
rect 15970 -1679 16008 -1645
rect 16042 -1679 16080 -1645
rect 16114 -1679 16152 -1645
rect 16186 -1679 16224 -1645
rect 16258 -1679 16296 -1645
rect 16330 -1679 16368 -1645
rect 16402 -1679 16440 -1645
rect 16474 -1679 16512 -1645
rect 16546 -1679 16575 -1645
rect 15619 -1691 16575 -1679
rect 2755 -1695 3041 -1691
rect 2757 -2191 3041 -2187
rect 2757 -2243 2763 -2191
rect 2815 -2243 2837 -2191
rect 2889 -2243 2910 -2191
rect 2962 -2243 2983 -2191
rect 3035 -2243 3041 -2191
rect 2757 -2255 3041 -2243
rect 2757 -2307 2763 -2255
rect 2815 -2307 2837 -2255
rect 2889 -2307 2910 -2255
rect 2962 -2307 2983 -2255
rect 3035 -2307 3041 -2255
rect 17162 -2301 17229 -2249
rect 2757 -2311 3041 -2307
rect 17162 -2393 17231 -2341
rect 17162 -2533 17259 -2481
rect 17162 -2613 17259 -2561
tri 25410 -2938 25486 -2862 se
rect 25486 -2868 25538 -2862
rect 25486 -2932 25538 -2920
tri 17969 -2990 18021 -2938 se
rect 18021 -2984 25486 -2938
rect 18021 -2990 25538 -2984
tri 17967 -2992 17969 -2990 se
rect 17969 -2992 18041 -2990
tri 18041 -2992 18043 -2990 nw
rect 17432 -3044 17438 -2992
rect 17490 -3044 17502 -2992
rect 17554 -3044 17989 -2992
tri 17989 -3044 18041 -2992 nw
rect 16911 -3782 16963 -3736
<< via1 >>
rect 24087 26762 24139 26814
rect 24181 26762 24233 26814
rect 24274 26762 24326 26814
rect 24087 26698 24139 26750
rect 24181 26698 24233 26750
rect 24274 26698 24326 26750
rect 19271 22193 19323 22245
rect 19341 22193 19393 22245
rect 19411 22193 19463 22245
rect 19480 22193 19532 22245
rect 19549 22193 19601 22245
rect 19618 22193 19670 22245
rect 19687 22193 19739 22245
rect 19756 22193 19808 22245
rect 19825 22193 19877 22245
rect 19271 22129 19323 22181
rect 19341 22129 19393 22181
rect 19411 22129 19463 22181
rect 19480 22129 19532 22181
rect 19549 22129 19601 22181
rect 19618 22129 19670 22181
rect 19687 22129 19739 22181
rect 19756 22129 19808 22181
rect 19825 22129 19877 22181
rect 21012 22193 21064 22245
rect 21079 22193 21131 22245
rect 21146 22193 21198 22245
rect 21213 22193 21265 22245
rect 21280 22193 21332 22245
rect 21347 22193 21399 22245
rect 21414 22193 21466 22245
rect 21481 22193 21533 22245
rect 21548 22193 21600 22245
rect 21615 22193 21667 22245
rect 21681 22193 21733 22245
rect 21747 22193 21799 22245
rect 21813 22193 21865 22245
rect 21012 22129 21064 22181
rect 21079 22129 21131 22181
rect 21146 22129 21198 22181
rect 21213 22129 21265 22181
rect 21280 22129 21332 22181
rect 21347 22129 21399 22181
rect 21414 22129 21466 22181
rect 21481 22129 21533 22181
rect 21548 22129 21600 22181
rect 21615 22129 21667 22181
rect 21681 22129 21733 22181
rect 21747 22129 21799 22181
rect 21813 22129 21865 22181
rect 17327 21955 17443 22071
rect 17482 21961 17598 22077
rect 17636 21961 17752 22077
rect 19347 21961 19463 22077
rect 20266 21827 20318 21879
rect 20355 21827 20407 21879
rect 20443 21827 20495 21879
rect 20266 21763 20318 21815
rect 20355 21763 20407 21815
rect 20443 21763 20495 21815
rect 23742 19733 23794 19785
rect 23806 19733 23858 19785
rect 20266 19649 20318 19701
rect 20355 19649 20407 19701
rect 20444 19649 20496 19701
rect 20266 19585 20318 19637
rect 20355 19585 20407 19637
rect 20444 19585 20496 19637
rect 19227 18730 19279 18782
rect 19294 18730 19346 18782
rect 19361 18730 19413 18782
rect 19428 18730 19480 18782
rect 19495 18730 19547 18782
rect 19562 18730 19614 18782
rect 19629 18730 19681 18782
rect 19696 18730 19748 18782
rect 19763 18730 19815 18782
rect 19830 18730 19882 18782
rect 19897 18730 19949 18782
rect 19964 18730 20016 18782
rect 20031 18730 20083 18782
rect 20098 18730 20150 18782
rect 20165 18730 20217 18782
rect 20232 18730 20284 18782
rect 20299 18730 20351 18782
rect 20366 18730 20418 18782
rect 20433 18730 20485 18782
rect 20500 18730 20552 18782
rect 19227 18666 19279 18718
rect 19294 18666 19346 18718
rect 19361 18666 19413 18718
rect 19428 18666 19480 18718
rect 19495 18666 19547 18718
rect 19562 18666 19614 18718
rect 19629 18666 19681 18718
rect 19696 18666 19748 18718
rect 19763 18666 19815 18718
rect 19830 18666 19882 18718
rect 19897 18666 19949 18718
rect 19964 18666 20016 18718
rect 20031 18666 20083 18718
rect 20098 18666 20150 18718
rect 20165 18666 20217 18718
rect 20232 18666 20284 18718
rect 20299 18666 20351 18718
rect 20366 18666 20418 18718
rect 20433 18666 20485 18718
rect 20500 18666 20552 18718
rect 19227 18602 19279 18654
rect 19294 18602 19346 18654
rect 19361 18602 19413 18654
rect 19428 18602 19480 18654
rect 19495 18602 19547 18654
rect 19562 18602 19614 18654
rect 19629 18602 19681 18654
rect 19696 18602 19748 18654
rect 19763 18602 19815 18654
rect 19830 18602 19882 18654
rect 19897 18602 19949 18654
rect 19964 18602 20016 18654
rect 20031 18602 20083 18654
rect 20098 18602 20150 18654
rect 20165 18602 20217 18654
rect 20232 18602 20284 18654
rect 20299 18602 20351 18654
rect 20366 18602 20418 18654
rect 20433 18602 20485 18654
rect 20500 18602 20552 18654
rect 19227 18538 19279 18590
rect 19294 18538 19346 18590
rect 19361 18538 19413 18590
rect 19428 18538 19480 18590
rect 19495 18538 19547 18590
rect 19562 18538 19614 18590
rect 19629 18538 19681 18590
rect 19696 18538 19748 18590
rect 19763 18538 19815 18590
rect 19830 18538 19882 18590
rect 19897 18538 19949 18590
rect 19964 18538 20016 18590
rect 20031 18538 20083 18590
rect 20098 18538 20150 18590
rect 20165 18538 20217 18590
rect 20232 18538 20284 18590
rect 20299 18538 20351 18590
rect 20366 18538 20418 18590
rect 20433 18538 20485 18590
rect 20500 18538 20552 18590
rect 21048 18729 21100 18781
rect 21117 18729 21169 18781
rect 21186 18729 21238 18781
rect 21254 18729 21306 18781
rect 21322 18729 21374 18781
rect 21390 18729 21442 18781
rect 21458 18729 21510 18781
rect 21526 18729 21578 18781
rect 21594 18729 21646 18781
rect 21662 18729 21714 18781
rect 21048 18665 21100 18717
rect 21117 18665 21169 18717
rect 21186 18665 21238 18717
rect 21254 18665 21306 18717
rect 21322 18665 21374 18717
rect 21390 18665 21442 18717
rect 21458 18665 21510 18717
rect 21526 18665 21578 18717
rect 21594 18665 21646 18717
rect 21662 18665 21714 18717
rect 21048 18601 21100 18653
rect 21117 18601 21169 18653
rect 21186 18601 21238 18653
rect 21254 18601 21306 18653
rect 21322 18601 21374 18653
rect 21390 18601 21442 18653
rect 21458 18601 21510 18653
rect 21526 18601 21578 18653
rect 21594 18601 21646 18653
rect 21662 18601 21714 18653
rect 21048 18537 21100 18589
rect 21117 18537 21169 18589
rect 21186 18537 21238 18589
rect 21254 18537 21306 18589
rect 21322 18537 21374 18589
rect 21390 18537 21442 18589
rect 21458 18537 21510 18589
rect 21526 18537 21578 18589
rect 21594 18537 21646 18589
rect 21662 18537 21714 18589
rect 31029 18739 31081 18791
rect 31093 18739 31145 18791
rect 31157 18739 31209 18791
rect 31221 18739 31273 18791
rect 31285 18739 31337 18791
rect 31349 18739 31401 18791
rect 31029 18672 31081 18724
rect 31093 18672 31145 18724
rect 31157 18672 31209 18724
rect 31221 18672 31273 18724
rect 31285 18672 31337 18724
rect 31349 18672 31401 18724
rect 31029 18605 31081 18657
rect 31093 18605 31145 18657
rect 31157 18605 31209 18657
rect 31221 18605 31273 18657
rect 31285 18605 31337 18657
rect 31349 18605 31401 18657
rect 31029 18538 31081 18590
rect 31093 18538 31145 18590
rect 31157 18538 31209 18590
rect 31221 18538 31273 18590
rect 31285 18538 31337 18590
rect 31349 18538 31401 18590
rect 31029 18471 31081 18523
rect 31093 18471 31145 18523
rect 31157 18471 31209 18523
rect 31221 18471 31273 18523
rect 31285 18471 31337 18523
rect 31349 18471 31401 18523
rect 31029 18404 31081 18456
rect 31093 18404 31145 18456
rect 31157 18404 31209 18456
rect 31221 18404 31273 18456
rect 31285 18404 31337 18456
rect 31349 18404 31401 18456
rect 31029 18337 31081 18389
rect 31093 18337 31145 18389
rect 31157 18337 31209 18389
rect 31221 18337 31273 18389
rect 31285 18337 31337 18389
rect 31349 18337 31401 18389
rect 31029 18270 31081 18322
rect 31093 18270 31145 18322
rect 31157 18270 31209 18322
rect 31221 18270 31273 18322
rect 31285 18270 31337 18322
rect 31349 18270 31401 18322
rect 31029 18203 31081 18255
rect 31093 18203 31145 18255
rect 31157 18203 31209 18255
rect 31221 18203 31273 18255
rect 31285 18203 31337 18255
rect 31349 18203 31401 18255
rect 31029 18136 31081 18188
rect 31093 18136 31145 18188
rect 31157 18136 31209 18188
rect 31221 18136 31273 18188
rect 31285 18136 31337 18188
rect 31349 18136 31401 18188
rect 31029 18069 31081 18121
rect 31093 18069 31145 18121
rect 31157 18069 31209 18121
rect 31221 18069 31273 18121
rect 31285 18069 31337 18121
rect 31349 18069 31401 18121
rect 23038 14365 23090 14417
rect 23102 14365 23154 14417
rect 23761 14365 23813 14417
rect 23825 14365 23877 14417
rect 19435 8031 19487 8083
rect 19503 8031 19555 8083
rect 19571 8031 19623 8083
rect 19639 8031 19691 8083
rect 19707 8031 19759 8083
rect 19775 8031 19827 8083
rect 19842 8031 19894 8083
rect 20844 8031 20896 8083
rect 20926 8031 20978 8083
rect 21008 8031 21060 8083
rect 21090 8031 21142 8083
rect 21634 8031 21686 8083
rect 21701 8031 21753 8083
rect 21768 8031 21820 8083
rect 21834 8031 21886 8083
rect 21900 8031 21952 8083
rect 21966 8031 22018 8083
rect 22239 8031 22291 8083
rect 22309 8031 22361 8083
rect 22379 8031 22431 8083
rect 22448 8031 22500 8083
rect 22517 8031 22569 8083
rect 22586 8031 22638 8083
rect 22655 8031 22707 8083
rect 19435 7967 19487 8019
rect 19503 7967 19555 8019
rect 19571 7967 19623 8019
rect 19639 7967 19691 8019
rect 19707 7967 19759 8019
rect 19775 7967 19827 8019
rect 19842 7967 19894 8019
rect 20844 7967 20896 8019
rect 20926 7967 20978 8019
rect 21008 7967 21060 8019
rect 21090 7967 21142 8019
rect 21634 7967 21686 8019
rect 21701 7967 21753 8019
rect 21768 7967 21820 8019
rect 21834 7967 21886 8019
rect 21900 7967 21952 8019
rect 21966 7967 22018 8019
rect 22239 7967 22291 8019
rect 22309 7967 22361 8019
rect 22379 7967 22431 8019
rect 22448 7967 22500 8019
rect 22517 7967 22569 8019
rect 22586 7967 22638 8019
rect 22655 7967 22707 8019
rect 19435 7903 19487 7955
rect 19503 7903 19555 7955
rect 19571 7903 19623 7955
rect 19639 7903 19691 7955
rect 19707 7903 19759 7955
rect 19775 7903 19827 7955
rect 19842 7903 19894 7955
rect 20844 7903 20896 7955
rect 20926 7903 20978 7955
rect 21008 7903 21060 7955
rect 21090 7903 21142 7955
rect 21634 7903 21686 7955
rect 21701 7903 21753 7955
rect 21768 7903 21820 7955
rect 21834 7903 21886 7955
rect 21900 7903 21952 7955
rect 21966 7903 22018 7955
rect 22239 7903 22291 7955
rect 22309 7903 22361 7955
rect 22379 7903 22431 7955
rect 22448 7903 22500 7955
rect 22517 7903 22569 7955
rect 22586 7903 22638 7955
rect 22655 7903 22707 7955
rect 22466 6184 22582 6300
rect -3209 4508 -3157 4560
rect -3209 4444 -3157 4496
rect -2889 4500 -2837 4552
rect -2889 4436 -2837 4488
rect -2809 4500 -2757 4552
rect -2809 4436 -2757 4488
rect -2729 4487 -2677 4539
rect -2729 4423 -2677 4475
rect -2569 4487 -2517 4539
rect -2569 4423 -2517 4475
rect 4126 4467 4153 4497
rect 4153 4467 4178 4497
rect 4196 4467 4229 4497
rect 4229 4467 4248 4497
rect 4126 4445 4178 4467
rect 4196 4445 4248 4467
rect 4266 4467 4271 4497
rect 4271 4467 4305 4497
rect 4305 4467 4318 4497
rect 4266 4445 4318 4467
rect 4336 4467 4347 4497
rect 4347 4467 4381 4497
rect 4381 4467 4388 4497
rect 4336 4445 4388 4467
rect 4406 4467 4423 4497
rect 4423 4467 4457 4497
rect 4457 4467 4458 4497
rect 4406 4445 4458 4467
rect 4476 4467 4499 4497
rect 4499 4467 4528 4497
rect 4476 4445 4528 4467
rect 4126 4425 4178 4432
rect 4196 4425 4248 4432
rect 4126 4391 4153 4425
rect 4153 4391 4178 4425
rect 4196 4391 4229 4425
rect 4229 4391 4248 4425
rect 4126 4380 4178 4391
rect 4196 4380 4248 4391
rect 4266 4425 4318 4432
rect 4266 4391 4271 4425
rect 4271 4391 4305 4425
rect 4305 4391 4318 4425
rect 4266 4380 4318 4391
rect 4336 4425 4388 4432
rect 4336 4391 4347 4425
rect 4347 4391 4381 4425
rect 4381 4391 4388 4425
rect 4336 4380 4388 4391
rect 4406 4425 4458 4432
rect 4406 4391 4423 4425
rect 4423 4391 4457 4425
rect 4457 4391 4458 4425
rect 4406 4380 4458 4391
rect 4476 4425 4528 4432
rect 4476 4391 4499 4425
rect 4499 4391 4528 4425
rect 4476 4380 4528 4391
rect 4126 4349 4178 4367
rect 4196 4349 4248 4367
rect 4126 4315 4153 4349
rect 4153 4315 4178 4349
rect 4196 4315 4229 4349
rect 4229 4315 4248 4349
rect 4266 4349 4318 4367
rect 4266 4315 4271 4349
rect 4271 4315 4305 4349
rect 4305 4315 4318 4349
rect 4336 4349 4388 4367
rect 4336 4315 4347 4349
rect 4347 4315 4381 4349
rect 4381 4315 4388 4349
rect 4406 4349 4458 4367
rect 4406 4315 4423 4349
rect 4423 4315 4457 4349
rect 4457 4315 4458 4349
rect 4476 4349 4528 4367
rect 4476 4315 4499 4349
rect 4499 4315 4528 4349
rect 4126 4273 4178 4302
rect 4196 4273 4248 4302
rect 4126 4250 4153 4273
rect 4153 4250 4178 4273
rect 4196 4250 4229 4273
rect 4229 4250 4248 4273
rect 4266 4273 4318 4302
rect 4266 4250 4271 4273
rect 4271 4250 4305 4273
rect 4305 4250 4318 4273
rect 4336 4273 4388 4302
rect 4336 4250 4347 4273
rect 4347 4250 4381 4273
rect 4381 4250 4388 4273
rect 4406 4273 4458 4302
rect 4406 4250 4423 4273
rect 4423 4250 4457 4273
rect 4457 4250 4458 4273
rect 4476 4273 4528 4302
rect 4476 4250 4499 4273
rect 4499 4250 4528 4273
rect 4126 4197 4178 4237
rect 4196 4197 4248 4237
rect 4126 4185 4153 4197
rect 4153 4185 4178 4197
rect 4196 4185 4229 4197
rect 4229 4185 4248 4197
rect 4266 4197 4318 4237
rect 4266 4185 4271 4197
rect 4271 4185 4305 4197
rect 4305 4185 4318 4197
rect 4336 4197 4388 4237
rect 4336 4185 4347 4197
rect 4347 4185 4381 4197
rect 4381 4185 4388 4197
rect 4406 4197 4458 4237
rect 4406 4185 4423 4197
rect 4423 4185 4457 4197
rect 4457 4185 4458 4197
rect 4476 4197 4528 4237
rect 4476 4185 4499 4197
rect 4499 4185 4528 4197
rect 4126 4163 4153 4171
rect 4153 4163 4178 4171
rect 4196 4163 4229 4171
rect 4229 4163 4248 4171
rect 4126 4121 4178 4163
rect 4196 4121 4248 4163
rect 4126 4119 4153 4121
rect 4153 4119 4178 4121
rect 4196 4119 4229 4121
rect 4229 4119 4248 4121
rect 4266 4163 4271 4171
rect 4271 4163 4305 4171
rect 4305 4163 4318 4171
rect 4266 4121 4318 4163
rect 4266 4119 4271 4121
rect 4271 4119 4305 4121
rect 4305 4119 4318 4121
rect 4336 4163 4347 4171
rect 4347 4163 4381 4171
rect 4381 4163 4388 4171
rect 4336 4121 4388 4163
rect 4336 4119 4347 4121
rect 4347 4119 4381 4121
rect 4381 4119 4388 4121
rect 4406 4163 4423 4171
rect 4423 4163 4457 4171
rect 4457 4163 4458 4171
rect 4406 4121 4458 4163
rect 4406 4119 4423 4121
rect 4423 4119 4457 4121
rect 4457 4119 4458 4121
rect 4476 4163 4499 4171
rect 4499 4163 4528 4171
rect 4476 4121 4528 4163
rect 4476 4119 4499 4121
rect 4499 4119 4528 4121
rect 4126 4087 4153 4105
rect 4153 4087 4178 4105
rect 4196 4087 4229 4105
rect 4229 4087 4248 4105
rect -8 4031 44 4043
rect -8 3997 -4 4031
rect -4 3997 30 4031
rect 30 3997 44 4031
rect -8 3991 44 3997
rect 56 4031 108 4043
rect 56 3997 68 4031
rect 68 3997 102 4031
rect 102 3997 108 4031
rect 56 3991 108 3997
rect 1627 4015 1679 4067
rect 1708 4015 1760 4067
rect 4126 4053 4178 4087
rect 4196 4053 4248 4087
rect 4266 4087 4271 4105
rect 4271 4087 4305 4105
rect 4305 4087 4318 4105
rect 4266 4053 4318 4087
rect 4336 4087 4347 4105
rect 4347 4087 4381 4105
rect 4381 4087 4388 4105
rect 4336 4053 4388 4087
rect 4406 4087 4423 4105
rect 4423 4087 4457 4105
rect 4457 4087 4458 4105
rect 4406 4053 4458 4087
rect 4476 4087 4499 4105
rect 4499 4087 4528 4105
rect 4476 4053 4528 4087
rect 6268 4083 6320 4135
rect 6344 4083 6396 4135
rect 8408 4083 8460 4135
rect 8472 4083 8524 4135
rect 4126 4011 4153 4039
rect 4153 4011 4178 4039
rect 4196 4011 4229 4039
rect 4229 4011 4248 4039
rect 4126 3987 4178 4011
rect 4196 3987 4248 4011
rect 4266 4011 4271 4039
rect 4271 4011 4305 4039
rect 4305 4011 4318 4039
rect 4266 3987 4318 4011
rect 4336 4011 4347 4039
rect 4347 4011 4381 4039
rect 4381 4011 4388 4039
rect 4336 3987 4388 4011
rect 4406 4011 4423 4039
rect 4423 4011 4457 4039
rect 4457 4011 4458 4039
rect 4406 3987 4458 4011
rect 4476 4011 4499 4039
rect 4499 4011 4528 4039
rect 4476 3987 4528 4011
rect 4126 3968 4178 3973
rect 4196 3968 4248 3973
rect 4126 3934 4153 3968
rect 4153 3934 4178 3968
rect 4196 3934 4229 3968
rect 4229 3934 4248 3968
rect 4126 3921 4178 3934
rect 4196 3921 4248 3934
rect 4266 3968 4318 3973
rect 4266 3934 4271 3968
rect 4271 3934 4305 3968
rect 4305 3934 4318 3968
rect 4266 3921 4318 3934
rect 4336 3968 4388 3973
rect 4336 3934 4347 3968
rect 4347 3934 4381 3968
rect 4381 3934 4388 3968
rect 4336 3921 4388 3934
rect 4406 3968 4458 3973
rect 4406 3934 4423 3968
rect 4423 3934 4457 3968
rect 4457 3934 4458 3968
rect 4406 3921 4458 3934
rect 4476 3968 4528 3973
rect 4476 3934 4499 3968
rect 4499 3934 4528 3968
rect 4476 3921 4528 3934
rect 4126 3891 4178 3907
rect 4196 3891 4248 3907
rect 4126 3857 4153 3891
rect 4153 3857 4178 3891
rect 4196 3857 4229 3891
rect 4229 3857 4248 3891
rect 4126 3855 4178 3857
rect 4196 3855 4248 3857
rect 4266 3891 4318 3907
rect 4266 3857 4271 3891
rect 4271 3857 4305 3891
rect 4305 3857 4318 3891
rect 4266 3855 4318 3857
rect 4336 3891 4388 3907
rect 4336 3857 4347 3891
rect 4347 3857 4381 3891
rect 4381 3857 4388 3891
rect 4336 3855 4388 3857
rect 4406 3891 4458 3907
rect 4406 3857 4423 3891
rect 4423 3857 4457 3891
rect 4457 3857 4458 3891
rect 4406 3855 4458 3857
rect 4476 3891 4528 3907
rect 4476 3857 4499 3891
rect 4499 3857 4528 3891
rect 4476 3855 4528 3857
rect 6319 3609 6371 3661
rect 6383 3609 6435 3661
rect 9392 3609 9444 3661
rect 9456 3609 9508 3661
rect 8240 3523 8292 3575
rect 8304 3523 8356 3575
rect 10440 3438 10492 3490
rect 10504 3438 10556 3490
rect -3049 3367 -2997 3419
rect -203 3373 -151 3425
rect -139 3373 -87 3425
rect 39 3408 91 3410
rect 39 3374 45 3408
rect 45 3374 79 3408
rect 79 3374 91 3408
rect -3049 3303 -2997 3355
rect 39 3358 91 3374
rect 39 3336 91 3346
rect 39 3302 45 3336
rect 45 3302 79 3336
rect 79 3302 91 3336
rect 6330 3358 6382 3410
rect 6394 3358 6446 3410
rect 39 3294 91 3302
rect 9195 3121 9247 3173
rect 9259 3121 9311 3173
rect 1128 1780 1180 1832
rect 1192 1780 1244 1832
rect 1256 1780 1308 1832
rect 1320 1780 1372 1832
rect 1128 1712 1180 1764
rect 1192 1712 1244 1764
rect 1256 1712 1308 1764
rect 1320 1712 1372 1764
rect 4243 1698 4295 1750
rect 4307 1698 4359 1750
rect 4371 1698 4423 1750
rect 4435 1698 4487 1750
rect 4499 1698 4551 1750
rect 4563 1698 4615 1750
rect 4627 1746 4650 1750
rect 4650 1746 4679 1750
rect 4691 1746 4722 1750
rect 4722 1746 4743 1750
rect 4627 1702 4679 1746
rect 4691 1702 4743 1746
rect 4627 1698 4650 1702
rect 4650 1698 4679 1702
rect 4691 1698 4722 1702
rect 4722 1698 4743 1702
rect 1128 1644 1180 1696
rect 1192 1644 1244 1696
rect 1256 1644 1308 1696
rect 1320 1644 1372 1696
rect 4243 1630 4295 1682
rect 4307 1630 4359 1682
rect 4371 1630 4423 1682
rect 4435 1630 4487 1682
rect 4499 1630 4551 1682
rect 4563 1630 4615 1682
rect 4627 1668 4650 1682
rect 4650 1668 4679 1682
rect 4691 1668 4722 1682
rect 4722 1668 4743 1682
rect 4627 1630 4679 1668
rect 4691 1630 4743 1668
rect 1128 1575 1180 1627
rect 1192 1575 1244 1627
rect 1256 1575 1308 1627
rect 1320 1575 1372 1627
rect 4243 1562 4295 1614
rect 4307 1562 4359 1614
rect 4371 1562 4423 1614
rect 4435 1562 4487 1614
rect 4499 1562 4551 1614
rect 4563 1562 4615 1614
rect 4627 1590 4650 1614
rect 4650 1590 4679 1614
rect 4691 1590 4722 1614
rect 4722 1590 4743 1614
rect 4627 1562 4679 1590
rect 4691 1562 4743 1590
rect 1128 1506 1180 1558
rect 1192 1506 1244 1558
rect 1256 1506 1308 1558
rect 1320 1506 1372 1558
rect 19435 1719 19487 1771
rect 19504 1719 19556 1771
rect 19572 1719 19624 1771
rect 19640 1719 19692 1771
rect 19708 1719 19760 1771
rect 19776 1719 19828 1771
rect 19844 1719 19896 1771
rect 19912 1719 19964 1771
rect 19980 1719 20032 1771
rect 20048 1719 20100 1771
rect 20116 1719 20168 1771
rect 20184 1719 20236 1771
rect 20252 1719 20304 1771
rect 20844 1719 20896 1771
rect 20926 1719 20978 1771
rect 21008 1719 21060 1771
rect 21090 1719 21142 1771
rect 21550 1719 21602 1771
rect 21620 1719 21672 1771
rect 21690 1719 21742 1771
rect 21759 1719 21811 1771
rect 21828 1719 21880 1771
rect 21897 1719 21949 1771
rect 21966 1719 22018 1771
rect 22239 1719 22291 1771
rect 22309 1719 22361 1771
rect 22379 1719 22431 1771
rect 22448 1719 22500 1771
rect 22517 1719 22569 1771
rect 22586 1719 22638 1771
rect 22655 1719 22707 1771
rect 19435 1655 19487 1707
rect 19504 1655 19556 1707
rect 19572 1655 19624 1707
rect 19640 1655 19692 1707
rect 19708 1655 19760 1707
rect 19776 1655 19828 1707
rect 19844 1655 19896 1707
rect 19912 1655 19964 1707
rect 19980 1655 20032 1707
rect 20048 1655 20100 1707
rect 20116 1655 20168 1707
rect 20184 1655 20236 1707
rect 20252 1655 20304 1707
rect 20844 1655 20896 1707
rect 20926 1655 20978 1707
rect 21008 1655 21060 1707
rect 21090 1655 21142 1707
rect 21550 1655 21602 1707
rect 21620 1655 21672 1707
rect 21690 1655 21742 1707
rect 21759 1655 21811 1707
rect 21828 1655 21880 1707
rect 21897 1655 21949 1707
rect 21966 1655 22018 1707
rect 22239 1655 22291 1707
rect 22309 1655 22361 1707
rect 22379 1655 22431 1707
rect 22448 1655 22500 1707
rect 22517 1655 22569 1707
rect 22586 1655 22638 1707
rect 22655 1655 22707 1707
rect 19435 1591 19487 1643
rect 19504 1591 19556 1643
rect 19572 1591 19624 1643
rect 19640 1591 19692 1643
rect 19708 1591 19760 1643
rect 19776 1591 19828 1643
rect 19844 1591 19896 1643
rect 19912 1591 19964 1643
rect 19980 1591 20032 1643
rect 20048 1591 20100 1643
rect 20116 1591 20168 1643
rect 20184 1591 20236 1643
rect 20252 1591 20304 1643
rect 20844 1591 20896 1643
rect 20926 1591 20978 1643
rect 21008 1591 21060 1643
rect 21090 1591 21142 1643
rect 21550 1591 21602 1643
rect 21620 1591 21672 1643
rect 21690 1591 21742 1643
rect 21759 1591 21811 1643
rect 21828 1591 21880 1643
rect 21897 1591 21949 1643
rect 21966 1591 22018 1643
rect 22239 1591 22291 1643
rect 22309 1591 22361 1643
rect 22379 1591 22431 1643
rect 22448 1591 22500 1643
rect 22517 1591 22569 1643
rect 22586 1591 22638 1643
rect 22655 1591 22707 1643
rect 4243 1493 4295 1545
rect 4307 1493 4359 1545
rect 4371 1493 4423 1545
rect 4435 1493 4487 1545
rect 4499 1493 4551 1545
rect 4563 1493 4615 1545
rect 4627 1512 4650 1545
rect 4650 1512 4679 1545
rect 4691 1512 4722 1545
rect 4722 1512 4743 1545
rect 4627 1493 4679 1512
rect 4691 1493 4743 1512
rect 1128 1437 1180 1489
rect 1192 1437 1244 1489
rect 1256 1437 1308 1489
rect 1320 1437 1372 1489
rect 4243 1424 4295 1476
rect 4307 1424 4359 1476
rect 4371 1424 4423 1476
rect 4435 1424 4487 1476
rect 4499 1424 4551 1476
rect 4563 1424 4615 1476
rect 4627 1468 4679 1476
rect 4691 1468 4743 1476
rect 4627 1434 4650 1468
rect 4650 1434 4679 1468
rect 4691 1434 4722 1468
rect 4722 1434 4743 1468
rect 4627 1424 4679 1434
rect 4691 1424 4743 1434
rect 1128 1368 1180 1420
rect 1192 1368 1244 1420
rect 1256 1368 1308 1420
rect 1320 1368 1372 1420
rect 4243 1355 4295 1407
rect 4307 1355 4359 1407
rect 4371 1355 4423 1407
rect 4435 1355 4487 1407
rect 4499 1355 4551 1407
rect 4563 1355 4615 1407
rect 4627 1355 4679 1407
rect 4691 1392 4743 1407
rect 4691 1355 4721 1392
rect 4721 1355 4743 1392
rect 1128 1299 1180 1351
rect 1192 1299 1244 1351
rect 1256 1299 1308 1351
rect 1320 1299 1372 1351
rect 4243 1286 4295 1338
rect 4307 1286 4359 1338
rect 4371 1286 4423 1338
rect 4435 1286 4487 1338
rect 4499 1286 4551 1338
rect 4563 1286 4615 1338
rect 4627 1286 4679 1338
rect 4691 1286 4721 1338
rect 4721 1286 4743 1338
rect 1128 1231 1180 1282
rect 1192 1231 1244 1282
rect 1256 1231 1308 1282
rect 1320 1231 1372 1282
rect 4243 1231 4295 1269
rect 4307 1231 4359 1269
rect 4371 1231 4423 1269
rect 4435 1231 4487 1269
rect 4499 1231 4551 1269
rect 1128 1230 1180 1231
rect 1192 1230 1244 1231
rect 1256 1230 1308 1231
rect 1320 1230 1372 1231
rect 4243 1217 4295 1231
rect 4307 1217 4359 1231
rect 4371 1217 4423 1231
rect 4435 1217 4487 1231
rect 4499 1217 4551 1231
rect 4563 1217 4615 1269
rect 4627 1217 4679 1269
rect 4691 1217 4721 1269
rect 4721 1217 4743 1269
rect 13919 1139 13971 1191
rect 6930 1068 6982 1120
rect 6996 1068 7048 1120
rect 13919 1075 13971 1127
rect 14004 1139 14056 1191
rect 14726 1151 14778 1203
rect 14790 1151 14842 1203
rect 14004 1075 14056 1127
rect 14178 1068 14230 1120
rect 14242 1068 14294 1120
rect 14602 1068 14654 1120
rect 14666 1068 14718 1120
rect -203 815 -151 867
rect -139 815 -87 867
rect 8639 813 8691 822
rect 8722 813 8774 822
rect 8805 813 8857 822
rect 8888 813 8940 822
rect 8971 813 9023 822
rect 9053 813 9105 822
rect 8639 779 8644 813
rect 8644 779 8678 813
rect 8678 779 8691 813
rect 8722 779 8752 813
rect 8752 779 8774 813
rect 8805 779 8826 813
rect 8826 779 8857 813
rect 8888 779 8900 813
rect 8900 779 8940 813
rect 8971 779 8974 813
rect 8974 779 9014 813
rect 9014 779 9023 813
rect 9053 779 9088 813
rect 9088 779 9105 813
rect 8639 770 8691 779
rect 8722 770 8774 779
rect 8805 770 8857 779
rect 8888 770 8940 779
rect 8971 770 9023 779
rect 9053 770 9105 779
rect 14678 794 14730 803
rect 14678 760 14682 794
rect 14682 760 14716 794
rect 14716 760 14730 794
rect 14678 751 14730 760
rect 14742 794 14794 803
rect 14742 760 14754 794
rect 14754 760 14788 794
rect 14788 760 14794 794
rect 14742 751 14794 760
rect 6930 590 6982 642
rect 6996 590 7048 642
rect 7429 508 7481 560
rect 7493 508 7545 560
rect 14678 596 14730 605
rect 14678 562 14682 596
rect 14682 562 14716 596
rect 14716 562 14730 596
rect 14678 553 14730 562
rect 14742 596 14794 605
rect 14742 562 14754 596
rect 14754 562 14788 596
rect 14788 562 14794 596
rect 14742 553 14794 562
rect 9175 428 9227 480
rect 9239 428 9291 480
rect 13783 -252 13835 -200
rect 13783 -333 13835 -281
rect 2764 -1146 2816 -1094
rect 2837 -1146 2889 -1094
rect 2910 -1146 2962 -1094
rect 2982 -1146 3034 -1094
rect 2764 -1210 2816 -1158
rect 2837 -1210 2889 -1158
rect 2910 -1210 2962 -1158
rect 2982 -1210 3034 -1158
rect 2764 -1274 2816 -1222
rect 2837 -1274 2889 -1222
rect 2910 -1274 2962 -1222
rect 2982 -1274 3034 -1222
rect 19443 384 19495 436
rect 19510 384 19562 436
rect 19577 384 19629 436
rect 19644 384 19696 436
rect 19711 384 19763 436
rect 19778 384 19830 436
rect 19845 384 19897 436
rect 19912 384 19964 436
rect 19979 384 20031 436
rect 20046 384 20098 436
rect 20113 384 20165 436
rect 20179 384 20231 436
rect 20245 384 20297 436
rect 20931 384 20983 436
rect 21011 384 21063 436
rect 21091 384 21143 436
rect 21171 384 21223 436
rect 21550 384 21602 436
rect 21619 384 21671 436
rect 21688 384 21740 436
rect 21757 384 21809 436
rect 21826 384 21878 436
rect 21895 384 21947 436
rect 21964 384 22016 436
rect 22235 384 22287 436
rect 22304 384 22356 436
rect 22373 384 22425 436
rect 22442 384 22494 436
rect 22511 384 22563 436
rect 22580 384 22632 436
rect 22649 384 22701 436
rect 19443 320 19495 372
rect 19510 320 19562 372
rect 19577 320 19629 372
rect 19644 320 19696 372
rect 19711 320 19763 372
rect 19778 320 19830 372
rect 19845 320 19897 372
rect 19912 320 19964 372
rect 19979 320 20031 372
rect 20046 320 20098 372
rect 20113 320 20165 372
rect 20179 320 20231 372
rect 20245 320 20297 372
rect 20931 320 20983 372
rect 21011 320 21063 372
rect 21091 320 21143 372
rect 21171 320 21223 372
rect 21550 320 21602 372
rect 21619 320 21671 372
rect 21688 320 21740 372
rect 21757 320 21809 372
rect 21826 320 21878 372
rect 21895 320 21947 372
rect 21964 320 22016 372
rect 22235 320 22287 372
rect 22304 320 22356 372
rect 22373 320 22425 372
rect 22442 320 22494 372
rect 22511 320 22563 372
rect 22580 320 22632 372
rect 22649 320 22701 372
rect 19443 256 19495 308
rect 19510 256 19562 308
rect 19577 256 19629 308
rect 19644 256 19696 308
rect 19711 256 19763 308
rect 19778 256 19830 308
rect 19845 256 19897 308
rect 19912 256 19964 308
rect 19979 256 20031 308
rect 20046 256 20098 308
rect 20113 256 20165 308
rect 20179 256 20231 308
rect 20245 256 20297 308
rect 20931 256 20983 308
rect 21011 256 21063 308
rect 21091 256 21143 308
rect 21171 256 21223 308
rect 21550 256 21602 308
rect 21619 256 21671 308
rect 21688 256 21740 308
rect 21757 256 21809 308
rect 21826 256 21878 308
rect 21895 256 21947 308
rect 21964 256 22016 308
rect 22235 256 22287 308
rect 22304 256 22356 308
rect 22373 256 22425 308
rect 22442 256 22494 308
rect 22511 256 22563 308
rect 22580 256 22632 308
rect 22649 256 22701 308
rect 19443 192 19495 244
rect 19510 192 19562 244
rect 19577 192 19629 244
rect 19644 192 19696 244
rect 19711 192 19763 244
rect 19778 192 19830 244
rect 19845 192 19897 244
rect 19912 192 19964 244
rect 19979 192 20031 244
rect 20046 192 20098 244
rect 20113 192 20165 244
rect 20179 192 20231 244
rect 20245 192 20297 244
rect 20931 192 20983 244
rect 21011 192 21063 244
rect 21091 192 21143 244
rect 21171 192 21223 244
rect 21550 192 21602 244
rect 21619 192 21671 244
rect 21688 192 21740 244
rect 21757 192 21809 244
rect 21826 192 21878 244
rect 21895 192 21947 244
rect 21964 192 22016 244
rect 22235 192 22287 244
rect 22304 192 22356 244
rect 22373 192 22425 244
rect 22442 192 22494 244
rect 22511 192 22563 244
rect 22580 192 22632 244
rect 22649 192 22701 244
rect 23822 177 23874 229
rect 23822 113 23874 165
rect 2761 -1627 2813 -1575
rect 2835 -1627 2887 -1575
rect 2909 -1627 2961 -1575
rect 2983 -1627 3035 -1575
rect 2761 -1691 2813 -1639
rect 2835 -1691 2887 -1639
rect 2909 -1691 2961 -1639
rect 2983 -1691 3035 -1639
rect 2763 -2243 2815 -2191
rect 2837 -2243 2889 -2191
rect 2910 -2243 2962 -2191
rect 2983 -2243 3035 -2191
rect 2763 -2307 2815 -2255
rect 2837 -2307 2889 -2255
rect 2910 -2307 2962 -2255
rect 2983 -2307 3035 -2255
rect 25486 -2920 25538 -2868
rect 25486 -2984 25538 -2932
rect 17438 -3044 17490 -2992
rect 17502 -3044 17554 -2992
<< metal2 >>
rect 29198 27541 29541 28480
rect 24078 27046 25734 27186
rect 24078 26845 24437 27046
tri 24437 26845 24638 27046 nw
rect 24078 26814 24334 26845
rect 24078 26762 24087 26814
rect 24139 26762 24181 26814
rect 24233 26762 24274 26814
rect 24326 26762 24334 26814
rect 24078 26750 24334 26762
rect 24078 26698 24087 26750
rect 24139 26698 24181 26750
rect 24233 26698 24274 26750
rect 24326 26698 24334 26750
tri 24334 26742 24437 26845 nw
tri 26660 26742 26763 26845 se
rect 26763 26742 26963 26845
tri 20022 24298 20050 24326 ne
rect 20050 24298 20618 24326
tri 20618 24298 20646 24326 nw
tri 20050 24090 20258 24298 ne
tri 4651 22257 5002 22608 se
rect 5002 22492 6565 22608
rect 5002 22257 6330 22492
tri 6330 22257 6565 22492 nw
tri 4639 22245 4651 22257 se
rect 4651 22245 6318 22257
tri 6318 22245 6330 22257 nw
tri 4597 22203 4639 22245 se
rect 4639 22203 6276 22245
tri 6276 22203 6318 22245 nw
tri 3969 22193 3979 22203 se
rect 3979 22193 6266 22203
tri 6266 22193 6276 22203 nw
rect 19254 22201 19263 22257
rect 19319 22245 19357 22257
rect 19413 22245 19450 22257
rect 19506 22245 19543 22257
rect 19599 22245 19636 22257
rect 19692 22245 19729 22257
rect 19785 22245 19822 22257
rect 19254 22193 19271 22201
rect 19323 22193 19341 22245
rect 19532 22201 19543 22245
rect 19393 22193 19411 22201
rect 19463 22193 19480 22201
rect 19532 22193 19549 22201
rect 19601 22193 19618 22245
rect 19808 22201 19822 22245
rect 19878 22201 19887 22257
rect 19670 22193 19687 22201
rect 19739 22193 19756 22201
rect 19808 22193 19825 22201
rect 19877 22193 19887 22201
tri 3957 22181 3969 22193 se
rect 3969 22181 6254 22193
tri 6254 22181 6266 22193 nw
rect 19254 22181 19887 22193
tri 3905 22129 3957 22181 se
rect 3957 22129 6202 22181
tri 6202 22129 6254 22181 nw
rect 19254 22177 19271 22181
tri 3853 22077 3905 22129 se
rect 3905 22077 6150 22129
tri 6150 22077 6202 22129 nw
tri 17423 22077 17475 22129 se
rect 17475 22077 17603 22129
rect 19254 22121 19263 22177
rect 19323 22129 19341 22181
rect 19393 22177 19411 22181
rect 19463 22177 19480 22181
rect 19532 22177 19549 22181
rect 19532 22129 19543 22177
rect 19601 22129 19618 22181
rect 19670 22177 19687 22181
rect 19739 22177 19756 22181
rect 19808 22177 19825 22181
rect 19877 22177 19887 22181
rect 19808 22129 19822 22177
rect 19319 22121 19357 22129
rect 19413 22121 19450 22129
rect 19506 22121 19543 22129
rect 19599 22121 19636 22129
rect 19692 22121 19729 22129
rect 19785 22121 19822 22129
rect 19878 22121 19887 22177
tri 3847 22071 3853 22077 se
rect 3853 22071 6144 22077
tri 6144 22071 6150 22077 nw
rect 17327 22071 17482 22077
tri 3731 21955 3847 22071 se
rect 3847 21955 6028 22071
tri 6028 21955 6144 22071 nw
rect 17443 21961 17482 22071
rect 17598 21961 17603 22077
rect 17443 21955 17603 21961
rect 17636 22077 17752 22083
rect 19341 21961 19347 22077
rect 19463 21961 19469 22077
rect 17636 21955 17752 21961
tri 3725 21949 3731 21955 se
rect 3731 21949 6022 21955
tri 6022 21949 6028 21955 nw
rect 17327 21949 17603 21955
tri 3655 21879 3725 21949 se
rect 3725 21879 5952 21949
tri 5952 21879 6022 21949 nw
rect 20258 21879 20504 24298
tri 20504 24184 20618 24298 nw
tri 3603 21827 3655 21879 se
rect 3655 21827 5900 21879
tri 5900 21827 5952 21879 nw
rect 20258 21827 20266 21879
rect 20318 21827 20355 21879
rect 20407 21827 20443 21879
rect 20495 21827 20504 21879
tri 3602 21826 3603 21827 se
rect 3603 21826 5899 21827
tri 5899 21826 5900 21827 nw
rect 3602 21815 5888 21826
tri 5888 21815 5899 21826 nw
rect 20258 21815 20504 21827
rect 3602 21763 5836 21815
tri 5836 21763 5888 21815 nw
rect 20258 21763 20266 21815
rect 20318 21763 20355 21815
rect 20407 21763 20443 21815
rect 20495 21763 20504 21815
rect 3602 21656 5729 21763
tri 5729 21656 5836 21763 nw
rect 17782 21612 18092 21652
rect 20258 19701 20504 21763
rect 20258 19649 20266 19701
rect 20318 19649 20355 19701
rect 20407 19649 20444 19701
rect 20496 19649 20504 19701
rect 20258 19637 20504 19649
rect 20258 19585 20266 19637
rect 20318 19585 20355 19637
rect 20407 19585 20444 19637
rect 20496 19585 20504 19637
rect 20258 19583 20504 19585
rect 19208 18807 20570 18809
rect 19208 18751 19217 18807
rect 19273 18782 19298 18807
rect 19354 18782 19379 18807
rect 19435 18782 19460 18807
rect 19516 18782 19541 18807
rect 19597 18782 19622 18807
rect 19678 18782 19703 18807
rect 19759 18782 19784 18807
rect 19840 18782 19865 18807
rect 19208 18730 19227 18751
rect 19279 18730 19294 18782
rect 19354 18751 19361 18782
rect 19614 18751 19622 18782
rect 19346 18730 19361 18751
rect 19413 18730 19428 18751
rect 19480 18730 19495 18751
rect 19547 18730 19562 18751
rect 19614 18730 19629 18751
rect 19681 18730 19696 18782
rect 19759 18751 19763 18782
rect 19748 18730 19763 18751
rect 19815 18730 19830 18751
rect 19208 18727 19865 18730
rect 19208 18671 19217 18727
rect 19273 18718 19298 18727
rect 19354 18718 19379 18727
rect 19435 18718 19460 18727
rect 19516 18718 19541 18727
rect 19597 18718 19622 18727
rect 19678 18718 19703 18727
rect 19759 18718 19784 18727
rect 19840 18718 19865 18727
rect 19208 18666 19227 18671
rect 19279 18666 19294 18718
rect 19354 18671 19361 18718
rect 19614 18671 19622 18718
rect 19346 18666 19361 18671
rect 19413 18666 19428 18671
rect 19480 18666 19495 18671
rect 19547 18666 19562 18671
rect 19614 18666 19629 18671
rect 19681 18666 19696 18718
rect 19759 18671 19763 18718
rect 19748 18666 19763 18671
rect 19815 18666 19830 18671
rect 19208 18654 19865 18666
rect 19208 18647 19227 18654
rect 19208 18591 19217 18647
rect 19279 18602 19294 18654
rect 19346 18647 19361 18654
rect 19413 18647 19428 18654
rect 19480 18647 19495 18654
rect 19547 18647 19562 18654
rect 19614 18647 19629 18654
rect 19354 18602 19361 18647
rect 19614 18602 19622 18647
rect 19681 18602 19696 18654
rect 19748 18647 19763 18654
rect 19815 18647 19830 18654
rect 19759 18602 19763 18647
rect 19273 18591 19298 18602
rect 19354 18591 19379 18602
rect 19435 18591 19460 18602
rect 19516 18591 19541 18602
rect 19597 18591 19622 18602
rect 19678 18591 19703 18602
rect 19759 18591 19784 18602
rect 19840 18591 19865 18602
rect 19208 18590 19865 18591
rect 19208 18567 19227 18590
rect 19208 18511 19217 18567
rect 19279 18538 19294 18590
rect 19346 18567 19361 18590
rect 19413 18567 19428 18590
rect 19480 18567 19495 18590
rect 19547 18567 19562 18590
rect 19614 18567 19629 18590
rect 19354 18538 19361 18567
rect 19614 18538 19622 18567
rect 19681 18538 19696 18590
rect 19748 18567 19763 18590
rect 19815 18567 19830 18590
rect 19759 18538 19763 18567
rect 19273 18511 19298 18538
rect 19354 18511 19379 18538
rect 19435 18511 19460 18538
rect 19516 18511 19541 18538
rect 19597 18511 19622 18538
rect 19678 18511 19703 18538
rect 19759 18511 19784 18538
rect 19840 18511 19865 18538
rect 20561 18511 20570 18807
rect 19208 18509 20570 18511
rect 20658 18157 20968 24298
rect 21002 22258 21874 22266
rect 21002 22202 21011 22258
rect 21067 22245 21100 22258
rect 21156 22245 21189 22258
rect 21245 22245 21278 22258
rect 21334 22245 21367 22258
rect 21423 22245 21456 22258
rect 21512 22245 21545 22258
rect 21601 22245 21633 22258
rect 21689 22245 21721 22258
rect 21777 22245 21809 22258
rect 21067 22202 21079 22245
rect 21265 22202 21278 22245
rect 21334 22202 21347 22245
rect 21533 22202 21545 22245
rect 21601 22202 21615 22245
rect 21799 22202 21809 22245
rect 21002 22193 21012 22202
rect 21064 22193 21079 22202
rect 21131 22193 21146 22202
rect 21198 22193 21213 22202
rect 21265 22193 21280 22202
rect 21332 22193 21347 22202
rect 21399 22193 21414 22202
rect 21466 22193 21481 22202
rect 21533 22193 21548 22202
rect 21600 22193 21615 22202
rect 21667 22193 21681 22202
rect 21733 22193 21747 22202
rect 21799 22193 21813 22202
rect 21865 22193 21874 22258
rect 21002 22181 21874 22193
rect 21002 22178 21012 22181
rect 21064 22178 21079 22181
rect 21131 22178 21146 22181
rect 21198 22178 21213 22181
rect 21265 22178 21280 22181
rect 21332 22178 21347 22181
rect 21399 22178 21414 22181
rect 21466 22178 21481 22181
rect 21533 22178 21548 22181
rect 21600 22178 21615 22181
rect 21667 22178 21681 22181
rect 21733 22178 21747 22181
rect 21799 22178 21813 22181
rect 21002 22122 21011 22178
rect 21067 22129 21079 22178
rect 21265 22129 21278 22178
rect 21334 22129 21347 22178
rect 21533 22129 21545 22178
rect 21601 22129 21615 22178
rect 21799 22129 21809 22178
rect 21067 22122 21100 22129
rect 21156 22122 21189 22129
rect 21245 22122 21278 22129
rect 21334 22122 21367 22129
rect 21423 22122 21456 22129
rect 21512 22122 21545 22129
rect 21601 22122 21633 22129
rect 21689 22122 21721 22129
rect 21777 22122 21809 22129
rect 21865 22122 21874 22181
rect 21002 22114 21874 22122
rect 23423 21185 23683 24270
rect 24078 22244 24334 26698
tri 26381 26463 26660 26742 se
rect 26660 26463 26963 26742
rect 23736 19733 23742 19785
rect 23794 19733 23806 19785
rect 23858 19733 23864 19785
tri 23736 19696 23773 19733 ne
rect 21039 18807 21724 18809
rect 21039 18729 21048 18807
rect 21104 18781 21136 18807
rect 21192 18781 21224 18807
rect 21280 18781 21311 18807
rect 21367 18781 21398 18807
rect 21454 18781 21485 18807
rect 21541 18781 21572 18807
rect 21628 18781 21659 18807
rect 21104 18751 21117 18781
rect 21306 18751 21311 18781
rect 21100 18729 21117 18751
rect 21169 18729 21186 18751
rect 21238 18729 21254 18751
rect 21306 18729 21322 18751
rect 21374 18729 21390 18781
rect 21454 18751 21458 18781
rect 21646 18751 21659 18781
rect 21715 18751 21724 18807
rect 21442 18729 21458 18751
rect 21510 18729 21526 18751
rect 21578 18729 21594 18751
rect 21646 18729 21662 18751
rect 21714 18729 21724 18751
rect 21039 18727 21724 18729
rect 21039 18665 21048 18727
rect 21104 18717 21136 18727
rect 21192 18717 21224 18727
rect 21280 18717 21311 18727
rect 21367 18717 21398 18727
rect 21454 18717 21485 18727
rect 21541 18717 21572 18727
rect 21628 18717 21659 18727
rect 21104 18671 21117 18717
rect 21306 18671 21311 18717
rect 21100 18665 21117 18671
rect 21169 18665 21186 18671
rect 21238 18665 21254 18671
rect 21306 18665 21322 18671
rect 21374 18665 21390 18717
rect 21454 18671 21458 18717
rect 21646 18671 21659 18717
rect 21715 18671 21724 18727
tri 23755 18683 23773 18701 se
rect 23773 18683 23813 19733
tri 23813 19696 23850 19733 nw
tri 23744 18672 23755 18683 se
rect 23755 18672 23802 18683
tri 23802 18672 23813 18683 nw
rect 24083 18802 24317 18811
rect 24083 18746 24092 18802
rect 24148 18746 24172 18802
rect 24228 18746 24252 18802
rect 24308 18746 24317 18802
rect 30985 18804 31435 18813
rect 24083 18689 24317 18746
rect 21442 18665 21458 18671
rect 21510 18665 21526 18671
rect 21578 18665 21594 18671
rect 21646 18665 21662 18671
rect 21714 18665 21724 18671
rect 21039 18653 21724 18665
tri 23729 18657 23744 18672 se
rect 23744 18657 23787 18672
tri 23787 18657 23802 18672 nw
rect 21039 18591 21048 18653
rect 21100 18647 21117 18653
rect 21169 18647 21186 18653
rect 21238 18647 21254 18653
rect 21306 18647 21322 18653
rect 21104 18601 21117 18647
rect 21306 18601 21311 18647
rect 21374 18601 21390 18653
rect 21442 18647 21458 18653
rect 21510 18647 21526 18653
rect 21578 18647 21594 18653
rect 21646 18647 21662 18653
rect 21714 18647 21724 18653
rect 21454 18601 21458 18647
rect 21646 18601 21659 18647
rect 21104 18591 21136 18601
rect 21192 18591 21224 18601
rect 21280 18591 21311 18601
rect 21367 18591 21398 18601
rect 21454 18591 21485 18601
rect 21541 18591 21572 18601
rect 21628 18591 21659 18601
rect 21715 18591 21724 18647
tri 23710 18638 23729 18657 se
rect 23729 18638 23768 18657
tri 23768 18638 23787 18657 nw
tri 23677 18605 23710 18638 se
rect 23710 18605 23735 18638
tri 23735 18605 23768 18638 nw
rect 24083 18633 24092 18689
rect 24148 18633 24172 18689
rect 24228 18633 24252 18689
rect 24308 18633 24317 18689
rect 21039 18589 21724 18591
tri 23662 18590 23677 18605 se
rect 23677 18590 23720 18605
tri 23720 18590 23735 18605 nw
rect 21039 18511 21048 18589
rect 21100 18567 21117 18589
rect 21169 18567 21186 18589
rect 21238 18567 21254 18589
rect 21306 18567 21322 18589
rect 21104 18537 21117 18567
rect 21306 18537 21311 18567
rect 21374 18537 21390 18589
rect 21442 18567 21458 18589
rect 21510 18567 21526 18589
rect 21578 18567 21594 18589
rect 21646 18567 21662 18589
rect 21714 18567 21724 18589
tri 23652 18580 23662 18590 se
rect 23662 18580 23710 18590
tri 23710 18580 23720 18590 nw
rect 21454 18537 21458 18567
rect 21646 18537 21659 18567
rect 21104 18511 21136 18537
rect 21192 18511 21224 18537
rect 21280 18511 21311 18537
rect 21367 18511 21398 18537
rect 21454 18511 21485 18537
rect 21541 18511 21572 18537
rect 21628 18511 21659 18537
rect 21715 18511 21724 18567
tri 23610 18538 23652 18580 se
rect 23652 18538 23668 18580
tri 23668 18538 23710 18580 nw
rect 24083 18575 24317 18633
tri 23595 18523 23610 18538 se
rect 23610 18523 23653 18538
tri 23653 18523 23668 18538 nw
tri 23594 18522 23595 18523 se
rect 23595 18522 23652 18523
tri 23652 18522 23653 18523 nw
rect 21039 18509 21724 18511
tri 23581 18509 23594 18522 se
rect 23594 18510 23640 18522
tri 23640 18510 23652 18522 nw
rect 24083 18519 24092 18575
rect 24148 18519 24172 18575
rect 24228 18519 24252 18575
rect 24308 18519 24317 18575
rect 24083 18510 24317 18519
rect 29456 18791 29816 18800
rect 29456 18735 29488 18791
rect 29544 18735 29568 18791
rect 29624 18735 29648 18791
rect 29704 18735 29728 18791
rect 29784 18735 29816 18791
rect 29456 18705 29816 18735
rect 29456 18649 29488 18705
rect 29544 18649 29568 18705
rect 29624 18649 29648 18705
rect 29704 18649 29728 18705
rect 29784 18649 29816 18705
rect 29456 18618 29816 18649
rect 29456 18562 29488 18618
rect 29544 18562 29568 18618
rect 29624 18562 29648 18618
rect 29704 18562 29728 18618
rect 29784 18562 29816 18618
rect 29456 18531 29816 18562
rect 23594 18509 23639 18510
tri 23639 18509 23640 18510 nw
tri 23543 18471 23581 18509 se
rect 23581 18471 23601 18509
tri 23601 18471 23639 18509 nw
rect 29456 18475 29488 18531
rect 29544 18475 29568 18531
rect 29624 18475 29648 18531
rect 29704 18475 29728 18531
rect 29784 18475 29816 18531
tri 23536 18464 23543 18471 se
rect 23543 18464 23594 18471
tri 23594 18464 23601 18471 nw
tri 23528 18456 23536 18464 se
rect 23536 18456 23586 18464
tri 23586 18456 23594 18464 nw
tri 23478 18406 23528 18456 se
rect 23528 18406 23536 18456
tri 23536 18406 23586 18456 nw
rect 29456 18444 29816 18475
tri 23476 18404 23478 18406 se
rect 23478 18404 23534 18406
tri 23534 18404 23536 18406 nw
tri 23461 18389 23476 18404 se
rect 23476 18389 23519 18404
tri 23519 18389 23534 18404 nw
tri 23420 18348 23461 18389 se
rect 23461 18348 23478 18389
tri 23478 18348 23519 18389 nw
rect 29456 18388 29488 18444
rect 29544 18388 29568 18444
rect 29624 18388 29648 18444
rect 29704 18388 29728 18444
rect 29784 18388 29816 18444
rect 29456 18357 29816 18388
tri 23409 18337 23420 18348 se
rect 23420 18337 23467 18348
tri 23467 18337 23478 18348 nw
tri 23394 18322 23409 18337 se
rect 23409 18322 23452 18337
tri 23452 18322 23467 18337 nw
tri 23362 18290 23394 18322 se
rect 23394 18290 23420 18322
tri 23420 18290 23452 18322 nw
rect 29456 18301 29488 18357
rect 29544 18301 29568 18357
rect 29624 18301 29648 18357
rect 29704 18301 29728 18357
rect 29784 18301 29816 18357
tri 23342 18270 23362 18290 se
rect 23362 18270 23400 18290
tri 23400 18270 23420 18290 nw
rect 29456 18270 29816 18301
tri 23327 18255 23342 18270 se
rect 23342 18255 23385 18270
tri 23385 18255 23400 18270 nw
tri 23304 18232 23327 18255 se
rect 23327 18232 23362 18255
tri 23362 18232 23385 18255 nw
tri 23275 18203 23304 18232 se
rect 23304 18203 23333 18232
tri 23333 18203 23362 18232 nw
rect 29456 18214 29488 18270
rect 29544 18214 29568 18270
rect 29624 18214 29648 18270
rect 29704 18214 29728 18270
rect 29784 18214 29816 18270
tri 23260 18188 23275 18203 se
rect 23275 18188 23318 18203
tri 23318 18188 23333 18203 nw
tri 23246 18174 23260 18188 se
rect 23260 18174 23304 18188
tri 23304 18174 23318 18188 nw
rect 29456 18183 29816 18214
tri 23229 18157 23246 18174 se
rect 23246 18157 23287 18174
tri 23287 18157 23304 18174 nw
tri 23208 18136 23229 18157 se
rect 23229 18136 23266 18157
tri 23266 18136 23287 18157 nw
tri 23193 18121 23208 18136 se
rect 23208 18121 23251 18136
tri 23251 18121 23266 18136 nw
rect 29456 18127 29488 18183
rect 29544 18127 29568 18183
rect 29624 18127 29648 18183
rect 29704 18127 29728 18183
rect 29784 18127 29816 18183
tri 23188 18116 23193 18121 se
rect 23193 18116 23246 18121
tri 23246 18116 23251 18121 nw
tri 23141 18069 23188 18116 se
rect 23188 18069 23199 18116
tri 23199 18069 23246 18116 nw
rect 29456 18096 29816 18127
tri 23130 18058 23141 18069 se
rect 23141 18058 23188 18069
tri 23188 18058 23199 18069 nw
tri 23072 18000 23130 18058 se
tri 23130 18000 23188 18058 nw
rect 29456 18040 29488 18096
rect 29544 18040 29568 18096
rect 29624 18040 29648 18096
rect 29704 18040 29728 18096
rect 29784 18040 29816 18096
rect 29456 18009 29816 18040
tri 23032 17960 23072 18000 se
rect 20284 14889 20506 14963
rect 19429 14775 19911 14828
rect 19429 14719 19471 14775
rect 19527 14719 19551 14775
rect 19607 14719 19631 14775
rect 19687 14719 19711 14775
rect 19767 14719 19791 14775
rect 19847 14719 19911 14775
rect 19429 14694 19911 14719
rect 19429 14638 19471 14694
rect 19527 14638 19551 14694
rect 19607 14638 19631 14694
rect 19687 14638 19711 14694
rect 19767 14638 19791 14694
rect 19847 14638 19911 14694
rect 19429 14613 19911 14638
rect 19429 14557 19471 14613
rect 19527 14557 19551 14613
rect 19607 14557 19631 14613
rect 19687 14557 19711 14613
rect 19767 14557 19791 14613
rect 19847 14557 19911 14613
rect 19429 14532 19911 14557
rect 19429 14476 19471 14532
rect 19527 14476 19551 14532
rect 19607 14476 19631 14532
rect 19687 14476 19711 14532
rect 19767 14476 19791 14532
rect 19847 14476 19911 14532
rect 19429 14451 19911 14476
rect 19429 14395 19471 14451
rect 19527 14395 19551 14451
rect 19607 14395 19631 14451
rect 19687 14395 19711 14451
rect 19767 14395 19791 14451
rect 19847 14395 19911 14451
rect 19429 14370 19911 14395
rect 19429 14314 19471 14370
rect 19527 14314 19551 14370
rect 19607 14314 19631 14370
rect 19687 14314 19711 14370
rect 19767 14314 19791 14370
rect 19847 14314 19911 14370
rect 19429 14289 19911 14314
rect 19429 14233 19471 14289
rect 19527 14233 19551 14289
rect 19607 14233 19631 14289
rect 19687 14233 19711 14289
rect 19767 14233 19791 14289
rect 19847 14233 19911 14289
rect 19429 14208 19911 14233
rect 19429 14152 19471 14208
rect 19527 14152 19551 14208
rect 19607 14152 19631 14208
rect 19687 14152 19711 14208
rect 19767 14152 19791 14208
rect 19847 14152 19911 14208
rect 19429 14127 19911 14152
rect 19429 14071 19471 14127
rect 19527 14071 19551 14127
rect 19607 14071 19631 14127
rect 19687 14071 19711 14127
rect 19767 14071 19791 14127
rect 19847 14071 19911 14127
rect 19429 14046 19911 14071
rect 19429 13990 19471 14046
rect 19527 13990 19551 14046
rect 19607 13990 19631 14046
rect 19687 13990 19711 14046
rect 19767 13990 19791 14046
rect 19847 13990 19911 14046
rect 19429 13965 19911 13990
rect 19429 13909 19471 13965
rect 19527 13909 19551 13965
rect 19607 13909 19631 13965
rect 19687 13909 19711 13965
rect 19767 13909 19791 13965
rect 19847 13909 19911 13965
rect 19429 13884 19911 13909
rect 19429 13828 19471 13884
rect 19527 13828 19551 13884
rect 19607 13828 19631 13884
rect 19687 13828 19711 13884
rect 19767 13828 19791 13884
rect 19847 13828 19911 13884
rect 19429 13803 19911 13828
rect 19429 13747 19471 13803
rect 19527 13747 19551 13803
rect 19607 13747 19631 13803
rect 19687 13747 19711 13803
rect 19767 13747 19791 13803
rect 19847 13747 19911 13803
rect 19429 13722 19911 13747
rect 19429 13666 19471 13722
rect 19527 13666 19551 13722
rect 19607 13666 19631 13722
rect 19687 13666 19711 13722
rect 19767 13666 19791 13722
rect 19847 13666 19911 13722
rect 19429 13641 19911 13666
rect 19429 13585 19471 13641
rect 19527 13585 19551 13641
rect 19607 13585 19631 13641
rect 19687 13585 19711 13641
rect 19767 13585 19791 13641
rect 19847 13585 19911 13641
rect 19429 13560 19911 13585
rect 19429 13504 19471 13560
rect 19527 13504 19551 13560
rect 19607 13504 19631 13560
rect 19687 13504 19711 13560
rect 19767 13504 19791 13560
rect 19847 13504 19911 13560
rect 19429 13479 19911 13504
rect 19429 13423 19471 13479
rect 19527 13423 19551 13479
rect 19607 13423 19631 13479
rect 19687 13423 19711 13479
rect 19767 13423 19791 13479
rect 19847 13423 19911 13479
rect 19429 13398 19911 13423
rect 19429 13342 19471 13398
rect 19527 13342 19551 13398
rect 19607 13342 19631 13398
rect 19687 13342 19711 13398
rect 19767 13342 19791 13398
rect 19847 13342 19911 13398
rect 19429 13317 19911 13342
rect 19429 13261 19471 13317
rect 19527 13261 19551 13317
rect 19607 13261 19631 13317
rect 19687 13261 19711 13317
rect 19767 13261 19791 13317
rect 19847 13261 19911 13317
rect 19429 13236 19911 13261
rect 19429 13180 19471 13236
rect 19527 13180 19551 13236
rect 19607 13180 19631 13236
rect 19687 13180 19711 13236
rect 19767 13180 19791 13236
rect 19847 13180 19911 13236
rect 19429 13155 19911 13180
rect 19429 13099 19471 13155
rect 19527 13099 19551 13155
rect 19607 13099 19631 13155
rect 19687 13099 19711 13155
rect 19767 13099 19791 13155
rect 19847 13099 19911 13155
rect 19429 13074 19911 13099
rect 19429 13018 19471 13074
rect 19527 13018 19551 13074
rect 19607 13018 19631 13074
rect 19687 13018 19711 13074
rect 19767 13018 19791 13074
rect 19847 13018 19911 13074
rect 19429 12993 19911 13018
rect 19429 12937 19471 12993
rect 19527 12937 19551 12993
rect 19607 12937 19631 12993
rect 19687 12937 19711 12993
rect 19767 12937 19791 12993
rect 19847 12937 19911 12993
rect 19429 12912 19911 12937
rect 19429 12856 19471 12912
rect 19527 12856 19551 12912
rect 19607 12856 19631 12912
rect 19687 12856 19711 12912
rect 19767 12856 19791 12912
rect 19847 12856 19911 12912
rect 19429 12831 19911 12856
rect 19429 12775 19471 12831
rect 19527 12775 19551 12831
rect 19607 12775 19631 12831
rect 19687 12775 19711 12831
rect 19767 12775 19791 12831
rect 19847 12775 19911 12831
rect 19429 12750 19911 12775
rect 19429 12694 19471 12750
rect 19527 12694 19551 12750
rect 19607 12694 19631 12750
rect 19687 12694 19711 12750
rect 19767 12694 19791 12750
rect 19847 12694 19911 12750
rect 19429 12669 19911 12694
rect 19429 12613 19471 12669
rect 19527 12613 19551 12669
rect 19607 12613 19631 12669
rect 19687 12613 19711 12669
rect 19767 12613 19791 12669
rect 19847 12613 19911 12669
rect 19429 12588 19911 12613
rect 19429 12532 19471 12588
rect 19527 12532 19551 12588
rect 19607 12532 19631 12588
rect 19687 12532 19711 12588
rect 19767 12532 19791 12588
rect 19847 12532 19911 12588
rect 19429 12507 19911 12532
rect 19429 12451 19471 12507
rect 19527 12451 19551 12507
rect 19607 12451 19631 12507
rect 19687 12451 19711 12507
rect 19767 12451 19791 12507
rect 19847 12451 19911 12507
rect 19429 12426 19911 12451
rect 19429 12370 19471 12426
rect 19527 12370 19551 12426
rect 19607 12370 19631 12426
rect 19687 12370 19711 12426
rect 19767 12370 19791 12426
rect 19847 12370 19911 12426
rect 19429 12345 19911 12370
rect 19429 12289 19471 12345
rect 19527 12289 19551 12345
rect 19607 12289 19631 12345
rect 19687 12289 19711 12345
rect 19767 12289 19791 12345
rect 19847 12289 19911 12345
rect 19429 12264 19911 12289
rect 19429 12208 19471 12264
rect 19527 12208 19551 12264
rect 19607 12208 19631 12264
rect 19687 12208 19711 12264
rect 19767 12208 19791 12264
rect 19847 12208 19911 12264
rect 19429 12183 19911 12208
rect 19429 12127 19471 12183
rect 19527 12127 19551 12183
rect 19607 12127 19631 12183
rect 19687 12127 19711 12183
rect 19767 12127 19791 12183
rect 19847 12127 19911 12183
rect 19429 12102 19911 12127
rect 19429 12046 19471 12102
rect 19527 12046 19551 12102
rect 19607 12046 19631 12102
rect 19687 12046 19711 12102
rect 19767 12046 19791 12102
rect 19847 12046 19911 12102
rect 19429 12021 19911 12046
rect 19429 11965 19471 12021
rect 19527 11965 19551 12021
rect 19607 11965 19631 12021
rect 19687 11965 19711 12021
rect 19767 11965 19791 12021
rect 19847 11965 19911 12021
rect 19429 11939 19911 11965
rect 19429 11883 19471 11939
rect 19527 11883 19551 11939
rect 19607 11883 19631 11939
rect 19687 11883 19711 11939
rect 19767 11883 19791 11939
rect 19847 11883 19911 11939
rect 19429 11857 19911 11883
rect 19429 11801 19471 11857
rect 19527 11801 19551 11857
rect 19607 11801 19631 11857
rect 19687 11801 19711 11857
rect 19767 11801 19791 11857
rect 19847 11801 19911 11857
rect 19429 11775 19911 11801
rect 19429 11719 19471 11775
rect 19527 11719 19551 11775
rect 19607 11719 19631 11775
rect 19687 11719 19711 11775
rect 19767 11719 19791 11775
rect 19847 11719 19911 11775
rect 19429 11693 19911 11719
rect 19429 11637 19471 11693
rect 19527 11637 19551 11693
rect 19607 11637 19631 11693
rect 19687 11637 19711 11693
rect 19767 11637 19791 11693
rect 19847 11637 19911 11693
rect 19429 11611 19911 11637
rect 19429 11555 19471 11611
rect 19527 11555 19551 11611
rect 19607 11555 19631 11611
rect 19687 11555 19711 11611
rect 19767 11555 19791 11611
rect 19847 11555 19911 11611
rect 19429 11529 19911 11555
rect 19429 11473 19471 11529
rect 19527 11473 19551 11529
rect 19607 11473 19631 11529
rect 19687 11473 19711 11529
rect 19767 11473 19791 11529
rect 19847 11473 19911 11529
rect 19429 11447 19911 11473
rect 19429 11391 19471 11447
rect 19527 11391 19551 11447
rect 19607 11391 19631 11447
rect 19687 11391 19711 11447
rect 19767 11391 19791 11447
rect 19847 11391 19911 11447
rect 19429 11365 19911 11391
rect 19429 11336 19551 11365
tri 19551 11340 19576 11365 nw
tri 19634 11340 19659 11365 ne
rect 19429 11280 19462 11336
rect 19518 11280 19551 11336
rect 19429 11256 19551 11280
rect 19429 11200 19462 11256
rect 19518 11200 19551 11256
rect 19429 11176 19551 11200
rect 19429 11120 19462 11176
rect 19518 11120 19551 11176
rect 19429 11096 19551 11120
rect 19429 11040 19462 11096
rect 19518 11040 19551 11096
rect 19429 11015 19551 11040
rect 19429 10959 19462 11015
rect 19518 10959 19551 11015
rect 19429 10934 19551 10959
rect 19429 10878 19462 10934
rect 19518 10878 19551 10934
rect 19429 10853 19551 10878
rect 19429 10797 19462 10853
rect 19518 10797 19551 10853
rect 19429 10772 19551 10797
rect 19429 10716 19462 10772
rect 19518 10716 19551 10772
rect 19429 10691 19551 10716
rect 19429 10635 19462 10691
rect 19518 10635 19551 10691
rect 19429 10610 19551 10635
rect 19429 10554 19462 10610
rect 19518 10554 19551 10610
rect 19429 10529 19551 10554
rect 19429 10473 19462 10529
rect 19518 10473 19551 10529
rect 19429 10448 19551 10473
rect 19429 10392 19462 10448
rect 19518 10392 19551 10448
rect 19429 10367 19551 10392
rect 19429 10311 19462 10367
rect 19518 10311 19551 10367
rect 19429 10286 19551 10311
rect 19429 10230 19462 10286
rect 19518 10230 19551 10286
rect 19429 10205 19551 10230
rect 19429 10149 19462 10205
rect 19518 10149 19551 10205
rect 19429 10124 19551 10149
rect 19429 10068 19462 10124
rect 19518 10068 19551 10124
rect 19429 10043 19551 10068
rect 19429 9987 19462 10043
rect 19518 9987 19551 10043
rect 19429 9962 19551 9987
rect 19429 9906 19462 9962
rect 19518 9906 19551 9962
rect 19429 9881 19551 9906
rect 19429 9825 19462 9881
rect 19518 9825 19551 9881
rect 19429 9800 19551 9825
rect 19429 9744 19462 9800
rect 19518 9744 19551 9800
rect 19429 9719 19551 9744
rect 19429 9663 19462 9719
rect 19518 9663 19551 9719
rect 19429 9638 19551 9663
rect 19429 9582 19462 9638
rect 19518 9582 19551 9638
rect 19429 9557 19551 9582
rect 19429 9501 19462 9557
rect 19518 9501 19551 9557
rect 19429 9476 19551 9501
rect 19429 9420 19462 9476
rect 19518 9420 19551 9476
rect 19429 9395 19551 9420
rect 19429 9339 19462 9395
rect 19518 9339 19551 9395
rect 19429 9314 19551 9339
rect 19429 9258 19462 9314
rect 19518 9258 19551 9314
rect 19429 9233 19551 9258
rect 19429 9177 19462 9233
rect 19518 9177 19551 9233
rect 19429 9152 19551 9177
rect 19429 9096 19462 9152
rect 19518 9096 19551 9152
rect 19429 9071 19551 9096
rect 19429 9015 19462 9071
rect 19518 9015 19551 9071
rect 19429 8990 19551 9015
rect 19429 8934 19462 8990
rect 19518 8934 19551 8990
rect 19429 8909 19551 8934
rect 19429 8853 19462 8909
rect 19518 8853 19551 8909
rect 19429 8828 19551 8853
rect 19429 8772 19462 8828
rect 19518 8772 19551 8828
rect 19429 8732 19551 8772
rect 19659 11333 19911 11365
rect 19659 11277 19720 11333
rect 19776 11277 19800 11333
rect 19856 11277 19911 11333
rect 19659 11252 19911 11277
rect 19659 11196 19720 11252
rect 19776 11196 19800 11252
rect 19856 11196 19911 11252
rect 19659 11171 19911 11196
rect 19659 11115 19720 11171
rect 19776 11115 19800 11171
rect 19856 11115 19911 11171
rect 19659 11090 19911 11115
rect 19659 11034 19720 11090
rect 19776 11034 19800 11090
rect 19856 11034 19911 11090
rect 19659 11009 19911 11034
rect 19659 10953 19720 11009
rect 19776 10953 19800 11009
rect 19856 10953 19911 11009
rect 19659 10928 19911 10953
rect 19659 10872 19720 10928
rect 19776 10872 19800 10928
rect 19856 10872 19911 10928
rect 19659 10847 19911 10872
rect 19659 10791 19720 10847
rect 19776 10791 19800 10847
rect 19856 10791 19911 10847
rect 19659 10766 19911 10791
rect 19659 10710 19720 10766
rect 19776 10710 19800 10766
rect 19856 10710 19911 10766
rect 19659 10685 19911 10710
rect 19659 10629 19720 10685
rect 19776 10629 19800 10685
rect 19856 10629 19911 10685
rect 19659 10604 19911 10629
rect 19659 10548 19720 10604
rect 19776 10548 19800 10604
rect 19856 10548 19911 10604
rect 19659 10523 19911 10548
rect 19659 10467 19720 10523
rect 19776 10467 19800 10523
rect 19856 10467 19911 10523
rect 19659 10442 19911 10467
rect 19659 10386 19720 10442
rect 19776 10386 19800 10442
rect 19856 10386 19911 10442
rect 19659 10361 19911 10386
rect 19659 10305 19720 10361
rect 19776 10305 19800 10361
rect 19856 10305 19911 10361
rect 19659 10280 19911 10305
rect 19659 10224 19720 10280
rect 19776 10224 19800 10280
rect 19856 10224 19911 10280
rect 19659 10199 19911 10224
rect 19659 10143 19720 10199
rect 19776 10143 19800 10199
rect 19856 10143 19911 10199
rect 19659 10118 19911 10143
rect 19659 10062 19720 10118
rect 19776 10062 19800 10118
rect 19856 10062 19911 10118
rect 19659 10037 19911 10062
rect 19659 9981 19720 10037
rect 19776 9981 19800 10037
rect 19856 9981 19911 10037
rect 19659 9956 19911 9981
rect 19659 9900 19720 9956
rect 19776 9900 19800 9956
rect 19856 9900 19911 9956
rect 19659 9875 19911 9900
rect 19659 9819 19720 9875
rect 19776 9819 19800 9875
rect 19856 9819 19911 9875
rect 19659 9794 19911 9819
rect 19659 9738 19720 9794
rect 19776 9738 19800 9794
rect 19856 9738 19911 9794
rect 19659 9713 19911 9738
rect 19659 9657 19720 9713
rect 19776 9657 19800 9713
rect 19856 9657 19911 9713
rect 19659 9631 19911 9657
rect 19659 9575 19720 9631
rect 19776 9575 19800 9631
rect 19856 9575 19911 9631
rect 19659 9549 19911 9575
rect 19659 9493 19720 9549
rect 19776 9493 19800 9549
rect 19856 9493 19911 9549
rect 19659 9467 19911 9493
rect 19659 9411 19720 9467
rect 19776 9411 19800 9467
rect 19856 9411 19911 9467
rect 19659 9385 19911 9411
rect 19659 9329 19720 9385
rect 19776 9329 19800 9385
rect 19856 9329 19911 9385
rect 19659 9303 19911 9329
rect 19659 9247 19720 9303
rect 19776 9247 19800 9303
rect 19856 9247 19911 9303
rect 19659 9221 19911 9247
rect 19659 9165 19720 9221
rect 19776 9165 19800 9221
rect 19856 9165 19911 9221
rect 19659 9139 19911 9165
rect 19659 9083 19720 9139
rect 19776 9083 19800 9139
rect 19856 9083 19911 9139
rect 19659 9057 19911 9083
rect 19659 9001 19720 9057
rect 19776 9001 19800 9057
rect 19856 9001 19911 9057
rect 19659 8975 19911 9001
rect 19659 8919 19720 8975
rect 19776 8919 19800 8975
rect 19856 8919 19911 8975
rect 19659 8893 19911 8919
rect 19659 8837 19720 8893
rect 19776 8837 19800 8893
rect 19856 8837 19911 8893
rect 19659 8811 19911 8837
tri 19551 8732 19576 8757 sw
tri 19634 8732 19659 8757 se
rect 19659 8755 19720 8811
rect 19776 8755 19800 8811
rect 19856 8755 19911 8811
rect 19659 8732 19911 8755
rect 19429 8669 19911 8732
rect 19429 8613 19482 8669
rect 19538 8613 19562 8669
rect 19618 8613 19642 8669
rect 19698 8613 19722 8669
rect 19778 8613 19802 8669
rect 19858 8613 19911 8669
rect 19429 8584 19911 8613
rect 19429 8528 19482 8584
rect 19538 8528 19562 8584
rect 19618 8528 19642 8584
rect 19698 8528 19722 8584
rect 19778 8528 19802 8584
rect 19858 8528 19911 8584
rect 19429 8498 19911 8528
rect 19429 8442 19482 8498
rect 19538 8442 19562 8498
rect 19618 8442 19642 8498
rect 19698 8442 19722 8498
rect 19778 8442 19802 8498
rect 19858 8442 19911 8498
rect 19429 8412 19911 8442
rect 19429 8356 19482 8412
rect 19538 8356 19562 8412
rect 19618 8356 19642 8412
rect 19698 8356 19722 8412
rect 19778 8356 19802 8412
rect 19858 8356 19911 8412
rect 19429 8326 19911 8356
rect 19429 8270 19482 8326
rect 19538 8270 19562 8326
rect 19618 8270 19642 8326
rect 19698 8270 19722 8326
rect 19778 8270 19802 8326
rect 19858 8270 19911 8326
rect 19429 8240 19911 8270
rect 19429 8184 19482 8240
rect 19538 8184 19562 8240
rect 19618 8184 19642 8240
rect 19698 8184 19722 8240
rect 19778 8184 19802 8240
rect 19858 8184 19911 8240
rect 19429 8154 19911 8184
rect 19429 8098 19482 8154
rect 19538 8098 19562 8154
rect 19618 8098 19642 8154
rect 19698 8098 19722 8154
rect 19778 8098 19802 8154
rect 19858 8098 19911 8154
rect 19429 8083 19911 8098
rect 19429 8031 19435 8083
rect 19487 8068 19503 8083
rect 19555 8068 19571 8083
rect 19555 8031 19562 8068
rect 19623 8031 19639 8083
rect 19691 8068 19707 8083
rect 19759 8068 19775 8083
rect 19827 8068 19842 8083
rect 19698 8031 19707 8068
rect 19894 8031 19911 8083
rect 19429 8019 19482 8031
rect 19538 8019 19562 8031
rect 19618 8019 19642 8031
rect 19698 8019 19722 8031
rect 19778 8019 19802 8031
rect 19858 8019 19911 8031
rect 19429 7967 19435 8019
rect 19555 8012 19562 8019
rect 19487 7982 19503 8012
rect 19555 7982 19571 8012
rect 19555 7967 19562 7982
rect 19623 7967 19639 8019
rect 19698 8012 19707 8019
rect 19691 7982 19707 8012
rect 19759 7982 19775 8012
rect 19827 7982 19842 8012
rect 19698 7967 19707 7982
rect 19894 7967 19911 8019
rect 19429 7955 19482 7967
rect 19538 7955 19562 7967
rect 19618 7955 19642 7967
rect 19698 7955 19722 7967
rect 19778 7955 19802 7967
rect 19858 7955 19911 7967
rect 19429 7903 19435 7955
rect 19555 7926 19562 7955
rect 19487 7903 19503 7926
rect 19555 7903 19571 7926
rect 19623 7903 19639 7955
rect 19698 7926 19707 7955
rect 19691 7903 19707 7926
rect 19759 7903 19775 7926
rect 19827 7903 19842 7926
rect 19894 7903 19911 7955
rect -1954 5550 -1418 5559
rect -1954 5069 -1418 5094
rect -1898 5013 -1874 5069
rect -1818 5013 -1794 5069
rect -1738 5013 -1714 5069
rect -1658 5013 -1634 5069
rect -1578 5013 -1554 5069
rect -1498 5013 -1474 5069
rect -1954 4988 -1418 5013
rect -1898 4932 -1874 4988
rect -1818 4932 -1794 4988
rect -1738 4932 -1714 4988
rect -1658 4932 -1634 4988
rect -1578 4932 -1554 4988
rect -1498 4932 -1474 4988
rect -1954 4907 -1418 4932
rect -1898 4851 -1874 4907
rect -1818 4851 -1794 4907
rect -1738 4851 -1714 4907
rect -1658 4851 -1634 4907
rect -1578 4851 -1554 4907
rect -1498 4851 -1474 4907
rect -1954 4826 -1418 4851
rect -1898 4770 -1874 4826
rect -1818 4770 -1794 4826
rect -1738 4770 -1714 4826
rect -1658 4770 -1634 4826
rect -1578 4770 -1554 4826
rect -1498 4770 -1474 4826
rect -1954 4745 -1418 4770
rect -1898 4689 -1874 4745
rect -1818 4689 -1794 4745
rect -1738 4689 -1714 4745
rect -1658 4689 -1634 4745
rect -1578 4689 -1554 4745
rect -1498 4689 -1474 4745
rect -1954 4664 -1418 4689
rect -1898 4608 -1874 4664
rect -1818 4608 -1794 4664
rect -1738 4608 -1714 4664
rect -1658 4608 -1634 4664
rect -1578 4608 -1554 4664
rect -1498 4608 -1474 4664
rect -1954 4583 -1418 4608
rect -3209 4560 -3157 4566
rect -3209 4496 -3157 4508
rect -3209 4438 -3157 4444
rect -2889 4552 -2837 4558
rect -2889 4488 -2837 4500
rect -2889 4430 -2837 4436
rect -2809 4552 -2757 4558
rect -2809 4488 -2757 4500
rect -2809 4430 -2757 4436
rect -2729 4539 -2677 4545
rect -2729 4475 -2677 4487
rect -2729 4417 -2677 4423
rect -2569 4539 -2517 4545
rect -1898 4527 -1874 4583
rect -1818 4527 -1794 4583
rect -1738 4527 -1714 4583
rect -1658 4527 -1634 4583
rect -1578 4527 -1554 4583
rect -1498 4527 -1474 4583
rect -1954 4502 -1418 4527
rect -2569 4475 -2517 4487
rect -2409 4464 -2357 4498
rect -1898 4446 -1874 4502
rect -1818 4446 -1794 4502
rect -1738 4446 -1714 4502
rect -1658 4446 -1634 4502
rect -1578 4446 -1554 4502
rect -1498 4446 -1474 4502
rect -1954 4437 -1418 4446
rect -163 5550 373 5559
rect -163 5069 373 5094
rect -107 5013 -83 5069
rect -27 5013 -3 5069
rect 53 5013 77 5069
rect 133 5013 157 5069
rect 213 5013 237 5069
rect 293 5013 317 5069
rect -163 4988 373 5013
rect -107 4932 -83 4988
rect -27 4932 -3 4988
rect 53 4932 77 4988
rect 133 4932 157 4988
rect 213 4932 237 4988
rect 293 4932 317 4988
rect -163 4907 373 4932
rect -107 4851 -83 4907
rect -27 4851 -3 4907
rect 53 4851 77 4907
rect 133 4851 157 4907
rect 213 4851 237 4907
rect 293 4851 317 4907
rect -163 4826 373 4851
rect -107 4770 -83 4826
rect -27 4770 -3 4826
rect 53 4770 77 4826
rect 133 4770 157 4826
rect 213 4770 237 4826
rect 293 4770 317 4826
rect -163 4745 373 4770
rect -107 4689 -83 4745
rect -27 4689 -3 4745
rect 53 4689 77 4745
rect 133 4689 157 4745
rect 213 4689 237 4745
rect 293 4689 317 4745
rect -163 4664 373 4689
rect -107 4608 -83 4664
rect -27 4608 -3 4664
rect 53 4608 77 4664
rect 133 4608 157 4664
rect 213 4608 237 4664
rect 293 4608 317 4664
rect -163 4583 373 4608
rect -107 4527 -83 4583
rect -27 4527 -3 4583
rect 53 4527 77 4583
rect 133 4527 157 4583
rect 213 4527 237 4583
rect 293 4527 317 4583
rect -163 4502 373 4527
rect -107 4446 -83 4502
rect -27 4446 -3 4502
rect 53 4446 77 4502
rect 133 4446 157 4502
rect 213 4446 237 4502
rect 293 4446 317 4502
rect -163 4437 373 4446
rect 1657 5550 2193 5559
rect 1657 5069 2193 5094
rect 1713 5013 1737 5069
rect 1793 5013 1817 5069
rect 1873 5013 1897 5069
rect 1953 5013 1977 5069
rect 2033 5013 2057 5069
rect 2113 5013 2137 5069
rect 1657 4988 2193 5013
rect 1713 4932 1737 4988
rect 1793 4932 1817 4988
rect 1873 4932 1897 4988
rect 1953 4932 1977 4988
rect 2033 4932 2057 4988
rect 2113 4932 2137 4988
rect 1657 4907 2193 4932
rect 1713 4851 1737 4907
rect 1793 4851 1817 4907
rect 1873 4851 1897 4907
rect 1953 4851 1977 4907
rect 2033 4851 2057 4907
rect 2113 4851 2137 4907
rect 1657 4826 2193 4851
rect 1713 4770 1737 4826
rect 1793 4770 1817 4826
rect 1873 4770 1897 4826
rect 1953 4770 1977 4826
rect 2033 4770 2057 4826
rect 2113 4770 2137 4826
rect 1657 4745 2193 4770
rect 1713 4689 1737 4745
rect 1793 4689 1817 4745
rect 1873 4689 1897 4745
rect 1953 4689 1977 4745
rect 2033 4689 2057 4745
rect 2113 4689 2137 4745
rect 1657 4664 2193 4689
rect 1713 4608 1737 4664
rect 1793 4608 1817 4664
rect 1873 4608 1897 4664
rect 1953 4608 1977 4664
rect 2033 4608 2057 4664
rect 2113 4608 2137 4664
rect 1657 4583 2193 4608
rect 1713 4527 1737 4583
rect 1793 4527 1817 4583
rect 1873 4527 1897 4583
rect 1953 4527 1977 4583
rect 2033 4527 2057 4583
rect 2113 4527 2137 4583
rect 3458 5550 3994 5559
rect 3458 5069 3994 5094
rect 3514 5013 3538 5069
rect 3594 5013 3618 5069
rect 3674 5013 3698 5069
rect 3754 5013 3778 5069
rect 3834 5013 3858 5069
rect 3914 5013 3938 5069
rect 3458 4988 3994 5013
rect 3514 4932 3538 4988
rect 3594 4932 3618 4988
rect 3674 4932 3698 4988
rect 3754 4932 3778 4988
rect 3834 4932 3858 4988
rect 3914 4932 3938 4988
rect 3458 4907 3994 4932
rect 3514 4851 3538 4907
rect 3594 4851 3618 4907
rect 3674 4851 3698 4907
rect 3754 4851 3778 4907
rect 3834 4851 3858 4907
rect 3914 4851 3938 4907
rect 3458 4826 3994 4851
rect 3514 4770 3538 4826
rect 3594 4770 3618 4826
rect 3674 4770 3698 4826
rect 3754 4770 3778 4826
rect 3834 4770 3858 4826
rect 3914 4770 3938 4826
rect 3458 4745 3994 4770
rect 3514 4689 3538 4745
rect 3594 4689 3618 4745
rect 3674 4689 3698 4745
rect 3754 4689 3778 4745
rect 3834 4689 3858 4745
rect 3914 4689 3938 4745
rect 3458 4664 3994 4689
rect 3514 4608 3538 4664
rect 3594 4608 3618 4664
rect 3674 4608 3698 4664
rect 3754 4608 3778 4664
rect 3834 4608 3858 4664
rect 3914 4608 3938 4664
rect 3458 4583 3994 4608
rect 1657 4502 2193 4527
rect 1713 4446 1737 4502
rect 1793 4446 1817 4502
rect 1873 4446 1897 4502
rect 1953 4446 1977 4502
rect 2033 4446 2057 4502
rect 2113 4446 2137 4502
rect 2409 4464 2591 4538
rect 3514 4527 3538 4583
rect 3594 4527 3618 4583
rect 3674 4527 3698 4583
rect 3754 4527 3778 4583
rect 3834 4527 3858 4583
rect 3914 4527 3938 4583
rect 5266 5550 5802 5559
rect 5266 5069 5802 5094
rect 5322 5013 5346 5069
rect 5402 5013 5426 5069
rect 5482 5013 5506 5069
rect 5562 5013 5586 5069
rect 5642 5013 5666 5069
rect 5722 5013 5746 5069
rect 5266 4988 5802 5013
rect 5322 4932 5346 4988
rect 5402 4932 5426 4988
rect 5482 4932 5506 4988
rect 5562 4932 5586 4988
rect 5642 4932 5666 4988
rect 5722 4932 5746 4988
rect 5266 4907 5802 4932
rect 5322 4851 5346 4907
rect 5402 4851 5426 4907
rect 5482 4851 5506 4907
rect 5562 4851 5586 4907
rect 5642 4851 5666 4907
rect 5722 4851 5746 4907
rect 5266 4826 5802 4851
rect 5322 4770 5346 4826
rect 5402 4770 5426 4826
rect 5482 4770 5506 4826
rect 5562 4770 5586 4826
rect 5642 4770 5666 4826
rect 5722 4770 5746 4826
rect 5266 4745 5802 4770
rect 5322 4689 5346 4745
rect 5402 4689 5426 4745
rect 5482 4689 5506 4745
rect 5562 4689 5586 4745
rect 5642 4689 5666 4745
rect 5722 4689 5746 4745
rect 7061 5550 7597 5559
rect 7117 5494 7141 5550
rect 7197 5494 7221 5550
rect 7277 5494 7301 5550
rect 7357 5494 7381 5550
rect 7437 5494 7461 5550
rect 7517 5494 7541 5550
rect 10660 5558 11196 5567
rect 7061 5467 7597 5494
rect 7117 5411 7141 5467
rect 7197 5411 7221 5467
rect 7277 5411 7301 5467
rect 7357 5411 7381 5467
rect 7437 5411 7461 5467
rect 7517 5411 7541 5467
rect 7061 5384 7597 5411
rect 7117 5328 7141 5384
rect 7197 5328 7221 5384
rect 7277 5328 7301 5384
rect 7357 5328 7381 5384
rect 7437 5328 7461 5384
rect 7517 5328 7541 5384
rect 7061 5301 7597 5328
rect 7117 5245 7141 5301
rect 7197 5245 7221 5301
rect 7277 5245 7301 5301
rect 7357 5245 7381 5301
rect 7437 5245 7461 5301
rect 7517 5245 7541 5301
rect 7061 5218 7597 5245
rect 7117 5162 7141 5218
rect 7197 5162 7221 5218
rect 7277 5162 7301 5218
rect 7357 5162 7381 5218
rect 7437 5162 7461 5218
rect 7517 5162 7541 5218
rect 7061 5134 7597 5162
rect 7117 5078 7141 5134
rect 7197 5078 7221 5134
rect 7277 5078 7301 5134
rect 7357 5078 7381 5134
rect 7437 5078 7461 5134
rect 7517 5078 7541 5134
rect 7061 5050 7597 5078
rect 7117 4994 7141 5050
rect 7197 4994 7221 5050
rect 7277 4994 7301 5050
rect 7357 4994 7381 5050
rect 7437 4994 7461 5050
rect 7517 4994 7541 5050
rect 7061 4966 7597 4994
rect 7117 4910 7141 4966
rect 7197 4910 7221 4966
rect 7277 4910 7301 4966
rect 7357 4910 7381 4966
rect 7437 4910 7461 4966
rect 7517 4910 7541 4966
rect 7061 4882 7597 4910
rect 7117 4826 7141 4882
rect 7197 4826 7221 4882
rect 7277 4826 7301 4882
rect 7357 4826 7381 4882
rect 7437 4826 7461 4882
rect 7517 4826 7541 4882
rect 7061 4798 7597 4826
rect 7117 4742 7141 4798
rect 7197 4742 7221 4798
rect 7277 4742 7301 4798
rect 7357 4742 7381 4798
rect 7437 4742 7461 4798
rect 7517 4742 7541 4798
rect 7061 4733 7597 4742
rect 8868 5530 9412 5539
rect 8868 5474 8872 5530
rect 8928 5474 8952 5530
rect 9008 5474 9032 5530
rect 9088 5474 9112 5530
rect 9168 5474 9192 5530
rect 9248 5474 9272 5530
rect 9328 5474 9352 5530
rect 9408 5474 9412 5530
rect 8868 5449 9412 5474
rect 8868 5393 8872 5449
rect 8928 5393 8952 5449
rect 9008 5393 9032 5449
rect 9088 5393 9112 5449
rect 9168 5393 9192 5449
rect 9248 5393 9272 5449
rect 9328 5393 9352 5449
rect 9408 5393 9412 5449
rect 8868 5368 9412 5393
rect 8868 5312 8872 5368
rect 8928 5312 8952 5368
rect 9008 5312 9032 5368
rect 9088 5312 9112 5368
rect 9168 5312 9192 5368
rect 9248 5312 9272 5368
rect 9328 5312 9352 5368
rect 9408 5312 9412 5368
rect 8868 5287 9412 5312
rect 8868 5231 8872 5287
rect 8928 5231 8952 5287
rect 9008 5231 9032 5287
rect 9088 5231 9112 5287
rect 9168 5231 9192 5287
rect 9248 5231 9272 5287
rect 9328 5231 9352 5287
rect 9408 5231 9412 5287
rect 8868 5206 9412 5231
rect 8868 5150 8872 5206
rect 8928 5150 8952 5206
rect 9008 5150 9032 5206
rect 9088 5150 9112 5206
rect 9168 5150 9192 5206
rect 9248 5150 9272 5206
rect 9328 5150 9352 5206
rect 9408 5150 9412 5206
rect 8868 5125 9412 5150
rect 8868 5069 8872 5125
rect 8928 5069 8952 5125
rect 9008 5069 9032 5125
rect 9088 5069 9112 5125
rect 9168 5069 9192 5125
rect 9248 5069 9272 5125
rect 9328 5069 9352 5125
rect 9408 5069 9412 5125
rect 8868 5044 9412 5069
rect 8868 4988 8872 5044
rect 8928 4988 8952 5044
rect 9008 4988 9032 5044
rect 9088 4988 9112 5044
rect 9168 4988 9192 5044
rect 9248 4988 9272 5044
rect 9328 4988 9352 5044
rect 9408 4988 9412 5044
rect 8868 4963 9412 4988
rect 8868 4907 8872 4963
rect 8928 4907 8952 4963
rect 9008 4907 9032 4963
rect 9088 4907 9112 4963
rect 9168 4907 9192 4963
rect 9248 4907 9272 4963
rect 9328 4907 9352 4963
rect 9408 4907 9412 4963
rect 8868 4881 9412 4907
rect 8868 4825 8872 4881
rect 8928 4825 8952 4881
rect 9008 4825 9032 4881
rect 9088 4825 9112 4881
rect 9168 4825 9192 4881
rect 9248 4825 9272 4881
rect 9328 4825 9352 4881
rect 9408 4825 9412 4881
rect 8868 4799 9412 4825
rect 8868 4743 8872 4799
rect 8928 4743 8952 4799
rect 9008 4743 9032 4799
rect 9088 4743 9112 4799
rect 9168 4743 9192 4799
rect 9248 4743 9272 4799
rect 9328 4743 9352 4799
rect 9408 4743 9412 4799
rect 5266 4664 5802 4689
rect 5322 4608 5346 4664
rect 5402 4608 5426 4664
rect 5482 4608 5506 4664
rect 5562 4608 5586 4664
rect 5642 4608 5666 4664
rect 5722 4608 5746 4664
rect 8868 4717 9412 4743
rect 8868 4661 8872 4717
rect 8928 4661 8952 4717
rect 9008 4661 9032 4717
rect 9088 4661 9112 4717
rect 9168 4661 9192 4717
rect 9248 4661 9272 4717
rect 9328 4661 9352 4717
rect 9408 4661 9412 4717
rect 8868 4635 9412 4661
tri 8723 4624 8725 4626 nw
rect 5266 4583 5802 4608
rect 3458 4504 3994 4527
rect 3427 4502 4027 4504
rect 1657 4437 2193 4446
tri 2295 4445 2314 4464 se
rect 2314 4445 3299 4464
tri 3299 4445 3318 4464 nw
rect 3427 4446 3458 4502
rect 3514 4446 3538 4502
rect 3594 4446 3618 4502
rect 3674 4446 3698 4502
rect 3754 4446 3778 4502
rect 3834 4446 3858 4502
rect 3914 4446 3938 4502
rect 3994 4446 4027 4502
rect 4124 4497 4530 4503
rect 4124 4464 4126 4497
tri 2287 4437 2295 4445 se
rect 2295 4437 3286 4445
tri 2282 4432 2287 4437 se
rect 2287 4432 3286 4437
tri 3286 4432 3299 4445 nw
rect -2569 4417 -2517 4423
tri 2267 4417 2282 4432 se
rect 2282 4417 3234 4432
tri 2230 4380 2267 4417 se
rect 2267 4380 3234 4417
tri 3234 4380 3286 4432 nw
tri 2217 4367 2230 4380 se
rect 2230 4367 3221 4380
tri 3221 4367 3234 4380 nw
tri 2215 4365 2217 4367 se
rect 2217 4365 3219 4367
tri 3219 4365 3221 4367 nw
rect 2215 4315 3169 4365
tri 3169 4315 3219 4365 nw
rect 2215 4302 3156 4315
tri 3156 4302 3169 4315 nw
rect 2215 4294 3148 4302
tri 3148 4294 3156 4302 nw
rect 2215 4293 3147 4294
tri 3147 4293 3148 4294 nw
tri 3426 4293 3427 4294 se
rect 3427 4293 4027 4446
rect 865 4284 1095 4293
rect 921 4228 945 4284
rect 1001 4228 1025 4284
rect 1081 4228 1095 4284
rect 865 4200 1095 4228
rect 921 4144 945 4200
rect 1001 4144 1025 4200
rect 1081 4144 1095 4200
rect 865 4116 1095 4144
rect 921 4060 945 4116
rect 1001 4060 1025 4116
rect 1081 4060 1095 4116
rect -14 3991 -8 4043
rect 44 3991 56 4043
rect 108 3991 114 4043
rect 865 4031 1095 4060
rect 1464 4067 1654 4096
tri 1654 4067 1683 4096 sw
rect 1464 4044 1627 4067
rect 921 3975 945 4031
rect 1001 3975 1025 4031
rect 1081 3975 1095 4031
tri 1592 4015 1621 4044 ne
rect 1621 4015 1627 4044
rect 1679 4015 1708 4067
rect 1760 4015 1766 4067
rect 865 3946 1095 3975
rect 921 3890 945 3946
rect 1001 3890 1025 3946
rect 1081 3890 1095 3946
rect 865 3861 1095 3890
rect 921 3805 945 3861
rect 1001 3805 1025 3861
rect 1081 3805 1095 3861
rect 865 3776 1095 3805
rect 921 3720 945 3776
rect 1001 3720 1025 3776
rect 1081 3720 1095 3776
tri 841 3687 865 3711 se
rect 865 3687 1095 3720
rect -3049 3419 -2997 3425
rect -3049 3355 -2997 3367
rect -209 3373 -203 3425
rect -151 3373 -139 3425
rect -87 3373 -81 3425
tri -209 3358 -194 3373 ne
rect -194 3358 -96 3373
tri -96 3358 -81 3373 nw
rect 39 3410 665 3416
tri 665 3410 671 3416 sw
rect 91 3390 671 3410
tri 671 3390 691 3410 sw
rect 91 3358 691 3390
tri -194 3346 -182 3358 ne
rect -182 3346 -108 3358
tri -108 3346 -96 3358 nw
rect 39 3346 691 3358
tri -182 3335 -171 3346 ne
rect -3049 3297 -2997 3303
tri -209 867 -171 905 se
rect -171 867 -119 3346
tri -119 3335 -108 3346 nw
rect 91 3294 691 3346
rect 39 3288 691 3294
tri 39 3236 91 3288 ne
rect 91 3183 691 3288
rect 91 1447 167 3183
rect 623 1447 691 3183
rect 91 1422 691 1447
rect 91 1366 167 1422
rect 223 1366 247 1422
rect 303 1366 327 1422
rect 383 1366 407 1422
rect 463 1366 487 1422
rect 543 1366 567 1422
rect 623 1366 691 1422
rect 91 1068 691 1366
tri 747 2545 841 2639 se
rect 841 2545 1095 3687
rect 747 2514 1095 2545
rect 747 2473 1054 2514
tri 1054 2473 1095 2514 nw
tri 1551 2473 1879 2801 se
rect 1879 2473 2159 4255
rect 747 2444 1025 2473
tri 1025 2444 1054 2473 nw
tri 1317 2444 1346 2473 se
rect 1346 2444 2159 2473
rect 2215 4250 3104 4293
tri 3104 4250 3147 4293 nw
tri 3383 4250 3426 4293 se
rect 3426 4250 4027 4293
rect 2215 4237 3091 4250
tri 3091 4237 3104 4250 nw
tri 3370 4237 3383 4250 se
rect 3383 4237 4027 4250
rect 2215 4185 3039 4237
tri 3039 4185 3091 4237 nw
tri 3318 4185 3370 4237 se
rect 3370 4185 4027 4237
rect 2215 4171 3025 4185
tri 3025 4171 3039 4185 nw
tri 3304 4171 3318 4185 se
rect 3318 4171 4027 4185
rect 2215 4156 3010 4171
tri 3010 4156 3025 4171 nw
tri 3289 4156 3304 4171 se
rect 3304 4156 4027 4171
rect 2215 4143 2997 4156
tri 2997 4143 3010 4156 nw
tri 3276 4143 3289 4156 se
rect 3289 4143 4027 4156
rect 2215 4119 2973 4143
tri 2973 4119 2997 4143 nw
tri 3252 4119 3276 4143 se
rect 3276 4119 4027 4143
rect 2215 4105 2959 4119
tri 2959 4105 2973 4119 nw
tri 3238 4105 3252 4119 se
rect 3252 4105 4027 4119
rect 2215 4096 2950 4105
tri 2950 4096 2959 4105 nw
tri 3229 4096 3238 4105 se
rect 3238 4096 4027 4105
rect 2215 4067 2921 4096
tri 2921 4067 2950 4096 nw
tri 3200 4067 3229 4096 se
rect 3229 4067 4027 4096
rect 2215 4053 2907 4067
tri 2907 4053 2921 4067 nw
tri 3186 4053 3200 4067 se
rect 3200 4053 4027 4067
rect 2215 4039 2893 4053
tri 2893 4039 2907 4053 nw
tri 3172 4039 3186 4053 se
rect 3186 4039 4027 4053
rect 2215 4015 2869 4039
tri 2869 4015 2893 4039 nw
tri 3148 4015 3172 4039 se
rect 3172 4015 4027 4039
rect 2215 3987 2841 4015
tri 2841 3987 2869 4015 nw
tri 3120 3987 3148 4015 se
rect 3148 3987 4027 4015
rect 2215 3973 2827 3987
tri 2827 3973 2841 3987 nw
tri 3106 3973 3120 3987 se
rect 3120 3973 4027 3987
rect 2215 3183 2815 3973
tri 2815 3961 2827 3973 nw
tri 3094 3961 3106 3973 se
rect 3106 3961 4027 3973
rect 2215 3127 2288 3183
rect 2344 3127 2368 3183
rect 2424 3127 2448 3183
rect 2504 3127 2528 3183
rect 2584 3127 2608 3183
rect 2664 3127 2688 3183
rect 2744 3127 2815 3183
rect 2215 3093 2815 3127
rect 2215 3037 2288 3093
rect 2344 3037 2368 3093
rect 2424 3037 2448 3093
rect 2504 3037 2528 3093
rect 2584 3037 2608 3093
rect 2664 3037 2688 3093
rect 2744 3037 2815 3093
rect 2215 3003 2815 3037
rect 2215 2947 2288 3003
rect 2344 2947 2368 3003
rect 2424 2947 2448 3003
rect 2504 2947 2528 3003
rect 2584 2947 2608 3003
rect 2664 2947 2688 3003
rect 2744 2947 2815 3003
rect 2215 2913 2815 2947
rect 2215 2857 2288 2913
rect 2344 2857 2368 2913
rect 2424 2857 2448 2913
rect 2504 2857 2528 2913
rect 2584 2857 2608 2913
rect 2664 2857 2688 2913
rect 2744 2857 2815 2913
rect 2215 2823 2815 2857
rect 2215 2767 2288 2823
rect 2344 2767 2368 2823
rect 2424 2767 2448 2823
rect 2504 2767 2528 2823
rect 2584 2767 2608 2823
rect 2664 2767 2688 2823
rect 2744 2767 2815 2823
rect 2215 2733 2815 2767
rect 2215 2677 2288 2733
rect 2344 2677 2368 2733
rect 2424 2677 2448 2733
rect 2504 2677 2528 2733
rect 2584 2677 2608 2733
rect 2664 2677 2688 2733
rect 2744 2677 2815 2733
rect 2215 2642 2815 2677
rect 2215 2586 2288 2642
rect 2344 2586 2368 2642
rect 2424 2586 2448 2642
rect 2504 2586 2528 2642
rect 2584 2586 2608 2642
rect 2664 2586 2688 2642
rect 2744 2586 2815 2642
rect 2215 2551 2815 2586
rect 2215 2495 2288 2551
rect 2344 2495 2368 2551
rect 2424 2495 2448 2551
rect 2504 2495 2528 2551
rect 2584 2495 2608 2551
rect 2664 2495 2688 2551
rect 2744 2495 2815 2551
tri 3085 3952 3094 3961 se
rect 3094 3952 4027 3961
rect 3085 3671 4027 3952
rect 3085 3661 4017 3671
tri 4017 3661 4027 3671 nw
rect 4121 4445 4126 4464
rect 4178 4445 4196 4497
rect 4248 4445 4266 4497
rect 4318 4445 4336 4497
rect 4388 4445 4406 4497
rect 4458 4445 4476 4497
rect 4528 4464 4530 4497
rect 4584 4464 4766 4538
rect 5322 4527 5346 4583
rect 5402 4527 5426 4583
rect 5482 4527 5506 4583
rect 5562 4527 5586 4583
rect 5642 4527 5666 4583
rect 5722 4527 5746 4583
rect 5266 4502 5802 4527
rect 4528 4445 5119 4464
tri 5119 4463 5120 4464 nw
rect 4121 4432 5119 4445
rect 4121 4380 4126 4432
rect 4178 4380 4196 4432
rect 4248 4380 4266 4432
rect 4318 4380 4336 4432
rect 4388 4380 4406 4432
rect 4458 4380 4476 4432
rect 4528 4380 5119 4432
rect 4121 4367 5119 4380
rect 4121 4315 4126 4367
rect 4178 4315 4196 4367
rect 4248 4315 4266 4367
rect 4318 4315 4336 4367
rect 4388 4315 4406 4367
rect 4458 4315 4476 4367
rect 4528 4315 5119 4367
rect 4121 4302 5119 4315
rect 4121 4250 4126 4302
rect 4178 4250 4196 4302
rect 4248 4250 4266 4302
rect 4318 4250 4336 4302
rect 4388 4250 4406 4302
rect 4458 4250 4476 4302
rect 4528 4250 5119 4302
rect 5231 4446 5266 4464
rect 5322 4446 5346 4502
rect 5402 4446 5426 4502
rect 5482 4446 5506 4502
rect 5562 4446 5586 4502
rect 5642 4446 5666 4502
rect 5722 4446 5746 4502
rect 6330 4464 6512 4538
rect 7725 4531 8190 4624
tri 8190 4531 8283 4624 nw
rect 8868 4579 8872 4635
rect 8928 4579 8952 4635
rect 9008 4579 9032 4635
rect 9088 4579 9112 4635
rect 9168 4579 9192 4635
rect 9248 4579 9272 4635
rect 9328 4579 9352 4635
rect 9408 4579 9412 4635
rect 8868 4553 9412 4579
tri 7682 4488 7725 4531 se
rect 7725 4488 8147 4531
tri 8147 4488 8190 4531 nw
rect 8868 4497 8872 4553
rect 8928 4497 8952 4553
rect 9008 4497 9032 4553
rect 9088 4497 9112 4553
rect 9168 4497 9192 4553
rect 9248 4497 9272 4553
rect 9328 4497 9352 4553
rect 9408 4497 9412 4553
rect 10716 5502 10740 5558
rect 10796 5502 10820 5558
rect 10876 5502 10900 5558
rect 10956 5502 10980 5558
rect 11036 5502 11060 5558
rect 11116 5502 11140 5558
rect 10660 5476 11196 5502
rect 10716 5420 10740 5476
rect 10796 5420 10820 5476
rect 10876 5420 10900 5476
rect 10956 5420 10980 5476
rect 11036 5420 11060 5476
rect 11116 5420 11140 5476
rect 12465 5558 13001 5567
rect 12521 5502 12545 5558
rect 12601 5502 12625 5558
rect 12681 5502 12705 5558
rect 12761 5502 12785 5558
rect 12841 5502 12865 5558
rect 12921 5502 12945 5558
rect 12465 5476 13001 5502
rect 10660 5393 11196 5420
tri 11320 5415 11350 5445 ne
tri 11402 5415 11432 5445 nw
rect 12521 5420 12545 5476
rect 12601 5420 12625 5476
rect 12681 5420 12705 5476
rect 12761 5420 12785 5476
rect 12841 5420 12865 5476
rect 12921 5420 12945 5476
rect 14278 5558 14814 5567
rect 14334 5502 14358 5558
rect 14414 5502 14438 5558
rect 14494 5502 14518 5558
rect 14574 5502 14598 5558
rect 14654 5502 14678 5558
rect 14734 5502 14758 5558
rect 14278 5476 14814 5502
rect 10716 5337 10740 5393
rect 10796 5337 10820 5393
rect 10876 5337 10900 5393
rect 10956 5337 10980 5393
rect 11036 5337 11060 5393
rect 11116 5337 11140 5393
rect 10660 5310 11196 5337
rect 10716 5254 10740 5310
rect 10796 5254 10820 5310
rect 10876 5254 10900 5310
rect 10956 5254 10980 5310
rect 11036 5254 11060 5310
rect 11116 5254 11140 5310
rect 10660 5227 11196 5254
rect 10716 5171 10740 5227
rect 10796 5171 10820 5227
rect 10876 5171 10900 5227
rect 10956 5171 10980 5227
rect 11036 5171 11060 5227
rect 11116 5171 11140 5227
rect 12465 5393 13001 5420
tri 13096 5415 13126 5445 ne
tri 13178 5415 13208 5445 nw
tri 14065 5415 14095 5445 ne
tri 14147 5415 14177 5445 nw
rect 14334 5420 14358 5476
rect 14414 5420 14438 5476
rect 14494 5420 14518 5476
rect 14574 5420 14598 5476
rect 14654 5420 14678 5476
rect 14734 5420 14758 5476
rect 12521 5337 12545 5393
rect 12601 5337 12625 5393
rect 12681 5337 12705 5393
rect 12761 5337 12785 5393
rect 12841 5337 12865 5393
rect 12921 5337 12945 5393
rect 12465 5310 13001 5337
rect 12521 5254 12545 5310
rect 12601 5254 12625 5310
rect 12681 5254 12705 5310
rect 12761 5254 12785 5310
rect 12841 5254 12865 5310
rect 12921 5254 12945 5310
rect 12465 5227 13001 5254
rect 10660 5144 11196 5171
tri 11320 5167 11350 5197 se
tri 11402 5167 11432 5197 sw
rect 12521 5171 12545 5227
rect 12601 5171 12625 5227
rect 12681 5171 12705 5227
rect 12761 5171 12785 5227
rect 12841 5171 12865 5227
rect 12921 5171 12945 5227
rect 14278 5393 14814 5420
rect 14334 5337 14358 5393
rect 14414 5337 14438 5393
rect 14494 5337 14518 5393
rect 14574 5337 14598 5393
rect 14654 5337 14678 5393
rect 14734 5337 14758 5393
rect 14278 5310 14814 5337
rect 14334 5254 14358 5310
rect 14414 5254 14438 5310
rect 14494 5254 14518 5310
rect 14574 5254 14598 5310
rect 14654 5254 14678 5310
rect 14734 5254 14758 5310
rect 14278 5227 14814 5254
rect 10716 5088 10740 5144
rect 10796 5088 10820 5144
rect 10876 5088 10900 5144
rect 10956 5088 10980 5144
rect 11036 5088 11060 5144
rect 11116 5088 11140 5144
rect 10660 5061 11196 5088
rect 10716 5005 10740 5061
rect 10796 5005 10820 5061
rect 10876 5005 10900 5061
rect 10956 5005 10980 5061
rect 11036 5005 11060 5061
rect 11116 5005 11140 5061
rect 10660 4978 11196 5005
rect 10716 4922 10740 4978
rect 10796 4922 10820 4978
rect 10876 4922 10900 4978
rect 10956 4922 10980 4978
rect 11036 4922 11060 4978
rect 11116 4922 11140 4978
rect 10660 4895 11196 4922
rect 10716 4839 10740 4895
rect 10796 4839 10820 4895
rect 10876 4839 10900 4895
rect 10956 4839 10980 4895
rect 11036 4839 11060 4895
rect 11116 4839 11140 4895
rect 10660 4812 11196 4839
rect 10716 4756 10740 4812
rect 10796 4756 10820 4812
rect 10876 4756 10900 4812
rect 10956 4756 10980 4812
rect 11036 4756 11060 4812
rect 11116 4756 11140 4812
rect 10660 4729 11196 4756
rect 10716 4673 10740 4729
rect 10796 4673 10820 4729
rect 10876 4673 10900 4729
rect 10956 4673 10980 4729
rect 11036 4673 11060 4729
rect 11116 4673 11140 4729
rect 10660 4646 11196 4673
rect 10716 4590 10740 4646
rect 10796 4590 10820 4646
rect 10876 4590 10900 4646
rect 10956 4590 10980 4646
rect 11036 4590 11060 4646
rect 11116 4590 11140 4646
rect 10660 4563 11196 4590
rect 8868 4488 9412 4497
tri 7658 4464 7682 4488 se
rect 7682 4464 8123 4488
tri 8123 4464 8147 4488 nw
rect 9024 4464 9246 4488
rect 9700 4464 9882 4538
rect 10716 4507 10740 4563
rect 10796 4507 10820 4563
rect 10876 4507 10900 4563
rect 10956 4507 10980 4563
rect 11036 4507 11060 4563
rect 11116 4507 11140 4563
rect 12465 5144 13001 5171
tri 13096 5167 13126 5197 se
tri 13178 5167 13208 5197 sw
tri 14065 5167 14095 5197 se
tri 14147 5167 14177 5197 sw
rect 14334 5171 14358 5227
rect 14414 5171 14438 5227
rect 14494 5171 14518 5227
rect 14574 5171 14598 5227
rect 14654 5171 14678 5227
rect 14734 5171 14758 5227
rect 12521 5088 12545 5144
rect 12601 5088 12625 5144
rect 12681 5088 12705 5144
rect 12761 5088 12785 5144
rect 12841 5088 12865 5144
rect 12921 5088 12945 5144
rect 12465 5061 13001 5088
rect 12521 5005 12545 5061
rect 12601 5005 12625 5061
rect 12681 5005 12705 5061
rect 12761 5005 12785 5061
rect 12841 5005 12865 5061
rect 12921 5005 12945 5061
rect 12465 4978 13001 5005
rect 12521 4922 12545 4978
rect 12601 4922 12625 4978
rect 12681 4922 12705 4978
rect 12761 4922 12785 4978
rect 12841 4922 12865 4978
rect 12921 4922 12945 4978
rect 12465 4895 13001 4922
rect 12521 4839 12545 4895
rect 12601 4839 12625 4895
rect 12681 4839 12705 4895
rect 12761 4839 12785 4895
rect 12841 4839 12865 4895
rect 12921 4839 12945 4895
rect 12465 4812 13001 4839
rect 12521 4756 12545 4812
rect 12601 4756 12625 4812
rect 12681 4756 12705 4812
rect 12761 4756 12785 4812
rect 12841 4756 12865 4812
rect 12921 4756 12945 4812
rect 12465 4729 13001 4756
rect 12521 4673 12545 4729
rect 12601 4673 12625 4729
rect 12681 4673 12705 4729
rect 12761 4673 12785 4729
rect 12841 4673 12865 4729
rect 12921 4673 12945 4729
rect 12465 4646 13001 4673
rect 12521 4590 12545 4646
rect 12601 4590 12625 4646
rect 12681 4590 12705 4646
rect 12761 4590 12785 4646
rect 12841 4590 12865 4646
rect 12921 4590 12945 4646
rect 12465 4563 13001 4590
rect 11196 4507 11243 4538
rect 11737 4535 11919 4538
rect 10660 4498 11243 4507
rect 11022 4464 11243 4498
rect 11338 4498 12338 4535
tri 12338 4498 12375 4535 sw
rect 12521 4507 12545 4563
rect 12601 4507 12625 4563
rect 12681 4507 12705 4563
rect 12761 4507 12785 4563
rect 12841 4507 12865 4563
rect 12921 4507 12945 4563
rect 12465 4498 13001 4507
rect 14278 5144 14814 5171
rect 14334 5088 14358 5144
rect 14414 5088 14438 5144
rect 14494 5088 14518 5144
rect 14574 5088 14598 5144
rect 14654 5088 14678 5144
rect 14734 5088 14758 5144
rect 14278 5061 14814 5088
rect 14334 5005 14358 5061
rect 14414 5005 14438 5061
rect 14494 5005 14518 5061
rect 14574 5005 14598 5061
rect 14654 5005 14678 5061
rect 14734 5005 14758 5061
rect 14278 4978 14814 5005
rect 14334 4922 14358 4978
rect 14414 4922 14438 4978
rect 14494 4922 14518 4978
rect 14574 4922 14598 4978
rect 14654 4922 14678 4978
rect 14734 4922 14758 4978
rect 14278 4895 14814 4922
rect 14334 4839 14358 4895
rect 14414 4839 14438 4895
rect 14494 4839 14518 4895
rect 14574 4839 14598 4895
rect 14654 4839 14678 4895
rect 14734 4839 14758 4895
rect 14278 4812 14814 4839
rect 14334 4756 14358 4812
rect 14414 4756 14438 4812
rect 14494 4756 14518 4812
rect 14574 4756 14598 4812
rect 14654 4756 14678 4812
rect 14734 4756 14758 4812
rect 14278 4729 14814 4756
rect 14334 4673 14358 4729
rect 14414 4673 14438 4729
rect 14494 4673 14518 4729
rect 14574 4673 14598 4729
rect 14654 4673 14678 4729
rect 14734 4673 14758 4729
rect 14278 4646 14814 4673
rect 14334 4590 14358 4646
rect 14414 4590 14438 4646
rect 14494 4590 14518 4646
rect 14574 4590 14598 4646
rect 14654 4590 14678 4646
rect 14734 4590 14758 4646
rect 14278 4563 14814 4590
rect 14334 4507 14358 4563
rect 14414 4507 14438 4563
rect 14494 4507 14518 4563
rect 14574 4507 14598 4563
rect 14654 4507 14678 4563
rect 14734 4507 14758 4563
rect 16064 5556 16520 5565
rect 16120 5500 16144 5556
rect 16200 5500 16224 5556
rect 16280 5500 16304 5556
rect 16360 5500 16384 5556
rect 16440 5500 16464 5556
rect 16064 5474 16520 5500
rect 16120 5418 16144 5474
rect 16200 5418 16224 5474
rect 16280 5418 16304 5474
rect 16360 5418 16384 5474
rect 16440 5418 16464 5474
rect 16064 5392 16520 5418
rect 16120 5336 16144 5392
rect 16200 5336 16224 5392
rect 16280 5336 16304 5392
rect 16360 5336 16384 5392
rect 16440 5336 16464 5392
rect 16064 5310 16520 5336
rect 16120 5254 16144 5310
rect 16200 5254 16224 5310
rect 16280 5254 16304 5310
rect 16360 5254 16384 5310
rect 16440 5254 16464 5310
rect 16064 5228 16520 5254
rect 16120 5172 16144 5228
rect 16200 5172 16224 5228
rect 16280 5172 16304 5228
rect 16360 5172 16384 5228
rect 16440 5172 16464 5228
rect 16064 5146 16520 5172
rect 16120 5090 16144 5146
rect 16200 5090 16224 5146
rect 16280 5090 16304 5146
rect 16360 5090 16384 5146
rect 16440 5090 16464 5146
rect 16064 5064 16520 5090
rect 16120 5008 16144 5064
rect 16200 5008 16224 5064
rect 16280 5008 16304 5064
rect 16360 5008 16384 5064
rect 16440 5008 16464 5064
rect 16064 4982 16520 5008
rect 16120 4926 16144 4982
rect 16200 4926 16224 4982
rect 16280 4926 16304 4982
rect 16360 4926 16384 4982
rect 16440 4926 16464 4982
rect 16064 4900 16520 4926
rect 16120 4844 16144 4900
rect 16200 4844 16224 4900
rect 16280 4844 16304 4900
rect 16360 4844 16384 4900
rect 16440 4844 16464 4900
rect 16064 4818 16520 4844
rect 16120 4762 16144 4818
rect 16200 4762 16224 4818
rect 16280 4762 16304 4818
rect 16360 4762 16384 4818
rect 16440 4762 16464 4818
rect 16064 4735 16520 4762
rect 16120 4679 16144 4735
rect 16200 4679 16224 4735
rect 16280 4679 16304 4735
rect 16360 4679 16384 4735
rect 16440 4679 16464 4735
rect 16064 4652 16520 4679
rect 16120 4596 16144 4652
rect 16200 4596 16224 4652
rect 16280 4596 16304 4652
rect 16360 4596 16384 4652
rect 16440 4596 16464 4652
rect 16064 4569 16520 4596
rect 14278 4498 14814 4507
rect 11338 4488 12375 4498
tri 12375 4488 12385 4498 sw
rect 11338 4464 12385 4488
tri 12385 4464 12409 4488 sw
rect 14436 4464 14658 4498
rect 15306 4464 15488 4538
rect 5802 4446 5831 4464
rect 5231 4425 5831 4446
tri 6154 4437 6181 4464 ne
rect 6181 4437 6918 4464
tri 7631 4437 7658 4464 se
rect 7658 4437 8096 4464
tri 8096 4437 8123 4464 nw
rect 8839 4463 9439 4464
rect 8839 4444 9420 4463
tri 9420 4444 9439 4463 nw
tri 9535 4444 9555 4464 ne
rect 9555 4444 10494 4464
tri 8832 4437 8839 4444 se
rect 8839 4437 9413 4444
tri 9413 4437 9420 4444 nw
tri 9555 4437 9562 4444 ne
rect 9562 4437 10494 4444
tri 10494 4437 10521 4464 nw
tri 11338 4437 11365 4464 ne
rect 11365 4437 12409 4464
tri 12409 4437 12436 4464 sw
tri 6181 4435 6183 4437 ne
rect 6183 4435 6918 4437
tri 7629 4435 7631 4437 se
rect 7631 4435 8084 4437
tri 5831 4425 5841 4435 sw
tri 6183 4425 6193 4435 ne
rect 6193 4425 6918 4435
tri 7619 4425 7629 4435 se
rect 7629 4425 8084 4435
tri 8084 4425 8096 4437 nw
tri 8820 4425 8832 4437 se
rect 8832 4425 9401 4437
tri 9401 4425 9413 4437 nw
tri 9562 4425 9574 4437 ne
rect 9574 4425 10482 4437
tri 10482 4425 10494 4437 nw
tri 11365 4425 11377 4437 ne
rect 11377 4425 12436 4437
rect 5231 4417 5841 4425
tri 5841 4417 5849 4425 sw
tri 6193 4417 6201 4425 ne
rect 6201 4417 6918 4425
tri 7611 4417 7619 4425 se
rect 7619 4417 7898 4425
rect 5231 4346 5849 4417
tri 5231 4293 5284 4346 ne
rect 5284 4293 5849 4346
tri 5849 4293 5973 4417 sw
tri 6201 4389 6229 4417 ne
rect 6229 4389 6918 4417
tri 7583 4389 7611 4417 se
rect 7611 4389 7898 4417
tri 6229 4293 6325 4389 ne
rect 6325 4293 6918 4389
tri 6918 4293 7014 4389 sw
tri 7487 4293 7583 4389 se
rect 7583 4293 7898 4389
rect 4121 4237 5119 4250
rect 4121 4185 4126 4237
rect 4178 4185 4196 4237
rect 4248 4185 4266 4237
rect 4318 4185 4336 4237
rect 4388 4185 4406 4237
rect 4458 4185 4476 4237
rect 4528 4185 5119 4237
rect 4121 4171 5119 4185
rect 4121 4119 4126 4171
rect 4178 4119 4196 4171
rect 4248 4119 4266 4171
rect 4318 4119 4336 4171
rect 4388 4119 4406 4171
rect 4458 4119 4476 4171
rect 4528 4119 5119 4171
tri 5284 4143 5434 4293 ne
rect 4121 4105 5119 4119
rect 4121 4053 4126 4105
rect 4178 4053 4196 4105
rect 4248 4053 4266 4105
rect 4318 4053 4336 4105
rect 4388 4053 4406 4105
rect 4458 4053 4476 4105
rect 4528 4053 5119 4105
rect 4121 4039 5119 4053
rect 4121 3987 4126 4039
rect 4178 3987 4196 4039
rect 4248 3987 4266 4039
rect 4318 3987 4336 4039
rect 4388 3987 4406 4039
rect 4458 3987 4476 4039
rect 4528 3987 5119 4039
rect 4121 3973 5119 3987
rect 4121 3921 4126 3973
rect 4178 3921 4196 3973
rect 4248 3921 4266 3973
rect 4318 3921 4336 3973
rect 4388 3921 4406 3973
rect 4458 3921 4476 3973
rect 4528 3921 5119 3973
rect 4121 3907 5119 3921
rect 4121 3855 4126 3907
rect 4178 3855 4196 3907
rect 4248 3855 4266 3907
rect 4318 3855 4336 3907
rect 4388 3855 4406 3907
rect 4458 3855 4476 3907
rect 4528 3855 5119 3907
rect 3085 3609 3965 3661
tri 3965 3609 4017 3661 nw
rect 3085 3575 3931 3609
tri 3931 3575 3965 3609 nw
rect 2215 2444 2815 2495
tri 3075 2486 3085 2496 se
rect 3085 2486 3918 3575
tri 3918 3562 3931 3575 nw
rect 4121 3138 5119 3855
rect 4121 3082 4228 3138
rect 4284 3082 4308 3138
rect 4364 3082 4388 3138
rect 4444 3082 4468 3138
rect 4524 3082 4548 3138
rect 4604 3082 4628 3138
rect 4684 3082 4708 3138
rect 4764 3082 4788 3138
rect 4844 3082 4868 3138
rect 4924 3082 4948 3138
rect 5004 3082 5028 3138
rect 5084 3082 5119 3138
rect 4121 3057 5119 3082
rect 4121 3001 4228 3057
rect 4284 3001 4308 3057
rect 4364 3001 4388 3057
rect 4444 3001 4468 3057
rect 4524 3001 4548 3057
rect 4604 3001 4628 3057
rect 4684 3001 4708 3057
rect 4764 3001 4788 3057
rect 4844 3001 4868 3057
rect 4924 3001 4948 3057
rect 5004 3001 5028 3057
rect 5084 3001 5119 3057
rect 4121 2976 5119 3001
rect 4121 2920 4228 2976
rect 4284 2920 4308 2976
rect 4364 2920 4388 2976
rect 4444 2920 4468 2976
rect 4524 2920 4548 2976
rect 4604 2920 4628 2976
rect 4684 2920 4708 2976
rect 4764 2920 4788 2976
rect 4844 2920 4868 2976
rect 4924 2920 4948 2976
rect 5004 2920 5028 2976
rect 5084 2920 5119 2976
rect 4121 2895 5119 2920
rect 4121 2839 4228 2895
rect 4284 2839 4308 2895
rect 4364 2839 4388 2895
rect 4444 2839 4468 2895
rect 4524 2839 4548 2895
rect 4604 2839 4628 2895
rect 4684 2839 4708 2895
rect 4764 2839 4788 2895
rect 4844 2839 4868 2895
rect 4924 2839 4948 2895
rect 5004 2839 5028 2895
rect 5084 2839 5119 2895
rect 4121 2814 5119 2839
rect 4121 2758 4228 2814
rect 4284 2758 4308 2814
rect 4364 2758 4388 2814
rect 4444 2758 4468 2814
rect 4524 2758 4548 2814
rect 4604 2758 4628 2814
rect 4684 2758 4708 2814
rect 4764 2758 4788 2814
rect 4844 2758 4868 2814
rect 4924 2758 4948 2814
rect 5004 2758 5028 2814
rect 5084 2758 5119 2814
rect 4121 2740 5119 2758
tri 4121 2668 4193 2740 ne
rect 4193 2733 5119 2740
rect 4193 2677 4228 2733
rect 4284 2677 4308 2733
rect 4364 2677 4388 2733
rect 4444 2677 4468 2733
rect 4524 2677 4548 2733
rect 4604 2677 4628 2733
rect 4684 2677 4708 2733
rect 4764 2677 4788 2733
rect 4844 2677 4868 2733
rect 4924 2677 4948 2733
rect 5004 2677 5028 2733
rect 5084 2677 5119 2733
tri 3033 2444 3075 2486 se
rect 3075 2444 3918 2486
rect 747 1203 1001 2444
tri 1001 2420 1025 2444 nw
tri 1293 2420 1317 2444 se
rect 1317 2420 2159 2444
tri 1081 2208 1293 2420 se
rect 1293 2208 2159 2420
rect 1081 2147 2159 2208
tri 2751 2162 3033 2444 se
rect 3033 2162 3918 2444
rect 1081 2034 1444 2147
tri 1444 2034 1557 2147 nw
rect 1081 2027 1437 2034
tri 1437 2027 1444 2034 nw
rect 1081 1832 1407 2027
tri 1407 1997 1437 2027 nw
rect 1583 2018 1903 2034
rect 1081 1780 1128 1832
rect 1180 1780 1192 1832
rect 1244 1780 1256 1832
rect 1308 1780 1320 1832
rect 1372 1780 1407 1832
rect 1081 1764 1407 1780
rect 1081 1712 1128 1764
rect 1180 1712 1192 1764
rect 1244 1712 1256 1764
rect 1308 1712 1320 1764
rect 1372 1712 1407 1764
rect 1081 1696 1407 1712
rect 1081 1644 1128 1696
rect 1180 1644 1192 1696
rect 1244 1644 1256 1696
rect 1308 1644 1320 1696
rect 1372 1644 1407 1696
rect 1081 1627 1407 1644
rect 1081 1575 1128 1627
rect 1180 1575 1192 1627
rect 1244 1575 1256 1627
rect 1308 1575 1320 1627
rect 1372 1575 1407 1627
rect 1081 1558 1407 1575
rect 1081 1506 1128 1558
rect 1180 1506 1192 1558
rect 1244 1506 1256 1558
rect 1308 1506 1320 1558
rect 1372 1506 1407 1558
rect 1081 1489 1407 1506
rect 1081 1437 1128 1489
rect 1180 1437 1192 1489
rect 1244 1437 1256 1489
rect 1308 1437 1320 1489
rect 1372 1437 1407 1489
rect 1081 1420 1407 1437
rect 1081 1368 1128 1420
rect 1180 1368 1192 1420
rect 1244 1368 1256 1420
rect 1308 1368 1320 1420
rect 1372 1368 1407 1420
rect 1583 1962 1594 2018
rect 1650 1962 1674 2018
rect 1730 1962 1754 2018
rect 1810 1962 1834 2018
rect 1890 1962 1903 2018
rect 1583 1932 1903 1962
rect 1583 1876 1594 1932
rect 1650 1876 1674 1932
rect 1730 1876 1754 1932
rect 1810 1876 1834 1932
rect 1890 1876 1903 1932
rect 1583 1846 1903 1876
rect 1583 1790 1594 1846
rect 1650 1790 1674 1846
rect 1730 1790 1754 1846
rect 1810 1790 1834 1846
rect 1890 1790 1903 1846
rect 1583 1760 1903 1790
rect 1583 1704 1594 1760
rect 1650 1704 1674 1760
rect 1730 1704 1754 1760
rect 1810 1704 1834 1760
rect 1890 1704 1903 1760
rect 1583 1674 1903 1704
rect 1583 1618 1594 1674
rect 1650 1618 1674 1674
rect 1730 1618 1754 1674
rect 1810 1618 1834 1674
rect 1890 1618 1903 1674
rect 1583 1587 1903 1618
rect 1583 1531 1594 1587
rect 1650 1531 1674 1587
rect 1730 1531 1754 1587
rect 1810 1531 1834 1587
rect 1890 1531 1903 1587
rect 1583 1500 1903 1531
rect 1583 1444 1594 1500
rect 1650 1444 1674 1500
rect 1730 1444 1754 1500
rect 1810 1444 1834 1500
rect 1890 1444 1903 1500
rect 1583 1413 1903 1444
rect 1583 1382 1594 1413
rect 1081 1351 1407 1368
rect 1081 1299 1128 1351
rect 1180 1299 1192 1351
rect 1244 1299 1256 1351
rect 1308 1299 1320 1351
rect 1372 1299 1407 1351
rect 1587 1357 1594 1382
rect 1650 1357 1674 1413
rect 1730 1357 1754 1413
rect 1810 1357 1834 1413
rect 1890 1382 1903 1413
rect 2403 2018 2723 2034
rect 2403 1962 2415 2018
rect 2471 1962 2495 2018
rect 2551 1962 2575 2018
rect 2631 1962 2655 2018
rect 2711 1962 2723 2018
rect 2403 1932 2723 1962
rect 2403 1876 2415 1932
rect 2471 1876 2495 1932
rect 2551 1876 2575 1932
rect 2631 1876 2655 1932
rect 2711 1876 2723 1932
rect 2403 1846 2723 1876
rect 2403 1790 2415 1846
rect 2471 1790 2495 1846
rect 2551 1790 2575 1846
rect 2631 1790 2655 1846
rect 2711 1790 2723 1846
rect 2403 1760 2723 1790
rect 2403 1704 2415 1760
rect 2471 1704 2495 1760
rect 2551 1704 2575 1760
rect 2631 1704 2655 1760
rect 2711 1704 2723 1760
rect 2403 1674 2723 1704
rect 2403 1618 2415 1674
rect 2471 1618 2495 1674
rect 2551 1618 2575 1674
rect 2631 1618 2655 1674
rect 2711 1618 2723 1674
rect 2403 1587 2723 1618
rect 2403 1531 2415 1587
rect 2471 1531 2495 1587
rect 2551 1531 2575 1587
rect 2631 1531 2655 1587
rect 2711 1531 2723 1587
rect 2403 1500 2723 1531
rect 2403 1444 2415 1500
rect 2471 1444 2495 1500
rect 2551 1444 2575 1500
rect 2631 1444 2655 1500
rect 2711 1444 2723 1500
rect 2403 1413 2723 1444
rect 2403 1382 2415 1413
rect 1890 1357 1897 1382
rect 1587 1348 1897 1357
rect 2408 1357 2415 1382
rect 2471 1357 2495 1413
rect 2551 1357 2575 1413
rect 2631 1357 2655 1413
rect 2711 1382 2723 1413
rect 2751 1851 3918 2162
rect 4193 2652 5119 2677
rect 4193 2596 4228 2652
rect 4284 2596 4308 2652
rect 4364 2596 4388 2652
rect 4444 2596 4468 2652
rect 4524 2596 4548 2652
rect 4604 2596 4628 2652
rect 4684 2596 4708 2652
rect 4764 2596 4788 2652
rect 4844 2596 4868 2652
rect 4924 2596 4948 2652
rect 5004 2596 5028 2652
rect 5084 2596 5119 2652
rect 4193 2571 5119 2596
rect 4193 2515 4228 2571
rect 4284 2515 4308 2571
rect 4364 2515 4388 2571
rect 4444 2515 4468 2571
rect 4524 2515 4548 2571
rect 4604 2515 4628 2571
rect 4684 2515 4708 2571
rect 4764 2515 4788 2571
rect 4844 2515 4868 2571
rect 4924 2515 4948 2571
rect 5004 2515 5028 2571
rect 5084 2515 5119 2571
rect 4193 2490 5119 2515
rect 4193 2434 4228 2490
rect 4284 2434 4308 2490
rect 4364 2434 4388 2490
rect 4444 2434 4468 2490
rect 4524 2434 4548 2490
rect 4604 2434 4628 2490
rect 4684 2434 4708 2490
rect 4764 2434 4788 2490
rect 4844 2434 4868 2490
rect 4924 2434 4948 2490
rect 5004 2434 5028 2490
rect 5084 2434 5119 2490
rect 4193 2408 5119 2434
rect 4193 2352 4228 2408
rect 4284 2352 4308 2408
rect 4364 2352 4388 2408
rect 4444 2352 4468 2408
rect 4524 2352 4548 2408
rect 4604 2352 4628 2408
rect 4684 2352 4708 2408
rect 4764 2352 4788 2408
rect 4844 2352 4868 2408
rect 4924 2352 4948 2408
rect 5004 2352 5028 2408
rect 5084 2352 5119 2408
rect 4193 2326 5119 2352
rect 4193 2270 4228 2326
rect 4284 2270 4308 2326
rect 4364 2270 4388 2326
rect 4444 2270 4468 2326
rect 4524 2270 4548 2326
rect 4604 2270 4628 2326
rect 4684 2270 4708 2326
rect 4764 2270 4788 2326
rect 4844 2270 4868 2326
rect 4924 2270 4948 2326
rect 5004 2270 5028 2326
rect 5084 2270 5119 2326
rect 4193 2244 5119 2270
rect 4193 2188 4228 2244
rect 4284 2188 4308 2244
rect 4364 2188 4388 2244
rect 4444 2188 4468 2244
rect 4524 2188 4548 2244
rect 4604 2188 4628 2244
rect 4684 2188 4708 2244
rect 4764 2188 4788 2244
rect 4844 2188 4868 2244
rect 4924 2188 4948 2244
rect 5004 2188 5028 2244
rect 5084 2188 5119 2244
rect 4193 2162 5119 2188
rect 4193 2106 4228 2162
rect 4284 2106 4308 2162
rect 4364 2106 4388 2162
rect 4444 2106 4468 2162
rect 4524 2106 4548 2162
rect 4604 2106 4628 2162
rect 4684 2106 4708 2162
rect 4764 2106 4788 2162
rect 4844 2106 4868 2162
rect 4924 2106 4948 2162
rect 5004 2106 5028 2162
rect 5084 2106 5119 2162
rect 4193 2080 5119 2106
rect 4193 2024 4228 2080
rect 4284 2024 4308 2080
rect 4364 2024 4388 2080
rect 4444 2024 4468 2080
rect 4524 2024 4548 2080
rect 4604 2024 4628 2080
rect 4684 2024 4708 2080
rect 4764 2024 4788 2080
rect 4844 2024 4868 2080
rect 4924 2024 4948 2080
rect 5004 2024 5028 2080
rect 5084 2024 5119 2080
rect 4193 1998 5119 2024
rect 4193 1942 4228 1998
rect 4284 1942 4308 1998
rect 4364 1942 4388 1998
rect 4444 1942 4468 1998
rect 4524 1942 4548 1998
rect 4604 1942 4628 1998
rect 4684 1942 4708 1998
rect 4764 1942 4788 1998
rect 4844 1942 4868 1998
rect 4924 1942 4948 1998
rect 5004 1942 5028 1998
rect 5084 1942 5119 1998
tri 3918 1851 3992 1925 sw
rect 4193 1916 5119 1942
rect 4193 1860 4228 1916
rect 4284 1860 4308 1916
rect 4364 1860 4388 1916
rect 4444 1860 4468 1916
rect 4524 1860 4548 1916
rect 4604 1860 4628 1916
rect 4684 1860 4708 1916
rect 4764 1860 4788 1916
rect 4844 1860 4868 1916
rect 4924 1860 4948 1916
rect 5004 1860 5028 1916
rect 5084 1860 5119 1916
rect 4193 1851 5119 1860
rect 5434 4141 5973 4293
tri 5973 4141 6125 4293 sw
tri 6325 4239 6379 4293 ne
rect 6379 4239 7014 4293
tri 7014 4239 7068 4293 sw
tri 7433 4239 7487 4293 se
rect 7487 4239 7898 4293
tri 7898 4239 8084 4425 nw
tri 8634 4239 8820 4425 se
rect 8820 4239 9213 4425
tri 6379 4141 6477 4239 ne
rect 6477 4141 7800 4239
tri 7800 4141 7898 4239 nw
tri 8632 4237 8634 4239 se
rect 8634 4237 9213 4239
tri 9213 4237 9401 4425 nw
rect 9574 4417 10474 4425
tri 10474 4417 10482 4425 nw
tri 11377 4417 11385 4425 ne
rect 11385 4417 12436 4425
tri 12436 4417 12456 4437 sw
rect 9574 4356 10413 4417
tri 10413 4356 10474 4417 nw
tri 11385 4356 11446 4417 ne
rect 11446 4356 12456 4417
rect 9574 4293 10350 4356
tri 10350 4293 10413 4356 nw
rect 10590 4340 10859 4356
tri 11446 4349 11453 4356 ne
rect 11453 4349 12456 4356
tri 12456 4349 12524 4417 sw
rect 8632 4141 9117 4237
tri 9117 4141 9213 4237 nw
rect 5434 4135 6125 4141
tri 6125 4135 6131 4141 sw
tri 6477 4135 6483 4141 ne
rect 6483 4135 7794 4141
tri 7794 4135 7800 4141 nw
rect 5434 4112 6131 4135
tri 6131 4112 6154 4135 sw
rect 5434 4083 6154 4112
tri 6154 4083 6183 4112 sw
rect 6262 4083 6268 4135
rect 6320 4083 6344 4135
rect 6396 4083 6402 4135
tri 6483 4112 6506 4135 ne
rect 6506 4112 7760 4135
tri 6506 4083 6535 4112 ne
rect 6535 4083 7760 4112
tri 7760 4101 7794 4135 nw
rect 8402 4083 8408 4135
rect 8460 4083 8472 4135
rect 8524 4083 8531 4135
rect 5434 4067 6183 4083
tri 6183 4067 6199 4083 sw
tri 6284 4067 6300 4083 ne
rect 6300 4067 6379 4083
tri 6379 4067 6395 4083 nw
tri 6535 4067 6551 4083 ne
rect 6551 4067 7760 4083
tri 8454 4067 8470 4083 ne
rect 8470 4067 8531 4083
rect 5434 4058 6199 4067
tri 6199 4058 6208 4067 sw
tri 6300 4058 6309 4067 ne
rect 6309 4058 6370 4067
tri 6370 4058 6379 4067 nw
tri 6551 4058 6560 4067 ne
rect 6560 4058 7760 4067
tri 8470 4058 8479 4067 ne
rect 5434 4050 6208 4058
tri 6208 4050 6216 4058 sw
tri 6309 4054 6313 4058 ne
rect 5434 1991 6216 4050
rect 6313 3661 6366 4058
tri 6366 4054 6370 4058 nw
tri 6560 4054 6564 4058 ne
rect 6564 4054 7760 4058
tri 6564 3978 6640 4054 ne
rect 6640 3978 7760 4054
tri 6640 3856 6762 3978 ne
tri 6366 3661 6399 3694 sw
rect 6313 3609 6319 3661
rect 6371 3609 6383 3661
rect 6435 3609 6441 3661
rect 6324 3358 6330 3410
rect 6382 3358 6394 3410
rect 6446 3358 6452 3410
tri 6377 3330 6405 3358 ne
rect 6405 2607 6452 3358
rect 6762 3149 7760 3978
rect 6762 3093 6798 3149
rect 6854 3093 6884 3149
rect 6940 3093 6970 3149
rect 7026 3093 7056 3149
rect 7112 3093 7142 3149
rect 7198 3093 7228 3149
rect 7284 3093 7314 3149
rect 7370 3093 7400 3149
rect 7456 3093 7486 3149
rect 7542 3093 7572 3149
rect 7628 3093 7657 3149
rect 7713 3093 7760 3149
rect 6762 3069 7760 3093
rect 6762 3013 6798 3069
rect 6854 3013 6884 3069
rect 6940 3013 6970 3069
rect 7026 3013 7056 3069
rect 7112 3013 7142 3069
rect 7198 3013 7228 3069
rect 7284 3013 7314 3069
rect 7370 3013 7400 3069
rect 7456 3013 7486 3069
rect 7542 3013 7572 3069
rect 7628 3013 7657 3069
rect 7713 3013 7760 3069
rect 6762 2989 7760 3013
rect 6762 2933 6798 2989
rect 6854 2933 6884 2989
rect 6940 2933 6970 2989
rect 7026 2933 7056 2989
rect 7112 2933 7142 2989
rect 7198 2933 7228 2989
rect 7284 2933 7314 2989
rect 7370 2933 7400 2989
rect 7456 2933 7486 2989
rect 7542 2933 7572 2989
rect 7628 2933 7657 2989
rect 7713 2933 7760 2989
rect 6762 2909 7760 2933
rect 6762 2853 6798 2909
rect 6854 2853 6884 2909
rect 6940 2853 6970 2909
rect 7026 2853 7056 2909
rect 7112 2853 7142 2909
rect 7198 2853 7228 2909
rect 7284 2853 7314 2909
rect 7370 2853 7400 2909
rect 7456 2853 7486 2909
rect 7542 2853 7572 2909
rect 7628 2853 7657 2909
rect 7713 2853 7760 2909
rect 6762 2829 7760 2853
rect 6762 2773 6798 2829
rect 6854 2773 6884 2829
rect 6940 2773 6970 2829
rect 7026 2773 7056 2829
rect 7112 2773 7142 2829
rect 7198 2773 7228 2829
rect 7284 2773 7314 2829
rect 7370 2773 7400 2829
rect 7456 2773 7486 2829
rect 7542 2773 7572 2829
rect 7628 2773 7657 2829
rect 7713 2773 7760 2829
rect 6762 2749 7760 2773
rect 6762 2693 6798 2749
rect 6854 2693 6884 2749
rect 6940 2693 6970 2749
rect 7026 2693 7056 2749
rect 7112 2693 7142 2749
rect 7198 2693 7228 2749
rect 7284 2693 7314 2749
rect 7370 2693 7400 2749
rect 7456 2693 7486 2749
rect 7542 2693 7572 2749
rect 7628 2693 7657 2749
rect 7713 2693 7760 2749
rect 6762 2669 7760 2693
tri 6405 2583 6429 2607 ne
rect 6429 2583 6452 2607
tri 6452 2583 6503 2634 sw
rect 6762 2613 6798 2669
rect 6854 2613 6884 2669
rect 6940 2613 6970 2669
rect 7026 2613 7056 2669
rect 7112 2613 7142 2669
rect 7198 2613 7228 2669
rect 7284 2613 7314 2669
rect 7370 2613 7400 2669
rect 7456 2613 7486 2669
rect 7542 2613 7572 2669
rect 7628 2613 7657 2669
rect 7713 2613 7760 2669
rect 8234 3523 8240 3575
rect 8292 3523 8304 3575
rect 8356 3523 8362 3575
rect 6762 2589 7760 2613
tri 6429 2560 6452 2583 ne
rect 6452 2560 6503 2583
tri 6452 2509 6503 2560 ne
tri 6503 2509 6577 2583 sw
rect 6762 2533 6798 2589
rect 6854 2533 6884 2589
rect 6940 2533 6970 2589
rect 7026 2533 7056 2589
rect 7112 2533 7142 2589
rect 7198 2533 7228 2589
rect 7284 2533 7314 2589
rect 7370 2533 7400 2589
rect 7456 2533 7486 2589
rect 7542 2533 7572 2589
rect 7628 2533 7657 2589
rect 7713 2533 7760 2589
tri 8160 2541 8234 2615 se
rect 8234 2593 8286 3523
tri 8286 3498 8311 3523 nw
tri 8234 2541 8286 2593 nw
tri 6503 2435 6577 2509 ne
tri 6577 2435 6651 2509 sw
rect 6762 2495 7760 2533
tri 8144 2525 8160 2541 se
tri 8128 2509 8144 2525 se
rect 8144 2509 8160 2525
tri 8114 2495 8128 2509 se
rect 8128 2495 8160 2509
tri 8086 2467 8114 2495 se
rect 8114 2467 8160 2495
tri 8160 2467 8234 2541 nw
tri 8054 2435 8086 2467 se
tri 6577 2361 6651 2435 ne
tri 6651 2361 6725 2435 sw
tri 8012 2393 8054 2435 se
rect 8054 2393 8086 2435
tri 8086 2393 8160 2467 nw
tri 7980 2361 8012 2393 se
tri 6651 2287 6725 2361 ne
tri 6725 2287 6799 2361 sw
tri 7938 2319 7980 2361 se
rect 7980 2319 8012 2361
tri 8012 2319 8086 2393 nw
tri 7906 2287 7938 2319 se
tri 6725 2213 6799 2287 ne
tri 6799 2213 6873 2287 sw
tri 7864 2245 7906 2287 se
rect 7906 2245 7938 2287
tri 7938 2245 8012 2319 nw
tri 7832 2213 7864 2245 se
tri 6799 2139 6873 2213 ne
tri 6873 2139 6947 2213 sw
tri 7790 2171 7832 2213 se
rect 7832 2171 7864 2213
tri 7864 2171 7938 2245 nw
tri 7758 2139 7790 2171 se
tri 6873 2065 6947 2139 ne
tri 6947 2065 7021 2139 sw
tri 7716 2097 7758 2139 se
rect 7758 2097 7790 2139
tri 7790 2097 7864 2171 nw
tri 7684 2065 7716 2097 se
tri 6947 2001 7011 2065 ne
rect 7011 2001 7021 2065
tri 6216 1991 6226 2001 sw
tri 7011 1991 7021 2001 ne
tri 7021 1991 7095 2065 sw
tri 7642 2023 7684 2065 se
rect 7684 2023 7716 2065
tri 7716 2023 7790 2097 nw
tri 7610 1991 7642 2023 se
rect 5434 1917 6226 1991
tri 6226 1917 6300 1991 sw
tri 7021 1917 7095 1991 ne
tri 7095 1917 7169 1991 sw
tri 7568 1949 7610 1991 se
rect 7610 1949 7642 1991
tri 7642 1949 7716 2023 nw
rect 5434 1895 6300 1917
tri 6300 1895 6322 1917 sw
tri 7095 1895 7117 1917 ne
rect 5434 1851 6322 1895
tri 6322 1851 6366 1895 sw
rect 2751 1849 3992 1851
rect 2751 1771 3121 1849
tri 3121 1771 3199 1849 nw
tri 3424 1771 3502 1849 ne
rect 3502 1771 3992 1849
tri 3992 1771 4072 1851 sw
rect 5434 1771 6366 1851
tri 6366 1771 6446 1851 sw
rect 2751 1750 3100 1771
tri 3100 1750 3121 1771 nw
tri 3502 1750 3523 1771 ne
rect 3523 1763 4072 1771
tri 4072 1763 4080 1771 sw
rect 3523 1750 4080 1763
tri 4080 1750 4093 1763 sw
rect 4235 1750 4755 1763
rect 2751 1744 3094 1750
tri 3094 1744 3100 1750 nw
tri 3523 1744 3529 1750 ne
rect 3529 1744 4093 1750
tri 4093 1744 4099 1750 sw
rect 2751 1702 3052 1744
tri 3052 1702 3094 1744 nw
tri 3529 1710 3563 1744 ne
rect 3563 1710 4099 1744
rect 3155 1702 3301 1710
tri 3301 1702 3309 1710 sw
tri 3563 1702 3571 1710 ne
rect 3571 1702 4099 1710
rect 2751 1698 3048 1702
tri 3048 1698 3052 1702 nw
rect 3155 1698 3309 1702
tri 3309 1698 3313 1702 sw
tri 3571 1698 3575 1702 ne
rect 3575 1698 4099 1702
rect 2711 1357 2718 1382
rect 2408 1348 2718 1357
rect 1081 1282 1407 1299
rect 1081 1230 1128 1282
rect 1180 1230 1192 1282
rect 1244 1230 1256 1282
rect 1308 1230 1320 1282
rect 1372 1230 1407 1282
rect 1081 1212 1407 1230
tri 1001 1203 1009 1211 sw
rect 747 1191 1009 1203
tri 1009 1191 1021 1203 sw
rect 747 1139 1021 1191
tri 1021 1139 1073 1191 sw
rect 747 1127 1073 1139
tri 1073 1127 1085 1139 sw
rect 747 1120 1085 1127
tri 1085 1120 1092 1127 sw
rect 747 1068 1092 1120
tri 1092 1068 1144 1120 sw
tri -119 867 -81 905 sw
rect -209 815 -203 867
rect -151 815 -139 867
rect -87 815 -81 867
rect 747 490 1041 1068
tri 747 480 757 490 ne
rect 757 480 1041 490
tri 757 428 809 480 ne
rect 809 428 1041 480
tri 809 384 853 428 ne
rect 853 384 1041 428
tri 853 372 865 384 ne
rect 865 372 1041 384
tri 865 320 917 372 ne
rect 917 320 1041 372
tri 917 308 929 320 ne
rect 929 308 1041 320
tri 929 276 961 308 ne
rect 961 276 1041 308
rect 2751 824 3047 1698
tri 3047 1697 3048 1698 nw
rect 3155 1693 3313 1698
rect 3155 1637 3161 1693
rect 3217 1637 3241 1693
rect 3297 1682 3313 1693
tri 3313 1682 3329 1698 sw
tri 3575 1682 3591 1698 ne
rect 3591 1682 4099 1698
rect 3297 1637 3329 1682
rect 3155 1630 3329 1637
tri 3329 1630 3381 1682 sw
tri 3591 1630 3643 1682 ne
rect 3643 1630 4099 1682
rect 3155 1614 3381 1630
tri 3381 1614 3397 1630 sw
tri 3643 1614 3659 1630 ne
rect 3659 1614 4099 1630
rect 3155 1601 3397 1614
rect 3155 1545 3161 1601
rect 3217 1545 3241 1601
rect 3297 1574 3397 1601
tri 3397 1574 3437 1614 sw
tri 3659 1574 3699 1614 ne
rect 3297 1562 3437 1574
tri 3437 1562 3449 1574 sw
rect 3297 1545 3449 1562
tri 3449 1545 3466 1562 sw
rect 3155 1539 3466 1545
tri 3466 1539 3472 1545 sw
rect 3155 1536 3472 1539
tri 3472 1536 3475 1539 sw
rect 3155 1530 3475 1536
rect 3155 1508 3321 1530
rect 3155 1452 3161 1508
rect 3217 1452 3241 1508
rect 3297 1474 3321 1508
rect 3377 1474 3401 1530
rect 3457 1474 3475 1530
rect 3297 1452 3475 1474
rect 3155 1418 3475 1452
rect 3155 1415 3321 1418
rect 3155 1382 3161 1415
rect 3159 1359 3161 1382
rect 3217 1359 3241 1415
rect 3297 1382 3321 1415
rect 3297 1359 3299 1382
rect 3159 1350 3299 1359
rect 3314 1362 3321 1382
rect 3377 1362 3401 1418
rect 3457 1382 3475 1418
rect 3699 1382 4099 1614
rect 4235 1698 4243 1750
rect 4295 1698 4307 1750
rect 4359 1698 4371 1750
rect 4423 1698 4435 1750
rect 4487 1698 4499 1750
rect 4551 1698 4563 1750
rect 4615 1698 4627 1750
rect 4679 1698 4691 1750
rect 4743 1698 4755 1750
rect 4235 1682 4755 1698
rect 4235 1630 4243 1682
rect 4295 1630 4307 1682
rect 4359 1630 4371 1682
rect 4423 1630 4435 1682
rect 4487 1630 4499 1682
rect 4551 1630 4563 1682
rect 4615 1630 4627 1682
rect 4679 1630 4691 1682
rect 4743 1630 4755 1682
rect 4235 1614 4755 1630
rect 4235 1562 4243 1614
rect 4295 1562 4307 1614
rect 4359 1562 4371 1614
rect 4423 1562 4435 1614
rect 4487 1562 4499 1614
rect 4551 1562 4563 1614
rect 4615 1562 4627 1614
rect 4679 1562 4691 1614
rect 4743 1562 4755 1614
rect 4235 1545 4755 1562
rect 4235 1493 4243 1545
rect 4295 1493 4307 1545
rect 4359 1493 4371 1545
rect 4423 1493 4435 1545
rect 4487 1493 4499 1545
rect 4551 1493 4563 1545
rect 4615 1493 4627 1545
rect 4679 1493 4691 1545
rect 4743 1493 4755 1545
rect 4235 1476 4755 1493
rect 4235 1424 4243 1476
rect 4295 1424 4307 1476
rect 4359 1424 4371 1476
rect 4423 1424 4435 1476
rect 4487 1424 4499 1476
rect 4551 1424 4563 1476
rect 4615 1424 4627 1476
rect 4679 1424 4691 1476
rect 4743 1424 4755 1476
rect 4235 1407 4755 1424
rect 3457 1362 3464 1382
rect 3314 1353 3464 1362
rect 4235 1355 4243 1407
rect 4295 1355 4307 1407
rect 4359 1355 4371 1407
rect 4423 1355 4435 1407
rect 4487 1355 4499 1407
rect 4551 1355 4563 1407
rect 4615 1355 4627 1407
rect 4679 1355 4691 1407
rect 4743 1355 4755 1407
rect 2751 -752 2787 824
rect 3003 -752 3047 824
rect 4235 1338 4755 1355
rect 4235 1286 4243 1338
rect 4295 1286 4307 1338
rect 4359 1286 4371 1338
rect 4423 1286 4435 1338
rect 4487 1286 4499 1338
rect 4551 1286 4563 1338
rect 4615 1286 4627 1338
rect 4679 1286 4691 1338
rect 4743 1286 4755 1338
rect 4235 1269 4755 1286
rect 4235 1217 4243 1269
rect 4295 1217 4307 1269
rect 4359 1217 4371 1269
rect 4423 1217 4435 1269
rect 4487 1217 4499 1269
rect 4551 1217 4563 1269
rect 4615 1217 4627 1269
rect 4679 1217 4691 1269
rect 4743 1217 4755 1269
rect 4235 291 4755 1217
rect 5434 1756 6446 1771
tri 6446 1756 6461 1771 sw
rect 5434 1719 6461 1756
tri 6461 1719 6498 1756 sw
rect 5434 1707 6498 1719
tri 6498 1707 6510 1719 sw
rect 5434 1655 6510 1707
tri 6510 1655 6562 1707 sw
rect 5434 1643 6562 1655
tri 6562 1643 6574 1655 sw
rect 5434 1600 6574 1643
tri 6574 1600 6617 1643 sw
tri 5420 1068 5434 1082 se
rect 5434 1068 6617 1600
rect 6924 1068 6930 1120
rect 6982 1068 6996 1120
rect 7048 1068 7054 1120
tri 5257 905 5420 1068 se
rect 5420 905 6617 1068
tri 6947 1041 6974 1068 ne
tri 5185 833 5257 905 se
rect 5257 833 6617 905
tri 5179 827 5185 833 se
rect 5185 827 6617 833
rect 5179 725 6617 827
tri 6947 642 6974 669 se
rect 6974 642 7027 1068
tri 7027 1041 7054 1068 nw
rect 7117 693 7169 1917
tri 7536 1917 7568 1949 se
rect 7568 1917 7610 1949
tri 7610 1917 7642 1949 nw
tri 7169 720 7194 745 sw
tri 7027 642 7054 669 sw
rect 6924 590 6930 642
rect 6982 590 6996 642
rect 7048 590 7054 642
tri 7511 560 7536 585 se
rect 7536 560 7588 1917
tri 7588 1895 7610 1917 nw
rect 7782 1831 8262 1842
rect 7782 1775 7794 1831
rect 7850 1775 7874 1831
rect 7930 1775 7954 1831
rect 8010 1775 8034 1831
rect 8090 1775 8114 1831
rect 8170 1775 8194 1831
rect 8250 1775 8262 1831
rect 7782 1748 8262 1775
rect 7782 1692 7794 1748
rect 7850 1692 7874 1748
rect 7930 1692 7954 1748
rect 8010 1692 8034 1748
rect 8090 1692 8114 1748
rect 8170 1692 8194 1748
rect 8250 1692 8262 1748
rect 7782 1665 8262 1692
rect 7782 1609 7794 1665
rect 7850 1609 7874 1665
rect 7930 1609 7954 1665
rect 8010 1609 8034 1665
rect 8090 1609 8114 1665
rect 8170 1609 8194 1665
rect 8250 1609 8262 1665
rect 7782 1582 8262 1609
rect 7782 1526 7794 1582
rect 7850 1526 7874 1582
rect 7930 1526 7954 1582
rect 8010 1526 8034 1582
rect 8090 1526 8114 1582
rect 8170 1526 8194 1582
rect 8250 1526 8262 1582
rect 7782 1498 8262 1526
rect 7782 1442 7794 1498
rect 7850 1442 7874 1498
rect 7930 1442 7954 1498
rect 8010 1442 8034 1498
rect 8090 1442 8114 1498
rect 8170 1442 8194 1498
rect 8250 1442 8262 1498
rect 7782 1414 8262 1442
rect 7782 1358 7794 1414
rect 7850 1358 7874 1414
rect 7930 1358 7954 1414
rect 8010 1358 8034 1414
rect 8090 1358 8114 1414
rect 8170 1358 8194 1414
rect 8250 1358 8262 1414
rect 7782 1065 8262 1358
rect 7423 508 7429 560
rect 7481 508 7493 560
rect 7545 508 7588 560
rect 8479 291 8531 4067
rect 8632 4132 9087 4141
rect 8632 4076 8675 4132
rect 8731 4076 8755 4132
rect 8811 4076 8835 4132
rect 8891 4076 8915 4132
rect 8971 4076 8995 4132
rect 9051 4076 9087 4132
tri 9087 4111 9117 4141 nw
rect 8632 4048 9087 4076
rect 8632 3992 8675 4048
rect 8731 3992 8755 4048
rect 8811 3992 8835 4048
rect 8891 3992 8915 4048
rect 8971 3992 8995 4048
rect 9051 3992 9087 4048
rect 8632 3964 9087 3992
rect 8632 3908 8675 3964
rect 8731 3908 8755 3964
rect 8811 3908 8835 3964
rect 8891 3908 8915 3964
rect 8971 3908 8995 3964
rect 9051 3908 9087 3964
rect 8632 3880 9087 3908
rect 8632 3824 8675 3880
rect 8731 3824 8755 3880
rect 8811 3824 8835 3880
rect 8891 3824 8915 3880
rect 8971 3824 8995 3880
rect 9051 3824 9087 3880
rect 8632 3795 9087 3824
rect 8632 3739 8675 3795
rect 8731 3739 8755 3795
rect 8811 3739 8835 3795
rect 8891 3739 8915 3795
rect 8971 3739 8995 3795
rect 9051 3739 9087 3795
rect 8632 2169 9087 3739
rect 9386 3609 9392 3661
rect 9444 3609 9456 3661
rect 9508 3609 9514 3661
tri 9437 3584 9462 3609 ne
rect 9189 3121 9195 3173
rect 9247 3121 9259 3173
rect 9311 3121 9317 3173
tri 9189 3091 9219 3121 ne
tri 9087 2169 9113 2195 sw
rect 8632 1301 9113 2169
rect 8633 822 9111 843
rect 8633 770 8639 822
rect 8691 770 8722 822
rect 8774 770 8805 822
rect 8857 770 8888 822
rect 8940 770 8971 822
rect 9023 770 9053 822
rect 9105 770 9111 822
rect 8633 749 9111 770
tri 9169 480 9219 530 se
rect 9219 480 9271 3121
tri 9271 3091 9301 3121 nw
tri 9271 480 9296 505 sw
rect 9169 428 9175 480
rect 9227 428 9239 480
rect 9291 428 9297 480
rect 9462 291 9514 3609
rect 9574 3145 10345 4293
tri 10345 4288 10350 4293 nw
rect 10590 3964 10609 4340
rect 10825 3964 10859 4340
tri 11453 4242 11560 4349 ne
rect 11560 4242 12524 4349
tri 12020 4204 12058 4242 ne
rect 12058 4204 12524 4242
tri 12524 4204 12669 4349 sw
tri 12058 4117 12145 4204 ne
rect 12145 4117 12669 4204
tri 12145 4085 12177 4117 ne
rect 10590 3939 10859 3964
rect 10590 3883 10609 3939
rect 10665 3883 10689 3939
rect 10745 3883 10769 3939
rect 10825 3883 10859 3939
rect 10590 3858 10859 3883
rect 10590 3802 10609 3858
rect 10665 3802 10689 3858
rect 10745 3802 10769 3858
rect 10825 3802 10859 3858
rect 10590 3777 10859 3802
rect 10590 3721 10609 3777
rect 10665 3721 10689 3777
rect 10745 3721 10769 3777
rect 10825 3721 10859 3777
rect 9574 3089 9602 3145
rect 9658 3089 9682 3145
rect 9738 3089 9762 3145
rect 9818 3089 9842 3145
rect 9898 3089 9922 3145
rect 9978 3089 10002 3145
rect 10058 3089 10082 3145
rect 10138 3089 10162 3145
rect 10218 3089 10242 3145
rect 10298 3089 10345 3145
rect 9574 3058 10345 3089
rect 9574 3002 9602 3058
rect 9658 3002 9682 3058
rect 9738 3002 9762 3058
rect 9818 3002 9842 3058
rect 9898 3002 9922 3058
rect 9978 3002 10002 3058
rect 10058 3002 10082 3058
rect 10138 3002 10162 3058
rect 10218 3002 10242 3058
rect 10298 3002 10345 3058
rect 9574 2971 10345 3002
rect 9574 2915 9602 2971
rect 9658 2915 9682 2971
rect 9738 2915 9762 2971
rect 9818 2915 9842 2971
rect 9898 2915 9922 2971
rect 9978 2915 10002 2971
rect 10058 2915 10082 2971
rect 10138 2915 10162 2971
rect 10218 2915 10242 2971
rect 10298 2915 10345 2971
rect 9574 2884 10345 2915
rect 9574 2828 9602 2884
rect 9658 2828 9682 2884
rect 9738 2828 9762 2884
rect 9818 2828 9842 2884
rect 9898 2828 9922 2884
rect 9978 2828 10002 2884
rect 10058 2828 10082 2884
rect 10138 2828 10162 2884
rect 10218 2828 10242 2884
rect 10298 2828 10345 2884
rect 9574 2797 10345 2828
rect 9574 2741 9602 2797
rect 9658 2741 9682 2797
rect 9738 2741 9762 2797
rect 9818 2741 9842 2797
rect 9898 2741 9922 2797
rect 9978 2741 10002 2797
rect 10058 2741 10082 2797
rect 10138 2741 10162 2797
rect 10218 2741 10242 2797
rect 10298 2741 10345 2797
rect 9574 2710 10345 2741
rect 9574 2654 9602 2710
rect 9658 2654 9682 2710
rect 9738 2654 9762 2710
rect 9818 2654 9842 2710
rect 9898 2654 9922 2710
rect 9978 2654 10002 2710
rect 10058 2654 10082 2710
rect 10138 2654 10162 2710
rect 10218 2654 10242 2710
rect 10298 2654 10345 2710
rect 9574 2623 10345 2654
rect 9574 2567 9602 2623
rect 9658 2567 9682 2623
rect 9738 2567 9762 2623
rect 9818 2567 9842 2623
rect 9898 2567 9922 2623
rect 9978 2567 10002 2623
rect 10058 2567 10082 2623
rect 10138 2567 10162 2623
rect 10218 2567 10242 2623
rect 10298 2567 10345 2623
rect 9574 2536 10345 2567
rect 9574 2480 9602 2536
rect 9658 2480 9682 2536
rect 9738 2480 9762 2536
rect 9818 2480 9842 2536
rect 9898 2480 9922 2536
rect 9978 2480 10002 2536
rect 10058 2480 10082 2536
rect 10138 2480 10162 2536
rect 10218 2480 10242 2536
rect 10298 2480 10345 2536
rect 9574 2448 10345 2480
rect 9574 2392 9602 2448
rect 9658 2392 9682 2448
rect 9738 2392 9762 2448
rect 9818 2392 9842 2448
rect 9898 2392 9922 2448
rect 9978 2392 10002 2448
rect 10058 2392 10082 2448
rect 10138 2392 10162 2448
rect 10218 2392 10242 2448
rect 10298 2392 10345 2448
rect 9574 2360 10345 2392
rect 9574 2304 9602 2360
rect 9658 2304 9682 2360
rect 9738 2304 9762 2360
rect 9818 2304 9842 2360
rect 9898 2304 9922 2360
rect 9978 2304 10002 2360
rect 10058 2304 10082 2360
rect 10138 2304 10162 2360
rect 10218 2304 10242 2360
rect 10298 2304 10345 2360
rect 9574 2272 10345 2304
rect 9574 2216 9602 2272
rect 9658 2216 9682 2272
rect 9738 2216 9762 2272
rect 9818 2216 9842 2272
rect 9898 2216 9922 2272
rect 9978 2216 10002 2272
rect 10058 2216 10082 2272
rect 10138 2216 10162 2272
rect 10218 2216 10242 2272
rect 10298 2216 10345 2272
rect 9574 2167 10345 2216
rect 10434 3438 10440 3490
rect 10492 3438 10504 3490
rect 10556 3438 10562 3490
tri 10407 2073 10434 2100 se
rect 10434 2073 10562 3438
rect 9698 2049 9989 2073
tri 10392 2058 10407 2073 se
rect 10407 2058 10562 2073
rect 9698 1993 9735 2049
rect 9791 1993 9815 2049
rect 9871 1993 9895 2049
rect 9951 1993 9989 2049
rect 9698 1959 9989 1993
tri 10299 1965 10392 2058 se
rect 10392 2046 10562 2058
rect 10392 1965 10481 2046
tri 10481 1965 10562 2046 nw
rect 9698 1903 9735 1959
rect 9791 1903 9815 1959
rect 9871 1903 9895 1959
rect 9951 1903 9989 1959
tri 10252 1918 10299 1965 se
rect 10299 1937 10453 1965
tri 10453 1937 10481 1965 nw
tri 10562 1937 10590 1965 se
rect 10590 1937 10859 3721
rect 10299 1918 10434 1937
tri 10434 1918 10453 1937 nw
tri 10543 1918 10562 1937 se
rect 10562 1918 10859 1937
rect 9698 1869 9989 1903
rect 9698 1813 9735 1869
rect 9791 1813 9815 1869
rect 9871 1813 9895 1869
rect 9951 1813 9989 1869
rect 9698 1779 9989 1813
rect 9698 1723 9735 1779
rect 9791 1723 9815 1779
rect 9871 1723 9895 1779
rect 9951 1723 9989 1779
rect 9698 1689 9989 1723
rect 9698 1633 9735 1689
rect 9791 1633 9815 1689
rect 9871 1633 9895 1689
rect 9951 1633 9989 1689
rect 9698 1599 9989 1633
rect 9698 1543 9735 1599
rect 9791 1543 9815 1599
rect 9871 1543 9895 1599
rect 9951 1543 9989 1599
rect 9698 1509 9989 1543
rect 9698 1453 9735 1509
rect 9791 1453 9815 1509
rect 9871 1453 9895 1509
rect 9951 1453 9989 1509
rect 9698 1418 9989 1453
rect 9698 1362 9735 1418
rect 9791 1362 9815 1418
rect 9871 1362 9895 1418
rect 9951 1362 9989 1418
rect 2751 -777 3047 -752
rect 2751 -833 2787 -777
rect 2843 -833 2867 -777
rect 2923 -833 2947 -777
rect 3003 -833 3047 -777
rect 2751 -858 3047 -833
rect 2751 -914 2787 -858
rect 2843 -914 2867 -858
rect 2923 -914 2947 -858
rect 3003 -914 3047 -858
rect 2751 -939 3047 -914
rect 2751 -995 2787 -939
rect 2843 -995 2867 -939
rect 2923 -995 2947 -939
rect 3003 -995 3047 -939
rect 2751 -1020 3047 -995
rect 2751 -1076 2787 -1020
rect 2843 -1076 2867 -1020
rect 2923 -1076 2947 -1020
rect 3003 -1076 3047 -1020
rect 2751 -1094 3047 -1076
rect 2751 -1146 2764 -1094
rect 2816 -1101 2837 -1094
rect 2889 -1101 2910 -1094
rect 2962 -1101 2982 -1094
rect 3034 -1146 3047 -1094
rect 2751 -1157 2787 -1146
rect 2843 -1157 2867 -1146
rect 2923 -1157 2947 -1146
rect 3003 -1157 3047 -1146
rect 2751 -1158 3047 -1157
rect 2751 -1210 2764 -1158
rect 2816 -1182 2837 -1158
rect 2889 -1182 2910 -1158
rect 2962 -1182 2982 -1158
rect 3034 -1210 3047 -1158
rect 2751 -1222 2787 -1210
rect 2843 -1222 2867 -1210
rect 2923 -1222 2947 -1210
rect 3003 -1222 3047 -1210
rect 2751 -1274 2764 -1222
rect 2816 -1263 2837 -1238
rect 2889 -1263 2910 -1238
rect 2962 -1263 2982 -1238
rect 3034 -1274 3047 -1222
rect 2751 -1319 2787 -1274
rect 2843 -1319 2867 -1274
rect 2923 -1319 2947 -1274
rect 3003 -1319 3047 -1274
rect 2751 -1344 3047 -1319
rect 2751 -1400 2787 -1344
rect 2843 -1400 2867 -1344
rect 2923 -1400 2947 -1344
rect 3003 -1400 3047 -1344
rect 2751 -1425 3047 -1400
rect 2751 -1481 2787 -1425
rect 2843 -1481 2867 -1425
rect 2923 -1481 2947 -1425
rect 3003 -1481 3047 -1425
rect 2751 -1506 3047 -1481
rect 2751 -1562 2787 -1506
rect 2843 -1562 2867 -1506
rect 2923 -1562 2947 -1506
rect 3003 -1562 3047 -1506
rect 2751 -1575 3047 -1562
rect 2751 -1627 2761 -1575
rect 2813 -1587 2835 -1575
rect 2887 -1587 2909 -1575
rect 2961 -1587 2983 -1575
rect 3035 -1627 3047 -1575
rect 2751 -1639 2787 -1627
rect 2843 -1639 2867 -1627
rect 2923 -1639 2947 -1627
rect 3003 -1639 3047 -1627
rect 2751 -1691 2761 -1639
rect 2813 -1668 2835 -1643
rect 2887 -1668 2909 -1643
rect 2961 -1668 2983 -1643
rect 3035 -1691 3047 -1639
rect 2751 -1724 2787 -1691
rect 2843 -1724 2867 -1691
rect 2923 -1724 2947 -1691
rect 3003 -1724 3047 -1691
rect 2751 -1749 3047 -1724
rect 2751 -1805 2787 -1749
rect 2843 -1805 2867 -1749
rect 2923 -1805 2947 -1749
rect 3003 -1805 3047 -1749
rect 2751 -1830 3047 -1805
rect 2751 -1886 2787 -1830
rect 2843 -1886 2867 -1830
rect 2923 -1886 2947 -1830
rect 3003 -1886 3047 -1830
rect 2751 -1911 3047 -1886
rect 9698 -813 9989 1362
tri 10145 1811 10252 1918 se
rect 10252 1811 10327 1918
tri 10327 1811 10434 1918 nw
tri 10436 1811 10543 1918 se
rect 10543 1811 10859 1918
rect 10145 1809 10325 1811
tri 10325 1809 10327 1811 nw
tri 10434 1809 10436 1811 se
rect 10436 1809 10859 1811
rect 10145 1771 10287 1809
tri 10287 1771 10325 1809 nw
tri 10396 1771 10434 1809 se
rect 10434 1771 10859 1809
rect 10145 588 10273 1771
tri 10273 1757 10287 1771 nw
tri 10382 1757 10396 1771 se
rect 10396 1757 10859 1771
tri 10369 1744 10382 1757 se
rect 10382 1744 10859 1757
rect 10369 827 10859 1744
rect 10369 771 10386 827
rect 10442 771 10466 827
rect 10522 771 10546 827
rect 10602 771 10626 827
rect 10682 771 10706 827
rect 10762 771 10786 827
rect 10842 771 10859 827
rect 10369 740 10859 771
rect 10369 684 10386 740
rect 10442 684 10466 740
rect 10522 684 10546 740
rect 10602 684 10626 740
rect 10682 684 10706 740
rect 10762 684 10786 740
rect 10842 684 10859 740
rect 10369 652 10859 684
rect 10369 596 10386 652
rect 10442 596 10466 652
rect 10522 596 10546 652
rect 10602 596 10626 652
rect 10682 596 10706 652
rect 10762 596 10786 652
rect 10842 596 10859 652
rect 10369 564 10859 596
rect 10369 508 10386 564
rect 10442 508 10466 564
rect 10522 508 10546 564
rect 10602 508 10626 564
rect 10682 508 10706 564
rect 10762 508 10786 564
rect 10842 508 10859 564
rect 10369 476 10859 508
rect 10369 420 10386 476
rect 10442 420 10466 476
rect 10522 420 10546 476
rect 10602 420 10626 476
rect 10682 420 10706 476
rect 10762 420 10786 476
rect 10842 420 10859 476
rect 10369 388 10859 420
rect 10369 332 10386 388
rect 10442 332 10466 388
rect 10522 332 10546 388
rect 10602 332 10626 388
rect 10682 332 10706 388
rect 10762 332 10786 388
rect 10842 332 10859 388
rect 10369 300 10859 332
rect 10369 244 10386 300
rect 10442 244 10466 300
rect 10522 244 10546 300
rect 10602 244 10626 300
rect 10682 244 10706 300
rect 10762 244 10786 300
rect 10842 244 10859 300
tri 10967 3730 11226 3989 se
rect 11226 3730 12069 3989
rect 10967 291 12069 3730
rect 12177 3190 12669 4117
rect 12177 2494 12194 3190
rect 12650 2494 12669 3190
rect 12177 2469 12669 2494
rect 12177 2413 12194 2469
rect 12250 2413 12274 2469
rect 12330 2413 12354 2469
rect 12410 2413 12434 2469
rect 12490 2413 12514 2469
rect 12570 2413 12594 2469
rect 12650 2413 12669 2469
rect 12177 2388 12669 2413
rect 12177 2332 12194 2388
rect 12250 2332 12274 2388
rect 12330 2332 12354 2388
rect 12410 2332 12434 2388
rect 12490 2332 12514 2388
rect 12570 2332 12594 2388
rect 12650 2332 12669 2388
rect 12177 2307 12669 2332
rect 12177 2251 12194 2307
rect 12250 2251 12274 2307
rect 12330 2251 12354 2307
rect 12410 2251 12434 2307
rect 12490 2251 12514 2307
rect 12570 2251 12594 2307
rect 12650 2251 12669 2307
rect 12177 2226 12669 2251
rect 12177 2170 12194 2226
rect 12250 2170 12274 2226
rect 12330 2170 12354 2226
rect 12410 2170 12434 2226
rect 12490 2170 12514 2226
rect 12570 2170 12594 2226
rect 12650 2170 12669 2226
rect 12177 2145 12669 2170
rect 12177 2089 12194 2145
rect 12250 2089 12274 2145
rect 12330 2089 12354 2145
rect 12410 2089 12434 2145
rect 12490 2089 12514 2145
rect 12570 2089 12594 2145
rect 12650 2089 12669 2145
rect 12177 2064 12669 2089
rect 12177 2008 12194 2064
rect 12250 2008 12274 2064
rect 12330 2008 12354 2064
rect 12410 2008 12434 2064
rect 12490 2008 12514 2064
rect 12570 2008 12594 2064
rect 12650 2008 12669 2064
rect 12177 1983 12669 2008
rect 12177 1927 12194 1983
rect 12250 1927 12274 1983
rect 12330 1927 12354 1983
rect 12410 1927 12434 1983
rect 12490 1927 12514 1983
rect 12570 1927 12594 1983
rect 12650 1927 12669 1983
rect 12177 1902 12669 1927
rect 12177 1846 12194 1902
rect 12250 1846 12274 1902
rect 12330 1846 12354 1902
rect 12410 1846 12434 1902
rect 12490 1846 12514 1902
rect 12570 1846 12594 1902
rect 12650 1846 12669 1902
rect 12177 1821 12669 1846
rect 12177 1765 12194 1821
rect 12250 1765 12274 1821
rect 12330 1765 12354 1821
rect 12410 1765 12434 1821
rect 12490 1765 12514 1821
rect 12570 1765 12594 1821
rect 12650 1765 12669 1821
rect 12177 1740 12669 1765
rect 12177 1684 12194 1740
rect 12250 1684 12274 1740
rect 12330 1684 12354 1740
rect 12410 1684 12434 1740
rect 12490 1684 12514 1740
rect 12570 1684 12594 1740
rect 12650 1684 12669 1740
rect 12177 1659 12669 1684
rect 12177 1603 12194 1659
rect 12250 1603 12274 1659
rect 12330 1603 12354 1659
rect 12410 1603 12434 1659
rect 12490 1603 12514 1659
rect 12570 1603 12594 1659
rect 12650 1603 12669 1659
rect 12177 1578 12669 1603
rect 12177 1522 12194 1578
rect 12250 1522 12274 1578
rect 12330 1522 12354 1578
rect 12410 1522 12434 1578
rect 12490 1522 12514 1578
rect 12570 1522 12594 1578
rect 12650 1522 12669 1578
rect 12177 1497 12669 1522
rect 12177 1441 12194 1497
rect 12250 1441 12274 1497
rect 12330 1441 12354 1497
rect 12410 1441 12434 1497
rect 12490 1441 12514 1497
rect 12570 1441 12594 1497
rect 12650 1441 12669 1497
rect 12177 1416 12669 1441
rect 12177 1360 12194 1416
rect 12250 1360 12274 1416
rect 12330 1360 12354 1416
rect 12410 1360 12434 1416
rect 12490 1360 12514 1416
rect 12570 1360 12594 1416
rect 12650 1360 12669 1416
rect 12177 1346 12669 1360
rect 10369 228 10859 244
rect 2751 -1967 2787 -1911
rect 2843 -1967 2867 -1911
rect 2923 -1967 2947 -1911
rect 3003 -1967 3047 -1911
tri 7489 -1930 7515 -1904 sw
rect 2751 -2191 3047 -1967
tri 7498 -2030 7546 -1982 ne
rect 2751 -2243 2763 -2191
rect 2815 -2243 2837 -2191
rect 2889 -2243 2910 -2191
rect 2962 -2243 2983 -2191
rect 3035 -2243 3047 -2191
rect 2751 -2255 3047 -2243
rect 2751 -2307 2763 -2255
rect 2815 -2307 2837 -2255
rect 2889 -2307 2910 -2255
rect 2962 -2307 2983 -2255
rect 3035 -2307 3047 -2255
rect 2751 -2355 3047 -2307
rect 9698 -2187 9817 -813
tri 9817 -985 9989 -813 nw
rect 12725 -1242 13269 4117
rect 13297 4100 13886 4117
rect 13297 4044 13307 4100
rect 13363 4044 13392 4100
rect 13448 4044 13476 4100
rect 13532 4044 13560 4100
rect 13616 4044 13644 4100
rect 13700 4044 13728 4100
rect 13784 4044 13812 4100
rect 13868 4044 13886 4100
rect 13297 4020 13886 4044
rect 13297 3964 13307 4020
rect 13363 3964 13392 4020
rect 13448 3964 13476 4020
rect 13532 3964 13560 4020
rect 13616 3964 13644 4020
rect 13700 3964 13728 4020
rect 13784 3964 13812 4020
rect 13868 3964 13886 4020
rect 13297 3940 13886 3964
rect 13297 3884 13307 3940
rect 13363 3884 13392 3940
rect 13448 3884 13476 3940
rect 13532 3884 13560 3940
rect 13616 3884 13644 3940
rect 13700 3884 13728 3940
rect 13784 3884 13812 3940
rect 13868 3884 13886 3940
rect 13297 3860 13886 3884
rect 13297 3804 13307 3860
rect 13363 3804 13392 3860
rect 13448 3804 13476 3860
rect 13532 3804 13560 3860
rect 13616 3804 13644 3860
rect 13700 3804 13728 3860
rect 13784 3804 13812 3860
rect 13868 3804 13886 3860
rect 13297 3780 13886 3804
rect 13297 3724 13307 3780
rect 13363 3724 13392 3780
rect 13448 3724 13476 3780
rect 13532 3724 13560 3780
rect 13616 3724 13644 3780
rect 13700 3724 13728 3780
rect 13784 3724 13812 3780
rect 13868 3724 13886 3780
rect 13297 832 13886 3724
tri 14710 3712 14941 3943 se
rect 14941 3712 15794 4464
tri 14709 3711 14710 3712 se
rect 14710 3711 15794 3712
tri 14659 3661 14709 3711 se
rect 14709 3661 15794 3711
tri 14607 3609 14659 3661 se
rect 14659 3609 15794 3661
tri 14573 3575 14607 3609 se
rect 14607 3575 15794 3609
tri 14521 3523 14573 3575 se
rect 14573 3523 15794 3575
tri 14488 3490 14521 3523 se
rect 14521 3490 15794 3523
tri 14436 3438 14488 3490 se
rect 14488 3438 15794 3490
tri 14423 3425 14436 3438 se
rect 14436 3425 15794 3438
tri 14414 3416 14423 3425 se
rect 14423 3416 15794 3425
tri 14408 3410 14414 3416 se
rect 14414 3410 15794 3416
tri 14197 3199 14408 3410 se
rect 14408 3386 15794 3410
rect 14408 3199 15592 3386
tri 14182 3184 14197 3199 se
rect 14197 3184 15592 3199
tri 15592 3184 15794 3386 nw
rect 13942 3162 15570 3184
tri 15570 3162 15592 3184 nw
rect 13942 3159 15561 3162
rect 13942 3103 13972 3159
rect 14028 3103 14063 3159
rect 14119 3103 14154 3159
rect 14210 3103 14244 3159
rect 14300 3103 14334 3159
rect 14390 3103 14424 3159
rect 14480 3103 14514 3159
rect 14570 3153 15561 3159
tri 15561 3153 15570 3162 nw
rect 14570 3145 15249 3153
rect 14570 3103 14630 3145
rect 13942 3089 14630 3103
rect 14686 3089 14718 3145
rect 14774 3089 14806 3145
rect 14862 3089 14894 3145
rect 14950 3089 14982 3145
rect 15038 3089 15070 3145
rect 15126 3089 15158 3145
rect 15214 3089 15249 3145
rect 13942 3079 15249 3089
rect 13942 3023 13972 3079
rect 14028 3023 14063 3079
rect 14119 3023 14154 3079
rect 14210 3023 14244 3079
rect 14300 3023 14334 3079
rect 14390 3023 14424 3079
rect 14480 3023 14514 3079
rect 14570 3065 15249 3079
rect 14570 3023 14630 3065
rect 13942 3009 14630 3023
rect 14686 3009 14718 3065
rect 14774 3009 14806 3065
rect 14862 3009 14894 3065
rect 14950 3009 14982 3065
rect 15038 3009 15070 3065
rect 15126 3009 15158 3065
rect 15214 3009 15249 3065
rect 13942 2999 15249 3009
rect 13942 2943 13972 2999
rect 14028 2943 14063 2999
rect 14119 2943 14154 2999
rect 14210 2943 14244 2999
rect 14300 2943 14334 2999
rect 14390 2943 14424 2999
rect 14480 2943 14514 2999
rect 14570 2985 15249 2999
rect 14570 2943 14630 2985
rect 13942 2929 14630 2943
rect 14686 2929 14718 2985
rect 14774 2929 14806 2985
rect 14862 2929 14894 2985
rect 14950 2929 14982 2985
rect 15038 2929 15070 2985
rect 15126 2929 15158 2985
rect 15214 2929 15249 2985
rect 13942 2919 15249 2929
rect 13942 2863 13972 2919
rect 14028 2863 14063 2919
rect 14119 2863 14154 2919
rect 14210 2863 14244 2919
rect 14300 2863 14334 2919
rect 14390 2863 14424 2919
rect 14480 2863 14514 2919
rect 14570 2905 15249 2919
rect 14570 2863 14630 2905
rect 13942 2849 14630 2863
rect 14686 2849 14718 2905
rect 14774 2849 14806 2905
rect 14862 2849 14894 2905
rect 14950 2849 14982 2905
rect 15038 2849 15070 2905
rect 15126 2849 15158 2905
rect 15214 2849 15249 2905
rect 13942 2841 15249 2849
tri 15249 2841 15561 3153 nw
rect 13942 2839 15206 2841
rect 13942 2783 13972 2839
rect 14028 2783 14063 2839
rect 14119 2783 14154 2839
rect 14210 2783 14244 2839
rect 14300 2783 14334 2839
rect 14390 2783 14424 2839
rect 14480 2783 14514 2839
rect 14570 2798 15206 2839
tri 15206 2798 15249 2841 nw
rect 14570 2789 14907 2798
rect 14570 2783 14641 2789
rect 13942 2759 14641 2783
rect 13942 2703 13972 2759
rect 14028 2703 14063 2759
rect 14119 2703 14154 2759
rect 14210 2703 14244 2759
rect 14300 2703 14334 2759
rect 14390 2703 14424 2759
rect 14480 2703 14514 2759
rect 14570 2733 14641 2759
rect 14697 2733 14721 2789
rect 14777 2733 14801 2789
rect 14857 2733 14907 2789
rect 14570 2703 14907 2733
rect 13942 2679 14907 2703
rect 13942 2623 13972 2679
rect 14028 2623 14063 2679
rect 14119 2623 14154 2679
rect 14210 2623 14244 2679
rect 14300 2623 14334 2679
rect 14390 2623 14424 2679
rect 14480 2623 14514 2679
rect 14570 2677 14907 2679
rect 14570 2623 14641 2677
rect 13942 2621 14641 2623
rect 14697 2621 14721 2677
rect 14777 2621 14801 2677
rect 14857 2621 14907 2677
rect 13942 2599 14907 2621
rect 13942 2543 13972 2599
rect 14028 2543 14063 2599
rect 14119 2543 14154 2599
rect 14210 2543 14244 2599
rect 14300 2543 14334 2599
rect 14390 2543 14424 2599
rect 14480 2543 14514 2599
rect 14570 2564 14907 2599
rect 14570 2543 14641 2564
rect 13942 2519 14641 2543
rect 13942 2463 13972 2519
rect 14028 2463 14063 2519
rect 14119 2463 14154 2519
rect 14210 2463 14244 2519
rect 14300 2463 14334 2519
rect 14390 2463 14424 2519
rect 14480 2463 14514 2519
rect 14570 2508 14641 2519
rect 14697 2508 14721 2564
rect 14777 2508 14801 2564
rect 14857 2508 14907 2564
rect 14570 2499 14907 2508
tri 14907 2499 15206 2798 nw
tri 15832 2764 15853 2785 se
rect 15853 2769 15911 4521
rect 16120 4513 16144 4569
rect 16200 4513 16224 4569
rect 16280 4513 16304 4569
rect 16360 4513 16384 4569
rect 16440 4513 16464 4569
rect 16064 4504 16520 4513
rect 16190 4464 16412 4504
tri 16573 3356 16633 3416 se
rect 16633 3392 16691 4521
rect 16633 3356 16655 3392
tri 16655 3356 16691 3392 nw
tri 16712 3356 16786 3430 se
rect 16786 3414 16844 4522
rect 17012 4464 17332 4529
rect 16786 3402 16832 3414
tri 16832 3402 16844 3414 nw
rect 16786 3368 16798 3402
tri 16798 3368 16832 3402 nw
tri 16838 3368 16872 3402 se
rect 16872 3386 16930 4464
tri 16786 3356 16798 3368 nw
tri 16826 3356 16838 3368 se
rect 16838 3356 16872 3368
tri 16551 3334 16573 3356 se
rect 16573 3335 16634 3356
tri 16634 3335 16655 3356 nw
tri 16691 3335 16712 3356 se
rect 16712 3335 16758 3356
rect 16573 3334 16633 3335
tri 16633 3334 16634 3335 nw
tri 16690 3334 16691 3335 se
rect 16691 3334 16758 3335
tri 16499 3282 16551 3334 se
rect 16551 3282 16581 3334
tri 16581 3282 16633 3334 nw
tri 16638 3282 16690 3334 se
rect 16690 3328 16758 3334
tri 16758 3328 16786 3356 nw
tri 16798 3328 16826 3356 se
rect 16826 3328 16872 3356
tri 16872 3328 16930 3386 nw
rect 16690 3294 16724 3328
tri 16724 3294 16758 3328 nw
tri 16764 3294 16798 3328 se
rect 16690 3282 16712 3294
tri 16712 3282 16724 3294 nw
tri 16752 3282 16764 3294 se
rect 16764 3282 16798 3294
tri 16469 3252 16499 3282 se
rect 16499 3277 16576 3282
tri 16576 3277 16581 3282 nw
tri 16633 3277 16638 3282 se
rect 16638 3277 16684 3282
rect 16499 3252 16551 3277
tri 16551 3252 16576 3277 nw
tri 16608 3252 16633 3277 se
rect 16633 3254 16684 3277
tri 16684 3254 16712 3282 nw
tri 16724 3254 16752 3282 se
rect 16752 3254 16798 3282
tri 16798 3254 16872 3328 nw
rect 16633 3252 16650 3254
tri 16425 3208 16469 3252 se
rect 16469 3208 16507 3252
tri 16507 3208 16551 3252 nw
tri 16564 3208 16608 3252 se
rect 16608 3220 16650 3252
tri 16650 3220 16684 3254 nw
tri 16690 3220 16724 3254 se
rect 16608 3208 16638 3220
tri 16638 3208 16650 3220 nw
tri 16678 3208 16690 3220 se
rect 16690 3208 16724 3220
tri 16401 3184 16425 3208 se
rect 16425 3195 16494 3208
tri 16494 3195 16507 3208 nw
tri 16551 3195 16564 3208 se
rect 16564 3195 16610 3208
rect 16425 3184 16483 3195
tri 16483 3184 16494 3195 nw
tri 16540 3184 16551 3195 se
rect 16551 3184 16610 3195
tri 16387 3170 16401 3184 se
rect 16401 3170 16469 3184
tri 16469 3170 16483 3184 nw
tri 16526 3170 16540 3184 se
rect 16540 3180 16610 3184
tri 16610 3180 16638 3208 nw
tri 16650 3180 16678 3208 se
rect 16678 3180 16724 3208
tri 16724 3180 16798 3254 nw
rect 16540 3170 16576 3180
tri 16379 3162 16387 3170 se
rect 16387 3162 16461 3170
tri 16461 3162 16469 3170 nw
tri 16518 3162 16526 3170 se
rect 16526 3162 16576 3170
tri 16370 3153 16379 3162 se
rect 16379 3153 16452 3162
tri 16452 3153 16461 3162 nw
tri 16509 3153 16518 3162 se
rect 16518 3153 16576 3162
tri 16351 3134 16370 3153 se
rect 16370 3134 16433 3153
tri 16433 3134 16452 3153 nw
tri 16490 3134 16509 3153 se
rect 16509 3146 16576 3153
tri 16576 3146 16610 3180 nw
tri 16616 3146 16650 3180 se
rect 16509 3134 16564 3146
tri 16564 3134 16576 3146 nw
tri 16604 3134 16616 3146 se
rect 16616 3134 16650 3146
tri 16305 3088 16351 3134 se
rect 16351 3113 16412 3134
tri 16412 3113 16433 3134 nw
tri 16469 3113 16490 3134 se
rect 16490 3113 16536 3134
rect 16351 3088 16387 3113
tri 16387 3088 16412 3113 nw
tri 16444 3088 16469 3113 se
rect 16469 3106 16536 3113
tri 16536 3106 16564 3134 nw
tri 16576 3106 16604 3134 se
rect 16604 3106 16650 3134
tri 16650 3106 16724 3180 nw
rect 19429 3173 19911 7903
rect 20833 14803 21151 14827
rect 20833 13307 20888 14803
rect 21104 13307 21151 14803
rect 20833 13282 21151 13307
rect 20833 13226 20888 13282
rect 20944 13226 20968 13282
rect 21024 13226 21048 13282
rect 21104 13226 21151 13282
rect 20833 13201 21151 13226
rect 20833 13145 20888 13201
rect 20944 13145 20968 13201
rect 21024 13145 21048 13201
rect 21104 13145 21151 13201
rect 20833 13120 21151 13145
rect 20833 13064 20888 13120
rect 20944 13064 20968 13120
rect 21024 13064 21048 13120
rect 21104 13064 21151 13120
rect 20833 13039 21151 13064
rect 20833 12983 20888 13039
rect 20944 12983 20968 13039
rect 21024 12983 21048 13039
rect 21104 12983 21151 13039
rect 20833 12958 21151 12983
rect 20833 12902 20888 12958
rect 20944 12902 20968 12958
rect 21024 12902 21048 12958
rect 21104 12902 21151 12958
rect 20833 12877 21151 12902
rect 20833 12821 20888 12877
rect 20944 12821 20968 12877
rect 21024 12821 21048 12877
rect 21104 12821 21151 12877
rect 20833 12796 21151 12821
rect 20833 12740 20888 12796
rect 20944 12740 20968 12796
rect 21024 12740 21048 12796
rect 21104 12740 21151 12796
rect 20833 12715 21151 12740
rect 20833 12659 20888 12715
rect 20944 12659 20968 12715
rect 21024 12659 21048 12715
rect 21104 12659 21151 12715
rect 20833 12634 21151 12659
rect 20833 12578 20888 12634
rect 20944 12578 20968 12634
rect 21024 12578 21048 12634
rect 21104 12578 21151 12634
rect 20833 12553 21151 12578
rect 20833 12497 20888 12553
rect 20944 12497 20968 12553
rect 21024 12497 21048 12553
rect 21104 12497 21151 12553
rect 20833 12472 21151 12497
rect 20833 12416 20888 12472
rect 20944 12416 20968 12472
rect 21024 12416 21048 12472
rect 21104 12416 21151 12472
rect 20833 12391 21151 12416
rect 20833 12335 20888 12391
rect 20944 12335 20968 12391
rect 21024 12335 21048 12391
rect 21104 12335 21151 12391
rect 20833 12310 21151 12335
rect 20833 12254 20888 12310
rect 20944 12254 20968 12310
rect 21024 12254 21048 12310
rect 21104 12254 21151 12310
rect 20833 12229 21151 12254
rect 20833 12173 20888 12229
rect 20944 12173 20968 12229
rect 21024 12173 21048 12229
rect 21104 12173 21151 12229
rect 20833 12148 21151 12173
rect 20833 12092 20888 12148
rect 20944 12092 20968 12148
rect 21024 12092 21048 12148
rect 21104 12092 21151 12148
rect 20833 12067 21151 12092
rect 20833 12011 20888 12067
rect 20944 12011 20968 12067
rect 21024 12011 21048 12067
rect 21104 12011 21151 12067
rect 20833 11986 21151 12011
rect 20833 11930 20888 11986
rect 20944 11930 20968 11986
rect 21024 11930 21048 11986
rect 21104 11930 21151 11986
rect 20833 11905 21151 11930
rect 20833 11849 20888 11905
rect 20944 11849 20968 11905
rect 21024 11849 21048 11905
rect 21104 11849 21151 11905
rect 20833 11824 21151 11849
rect 20833 11768 20888 11824
rect 20944 11768 20968 11824
rect 21024 11768 21048 11824
rect 21104 11768 21151 11824
rect 20833 11743 21151 11768
rect 20833 11687 20888 11743
rect 20944 11687 20968 11743
rect 21024 11687 21048 11743
rect 21104 11687 21151 11743
rect 20833 11662 21151 11687
rect 20833 11606 20888 11662
rect 20944 11606 20968 11662
rect 21024 11606 21048 11662
rect 21104 11606 21151 11662
rect 20833 11581 21151 11606
rect 20833 11525 20888 11581
rect 20944 11525 20968 11581
rect 21024 11525 21048 11581
rect 21104 11525 21151 11581
rect 20833 11500 21151 11525
rect 20833 11444 20888 11500
rect 20944 11444 20968 11500
rect 21024 11444 21048 11500
rect 21104 11444 21151 11500
rect 20833 11419 21151 11444
rect 20833 11363 20888 11419
rect 20944 11363 20968 11419
rect 21024 11363 21048 11419
rect 21104 11363 21151 11419
rect 20833 11338 21151 11363
rect 20833 11282 20888 11338
rect 20944 11282 20968 11338
rect 21024 11282 21048 11338
rect 21104 11282 21151 11338
rect 20833 11257 21151 11282
rect 20833 11201 20888 11257
rect 20944 11201 20968 11257
rect 21024 11201 21048 11257
rect 21104 11201 21151 11257
rect 20833 11176 21151 11201
rect 20833 11120 20888 11176
rect 20944 11120 20968 11176
rect 21024 11120 21048 11176
rect 21104 11120 21151 11176
rect 20833 11095 21151 11120
rect 20833 11039 20888 11095
rect 20944 11039 20968 11095
rect 21024 11039 21048 11095
rect 21104 11039 21151 11095
rect 20833 11014 21151 11039
rect 20833 10958 20888 11014
rect 20944 10958 20968 11014
rect 21024 10958 21048 11014
rect 21104 10958 21151 11014
rect 20833 10933 21151 10958
rect 20833 10877 20888 10933
rect 20944 10877 20968 10933
rect 21024 10877 21048 10933
rect 21104 10877 21151 10933
rect 20833 10852 21151 10877
rect 20833 10796 20888 10852
rect 20944 10796 20968 10852
rect 21024 10796 21048 10852
rect 21104 10796 21151 10852
rect 20833 10771 21151 10796
rect 20833 10715 20888 10771
rect 20944 10715 20968 10771
rect 21024 10715 21048 10771
rect 21104 10715 21151 10771
rect 20833 10690 21151 10715
rect 20833 10634 20888 10690
rect 20944 10634 20968 10690
rect 21024 10634 21048 10690
rect 21104 10634 21151 10690
rect 20833 10609 21151 10634
rect 20833 10553 20888 10609
rect 20944 10553 20968 10609
rect 21024 10553 21048 10609
rect 21104 10553 21151 10609
rect 20833 10528 21151 10553
rect 20833 10472 20888 10528
rect 20944 10472 20968 10528
rect 21024 10472 21048 10528
rect 21104 10472 21151 10528
rect 20833 10447 21151 10472
rect 20833 10391 20888 10447
rect 20944 10391 20968 10447
rect 21024 10391 21048 10447
rect 21104 10391 21151 10447
rect 20833 10366 21151 10391
rect 20833 10310 20888 10366
rect 20944 10310 20968 10366
rect 21024 10310 21048 10366
rect 21104 10310 21151 10366
rect 20833 10285 21151 10310
rect 20833 10229 20888 10285
rect 20944 10229 20968 10285
rect 21024 10229 21048 10285
rect 21104 10229 21151 10285
rect 20833 10204 21151 10229
rect 20833 10148 20888 10204
rect 20944 10148 20968 10204
rect 21024 10148 21048 10204
rect 21104 10148 21151 10204
rect 20833 10123 21151 10148
rect 20833 10067 20888 10123
rect 20944 10067 20968 10123
rect 21024 10067 21048 10123
rect 21104 10067 21151 10123
rect 21538 14801 21963 14827
rect 21538 10185 21641 14801
tri 21538 10106 21617 10185 ne
rect 20833 10042 21151 10067
rect 20833 9986 20888 10042
rect 20944 9986 20968 10042
rect 21024 9986 21048 10042
rect 21104 9986 21151 10042
rect 20833 9961 21151 9986
rect 20833 9905 20888 9961
rect 20944 9905 20968 9961
rect 21024 9905 21048 9961
rect 21104 9905 21151 9961
rect 20833 9880 21151 9905
rect 20833 9824 20888 9880
rect 20944 9824 20968 9880
rect 21024 9824 21048 9880
rect 21104 9824 21151 9880
rect 20833 9799 21151 9824
rect 20833 9743 20888 9799
rect 20944 9743 20968 9799
rect 21024 9743 21048 9799
rect 21104 9743 21151 9799
rect 20833 9718 21151 9743
rect 20833 9662 20888 9718
rect 20944 9662 20968 9718
rect 21024 9662 21048 9718
rect 21104 9662 21151 9718
rect 20833 9637 21151 9662
rect 20833 9581 20888 9637
rect 20944 9581 20968 9637
rect 21024 9581 21048 9637
rect 21104 9581 21151 9637
rect 20833 9556 21151 9581
rect 20833 9500 20888 9556
rect 20944 9500 20968 9556
rect 21024 9500 21048 9556
rect 21104 9500 21151 9556
rect 20833 9475 21151 9500
rect 20833 9419 20888 9475
rect 20944 9419 20968 9475
rect 21024 9419 21048 9475
rect 21104 9419 21151 9475
rect 20833 9394 21151 9419
rect 20833 9338 20888 9394
rect 20944 9338 20968 9394
rect 21024 9338 21048 9394
rect 21104 9338 21151 9394
rect 20833 9313 21151 9338
rect 20833 9257 20888 9313
rect 20944 9257 20968 9313
rect 21024 9257 21048 9313
rect 21104 9257 21151 9313
rect 20833 9232 21151 9257
rect 20833 9176 20888 9232
rect 20944 9176 20968 9232
rect 21024 9176 21048 9232
rect 21104 9176 21151 9232
rect 20833 9151 21151 9176
rect 20833 9095 20888 9151
rect 20944 9095 20968 9151
rect 21024 9095 21048 9151
rect 21104 9095 21151 9151
rect 20833 9070 21151 9095
rect 20833 9014 20888 9070
rect 20944 9014 20968 9070
rect 21024 9014 21048 9070
rect 21104 9014 21151 9070
rect 20833 8989 21151 9014
rect 20833 8933 20888 8989
rect 20944 8933 20968 8989
rect 21024 8933 21048 8989
rect 21104 8933 21151 8989
rect 20833 8908 21151 8933
rect 20833 8852 20888 8908
rect 20944 8852 20968 8908
rect 21024 8852 21048 8908
rect 21104 8852 21151 8908
rect 20833 8827 21151 8852
rect 20833 8771 20888 8827
rect 20944 8771 20968 8827
rect 21024 8771 21048 8827
rect 21104 8771 21151 8827
rect 20833 8746 21151 8771
rect 20833 8690 20888 8746
rect 20944 8690 20968 8746
rect 21024 8690 21048 8746
rect 21104 8690 21151 8746
rect 20833 8665 21151 8690
rect 20833 8609 20888 8665
rect 20944 8609 20968 8665
rect 21024 8609 21048 8665
rect 21104 8609 21151 8665
rect 20833 8584 21151 8609
rect 20833 8528 20888 8584
rect 20944 8528 20968 8584
rect 21024 8528 21048 8584
rect 21104 8528 21151 8584
rect 20833 8503 21151 8528
rect 20833 8447 20888 8503
rect 20944 8447 20968 8503
rect 21024 8447 21048 8503
rect 21104 8447 21151 8503
rect 20833 8422 21151 8447
rect 20833 8366 20888 8422
rect 20944 8366 20968 8422
rect 21024 8366 21048 8422
rect 21104 8366 21151 8422
rect 20833 8341 21151 8366
rect 20833 8285 20888 8341
rect 20944 8285 20968 8341
rect 21024 8285 21048 8341
rect 21104 8285 21151 8341
rect 20833 8260 21151 8285
rect 20833 8204 20888 8260
rect 20944 8204 20968 8260
rect 21024 8204 21048 8260
rect 21104 8204 21151 8260
rect 20833 8179 21151 8204
rect 20833 8123 20888 8179
rect 20944 8123 20968 8179
rect 21024 8123 21048 8179
rect 21104 8123 21151 8179
rect 20833 8098 21151 8123
rect 20833 8083 20888 8098
rect 20944 8083 20968 8098
rect 21024 8083 21048 8098
rect 21104 8083 21151 8098
rect 20833 8031 20844 8083
rect 20896 8031 20926 8042
rect 20978 8031 21008 8042
rect 21060 8031 21090 8042
rect 21142 8031 21151 8083
rect 20833 8019 21151 8031
rect 20833 7967 20844 8019
rect 20896 8017 20926 8019
rect 20978 8017 21008 8019
rect 21060 8017 21090 8019
rect 21142 7967 21151 8019
rect 20833 7961 20888 7967
rect 20944 7961 20968 7967
rect 21024 7961 21048 7967
rect 21104 7961 21151 7967
rect 20833 7955 21151 7961
rect 20833 7903 20844 7955
rect 20896 7936 20926 7955
rect 20978 7936 21008 7955
rect 21060 7936 21090 7955
rect 21142 7903 21151 7955
rect 20833 7880 20888 7903
rect 20944 7880 20968 7903
rect 21024 7880 21048 7903
rect 21104 7880 21151 7903
tri 19911 3173 19942 3204 sw
rect 19429 3121 19942 3173
tri 19942 3121 19994 3173 sw
rect 16469 3088 16502 3106
tri 16277 3060 16305 3088 se
rect 16305 3060 16359 3088
tri 16359 3060 16387 3088 nw
tri 16416 3060 16444 3088 se
rect 16444 3072 16502 3088
tri 16502 3072 16536 3106 nw
tri 16542 3072 16576 3106 se
rect 16444 3060 16490 3072
tri 16490 3060 16502 3072 nw
tri 16530 3060 16542 3072 se
rect 16542 3060 16576 3072
tri 16223 3006 16277 3060 se
rect 16277 3031 16330 3060
tri 16330 3031 16359 3060 nw
tri 16387 3031 16416 3060 se
rect 16416 3032 16462 3060
tri 16462 3032 16490 3060 nw
tri 16502 3032 16530 3060 se
rect 16530 3032 16576 3060
tri 16576 3032 16650 3106 nw
rect 19429 3091 19994 3121
tri 19994 3091 20024 3121 sw
rect 16416 3031 16428 3032
rect 16277 3006 16305 3031
tri 16305 3006 16330 3031 nw
tri 16362 3006 16387 3031 se
rect 16387 3006 16428 3031
tri 16203 2986 16223 3006 se
rect 16223 2986 16285 3006
tri 16285 2986 16305 3006 nw
tri 16342 2986 16362 3006 se
rect 16362 2998 16428 3006
tri 16428 2998 16462 3032 nw
tri 16468 2998 16502 3032 se
rect 16362 2986 16416 2998
tri 16416 2986 16428 2998 nw
tri 16456 2986 16468 2998 se
rect 16468 2986 16502 2998
tri 16141 2924 16203 2986 se
rect 16203 2949 16248 2986
tri 16248 2949 16285 2986 nw
tri 16305 2949 16342 2986 se
rect 16342 2958 16388 2986
tri 16388 2958 16416 2986 nw
tri 16428 2958 16456 2986 se
rect 16456 2958 16502 2986
tri 16502 2958 16576 3032 nw
rect 16342 2949 16354 2958
rect 16203 2924 16223 2949
tri 16223 2924 16248 2949 nw
tri 16280 2924 16305 2949 se
rect 16305 2924 16354 2949
tri 16354 2924 16388 2958 nw
tri 16394 2924 16428 2958 se
tri 16129 2912 16141 2924 se
rect 16141 2912 16211 2924
tri 16211 2912 16223 2924 nw
tri 16268 2912 16280 2924 se
rect 16280 2912 16342 2924
tri 16342 2912 16354 2924 nw
tri 16382 2912 16394 2924 se
rect 16394 2912 16428 2924
tri 16059 2842 16129 2912 se
rect 16129 2867 16166 2912
tri 16166 2867 16211 2912 nw
tri 16223 2867 16268 2912 se
rect 16268 2884 16314 2912
tri 16314 2884 16342 2912 nw
tri 16354 2884 16382 2912 se
rect 16382 2884 16428 2912
tri 16428 2884 16502 2958 nw
rect 16268 2867 16280 2884
rect 16129 2842 16141 2867
tri 16141 2842 16166 2867 nw
tri 16198 2842 16223 2867 se
rect 16223 2850 16280 2867
tri 16280 2850 16314 2884 nw
tri 16320 2850 16354 2884 se
rect 16223 2842 16268 2850
tri 16058 2841 16059 2842 se
rect 16059 2841 16140 2842
tri 16140 2841 16141 2842 nw
tri 16197 2841 16198 2842 se
rect 16198 2841 16268 2842
tri 16055 2838 16058 2841 se
rect 16058 2838 16137 2841
tri 16137 2838 16140 2841 nw
tri 16194 2838 16197 2841 se
rect 16197 2838 16268 2841
tri 16268 2838 16280 2850 nw
tri 16308 2838 16320 2850 se
rect 16320 2838 16354 2850
tri 16015 2798 16055 2838 se
rect 16055 2798 16097 2838
tri 16097 2798 16137 2838 nw
tri 16154 2798 16194 2838 se
rect 16194 2810 16240 2838
tri 16240 2810 16268 2838 nw
tri 16280 2810 16308 2838 se
rect 16308 2810 16354 2838
tri 16354 2810 16428 2884 nw
rect 16194 2798 16206 2810
rect 15853 2764 15906 2769
tri 15906 2764 15911 2769 nw
tri 15981 2764 16015 2798 se
rect 16015 2785 16084 2798
tri 16084 2785 16097 2798 nw
tri 16141 2785 16154 2798 se
rect 16154 2785 16206 2798
rect 16015 2764 16063 2785
tri 16063 2764 16084 2785 nw
tri 16120 2764 16141 2785 se
rect 16141 2776 16206 2785
tri 16206 2776 16240 2810 nw
tri 16246 2776 16280 2810 se
rect 16141 2764 16194 2776
tri 16194 2764 16206 2776 nw
tri 16234 2764 16246 2776 se
rect 16246 2764 16280 2776
tri 15828 2760 15832 2764 se
rect 15832 2760 15902 2764
tri 15902 2760 15906 2764 nw
tri 15977 2760 15981 2764 se
rect 15981 2760 16059 2764
tri 16059 2760 16063 2764 nw
tri 16116 2760 16120 2764 se
rect 16120 2760 16190 2764
tri 16190 2760 16194 2764 nw
tri 16230 2760 16234 2764 se
rect 16234 2760 16280 2764
tri 15779 2711 15828 2760 se
rect 15828 2711 15853 2760
tri 15853 2711 15902 2760 nw
tri 15928 2711 15977 2760 se
rect 15977 2711 16002 2760
tri 15758 2690 15779 2711 se
rect 15779 2690 15832 2711
tri 15832 2690 15853 2711 nw
tri 15907 2690 15928 2711 se
rect 15928 2703 16002 2711
tri 16002 2703 16059 2760 nw
tri 16059 2703 16116 2760 se
rect 16116 2736 16166 2760
tri 16166 2736 16190 2760 nw
tri 16206 2736 16230 2760 se
rect 16230 2736 16280 2760
tri 16280 2736 16354 2810 nw
rect 19429 2805 20024 3091
tri 20024 2805 20310 3091 sw
rect 16116 2703 16132 2736
rect 15928 2690 15989 2703
tri 15989 2690 16002 2703 nw
tri 16046 2690 16059 2703 se
rect 16059 2702 16132 2703
tri 16132 2702 16166 2736 nw
tri 16172 2702 16206 2736 se
rect 16059 2690 16120 2702
tri 16120 2690 16132 2702 nw
tri 16160 2690 16172 2702 se
rect 16172 2690 16206 2702
tri 15746 2678 15758 2690 se
rect 15758 2678 15820 2690
tri 15820 2678 15832 2690 nw
tri 15895 2678 15907 2690 se
rect 15907 2678 15977 2690
tri 15977 2678 15989 2690 nw
tri 16034 2678 16046 2690 se
rect 16046 2678 16108 2690
tri 16108 2678 16120 2690 nw
tri 16148 2678 16160 2690 se
rect 16160 2678 16206 2690
tri 15705 2637 15746 2678 se
rect 15746 2637 15779 2678
tri 15779 2637 15820 2678 nw
tri 15854 2637 15895 2678 se
rect 15895 2637 15920 2678
tri 15684 2616 15705 2637 se
rect 15705 2616 15758 2637
tri 15758 2616 15779 2637 nw
tri 15833 2616 15854 2637 se
rect 15854 2621 15920 2637
tri 15920 2621 15977 2678 nw
tri 15977 2621 16034 2678 se
rect 16034 2662 16092 2678
tri 16092 2662 16108 2678 nw
tri 16132 2662 16148 2678 se
rect 16148 2662 16206 2678
tri 16206 2662 16280 2736 nw
rect 16034 2628 16058 2662
tri 16058 2628 16092 2662 nw
tri 16098 2628 16132 2662 se
rect 16034 2621 16046 2628
rect 15854 2616 15915 2621
tri 15915 2616 15920 2621 nw
tri 15972 2616 15977 2621 se
rect 15977 2616 16046 2621
tri 16046 2616 16058 2628 nw
tri 16086 2616 16098 2628 se
rect 16098 2616 16132 2628
tri 15664 2596 15684 2616 se
rect 15684 2596 15738 2616
tri 15738 2596 15758 2616 nw
tri 15813 2596 15833 2616 se
rect 15833 2596 15895 2616
tri 15895 2596 15915 2616 nw
tri 15952 2596 15972 2616 se
rect 15972 2596 16026 2616
tri 16026 2596 16046 2616 nw
tri 16066 2596 16086 2616 se
rect 16086 2596 16132 2616
tri 15631 2563 15664 2596 se
rect 15664 2563 15705 2596
tri 15705 2563 15738 2596 nw
tri 15780 2563 15813 2596 se
rect 15813 2563 15841 2596
tri 15610 2542 15631 2563 se
rect 15631 2542 15684 2563
tri 15684 2542 15705 2563 nw
tri 15759 2542 15780 2563 se
rect 15780 2542 15841 2563
tri 15841 2542 15895 2596 nw
tri 15898 2542 15952 2596 se
rect 15952 2588 16018 2596
tri 16018 2588 16026 2596 nw
tri 16058 2588 16066 2596 se
rect 16066 2588 16132 2596
tri 16132 2588 16206 2662 nw
rect 15952 2554 15984 2588
tri 15984 2554 16018 2588 nw
tri 16024 2554 16058 2588 se
rect 15952 2542 15972 2554
tri 15972 2542 15984 2554 nw
tri 16012 2542 16024 2554 se
rect 16024 2542 16058 2554
tri 15582 2514 15610 2542 se
rect 15610 2514 15656 2542
tri 15656 2514 15684 2542 nw
tri 15731 2514 15759 2542 se
rect 15759 2539 15838 2542
tri 15838 2539 15841 2542 nw
tri 15895 2539 15898 2542 se
rect 15898 2539 15944 2542
rect 15759 2514 15813 2539
tri 15813 2514 15838 2539 nw
tri 15870 2514 15895 2539 se
rect 15895 2514 15944 2539
tri 15944 2514 15972 2542 nw
tri 15984 2514 16012 2542 se
rect 16012 2514 16058 2542
tri 16058 2514 16132 2588 nw
tri 15567 2499 15582 2514 se
rect 15582 2499 15641 2514
tri 15641 2499 15656 2514 nw
tri 15716 2499 15731 2514 se
rect 15731 2499 15798 2514
tri 15798 2499 15813 2514 nw
tri 15855 2499 15870 2514 se
rect 15870 2499 15910 2514
rect 14570 2463 14628 2499
rect 13942 2439 14628 2463
rect 13942 2383 13972 2439
rect 14028 2383 14063 2439
rect 14119 2383 14154 2439
rect 14210 2383 14244 2439
rect 14300 2383 14334 2439
rect 14390 2383 14424 2439
rect 14480 2383 14514 2439
rect 14570 2383 14628 2439
rect 13942 2359 14628 2383
rect 13942 2303 13972 2359
rect 14028 2303 14063 2359
rect 14119 2303 14154 2359
rect 14210 2303 14244 2359
rect 14300 2303 14334 2359
rect 14390 2303 14424 2359
rect 14480 2303 14514 2359
rect 14570 2303 14628 2359
rect 13942 2279 14628 2303
rect 13942 2223 13972 2279
rect 14028 2223 14063 2279
rect 14119 2223 14154 2279
rect 14210 2223 14244 2279
rect 14300 2223 14334 2279
rect 14390 2223 14424 2279
rect 14480 2223 14514 2279
rect 14570 2223 14628 2279
rect 13942 2220 14628 2223
tri 14628 2220 14907 2499 nw
tri 15557 2489 15567 2499 se
rect 15567 2489 15631 2499
tri 15631 2489 15641 2499 nw
tri 15706 2489 15716 2499 se
rect 15716 2489 15767 2499
tri 15536 2468 15557 2489 se
rect 15557 2468 15610 2489
tri 15610 2468 15631 2489 nw
tri 15685 2468 15706 2489 se
rect 15706 2468 15767 2489
tri 15767 2468 15798 2499 nw
tri 15824 2468 15855 2499 se
rect 15855 2480 15910 2499
tri 15910 2480 15944 2514 nw
tri 15950 2480 15984 2514 se
rect 15855 2468 15898 2480
tri 15898 2468 15910 2480 nw
tri 15938 2468 15950 2480 se
rect 15950 2468 15984 2480
tri 15500 2432 15536 2468 se
rect 15536 2432 15574 2468
tri 15574 2432 15610 2468 nw
tri 15649 2432 15685 2468 se
rect 15685 2457 15756 2468
tri 15756 2457 15767 2468 nw
tri 15813 2457 15824 2468 se
rect 15824 2457 15870 2468
rect 15685 2432 15731 2457
tri 15731 2432 15756 2457 nw
tri 15788 2432 15813 2457 se
rect 15813 2440 15870 2457
tri 15870 2440 15898 2468 nw
tri 15910 2440 15938 2468 se
rect 15938 2440 15984 2468
tri 15984 2440 16058 2514 nw
rect 15813 2432 15836 2440
tri 15483 2415 15500 2432 se
rect 15500 2415 15557 2432
tri 15557 2415 15574 2432 nw
tri 15632 2415 15649 2432 se
rect 15649 2415 15693 2432
tri 15462 2394 15483 2415 se
rect 15483 2394 15536 2415
tri 15536 2394 15557 2415 nw
tri 15611 2394 15632 2415 se
rect 15632 2394 15693 2415
tri 15693 2394 15731 2432 nw
tri 15750 2394 15788 2432 se
rect 15788 2406 15836 2432
tri 15836 2406 15870 2440 nw
tri 15876 2406 15910 2440 se
rect 15788 2394 15824 2406
tri 15824 2394 15836 2406 nw
tri 15864 2394 15876 2406 se
rect 15876 2394 15910 2406
tri 15418 2350 15462 2394 se
rect 15462 2350 15492 2394
tri 15492 2350 15536 2394 nw
tri 15567 2350 15611 2394 se
rect 15611 2375 15674 2394
tri 15674 2375 15693 2394 nw
tri 15731 2375 15750 2394 se
rect 15750 2375 15796 2394
rect 15611 2350 15649 2375
tri 15649 2350 15674 2375 nw
tri 15706 2350 15731 2375 se
rect 15731 2366 15796 2375
tri 15796 2366 15824 2394 nw
tri 15836 2366 15864 2394 se
rect 15864 2366 15910 2394
tri 15910 2366 15984 2440 nw
rect 15731 2350 15762 2366
tri 15409 2341 15418 2350 se
rect 15418 2341 15483 2350
tri 15483 2341 15492 2350 nw
tri 15558 2341 15567 2350 se
rect 15567 2341 15619 2350
tri 15388 2320 15409 2341 se
rect 15409 2320 15462 2341
tri 15462 2320 15483 2341 nw
tri 15537 2320 15558 2341 se
rect 15558 2320 15619 2341
tri 15619 2320 15649 2350 nw
tri 15676 2320 15706 2350 se
rect 15706 2332 15762 2350
tri 15762 2332 15796 2366 nw
tri 15802 2332 15836 2366 se
rect 15706 2320 15750 2332
tri 15750 2320 15762 2332 nw
tri 15790 2320 15802 2332 se
rect 15802 2320 15836 2332
tri 15336 2268 15388 2320 se
rect 15388 2268 15410 2320
tri 15410 2268 15462 2320 nw
tri 15485 2268 15537 2320 se
rect 15537 2293 15592 2320
tri 15592 2293 15619 2320 nw
tri 15649 2293 15676 2320 se
rect 15676 2293 15722 2320
rect 15537 2268 15567 2293
tri 15567 2268 15592 2293 nw
tri 15624 2268 15649 2293 se
rect 15649 2292 15722 2293
tri 15722 2292 15750 2320 nw
tri 15762 2292 15790 2320 se
rect 15790 2292 15836 2320
tri 15836 2292 15910 2366 nw
rect 15649 2268 15688 2292
tri 15335 2267 15336 2268 se
rect 15336 2267 15409 2268
tri 15409 2267 15410 2268 nw
tri 15484 2267 15485 2268 se
rect 15485 2267 15545 2268
tri 15314 2246 15335 2267 se
rect 15335 2246 15388 2267
tri 15388 2246 15409 2267 nw
tri 15463 2246 15484 2267 se
rect 15484 2246 15545 2267
tri 15545 2246 15567 2268 nw
tri 15602 2246 15624 2268 se
rect 15624 2258 15688 2268
tri 15688 2258 15722 2292 nw
tri 15728 2258 15762 2292 se
rect 15624 2246 15676 2258
tri 15676 2246 15688 2258 nw
tri 15716 2246 15728 2258 se
rect 15728 2246 15762 2258
tri 15288 2220 15314 2246 se
rect 15314 2220 15362 2246
tri 15362 2220 15388 2246 nw
tri 15437 2220 15463 2246 se
rect 15463 2220 15519 2246
tri 15519 2220 15545 2246 nw
tri 15576 2220 15602 2246 se
rect 15602 2220 15648 2246
rect 13942 2186 14594 2220
tri 14594 2186 14628 2220 nw
tri 15261 2193 15288 2220 se
rect 15288 2193 15335 2220
tri 15335 2193 15362 2220 nw
tri 15410 2193 15437 2220 se
rect 15437 2211 15510 2220
tri 15510 2211 15519 2220 nw
tri 15567 2211 15576 2220 se
rect 15576 2218 15648 2220
tri 15648 2218 15676 2246 nw
tri 15688 2218 15716 2246 se
rect 15716 2218 15762 2246
tri 15762 2218 15836 2292 nw
rect 15576 2211 15614 2218
rect 15437 2193 15485 2211
tri 15254 2186 15261 2193 se
rect 15261 2186 15328 2193
tri 15328 2186 15335 2193 nw
tri 15403 2186 15410 2193 se
rect 15410 2186 15485 2193
tri 15485 2186 15510 2211 nw
tri 15542 2186 15567 2211 se
rect 15567 2186 15614 2211
tri 15240 2172 15254 2186 se
rect 15254 2172 15314 2186
tri 15314 2172 15328 2186 nw
tri 15389 2172 15403 2186 se
rect 15403 2172 15471 2186
tri 15471 2172 15485 2186 nw
tri 15528 2172 15542 2186 se
rect 15542 2184 15614 2186
tri 15614 2184 15648 2218 nw
tri 15654 2184 15688 2218 se
rect 15542 2172 15602 2184
tri 15602 2172 15614 2184 nw
tri 15642 2172 15654 2184 se
rect 15654 2172 15688 2184
tri 15187 2119 15240 2172 se
rect 15240 2119 15261 2172
tri 15261 2119 15314 2172 nw
tri 15336 2119 15389 2172 se
rect 15389 2129 15428 2172
tri 15428 2129 15471 2172 nw
tri 15485 2129 15528 2172 se
rect 15528 2144 15574 2172
tri 15574 2144 15602 2172 nw
tri 15614 2144 15642 2172 se
rect 15642 2144 15688 2172
tri 15688 2144 15762 2218 nw
rect 15528 2129 15540 2144
rect 15389 2119 15403 2129
tri 15172 2104 15187 2119 se
rect 15187 2104 15246 2119
tri 15246 2104 15261 2119 nw
tri 15321 2104 15336 2119 se
rect 15336 2104 15403 2119
tri 15403 2104 15428 2129 nw
tri 15460 2104 15485 2129 se
rect 15485 2110 15540 2129
tri 15540 2110 15574 2144 nw
tri 15580 2110 15614 2144 se
rect 15485 2104 15528 2110
tri 15166 2098 15172 2104 se
rect 15172 2098 15240 2104
tri 15240 2098 15246 2104 nw
tri 15315 2098 15321 2104 se
rect 15321 2098 15397 2104
tri 15397 2098 15403 2104 nw
tri 15454 2098 15460 2104 se
rect 15460 2098 15528 2104
tri 15528 2098 15540 2110 nw
tri 15568 2098 15580 2110 se
rect 15580 2098 15614 2110
tri 15113 2045 15166 2098 se
rect 15166 2045 15187 2098
tri 15187 2045 15240 2098 nw
tri 15262 2045 15315 2098 se
rect 15315 2047 15346 2098
tri 15346 2047 15397 2098 nw
tri 15403 2047 15454 2098 se
rect 15454 2070 15500 2098
tri 15500 2070 15528 2098 nw
tri 15540 2070 15568 2098 se
rect 15568 2070 15614 2098
tri 15614 2070 15688 2144 nw
rect 15454 2047 15466 2070
rect 15315 2045 15323 2047
tri 15092 2024 15113 2045 se
rect 15113 2024 15166 2045
tri 15166 2024 15187 2045 nw
tri 15241 2024 15262 2045 se
rect 15262 2024 15323 2045
tri 15323 2024 15346 2047 nw
tri 15380 2024 15403 2047 se
rect 15403 2036 15466 2047
tri 15466 2036 15500 2070 nw
tri 15506 2036 15540 2070 se
rect 15403 2024 15454 2036
tri 15454 2024 15466 2036 nw
tri 15494 2024 15506 2036 se
rect 15506 2024 15540 2036
tri 15090 2022 15092 2024 se
rect 15092 2022 15164 2024
tri 15164 2022 15166 2024 nw
tri 15239 2022 15241 2024 se
rect 15241 2022 15321 2024
tri 15321 2022 15323 2024 nw
tri 15378 2022 15380 2024 se
rect 15380 2022 15452 2024
tri 15452 2022 15454 2024 nw
tri 15492 2022 15494 2024 se
rect 15494 2022 15540 2024
tri 15047 1979 15090 2022 se
rect 15090 1979 15121 2022
tri 15121 1979 15164 2022 nw
tri 15196 1979 15239 2022 se
rect 15239 1979 15264 2022
tri 14103 1950 14132 1979 se
rect 14132 1950 15092 1979
tri 15092 1950 15121 1979 nw
tri 15167 1950 15196 1979 se
rect 15196 1965 15264 1979
tri 15264 1965 15321 2022 nw
tri 15321 1965 15378 2022 se
rect 15378 1996 15426 2022
tri 15426 1996 15452 2022 nw
tri 15466 1996 15492 2022 se
rect 15492 1996 15540 2022
tri 15540 1996 15614 2070 nw
rect 15378 1965 15392 1996
rect 15196 1950 15249 1965
tri 15249 1950 15264 1965 nw
tri 15306 1950 15321 1965 se
rect 15321 1962 15392 1965
tri 15392 1962 15426 1996 nw
tri 15432 1962 15466 1996 se
rect 15321 1950 15380 1962
tri 15380 1950 15392 1962 nw
tri 15420 1950 15432 1962 se
rect 15432 1950 15466 1962
tri 14093 1940 14103 1950 se
rect 14103 1940 15082 1950
tri 15082 1940 15092 1950 nw
tri 15157 1940 15167 1950 se
rect 15167 1940 15239 1950
tri 15239 1940 15249 1950 nw
tri 15296 1940 15306 1950 se
rect 15306 1940 15352 1950
tri 14066 1913 14093 1940 se
rect 14093 1927 15069 1940
tri 15069 1927 15082 1940 nw
tri 15144 1927 15157 1940 se
rect 15157 1927 15212 1940
rect 14093 1913 14140 1927
tri 14140 1913 14154 1927 nw
tri 15130 1913 15144 1927 se
rect 15144 1913 15212 1927
tri 15212 1913 15239 1940 nw
tri 15269 1913 15296 1940 se
rect 15296 1922 15352 1940
tri 15352 1922 15380 1950 nw
tri 15392 1922 15420 1950 se
rect 15420 1922 15466 1950
tri 15466 1922 15540 1996 nw
rect 15296 1913 15343 1922
tri 15343 1913 15352 1922 nw
tri 15383 1913 15392 1922 se
rect 15392 1913 15457 1922
tri 15457 1913 15466 1922 nw
tri 14058 1905 14066 1913 se
rect 14066 1905 14132 1913
tri 14132 1905 14140 1913 nw
tri 15122 1905 15130 1913 se
rect 15130 1905 15203 1913
tri 14057 1904 14058 1905 se
rect 14058 1904 14131 1905
tri 14131 1904 14132 1905 nw
tri 15121 1904 15122 1905 se
rect 15122 1904 15203 1905
tri 15203 1904 15212 1913 nw
tri 15260 1904 15269 1913 se
rect 15269 1904 15334 1913
tri 15334 1904 15343 1913 nw
tri 15374 1904 15383 1913 se
rect 15383 1904 15448 1913
tri 15448 1904 15457 1913 nw
tri 15612 1904 15621 1913 se
rect 15621 1904 15984 1913
tri 14047 1894 14057 1904 se
rect 14057 1894 14121 1904
tri 14121 1894 14131 1904 nw
tri 15111 1894 15121 1904 se
rect 15121 1894 15193 1904
tri 15193 1894 15203 1904 nw
tri 15250 1894 15260 1904 se
rect 15260 1894 15318 1904
tri 14029 1876 14047 1894 se
rect 14047 1876 14103 1894
tri 14103 1876 14121 1894 nw
tri 14159 1876 14177 1894 se
rect 14177 1876 15175 1894
tri 15175 1876 15193 1894 nw
tri 15232 1876 15250 1894 se
rect 15250 1888 15318 1894
tri 15318 1888 15334 1904 nw
tri 15358 1888 15374 1904 se
rect 15374 1888 15420 1904
rect 15250 1876 15306 1888
tri 15306 1876 15318 1888 nw
tri 15346 1876 15358 1888 se
rect 15358 1876 15420 1888
tri 15420 1876 15448 1904 nw
tri 15584 1876 15612 1904 se
rect 15612 1895 15984 1904
rect 15612 1876 15650 1895
tri 13984 1831 14029 1876 se
rect 14029 1849 14076 1876
tri 14076 1849 14103 1876 nw
tri 14132 1849 14159 1876 se
rect 14159 1849 15141 1876
rect 14029 1831 14058 1849
tri 14058 1831 14076 1849 nw
tri 14114 1831 14132 1849 se
rect 14132 1842 15141 1849
tri 15141 1842 15175 1876 nw
tri 15198 1842 15232 1876 se
rect 15232 1848 15278 1876
tri 15278 1848 15306 1876 nw
tri 15318 1848 15346 1876 se
rect 15346 1848 15392 1876
tri 15392 1848 15420 1876 nw
tri 15556 1848 15584 1876 se
rect 15584 1848 15650 1876
rect 15232 1842 15244 1848
rect 14132 1831 14177 1842
tri 13973 1820 13984 1831 se
rect 13984 1820 14047 1831
tri 14047 1820 14058 1831 nw
tri 14103 1820 14114 1831 se
rect 14114 1820 14177 1831
tri 14177 1820 14199 1842 nw
tri 15176 1820 15198 1842 se
rect 15198 1820 15244 1842
tri 13962 1809 13973 1820 se
rect 13973 1809 14036 1820
tri 14036 1809 14047 1820 nw
tri 14092 1809 14103 1820 se
rect 14103 1809 14166 1820
tri 14166 1809 14177 1820 nw
tri 15165 1809 15176 1820 se
rect 15176 1814 15244 1820
tri 15244 1814 15278 1848 nw
tri 15284 1814 15318 1848 se
rect 15176 1809 15239 1814
tri 15239 1809 15244 1814 nw
tri 15279 1809 15284 1814 se
rect 15284 1809 15318 1814
tri 13924 1771 13962 1809 se
rect 13962 1775 14002 1809
tri 14002 1775 14036 1809 nw
tri 14058 1775 14092 1809 se
rect 14092 1775 14128 1809
rect 13962 1771 13998 1775
tri 13998 1771 14002 1775 nw
tri 14054 1771 14058 1775 se
rect 14058 1771 14128 1775
tri 14128 1771 14166 1809 nw
tri 14190 1771 14228 1809 se
rect 14228 1774 15204 1809
tri 15204 1774 15239 1809 nw
tri 15244 1774 15279 1809 se
rect 15279 1774 15318 1809
tri 15318 1774 15392 1848 nw
tri 15482 1774 15556 1848 se
rect 15556 1774 15650 1848
rect 14228 1771 15201 1774
tri 15201 1771 15204 1774 nw
tri 15241 1771 15244 1774 se
rect 15244 1771 15315 1774
tri 15315 1771 15318 1774 nw
tri 15479 1771 15482 1774 se
rect 15482 1771 15650 1774
rect 13297 776 13320 832
rect 13376 776 13400 832
rect 13456 776 13480 832
rect 13536 776 13560 832
rect 13616 776 13640 832
rect 13696 823 13886 832
rect 13696 815 13878 823
tri 13878 815 13886 823 nw
tri 13919 1766 13924 1771 se
rect 13924 1766 13993 1771
tri 13993 1766 13998 1771 nw
tri 14049 1766 14054 1771 se
rect 14054 1766 14115 1771
rect 13919 1746 13973 1766
tri 13973 1746 13993 1766 nw
tri 14029 1746 14049 1766 se
rect 14049 1758 14115 1766
tri 14115 1758 14128 1771 nw
tri 14177 1758 14190 1771 se
rect 14190 1764 15194 1771
tri 15194 1764 15201 1771 nw
tri 15234 1764 15241 1771 se
rect 15241 1764 15268 1771
rect 14190 1758 15187 1764
rect 14049 1746 14103 1758
tri 14103 1746 14115 1758 nw
tri 14165 1746 14177 1758 se
rect 14177 1757 15187 1758
tri 15187 1757 15194 1764 nw
tri 15227 1757 15234 1764 se
rect 15234 1757 15268 1764
rect 14177 1746 14228 1757
rect 13919 1191 13971 1746
tri 13971 1744 13973 1746 nw
tri 14027 1744 14029 1746 se
rect 14029 1744 14092 1746
tri 14018 1735 14027 1744 se
rect 14027 1735 14092 1744
tri 14092 1735 14103 1746 nw
tri 14154 1735 14165 1746 se
rect 14165 1735 14228 1746
tri 14228 1735 14250 1757 nw
tri 15205 1735 15227 1757 se
rect 15227 1735 15268 1757
rect 13919 1127 13971 1139
rect 13696 803 13866 815
tri 13866 803 13878 815 nw
tri 13907 803 13919 815 se
rect 13919 803 13971 1075
rect 13696 794 13845 803
rect 13696 776 13720 794
rect 13297 746 13720 776
rect 13297 690 13320 746
rect 13376 690 13400 746
rect 13456 738 13720 746
rect 13776 782 13845 794
tri 13845 782 13866 803 nw
tri 13886 782 13907 803 se
rect 13907 793 13971 803
rect 13907 785 13963 793
tri 13963 785 13971 793 nw
tri 14004 1721 14018 1735 se
rect 14018 1721 14078 1735
tri 14078 1721 14092 1735 nw
tri 14140 1721 14154 1735 se
rect 14154 1724 14217 1735
tri 14217 1724 14228 1735 nw
tri 15194 1724 15205 1735 se
rect 15205 1724 15268 1735
tri 15268 1724 15315 1771 nw
tri 15432 1724 15479 1771 se
rect 15479 1724 15650 1771
rect 14154 1721 14212 1724
rect 14004 1719 14076 1721
tri 14076 1719 14078 1721 nw
tri 14138 1719 14140 1721 se
rect 14140 1719 14212 1721
tri 14212 1719 14217 1724 nw
tri 14268 1719 14273 1724 se
rect 14273 1719 15263 1724
tri 15263 1719 15268 1724 nw
tri 15427 1719 15432 1724 se
rect 15432 1719 15650 1724
rect 14004 1707 14064 1719
tri 14064 1707 14076 1719 nw
tri 14126 1707 14138 1719 se
rect 14138 1707 14200 1719
tri 14200 1707 14212 1719 nw
tri 14256 1707 14268 1719 se
rect 14268 1707 15251 1719
tri 15251 1707 15263 1719 nw
tri 15415 1707 15427 1719 se
rect 15427 1707 15650 1719
rect 14004 1191 14056 1707
tri 14056 1699 14064 1707 nw
tri 14118 1699 14126 1707 se
rect 14126 1706 14199 1707
tri 14199 1706 14200 1707 nw
tri 14255 1706 14256 1707 se
rect 14256 1706 15216 1707
rect 14126 1699 14160 1706
rect 14004 1127 14056 1139
rect 13907 782 13930 785
rect 13776 751 13814 782
tri 13814 751 13845 782 nw
tri 13855 751 13886 782 se
rect 13886 752 13930 782
tri 13930 752 13963 785 nw
tri 13971 752 14004 785 se
rect 14004 763 14056 1075
rect 14004 752 14044 763
rect 13886 751 13929 752
tri 13929 751 13930 752 nw
tri 13970 751 13971 752 se
rect 13971 751 14044 752
tri 14044 751 14056 763 nw
tri 14086 1667 14118 1699 se
rect 14118 1667 14160 1699
tri 14160 1667 14199 1706 nw
tri 14216 1667 14255 1706 se
rect 14255 1672 15216 1706
tri 15216 1672 15251 1707 nw
tri 15380 1672 15415 1707 se
rect 15415 1672 15650 1707
rect 14255 1667 14278 1672
rect 14086 1655 14148 1667
tri 14148 1655 14160 1667 nw
tri 14204 1655 14216 1667 se
rect 14216 1655 14278 1667
tri 14278 1655 14295 1672 nw
tri 15363 1655 15380 1672 se
rect 15380 1655 15650 1672
rect 13776 741 13804 751
tri 13804 741 13814 751 nw
tri 13845 741 13855 751 se
rect 13855 741 13919 751
tri 13919 741 13929 751 nw
tri 13960 741 13970 751 se
rect 13970 741 14023 751
rect 13776 738 13792 741
rect 13456 737 13792 738
rect 13456 690 13480 737
rect 13297 681 13480 690
rect 13536 730 13792 737
rect 13536 681 13560 730
rect 13297 674 13560 681
rect 13616 729 13792 730
tri 13792 729 13804 741 nw
tri 13833 729 13845 741 se
rect 13845 729 13889 741
rect 13616 708 13771 729
tri 13771 708 13792 729 nw
tri 13812 708 13833 729 se
rect 13833 711 13889 729
tri 13889 711 13919 741 nw
tri 13949 730 13960 741 se
rect 13960 730 14023 741
tri 14023 730 14044 751 nw
tri 13930 711 13949 730 se
rect 13949 711 14004 730
tri 14004 711 14023 730 nw
tri 14067 711 14086 730 se
rect 14086 713 14143 1655
tri 14143 1650 14148 1655 nw
tri 14199 1650 14204 1655 se
rect 14204 1650 14273 1655
tri 14273 1650 14278 1655 nw
tri 15358 1650 15363 1655 se
rect 15363 1650 15650 1655
tri 14196 1647 14199 1650 se
rect 14199 1647 14270 1650
tri 14270 1647 14273 1650 nw
tri 15355 1647 15358 1650 se
rect 15358 1647 15650 1650
tri 14192 1643 14196 1647 se
rect 14196 1643 14266 1647
tri 14266 1643 14270 1647 nw
tri 15351 1643 15355 1647 se
rect 15355 1643 15650 1647
rect 14086 711 14131 713
rect 13833 708 13886 711
tri 13886 708 13889 711 nw
tri 13927 708 13930 711 se
rect 13930 708 13960 711
rect 13616 706 13730 708
rect 13616 674 13640 706
rect 13297 660 13640 674
rect 13297 604 13320 660
rect 13376 604 13400 660
rect 13456 650 13640 660
rect 13696 667 13730 706
tri 13730 667 13771 708 nw
tri 13771 667 13812 708 se
rect 13812 678 13856 708
tri 13856 678 13886 708 nw
tri 13897 678 13927 708 se
rect 13927 678 13960 708
rect 13812 667 13845 678
tri 13845 667 13856 678 nw
tri 13886 667 13897 678 se
rect 13897 667 13960 678
tri 13960 667 14004 711 nw
tri 14023 667 14067 711 se
rect 14067 701 14131 711
tri 14131 701 14143 713 nw
tri 14171 1622 14192 1643 se
rect 14192 1622 14245 1643
tri 14245 1622 14266 1643 nw
tri 15330 1622 15351 1643 se
rect 15351 1638 15650 1643
rect 15351 1622 15380 1638
rect 14171 1151 14228 1622
tri 14228 1605 14245 1622 nw
tri 15313 1605 15330 1622 se
rect 15330 1605 15380 1622
tri 15299 1591 15313 1605 se
rect 15313 1591 15380 1605
tri 15064 1356 15299 1591 se
rect 15299 1582 15380 1591
rect 15436 1582 15460 1638
rect 15516 1582 15540 1638
rect 15596 1582 15650 1638
rect 15299 1530 15650 1582
rect 15299 1474 15380 1530
rect 15436 1474 15460 1530
rect 15516 1474 15540 1530
rect 15596 1474 15650 1530
rect 15299 1421 15650 1474
rect 15299 1365 15380 1421
rect 15436 1365 15460 1421
rect 15516 1365 15540 1421
rect 15596 1365 15650 1421
rect 15299 1359 15650 1365
rect 15946 1359 15984 1895
rect 15299 1356 15984 1359
tri 15059 1351 15064 1356 se
rect 15064 1351 15984 1356
tri 15058 1350 15059 1351 se
rect 15059 1350 15984 1351
tri 14986 1278 15058 1350 se
rect 15058 1278 15984 1350
tri 14228 1151 14242 1165 sw
rect 14720 1151 14726 1203
rect 14778 1151 14790 1203
rect 14842 1151 14883 1203
rect 14171 1120 14242 1151
tri 14242 1120 14273 1151 sw
tri 14797 1120 14828 1151 ne
rect 14828 1120 14883 1151
rect 14171 1068 14178 1120
rect 14230 1068 14242 1120
rect 14294 1068 14300 1120
rect 14596 1068 14602 1120
rect 14654 1068 14666 1120
rect 14718 1068 14724 1120
tri 14828 1117 14831 1120 ne
rect 14067 667 14097 701
tri 14097 667 14131 701 nw
tri 14137 667 14171 701 se
rect 14171 684 14228 1068
tri 14228 1023 14273 1068 nw
tri 14631 1027 14672 1068 ne
rect 14672 803 14724 1068
tri 14724 803 14765 844 sw
rect 14672 751 14678 803
rect 14730 751 14742 803
rect 14794 751 14800 803
rect 14171 667 14180 684
rect 13696 650 13697 667
rect 13456 641 13697 650
rect 13456 604 13480 641
rect 13297 585 13480 604
rect 13536 634 13697 641
tri 13697 634 13730 667 nw
tri 13738 634 13771 667 se
rect 13771 637 13815 667
tri 13815 637 13845 667 nw
tri 13875 656 13886 667 se
rect 13886 656 13949 667
tri 13949 656 13960 667 nw
tri 14012 656 14023 667 se
rect 14023 656 14086 667
tri 14086 656 14097 667 nw
tri 14126 656 14137 667 se
rect 14137 656 14180 667
tri 13856 637 13875 656 se
rect 13875 648 13941 656
tri 13941 648 13949 656 nw
tri 14004 648 14012 656 se
rect 14012 648 14057 656
rect 13875 637 13930 648
tri 13930 637 13941 648 nw
tri 13993 637 14004 648 se
rect 14004 637 14057 648
rect 13771 634 13783 637
rect 13536 628 13668 634
rect 13536 585 13560 628
rect 13297 574 13560 585
rect 13297 518 13320 574
rect 13376 518 13400 574
rect 13456 572 13560 574
rect 13616 605 13668 628
tri 13668 605 13697 634 nw
tri 13709 605 13738 634 se
rect 13738 605 13783 634
tri 13783 605 13815 637 nw
tri 13824 605 13856 637 se
rect 13856 605 13898 637
tri 13898 605 13930 637 nw
tri 13961 605 13993 637 se
rect 13993 627 14057 637
tri 14057 627 14086 656 nw
tri 14106 636 14126 656 se
rect 14126 636 14180 656
tri 14180 636 14228 684 nw
tri 14097 627 14106 636 se
rect 14106 627 14171 636
tri 14171 627 14180 636 nw
tri 14822 627 14831 636 se
rect 14831 627 14883 1120
rect 13993 605 14035 627
tri 14035 605 14057 627 nw
tri 14075 605 14097 627 se
rect 14097 605 14149 627
tri 14149 605 14171 627 nw
tri 14800 605 14822 627 se
rect 14822 605 14883 627
rect 13616 593 13656 605
tri 13656 593 13668 605 nw
tri 13697 593 13709 605 se
rect 13709 604 13782 605
tri 13782 604 13783 605 nw
tri 13823 604 13824 605 se
rect 13824 604 13886 605
rect 13709 593 13771 604
tri 13771 593 13782 604 nw
tri 13812 593 13823 604 se
rect 13823 593 13886 604
tri 13886 593 13898 605 nw
tri 13949 593 13961 605 se
rect 13961 593 14023 605
tri 14023 593 14035 605 nw
tri 14063 593 14075 605 se
rect 14075 593 14097 605
rect 13616 572 13623 593
rect 13456 560 13623 572
tri 13623 560 13656 593 nw
tri 13664 560 13697 593 se
rect 13697 563 13741 593
tri 13741 563 13771 593 nw
tri 13801 582 13812 593 se
rect 13812 582 13875 593
tri 13875 582 13886 593 nw
tri 13938 582 13949 593 se
rect 13949 582 14012 593
tri 14012 582 14023 593 nw
tri 14052 582 14063 593 se
rect 14063 582 14097 593
tri 13782 563 13801 582 se
rect 13801 574 13867 582
tri 13867 574 13875 582 nw
tri 13930 574 13938 582 se
rect 13938 574 13983 582
rect 13801 563 13856 574
tri 13856 563 13867 574 nw
tri 13919 563 13930 574 se
rect 13930 563 13983 574
rect 13697 560 13731 563
rect 13456 553 13616 560
tri 13616 553 13623 560 nw
tri 13657 553 13664 560 se
rect 13664 553 13731 560
tri 13731 553 13741 563 nw
tri 13772 553 13782 563 se
rect 13782 553 13846 563
tri 13846 553 13856 563 nw
tri 13909 553 13919 563 se
rect 13919 553 13983 563
tri 13983 553 14012 582 nw
tri 14023 553 14052 582 se
rect 14052 553 14097 582
tri 14097 553 14149 605 nw
rect 14672 553 14678 605
rect 14730 553 14742 605
rect 14794 553 14883 605
rect 13456 545 13582 553
rect 13456 518 13480 545
rect 13297 489 13480 518
rect 13536 519 13582 545
tri 13582 519 13616 553 nw
tri 13623 519 13657 553 se
rect 13657 530 13708 553
tri 13708 530 13731 553 nw
tri 13749 530 13772 553 se
rect 13772 530 13823 553
tri 13823 530 13846 553 nw
tri 13886 530 13909 553 se
rect 13909 530 13949 553
rect 13657 519 13697 530
tri 13697 519 13708 530 nw
tri 13738 519 13749 530 se
rect 13749 519 13812 530
tri 13812 519 13823 530 nw
tri 13875 519 13886 530 se
rect 13886 519 13949 530
tri 13949 519 13983 553 nw
tri 13989 519 14023 553 se
rect 13536 489 13549 519
rect 13297 487 13549 489
rect 13297 431 13320 487
rect 13376 431 13400 487
rect 13456 486 13549 487
tri 13549 486 13582 519 nw
tri 13590 486 13623 519 se
rect 13623 489 13667 519
tri 13667 489 13697 519 nw
tri 13727 508 13738 519 se
rect 13738 508 13801 519
tri 13801 508 13812 519 nw
tri 13864 508 13875 519 se
rect 13875 508 13938 519
tri 13938 508 13949 519 nw
tri 13978 508 13989 519 se
rect 13989 508 14023 519
tri 13708 489 13727 508 se
rect 13727 500 13793 508
tri 13793 500 13801 508 nw
tri 13856 500 13864 508 se
rect 13864 500 13909 508
rect 13727 489 13782 500
tri 13782 489 13793 500 nw
tri 13845 489 13856 500 se
rect 13856 489 13909 500
rect 13623 486 13634 489
rect 13456 480 13543 486
tri 13543 480 13549 486 nw
tri 13584 480 13590 486 se
rect 13590 480 13634 486
rect 13456 445 13508 480
tri 13508 445 13543 480 nw
tri 13549 445 13584 480 se
rect 13584 456 13634 480
tri 13634 456 13667 489 nw
tri 13675 456 13708 489 se
rect 13708 456 13738 489
rect 13584 445 13623 456
tri 13623 445 13634 456 nw
tri 13664 445 13675 456 se
rect 13675 445 13738 456
tri 13738 445 13782 489 nw
tri 13801 445 13845 489 se
rect 13845 479 13909 489
tri 13909 479 13938 508 nw
tri 13949 479 13978 508 se
rect 13978 479 14023 508
tri 14023 479 14097 553 nw
rect 13845 456 13886 479
tri 13886 456 13909 479 nw
tri 13926 456 13949 479 se
rect 13949 456 13980 479
rect 13845 445 13875 456
tri 13875 445 13886 456 nw
tri 13915 445 13926 456 se
rect 13926 445 13980 456
rect 13456 436 13499 445
tri 13499 436 13508 445 nw
tri 13540 436 13549 445 se
rect 13549 436 13614 445
tri 13614 436 13623 445 nw
tri 13655 436 13664 445 se
rect 13664 436 13729 445
tri 13729 436 13738 445 nw
tri 13792 436 13801 445 se
rect 13801 436 13866 445
tri 13866 436 13875 445 nw
tri 13906 436 13915 445 se
rect 13915 436 13980 445
tri 13980 436 14023 479 nw
rect 13456 431 13480 436
rect 13297 417 13480 431
tri 13480 417 13499 436 nw
tri 13537 433 13540 436 se
rect 13540 433 13611 436
tri 13611 433 13614 436 nw
tri 13653 434 13655 436 se
rect 13655 434 13727 436
tri 13727 434 13729 436 nw
tri 13790 434 13792 436 se
rect 13792 434 13864 436
tri 13864 434 13866 436 nw
tri 13904 434 13906 436 se
rect 13906 434 13949 436
tri 13652 433 13653 434 se
rect 13653 433 13726 434
tri 13726 433 13727 434 nw
tri 13789 433 13790 434 se
rect 13790 433 13847 434
rect 13537 417 13595 433
tri 13595 417 13611 433 nw
tri 13636 417 13652 433 se
rect 13652 426 13719 433
tri 13719 426 13726 433 nw
tri 13782 426 13789 433 se
rect 13789 426 13847 433
rect 13652 417 13710 426
tri 13710 417 13719 426 nw
tri 13773 417 13782 426 se
rect 13782 417 13847 426
tri 13847 417 13864 434 nw
tri 13887 417 13904 434 se
rect 13904 417 13949 434
rect 13537 291 13589 417
tri 13589 411 13595 417 nw
tri 13634 415 13636 417 se
rect 13636 415 13708 417
tri 13708 415 13710 417 nw
tri 13771 415 13773 417 se
rect 13773 415 13835 417
tri 13630 411 13634 415 se
rect 13634 411 13704 415
tri 13704 411 13708 415 nw
tri 13767 411 13771 415 se
rect 13771 411 13835 415
tri 13620 401 13630 411 se
rect 13630 401 13694 411
tri 13694 401 13704 411 nw
tri 13757 401 13767 411 se
rect 13767 405 13835 411
tri 13835 405 13847 417 nw
tri 13875 405 13887 417 se
rect 13887 405 13949 417
tri 13949 405 13980 436 nw
rect 13767 401 13814 405
rect 13620 384 13677 401
tri 13677 384 13694 401 nw
tri 13740 384 13757 401 se
rect 13757 384 13814 401
tri 13814 384 13835 405 nw
tri 13854 384 13875 405 se
rect 13875 384 13928 405
tri 13928 384 13949 405 nw
rect 13620 -630 13672 384
tri 13672 379 13677 384 nw
tri 13735 379 13740 384 se
rect 13740 379 13802 384
tri 13728 372 13735 379 se
rect 13735 372 13802 379
tri 13802 372 13814 384 nw
tri 13842 372 13854 384 se
rect 13854 372 13916 384
tri 13916 372 13928 384 nw
tri 13716 360 13728 372 se
rect 13728 371 13801 372
tri 13801 371 13802 372 nw
tri 13841 371 13842 372 se
rect 13842 371 13875 372
rect 13728 360 13790 371
tri 13790 360 13801 371 nw
tri 13830 360 13841 371 se
rect 13841 360 13875 371
tri 13703 347 13716 360 se
rect 13716 347 13777 360
tri 13777 347 13790 360 nw
tri 13817 347 13830 360 se
rect 13830 347 13875 360
rect 12725 -1281 13230 -1242
tri 13230 -1281 13269 -1242 nw
rect 12725 -1373 13167 -1281
tri 13167 -1344 13230 -1281 nw
tri 13629 -1933 13703 -1859 se
rect 13703 -1881 13755 347
tri 13755 325 13777 347 nw
tri 13801 331 13817 347 se
rect 13817 331 13875 347
tri 13875 331 13916 372 nw
tri 13795 325 13801 331 se
rect 13801 325 13864 331
tri 13790 320 13795 325 se
rect 13795 320 13864 325
tri 13864 320 13875 331 nw
tri 13783 313 13790 320 se
rect 13790 313 13857 320
tri 13857 313 13864 320 nw
rect 13783 308 13852 313
tri 13852 308 13857 313 nw
rect 13783 -200 13835 308
tri 13835 291 13852 308 nw
rect 13783 -281 13835 -252
rect 13783 -339 13835 -333
tri 14833 -463 14849 -447 nw
tri 14770 -1381 14797 -1354 se
tri 13703 -1933 13755 -1881 nw
tri 13586 -1976 13629 -1933 se
tri 13555 -2007 13586 -1976 se
rect 13586 -2007 13629 -1976
tri 13629 -2007 13703 -1933 nw
tri 13481 -2081 13555 -2007 se
tri 13555 -2081 13629 -2007 nw
tri 13407 -2155 13481 -2081 se
tri 13481 -2155 13555 -2081 nw
tri 13388 -2174 13407 -2155 se
rect 13407 -2174 13451 -2155
tri 9817 -2187 9830 -2174 sw
tri 13377 -2185 13388 -2174 se
rect 13388 -2185 13451 -2174
tri 13451 -2185 13481 -2155 nw
rect 13377 -2187 13449 -2185
tri 13449 -2187 13451 -2185 nw
rect 9698 -2311 9830 -2187
tri 9830 -2311 9954 -2187 sw
rect 9698 -2346 9954 -2311
tri 9954 -2346 9989 -2311 sw
rect 9698 -2871 9989 -2346
rect 9698 -2927 9728 -2871
rect 9784 -2927 9808 -2871
rect 9864 -2927 9888 -2871
rect 9944 -2927 9989 -2871
rect 9698 -2955 9989 -2927
rect 9698 -3011 9728 -2955
rect 9784 -3011 9808 -2955
rect 9864 -3011 9888 -2955
rect 9944 -3011 9989 -2955
rect 9698 -3039 9989 -3011
rect 9698 -3095 9728 -3039
rect 9784 -3095 9808 -3039
rect 9864 -3095 9888 -3039
rect 9944 -3095 9989 -3039
rect 9698 -3123 9989 -3095
rect 9698 -3179 9728 -3123
rect 9784 -3179 9808 -3123
rect 9864 -3179 9888 -3123
rect 9944 -3179 9989 -3123
rect 9698 -3207 9989 -3179
rect 9698 -3263 9728 -3207
rect 9784 -3263 9808 -3207
rect 9864 -3263 9888 -3207
rect 9944 -3263 9989 -3207
rect 9698 -3291 9989 -3263
rect 9698 -3347 9728 -3291
rect 9784 -3347 9808 -3291
rect 9864 -3347 9888 -3291
rect 9944 -3347 9989 -3291
rect 9698 -3375 9989 -3347
rect 9698 -3431 9728 -3375
rect 9784 -3431 9808 -3375
rect 9864 -3431 9888 -3375
rect 9944 -3431 9989 -3375
rect 9698 -3459 9989 -3431
rect 9698 -3515 9728 -3459
rect 9784 -3515 9808 -3459
rect 9864 -3515 9888 -3459
rect 9944 -3515 9989 -3459
rect 9698 -3543 9989 -3515
rect 9698 -3599 9728 -3543
rect 9784 -3599 9808 -3543
rect 9864 -3599 9888 -3543
rect 9944 -3599 9989 -3543
rect 9698 -3628 9989 -3599
rect 9698 -3684 9728 -3628
rect 9784 -3684 9808 -3628
rect 9864 -3684 9888 -3628
rect 9944 -3684 9989 -3628
rect 9698 -3699 9989 -3684
rect 13377 -5730 13429 -2187
tri 13429 -2207 13449 -2187 nw
rect 14986 -2881 15984 1278
rect 16121 249 16633 1792
rect 19429 1771 20310 2805
rect 19429 1719 19435 1771
rect 19487 1719 19504 1771
rect 19556 1719 19572 1771
rect 19624 1719 19640 1771
rect 19692 1719 19708 1771
rect 19760 1719 19776 1771
rect 19828 1719 19844 1771
rect 19896 1719 19912 1771
rect 19964 1719 19980 1771
rect 20032 1719 20048 1771
rect 20100 1719 20116 1771
rect 20168 1719 20184 1771
rect 20236 1719 20252 1771
rect 20304 1719 20310 1771
rect 19429 1707 20310 1719
rect 19429 1655 19435 1707
rect 19487 1655 19504 1707
rect 19556 1655 19572 1707
rect 19624 1655 19640 1707
rect 19692 1655 19708 1707
rect 19760 1655 19776 1707
rect 19828 1655 19844 1707
rect 19896 1655 19912 1707
rect 19964 1655 19980 1707
rect 20032 1655 20048 1707
rect 20100 1655 20116 1707
rect 20168 1655 20184 1707
rect 20236 1655 20252 1707
rect 20304 1655 20310 1707
rect 19429 1643 20310 1655
rect 19429 1591 19435 1643
rect 19487 1591 19504 1643
rect 19556 1591 19572 1643
rect 19624 1591 19640 1643
rect 19692 1591 19708 1643
rect 19760 1591 19776 1643
rect 19828 1591 19844 1643
rect 19896 1591 19912 1643
rect 19964 1591 19980 1643
rect 20032 1591 20048 1643
rect 20100 1591 20116 1643
rect 20168 1591 20184 1643
rect 20236 1591 20252 1643
rect 20304 1591 20310 1643
rect 19429 436 20310 1591
rect 20833 1771 21151 7880
rect 21617 8425 21641 10185
rect 21937 11545 21963 14801
rect 23032 14417 23072 17960
tri 23072 17942 23130 18000 nw
rect 29456 17953 29488 18009
rect 29544 17953 29568 18009
rect 29624 17953 29648 18009
rect 29704 17953 29728 18009
rect 29784 17953 29816 18009
rect 26316 17914 26572 17940
rect 26316 17858 26328 17914
rect 26384 17858 26416 17914
rect 26472 17858 26504 17914
rect 26560 17858 26572 17914
rect 26316 17834 26572 17858
rect 26316 17778 26328 17834
rect 26384 17778 26416 17834
rect 26472 17778 26504 17834
rect 26560 17778 26572 17834
rect 26316 17737 26572 17778
rect 29456 17922 29816 17953
rect 29456 17866 29488 17922
rect 29544 17866 29568 17922
rect 29624 17866 29648 17922
rect 29704 17866 29728 17922
rect 29784 17866 29816 17922
rect 29456 17835 29816 17866
rect 29456 17779 29488 17835
rect 29544 17779 29568 17835
rect 29624 17779 29648 17835
rect 29704 17779 29728 17835
rect 29784 17779 29816 17835
rect 29456 17770 29816 17779
rect 30985 18748 31022 18804
rect 31078 18791 31102 18804
rect 31158 18791 31182 18804
rect 31238 18791 31262 18804
rect 31318 18791 31342 18804
rect 31398 18791 31435 18804
rect 30985 18739 31029 18748
rect 31081 18739 31093 18791
rect 31337 18748 31342 18791
rect 31145 18739 31157 18748
rect 31209 18739 31221 18748
rect 31273 18739 31285 18748
rect 31337 18739 31349 18748
rect 31401 18739 31435 18791
rect 30985 18724 31435 18739
rect 30985 18723 31029 18724
rect 30985 18667 31022 18723
rect 31081 18672 31093 18724
rect 31145 18723 31157 18724
rect 31209 18723 31221 18724
rect 31273 18723 31285 18724
rect 31337 18723 31349 18724
rect 31337 18672 31342 18723
rect 31401 18672 31435 18724
rect 31078 18667 31102 18672
rect 31158 18667 31182 18672
rect 31238 18667 31262 18672
rect 31318 18667 31342 18672
rect 31398 18667 31435 18672
rect 30985 18657 31435 18667
rect 30985 18642 31029 18657
rect 30985 18586 31022 18642
rect 31081 18605 31093 18657
rect 31145 18642 31157 18657
rect 31209 18642 31221 18657
rect 31273 18642 31285 18657
rect 31337 18642 31349 18657
rect 31337 18605 31342 18642
rect 31401 18605 31435 18657
rect 31078 18590 31102 18605
rect 31158 18590 31182 18605
rect 31238 18590 31262 18605
rect 31318 18590 31342 18605
rect 31398 18590 31435 18605
rect 30985 18561 31029 18586
rect 30985 18505 31022 18561
rect 31081 18538 31093 18590
rect 31337 18586 31342 18590
rect 31145 18561 31157 18586
rect 31209 18561 31221 18586
rect 31273 18561 31285 18586
rect 31337 18561 31349 18586
rect 31337 18538 31342 18561
rect 31401 18538 31435 18590
rect 31078 18523 31102 18538
rect 31158 18523 31182 18538
rect 31238 18523 31262 18538
rect 31318 18523 31342 18538
rect 31398 18523 31435 18538
rect 30985 18480 31029 18505
rect 30985 18424 31022 18480
rect 31081 18471 31093 18523
rect 31337 18505 31342 18523
rect 31145 18480 31157 18505
rect 31209 18480 31221 18505
rect 31273 18480 31285 18505
rect 31337 18480 31349 18505
rect 31337 18471 31342 18480
rect 31401 18471 31435 18523
rect 31078 18456 31102 18471
rect 31158 18456 31182 18471
rect 31238 18456 31262 18471
rect 31318 18456 31342 18471
rect 31398 18456 31435 18471
rect 30985 18404 31029 18424
rect 31081 18404 31093 18456
rect 31337 18424 31342 18456
rect 31145 18404 31157 18424
rect 31209 18404 31221 18424
rect 31273 18404 31285 18424
rect 31337 18404 31349 18424
rect 31401 18404 31435 18456
rect 30985 18398 31435 18404
rect 30985 18342 31022 18398
rect 31078 18389 31102 18398
rect 31158 18389 31182 18398
rect 31238 18389 31262 18398
rect 31318 18389 31342 18398
rect 31398 18389 31435 18398
rect 30985 18337 31029 18342
rect 31081 18337 31093 18389
rect 31337 18342 31342 18389
rect 31145 18337 31157 18342
rect 31209 18337 31221 18342
rect 31273 18337 31285 18342
rect 31337 18337 31349 18342
rect 31401 18337 31435 18389
rect 30985 18322 31435 18337
rect 30985 18316 31029 18322
rect 30985 18260 31022 18316
rect 31081 18270 31093 18322
rect 31145 18316 31157 18322
rect 31209 18316 31221 18322
rect 31273 18316 31285 18322
rect 31337 18316 31349 18322
rect 31337 18270 31342 18316
rect 31401 18270 31435 18322
rect 31078 18260 31102 18270
rect 31158 18260 31182 18270
rect 31238 18260 31262 18270
rect 31318 18260 31342 18270
rect 31398 18260 31435 18270
rect 30985 18255 31435 18260
rect 30985 18234 31029 18255
rect 30985 18178 31022 18234
rect 31081 18203 31093 18255
rect 31145 18234 31157 18255
rect 31209 18234 31221 18255
rect 31273 18234 31285 18255
rect 31337 18234 31349 18255
rect 31337 18203 31342 18234
rect 31401 18203 31435 18255
rect 31078 18188 31102 18203
rect 31158 18188 31182 18203
rect 31238 18188 31262 18203
rect 31318 18188 31342 18203
rect 31398 18188 31435 18203
rect 30985 18152 31029 18178
rect 30985 18096 31022 18152
rect 31081 18136 31093 18188
rect 31337 18178 31342 18188
rect 31145 18152 31157 18178
rect 31209 18152 31221 18178
rect 31273 18152 31285 18178
rect 31337 18152 31349 18178
rect 31337 18136 31342 18152
rect 31401 18136 31435 18188
rect 31078 18121 31102 18136
rect 31158 18121 31182 18136
rect 31238 18121 31262 18136
rect 31318 18121 31342 18136
rect 31398 18121 31435 18136
rect 30985 18070 31029 18096
rect 30985 18014 31022 18070
rect 31081 18069 31093 18121
rect 31337 18096 31342 18121
rect 31145 18070 31157 18096
rect 31209 18070 31221 18096
rect 31273 18070 31285 18096
rect 31337 18070 31349 18096
rect 31337 18069 31342 18070
rect 31401 18069 31435 18121
rect 31078 18014 31102 18069
rect 31158 18014 31182 18069
rect 31238 18014 31262 18069
rect 31318 18014 31342 18069
rect 31398 18014 31435 18069
rect 30985 17988 31435 18014
rect 30985 17932 31022 17988
rect 31078 17932 31102 17988
rect 31158 17932 31182 17988
rect 31238 17932 31262 17988
rect 31318 17932 31342 17988
rect 31398 17932 31435 17988
rect 30985 17906 31435 17932
rect 30985 17850 31022 17906
rect 31078 17850 31102 17906
rect 31158 17850 31182 17906
rect 31238 17850 31262 17906
rect 31318 17850 31342 17906
rect 31398 17850 31435 17906
rect 30985 17824 31435 17850
rect 30985 17768 31022 17824
rect 31078 17768 31102 17824
rect 31158 17768 31182 17824
rect 31238 17768 31262 17824
rect 31318 17768 31342 17824
rect 31398 17768 31435 17824
rect 30985 17759 31435 17768
tri 23072 14417 23105 14450 sw
rect 23032 14365 23038 14417
rect 23090 14365 23102 14417
rect 23154 14365 23160 14417
rect 23755 14365 23761 14417
rect 23813 14365 23825 14417
rect 23877 14365 23883 14417
tri 23798 14336 23827 14365 ne
tri 21963 11545 22028 11610 sw
rect 21937 8425 22028 11545
rect 21617 8400 22028 8425
rect 21617 8344 21641 8400
rect 21697 8344 21721 8400
rect 21777 8344 21801 8400
rect 21857 8344 21881 8400
rect 21937 8344 22028 8400
rect 21617 8319 22028 8344
rect 21617 8263 21641 8319
rect 21697 8263 21721 8319
rect 21777 8263 21801 8319
rect 21857 8263 21881 8319
rect 21937 8263 22028 8319
rect 21617 8238 22028 8263
rect 21617 8182 21641 8238
rect 21697 8182 21721 8238
rect 21777 8182 21801 8238
rect 21857 8182 21881 8238
rect 21937 8182 22028 8238
rect 21617 8157 22028 8182
rect 21617 8101 21641 8157
rect 21697 8101 21721 8157
rect 21777 8101 21801 8157
rect 21857 8101 21881 8157
rect 21937 8101 22028 8157
rect 21617 8083 22028 8101
rect 21617 8031 21634 8083
rect 21686 8076 21701 8083
rect 21753 8076 21768 8083
rect 21820 8076 21834 8083
rect 21886 8076 21900 8083
rect 21697 8031 21701 8076
rect 21952 8031 21966 8083
rect 22018 8031 22028 8083
rect 21617 8020 21641 8031
rect 21697 8020 21721 8031
rect 21777 8020 21801 8031
rect 21857 8020 21881 8031
rect 21937 8020 22028 8031
rect 21617 8019 22028 8020
rect 21617 7967 21634 8019
rect 21686 7995 21701 8019
rect 21753 7995 21768 8019
rect 21820 7995 21834 8019
rect 21886 7995 21900 8019
rect 21697 7967 21701 7995
rect 21952 7967 21966 8019
rect 22018 7967 22028 8019
rect 21617 7955 21641 7967
rect 21697 7955 21721 7967
rect 21777 7955 21801 7967
rect 21857 7955 21881 7967
rect 21937 7955 22028 7967
rect 21617 7903 21634 7955
rect 21697 7939 21701 7955
rect 21686 7914 21701 7939
rect 21753 7914 21768 7939
rect 21820 7914 21834 7939
rect 21886 7914 21900 7939
rect 21697 7903 21701 7914
rect 21952 7903 21966 7955
rect 22018 7903 22028 7955
rect 21617 7858 21641 7903
rect 21697 7858 21721 7903
rect 21777 7858 21801 7903
rect 21857 7858 21881 7903
rect 21937 7858 22028 7903
rect 20833 1719 20844 1771
rect 20896 1719 20926 1771
rect 20978 1719 21008 1771
rect 21060 1719 21090 1771
rect 21142 1719 21151 1771
rect 20833 1707 21151 1719
rect 20833 1655 20844 1707
rect 20896 1655 20926 1707
rect 20978 1655 21008 1707
rect 21060 1655 21090 1707
rect 21142 1655 21151 1707
rect 20833 1643 21151 1655
rect 20833 1591 20844 1643
rect 20896 1591 20926 1643
rect 20978 1591 21008 1643
rect 21060 1591 21090 1643
rect 21142 1591 21151 1643
rect 20833 1350 21151 1591
tri 21538 6079 21617 6158 se
rect 21617 6079 22028 7858
rect 21538 1771 22028 6079
rect 22215 8095 22725 8139
rect 22215 8039 22231 8095
rect 22287 8083 22316 8095
rect 22372 8083 22400 8095
rect 22456 8083 22484 8095
rect 22540 8083 22568 8095
rect 22624 8083 22652 8095
rect 22215 8031 22239 8039
rect 22291 8031 22309 8083
rect 22372 8039 22379 8083
rect 22638 8039 22652 8083
rect 22708 8039 22725 8095
rect 22361 8031 22379 8039
rect 22431 8031 22448 8039
rect 22500 8031 22517 8039
rect 22569 8031 22586 8039
rect 22638 8031 22655 8039
rect 22707 8031 22725 8039
rect 22215 8019 22725 8031
rect 22215 8015 22239 8019
rect 22215 7959 22231 8015
rect 22291 7967 22309 8019
rect 22361 8015 22379 8019
rect 22431 8015 22448 8019
rect 22500 8015 22517 8019
rect 22569 8015 22586 8019
rect 22638 8015 22655 8019
rect 22707 8015 22725 8019
rect 22372 7967 22379 8015
rect 22638 7967 22652 8015
rect 22287 7959 22316 7967
rect 22372 7959 22400 7967
rect 22456 7959 22484 7967
rect 22540 7959 22568 7967
rect 22624 7959 22652 7967
rect 22708 7959 22725 8015
rect 22215 7955 22725 7959
rect 22215 7935 22239 7955
rect 22215 7879 22231 7935
rect 22291 7903 22309 7955
rect 22361 7935 22379 7955
rect 22431 7935 22448 7955
rect 22500 7935 22517 7955
rect 22569 7935 22586 7955
rect 22638 7935 22655 7955
rect 22707 7935 22725 7955
rect 22372 7903 22379 7935
rect 22638 7903 22652 7935
rect 22287 7879 22316 7903
rect 22372 7879 22400 7903
rect 22456 7879 22484 7903
rect 22540 7879 22568 7903
rect 22624 7879 22652 7903
rect 22708 7879 22725 7935
rect 22215 6404 22725 7879
rect 21538 1719 21550 1771
rect 21602 1719 21620 1771
rect 21672 1719 21690 1771
rect 21742 1719 21759 1771
rect 21811 1719 21828 1771
rect 21880 1719 21897 1771
rect 21949 1719 21966 1771
rect 22018 1719 22028 1771
rect 21538 1707 22028 1719
rect 21538 1655 21550 1707
rect 21602 1655 21620 1707
rect 21672 1655 21690 1707
rect 21742 1655 21759 1707
rect 21811 1655 21828 1707
rect 21880 1655 21897 1707
rect 21949 1655 21966 1707
rect 22018 1655 22028 1707
rect 21538 1643 22028 1655
rect 21538 1591 21550 1643
rect 21602 1591 21620 1643
rect 21672 1591 21690 1643
rect 21742 1591 21759 1643
rect 21811 1591 21828 1643
rect 21880 1591 21897 1643
rect 21949 1591 21966 1643
rect 22018 1591 22028 1643
tri 21151 1350 21162 1361 sw
rect 20833 1274 21162 1350
tri 21162 1274 21238 1350 sw
rect 20833 1229 21238 1274
tri 20833 1142 20920 1229 ne
rect 19429 384 19443 436
rect 19495 384 19510 436
rect 19562 384 19577 436
rect 19629 384 19644 436
rect 19696 384 19711 436
rect 19763 384 19778 436
rect 19830 384 19845 436
rect 19897 384 19912 436
rect 19964 384 19979 436
rect 20031 384 20046 436
rect 20098 384 20113 436
rect 20165 384 20179 436
rect 20231 384 20245 436
rect 20297 384 20310 436
rect 19429 372 20310 384
rect 19429 320 19443 372
rect 19495 320 19510 372
rect 19562 320 19577 372
rect 19629 320 19644 372
rect 19696 320 19711 372
rect 19763 320 19778 372
rect 19830 320 19845 372
rect 19897 320 19912 372
rect 19964 320 19979 372
rect 20031 320 20046 372
rect 20098 320 20113 372
rect 20165 320 20179 372
rect 20231 320 20245 372
rect 20297 320 20310 372
rect 19429 308 20310 320
rect 19429 256 19443 308
rect 19495 256 19510 308
rect 19562 256 19577 308
rect 19629 256 19644 308
rect 19696 256 19711 308
rect 19763 256 19778 308
rect 19830 256 19845 308
rect 19897 256 19912 308
rect 19964 256 19979 308
rect 20031 256 20046 308
rect 20098 256 20113 308
rect 20165 256 20179 308
rect 20231 256 20245 308
rect 20297 256 20310 308
rect 19429 244 20310 256
rect 19429 192 19443 244
rect 19495 192 19510 244
rect 19562 192 19577 244
rect 19629 192 19644 244
rect 19696 192 19711 244
rect 19763 192 19778 244
rect 19830 192 19845 244
rect 19897 192 19912 244
rect 19964 192 19979 244
rect 20031 192 20046 244
rect 20098 192 20113 244
rect 20165 192 20179 244
rect 20231 192 20245 244
rect 20297 192 20310 244
rect 19429 -2452 20310 192
rect 20920 436 21238 1229
rect 20920 384 20931 436
rect 20983 384 21011 436
rect 21063 384 21091 436
rect 21143 384 21171 436
rect 21223 384 21238 436
rect 20920 372 21238 384
rect 20920 320 20931 372
rect 20983 320 21011 372
rect 21063 320 21091 372
rect 21143 320 21171 372
rect 21223 320 21238 372
rect 20920 308 21238 320
rect 20920 256 20931 308
rect 20983 256 21011 308
rect 21063 256 21091 308
rect 21143 256 21171 308
rect 21223 256 21238 308
rect 20920 244 21238 256
rect 20920 192 20931 244
rect 20983 192 21011 244
rect 21063 192 21091 244
rect 21143 192 21171 244
rect 21223 192 21238 244
tri 20855 -2366 20920 -2301 se
rect 20920 -2366 21238 192
tri 19429 -2512 19489 -2452 ne
rect 19489 -2512 20310 -2452
tri 20310 -2512 20456 -2366 sw
tri 20709 -2512 20855 -2366 se
rect 20855 -2370 21238 -2366
rect 20855 -2512 21096 -2370
tri 21096 -2512 21238 -2370 nw
rect 21538 436 22028 1591
rect 22090 3063 22146 3072
rect 22090 2983 22146 3007
rect 22090 2903 22146 2927
rect 22090 2823 22146 2847
rect 22090 2743 22146 2767
rect 22090 2663 22146 2687
rect 22090 2583 22146 2607
rect 22090 2503 22146 2527
rect 22090 2423 22146 2447
rect 22090 2343 22146 2367
rect 22090 2263 22146 2287
rect 22090 2183 22146 2207
rect 22090 2103 22146 2127
rect 22090 2023 22146 2047
rect 22090 1943 22146 1967
rect 22090 1863 22146 1887
rect 22090 1782 22146 1807
rect 22090 1701 22146 1726
rect 22090 1620 22146 1645
rect 22090 1539 22146 1564
rect 22090 1474 22146 1483
rect 22215 2470 22431 6404
tri 22431 6349 22486 6404 nw
tri 22562 6349 22617 6404 ne
rect 22459 6300 22589 6309
rect 22459 6184 22466 6300
rect 22582 6184 22589 6300
rect 22459 4431 22589 6184
tri 22431 2470 22486 2525 sw
tri 22562 2470 22617 2525 se
rect 22617 2470 22725 6404
rect 22215 1771 22725 2470
rect 22215 1719 22239 1771
rect 22291 1719 22309 1771
rect 22361 1719 22379 1771
rect 22431 1719 22448 1771
rect 22500 1719 22517 1771
rect 22569 1719 22586 1771
rect 22638 1719 22655 1771
rect 22707 1719 22725 1771
rect 22215 1707 22725 1719
rect 22215 1655 22239 1707
rect 22291 1655 22309 1707
rect 22361 1655 22379 1707
rect 22431 1655 22448 1707
rect 22500 1655 22517 1707
rect 22569 1655 22586 1707
rect 22638 1655 22655 1707
rect 22707 1655 22725 1707
rect 22215 1643 22725 1655
rect 22215 1591 22239 1643
rect 22291 1591 22309 1643
rect 22361 1591 22379 1643
rect 22431 1591 22448 1643
rect 22500 1591 22517 1643
rect 22569 1591 22586 1643
rect 22638 1591 22655 1643
rect 22707 1591 22725 1643
rect 21538 384 21550 436
rect 21602 384 21619 436
rect 21671 384 21688 436
rect 21740 384 21757 436
rect 21809 384 21826 436
rect 21878 384 21895 436
rect 21947 384 21964 436
rect 22016 384 22028 436
rect 21538 372 22028 384
rect 21538 320 21550 372
rect 21602 320 21619 372
rect 21671 320 21688 372
rect 21740 320 21757 372
rect 21809 320 21826 372
rect 21878 320 21895 372
rect 21947 320 21964 372
rect 22016 320 22028 372
rect 21538 308 22028 320
rect 21538 256 21550 308
rect 21602 256 21619 308
rect 21671 256 21688 308
rect 21740 256 21757 308
rect 21809 256 21826 308
rect 21878 256 21895 308
rect 21947 256 21964 308
rect 22016 256 22028 308
rect 21538 244 22028 256
rect 21538 192 21550 244
rect 21602 192 21619 244
rect 21671 192 21688 244
rect 21740 192 21757 244
rect 21809 192 21826 244
rect 21878 192 21895 244
rect 21947 192 21964 244
rect 22016 192 22028 244
tri 19489 -2862 19839 -2512 ne
rect 19839 -2862 20750 -2512
tri 20750 -2858 21096 -2512 nw
rect 21538 -2685 22028 192
tri 19839 -2868 19845 -2862 ne
rect 19845 -2868 20750 -2862
tri 19845 -2872 19849 -2868 ne
rect 19849 -2872 20750 -2868
rect 14986 -2937 15246 -2881
rect 15302 -2937 15326 -2881
rect 15382 -2937 15406 -2881
rect 15462 -2937 15486 -2881
rect 15542 -2937 15566 -2881
rect 15622 -2937 15646 -2881
rect 15702 -2937 15726 -2881
rect 15782 -2937 15806 -2881
rect 15862 -2937 15886 -2881
rect 15942 -2937 15984 -2881
tri 19849 -2920 19897 -2872 ne
rect 19897 -2920 20750 -2872
tri 19897 -2932 19909 -2920 ne
rect 19909 -2932 20750 -2920
rect 14986 -2964 15984 -2937
rect 14986 -3020 15246 -2964
rect 15302 -3020 15326 -2964
rect 15382 -3020 15406 -2964
rect 15462 -3020 15486 -2964
rect 15542 -3020 15566 -2964
rect 15622 -3020 15646 -2964
rect 15702 -3020 15726 -2964
rect 15782 -3020 15806 -2964
rect 15862 -3020 15886 -2964
rect 15942 -3020 15984 -2964
tri 19909 -2984 19961 -2932 ne
rect 19961 -2984 20750 -2932
tri 19961 -2992 19969 -2984 ne
rect 19969 -2992 20750 -2984
rect 14986 -3047 15984 -3020
rect 14986 -3103 15246 -3047
rect 15302 -3103 15326 -3047
rect 15382 -3103 15406 -3047
rect 15462 -3103 15486 -3047
rect 15542 -3103 15566 -3047
rect 15622 -3103 15646 -3047
rect 15702 -3103 15726 -3047
rect 15782 -3103 15806 -3047
rect 15862 -3103 15886 -3047
rect 15942 -3103 15984 -3047
rect 14986 -3131 15984 -3103
rect 14986 -3187 15246 -3131
rect 15302 -3187 15326 -3131
rect 15382 -3187 15406 -3131
rect 15462 -3187 15486 -3131
rect 15542 -3187 15566 -3131
rect 15622 -3187 15646 -3131
rect 15702 -3187 15726 -3131
rect 15782 -3187 15806 -3131
rect 15862 -3187 15886 -3131
rect 15942 -3187 15984 -3131
rect 14986 -3215 15984 -3187
rect 14986 -3271 15246 -3215
rect 15302 -3271 15326 -3215
rect 15382 -3271 15406 -3215
rect 15462 -3271 15486 -3215
rect 15542 -3271 15566 -3215
rect 15622 -3271 15646 -3215
rect 15702 -3271 15726 -3215
rect 15782 -3271 15806 -3215
rect 15862 -3271 15886 -3215
rect 15942 -3271 15984 -3215
rect 14986 -3299 15984 -3271
rect 14986 -3355 15246 -3299
rect 15302 -3355 15326 -3299
rect 15382 -3355 15406 -3299
rect 15462 -3355 15486 -3299
rect 15542 -3355 15566 -3299
rect 15622 -3355 15646 -3299
rect 15702 -3355 15726 -3299
rect 15782 -3355 15806 -3299
rect 15862 -3355 15886 -3299
rect 15942 -3355 15984 -3299
rect 14986 -3383 15984 -3355
rect 14986 -3439 15246 -3383
rect 15302 -3439 15326 -3383
rect 15382 -3439 15406 -3383
rect 15462 -3439 15486 -3383
rect 15542 -3439 15566 -3383
rect 15622 -3439 15646 -3383
rect 15702 -3439 15726 -3383
rect 15782 -3439 15806 -3383
rect 15862 -3439 15886 -3383
rect 15942 -3439 15984 -3383
rect 14986 -3467 15984 -3439
rect 14986 -3523 15246 -3467
rect 15302 -3523 15326 -3467
rect 15382 -3523 15406 -3467
rect 15462 -3523 15486 -3467
rect 15542 -3523 15566 -3467
rect 15622 -3523 15646 -3467
rect 15702 -3523 15726 -3467
rect 15782 -3523 15806 -3467
rect 15862 -3523 15886 -3467
rect 15942 -3523 15984 -3467
rect 14986 -3551 15984 -3523
rect 14986 -3607 15246 -3551
rect 15302 -3607 15326 -3551
rect 15382 -3607 15406 -3551
rect 15462 -3607 15486 -3551
rect 15542 -3607 15566 -3551
rect 15622 -3607 15646 -3551
rect 15702 -3607 15726 -3551
rect 15782 -3607 15806 -3551
rect 15862 -3607 15886 -3551
rect 15942 -3607 15984 -3551
rect 14986 -3635 15984 -3607
rect 14986 -3691 15246 -3635
rect 15302 -3691 15326 -3635
rect 15382 -3691 15406 -3635
rect 15462 -3691 15486 -3635
rect 15542 -3691 15566 -3635
rect 15622 -3691 15646 -3635
rect 15702 -3691 15726 -3635
rect 15782 -3691 15806 -3635
rect 15862 -3691 15886 -3635
rect 15942 -3691 15984 -3635
rect 14986 -3721 15984 -3691
rect 17432 -3044 17438 -2992
rect 17490 -3044 17502 -2992
rect 17554 -3044 17560 -2992
tri 19969 -3044 20021 -2992 ne
rect 20021 -3044 20750 -2992
tri 13429 -5730 13451 -5708 sw
tri 13377 -5804 13451 -5730 ne
tri 13451 -5804 13525 -5730 sw
tri 13451 -5878 13525 -5804 ne
tri 13525 -5870 13591 -5804 sw
rect 13525 -5878 13591 -5870
tri 13525 -5892 13539 -5878 ne
rect 13539 -7454 13591 -5878
rect 17012 -6078 17332 -6068
rect 17432 -6078 17484 -3044
tri 20021 -3333 20310 -3044 ne
rect 20310 -3333 20750 -3044
tri 20310 -3519 20496 -3333 ne
rect 20496 -3519 20750 -3333
rect 21538 -2862 21851 -2685
tri 21851 -2862 22028 -2685 nw
rect 22215 436 22725 1591
rect 22215 384 22235 436
rect 22287 384 22304 436
rect 22356 384 22373 436
rect 22425 384 22442 436
rect 22494 384 22511 436
rect 22563 384 22580 436
rect 22632 384 22649 436
rect 22701 384 22725 436
rect 22215 372 22725 384
rect 22215 320 22235 372
rect 22287 320 22304 372
rect 22356 320 22373 372
rect 22425 320 22442 372
rect 22494 320 22511 372
rect 22563 320 22580 372
rect 22632 320 22649 372
rect 22701 320 22725 372
rect 22215 308 22725 320
rect 22215 256 22235 308
rect 22287 256 22304 308
rect 22356 256 22373 308
rect 22425 256 22442 308
rect 22494 256 22511 308
rect 22563 256 22580 308
rect 22632 256 22649 308
rect 22701 256 22725 308
rect 22215 244 22725 256
rect 22215 192 22235 244
rect 22287 192 22304 244
rect 22356 192 22373 244
rect 22425 192 22442 244
rect 22494 192 22511 244
rect 22563 192 22580 244
rect 22632 192 22649 244
rect 22701 192 22725 244
rect 21538 -2868 21845 -2862
tri 21845 -2868 21851 -2862 nw
rect 21538 -4060 21843 -2868
tri 21843 -2870 21845 -2868 nw
tri 22204 -3800 22215 -3789 se
rect 22215 -3800 22725 192
rect 23413 3189 23623 3204
rect 23413 2493 23450 3189
rect 23586 2493 23623 3189
rect 23413 2468 23623 2493
rect 23413 2412 23450 2468
rect 23506 2412 23530 2468
rect 23586 2412 23623 2468
rect 23413 2387 23623 2412
rect 23413 2331 23450 2387
rect 23506 2331 23530 2387
rect 23586 2331 23623 2387
rect 23413 2306 23623 2331
rect 23413 2250 23450 2306
rect 23506 2250 23530 2306
rect 23586 2250 23623 2306
rect 23413 2225 23623 2250
rect 23413 2169 23450 2225
rect 23506 2169 23530 2225
rect 23586 2169 23623 2225
rect 23413 2144 23623 2169
rect 23413 2088 23450 2144
rect 23506 2088 23530 2144
rect 23586 2088 23623 2144
rect 23413 2063 23623 2088
rect 23413 2007 23450 2063
rect 23506 2007 23530 2063
rect 23586 2007 23623 2063
rect 23413 1982 23623 2007
rect 23413 1926 23450 1982
rect 23506 1926 23530 1982
rect 23586 1926 23623 1982
rect 23413 1901 23623 1926
rect 23413 1845 23450 1901
rect 23506 1845 23530 1901
rect 23586 1845 23623 1901
rect 23413 1820 23623 1845
rect 23413 1764 23450 1820
rect 23506 1764 23530 1820
rect 23586 1764 23623 1820
rect 23413 1739 23623 1764
rect 23413 1683 23450 1739
rect 23506 1683 23530 1739
rect 23586 1683 23623 1739
rect 23413 1658 23623 1683
rect 23413 1602 23450 1658
rect 23506 1602 23530 1658
rect 23586 1602 23623 1658
rect 23413 1577 23623 1602
rect 23413 1521 23450 1577
rect 23506 1521 23530 1577
rect 23586 1521 23623 1577
rect 23413 1496 23623 1521
rect 23413 1440 23450 1496
rect 23506 1440 23530 1496
rect 23586 1440 23623 1496
rect 23413 1415 23623 1440
rect 23413 1359 23450 1415
rect 23506 1359 23530 1415
rect 23586 1359 23623 1415
rect 23413 -2873 23623 1359
tri 23822 235 23827 240 se
rect 23827 235 23867 14365
tri 23867 14349 23883 14365 nw
rect 24154 3190 24428 3204
rect 24154 2734 24182 3190
rect 24398 2734 24428 3190
rect 24154 2709 24428 2734
rect 24154 2653 24182 2709
rect 24238 2653 24262 2709
rect 24318 2653 24342 2709
rect 24398 2653 24428 2709
rect 24154 2628 24428 2653
rect 24154 2572 24182 2628
rect 24238 2572 24262 2628
rect 24318 2572 24342 2628
rect 24398 2572 24428 2628
rect 24154 2547 24428 2572
rect 24154 2491 24182 2547
rect 24238 2491 24262 2547
rect 24318 2491 24342 2547
rect 24398 2491 24428 2547
rect 24154 2466 24428 2491
rect 24154 2410 24182 2466
rect 24238 2410 24262 2466
rect 24318 2410 24342 2466
rect 24398 2410 24428 2466
rect 24154 2385 24428 2410
rect 24154 2329 24182 2385
rect 24238 2329 24262 2385
rect 24318 2329 24342 2385
rect 24398 2329 24428 2385
rect 24154 2304 24428 2329
rect 24154 2248 24182 2304
rect 24238 2248 24262 2304
rect 24318 2248 24342 2304
rect 24398 2248 24428 2304
rect 24154 2223 24428 2248
rect 24154 2167 24182 2223
rect 24238 2167 24262 2223
rect 24318 2167 24342 2223
rect 24398 2167 24428 2223
rect 24154 2142 24428 2167
rect 24154 2086 24182 2142
rect 24238 2086 24262 2142
rect 24318 2086 24342 2142
rect 24398 2086 24428 2142
rect 24154 2061 24428 2086
rect 24154 2005 24182 2061
rect 24238 2005 24262 2061
rect 24318 2005 24342 2061
rect 24398 2005 24428 2061
rect 24154 1980 24428 2005
rect 24154 1924 24182 1980
rect 24238 1924 24262 1980
rect 24318 1924 24342 1980
rect 24398 1924 24428 1980
rect 24154 1899 24428 1924
rect 24154 1843 24182 1899
rect 24238 1843 24262 1899
rect 24318 1843 24342 1899
rect 24398 1843 24428 1899
rect 24154 1818 24428 1843
rect 24154 1762 24182 1818
rect 24238 1762 24262 1818
rect 24318 1762 24342 1818
rect 24398 1762 24428 1818
rect 24154 1737 24428 1762
rect 24154 1681 24182 1737
rect 24238 1681 24262 1737
rect 24318 1681 24342 1737
rect 24398 1681 24428 1737
rect 24154 1656 24428 1681
rect 24154 1600 24182 1656
rect 24238 1600 24262 1656
rect 24318 1600 24342 1656
rect 24398 1600 24428 1656
rect 24154 1575 24428 1600
rect 24154 1519 24182 1575
rect 24238 1519 24262 1575
rect 24318 1519 24342 1575
rect 24398 1519 24428 1575
rect 24154 1494 24428 1519
rect 24154 1438 24182 1494
rect 24238 1438 24262 1494
rect 24318 1438 24342 1494
rect 24398 1438 24428 1494
rect 24154 1413 24428 1438
rect 24154 1357 24182 1413
rect 24238 1357 24262 1413
rect 24318 1357 24342 1413
rect 24398 1357 24428 1413
tri 23867 235 23874 242 sw
rect 23822 229 23874 235
rect 23822 165 23874 177
rect 23822 107 23874 113
rect 23413 -2929 23449 -2873
rect 23505 -2929 23529 -2873
rect 23585 -2929 23623 -2873
rect 23413 -2958 23623 -2929
rect 23413 -3014 23449 -2958
rect 23505 -3014 23529 -2958
rect 23585 -3014 23623 -2958
rect 23413 -3043 23623 -3014
rect 23413 -3099 23449 -3043
rect 23505 -3099 23529 -3043
rect 23585 -3099 23623 -3043
rect 23413 -3128 23623 -3099
rect 23413 -3184 23449 -3128
rect 23505 -3184 23529 -3128
rect 23585 -3184 23623 -3128
rect 23413 -3214 23623 -3184
rect 23413 -3270 23449 -3214
rect 23505 -3270 23529 -3214
rect 23585 -3270 23623 -3214
rect 23413 -3300 23623 -3270
rect 23413 -3356 23449 -3300
rect 23505 -3356 23529 -3300
rect 23585 -3356 23623 -3300
rect 23413 -3386 23623 -3356
rect 23413 -3442 23449 -3386
rect 23505 -3442 23529 -3386
rect 23585 -3442 23623 -3386
rect 23413 -3472 23623 -3442
rect 23413 -3528 23449 -3472
rect 23505 -3528 23529 -3472
rect 23585 -3528 23623 -3472
rect 23413 -3558 23623 -3528
rect 23413 -3614 23449 -3558
rect 23505 -3614 23529 -3558
rect 23585 -3614 23623 -3558
rect 23413 -3644 23623 -3614
rect 23413 -3700 23449 -3644
rect 23505 -3700 23529 -3644
rect 23585 -3700 23623 -3644
rect 23413 -3716 23623 -3700
rect 24154 -2871 24428 1357
rect 24154 -2927 24183 -2871
rect 24239 -2927 24263 -2871
rect 24319 -2927 24343 -2871
rect 24399 -2927 24428 -2871
rect 24154 -2957 24428 -2927
rect 24154 -3013 24183 -2957
rect 24239 -3013 24263 -2957
rect 24319 -3013 24343 -2957
rect 24399 -3013 24428 -2957
rect 25486 -2868 25538 15069
rect 31290 14732 31434 14867
rect 31514 14727 31642 14867
rect 31700 14727 31828 14867
rect 27578 4679 28008 4708
rect 27578 4623 27606 4679
rect 27662 4623 27686 4679
rect 27742 4623 27766 4679
rect 27822 4623 27846 4679
rect 27902 4623 27926 4679
rect 27982 4623 28008 4679
rect 27578 4598 28008 4623
rect 27578 4542 27606 4598
rect 27662 4542 27686 4598
rect 27742 4542 27766 4598
rect 27822 4542 27846 4598
rect 27902 4542 27926 4598
rect 27982 4542 28008 4598
rect 27578 4517 28008 4542
rect 27578 4461 27606 4517
rect 27662 4461 27686 4517
rect 27742 4461 27766 4517
rect 27822 4461 27846 4517
rect 27902 4461 27926 4517
rect 27982 4461 28008 4517
rect 27578 4435 28008 4461
rect 27578 4379 27606 4435
rect 27662 4379 27686 4435
rect 27742 4379 27766 4435
rect 27822 4379 27846 4435
rect 27902 4379 27926 4435
rect 27982 4379 28008 4435
rect 27578 4353 28008 4379
rect 27578 4297 27606 4353
rect 27662 4297 27686 4353
rect 27742 4297 27766 4353
rect 27822 4297 27846 4353
rect 27902 4297 27926 4353
rect 27982 4297 28008 4353
rect 27578 4271 28008 4297
rect 27578 4215 27606 4271
rect 27662 4215 27686 4271
rect 27742 4215 27766 4271
rect 27822 4215 27846 4271
rect 27902 4215 27926 4271
rect 27982 4215 28008 4271
rect 27578 4189 28008 4215
rect 27578 4133 27606 4189
rect 27662 4133 27686 4189
rect 27742 4133 27766 4189
rect 27822 4133 27846 4189
rect 27902 4133 27926 4189
rect 27982 4133 28008 4189
rect 27578 4107 28008 4133
rect 27578 4051 27606 4107
rect 27662 4051 27686 4107
rect 27742 4051 27766 4107
rect 27822 4051 27846 4107
rect 27902 4051 27926 4107
rect 27982 4051 28008 4107
rect 27578 4025 28008 4051
rect 27578 3969 27606 4025
rect 27662 3969 27686 4025
rect 27742 3969 27766 4025
rect 27822 3969 27846 4025
rect 27902 3969 27926 4025
rect 27982 3969 28008 4025
rect 27578 3943 28008 3969
rect 27578 3887 27606 3943
rect 27662 3887 27686 3943
rect 27742 3887 27766 3943
rect 27822 3887 27846 3943
rect 27902 3887 27926 3943
rect 27982 3887 28008 3943
rect 27578 3861 28008 3887
rect 27578 3805 27606 3861
rect 27662 3805 27686 3861
rect 27742 3805 27766 3861
rect 27822 3805 27846 3861
rect 27902 3805 27926 3861
rect 27982 3805 28008 3861
rect 27578 3779 28008 3805
rect 27578 3723 27606 3779
rect 27662 3723 27686 3779
rect 27742 3723 27766 3779
rect 27822 3723 27846 3779
rect 27902 3723 27926 3779
rect 27982 3723 28008 3779
rect 25486 -2932 25538 -2920
rect 25486 -2992 25538 -2984
rect 25875 2436 26397 2465
rect 25875 2380 25907 2436
rect 25963 2380 25987 2436
rect 26043 2380 26067 2436
rect 26123 2380 26147 2436
rect 26203 2380 26227 2436
rect 26283 2380 26307 2436
rect 26363 2380 26397 2436
rect 25875 2353 26397 2380
rect 25875 2297 25907 2353
rect 25963 2297 25987 2353
rect 26043 2297 26067 2353
rect 26123 2297 26147 2353
rect 26203 2297 26227 2353
rect 26283 2297 26307 2353
rect 26363 2297 26397 2353
rect 25875 2270 26397 2297
rect 25875 2214 25907 2270
rect 25963 2214 25987 2270
rect 26043 2214 26067 2270
rect 26123 2214 26147 2270
rect 26203 2214 26227 2270
rect 26283 2214 26307 2270
rect 26363 2214 26397 2270
rect 25875 2187 26397 2214
rect 25875 2131 25907 2187
rect 25963 2131 25987 2187
rect 26043 2131 26067 2187
rect 26123 2131 26147 2187
rect 26203 2131 26227 2187
rect 26283 2131 26307 2187
rect 26363 2131 26397 2187
rect 25875 2104 26397 2131
rect 25875 2048 25907 2104
rect 25963 2048 25987 2104
rect 26043 2048 26067 2104
rect 26123 2048 26147 2104
rect 26203 2048 26227 2104
rect 26283 2048 26307 2104
rect 26363 2048 26397 2104
rect 25875 2021 26397 2048
rect 25875 1965 25907 2021
rect 25963 1965 25987 2021
rect 26043 1965 26067 2021
rect 26123 1965 26147 2021
rect 26203 1965 26227 2021
rect 26283 1965 26307 2021
rect 26363 1965 26397 2021
rect 25875 1938 26397 1965
rect 25875 1882 25907 1938
rect 25963 1882 25987 1938
rect 26043 1882 26067 1938
rect 26123 1882 26147 1938
rect 26203 1882 26227 1938
rect 26283 1882 26307 1938
rect 26363 1882 26397 1938
rect 25875 1855 26397 1882
rect 25875 1799 25907 1855
rect 25963 1799 25987 1855
rect 26043 1799 26067 1855
rect 26123 1799 26147 1855
rect 26203 1799 26227 1855
rect 26283 1799 26307 1855
rect 26363 1799 26397 1855
rect 25875 1771 26397 1799
rect 25875 1715 25907 1771
rect 25963 1715 25987 1771
rect 26043 1715 26067 1771
rect 26123 1715 26147 1771
rect 26203 1715 26227 1771
rect 26283 1715 26307 1771
rect 26363 1715 26397 1771
rect 25875 1687 26397 1715
rect 25875 1631 25907 1687
rect 25963 1631 25987 1687
rect 26043 1631 26067 1687
rect 26123 1631 26147 1687
rect 26203 1631 26227 1687
rect 26283 1631 26307 1687
rect 26363 1631 26397 1687
rect 25875 1603 26397 1631
rect 25875 1547 25907 1603
rect 25963 1547 25987 1603
rect 26043 1547 26067 1603
rect 26123 1547 26147 1603
rect 26203 1547 26227 1603
rect 26283 1547 26307 1603
rect 26363 1547 26397 1603
rect 25875 1519 26397 1547
rect 25875 1463 25907 1519
rect 25963 1463 25987 1519
rect 26043 1463 26067 1519
rect 26123 1463 26147 1519
rect 26203 1463 26227 1519
rect 26283 1463 26307 1519
rect 26363 1463 26397 1519
rect 25875 1435 26397 1463
rect 25875 1379 25907 1435
rect 25963 1379 25987 1435
rect 26043 1379 26067 1435
rect 26123 1379 26147 1435
rect 26203 1379 26227 1435
rect 26283 1379 26307 1435
rect 26363 1379 26397 1435
rect 25875 -2198 26397 1379
rect 27578 822 28008 3723
rect 27578 766 27606 822
rect 27662 766 27686 822
rect 27742 766 27766 822
rect 27822 766 27846 822
rect 27902 766 27926 822
rect 27982 766 28008 822
rect 27578 741 28008 766
rect 27578 685 27606 741
rect 27662 685 27686 741
rect 27742 685 27766 741
rect 27822 685 27846 741
rect 27902 685 27926 741
rect 27982 685 28008 741
rect 27578 660 28008 685
rect 27578 604 27606 660
rect 27662 604 27686 660
rect 27742 604 27766 660
rect 27822 604 27846 660
rect 27902 604 27926 660
rect 27982 604 28008 660
rect 27578 579 28008 604
rect 27578 523 27606 579
rect 27662 523 27686 579
rect 27742 523 27766 579
rect 27822 523 27846 579
rect 27902 523 27926 579
rect 27982 523 28008 579
rect 27578 498 28008 523
rect 27578 442 27606 498
rect 27662 442 27686 498
rect 27742 442 27766 498
rect 27822 442 27846 498
rect 27902 442 27926 498
rect 27982 442 28008 498
rect 27578 417 28008 442
rect 27578 361 27606 417
rect 27662 361 27686 417
rect 27742 361 27766 417
rect 27822 361 27846 417
rect 27902 361 27926 417
rect 27982 361 28008 417
rect 27578 335 28008 361
rect 27578 279 27606 335
rect 27662 279 27686 335
rect 27742 279 27766 335
rect 27822 279 27846 335
rect 27902 279 27926 335
rect 27982 279 28008 335
rect 27578 253 28008 279
rect 27578 197 27606 253
rect 27662 197 27686 253
rect 27742 197 27766 253
rect 27822 197 27846 253
rect 27902 197 27926 253
rect 27982 197 28008 253
rect 27578 171 28008 197
rect 27578 115 27606 171
rect 27662 115 27686 171
rect 27742 115 27766 171
rect 27822 115 27846 171
rect 27902 115 27926 171
rect 27982 115 28008 171
rect 27578 89 28008 115
rect 27578 33 27606 89
rect 27662 33 27686 89
rect 27742 33 27766 89
rect 27822 33 27846 89
rect 27902 33 27926 89
rect 27982 33 28008 89
rect 27578 7 28008 33
rect 27578 -49 27606 7
rect 27662 -49 27686 7
rect 27742 -49 27766 7
rect 27822 -49 27846 7
rect 27902 -49 27926 7
rect 27982 -49 28008 7
rect 27578 -75 28008 -49
rect 27578 -131 27606 -75
rect 27662 -131 27686 -75
rect 27742 -131 27766 -75
rect 27822 -131 27846 -75
rect 27902 -131 27926 -75
rect 27982 -131 28008 -75
rect 27578 -157 28008 -131
rect 27578 -213 27606 -157
rect 27662 -213 27686 -157
rect 27742 -213 27766 -157
rect 27822 -213 27846 -157
rect 27902 -213 27926 -157
rect 27982 -213 28008 -157
rect 27578 -239 28008 -213
rect 27578 -295 27606 -239
rect 27662 -295 27686 -239
rect 27742 -295 27766 -239
rect 27822 -295 27846 -239
rect 27902 -295 27926 -239
rect 27982 -295 28008 -239
rect 27578 -321 28008 -295
rect 27578 -377 27606 -321
rect 27662 -377 27686 -321
rect 27742 -377 27766 -321
rect 27822 -377 27846 -321
rect 27902 -377 27926 -321
rect 27982 -377 28008 -321
rect 25875 -2689 26294 -2198
tri 26294 -2301 26397 -2198 nw
tri 26294 -2689 26397 -2586 sw
rect 25875 -2878 26397 -2689
rect 25875 -2934 25905 -2878
rect 25961 -2934 25985 -2878
rect 26041 -2934 26065 -2878
rect 26121 -2934 26145 -2878
rect 26201 -2934 26225 -2878
rect 26281 -2934 26305 -2878
rect 26361 -2934 26397 -2878
rect 25875 -2962 26397 -2934
rect 24154 -3043 24428 -3013
rect 24154 -3099 24183 -3043
rect 24239 -3099 24263 -3043
rect 24319 -3099 24343 -3043
rect 24399 -3099 24428 -3043
rect 24154 -3129 24428 -3099
rect 24154 -3185 24183 -3129
rect 24239 -3185 24263 -3129
rect 24319 -3185 24343 -3129
rect 24399 -3185 24428 -3129
rect 24154 -3215 24428 -3185
rect 24154 -3271 24183 -3215
rect 24239 -3271 24263 -3215
rect 24319 -3271 24343 -3215
rect 24399 -3271 24428 -3215
rect 24154 -3301 24428 -3271
rect 24154 -3357 24183 -3301
rect 24239 -3357 24263 -3301
rect 24319 -3357 24343 -3301
rect 24399 -3357 24428 -3301
rect 24154 -3387 24428 -3357
rect 24154 -3443 24183 -3387
rect 24239 -3443 24263 -3387
rect 24319 -3443 24343 -3387
rect 24399 -3443 24428 -3387
rect 24154 -3473 24428 -3443
rect 24154 -3529 24183 -3473
rect 24239 -3529 24263 -3473
rect 24319 -3529 24343 -3473
rect 24399 -3529 24428 -3473
rect 24154 -3559 24428 -3529
rect 24154 -3615 24183 -3559
rect 24239 -3615 24263 -3559
rect 24319 -3615 24343 -3559
rect 24399 -3615 24428 -3559
rect 24154 -3646 24428 -3615
rect 24154 -3702 24183 -3646
rect 24239 -3702 24263 -3646
rect 24319 -3702 24343 -3646
rect 24399 -3702 24428 -3646
rect 24154 -3716 24428 -3702
rect 25875 -3018 25905 -2962
rect 25961 -3018 25985 -2962
rect 26041 -3018 26065 -2962
rect 26121 -3018 26145 -2962
rect 26201 -3018 26225 -2962
rect 26281 -3018 26305 -2962
rect 26361 -3018 26397 -2962
rect 25875 -3046 26397 -3018
rect 25875 -3102 25905 -3046
rect 25961 -3102 25985 -3046
rect 26041 -3102 26065 -3046
rect 26121 -3102 26145 -3046
rect 26201 -3102 26225 -3046
rect 26281 -3102 26305 -3046
rect 26361 -3102 26397 -3046
rect 25875 -3131 26397 -3102
rect 25875 -3187 25905 -3131
rect 25961 -3187 25985 -3131
rect 26041 -3187 26065 -3131
rect 26121 -3187 26145 -3131
rect 26201 -3187 26225 -3131
rect 26281 -3187 26305 -3131
rect 26361 -3187 26397 -3131
rect 25875 -3216 26397 -3187
rect 25875 -3272 25905 -3216
rect 25961 -3272 25985 -3216
rect 26041 -3272 26065 -3216
rect 26121 -3272 26145 -3216
rect 26201 -3272 26225 -3216
rect 26281 -3272 26305 -3216
rect 26361 -3272 26397 -3216
rect 25875 -3301 26397 -3272
rect 25875 -3357 25905 -3301
rect 25961 -3357 25985 -3301
rect 26041 -3357 26065 -3301
rect 26121 -3357 26145 -3301
rect 26201 -3357 26225 -3301
rect 26281 -3357 26305 -3301
rect 26361 -3357 26397 -3301
rect 25875 -3386 26397 -3357
rect 25875 -3442 25905 -3386
rect 25961 -3442 25985 -3386
rect 26041 -3442 26065 -3386
rect 26121 -3442 26145 -3386
rect 26201 -3442 26225 -3386
rect 26281 -3442 26305 -3386
rect 26361 -3442 26397 -3386
rect 25875 -3471 26397 -3442
rect 25875 -3527 25905 -3471
rect 25961 -3527 25985 -3471
rect 26041 -3527 26065 -3471
rect 26121 -3527 26145 -3471
rect 26201 -3527 26225 -3471
rect 26281 -3527 26305 -3471
rect 26361 -3527 26397 -3471
rect 25875 -3556 26397 -3527
rect 25875 -3612 25905 -3556
rect 25961 -3612 25985 -3556
rect 26041 -3612 26065 -3556
rect 26121 -3612 26145 -3556
rect 26201 -3612 26225 -3556
rect 26281 -3612 26305 -3556
rect 26361 -3612 26397 -3556
rect 25875 -3641 26397 -3612
rect 25875 -3697 25905 -3641
rect 25961 -3697 25985 -3641
rect 26041 -3697 26065 -3641
rect 26121 -3697 26145 -3641
rect 26201 -3697 26225 -3641
rect 26281 -3697 26305 -3641
rect 26361 -3697 26397 -3641
rect 25875 -3714 26397 -3697
tri 21843 -4060 22094 -3809 sw
rect 21538 -4231 22094 -4060
rect 21538 -4287 21547 -4231
rect 21603 -4287 21627 -4231
rect 21683 -4287 21707 -4231
rect 21763 -4287 21787 -4231
rect 21843 -4287 21867 -4231
rect 21923 -4287 21947 -4231
rect 22003 -4287 22027 -4231
rect 22083 -4287 22094 -4231
rect 21538 -4321 22094 -4287
rect 21538 -4377 21547 -4321
rect 21603 -4377 21627 -4321
rect 21683 -4377 21707 -4321
rect 21763 -4377 21787 -4321
rect 21843 -4377 21867 -4321
rect 21923 -4377 21947 -4321
rect 22003 -4377 22027 -4321
rect 22083 -4377 22094 -4321
rect 21538 -4411 22094 -4377
rect 21538 -4467 21547 -4411
rect 21603 -4467 21627 -4411
rect 21683 -4467 21707 -4411
rect 21763 -4467 21787 -4411
rect 21843 -4467 21867 -4411
rect 21923 -4467 21947 -4411
rect 22003 -4467 22027 -4411
rect 22083 -4467 22094 -4411
rect 21538 -4502 22094 -4467
rect 21538 -4558 21547 -4502
rect 21603 -4558 21627 -4502
rect 21683 -4558 21707 -4502
rect 21763 -4558 21787 -4502
rect 21843 -4558 21867 -4502
rect 21923 -4558 21947 -4502
rect 22003 -4558 22027 -4502
rect 22083 -4558 22094 -4502
rect 21538 -4593 22094 -4558
rect 21538 -4649 21547 -4593
rect 21603 -4649 21627 -4593
rect 21683 -4649 21707 -4593
rect 21763 -4649 21787 -4593
rect 21843 -4649 21867 -4593
rect 21923 -4649 21947 -4593
rect 22003 -4649 22027 -4593
rect 22083 -4649 22094 -4593
rect 21538 -4684 22094 -4649
rect 21538 -4740 21547 -4684
rect 21603 -4740 21627 -4684
rect 21683 -4740 21707 -4684
rect 21763 -4740 21787 -4684
rect 21843 -4740 21867 -4684
rect 21923 -4740 21947 -4684
rect 22003 -4740 22027 -4684
rect 22083 -4740 22094 -4684
rect 21538 -4775 22094 -4740
rect 21538 -4831 21547 -4775
rect 21603 -4831 21627 -4775
rect 21683 -4831 21707 -4775
rect 21763 -4831 21787 -4775
rect 21843 -4831 21867 -4775
rect 21923 -4831 21947 -4775
rect 22003 -4831 22027 -4775
rect 22083 -4831 22094 -4775
rect 21538 -4840 22094 -4831
rect 22204 -5069 22725 -3800
rect 26659 -5046 26687 -388
rect 27578 -403 28008 -377
rect 27578 -459 27606 -403
rect 27662 -459 27686 -403
rect 27742 -459 27766 -403
rect 27822 -459 27846 -403
rect 27902 -459 27926 -403
rect 27982 -459 28008 -403
rect 27578 -494 28008 -459
rect 28302 4685 28682 4708
rect 28302 4629 28345 4685
rect 28401 4629 28425 4685
rect 28481 4629 28505 4685
rect 28561 4629 28585 4685
rect 28641 4629 28682 4685
rect 28302 4603 28682 4629
rect 28302 4547 28345 4603
rect 28401 4547 28425 4603
rect 28481 4547 28505 4603
rect 28561 4547 28585 4603
rect 28641 4547 28682 4603
rect 28302 4521 28682 4547
rect 28302 4465 28345 4521
rect 28401 4465 28425 4521
rect 28481 4465 28505 4521
rect 28561 4465 28585 4521
rect 28641 4465 28682 4521
rect 28302 4439 28682 4465
rect 28302 4383 28345 4439
rect 28401 4383 28425 4439
rect 28481 4383 28505 4439
rect 28561 4383 28585 4439
rect 28641 4383 28682 4439
rect 28302 4357 28682 4383
rect 28302 4301 28345 4357
rect 28401 4301 28425 4357
rect 28481 4301 28505 4357
rect 28561 4301 28585 4357
rect 28641 4301 28682 4357
rect 28302 4275 28682 4301
rect 28302 4219 28345 4275
rect 28401 4219 28425 4275
rect 28481 4219 28505 4275
rect 28561 4219 28585 4275
rect 28641 4219 28682 4275
rect 28302 4193 28682 4219
rect 28302 4137 28345 4193
rect 28401 4137 28425 4193
rect 28481 4137 28505 4193
rect 28561 4137 28585 4193
rect 28641 4137 28682 4193
rect 28302 4111 28682 4137
rect 28302 4055 28345 4111
rect 28401 4055 28425 4111
rect 28481 4055 28505 4111
rect 28561 4055 28585 4111
rect 28641 4055 28682 4111
rect 28302 4028 28682 4055
rect 28302 3972 28345 4028
rect 28401 3972 28425 4028
rect 28481 3972 28505 4028
rect 28561 3972 28585 4028
rect 28641 3972 28682 4028
rect 28302 3945 28682 3972
rect 28302 3889 28345 3945
rect 28401 3889 28425 3945
rect 28481 3889 28505 3945
rect 28561 3889 28585 3945
rect 28641 3889 28682 3945
rect 28302 3862 28682 3889
rect 28302 3806 28345 3862
rect 28401 3806 28425 3862
rect 28481 3806 28505 3862
rect 28561 3806 28585 3862
rect 28641 3806 28682 3862
rect 28302 3779 28682 3806
rect 28302 3723 28345 3779
rect 28401 3723 28425 3779
rect 28481 3723 28505 3779
rect 28561 3723 28585 3779
rect 28641 3723 28682 3779
rect 28302 806 28682 3723
rect 28302 270 28345 806
rect 28641 270 28682 806
rect 28302 245 28682 270
rect 28302 189 28345 245
rect 28401 189 28425 245
rect 28481 189 28505 245
rect 28561 189 28585 245
rect 28641 189 28682 245
rect 28302 164 28682 189
rect 28302 108 28345 164
rect 28401 108 28425 164
rect 28481 108 28505 164
rect 28561 108 28585 164
rect 28641 108 28682 164
rect 28302 83 28682 108
rect 28302 27 28345 83
rect 28401 27 28425 83
rect 28481 27 28505 83
rect 28561 27 28585 83
rect 28641 27 28682 83
rect 28302 2 28682 27
rect 28302 -54 28345 2
rect 28401 -54 28425 2
rect 28481 -54 28505 2
rect 28561 -54 28585 2
rect 28641 -54 28682 2
rect 28302 -79 28682 -54
rect 28302 -135 28345 -79
rect 28401 -135 28425 -79
rect 28481 -135 28505 -79
rect 28561 -135 28585 -79
rect 28641 -135 28682 -79
rect 28302 -160 28682 -135
rect 28302 -216 28345 -160
rect 28401 -216 28425 -160
rect 28481 -216 28505 -160
rect 28561 -216 28585 -160
rect 28641 -216 28682 -160
rect 28302 -241 28682 -216
rect 28302 -297 28345 -241
rect 28401 -297 28425 -241
rect 28481 -297 28505 -241
rect 28561 -297 28585 -241
rect 28641 -297 28682 -241
rect 28302 -322 28682 -297
rect 28302 -378 28345 -322
rect 28401 -378 28425 -322
rect 28481 -378 28505 -322
rect 28561 -378 28585 -322
rect 28641 -378 28682 -322
rect 28302 -403 28682 -378
rect 28302 -459 28345 -403
rect 28401 -459 28425 -403
rect 28481 -459 28505 -403
rect 28561 -459 28585 -403
rect 28641 -459 28682 -403
rect 28302 -494 28682 -459
tri 22615 -5179 22725 -5069 nw
rect 17714 -6078 18524 -6062
rect 19925 -6078 20750 -6062
rect 22204 -6078 22615 -6068
rect 22753 -6078 22945 -6068
rect 23241 -6078 23293 -6008
rect 23393 -6078 23844 -6068
rect 23934 -6078 24126 -6068
rect 24516 -6078 24698 -6068
rect 24754 -6078 25461 -6068
rect 25519 -6078 25658 -6068
rect 25947 -6078 26360 -6068
rect 26818 -6078 27267 -6068
rect 28391 -6096 28865 -6068
rect 28978 -6096 29298 -6068
rect 31477 -6096 31828 -6068
<< via2 >>
rect 19263 22245 19319 22257
rect 19357 22245 19413 22257
rect 19450 22245 19506 22257
rect 19543 22245 19599 22257
rect 19636 22245 19692 22257
rect 19729 22245 19785 22257
rect 19822 22245 19878 22257
rect 19263 22201 19271 22245
rect 19271 22201 19319 22245
rect 19357 22201 19393 22245
rect 19393 22201 19411 22245
rect 19411 22201 19413 22245
rect 19450 22201 19463 22245
rect 19463 22201 19480 22245
rect 19480 22201 19506 22245
rect 19543 22201 19549 22245
rect 19549 22201 19599 22245
rect 19636 22201 19670 22245
rect 19670 22201 19687 22245
rect 19687 22201 19692 22245
rect 19729 22201 19739 22245
rect 19739 22201 19756 22245
rect 19756 22201 19785 22245
rect 19822 22201 19825 22245
rect 19825 22201 19877 22245
rect 19877 22201 19878 22245
rect 19263 22129 19271 22177
rect 19271 22129 19319 22177
rect 19357 22129 19393 22177
rect 19393 22129 19411 22177
rect 19411 22129 19413 22177
rect 19450 22129 19463 22177
rect 19463 22129 19480 22177
rect 19480 22129 19506 22177
rect 19543 22129 19549 22177
rect 19549 22129 19599 22177
rect 19636 22129 19670 22177
rect 19670 22129 19687 22177
rect 19687 22129 19692 22177
rect 19729 22129 19739 22177
rect 19739 22129 19756 22177
rect 19756 22129 19785 22177
rect 19822 22129 19825 22177
rect 19825 22129 19877 22177
rect 19877 22129 19878 22177
rect 19263 22121 19319 22129
rect 19357 22121 19413 22129
rect 19450 22121 19506 22129
rect 19543 22121 19599 22129
rect 19636 22121 19692 22129
rect 19729 22121 19785 22129
rect 19822 22121 19878 22129
rect 19217 18782 19273 18807
rect 19298 18782 19354 18807
rect 19379 18782 19435 18807
rect 19460 18782 19516 18807
rect 19541 18782 19597 18807
rect 19622 18782 19678 18807
rect 19703 18782 19759 18807
rect 19784 18782 19840 18807
rect 19865 18782 20561 18807
rect 19217 18751 19227 18782
rect 19227 18751 19273 18782
rect 19298 18751 19346 18782
rect 19346 18751 19354 18782
rect 19379 18751 19413 18782
rect 19413 18751 19428 18782
rect 19428 18751 19435 18782
rect 19460 18751 19480 18782
rect 19480 18751 19495 18782
rect 19495 18751 19516 18782
rect 19541 18751 19547 18782
rect 19547 18751 19562 18782
rect 19562 18751 19597 18782
rect 19622 18751 19629 18782
rect 19629 18751 19678 18782
rect 19703 18751 19748 18782
rect 19748 18751 19759 18782
rect 19784 18751 19815 18782
rect 19815 18751 19830 18782
rect 19830 18751 19840 18782
rect 19865 18730 19882 18782
rect 19882 18730 19897 18782
rect 19897 18730 19949 18782
rect 19949 18730 19964 18782
rect 19964 18730 20016 18782
rect 20016 18730 20031 18782
rect 20031 18730 20083 18782
rect 20083 18730 20098 18782
rect 20098 18730 20150 18782
rect 20150 18730 20165 18782
rect 20165 18730 20217 18782
rect 20217 18730 20232 18782
rect 20232 18730 20284 18782
rect 20284 18730 20299 18782
rect 20299 18730 20351 18782
rect 20351 18730 20366 18782
rect 20366 18730 20418 18782
rect 20418 18730 20433 18782
rect 20433 18730 20485 18782
rect 20485 18730 20500 18782
rect 20500 18730 20552 18782
rect 20552 18730 20561 18782
rect 19217 18718 19273 18727
rect 19298 18718 19354 18727
rect 19379 18718 19435 18727
rect 19460 18718 19516 18727
rect 19541 18718 19597 18727
rect 19622 18718 19678 18727
rect 19703 18718 19759 18727
rect 19784 18718 19840 18727
rect 19865 18718 20561 18730
rect 19217 18671 19227 18718
rect 19227 18671 19273 18718
rect 19298 18671 19346 18718
rect 19346 18671 19354 18718
rect 19379 18671 19413 18718
rect 19413 18671 19428 18718
rect 19428 18671 19435 18718
rect 19460 18671 19480 18718
rect 19480 18671 19495 18718
rect 19495 18671 19516 18718
rect 19541 18671 19547 18718
rect 19547 18671 19562 18718
rect 19562 18671 19597 18718
rect 19622 18671 19629 18718
rect 19629 18671 19678 18718
rect 19703 18671 19748 18718
rect 19748 18671 19759 18718
rect 19784 18671 19815 18718
rect 19815 18671 19830 18718
rect 19830 18671 19840 18718
rect 19865 18666 19882 18718
rect 19882 18666 19897 18718
rect 19897 18666 19949 18718
rect 19949 18666 19964 18718
rect 19964 18666 20016 18718
rect 20016 18666 20031 18718
rect 20031 18666 20083 18718
rect 20083 18666 20098 18718
rect 20098 18666 20150 18718
rect 20150 18666 20165 18718
rect 20165 18666 20217 18718
rect 20217 18666 20232 18718
rect 20232 18666 20284 18718
rect 20284 18666 20299 18718
rect 20299 18666 20351 18718
rect 20351 18666 20366 18718
rect 20366 18666 20418 18718
rect 20418 18666 20433 18718
rect 20433 18666 20485 18718
rect 20485 18666 20500 18718
rect 20500 18666 20552 18718
rect 20552 18666 20561 18718
rect 19865 18654 20561 18666
rect 19217 18602 19227 18647
rect 19227 18602 19273 18647
rect 19298 18602 19346 18647
rect 19346 18602 19354 18647
rect 19379 18602 19413 18647
rect 19413 18602 19428 18647
rect 19428 18602 19435 18647
rect 19460 18602 19480 18647
rect 19480 18602 19495 18647
rect 19495 18602 19516 18647
rect 19541 18602 19547 18647
rect 19547 18602 19562 18647
rect 19562 18602 19597 18647
rect 19622 18602 19629 18647
rect 19629 18602 19678 18647
rect 19703 18602 19748 18647
rect 19748 18602 19759 18647
rect 19784 18602 19815 18647
rect 19815 18602 19830 18647
rect 19830 18602 19840 18647
rect 19865 18602 19882 18654
rect 19882 18602 19897 18654
rect 19897 18602 19949 18654
rect 19949 18602 19964 18654
rect 19964 18602 20016 18654
rect 20016 18602 20031 18654
rect 20031 18602 20083 18654
rect 20083 18602 20098 18654
rect 20098 18602 20150 18654
rect 20150 18602 20165 18654
rect 20165 18602 20217 18654
rect 20217 18602 20232 18654
rect 20232 18602 20284 18654
rect 20284 18602 20299 18654
rect 20299 18602 20351 18654
rect 20351 18602 20366 18654
rect 20366 18602 20418 18654
rect 20418 18602 20433 18654
rect 20433 18602 20485 18654
rect 20485 18602 20500 18654
rect 20500 18602 20552 18654
rect 20552 18602 20561 18654
rect 19217 18591 19273 18602
rect 19298 18591 19354 18602
rect 19379 18591 19435 18602
rect 19460 18591 19516 18602
rect 19541 18591 19597 18602
rect 19622 18591 19678 18602
rect 19703 18591 19759 18602
rect 19784 18591 19840 18602
rect 19865 18590 20561 18602
rect 19217 18538 19227 18567
rect 19227 18538 19273 18567
rect 19298 18538 19346 18567
rect 19346 18538 19354 18567
rect 19379 18538 19413 18567
rect 19413 18538 19428 18567
rect 19428 18538 19435 18567
rect 19460 18538 19480 18567
rect 19480 18538 19495 18567
rect 19495 18538 19516 18567
rect 19541 18538 19547 18567
rect 19547 18538 19562 18567
rect 19562 18538 19597 18567
rect 19622 18538 19629 18567
rect 19629 18538 19678 18567
rect 19703 18538 19748 18567
rect 19748 18538 19759 18567
rect 19784 18538 19815 18567
rect 19815 18538 19830 18567
rect 19830 18538 19840 18567
rect 19865 18538 19882 18590
rect 19882 18538 19897 18590
rect 19897 18538 19949 18590
rect 19949 18538 19964 18590
rect 19964 18538 20016 18590
rect 20016 18538 20031 18590
rect 20031 18538 20083 18590
rect 20083 18538 20098 18590
rect 20098 18538 20150 18590
rect 20150 18538 20165 18590
rect 20165 18538 20217 18590
rect 20217 18538 20232 18590
rect 20232 18538 20284 18590
rect 20284 18538 20299 18590
rect 20299 18538 20351 18590
rect 20351 18538 20366 18590
rect 20366 18538 20418 18590
rect 20418 18538 20433 18590
rect 20433 18538 20485 18590
rect 20485 18538 20500 18590
rect 20500 18538 20552 18590
rect 20552 18538 20561 18590
rect 19217 18511 19273 18538
rect 19298 18511 19354 18538
rect 19379 18511 19435 18538
rect 19460 18511 19516 18538
rect 19541 18511 19597 18538
rect 19622 18511 19678 18538
rect 19703 18511 19759 18538
rect 19784 18511 19840 18538
rect 19865 18511 20561 18538
rect 21011 22245 21067 22258
rect 21100 22245 21156 22258
rect 21189 22245 21245 22258
rect 21278 22245 21334 22258
rect 21367 22245 21423 22258
rect 21456 22245 21512 22258
rect 21545 22245 21601 22258
rect 21633 22245 21689 22258
rect 21721 22245 21777 22258
rect 21809 22245 21865 22258
rect 21011 22202 21012 22245
rect 21012 22202 21064 22245
rect 21064 22202 21067 22245
rect 21100 22202 21131 22245
rect 21131 22202 21146 22245
rect 21146 22202 21156 22245
rect 21189 22202 21198 22245
rect 21198 22202 21213 22245
rect 21213 22202 21245 22245
rect 21278 22202 21280 22245
rect 21280 22202 21332 22245
rect 21332 22202 21334 22245
rect 21367 22202 21399 22245
rect 21399 22202 21414 22245
rect 21414 22202 21423 22245
rect 21456 22202 21466 22245
rect 21466 22202 21481 22245
rect 21481 22202 21512 22245
rect 21545 22202 21548 22245
rect 21548 22202 21600 22245
rect 21600 22202 21601 22245
rect 21633 22202 21667 22245
rect 21667 22202 21681 22245
rect 21681 22202 21689 22245
rect 21721 22202 21733 22245
rect 21733 22202 21747 22245
rect 21747 22202 21777 22245
rect 21809 22202 21813 22245
rect 21813 22202 21865 22245
rect 21011 22129 21012 22178
rect 21012 22129 21064 22178
rect 21064 22129 21067 22178
rect 21100 22129 21131 22178
rect 21131 22129 21146 22178
rect 21146 22129 21156 22178
rect 21189 22129 21198 22178
rect 21198 22129 21213 22178
rect 21213 22129 21245 22178
rect 21278 22129 21280 22178
rect 21280 22129 21332 22178
rect 21332 22129 21334 22178
rect 21367 22129 21399 22178
rect 21399 22129 21414 22178
rect 21414 22129 21423 22178
rect 21456 22129 21466 22178
rect 21466 22129 21481 22178
rect 21481 22129 21512 22178
rect 21545 22129 21548 22178
rect 21548 22129 21600 22178
rect 21600 22129 21601 22178
rect 21633 22129 21667 22178
rect 21667 22129 21681 22178
rect 21681 22129 21689 22178
rect 21721 22129 21733 22178
rect 21733 22129 21747 22178
rect 21747 22129 21777 22178
rect 21809 22129 21813 22178
rect 21813 22129 21865 22178
rect 21011 22122 21067 22129
rect 21100 22122 21156 22129
rect 21189 22122 21245 22129
rect 21278 22122 21334 22129
rect 21367 22122 21423 22129
rect 21456 22122 21512 22129
rect 21545 22122 21601 22129
rect 21633 22122 21689 22129
rect 21721 22122 21777 22129
rect 21809 22122 21865 22129
rect 21048 18781 21104 18807
rect 21136 18781 21192 18807
rect 21224 18781 21280 18807
rect 21311 18781 21367 18807
rect 21398 18781 21454 18807
rect 21485 18781 21541 18807
rect 21572 18781 21628 18807
rect 21659 18781 21715 18807
rect 21048 18751 21100 18781
rect 21100 18751 21104 18781
rect 21136 18751 21169 18781
rect 21169 18751 21186 18781
rect 21186 18751 21192 18781
rect 21224 18751 21238 18781
rect 21238 18751 21254 18781
rect 21254 18751 21280 18781
rect 21311 18751 21322 18781
rect 21322 18751 21367 18781
rect 21398 18751 21442 18781
rect 21442 18751 21454 18781
rect 21485 18751 21510 18781
rect 21510 18751 21526 18781
rect 21526 18751 21541 18781
rect 21572 18751 21578 18781
rect 21578 18751 21594 18781
rect 21594 18751 21628 18781
rect 21659 18751 21662 18781
rect 21662 18751 21714 18781
rect 21714 18751 21715 18781
rect 21048 18717 21104 18727
rect 21136 18717 21192 18727
rect 21224 18717 21280 18727
rect 21311 18717 21367 18727
rect 21398 18717 21454 18727
rect 21485 18717 21541 18727
rect 21572 18717 21628 18727
rect 21659 18717 21715 18727
rect 21048 18671 21100 18717
rect 21100 18671 21104 18717
rect 21136 18671 21169 18717
rect 21169 18671 21186 18717
rect 21186 18671 21192 18717
rect 21224 18671 21238 18717
rect 21238 18671 21254 18717
rect 21254 18671 21280 18717
rect 21311 18671 21322 18717
rect 21322 18671 21367 18717
rect 21398 18671 21442 18717
rect 21442 18671 21454 18717
rect 21485 18671 21510 18717
rect 21510 18671 21526 18717
rect 21526 18671 21541 18717
rect 21572 18671 21578 18717
rect 21578 18671 21594 18717
rect 21594 18671 21628 18717
rect 21659 18671 21662 18717
rect 21662 18671 21714 18717
rect 21714 18671 21715 18717
rect 24092 18746 24148 18802
rect 24172 18746 24228 18802
rect 24252 18746 24308 18802
rect 21048 18601 21100 18647
rect 21100 18601 21104 18647
rect 21136 18601 21169 18647
rect 21169 18601 21186 18647
rect 21186 18601 21192 18647
rect 21224 18601 21238 18647
rect 21238 18601 21254 18647
rect 21254 18601 21280 18647
rect 21311 18601 21322 18647
rect 21322 18601 21367 18647
rect 21398 18601 21442 18647
rect 21442 18601 21454 18647
rect 21485 18601 21510 18647
rect 21510 18601 21526 18647
rect 21526 18601 21541 18647
rect 21572 18601 21578 18647
rect 21578 18601 21594 18647
rect 21594 18601 21628 18647
rect 21659 18601 21662 18647
rect 21662 18601 21714 18647
rect 21714 18601 21715 18647
rect 21048 18591 21104 18601
rect 21136 18591 21192 18601
rect 21224 18591 21280 18601
rect 21311 18591 21367 18601
rect 21398 18591 21454 18601
rect 21485 18591 21541 18601
rect 21572 18591 21628 18601
rect 21659 18591 21715 18601
rect 24092 18633 24148 18689
rect 24172 18633 24228 18689
rect 24252 18633 24308 18689
rect 21048 18537 21100 18567
rect 21100 18537 21104 18567
rect 21136 18537 21169 18567
rect 21169 18537 21186 18567
rect 21186 18537 21192 18567
rect 21224 18537 21238 18567
rect 21238 18537 21254 18567
rect 21254 18537 21280 18567
rect 21311 18537 21322 18567
rect 21322 18537 21367 18567
rect 21398 18537 21442 18567
rect 21442 18537 21454 18567
rect 21485 18537 21510 18567
rect 21510 18537 21526 18567
rect 21526 18537 21541 18567
rect 21572 18537 21578 18567
rect 21578 18537 21594 18567
rect 21594 18537 21628 18567
rect 21659 18537 21662 18567
rect 21662 18537 21714 18567
rect 21714 18537 21715 18567
rect 21048 18511 21104 18537
rect 21136 18511 21192 18537
rect 21224 18511 21280 18537
rect 21311 18511 21367 18537
rect 21398 18511 21454 18537
rect 21485 18511 21541 18537
rect 21572 18511 21628 18537
rect 21659 18511 21715 18537
rect 24092 18519 24148 18575
rect 24172 18519 24228 18575
rect 24252 18519 24308 18575
rect 29488 18735 29544 18791
rect 29568 18735 29624 18791
rect 29648 18735 29704 18791
rect 29728 18735 29784 18791
rect 29488 18649 29544 18705
rect 29568 18649 29624 18705
rect 29648 18649 29704 18705
rect 29728 18649 29784 18705
rect 29488 18562 29544 18618
rect 29568 18562 29624 18618
rect 29648 18562 29704 18618
rect 29728 18562 29784 18618
rect 29488 18475 29544 18531
rect 29568 18475 29624 18531
rect 29648 18475 29704 18531
rect 29728 18475 29784 18531
rect 29488 18388 29544 18444
rect 29568 18388 29624 18444
rect 29648 18388 29704 18444
rect 29728 18388 29784 18444
rect 29488 18301 29544 18357
rect 29568 18301 29624 18357
rect 29648 18301 29704 18357
rect 29728 18301 29784 18357
rect 29488 18214 29544 18270
rect 29568 18214 29624 18270
rect 29648 18214 29704 18270
rect 29728 18214 29784 18270
rect 29488 18127 29544 18183
rect 29568 18127 29624 18183
rect 29648 18127 29704 18183
rect 29728 18127 29784 18183
rect 29488 18040 29544 18096
rect 29568 18040 29624 18096
rect 29648 18040 29704 18096
rect 29728 18040 29784 18096
rect 19471 14719 19527 14775
rect 19551 14719 19607 14775
rect 19631 14719 19687 14775
rect 19711 14719 19767 14775
rect 19791 14719 19847 14775
rect 19471 14638 19527 14694
rect 19551 14638 19607 14694
rect 19631 14638 19687 14694
rect 19711 14638 19767 14694
rect 19791 14638 19847 14694
rect 19471 14557 19527 14613
rect 19551 14557 19607 14613
rect 19631 14557 19687 14613
rect 19711 14557 19767 14613
rect 19791 14557 19847 14613
rect 19471 14476 19527 14532
rect 19551 14476 19607 14532
rect 19631 14476 19687 14532
rect 19711 14476 19767 14532
rect 19791 14476 19847 14532
rect 19471 14395 19527 14451
rect 19551 14395 19607 14451
rect 19631 14395 19687 14451
rect 19711 14395 19767 14451
rect 19791 14395 19847 14451
rect 19471 14314 19527 14370
rect 19551 14314 19607 14370
rect 19631 14314 19687 14370
rect 19711 14314 19767 14370
rect 19791 14314 19847 14370
rect 19471 14233 19527 14289
rect 19551 14233 19607 14289
rect 19631 14233 19687 14289
rect 19711 14233 19767 14289
rect 19791 14233 19847 14289
rect 19471 14152 19527 14208
rect 19551 14152 19607 14208
rect 19631 14152 19687 14208
rect 19711 14152 19767 14208
rect 19791 14152 19847 14208
rect 19471 14071 19527 14127
rect 19551 14071 19607 14127
rect 19631 14071 19687 14127
rect 19711 14071 19767 14127
rect 19791 14071 19847 14127
rect 19471 13990 19527 14046
rect 19551 13990 19607 14046
rect 19631 13990 19687 14046
rect 19711 13990 19767 14046
rect 19791 13990 19847 14046
rect 19471 13909 19527 13965
rect 19551 13909 19607 13965
rect 19631 13909 19687 13965
rect 19711 13909 19767 13965
rect 19791 13909 19847 13965
rect 19471 13828 19527 13884
rect 19551 13828 19607 13884
rect 19631 13828 19687 13884
rect 19711 13828 19767 13884
rect 19791 13828 19847 13884
rect 19471 13747 19527 13803
rect 19551 13747 19607 13803
rect 19631 13747 19687 13803
rect 19711 13747 19767 13803
rect 19791 13747 19847 13803
rect 19471 13666 19527 13722
rect 19551 13666 19607 13722
rect 19631 13666 19687 13722
rect 19711 13666 19767 13722
rect 19791 13666 19847 13722
rect 19471 13585 19527 13641
rect 19551 13585 19607 13641
rect 19631 13585 19687 13641
rect 19711 13585 19767 13641
rect 19791 13585 19847 13641
rect 19471 13504 19527 13560
rect 19551 13504 19607 13560
rect 19631 13504 19687 13560
rect 19711 13504 19767 13560
rect 19791 13504 19847 13560
rect 19471 13423 19527 13479
rect 19551 13423 19607 13479
rect 19631 13423 19687 13479
rect 19711 13423 19767 13479
rect 19791 13423 19847 13479
rect 19471 13342 19527 13398
rect 19551 13342 19607 13398
rect 19631 13342 19687 13398
rect 19711 13342 19767 13398
rect 19791 13342 19847 13398
rect 19471 13261 19527 13317
rect 19551 13261 19607 13317
rect 19631 13261 19687 13317
rect 19711 13261 19767 13317
rect 19791 13261 19847 13317
rect 19471 13180 19527 13236
rect 19551 13180 19607 13236
rect 19631 13180 19687 13236
rect 19711 13180 19767 13236
rect 19791 13180 19847 13236
rect 19471 13099 19527 13155
rect 19551 13099 19607 13155
rect 19631 13099 19687 13155
rect 19711 13099 19767 13155
rect 19791 13099 19847 13155
rect 19471 13018 19527 13074
rect 19551 13018 19607 13074
rect 19631 13018 19687 13074
rect 19711 13018 19767 13074
rect 19791 13018 19847 13074
rect 19471 12937 19527 12993
rect 19551 12937 19607 12993
rect 19631 12937 19687 12993
rect 19711 12937 19767 12993
rect 19791 12937 19847 12993
rect 19471 12856 19527 12912
rect 19551 12856 19607 12912
rect 19631 12856 19687 12912
rect 19711 12856 19767 12912
rect 19791 12856 19847 12912
rect 19471 12775 19527 12831
rect 19551 12775 19607 12831
rect 19631 12775 19687 12831
rect 19711 12775 19767 12831
rect 19791 12775 19847 12831
rect 19471 12694 19527 12750
rect 19551 12694 19607 12750
rect 19631 12694 19687 12750
rect 19711 12694 19767 12750
rect 19791 12694 19847 12750
rect 19471 12613 19527 12669
rect 19551 12613 19607 12669
rect 19631 12613 19687 12669
rect 19711 12613 19767 12669
rect 19791 12613 19847 12669
rect 19471 12532 19527 12588
rect 19551 12532 19607 12588
rect 19631 12532 19687 12588
rect 19711 12532 19767 12588
rect 19791 12532 19847 12588
rect 19471 12451 19527 12507
rect 19551 12451 19607 12507
rect 19631 12451 19687 12507
rect 19711 12451 19767 12507
rect 19791 12451 19847 12507
rect 19471 12370 19527 12426
rect 19551 12370 19607 12426
rect 19631 12370 19687 12426
rect 19711 12370 19767 12426
rect 19791 12370 19847 12426
rect 19471 12289 19527 12345
rect 19551 12289 19607 12345
rect 19631 12289 19687 12345
rect 19711 12289 19767 12345
rect 19791 12289 19847 12345
rect 19471 12208 19527 12264
rect 19551 12208 19607 12264
rect 19631 12208 19687 12264
rect 19711 12208 19767 12264
rect 19791 12208 19847 12264
rect 19471 12127 19527 12183
rect 19551 12127 19607 12183
rect 19631 12127 19687 12183
rect 19711 12127 19767 12183
rect 19791 12127 19847 12183
rect 19471 12046 19527 12102
rect 19551 12046 19607 12102
rect 19631 12046 19687 12102
rect 19711 12046 19767 12102
rect 19791 12046 19847 12102
rect 19471 11965 19527 12021
rect 19551 11965 19607 12021
rect 19631 11965 19687 12021
rect 19711 11965 19767 12021
rect 19791 11965 19847 12021
rect 19471 11883 19527 11939
rect 19551 11883 19607 11939
rect 19631 11883 19687 11939
rect 19711 11883 19767 11939
rect 19791 11883 19847 11939
rect 19471 11801 19527 11857
rect 19551 11801 19607 11857
rect 19631 11801 19687 11857
rect 19711 11801 19767 11857
rect 19791 11801 19847 11857
rect 19471 11719 19527 11775
rect 19551 11719 19607 11775
rect 19631 11719 19687 11775
rect 19711 11719 19767 11775
rect 19791 11719 19847 11775
rect 19471 11637 19527 11693
rect 19551 11637 19607 11693
rect 19631 11637 19687 11693
rect 19711 11637 19767 11693
rect 19791 11637 19847 11693
rect 19471 11555 19527 11611
rect 19551 11555 19607 11611
rect 19631 11555 19687 11611
rect 19711 11555 19767 11611
rect 19791 11555 19847 11611
rect 19471 11473 19527 11529
rect 19551 11473 19607 11529
rect 19631 11473 19687 11529
rect 19711 11473 19767 11529
rect 19791 11473 19847 11529
rect 19471 11391 19527 11447
rect 19551 11391 19607 11447
rect 19631 11391 19687 11447
rect 19711 11391 19767 11447
rect 19791 11391 19847 11447
rect 19462 11280 19518 11336
rect 19462 11200 19518 11256
rect 19462 11120 19518 11176
rect 19462 11040 19518 11096
rect 19462 10959 19518 11015
rect 19462 10878 19518 10934
rect 19462 10797 19518 10853
rect 19462 10716 19518 10772
rect 19462 10635 19518 10691
rect 19462 10554 19518 10610
rect 19462 10473 19518 10529
rect 19462 10392 19518 10448
rect 19462 10311 19518 10367
rect 19462 10230 19518 10286
rect 19462 10149 19518 10205
rect 19462 10068 19518 10124
rect 19462 9987 19518 10043
rect 19462 9906 19518 9962
rect 19462 9825 19518 9881
rect 19462 9744 19518 9800
rect 19462 9663 19518 9719
rect 19462 9582 19518 9638
rect 19462 9501 19518 9557
rect 19462 9420 19518 9476
rect 19462 9339 19518 9395
rect 19462 9258 19518 9314
rect 19462 9177 19518 9233
rect 19462 9096 19518 9152
rect 19462 9015 19518 9071
rect 19462 8934 19518 8990
rect 19462 8853 19518 8909
rect 19462 8772 19518 8828
rect 19720 11277 19776 11333
rect 19800 11277 19856 11333
rect 19720 11196 19776 11252
rect 19800 11196 19856 11252
rect 19720 11115 19776 11171
rect 19800 11115 19856 11171
rect 19720 11034 19776 11090
rect 19800 11034 19856 11090
rect 19720 10953 19776 11009
rect 19800 10953 19856 11009
rect 19720 10872 19776 10928
rect 19800 10872 19856 10928
rect 19720 10791 19776 10847
rect 19800 10791 19856 10847
rect 19720 10710 19776 10766
rect 19800 10710 19856 10766
rect 19720 10629 19776 10685
rect 19800 10629 19856 10685
rect 19720 10548 19776 10604
rect 19800 10548 19856 10604
rect 19720 10467 19776 10523
rect 19800 10467 19856 10523
rect 19720 10386 19776 10442
rect 19800 10386 19856 10442
rect 19720 10305 19776 10361
rect 19800 10305 19856 10361
rect 19720 10224 19776 10280
rect 19800 10224 19856 10280
rect 19720 10143 19776 10199
rect 19800 10143 19856 10199
rect 19720 10062 19776 10118
rect 19800 10062 19856 10118
rect 19720 9981 19776 10037
rect 19800 9981 19856 10037
rect 19720 9900 19776 9956
rect 19800 9900 19856 9956
rect 19720 9819 19776 9875
rect 19800 9819 19856 9875
rect 19720 9738 19776 9794
rect 19800 9738 19856 9794
rect 19720 9657 19776 9713
rect 19800 9657 19856 9713
rect 19720 9575 19776 9631
rect 19800 9575 19856 9631
rect 19720 9493 19776 9549
rect 19800 9493 19856 9549
rect 19720 9411 19776 9467
rect 19800 9411 19856 9467
rect 19720 9329 19776 9385
rect 19800 9329 19856 9385
rect 19720 9247 19776 9303
rect 19800 9247 19856 9303
rect 19720 9165 19776 9221
rect 19800 9165 19856 9221
rect 19720 9083 19776 9139
rect 19800 9083 19856 9139
rect 19720 9001 19776 9057
rect 19800 9001 19856 9057
rect 19720 8919 19776 8975
rect 19800 8919 19856 8975
rect 19720 8837 19776 8893
rect 19800 8837 19856 8893
rect 19720 8755 19776 8811
rect 19800 8755 19856 8811
rect 19482 8613 19538 8669
rect 19562 8613 19618 8669
rect 19642 8613 19698 8669
rect 19722 8613 19778 8669
rect 19802 8613 19858 8669
rect 19482 8528 19538 8584
rect 19562 8528 19618 8584
rect 19642 8528 19698 8584
rect 19722 8528 19778 8584
rect 19802 8528 19858 8584
rect 19482 8442 19538 8498
rect 19562 8442 19618 8498
rect 19642 8442 19698 8498
rect 19722 8442 19778 8498
rect 19802 8442 19858 8498
rect 19482 8356 19538 8412
rect 19562 8356 19618 8412
rect 19642 8356 19698 8412
rect 19722 8356 19778 8412
rect 19802 8356 19858 8412
rect 19482 8270 19538 8326
rect 19562 8270 19618 8326
rect 19642 8270 19698 8326
rect 19722 8270 19778 8326
rect 19802 8270 19858 8326
rect 19482 8184 19538 8240
rect 19562 8184 19618 8240
rect 19642 8184 19698 8240
rect 19722 8184 19778 8240
rect 19802 8184 19858 8240
rect 19482 8098 19538 8154
rect 19562 8098 19618 8154
rect 19642 8098 19698 8154
rect 19722 8098 19778 8154
rect 19802 8098 19858 8154
rect 19482 8031 19487 8068
rect 19487 8031 19503 8068
rect 19503 8031 19538 8068
rect 19562 8031 19571 8068
rect 19571 8031 19618 8068
rect 19642 8031 19691 8068
rect 19691 8031 19698 8068
rect 19722 8031 19759 8068
rect 19759 8031 19775 8068
rect 19775 8031 19778 8068
rect 19802 8031 19827 8068
rect 19827 8031 19842 8068
rect 19842 8031 19858 8068
rect 19482 8019 19538 8031
rect 19562 8019 19618 8031
rect 19642 8019 19698 8031
rect 19722 8019 19778 8031
rect 19802 8019 19858 8031
rect 19482 8012 19487 8019
rect 19487 8012 19503 8019
rect 19503 8012 19538 8019
rect 19562 8012 19571 8019
rect 19571 8012 19618 8019
rect 19482 7967 19487 7982
rect 19487 7967 19503 7982
rect 19503 7967 19538 7982
rect 19562 7967 19571 7982
rect 19571 7967 19618 7982
rect 19642 8012 19691 8019
rect 19691 8012 19698 8019
rect 19722 8012 19759 8019
rect 19759 8012 19775 8019
rect 19775 8012 19778 8019
rect 19802 8012 19827 8019
rect 19827 8012 19842 8019
rect 19842 8012 19858 8019
rect 19642 7967 19691 7982
rect 19691 7967 19698 7982
rect 19722 7967 19759 7982
rect 19759 7967 19775 7982
rect 19775 7967 19778 7982
rect 19802 7967 19827 7982
rect 19827 7967 19842 7982
rect 19842 7967 19858 7982
rect 19482 7955 19538 7967
rect 19562 7955 19618 7967
rect 19642 7955 19698 7967
rect 19722 7955 19778 7967
rect 19802 7955 19858 7967
rect 19482 7926 19487 7955
rect 19487 7926 19503 7955
rect 19503 7926 19538 7955
rect 19562 7926 19571 7955
rect 19571 7926 19618 7955
rect 19642 7926 19691 7955
rect 19691 7926 19698 7955
rect 19722 7926 19759 7955
rect 19759 7926 19775 7955
rect 19775 7926 19778 7955
rect 19802 7926 19827 7955
rect 19827 7926 19842 7955
rect 19842 7926 19858 7955
rect -1954 5094 -1418 5550
rect -1954 5013 -1898 5069
rect -1874 5013 -1818 5069
rect -1794 5013 -1738 5069
rect -1714 5013 -1658 5069
rect -1634 5013 -1578 5069
rect -1554 5013 -1498 5069
rect -1474 5013 -1418 5069
rect -1954 4932 -1898 4988
rect -1874 4932 -1818 4988
rect -1794 4932 -1738 4988
rect -1714 4932 -1658 4988
rect -1634 4932 -1578 4988
rect -1554 4932 -1498 4988
rect -1474 4932 -1418 4988
rect -1954 4851 -1898 4907
rect -1874 4851 -1818 4907
rect -1794 4851 -1738 4907
rect -1714 4851 -1658 4907
rect -1634 4851 -1578 4907
rect -1554 4851 -1498 4907
rect -1474 4851 -1418 4907
rect -1954 4770 -1898 4826
rect -1874 4770 -1818 4826
rect -1794 4770 -1738 4826
rect -1714 4770 -1658 4826
rect -1634 4770 -1578 4826
rect -1554 4770 -1498 4826
rect -1474 4770 -1418 4826
rect -1954 4689 -1898 4745
rect -1874 4689 -1818 4745
rect -1794 4689 -1738 4745
rect -1714 4689 -1658 4745
rect -1634 4689 -1578 4745
rect -1554 4689 -1498 4745
rect -1474 4689 -1418 4745
rect -1954 4608 -1898 4664
rect -1874 4608 -1818 4664
rect -1794 4608 -1738 4664
rect -1714 4608 -1658 4664
rect -1634 4608 -1578 4664
rect -1554 4608 -1498 4664
rect -1474 4608 -1418 4664
rect -1954 4527 -1898 4583
rect -1874 4527 -1818 4583
rect -1794 4527 -1738 4583
rect -1714 4527 -1658 4583
rect -1634 4527 -1578 4583
rect -1554 4527 -1498 4583
rect -1474 4527 -1418 4583
rect -1954 4446 -1898 4502
rect -1874 4446 -1818 4502
rect -1794 4446 -1738 4502
rect -1714 4446 -1658 4502
rect -1634 4446 -1578 4502
rect -1554 4446 -1498 4502
rect -1474 4446 -1418 4502
rect -163 5094 373 5550
rect -163 5013 -107 5069
rect -83 5013 -27 5069
rect -3 5013 53 5069
rect 77 5013 133 5069
rect 157 5013 213 5069
rect 237 5013 293 5069
rect 317 5013 373 5069
rect -163 4932 -107 4988
rect -83 4932 -27 4988
rect -3 4932 53 4988
rect 77 4932 133 4988
rect 157 4932 213 4988
rect 237 4932 293 4988
rect 317 4932 373 4988
rect -163 4851 -107 4907
rect -83 4851 -27 4907
rect -3 4851 53 4907
rect 77 4851 133 4907
rect 157 4851 213 4907
rect 237 4851 293 4907
rect 317 4851 373 4907
rect -163 4770 -107 4826
rect -83 4770 -27 4826
rect -3 4770 53 4826
rect 77 4770 133 4826
rect 157 4770 213 4826
rect 237 4770 293 4826
rect 317 4770 373 4826
rect -163 4689 -107 4745
rect -83 4689 -27 4745
rect -3 4689 53 4745
rect 77 4689 133 4745
rect 157 4689 213 4745
rect 237 4689 293 4745
rect 317 4689 373 4745
rect -163 4608 -107 4664
rect -83 4608 -27 4664
rect -3 4608 53 4664
rect 77 4608 133 4664
rect 157 4608 213 4664
rect 237 4608 293 4664
rect 317 4608 373 4664
rect -163 4527 -107 4583
rect -83 4527 -27 4583
rect -3 4527 53 4583
rect 77 4527 133 4583
rect 157 4527 213 4583
rect 237 4527 293 4583
rect 317 4527 373 4583
rect -163 4446 -107 4502
rect -83 4446 -27 4502
rect -3 4446 53 4502
rect 77 4446 133 4502
rect 157 4446 213 4502
rect 237 4446 293 4502
rect 317 4446 373 4502
rect 1657 5094 2193 5550
rect 1657 5013 1713 5069
rect 1737 5013 1793 5069
rect 1817 5013 1873 5069
rect 1897 5013 1953 5069
rect 1977 5013 2033 5069
rect 2057 5013 2113 5069
rect 2137 5013 2193 5069
rect 1657 4932 1713 4988
rect 1737 4932 1793 4988
rect 1817 4932 1873 4988
rect 1897 4932 1953 4988
rect 1977 4932 2033 4988
rect 2057 4932 2113 4988
rect 2137 4932 2193 4988
rect 1657 4851 1713 4907
rect 1737 4851 1793 4907
rect 1817 4851 1873 4907
rect 1897 4851 1953 4907
rect 1977 4851 2033 4907
rect 2057 4851 2113 4907
rect 2137 4851 2193 4907
rect 1657 4770 1713 4826
rect 1737 4770 1793 4826
rect 1817 4770 1873 4826
rect 1897 4770 1953 4826
rect 1977 4770 2033 4826
rect 2057 4770 2113 4826
rect 2137 4770 2193 4826
rect 1657 4689 1713 4745
rect 1737 4689 1793 4745
rect 1817 4689 1873 4745
rect 1897 4689 1953 4745
rect 1977 4689 2033 4745
rect 2057 4689 2113 4745
rect 2137 4689 2193 4745
rect 1657 4608 1713 4664
rect 1737 4608 1793 4664
rect 1817 4608 1873 4664
rect 1897 4608 1953 4664
rect 1977 4608 2033 4664
rect 2057 4608 2113 4664
rect 2137 4608 2193 4664
rect 1657 4527 1713 4583
rect 1737 4527 1793 4583
rect 1817 4527 1873 4583
rect 1897 4527 1953 4583
rect 1977 4527 2033 4583
rect 2057 4527 2113 4583
rect 2137 4527 2193 4583
rect 3458 5094 3994 5550
rect 3458 5013 3514 5069
rect 3538 5013 3594 5069
rect 3618 5013 3674 5069
rect 3698 5013 3754 5069
rect 3778 5013 3834 5069
rect 3858 5013 3914 5069
rect 3938 5013 3994 5069
rect 3458 4932 3514 4988
rect 3538 4932 3594 4988
rect 3618 4932 3674 4988
rect 3698 4932 3754 4988
rect 3778 4932 3834 4988
rect 3858 4932 3914 4988
rect 3938 4932 3994 4988
rect 3458 4851 3514 4907
rect 3538 4851 3594 4907
rect 3618 4851 3674 4907
rect 3698 4851 3754 4907
rect 3778 4851 3834 4907
rect 3858 4851 3914 4907
rect 3938 4851 3994 4907
rect 3458 4770 3514 4826
rect 3538 4770 3594 4826
rect 3618 4770 3674 4826
rect 3698 4770 3754 4826
rect 3778 4770 3834 4826
rect 3858 4770 3914 4826
rect 3938 4770 3994 4826
rect 3458 4689 3514 4745
rect 3538 4689 3594 4745
rect 3618 4689 3674 4745
rect 3698 4689 3754 4745
rect 3778 4689 3834 4745
rect 3858 4689 3914 4745
rect 3938 4689 3994 4745
rect 3458 4608 3514 4664
rect 3538 4608 3594 4664
rect 3618 4608 3674 4664
rect 3698 4608 3754 4664
rect 3778 4608 3834 4664
rect 3858 4608 3914 4664
rect 3938 4608 3994 4664
rect 1657 4446 1713 4502
rect 1737 4446 1793 4502
rect 1817 4446 1873 4502
rect 1897 4446 1953 4502
rect 1977 4446 2033 4502
rect 2057 4446 2113 4502
rect 2137 4446 2193 4502
rect 3458 4527 3514 4583
rect 3538 4527 3594 4583
rect 3618 4527 3674 4583
rect 3698 4527 3754 4583
rect 3778 4527 3834 4583
rect 3858 4527 3914 4583
rect 3938 4527 3994 4583
rect 5266 5094 5802 5550
rect 5266 5013 5322 5069
rect 5346 5013 5402 5069
rect 5426 5013 5482 5069
rect 5506 5013 5562 5069
rect 5586 5013 5642 5069
rect 5666 5013 5722 5069
rect 5746 5013 5802 5069
rect 5266 4932 5322 4988
rect 5346 4932 5402 4988
rect 5426 4932 5482 4988
rect 5506 4932 5562 4988
rect 5586 4932 5642 4988
rect 5666 4932 5722 4988
rect 5746 4932 5802 4988
rect 5266 4851 5322 4907
rect 5346 4851 5402 4907
rect 5426 4851 5482 4907
rect 5506 4851 5562 4907
rect 5586 4851 5642 4907
rect 5666 4851 5722 4907
rect 5746 4851 5802 4907
rect 5266 4770 5322 4826
rect 5346 4770 5402 4826
rect 5426 4770 5482 4826
rect 5506 4770 5562 4826
rect 5586 4770 5642 4826
rect 5666 4770 5722 4826
rect 5746 4770 5802 4826
rect 5266 4689 5322 4745
rect 5346 4689 5402 4745
rect 5426 4689 5482 4745
rect 5506 4689 5562 4745
rect 5586 4689 5642 4745
rect 5666 4689 5722 4745
rect 5746 4689 5802 4745
rect 7061 5494 7117 5550
rect 7141 5494 7197 5550
rect 7221 5494 7277 5550
rect 7301 5494 7357 5550
rect 7381 5494 7437 5550
rect 7461 5494 7517 5550
rect 7541 5494 7597 5550
rect 7061 5411 7117 5467
rect 7141 5411 7197 5467
rect 7221 5411 7277 5467
rect 7301 5411 7357 5467
rect 7381 5411 7437 5467
rect 7461 5411 7517 5467
rect 7541 5411 7597 5467
rect 7061 5328 7117 5384
rect 7141 5328 7197 5384
rect 7221 5328 7277 5384
rect 7301 5328 7357 5384
rect 7381 5328 7437 5384
rect 7461 5328 7517 5384
rect 7541 5328 7597 5384
rect 7061 5245 7117 5301
rect 7141 5245 7197 5301
rect 7221 5245 7277 5301
rect 7301 5245 7357 5301
rect 7381 5245 7437 5301
rect 7461 5245 7517 5301
rect 7541 5245 7597 5301
rect 7061 5162 7117 5218
rect 7141 5162 7197 5218
rect 7221 5162 7277 5218
rect 7301 5162 7357 5218
rect 7381 5162 7437 5218
rect 7461 5162 7517 5218
rect 7541 5162 7597 5218
rect 7061 5078 7117 5134
rect 7141 5078 7197 5134
rect 7221 5078 7277 5134
rect 7301 5078 7357 5134
rect 7381 5078 7437 5134
rect 7461 5078 7517 5134
rect 7541 5078 7597 5134
rect 7061 4994 7117 5050
rect 7141 4994 7197 5050
rect 7221 4994 7277 5050
rect 7301 4994 7357 5050
rect 7381 4994 7437 5050
rect 7461 4994 7517 5050
rect 7541 4994 7597 5050
rect 7061 4910 7117 4966
rect 7141 4910 7197 4966
rect 7221 4910 7277 4966
rect 7301 4910 7357 4966
rect 7381 4910 7437 4966
rect 7461 4910 7517 4966
rect 7541 4910 7597 4966
rect 7061 4826 7117 4882
rect 7141 4826 7197 4882
rect 7221 4826 7277 4882
rect 7301 4826 7357 4882
rect 7381 4826 7437 4882
rect 7461 4826 7517 4882
rect 7541 4826 7597 4882
rect 7061 4742 7117 4798
rect 7141 4742 7197 4798
rect 7221 4742 7277 4798
rect 7301 4742 7357 4798
rect 7381 4742 7437 4798
rect 7461 4742 7517 4798
rect 7541 4742 7597 4798
rect 8872 5474 8928 5530
rect 8952 5474 9008 5530
rect 9032 5474 9088 5530
rect 9112 5474 9168 5530
rect 9192 5474 9248 5530
rect 9272 5474 9328 5530
rect 9352 5474 9408 5530
rect 8872 5393 8928 5449
rect 8952 5393 9008 5449
rect 9032 5393 9088 5449
rect 9112 5393 9168 5449
rect 9192 5393 9248 5449
rect 9272 5393 9328 5449
rect 9352 5393 9408 5449
rect 8872 5312 8928 5368
rect 8952 5312 9008 5368
rect 9032 5312 9088 5368
rect 9112 5312 9168 5368
rect 9192 5312 9248 5368
rect 9272 5312 9328 5368
rect 9352 5312 9408 5368
rect 8872 5231 8928 5287
rect 8952 5231 9008 5287
rect 9032 5231 9088 5287
rect 9112 5231 9168 5287
rect 9192 5231 9248 5287
rect 9272 5231 9328 5287
rect 9352 5231 9408 5287
rect 8872 5150 8928 5206
rect 8952 5150 9008 5206
rect 9032 5150 9088 5206
rect 9112 5150 9168 5206
rect 9192 5150 9248 5206
rect 9272 5150 9328 5206
rect 9352 5150 9408 5206
rect 8872 5069 8928 5125
rect 8952 5069 9008 5125
rect 9032 5069 9088 5125
rect 9112 5069 9168 5125
rect 9192 5069 9248 5125
rect 9272 5069 9328 5125
rect 9352 5069 9408 5125
rect 8872 4988 8928 5044
rect 8952 4988 9008 5044
rect 9032 4988 9088 5044
rect 9112 4988 9168 5044
rect 9192 4988 9248 5044
rect 9272 4988 9328 5044
rect 9352 4988 9408 5044
rect 8872 4907 8928 4963
rect 8952 4907 9008 4963
rect 9032 4907 9088 4963
rect 9112 4907 9168 4963
rect 9192 4907 9248 4963
rect 9272 4907 9328 4963
rect 9352 4907 9408 4963
rect 8872 4825 8928 4881
rect 8952 4825 9008 4881
rect 9032 4825 9088 4881
rect 9112 4825 9168 4881
rect 9192 4825 9248 4881
rect 9272 4825 9328 4881
rect 9352 4825 9408 4881
rect 8872 4743 8928 4799
rect 8952 4743 9008 4799
rect 9032 4743 9088 4799
rect 9112 4743 9168 4799
rect 9192 4743 9248 4799
rect 9272 4743 9328 4799
rect 9352 4743 9408 4799
rect 5266 4608 5322 4664
rect 5346 4608 5402 4664
rect 5426 4608 5482 4664
rect 5506 4608 5562 4664
rect 5586 4608 5642 4664
rect 5666 4608 5722 4664
rect 5746 4608 5802 4664
rect 8872 4661 8928 4717
rect 8952 4661 9008 4717
rect 9032 4661 9088 4717
rect 9112 4661 9168 4717
rect 9192 4661 9248 4717
rect 9272 4661 9328 4717
rect 9352 4661 9408 4717
rect 3458 4446 3514 4502
rect 3538 4446 3594 4502
rect 3618 4446 3674 4502
rect 3698 4446 3754 4502
rect 3778 4446 3834 4502
rect 3858 4446 3914 4502
rect 3938 4446 3994 4502
rect 865 4228 921 4284
rect 945 4228 1001 4284
rect 1025 4228 1081 4284
rect 865 4144 921 4200
rect 945 4144 1001 4200
rect 1025 4144 1081 4200
rect 865 4060 921 4116
rect 945 4060 1001 4116
rect 1025 4060 1081 4116
rect 865 3975 921 4031
rect 945 3975 1001 4031
rect 1025 3975 1081 4031
rect 865 3890 921 3946
rect 945 3890 1001 3946
rect 1025 3890 1081 3946
rect 865 3805 921 3861
rect 945 3805 1001 3861
rect 1025 3805 1081 3861
rect 865 3720 921 3776
rect 945 3720 1001 3776
rect 1025 3720 1081 3776
rect 167 1447 623 3183
rect 167 1366 223 1422
rect 247 1366 303 1422
rect 327 1366 383 1422
rect 407 1366 463 1422
rect 487 1366 543 1422
rect 567 1366 623 1422
rect 2288 3127 2344 3183
rect 2368 3127 2424 3183
rect 2448 3127 2504 3183
rect 2528 3127 2584 3183
rect 2608 3127 2664 3183
rect 2688 3127 2744 3183
rect 2288 3037 2344 3093
rect 2368 3037 2424 3093
rect 2448 3037 2504 3093
rect 2528 3037 2584 3093
rect 2608 3037 2664 3093
rect 2688 3037 2744 3093
rect 2288 2947 2344 3003
rect 2368 2947 2424 3003
rect 2448 2947 2504 3003
rect 2528 2947 2584 3003
rect 2608 2947 2664 3003
rect 2688 2947 2744 3003
rect 2288 2857 2344 2913
rect 2368 2857 2424 2913
rect 2448 2857 2504 2913
rect 2528 2857 2584 2913
rect 2608 2857 2664 2913
rect 2688 2857 2744 2913
rect 2288 2767 2344 2823
rect 2368 2767 2424 2823
rect 2448 2767 2504 2823
rect 2528 2767 2584 2823
rect 2608 2767 2664 2823
rect 2688 2767 2744 2823
rect 2288 2677 2344 2733
rect 2368 2677 2424 2733
rect 2448 2677 2504 2733
rect 2528 2677 2584 2733
rect 2608 2677 2664 2733
rect 2688 2677 2744 2733
rect 2288 2586 2344 2642
rect 2368 2586 2424 2642
rect 2448 2586 2504 2642
rect 2528 2586 2584 2642
rect 2608 2586 2664 2642
rect 2688 2586 2744 2642
rect 2288 2495 2344 2551
rect 2368 2495 2424 2551
rect 2448 2495 2504 2551
rect 2528 2495 2584 2551
rect 2608 2495 2664 2551
rect 2688 2495 2744 2551
rect 5266 4527 5322 4583
rect 5346 4527 5402 4583
rect 5426 4527 5482 4583
rect 5506 4527 5562 4583
rect 5586 4527 5642 4583
rect 5666 4527 5722 4583
rect 5746 4527 5802 4583
rect 5266 4446 5322 4502
rect 5346 4446 5402 4502
rect 5426 4446 5482 4502
rect 5506 4446 5562 4502
rect 5586 4446 5642 4502
rect 5666 4446 5722 4502
rect 5746 4446 5802 4502
rect 8872 4579 8928 4635
rect 8952 4579 9008 4635
rect 9032 4579 9088 4635
rect 9112 4579 9168 4635
rect 9192 4579 9248 4635
rect 9272 4579 9328 4635
rect 9352 4579 9408 4635
rect 8872 4497 8928 4553
rect 8952 4497 9008 4553
rect 9032 4497 9088 4553
rect 9112 4497 9168 4553
rect 9192 4497 9248 4553
rect 9272 4497 9328 4553
rect 9352 4497 9408 4553
rect 10660 5502 10716 5558
rect 10740 5502 10796 5558
rect 10820 5502 10876 5558
rect 10900 5502 10956 5558
rect 10980 5502 11036 5558
rect 11060 5502 11116 5558
rect 11140 5502 11196 5558
rect 10660 5420 10716 5476
rect 10740 5420 10796 5476
rect 10820 5420 10876 5476
rect 10900 5420 10956 5476
rect 10980 5420 11036 5476
rect 11060 5420 11116 5476
rect 11140 5420 11196 5476
rect 12465 5502 12521 5558
rect 12545 5502 12601 5558
rect 12625 5502 12681 5558
rect 12705 5502 12761 5558
rect 12785 5502 12841 5558
rect 12865 5502 12921 5558
rect 12945 5502 13001 5558
rect 12465 5420 12521 5476
rect 12545 5420 12601 5476
rect 12625 5420 12681 5476
rect 12705 5420 12761 5476
rect 12785 5420 12841 5476
rect 12865 5420 12921 5476
rect 12945 5420 13001 5476
rect 14278 5502 14334 5558
rect 14358 5502 14414 5558
rect 14438 5502 14494 5558
rect 14518 5502 14574 5558
rect 14598 5502 14654 5558
rect 14678 5502 14734 5558
rect 14758 5502 14814 5558
rect 10660 5337 10716 5393
rect 10740 5337 10796 5393
rect 10820 5337 10876 5393
rect 10900 5337 10956 5393
rect 10980 5337 11036 5393
rect 11060 5337 11116 5393
rect 11140 5337 11196 5393
rect 10660 5254 10716 5310
rect 10740 5254 10796 5310
rect 10820 5254 10876 5310
rect 10900 5254 10956 5310
rect 10980 5254 11036 5310
rect 11060 5254 11116 5310
rect 11140 5254 11196 5310
rect 10660 5171 10716 5227
rect 10740 5171 10796 5227
rect 10820 5171 10876 5227
rect 10900 5171 10956 5227
rect 10980 5171 11036 5227
rect 11060 5171 11116 5227
rect 11140 5171 11196 5227
rect 14278 5420 14334 5476
rect 14358 5420 14414 5476
rect 14438 5420 14494 5476
rect 14518 5420 14574 5476
rect 14598 5420 14654 5476
rect 14678 5420 14734 5476
rect 14758 5420 14814 5476
rect 12465 5337 12521 5393
rect 12545 5337 12601 5393
rect 12625 5337 12681 5393
rect 12705 5337 12761 5393
rect 12785 5337 12841 5393
rect 12865 5337 12921 5393
rect 12945 5337 13001 5393
rect 12465 5254 12521 5310
rect 12545 5254 12601 5310
rect 12625 5254 12681 5310
rect 12705 5254 12761 5310
rect 12785 5254 12841 5310
rect 12865 5254 12921 5310
rect 12945 5254 13001 5310
rect 12465 5171 12521 5227
rect 12545 5171 12601 5227
rect 12625 5171 12681 5227
rect 12705 5171 12761 5227
rect 12785 5171 12841 5227
rect 12865 5171 12921 5227
rect 12945 5171 13001 5227
rect 14278 5337 14334 5393
rect 14358 5337 14414 5393
rect 14438 5337 14494 5393
rect 14518 5337 14574 5393
rect 14598 5337 14654 5393
rect 14678 5337 14734 5393
rect 14758 5337 14814 5393
rect 14278 5254 14334 5310
rect 14358 5254 14414 5310
rect 14438 5254 14494 5310
rect 14518 5254 14574 5310
rect 14598 5254 14654 5310
rect 14678 5254 14734 5310
rect 14758 5254 14814 5310
rect 10660 5088 10716 5144
rect 10740 5088 10796 5144
rect 10820 5088 10876 5144
rect 10900 5088 10956 5144
rect 10980 5088 11036 5144
rect 11060 5088 11116 5144
rect 11140 5088 11196 5144
rect 10660 5005 10716 5061
rect 10740 5005 10796 5061
rect 10820 5005 10876 5061
rect 10900 5005 10956 5061
rect 10980 5005 11036 5061
rect 11060 5005 11116 5061
rect 11140 5005 11196 5061
rect 10660 4922 10716 4978
rect 10740 4922 10796 4978
rect 10820 4922 10876 4978
rect 10900 4922 10956 4978
rect 10980 4922 11036 4978
rect 11060 4922 11116 4978
rect 11140 4922 11196 4978
rect 10660 4839 10716 4895
rect 10740 4839 10796 4895
rect 10820 4839 10876 4895
rect 10900 4839 10956 4895
rect 10980 4839 11036 4895
rect 11060 4839 11116 4895
rect 11140 4839 11196 4895
rect 10660 4756 10716 4812
rect 10740 4756 10796 4812
rect 10820 4756 10876 4812
rect 10900 4756 10956 4812
rect 10980 4756 11036 4812
rect 11060 4756 11116 4812
rect 11140 4756 11196 4812
rect 10660 4673 10716 4729
rect 10740 4673 10796 4729
rect 10820 4673 10876 4729
rect 10900 4673 10956 4729
rect 10980 4673 11036 4729
rect 11060 4673 11116 4729
rect 11140 4673 11196 4729
rect 10660 4590 10716 4646
rect 10740 4590 10796 4646
rect 10820 4590 10876 4646
rect 10900 4590 10956 4646
rect 10980 4590 11036 4646
rect 11060 4590 11116 4646
rect 11140 4590 11196 4646
rect 10660 4507 10716 4563
rect 10740 4507 10796 4563
rect 10820 4507 10876 4563
rect 10900 4507 10956 4563
rect 10980 4507 11036 4563
rect 11060 4507 11116 4563
rect 11140 4507 11196 4563
rect 14278 5171 14334 5227
rect 14358 5171 14414 5227
rect 14438 5171 14494 5227
rect 14518 5171 14574 5227
rect 14598 5171 14654 5227
rect 14678 5171 14734 5227
rect 14758 5171 14814 5227
rect 12465 5088 12521 5144
rect 12545 5088 12601 5144
rect 12625 5088 12681 5144
rect 12705 5088 12761 5144
rect 12785 5088 12841 5144
rect 12865 5088 12921 5144
rect 12945 5088 13001 5144
rect 12465 5005 12521 5061
rect 12545 5005 12601 5061
rect 12625 5005 12681 5061
rect 12705 5005 12761 5061
rect 12785 5005 12841 5061
rect 12865 5005 12921 5061
rect 12945 5005 13001 5061
rect 12465 4922 12521 4978
rect 12545 4922 12601 4978
rect 12625 4922 12681 4978
rect 12705 4922 12761 4978
rect 12785 4922 12841 4978
rect 12865 4922 12921 4978
rect 12945 4922 13001 4978
rect 12465 4839 12521 4895
rect 12545 4839 12601 4895
rect 12625 4839 12681 4895
rect 12705 4839 12761 4895
rect 12785 4839 12841 4895
rect 12865 4839 12921 4895
rect 12945 4839 13001 4895
rect 12465 4756 12521 4812
rect 12545 4756 12601 4812
rect 12625 4756 12681 4812
rect 12705 4756 12761 4812
rect 12785 4756 12841 4812
rect 12865 4756 12921 4812
rect 12945 4756 13001 4812
rect 12465 4673 12521 4729
rect 12545 4673 12601 4729
rect 12625 4673 12681 4729
rect 12705 4673 12761 4729
rect 12785 4673 12841 4729
rect 12865 4673 12921 4729
rect 12945 4673 13001 4729
rect 12465 4590 12521 4646
rect 12545 4590 12601 4646
rect 12625 4590 12681 4646
rect 12705 4590 12761 4646
rect 12785 4590 12841 4646
rect 12865 4590 12921 4646
rect 12945 4590 13001 4646
rect 12465 4507 12521 4563
rect 12545 4507 12601 4563
rect 12625 4507 12681 4563
rect 12705 4507 12761 4563
rect 12785 4507 12841 4563
rect 12865 4507 12921 4563
rect 12945 4507 13001 4563
rect 14278 5088 14334 5144
rect 14358 5088 14414 5144
rect 14438 5088 14494 5144
rect 14518 5088 14574 5144
rect 14598 5088 14654 5144
rect 14678 5088 14734 5144
rect 14758 5088 14814 5144
rect 14278 5005 14334 5061
rect 14358 5005 14414 5061
rect 14438 5005 14494 5061
rect 14518 5005 14574 5061
rect 14598 5005 14654 5061
rect 14678 5005 14734 5061
rect 14758 5005 14814 5061
rect 14278 4922 14334 4978
rect 14358 4922 14414 4978
rect 14438 4922 14494 4978
rect 14518 4922 14574 4978
rect 14598 4922 14654 4978
rect 14678 4922 14734 4978
rect 14758 4922 14814 4978
rect 14278 4839 14334 4895
rect 14358 4839 14414 4895
rect 14438 4839 14494 4895
rect 14518 4839 14574 4895
rect 14598 4839 14654 4895
rect 14678 4839 14734 4895
rect 14758 4839 14814 4895
rect 14278 4756 14334 4812
rect 14358 4756 14414 4812
rect 14438 4756 14494 4812
rect 14518 4756 14574 4812
rect 14598 4756 14654 4812
rect 14678 4756 14734 4812
rect 14758 4756 14814 4812
rect 14278 4673 14334 4729
rect 14358 4673 14414 4729
rect 14438 4673 14494 4729
rect 14518 4673 14574 4729
rect 14598 4673 14654 4729
rect 14678 4673 14734 4729
rect 14758 4673 14814 4729
rect 14278 4590 14334 4646
rect 14358 4590 14414 4646
rect 14438 4590 14494 4646
rect 14518 4590 14574 4646
rect 14598 4590 14654 4646
rect 14678 4590 14734 4646
rect 14758 4590 14814 4646
rect 14278 4507 14334 4563
rect 14358 4507 14414 4563
rect 14438 4507 14494 4563
rect 14518 4507 14574 4563
rect 14598 4507 14654 4563
rect 14678 4507 14734 4563
rect 14758 4507 14814 4563
rect 16064 5500 16120 5556
rect 16144 5500 16200 5556
rect 16224 5500 16280 5556
rect 16304 5500 16360 5556
rect 16384 5500 16440 5556
rect 16464 5500 16520 5556
rect 16064 5418 16120 5474
rect 16144 5418 16200 5474
rect 16224 5418 16280 5474
rect 16304 5418 16360 5474
rect 16384 5418 16440 5474
rect 16464 5418 16520 5474
rect 16064 5336 16120 5392
rect 16144 5336 16200 5392
rect 16224 5336 16280 5392
rect 16304 5336 16360 5392
rect 16384 5336 16440 5392
rect 16464 5336 16520 5392
rect 16064 5254 16120 5310
rect 16144 5254 16200 5310
rect 16224 5254 16280 5310
rect 16304 5254 16360 5310
rect 16384 5254 16440 5310
rect 16464 5254 16520 5310
rect 16064 5172 16120 5228
rect 16144 5172 16200 5228
rect 16224 5172 16280 5228
rect 16304 5172 16360 5228
rect 16384 5172 16440 5228
rect 16464 5172 16520 5228
rect 16064 5090 16120 5146
rect 16144 5090 16200 5146
rect 16224 5090 16280 5146
rect 16304 5090 16360 5146
rect 16384 5090 16440 5146
rect 16464 5090 16520 5146
rect 16064 5008 16120 5064
rect 16144 5008 16200 5064
rect 16224 5008 16280 5064
rect 16304 5008 16360 5064
rect 16384 5008 16440 5064
rect 16464 5008 16520 5064
rect 16064 4926 16120 4982
rect 16144 4926 16200 4982
rect 16224 4926 16280 4982
rect 16304 4926 16360 4982
rect 16384 4926 16440 4982
rect 16464 4926 16520 4982
rect 16064 4844 16120 4900
rect 16144 4844 16200 4900
rect 16224 4844 16280 4900
rect 16304 4844 16360 4900
rect 16384 4844 16440 4900
rect 16464 4844 16520 4900
rect 16064 4762 16120 4818
rect 16144 4762 16200 4818
rect 16224 4762 16280 4818
rect 16304 4762 16360 4818
rect 16384 4762 16440 4818
rect 16464 4762 16520 4818
rect 16064 4679 16120 4735
rect 16144 4679 16200 4735
rect 16224 4679 16280 4735
rect 16304 4679 16360 4735
rect 16384 4679 16440 4735
rect 16464 4679 16520 4735
rect 16064 4596 16120 4652
rect 16144 4596 16200 4652
rect 16224 4596 16280 4652
rect 16304 4596 16360 4652
rect 16384 4596 16440 4652
rect 16464 4596 16520 4652
rect 4228 3082 4284 3138
rect 4308 3082 4364 3138
rect 4388 3082 4444 3138
rect 4468 3082 4524 3138
rect 4548 3082 4604 3138
rect 4628 3082 4684 3138
rect 4708 3082 4764 3138
rect 4788 3082 4844 3138
rect 4868 3082 4924 3138
rect 4948 3082 5004 3138
rect 5028 3082 5084 3138
rect 4228 3001 4284 3057
rect 4308 3001 4364 3057
rect 4388 3001 4444 3057
rect 4468 3001 4524 3057
rect 4548 3001 4604 3057
rect 4628 3001 4684 3057
rect 4708 3001 4764 3057
rect 4788 3001 4844 3057
rect 4868 3001 4924 3057
rect 4948 3001 5004 3057
rect 5028 3001 5084 3057
rect 4228 2920 4284 2976
rect 4308 2920 4364 2976
rect 4388 2920 4444 2976
rect 4468 2920 4524 2976
rect 4548 2920 4604 2976
rect 4628 2920 4684 2976
rect 4708 2920 4764 2976
rect 4788 2920 4844 2976
rect 4868 2920 4924 2976
rect 4948 2920 5004 2976
rect 5028 2920 5084 2976
rect 4228 2839 4284 2895
rect 4308 2839 4364 2895
rect 4388 2839 4444 2895
rect 4468 2839 4524 2895
rect 4548 2839 4604 2895
rect 4628 2839 4684 2895
rect 4708 2839 4764 2895
rect 4788 2839 4844 2895
rect 4868 2839 4924 2895
rect 4948 2839 5004 2895
rect 5028 2839 5084 2895
rect 4228 2758 4284 2814
rect 4308 2758 4364 2814
rect 4388 2758 4444 2814
rect 4468 2758 4524 2814
rect 4548 2758 4604 2814
rect 4628 2758 4684 2814
rect 4708 2758 4764 2814
rect 4788 2758 4844 2814
rect 4868 2758 4924 2814
rect 4948 2758 5004 2814
rect 5028 2758 5084 2814
rect 4228 2677 4284 2733
rect 4308 2677 4364 2733
rect 4388 2677 4444 2733
rect 4468 2677 4524 2733
rect 4548 2677 4604 2733
rect 4628 2677 4684 2733
rect 4708 2677 4764 2733
rect 4788 2677 4844 2733
rect 4868 2677 4924 2733
rect 4948 2677 5004 2733
rect 5028 2677 5084 2733
rect 1594 1962 1650 2018
rect 1674 1962 1730 2018
rect 1754 1962 1810 2018
rect 1834 1962 1890 2018
rect 1594 1876 1650 1932
rect 1674 1876 1730 1932
rect 1754 1876 1810 1932
rect 1834 1876 1890 1932
rect 1594 1790 1650 1846
rect 1674 1790 1730 1846
rect 1754 1790 1810 1846
rect 1834 1790 1890 1846
rect 1594 1704 1650 1760
rect 1674 1704 1730 1760
rect 1754 1704 1810 1760
rect 1834 1704 1890 1760
rect 1594 1618 1650 1674
rect 1674 1618 1730 1674
rect 1754 1618 1810 1674
rect 1834 1618 1890 1674
rect 1594 1531 1650 1587
rect 1674 1531 1730 1587
rect 1754 1531 1810 1587
rect 1834 1531 1890 1587
rect 1594 1444 1650 1500
rect 1674 1444 1730 1500
rect 1754 1444 1810 1500
rect 1834 1444 1890 1500
rect 1594 1357 1650 1413
rect 1674 1357 1730 1413
rect 1754 1357 1810 1413
rect 1834 1357 1890 1413
rect 2415 1962 2471 2018
rect 2495 1962 2551 2018
rect 2575 1962 2631 2018
rect 2655 1962 2711 2018
rect 2415 1876 2471 1932
rect 2495 1876 2551 1932
rect 2575 1876 2631 1932
rect 2655 1876 2711 1932
rect 2415 1790 2471 1846
rect 2495 1790 2551 1846
rect 2575 1790 2631 1846
rect 2655 1790 2711 1846
rect 2415 1704 2471 1760
rect 2495 1704 2551 1760
rect 2575 1704 2631 1760
rect 2655 1704 2711 1760
rect 2415 1618 2471 1674
rect 2495 1618 2551 1674
rect 2575 1618 2631 1674
rect 2655 1618 2711 1674
rect 2415 1531 2471 1587
rect 2495 1531 2551 1587
rect 2575 1531 2631 1587
rect 2655 1531 2711 1587
rect 2415 1444 2471 1500
rect 2495 1444 2551 1500
rect 2575 1444 2631 1500
rect 2655 1444 2711 1500
rect 2415 1357 2471 1413
rect 2495 1357 2551 1413
rect 2575 1357 2631 1413
rect 2655 1357 2711 1413
rect 4228 2596 4284 2652
rect 4308 2596 4364 2652
rect 4388 2596 4444 2652
rect 4468 2596 4524 2652
rect 4548 2596 4604 2652
rect 4628 2596 4684 2652
rect 4708 2596 4764 2652
rect 4788 2596 4844 2652
rect 4868 2596 4924 2652
rect 4948 2596 5004 2652
rect 5028 2596 5084 2652
rect 4228 2515 4284 2571
rect 4308 2515 4364 2571
rect 4388 2515 4444 2571
rect 4468 2515 4524 2571
rect 4548 2515 4604 2571
rect 4628 2515 4684 2571
rect 4708 2515 4764 2571
rect 4788 2515 4844 2571
rect 4868 2515 4924 2571
rect 4948 2515 5004 2571
rect 5028 2515 5084 2571
rect 4228 2434 4284 2490
rect 4308 2434 4364 2490
rect 4388 2434 4444 2490
rect 4468 2434 4524 2490
rect 4548 2434 4604 2490
rect 4628 2434 4684 2490
rect 4708 2434 4764 2490
rect 4788 2434 4844 2490
rect 4868 2434 4924 2490
rect 4948 2434 5004 2490
rect 5028 2434 5084 2490
rect 4228 2352 4284 2408
rect 4308 2352 4364 2408
rect 4388 2352 4444 2408
rect 4468 2352 4524 2408
rect 4548 2352 4604 2408
rect 4628 2352 4684 2408
rect 4708 2352 4764 2408
rect 4788 2352 4844 2408
rect 4868 2352 4924 2408
rect 4948 2352 5004 2408
rect 5028 2352 5084 2408
rect 4228 2270 4284 2326
rect 4308 2270 4364 2326
rect 4388 2270 4444 2326
rect 4468 2270 4524 2326
rect 4548 2270 4604 2326
rect 4628 2270 4684 2326
rect 4708 2270 4764 2326
rect 4788 2270 4844 2326
rect 4868 2270 4924 2326
rect 4948 2270 5004 2326
rect 5028 2270 5084 2326
rect 4228 2188 4284 2244
rect 4308 2188 4364 2244
rect 4388 2188 4444 2244
rect 4468 2188 4524 2244
rect 4548 2188 4604 2244
rect 4628 2188 4684 2244
rect 4708 2188 4764 2244
rect 4788 2188 4844 2244
rect 4868 2188 4924 2244
rect 4948 2188 5004 2244
rect 5028 2188 5084 2244
rect 4228 2106 4284 2162
rect 4308 2106 4364 2162
rect 4388 2106 4444 2162
rect 4468 2106 4524 2162
rect 4548 2106 4604 2162
rect 4628 2106 4684 2162
rect 4708 2106 4764 2162
rect 4788 2106 4844 2162
rect 4868 2106 4924 2162
rect 4948 2106 5004 2162
rect 5028 2106 5084 2162
rect 4228 2024 4284 2080
rect 4308 2024 4364 2080
rect 4388 2024 4444 2080
rect 4468 2024 4524 2080
rect 4548 2024 4604 2080
rect 4628 2024 4684 2080
rect 4708 2024 4764 2080
rect 4788 2024 4844 2080
rect 4868 2024 4924 2080
rect 4948 2024 5004 2080
rect 5028 2024 5084 2080
rect 4228 1942 4284 1998
rect 4308 1942 4364 1998
rect 4388 1942 4444 1998
rect 4468 1942 4524 1998
rect 4548 1942 4604 1998
rect 4628 1942 4684 1998
rect 4708 1942 4764 1998
rect 4788 1942 4844 1998
rect 4868 1942 4924 1998
rect 4948 1942 5004 1998
rect 5028 1942 5084 1998
rect 4228 1860 4284 1916
rect 4308 1860 4364 1916
rect 4388 1860 4444 1916
rect 4468 1860 4524 1916
rect 4548 1860 4604 1916
rect 4628 1860 4684 1916
rect 4708 1860 4764 1916
rect 4788 1860 4844 1916
rect 4868 1860 4924 1916
rect 4948 1860 5004 1916
rect 5028 1860 5084 1916
rect 6798 3093 6854 3149
rect 6884 3093 6940 3149
rect 6970 3093 7026 3149
rect 7056 3093 7112 3149
rect 7142 3093 7198 3149
rect 7228 3093 7284 3149
rect 7314 3093 7370 3149
rect 7400 3093 7456 3149
rect 7486 3093 7542 3149
rect 7572 3093 7628 3149
rect 7657 3093 7713 3149
rect 6798 3013 6854 3069
rect 6884 3013 6940 3069
rect 6970 3013 7026 3069
rect 7056 3013 7112 3069
rect 7142 3013 7198 3069
rect 7228 3013 7284 3069
rect 7314 3013 7370 3069
rect 7400 3013 7456 3069
rect 7486 3013 7542 3069
rect 7572 3013 7628 3069
rect 7657 3013 7713 3069
rect 6798 2933 6854 2989
rect 6884 2933 6940 2989
rect 6970 2933 7026 2989
rect 7056 2933 7112 2989
rect 7142 2933 7198 2989
rect 7228 2933 7284 2989
rect 7314 2933 7370 2989
rect 7400 2933 7456 2989
rect 7486 2933 7542 2989
rect 7572 2933 7628 2989
rect 7657 2933 7713 2989
rect 6798 2853 6854 2909
rect 6884 2853 6940 2909
rect 6970 2853 7026 2909
rect 7056 2853 7112 2909
rect 7142 2853 7198 2909
rect 7228 2853 7284 2909
rect 7314 2853 7370 2909
rect 7400 2853 7456 2909
rect 7486 2853 7542 2909
rect 7572 2853 7628 2909
rect 7657 2853 7713 2909
rect 6798 2773 6854 2829
rect 6884 2773 6940 2829
rect 6970 2773 7026 2829
rect 7056 2773 7112 2829
rect 7142 2773 7198 2829
rect 7228 2773 7284 2829
rect 7314 2773 7370 2829
rect 7400 2773 7456 2829
rect 7486 2773 7542 2829
rect 7572 2773 7628 2829
rect 7657 2773 7713 2829
rect 6798 2693 6854 2749
rect 6884 2693 6940 2749
rect 6970 2693 7026 2749
rect 7056 2693 7112 2749
rect 7142 2693 7198 2749
rect 7228 2693 7284 2749
rect 7314 2693 7370 2749
rect 7400 2693 7456 2749
rect 7486 2693 7542 2749
rect 7572 2693 7628 2749
rect 7657 2693 7713 2749
rect 6798 2613 6854 2669
rect 6884 2613 6940 2669
rect 6970 2613 7026 2669
rect 7056 2613 7112 2669
rect 7142 2613 7198 2669
rect 7228 2613 7284 2669
rect 7314 2613 7370 2669
rect 7400 2613 7456 2669
rect 7486 2613 7542 2669
rect 7572 2613 7628 2669
rect 7657 2613 7713 2669
rect 6798 2533 6854 2589
rect 6884 2533 6940 2589
rect 6970 2533 7026 2589
rect 7056 2533 7112 2589
rect 7142 2533 7198 2589
rect 7228 2533 7284 2589
rect 7314 2533 7370 2589
rect 7400 2533 7456 2589
rect 7486 2533 7542 2589
rect 7572 2533 7628 2589
rect 7657 2533 7713 2589
rect 3161 1637 3217 1693
rect 3241 1637 3297 1693
rect 3161 1545 3217 1601
rect 3241 1545 3297 1601
rect 3161 1452 3217 1508
rect 3241 1452 3297 1508
rect 3321 1474 3377 1530
rect 3401 1474 3457 1530
rect 3161 1359 3217 1415
rect 3241 1359 3297 1415
rect 3321 1362 3377 1418
rect 3401 1362 3457 1418
rect 2787 -752 3003 824
rect 7794 1775 7850 1831
rect 7874 1775 7930 1831
rect 7954 1775 8010 1831
rect 8034 1775 8090 1831
rect 8114 1775 8170 1831
rect 8194 1775 8250 1831
rect 7794 1692 7850 1748
rect 7874 1692 7930 1748
rect 7954 1692 8010 1748
rect 8034 1692 8090 1748
rect 8114 1692 8170 1748
rect 8194 1692 8250 1748
rect 7794 1609 7850 1665
rect 7874 1609 7930 1665
rect 7954 1609 8010 1665
rect 8034 1609 8090 1665
rect 8114 1609 8170 1665
rect 8194 1609 8250 1665
rect 7794 1526 7850 1582
rect 7874 1526 7930 1582
rect 7954 1526 8010 1582
rect 8034 1526 8090 1582
rect 8114 1526 8170 1582
rect 8194 1526 8250 1582
rect 7794 1442 7850 1498
rect 7874 1442 7930 1498
rect 7954 1442 8010 1498
rect 8034 1442 8090 1498
rect 8114 1442 8170 1498
rect 8194 1442 8250 1498
rect 7794 1358 7850 1414
rect 7874 1358 7930 1414
rect 7954 1358 8010 1414
rect 8034 1358 8090 1414
rect 8114 1358 8170 1414
rect 8194 1358 8250 1414
rect 8675 4076 8731 4132
rect 8755 4076 8811 4132
rect 8835 4076 8891 4132
rect 8915 4076 8971 4132
rect 8995 4076 9051 4132
rect 8675 3992 8731 4048
rect 8755 3992 8811 4048
rect 8835 3992 8891 4048
rect 8915 3992 8971 4048
rect 8995 3992 9051 4048
rect 8675 3908 8731 3964
rect 8755 3908 8811 3964
rect 8835 3908 8891 3964
rect 8915 3908 8971 3964
rect 8995 3908 9051 3964
rect 8675 3824 8731 3880
rect 8755 3824 8811 3880
rect 8835 3824 8891 3880
rect 8915 3824 8971 3880
rect 8995 3824 9051 3880
rect 8675 3739 8731 3795
rect 8755 3739 8811 3795
rect 8835 3739 8891 3795
rect 8915 3739 8971 3795
rect 8995 3739 9051 3795
rect 10609 3964 10825 4340
rect 10609 3883 10665 3939
rect 10689 3883 10745 3939
rect 10769 3883 10825 3939
rect 10609 3802 10665 3858
rect 10689 3802 10745 3858
rect 10769 3802 10825 3858
rect 10609 3721 10665 3777
rect 10689 3721 10745 3777
rect 10769 3721 10825 3777
rect 9602 3089 9658 3145
rect 9682 3089 9738 3145
rect 9762 3089 9818 3145
rect 9842 3089 9898 3145
rect 9922 3089 9978 3145
rect 10002 3089 10058 3145
rect 10082 3089 10138 3145
rect 10162 3089 10218 3145
rect 10242 3089 10298 3145
rect 9602 3002 9658 3058
rect 9682 3002 9738 3058
rect 9762 3002 9818 3058
rect 9842 3002 9898 3058
rect 9922 3002 9978 3058
rect 10002 3002 10058 3058
rect 10082 3002 10138 3058
rect 10162 3002 10218 3058
rect 10242 3002 10298 3058
rect 9602 2915 9658 2971
rect 9682 2915 9738 2971
rect 9762 2915 9818 2971
rect 9842 2915 9898 2971
rect 9922 2915 9978 2971
rect 10002 2915 10058 2971
rect 10082 2915 10138 2971
rect 10162 2915 10218 2971
rect 10242 2915 10298 2971
rect 9602 2828 9658 2884
rect 9682 2828 9738 2884
rect 9762 2828 9818 2884
rect 9842 2828 9898 2884
rect 9922 2828 9978 2884
rect 10002 2828 10058 2884
rect 10082 2828 10138 2884
rect 10162 2828 10218 2884
rect 10242 2828 10298 2884
rect 9602 2741 9658 2797
rect 9682 2741 9738 2797
rect 9762 2741 9818 2797
rect 9842 2741 9898 2797
rect 9922 2741 9978 2797
rect 10002 2741 10058 2797
rect 10082 2741 10138 2797
rect 10162 2741 10218 2797
rect 10242 2741 10298 2797
rect 9602 2654 9658 2710
rect 9682 2654 9738 2710
rect 9762 2654 9818 2710
rect 9842 2654 9898 2710
rect 9922 2654 9978 2710
rect 10002 2654 10058 2710
rect 10082 2654 10138 2710
rect 10162 2654 10218 2710
rect 10242 2654 10298 2710
rect 9602 2567 9658 2623
rect 9682 2567 9738 2623
rect 9762 2567 9818 2623
rect 9842 2567 9898 2623
rect 9922 2567 9978 2623
rect 10002 2567 10058 2623
rect 10082 2567 10138 2623
rect 10162 2567 10218 2623
rect 10242 2567 10298 2623
rect 9602 2480 9658 2536
rect 9682 2480 9738 2536
rect 9762 2480 9818 2536
rect 9842 2480 9898 2536
rect 9922 2480 9978 2536
rect 10002 2480 10058 2536
rect 10082 2480 10138 2536
rect 10162 2480 10218 2536
rect 10242 2480 10298 2536
rect 9602 2392 9658 2448
rect 9682 2392 9738 2448
rect 9762 2392 9818 2448
rect 9842 2392 9898 2448
rect 9922 2392 9978 2448
rect 10002 2392 10058 2448
rect 10082 2392 10138 2448
rect 10162 2392 10218 2448
rect 10242 2392 10298 2448
rect 9602 2304 9658 2360
rect 9682 2304 9738 2360
rect 9762 2304 9818 2360
rect 9842 2304 9898 2360
rect 9922 2304 9978 2360
rect 10002 2304 10058 2360
rect 10082 2304 10138 2360
rect 10162 2304 10218 2360
rect 10242 2304 10298 2360
rect 9602 2216 9658 2272
rect 9682 2216 9738 2272
rect 9762 2216 9818 2272
rect 9842 2216 9898 2272
rect 9922 2216 9978 2272
rect 10002 2216 10058 2272
rect 10082 2216 10138 2272
rect 10162 2216 10218 2272
rect 10242 2216 10298 2272
rect 9735 1993 9791 2049
rect 9815 1993 9871 2049
rect 9895 1993 9951 2049
rect 9735 1903 9791 1959
rect 9815 1903 9871 1959
rect 9895 1903 9951 1959
rect 9735 1813 9791 1869
rect 9815 1813 9871 1869
rect 9895 1813 9951 1869
rect 9735 1723 9791 1779
rect 9815 1723 9871 1779
rect 9895 1723 9951 1779
rect 9735 1633 9791 1689
rect 9815 1633 9871 1689
rect 9895 1633 9951 1689
rect 9735 1543 9791 1599
rect 9815 1543 9871 1599
rect 9895 1543 9951 1599
rect 9735 1453 9791 1509
rect 9815 1453 9871 1509
rect 9895 1453 9951 1509
rect 9735 1362 9791 1418
rect 9815 1362 9871 1418
rect 9895 1362 9951 1418
rect 2787 -833 2843 -777
rect 2867 -833 2923 -777
rect 2947 -833 3003 -777
rect 2787 -914 2843 -858
rect 2867 -914 2923 -858
rect 2947 -914 3003 -858
rect 2787 -995 2843 -939
rect 2867 -995 2923 -939
rect 2947 -995 3003 -939
rect 2787 -1076 2843 -1020
rect 2867 -1076 2923 -1020
rect 2947 -1076 3003 -1020
rect 2787 -1146 2816 -1101
rect 2816 -1146 2837 -1101
rect 2837 -1146 2843 -1101
rect 2867 -1146 2889 -1101
rect 2889 -1146 2910 -1101
rect 2910 -1146 2923 -1101
rect 2947 -1146 2962 -1101
rect 2962 -1146 2982 -1101
rect 2982 -1146 3003 -1101
rect 2787 -1157 2843 -1146
rect 2867 -1157 2923 -1146
rect 2947 -1157 3003 -1146
rect 2787 -1210 2816 -1182
rect 2816 -1210 2837 -1182
rect 2837 -1210 2843 -1182
rect 2867 -1210 2889 -1182
rect 2889 -1210 2910 -1182
rect 2910 -1210 2923 -1182
rect 2947 -1210 2962 -1182
rect 2962 -1210 2982 -1182
rect 2982 -1210 3003 -1182
rect 2787 -1222 2843 -1210
rect 2867 -1222 2923 -1210
rect 2947 -1222 3003 -1210
rect 2787 -1238 2816 -1222
rect 2816 -1238 2837 -1222
rect 2837 -1238 2843 -1222
rect 2867 -1238 2889 -1222
rect 2889 -1238 2910 -1222
rect 2910 -1238 2923 -1222
rect 2947 -1238 2962 -1222
rect 2962 -1238 2982 -1222
rect 2982 -1238 3003 -1222
rect 2787 -1274 2816 -1263
rect 2816 -1274 2837 -1263
rect 2837 -1274 2843 -1263
rect 2867 -1274 2889 -1263
rect 2889 -1274 2910 -1263
rect 2910 -1274 2923 -1263
rect 2947 -1274 2962 -1263
rect 2962 -1274 2982 -1263
rect 2982 -1274 3003 -1263
rect 2787 -1319 2843 -1274
rect 2867 -1319 2923 -1274
rect 2947 -1319 3003 -1274
rect 2787 -1400 2843 -1344
rect 2867 -1400 2923 -1344
rect 2947 -1400 3003 -1344
rect 2787 -1481 2843 -1425
rect 2867 -1481 2923 -1425
rect 2947 -1481 3003 -1425
rect 2787 -1562 2843 -1506
rect 2867 -1562 2923 -1506
rect 2947 -1562 3003 -1506
rect 2787 -1627 2813 -1587
rect 2813 -1627 2835 -1587
rect 2835 -1627 2843 -1587
rect 2867 -1627 2887 -1587
rect 2887 -1627 2909 -1587
rect 2909 -1627 2923 -1587
rect 2947 -1627 2961 -1587
rect 2961 -1627 2983 -1587
rect 2983 -1627 3003 -1587
rect 2787 -1639 2843 -1627
rect 2867 -1639 2923 -1627
rect 2947 -1639 3003 -1627
rect 2787 -1643 2813 -1639
rect 2813 -1643 2835 -1639
rect 2835 -1643 2843 -1639
rect 2867 -1643 2887 -1639
rect 2887 -1643 2909 -1639
rect 2909 -1643 2923 -1639
rect 2947 -1643 2961 -1639
rect 2961 -1643 2983 -1639
rect 2983 -1643 3003 -1639
rect 2787 -1691 2813 -1668
rect 2813 -1691 2835 -1668
rect 2835 -1691 2843 -1668
rect 2867 -1691 2887 -1668
rect 2887 -1691 2909 -1668
rect 2909 -1691 2923 -1668
rect 2947 -1691 2961 -1668
rect 2961 -1691 2983 -1668
rect 2983 -1691 3003 -1668
rect 2787 -1724 2843 -1691
rect 2867 -1724 2923 -1691
rect 2947 -1724 3003 -1691
rect 2787 -1805 2843 -1749
rect 2867 -1805 2923 -1749
rect 2947 -1805 3003 -1749
rect 2787 -1886 2843 -1830
rect 2867 -1886 2923 -1830
rect 2947 -1886 3003 -1830
rect 10386 771 10442 827
rect 10466 771 10522 827
rect 10546 771 10602 827
rect 10626 771 10682 827
rect 10706 771 10762 827
rect 10786 771 10842 827
rect 10386 684 10442 740
rect 10466 684 10522 740
rect 10546 684 10602 740
rect 10626 684 10682 740
rect 10706 684 10762 740
rect 10786 684 10842 740
rect 10386 596 10442 652
rect 10466 596 10522 652
rect 10546 596 10602 652
rect 10626 596 10682 652
rect 10706 596 10762 652
rect 10786 596 10842 652
rect 10386 508 10442 564
rect 10466 508 10522 564
rect 10546 508 10602 564
rect 10626 508 10682 564
rect 10706 508 10762 564
rect 10786 508 10842 564
rect 10386 420 10442 476
rect 10466 420 10522 476
rect 10546 420 10602 476
rect 10626 420 10682 476
rect 10706 420 10762 476
rect 10786 420 10842 476
rect 10386 332 10442 388
rect 10466 332 10522 388
rect 10546 332 10602 388
rect 10626 332 10682 388
rect 10706 332 10762 388
rect 10786 332 10842 388
rect 10386 244 10442 300
rect 10466 244 10522 300
rect 10546 244 10602 300
rect 10626 244 10682 300
rect 10706 244 10762 300
rect 10786 244 10842 300
rect 12194 2494 12650 3190
rect 12194 2413 12250 2469
rect 12274 2413 12330 2469
rect 12354 2413 12410 2469
rect 12434 2413 12490 2469
rect 12514 2413 12570 2469
rect 12594 2413 12650 2469
rect 12194 2332 12250 2388
rect 12274 2332 12330 2388
rect 12354 2332 12410 2388
rect 12434 2332 12490 2388
rect 12514 2332 12570 2388
rect 12594 2332 12650 2388
rect 12194 2251 12250 2307
rect 12274 2251 12330 2307
rect 12354 2251 12410 2307
rect 12434 2251 12490 2307
rect 12514 2251 12570 2307
rect 12594 2251 12650 2307
rect 12194 2170 12250 2226
rect 12274 2170 12330 2226
rect 12354 2170 12410 2226
rect 12434 2170 12490 2226
rect 12514 2170 12570 2226
rect 12594 2170 12650 2226
rect 12194 2089 12250 2145
rect 12274 2089 12330 2145
rect 12354 2089 12410 2145
rect 12434 2089 12490 2145
rect 12514 2089 12570 2145
rect 12594 2089 12650 2145
rect 12194 2008 12250 2064
rect 12274 2008 12330 2064
rect 12354 2008 12410 2064
rect 12434 2008 12490 2064
rect 12514 2008 12570 2064
rect 12594 2008 12650 2064
rect 12194 1927 12250 1983
rect 12274 1927 12330 1983
rect 12354 1927 12410 1983
rect 12434 1927 12490 1983
rect 12514 1927 12570 1983
rect 12594 1927 12650 1983
rect 12194 1846 12250 1902
rect 12274 1846 12330 1902
rect 12354 1846 12410 1902
rect 12434 1846 12490 1902
rect 12514 1846 12570 1902
rect 12594 1846 12650 1902
rect 12194 1765 12250 1821
rect 12274 1765 12330 1821
rect 12354 1765 12410 1821
rect 12434 1765 12490 1821
rect 12514 1765 12570 1821
rect 12594 1765 12650 1821
rect 12194 1684 12250 1740
rect 12274 1684 12330 1740
rect 12354 1684 12410 1740
rect 12434 1684 12490 1740
rect 12514 1684 12570 1740
rect 12594 1684 12650 1740
rect 12194 1603 12250 1659
rect 12274 1603 12330 1659
rect 12354 1603 12410 1659
rect 12434 1603 12490 1659
rect 12514 1603 12570 1659
rect 12594 1603 12650 1659
rect 12194 1522 12250 1578
rect 12274 1522 12330 1578
rect 12354 1522 12410 1578
rect 12434 1522 12490 1578
rect 12514 1522 12570 1578
rect 12594 1522 12650 1578
rect 12194 1441 12250 1497
rect 12274 1441 12330 1497
rect 12354 1441 12410 1497
rect 12434 1441 12490 1497
rect 12514 1441 12570 1497
rect 12594 1441 12650 1497
rect 12194 1360 12250 1416
rect 12274 1360 12330 1416
rect 12354 1360 12410 1416
rect 12434 1360 12490 1416
rect 12514 1360 12570 1416
rect 12594 1360 12650 1416
rect 2787 -1967 2843 -1911
rect 2867 -1967 2923 -1911
rect 2947 -1967 3003 -1911
rect 13307 4044 13363 4100
rect 13392 4044 13448 4100
rect 13476 4044 13532 4100
rect 13560 4044 13616 4100
rect 13644 4044 13700 4100
rect 13728 4044 13784 4100
rect 13812 4044 13868 4100
rect 13307 3964 13363 4020
rect 13392 3964 13448 4020
rect 13476 3964 13532 4020
rect 13560 3964 13616 4020
rect 13644 3964 13700 4020
rect 13728 3964 13784 4020
rect 13812 3964 13868 4020
rect 13307 3884 13363 3940
rect 13392 3884 13448 3940
rect 13476 3884 13532 3940
rect 13560 3884 13616 3940
rect 13644 3884 13700 3940
rect 13728 3884 13784 3940
rect 13812 3884 13868 3940
rect 13307 3804 13363 3860
rect 13392 3804 13448 3860
rect 13476 3804 13532 3860
rect 13560 3804 13616 3860
rect 13644 3804 13700 3860
rect 13728 3804 13784 3860
rect 13812 3804 13868 3860
rect 13307 3724 13363 3780
rect 13392 3724 13448 3780
rect 13476 3724 13532 3780
rect 13560 3724 13616 3780
rect 13644 3724 13700 3780
rect 13728 3724 13784 3780
rect 13812 3724 13868 3780
rect 13972 3103 14028 3159
rect 14063 3103 14119 3159
rect 14154 3103 14210 3159
rect 14244 3103 14300 3159
rect 14334 3103 14390 3159
rect 14424 3103 14480 3159
rect 14514 3103 14570 3159
rect 14630 3089 14686 3145
rect 14718 3089 14774 3145
rect 14806 3089 14862 3145
rect 14894 3089 14950 3145
rect 14982 3089 15038 3145
rect 15070 3089 15126 3145
rect 15158 3089 15214 3145
rect 13972 3023 14028 3079
rect 14063 3023 14119 3079
rect 14154 3023 14210 3079
rect 14244 3023 14300 3079
rect 14334 3023 14390 3079
rect 14424 3023 14480 3079
rect 14514 3023 14570 3079
rect 14630 3009 14686 3065
rect 14718 3009 14774 3065
rect 14806 3009 14862 3065
rect 14894 3009 14950 3065
rect 14982 3009 15038 3065
rect 15070 3009 15126 3065
rect 15158 3009 15214 3065
rect 13972 2943 14028 2999
rect 14063 2943 14119 2999
rect 14154 2943 14210 2999
rect 14244 2943 14300 2999
rect 14334 2943 14390 2999
rect 14424 2943 14480 2999
rect 14514 2943 14570 2999
rect 14630 2929 14686 2985
rect 14718 2929 14774 2985
rect 14806 2929 14862 2985
rect 14894 2929 14950 2985
rect 14982 2929 15038 2985
rect 15070 2929 15126 2985
rect 15158 2929 15214 2985
rect 13972 2863 14028 2919
rect 14063 2863 14119 2919
rect 14154 2863 14210 2919
rect 14244 2863 14300 2919
rect 14334 2863 14390 2919
rect 14424 2863 14480 2919
rect 14514 2863 14570 2919
rect 14630 2849 14686 2905
rect 14718 2849 14774 2905
rect 14806 2849 14862 2905
rect 14894 2849 14950 2905
rect 14982 2849 15038 2905
rect 15070 2849 15126 2905
rect 15158 2849 15214 2905
rect 13972 2783 14028 2839
rect 14063 2783 14119 2839
rect 14154 2783 14210 2839
rect 14244 2783 14300 2839
rect 14334 2783 14390 2839
rect 14424 2783 14480 2839
rect 14514 2783 14570 2839
rect 13972 2703 14028 2759
rect 14063 2703 14119 2759
rect 14154 2703 14210 2759
rect 14244 2703 14300 2759
rect 14334 2703 14390 2759
rect 14424 2703 14480 2759
rect 14514 2703 14570 2759
rect 14641 2733 14697 2789
rect 14721 2733 14777 2789
rect 14801 2733 14857 2789
rect 13972 2623 14028 2679
rect 14063 2623 14119 2679
rect 14154 2623 14210 2679
rect 14244 2623 14300 2679
rect 14334 2623 14390 2679
rect 14424 2623 14480 2679
rect 14514 2623 14570 2679
rect 14641 2621 14697 2677
rect 14721 2621 14777 2677
rect 14801 2621 14857 2677
rect 13972 2543 14028 2599
rect 14063 2543 14119 2599
rect 14154 2543 14210 2599
rect 14244 2543 14300 2599
rect 14334 2543 14390 2599
rect 14424 2543 14480 2599
rect 14514 2543 14570 2599
rect 13972 2463 14028 2519
rect 14063 2463 14119 2519
rect 14154 2463 14210 2519
rect 14244 2463 14300 2519
rect 14334 2463 14390 2519
rect 14424 2463 14480 2519
rect 14514 2463 14570 2519
rect 14641 2508 14697 2564
rect 14721 2508 14777 2564
rect 14801 2508 14857 2564
rect 16064 4513 16120 4569
rect 16144 4513 16200 4569
rect 16224 4513 16280 4569
rect 16304 4513 16360 4569
rect 16384 4513 16440 4569
rect 16464 4513 16520 4569
rect 20888 13307 21104 14803
rect 20888 13226 20944 13282
rect 20968 13226 21024 13282
rect 21048 13226 21104 13282
rect 20888 13145 20944 13201
rect 20968 13145 21024 13201
rect 21048 13145 21104 13201
rect 20888 13064 20944 13120
rect 20968 13064 21024 13120
rect 21048 13064 21104 13120
rect 20888 12983 20944 13039
rect 20968 12983 21024 13039
rect 21048 12983 21104 13039
rect 20888 12902 20944 12958
rect 20968 12902 21024 12958
rect 21048 12902 21104 12958
rect 20888 12821 20944 12877
rect 20968 12821 21024 12877
rect 21048 12821 21104 12877
rect 20888 12740 20944 12796
rect 20968 12740 21024 12796
rect 21048 12740 21104 12796
rect 20888 12659 20944 12715
rect 20968 12659 21024 12715
rect 21048 12659 21104 12715
rect 20888 12578 20944 12634
rect 20968 12578 21024 12634
rect 21048 12578 21104 12634
rect 20888 12497 20944 12553
rect 20968 12497 21024 12553
rect 21048 12497 21104 12553
rect 20888 12416 20944 12472
rect 20968 12416 21024 12472
rect 21048 12416 21104 12472
rect 20888 12335 20944 12391
rect 20968 12335 21024 12391
rect 21048 12335 21104 12391
rect 20888 12254 20944 12310
rect 20968 12254 21024 12310
rect 21048 12254 21104 12310
rect 20888 12173 20944 12229
rect 20968 12173 21024 12229
rect 21048 12173 21104 12229
rect 20888 12092 20944 12148
rect 20968 12092 21024 12148
rect 21048 12092 21104 12148
rect 20888 12011 20944 12067
rect 20968 12011 21024 12067
rect 21048 12011 21104 12067
rect 20888 11930 20944 11986
rect 20968 11930 21024 11986
rect 21048 11930 21104 11986
rect 20888 11849 20944 11905
rect 20968 11849 21024 11905
rect 21048 11849 21104 11905
rect 20888 11768 20944 11824
rect 20968 11768 21024 11824
rect 21048 11768 21104 11824
rect 20888 11687 20944 11743
rect 20968 11687 21024 11743
rect 21048 11687 21104 11743
rect 20888 11606 20944 11662
rect 20968 11606 21024 11662
rect 21048 11606 21104 11662
rect 20888 11525 20944 11581
rect 20968 11525 21024 11581
rect 21048 11525 21104 11581
rect 20888 11444 20944 11500
rect 20968 11444 21024 11500
rect 21048 11444 21104 11500
rect 20888 11363 20944 11419
rect 20968 11363 21024 11419
rect 21048 11363 21104 11419
rect 20888 11282 20944 11338
rect 20968 11282 21024 11338
rect 21048 11282 21104 11338
rect 20888 11201 20944 11257
rect 20968 11201 21024 11257
rect 21048 11201 21104 11257
rect 20888 11120 20944 11176
rect 20968 11120 21024 11176
rect 21048 11120 21104 11176
rect 20888 11039 20944 11095
rect 20968 11039 21024 11095
rect 21048 11039 21104 11095
rect 20888 10958 20944 11014
rect 20968 10958 21024 11014
rect 21048 10958 21104 11014
rect 20888 10877 20944 10933
rect 20968 10877 21024 10933
rect 21048 10877 21104 10933
rect 20888 10796 20944 10852
rect 20968 10796 21024 10852
rect 21048 10796 21104 10852
rect 20888 10715 20944 10771
rect 20968 10715 21024 10771
rect 21048 10715 21104 10771
rect 20888 10634 20944 10690
rect 20968 10634 21024 10690
rect 21048 10634 21104 10690
rect 20888 10553 20944 10609
rect 20968 10553 21024 10609
rect 21048 10553 21104 10609
rect 20888 10472 20944 10528
rect 20968 10472 21024 10528
rect 21048 10472 21104 10528
rect 20888 10391 20944 10447
rect 20968 10391 21024 10447
rect 21048 10391 21104 10447
rect 20888 10310 20944 10366
rect 20968 10310 21024 10366
rect 21048 10310 21104 10366
rect 20888 10229 20944 10285
rect 20968 10229 21024 10285
rect 21048 10229 21104 10285
rect 20888 10148 20944 10204
rect 20968 10148 21024 10204
rect 21048 10148 21104 10204
rect 20888 10067 20944 10123
rect 20968 10067 21024 10123
rect 21048 10067 21104 10123
rect 20888 9986 20944 10042
rect 20968 9986 21024 10042
rect 21048 9986 21104 10042
rect 20888 9905 20944 9961
rect 20968 9905 21024 9961
rect 21048 9905 21104 9961
rect 20888 9824 20944 9880
rect 20968 9824 21024 9880
rect 21048 9824 21104 9880
rect 20888 9743 20944 9799
rect 20968 9743 21024 9799
rect 21048 9743 21104 9799
rect 20888 9662 20944 9718
rect 20968 9662 21024 9718
rect 21048 9662 21104 9718
rect 20888 9581 20944 9637
rect 20968 9581 21024 9637
rect 21048 9581 21104 9637
rect 20888 9500 20944 9556
rect 20968 9500 21024 9556
rect 21048 9500 21104 9556
rect 20888 9419 20944 9475
rect 20968 9419 21024 9475
rect 21048 9419 21104 9475
rect 20888 9338 20944 9394
rect 20968 9338 21024 9394
rect 21048 9338 21104 9394
rect 20888 9257 20944 9313
rect 20968 9257 21024 9313
rect 21048 9257 21104 9313
rect 20888 9176 20944 9232
rect 20968 9176 21024 9232
rect 21048 9176 21104 9232
rect 20888 9095 20944 9151
rect 20968 9095 21024 9151
rect 21048 9095 21104 9151
rect 20888 9014 20944 9070
rect 20968 9014 21024 9070
rect 21048 9014 21104 9070
rect 20888 8933 20944 8989
rect 20968 8933 21024 8989
rect 21048 8933 21104 8989
rect 20888 8852 20944 8908
rect 20968 8852 21024 8908
rect 21048 8852 21104 8908
rect 20888 8771 20944 8827
rect 20968 8771 21024 8827
rect 21048 8771 21104 8827
rect 20888 8690 20944 8746
rect 20968 8690 21024 8746
rect 21048 8690 21104 8746
rect 20888 8609 20944 8665
rect 20968 8609 21024 8665
rect 21048 8609 21104 8665
rect 20888 8528 20944 8584
rect 20968 8528 21024 8584
rect 21048 8528 21104 8584
rect 20888 8447 20944 8503
rect 20968 8447 21024 8503
rect 21048 8447 21104 8503
rect 20888 8366 20944 8422
rect 20968 8366 21024 8422
rect 21048 8366 21104 8422
rect 20888 8285 20944 8341
rect 20968 8285 21024 8341
rect 21048 8285 21104 8341
rect 20888 8204 20944 8260
rect 20968 8204 21024 8260
rect 21048 8204 21104 8260
rect 20888 8123 20944 8179
rect 20968 8123 21024 8179
rect 21048 8123 21104 8179
rect 20888 8083 20944 8098
rect 20968 8083 21024 8098
rect 21048 8083 21104 8098
rect 20888 8042 20896 8083
rect 20896 8042 20926 8083
rect 20926 8042 20944 8083
rect 20968 8042 20978 8083
rect 20978 8042 21008 8083
rect 21008 8042 21024 8083
rect 21048 8042 21060 8083
rect 21060 8042 21090 8083
rect 21090 8042 21104 8083
rect 20888 7967 20896 8017
rect 20896 7967 20926 8017
rect 20926 7967 20944 8017
rect 20968 7967 20978 8017
rect 20978 7967 21008 8017
rect 21008 7967 21024 8017
rect 21048 7967 21060 8017
rect 21060 7967 21090 8017
rect 21090 7967 21104 8017
rect 20888 7961 20944 7967
rect 20968 7961 21024 7967
rect 21048 7961 21104 7967
rect 20888 7903 20896 7936
rect 20896 7903 20926 7936
rect 20926 7903 20944 7936
rect 20968 7903 20978 7936
rect 20978 7903 21008 7936
rect 21008 7903 21024 7936
rect 21048 7903 21060 7936
rect 21060 7903 21090 7936
rect 21090 7903 21104 7936
rect 20888 7880 20944 7903
rect 20968 7880 21024 7903
rect 21048 7880 21104 7903
rect 13972 2383 14028 2439
rect 14063 2383 14119 2439
rect 14154 2383 14210 2439
rect 14244 2383 14300 2439
rect 14334 2383 14390 2439
rect 14424 2383 14480 2439
rect 14514 2383 14570 2439
rect 13972 2303 14028 2359
rect 14063 2303 14119 2359
rect 14154 2303 14210 2359
rect 14244 2303 14300 2359
rect 14334 2303 14390 2359
rect 14424 2303 14480 2359
rect 14514 2303 14570 2359
rect 13972 2223 14028 2279
rect 14063 2223 14119 2279
rect 14154 2223 14210 2279
rect 14244 2223 14300 2279
rect 14334 2223 14390 2279
rect 14424 2223 14480 2279
rect 14514 2223 14570 2279
rect 13320 776 13376 832
rect 13400 776 13456 832
rect 13480 776 13536 832
rect 13560 776 13616 832
rect 13640 776 13696 832
rect 13320 690 13376 746
rect 13400 690 13456 746
rect 13720 738 13776 794
rect 13480 681 13536 737
rect 13560 674 13616 730
rect 13320 604 13376 660
rect 13400 604 13456 660
rect 13640 650 13696 706
rect 15380 1582 15436 1638
rect 15460 1582 15516 1638
rect 15540 1582 15596 1638
rect 15380 1474 15436 1530
rect 15460 1474 15516 1530
rect 15540 1474 15596 1530
rect 15380 1365 15436 1421
rect 15460 1365 15516 1421
rect 15540 1365 15596 1421
rect 15650 1359 15946 1895
rect 13480 585 13536 641
rect 13320 518 13376 574
rect 13400 518 13456 574
rect 13560 572 13616 628
rect 13480 489 13536 545
rect 13320 431 13376 487
rect 13400 431 13456 487
rect 9728 -2927 9784 -2871
rect 9808 -2927 9864 -2871
rect 9888 -2927 9944 -2871
rect 9728 -3011 9784 -2955
rect 9808 -3011 9864 -2955
rect 9888 -3011 9944 -2955
rect 9728 -3095 9784 -3039
rect 9808 -3095 9864 -3039
rect 9888 -3095 9944 -3039
rect 9728 -3179 9784 -3123
rect 9808 -3179 9864 -3123
rect 9888 -3179 9944 -3123
rect 9728 -3263 9784 -3207
rect 9808 -3263 9864 -3207
rect 9888 -3263 9944 -3207
rect 9728 -3347 9784 -3291
rect 9808 -3347 9864 -3291
rect 9888 -3347 9944 -3291
rect 9728 -3431 9784 -3375
rect 9808 -3431 9864 -3375
rect 9888 -3431 9944 -3375
rect 9728 -3515 9784 -3459
rect 9808 -3515 9864 -3459
rect 9888 -3515 9944 -3459
rect 9728 -3599 9784 -3543
rect 9808 -3599 9864 -3543
rect 9888 -3599 9944 -3543
rect 9728 -3684 9784 -3628
rect 9808 -3684 9864 -3628
rect 9888 -3684 9944 -3628
rect 21641 8425 21937 14801
rect 29488 17953 29544 18009
rect 29568 17953 29624 18009
rect 29648 17953 29704 18009
rect 29728 17953 29784 18009
rect 26328 17858 26384 17914
rect 26416 17858 26472 17914
rect 26504 17858 26560 17914
rect 26328 17778 26384 17834
rect 26416 17778 26472 17834
rect 26504 17778 26560 17834
rect 29488 17866 29544 17922
rect 29568 17866 29624 17922
rect 29648 17866 29704 17922
rect 29728 17866 29784 17922
rect 29488 17779 29544 17835
rect 29568 17779 29624 17835
rect 29648 17779 29704 17835
rect 29728 17779 29784 17835
rect 31022 18791 31078 18804
rect 31102 18791 31158 18804
rect 31182 18791 31238 18804
rect 31262 18791 31318 18804
rect 31342 18791 31398 18804
rect 31022 18748 31029 18791
rect 31029 18748 31078 18791
rect 31102 18748 31145 18791
rect 31145 18748 31157 18791
rect 31157 18748 31158 18791
rect 31182 18748 31209 18791
rect 31209 18748 31221 18791
rect 31221 18748 31238 18791
rect 31262 18748 31273 18791
rect 31273 18748 31285 18791
rect 31285 18748 31318 18791
rect 31342 18748 31349 18791
rect 31349 18748 31398 18791
rect 31022 18672 31029 18723
rect 31029 18672 31078 18723
rect 31102 18672 31145 18723
rect 31145 18672 31157 18723
rect 31157 18672 31158 18723
rect 31182 18672 31209 18723
rect 31209 18672 31221 18723
rect 31221 18672 31238 18723
rect 31262 18672 31273 18723
rect 31273 18672 31285 18723
rect 31285 18672 31318 18723
rect 31342 18672 31349 18723
rect 31349 18672 31398 18723
rect 31022 18667 31078 18672
rect 31102 18667 31158 18672
rect 31182 18667 31238 18672
rect 31262 18667 31318 18672
rect 31342 18667 31398 18672
rect 31022 18605 31029 18642
rect 31029 18605 31078 18642
rect 31102 18605 31145 18642
rect 31145 18605 31157 18642
rect 31157 18605 31158 18642
rect 31182 18605 31209 18642
rect 31209 18605 31221 18642
rect 31221 18605 31238 18642
rect 31262 18605 31273 18642
rect 31273 18605 31285 18642
rect 31285 18605 31318 18642
rect 31342 18605 31349 18642
rect 31349 18605 31398 18642
rect 31022 18590 31078 18605
rect 31102 18590 31158 18605
rect 31182 18590 31238 18605
rect 31262 18590 31318 18605
rect 31342 18590 31398 18605
rect 31022 18586 31029 18590
rect 31029 18586 31078 18590
rect 31022 18538 31029 18561
rect 31029 18538 31078 18561
rect 31102 18586 31145 18590
rect 31145 18586 31157 18590
rect 31157 18586 31158 18590
rect 31182 18586 31209 18590
rect 31209 18586 31221 18590
rect 31221 18586 31238 18590
rect 31262 18586 31273 18590
rect 31273 18586 31285 18590
rect 31285 18586 31318 18590
rect 31342 18586 31349 18590
rect 31349 18586 31398 18590
rect 31102 18538 31145 18561
rect 31145 18538 31157 18561
rect 31157 18538 31158 18561
rect 31182 18538 31209 18561
rect 31209 18538 31221 18561
rect 31221 18538 31238 18561
rect 31262 18538 31273 18561
rect 31273 18538 31285 18561
rect 31285 18538 31318 18561
rect 31342 18538 31349 18561
rect 31349 18538 31398 18561
rect 31022 18523 31078 18538
rect 31102 18523 31158 18538
rect 31182 18523 31238 18538
rect 31262 18523 31318 18538
rect 31342 18523 31398 18538
rect 31022 18505 31029 18523
rect 31029 18505 31078 18523
rect 31022 18471 31029 18480
rect 31029 18471 31078 18480
rect 31102 18505 31145 18523
rect 31145 18505 31157 18523
rect 31157 18505 31158 18523
rect 31182 18505 31209 18523
rect 31209 18505 31221 18523
rect 31221 18505 31238 18523
rect 31262 18505 31273 18523
rect 31273 18505 31285 18523
rect 31285 18505 31318 18523
rect 31342 18505 31349 18523
rect 31349 18505 31398 18523
rect 31102 18471 31145 18480
rect 31145 18471 31157 18480
rect 31157 18471 31158 18480
rect 31182 18471 31209 18480
rect 31209 18471 31221 18480
rect 31221 18471 31238 18480
rect 31262 18471 31273 18480
rect 31273 18471 31285 18480
rect 31285 18471 31318 18480
rect 31342 18471 31349 18480
rect 31349 18471 31398 18480
rect 31022 18456 31078 18471
rect 31102 18456 31158 18471
rect 31182 18456 31238 18471
rect 31262 18456 31318 18471
rect 31342 18456 31398 18471
rect 31022 18424 31029 18456
rect 31029 18424 31078 18456
rect 31102 18424 31145 18456
rect 31145 18424 31157 18456
rect 31157 18424 31158 18456
rect 31182 18424 31209 18456
rect 31209 18424 31221 18456
rect 31221 18424 31238 18456
rect 31262 18424 31273 18456
rect 31273 18424 31285 18456
rect 31285 18424 31318 18456
rect 31342 18424 31349 18456
rect 31349 18424 31398 18456
rect 31022 18389 31078 18398
rect 31102 18389 31158 18398
rect 31182 18389 31238 18398
rect 31262 18389 31318 18398
rect 31342 18389 31398 18398
rect 31022 18342 31029 18389
rect 31029 18342 31078 18389
rect 31102 18342 31145 18389
rect 31145 18342 31157 18389
rect 31157 18342 31158 18389
rect 31182 18342 31209 18389
rect 31209 18342 31221 18389
rect 31221 18342 31238 18389
rect 31262 18342 31273 18389
rect 31273 18342 31285 18389
rect 31285 18342 31318 18389
rect 31342 18342 31349 18389
rect 31349 18342 31398 18389
rect 31022 18270 31029 18316
rect 31029 18270 31078 18316
rect 31102 18270 31145 18316
rect 31145 18270 31157 18316
rect 31157 18270 31158 18316
rect 31182 18270 31209 18316
rect 31209 18270 31221 18316
rect 31221 18270 31238 18316
rect 31262 18270 31273 18316
rect 31273 18270 31285 18316
rect 31285 18270 31318 18316
rect 31342 18270 31349 18316
rect 31349 18270 31398 18316
rect 31022 18260 31078 18270
rect 31102 18260 31158 18270
rect 31182 18260 31238 18270
rect 31262 18260 31318 18270
rect 31342 18260 31398 18270
rect 31022 18203 31029 18234
rect 31029 18203 31078 18234
rect 31102 18203 31145 18234
rect 31145 18203 31157 18234
rect 31157 18203 31158 18234
rect 31182 18203 31209 18234
rect 31209 18203 31221 18234
rect 31221 18203 31238 18234
rect 31262 18203 31273 18234
rect 31273 18203 31285 18234
rect 31285 18203 31318 18234
rect 31342 18203 31349 18234
rect 31349 18203 31398 18234
rect 31022 18188 31078 18203
rect 31102 18188 31158 18203
rect 31182 18188 31238 18203
rect 31262 18188 31318 18203
rect 31342 18188 31398 18203
rect 31022 18178 31029 18188
rect 31029 18178 31078 18188
rect 31022 18136 31029 18152
rect 31029 18136 31078 18152
rect 31102 18178 31145 18188
rect 31145 18178 31157 18188
rect 31157 18178 31158 18188
rect 31182 18178 31209 18188
rect 31209 18178 31221 18188
rect 31221 18178 31238 18188
rect 31262 18178 31273 18188
rect 31273 18178 31285 18188
rect 31285 18178 31318 18188
rect 31342 18178 31349 18188
rect 31349 18178 31398 18188
rect 31102 18136 31145 18152
rect 31145 18136 31157 18152
rect 31157 18136 31158 18152
rect 31182 18136 31209 18152
rect 31209 18136 31221 18152
rect 31221 18136 31238 18152
rect 31262 18136 31273 18152
rect 31273 18136 31285 18152
rect 31285 18136 31318 18152
rect 31342 18136 31349 18152
rect 31349 18136 31398 18152
rect 31022 18121 31078 18136
rect 31102 18121 31158 18136
rect 31182 18121 31238 18136
rect 31262 18121 31318 18136
rect 31342 18121 31398 18136
rect 31022 18096 31029 18121
rect 31029 18096 31078 18121
rect 31022 18069 31029 18070
rect 31029 18069 31078 18070
rect 31102 18096 31145 18121
rect 31145 18096 31157 18121
rect 31157 18096 31158 18121
rect 31182 18096 31209 18121
rect 31209 18096 31221 18121
rect 31221 18096 31238 18121
rect 31262 18096 31273 18121
rect 31273 18096 31285 18121
rect 31285 18096 31318 18121
rect 31342 18096 31349 18121
rect 31349 18096 31398 18121
rect 31102 18069 31145 18070
rect 31145 18069 31157 18070
rect 31157 18069 31158 18070
rect 31182 18069 31209 18070
rect 31209 18069 31221 18070
rect 31221 18069 31238 18070
rect 31262 18069 31273 18070
rect 31273 18069 31285 18070
rect 31285 18069 31318 18070
rect 31342 18069 31349 18070
rect 31349 18069 31398 18070
rect 31022 18014 31078 18069
rect 31102 18014 31158 18069
rect 31182 18014 31238 18069
rect 31262 18014 31318 18069
rect 31342 18014 31398 18069
rect 31022 17932 31078 17988
rect 31102 17932 31158 17988
rect 31182 17932 31238 17988
rect 31262 17932 31318 17988
rect 31342 17932 31398 17988
rect 31022 17850 31078 17906
rect 31102 17850 31158 17906
rect 31182 17850 31238 17906
rect 31262 17850 31318 17906
rect 31342 17850 31398 17906
rect 31022 17768 31078 17824
rect 31102 17768 31158 17824
rect 31182 17768 31238 17824
rect 31262 17768 31318 17824
rect 31342 17768 31398 17824
rect 21641 8344 21697 8400
rect 21721 8344 21777 8400
rect 21801 8344 21857 8400
rect 21881 8344 21937 8400
rect 21641 8263 21697 8319
rect 21721 8263 21777 8319
rect 21801 8263 21857 8319
rect 21881 8263 21937 8319
rect 21641 8182 21697 8238
rect 21721 8182 21777 8238
rect 21801 8182 21857 8238
rect 21881 8182 21937 8238
rect 21641 8101 21697 8157
rect 21721 8101 21777 8157
rect 21801 8101 21857 8157
rect 21881 8101 21937 8157
rect 21641 8031 21686 8076
rect 21686 8031 21697 8076
rect 21721 8031 21753 8076
rect 21753 8031 21768 8076
rect 21768 8031 21777 8076
rect 21801 8031 21820 8076
rect 21820 8031 21834 8076
rect 21834 8031 21857 8076
rect 21881 8031 21886 8076
rect 21886 8031 21900 8076
rect 21900 8031 21937 8076
rect 21641 8020 21697 8031
rect 21721 8020 21777 8031
rect 21801 8020 21857 8031
rect 21881 8020 21937 8031
rect 21641 7967 21686 7995
rect 21686 7967 21697 7995
rect 21721 7967 21753 7995
rect 21753 7967 21768 7995
rect 21768 7967 21777 7995
rect 21801 7967 21820 7995
rect 21820 7967 21834 7995
rect 21834 7967 21857 7995
rect 21881 7967 21886 7995
rect 21886 7967 21900 7995
rect 21900 7967 21937 7995
rect 21641 7955 21697 7967
rect 21721 7955 21777 7967
rect 21801 7955 21857 7967
rect 21881 7955 21937 7967
rect 21641 7939 21686 7955
rect 21686 7939 21697 7955
rect 21721 7939 21753 7955
rect 21753 7939 21768 7955
rect 21768 7939 21777 7955
rect 21801 7939 21820 7955
rect 21820 7939 21834 7955
rect 21834 7939 21857 7955
rect 21881 7939 21886 7955
rect 21886 7939 21900 7955
rect 21900 7939 21937 7955
rect 21641 7903 21686 7914
rect 21686 7903 21697 7914
rect 21721 7903 21753 7914
rect 21753 7903 21768 7914
rect 21768 7903 21777 7914
rect 21801 7903 21820 7914
rect 21820 7903 21834 7914
rect 21834 7903 21857 7914
rect 21881 7903 21886 7914
rect 21886 7903 21900 7914
rect 21900 7903 21937 7914
rect 21641 7858 21697 7903
rect 21721 7858 21777 7903
rect 21801 7858 21857 7903
rect 21881 7858 21937 7903
rect 22231 8083 22287 8095
rect 22316 8083 22372 8095
rect 22400 8083 22456 8095
rect 22484 8083 22540 8095
rect 22568 8083 22624 8095
rect 22652 8083 22708 8095
rect 22231 8039 22239 8083
rect 22239 8039 22287 8083
rect 22316 8039 22361 8083
rect 22361 8039 22372 8083
rect 22400 8039 22431 8083
rect 22431 8039 22448 8083
rect 22448 8039 22456 8083
rect 22484 8039 22500 8083
rect 22500 8039 22517 8083
rect 22517 8039 22540 8083
rect 22568 8039 22569 8083
rect 22569 8039 22586 8083
rect 22586 8039 22624 8083
rect 22652 8039 22655 8083
rect 22655 8039 22707 8083
rect 22707 8039 22708 8083
rect 22231 7967 22239 8015
rect 22239 7967 22287 8015
rect 22316 7967 22361 8015
rect 22361 7967 22372 8015
rect 22400 7967 22431 8015
rect 22431 7967 22448 8015
rect 22448 7967 22456 8015
rect 22484 7967 22500 8015
rect 22500 7967 22517 8015
rect 22517 7967 22540 8015
rect 22568 7967 22569 8015
rect 22569 7967 22586 8015
rect 22586 7967 22624 8015
rect 22652 7967 22655 8015
rect 22655 7967 22707 8015
rect 22707 7967 22708 8015
rect 22231 7959 22287 7967
rect 22316 7959 22372 7967
rect 22400 7959 22456 7967
rect 22484 7959 22540 7967
rect 22568 7959 22624 7967
rect 22652 7959 22708 7967
rect 22231 7903 22239 7935
rect 22239 7903 22287 7935
rect 22316 7903 22361 7935
rect 22361 7903 22372 7935
rect 22400 7903 22431 7935
rect 22431 7903 22448 7935
rect 22448 7903 22456 7935
rect 22484 7903 22500 7935
rect 22500 7903 22517 7935
rect 22517 7903 22540 7935
rect 22568 7903 22569 7935
rect 22569 7903 22586 7935
rect 22586 7903 22624 7935
rect 22652 7903 22655 7935
rect 22655 7903 22707 7935
rect 22707 7903 22708 7935
rect 22231 7879 22287 7903
rect 22316 7879 22372 7903
rect 22400 7879 22456 7903
rect 22484 7879 22540 7903
rect 22568 7879 22624 7903
rect 22652 7879 22708 7903
rect 22090 3007 22146 3063
rect 22090 2927 22146 2983
rect 22090 2847 22146 2903
rect 22090 2767 22146 2823
rect 22090 2687 22146 2743
rect 22090 2607 22146 2663
rect 22090 2527 22146 2583
rect 22090 2447 22146 2503
rect 22090 2367 22146 2423
rect 22090 2287 22146 2343
rect 22090 2207 22146 2263
rect 22090 2127 22146 2183
rect 22090 2047 22146 2103
rect 22090 1967 22146 2023
rect 22090 1887 22146 1943
rect 22090 1807 22146 1863
rect 22090 1726 22146 1782
rect 22090 1645 22146 1701
rect 22090 1564 22146 1620
rect 22090 1483 22146 1539
rect 15246 -2937 15302 -2881
rect 15326 -2937 15382 -2881
rect 15406 -2937 15462 -2881
rect 15486 -2937 15542 -2881
rect 15566 -2937 15622 -2881
rect 15646 -2937 15702 -2881
rect 15726 -2937 15782 -2881
rect 15806 -2937 15862 -2881
rect 15886 -2937 15942 -2881
rect 15246 -3020 15302 -2964
rect 15326 -3020 15382 -2964
rect 15406 -3020 15462 -2964
rect 15486 -3020 15542 -2964
rect 15566 -3020 15622 -2964
rect 15646 -3020 15702 -2964
rect 15726 -3020 15782 -2964
rect 15806 -3020 15862 -2964
rect 15886 -3020 15942 -2964
rect 15246 -3103 15302 -3047
rect 15326 -3103 15382 -3047
rect 15406 -3103 15462 -3047
rect 15486 -3103 15542 -3047
rect 15566 -3103 15622 -3047
rect 15646 -3103 15702 -3047
rect 15726 -3103 15782 -3047
rect 15806 -3103 15862 -3047
rect 15886 -3103 15942 -3047
rect 15246 -3187 15302 -3131
rect 15326 -3187 15382 -3131
rect 15406 -3187 15462 -3131
rect 15486 -3187 15542 -3131
rect 15566 -3187 15622 -3131
rect 15646 -3187 15702 -3131
rect 15726 -3187 15782 -3131
rect 15806 -3187 15862 -3131
rect 15886 -3187 15942 -3131
rect 15246 -3271 15302 -3215
rect 15326 -3271 15382 -3215
rect 15406 -3271 15462 -3215
rect 15486 -3271 15542 -3215
rect 15566 -3271 15622 -3215
rect 15646 -3271 15702 -3215
rect 15726 -3271 15782 -3215
rect 15806 -3271 15862 -3215
rect 15886 -3271 15942 -3215
rect 15246 -3355 15302 -3299
rect 15326 -3355 15382 -3299
rect 15406 -3355 15462 -3299
rect 15486 -3355 15542 -3299
rect 15566 -3355 15622 -3299
rect 15646 -3355 15702 -3299
rect 15726 -3355 15782 -3299
rect 15806 -3355 15862 -3299
rect 15886 -3355 15942 -3299
rect 15246 -3439 15302 -3383
rect 15326 -3439 15382 -3383
rect 15406 -3439 15462 -3383
rect 15486 -3439 15542 -3383
rect 15566 -3439 15622 -3383
rect 15646 -3439 15702 -3383
rect 15726 -3439 15782 -3383
rect 15806 -3439 15862 -3383
rect 15886 -3439 15942 -3383
rect 15246 -3523 15302 -3467
rect 15326 -3523 15382 -3467
rect 15406 -3523 15462 -3467
rect 15486 -3523 15542 -3467
rect 15566 -3523 15622 -3467
rect 15646 -3523 15702 -3467
rect 15726 -3523 15782 -3467
rect 15806 -3523 15862 -3467
rect 15886 -3523 15942 -3467
rect 15246 -3607 15302 -3551
rect 15326 -3607 15382 -3551
rect 15406 -3607 15462 -3551
rect 15486 -3607 15542 -3551
rect 15566 -3607 15622 -3551
rect 15646 -3607 15702 -3551
rect 15726 -3607 15782 -3551
rect 15806 -3607 15862 -3551
rect 15886 -3607 15942 -3551
rect 15246 -3691 15302 -3635
rect 15326 -3691 15382 -3635
rect 15406 -3691 15462 -3635
rect 15486 -3691 15542 -3635
rect 15566 -3691 15622 -3635
rect 15646 -3691 15702 -3635
rect 15726 -3691 15782 -3635
rect 15806 -3691 15862 -3635
rect 15886 -3691 15942 -3635
rect 23450 2493 23586 3189
rect 23450 2412 23506 2468
rect 23530 2412 23586 2468
rect 23450 2331 23506 2387
rect 23530 2331 23586 2387
rect 23450 2250 23506 2306
rect 23530 2250 23586 2306
rect 23450 2169 23506 2225
rect 23530 2169 23586 2225
rect 23450 2088 23506 2144
rect 23530 2088 23586 2144
rect 23450 2007 23506 2063
rect 23530 2007 23586 2063
rect 23450 1926 23506 1982
rect 23530 1926 23586 1982
rect 23450 1845 23506 1901
rect 23530 1845 23586 1901
rect 23450 1764 23506 1820
rect 23530 1764 23586 1820
rect 23450 1683 23506 1739
rect 23530 1683 23586 1739
rect 23450 1602 23506 1658
rect 23530 1602 23586 1658
rect 23450 1521 23506 1577
rect 23530 1521 23586 1577
rect 23450 1440 23506 1496
rect 23530 1440 23586 1496
rect 23450 1359 23506 1415
rect 23530 1359 23586 1415
rect 24182 2734 24398 3190
rect 24182 2653 24238 2709
rect 24262 2653 24318 2709
rect 24342 2653 24398 2709
rect 24182 2572 24238 2628
rect 24262 2572 24318 2628
rect 24342 2572 24398 2628
rect 24182 2491 24238 2547
rect 24262 2491 24318 2547
rect 24342 2491 24398 2547
rect 24182 2410 24238 2466
rect 24262 2410 24318 2466
rect 24342 2410 24398 2466
rect 24182 2329 24238 2385
rect 24262 2329 24318 2385
rect 24342 2329 24398 2385
rect 24182 2248 24238 2304
rect 24262 2248 24318 2304
rect 24342 2248 24398 2304
rect 24182 2167 24238 2223
rect 24262 2167 24318 2223
rect 24342 2167 24398 2223
rect 24182 2086 24238 2142
rect 24262 2086 24318 2142
rect 24342 2086 24398 2142
rect 24182 2005 24238 2061
rect 24262 2005 24318 2061
rect 24342 2005 24398 2061
rect 24182 1924 24238 1980
rect 24262 1924 24318 1980
rect 24342 1924 24398 1980
rect 24182 1843 24238 1899
rect 24262 1843 24318 1899
rect 24342 1843 24398 1899
rect 24182 1762 24238 1818
rect 24262 1762 24318 1818
rect 24342 1762 24398 1818
rect 24182 1681 24238 1737
rect 24262 1681 24318 1737
rect 24342 1681 24398 1737
rect 24182 1600 24238 1656
rect 24262 1600 24318 1656
rect 24342 1600 24398 1656
rect 24182 1519 24238 1575
rect 24262 1519 24318 1575
rect 24342 1519 24398 1575
rect 24182 1438 24238 1494
rect 24262 1438 24318 1494
rect 24342 1438 24398 1494
rect 24182 1357 24238 1413
rect 24262 1357 24318 1413
rect 24342 1357 24398 1413
rect 23449 -2929 23505 -2873
rect 23529 -2929 23585 -2873
rect 23449 -3014 23505 -2958
rect 23529 -3014 23585 -2958
rect 23449 -3099 23505 -3043
rect 23529 -3099 23585 -3043
rect 23449 -3184 23505 -3128
rect 23529 -3184 23585 -3128
rect 23449 -3270 23505 -3214
rect 23529 -3270 23585 -3214
rect 23449 -3356 23505 -3300
rect 23529 -3356 23585 -3300
rect 23449 -3442 23505 -3386
rect 23529 -3442 23585 -3386
rect 23449 -3528 23505 -3472
rect 23529 -3528 23585 -3472
rect 23449 -3614 23505 -3558
rect 23529 -3614 23585 -3558
rect 23449 -3700 23505 -3644
rect 23529 -3700 23585 -3644
rect 24183 -2927 24239 -2871
rect 24263 -2927 24319 -2871
rect 24343 -2927 24399 -2871
rect 24183 -3013 24239 -2957
rect 24263 -3013 24319 -2957
rect 24343 -3013 24399 -2957
rect 27606 4623 27662 4679
rect 27686 4623 27742 4679
rect 27766 4623 27822 4679
rect 27846 4623 27902 4679
rect 27926 4623 27982 4679
rect 27606 4542 27662 4598
rect 27686 4542 27742 4598
rect 27766 4542 27822 4598
rect 27846 4542 27902 4598
rect 27926 4542 27982 4598
rect 27606 4461 27662 4517
rect 27686 4461 27742 4517
rect 27766 4461 27822 4517
rect 27846 4461 27902 4517
rect 27926 4461 27982 4517
rect 27606 4379 27662 4435
rect 27686 4379 27742 4435
rect 27766 4379 27822 4435
rect 27846 4379 27902 4435
rect 27926 4379 27982 4435
rect 27606 4297 27662 4353
rect 27686 4297 27742 4353
rect 27766 4297 27822 4353
rect 27846 4297 27902 4353
rect 27926 4297 27982 4353
rect 27606 4215 27662 4271
rect 27686 4215 27742 4271
rect 27766 4215 27822 4271
rect 27846 4215 27902 4271
rect 27926 4215 27982 4271
rect 27606 4133 27662 4189
rect 27686 4133 27742 4189
rect 27766 4133 27822 4189
rect 27846 4133 27902 4189
rect 27926 4133 27982 4189
rect 27606 4051 27662 4107
rect 27686 4051 27742 4107
rect 27766 4051 27822 4107
rect 27846 4051 27902 4107
rect 27926 4051 27982 4107
rect 27606 3969 27662 4025
rect 27686 3969 27742 4025
rect 27766 3969 27822 4025
rect 27846 3969 27902 4025
rect 27926 3969 27982 4025
rect 27606 3887 27662 3943
rect 27686 3887 27742 3943
rect 27766 3887 27822 3943
rect 27846 3887 27902 3943
rect 27926 3887 27982 3943
rect 27606 3805 27662 3861
rect 27686 3805 27742 3861
rect 27766 3805 27822 3861
rect 27846 3805 27902 3861
rect 27926 3805 27982 3861
rect 27606 3723 27662 3779
rect 27686 3723 27742 3779
rect 27766 3723 27822 3779
rect 27846 3723 27902 3779
rect 27926 3723 27982 3779
rect 25907 2380 25963 2436
rect 25987 2380 26043 2436
rect 26067 2380 26123 2436
rect 26147 2380 26203 2436
rect 26227 2380 26283 2436
rect 26307 2380 26363 2436
rect 25907 2297 25963 2353
rect 25987 2297 26043 2353
rect 26067 2297 26123 2353
rect 26147 2297 26203 2353
rect 26227 2297 26283 2353
rect 26307 2297 26363 2353
rect 25907 2214 25963 2270
rect 25987 2214 26043 2270
rect 26067 2214 26123 2270
rect 26147 2214 26203 2270
rect 26227 2214 26283 2270
rect 26307 2214 26363 2270
rect 25907 2131 25963 2187
rect 25987 2131 26043 2187
rect 26067 2131 26123 2187
rect 26147 2131 26203 2187
rect 26227 2131 26283 2187
rect 26307 2131 26363 2187
rect 25907 2048 25963 2104
rect 25987 2048 26043 2104
rect 26067 2048 26123 2104
rect 26147 2048 26203 2104
rect 26227 2048 26283 2104
rect 26307 2048 26363 2104
rect 25907 1965 25963 2021
rect 25987 1965 26043 2021
rect 26067 1965 26123 2021
rect 26147 1965 26203 2021
rect 26227 1965 26283 2021
rect 26307 1965 26363 2021
rect 25907 1882 25963 1938
rect 25987 1882 26043 1938
rect 26067 1882 26123 1938
rect 26147 1882 26203 1938
rect 26227 1882 26283 1938
rect 26307 1882 26363 1938
rect 25907 1799 25963 1855
rect 25987 1799 26043 1855
rect 26067 1799 26123 1855
rect 26147 1799 26203 1855
rect 26227 1799 26283 1855
rect 26307 1799 26363 1855
rect 25907 1715 25963 1771
rect 25987 1715 26043 1771
rect 26067 1715 26123 1771
rect 26147 1715 26203 1771
rect 26227 1715 26283 1771
rect 26307 1715 26363 1771
rect 25907 1631 25963 1687
rect 25987 1631 26043 1687
rect 26067 1631 26123 1687
rect 26147 1631 26203 1687
rect 26227 1631 26283 1687
rect 26307 1631 26363 1687
rect 25907 1547 25963 1603
rect 25987 1547 26043 1603
rect 26067 1547 26123 1603
rect 26147 1547 26203 1603
rect 26227 1547 26283 1603
rect 26307 1547 26363 1603
rect 25907 1463 25963 1519
rect 25987 1463 26043 1519
rect 26067 1463 26123 1519
rect 26147 1463 26203 1519
rect 26227 1463 26283 1519
rect 26307 1463 26363 1519
rect 25907 1379 25963 1435
rect 25987 1379 26043 1435
rect 26067 1379 26123 1435
rect 26147 1379 26203 1435
rect 26227 1379 26283 1435
rect 26307 1379 26363 1435
rect 27606 766 27662 822
rect 27686 766 27742 822
rect 27766 766 27822 822
rect 27846 766 27902 822
rect 27926 766 27982 822
rect 27606 685 27662 741
rect 27686 685 27742 741
rect 27766 685 27822 741
rect 27846 685 27902 741
rect 27926 685 27982 741
rect 27606 604 27662 660
rect 27686 604 27742 660
rect 27766 604 27822 660
rect 27846 604 27902 660
rect 27926 604 27982 660
rect 27606 523 27662 579
rect 27686 523 27742 579
rect 27766 523 27822 579
rect 27846 523 27902 579
rect 27926 523 27982 579
rect 27606 442 27662 498
rect 27686 442 27742 498
rect 27766 442 27822 498
rect 27846 442 27902 498
rect 27926 442 27982 498
rect 27606 361 27662 417
rect 27686 361 27742 417
rect 27766 361 27822 417
rect 27846 361 27902 417
rect 27926 361 27982 417
rect 27606 279 27662 335
rect 27686 279 27742 335
rect 27766 279 27822 335
rect 27846 279 27902 335
rect 27926 279 27982 335
rect 27606 197 27662 253
rect 27686 197 27742 253
rect 27766 197 27822 253
rect 27846 197 27902 253
rect 27926 197 27982 253
rect 27606 115 27662 171
rect 27686 115 27742 171
rect 27766 115 27822 171
rect 27846 115 27902 171
rect 27926 115 27982 171
rect 27606 33 27662 89
rect 27686 33 27742 89
rect 27766 33 27822 89
rect 27846 33 27902 89
rect 27926 33 27982 89
rect 27606 -49 27662 7
rect 27686 -49 27742 7
rect 27766 -49 27822 7
rect 27846 -49 27902 7
rect 27926 -49 27982 7
rect 27606 -131 27662 -75
rect 27686 -131 27742 -75
rect 27766 -131 27822 -75
rect 27846 -131 27902 -75
rect 27926 -131 27982 -75
rect 27606 -213 27662 -157
rect 27686 -213 27742 -157
rect 27766 -213 27822 -157
rect 27846 -213 27902 -157
rect 27926 -213 27982 -157
rect 27606 -295 27662 -239
rect 27686 -295 27742 -239
rect 27766 -295 27822 -239
rect 27846 -295 27902 -239
rect 27926 -295 27982 -239
rect 27606 -377 27662 -321
rect 27686 -377 27742 -321
rect 27766 -377 27822 -321
rect 27846 -377 27902 -321
rect 27926 -377 27982 -321
rect 25905 -2934 25961 -2878
rect 25985 -2934 26041 -2878
rect 26065 -2934 26121 -2878
rect 26145 -2934 26201 -2878
rect 26225 -2934 26281 -2878
rect 26305 -2934 26361 -2878
rect 24183 -3099 24239 -3043
rect 24263 -3099 24319 -3043
rect 24343 -3099 24399 -3043
rect 24183 -3185 24239 -3129
rect 24263 -3185 24319 -3129
rect 24343 -3185 24399 -3129
rect 24183 -3271 24239 -3215
rect 24263 -3271 24319 -3215
rect 24343 -3271 24399 -3215
rect 24183 -3357 24239 -3301
rect 24263 -3357 24319 -3301
rect 24343 -3357 24399 -3301
rect 24183 -3443 24239 -3387
rect 24263 -3443 24319 -3387
rect 24343 -3443 24399 -3387
rect 24183 -3529 24239 -3473
rect 24263 -3529 24319 -3473
rect 24343 -3529 24399 -3473
rect 24183 -3615 24239 -3559
rect 24263 -3615 24319 -3559
rect 24343 -3615 24399 -3559
rect 24183 -3702 24239 -3646
rect 24263 -3702 24319 -3646
rect 24343 -3702 24399 -3646
rect 25905 -3018 25961 -2962
rect 25985 -3018 26041 -2962
rect 26065 -3018 26121 -2962
rect 26145 -3018 26201 -2962
rect 26225 -3018 26281 -2962
rect 26305 -3018 26361 -2962
rect 25905 -3102 25961 -3046
rect 25985 -3102 26041 -3046
rect 26065 -3102 26121 -3046
rect 26145 -3102 26201 -3046
rect 26225 -3102 26281 -3046
rect 26305 -3102 26361 -3046
rect 25905 -3187 25961 -3131
rect 25985 -3187 26041 -3131
rect 26065 -3187 26121 -3131
rect 26145 -3187 26201 -3131
rect 26225 -3187 26281 -3131
rect 26305 -3187 26361 -3131
rect 25905 -3272 25961 -3216
rect 25985 -3272 26041 -3216
rect 26065 -3272 26121 -3216
rect 26145 -3272 26201 -3216
rect 26225 -3272 26281 -3216
rect 26305 -3272 26361 -3216
rect 25905 -3357 25961 -3301
rect 25985 -3357 26041 -3301
rect 26065 -3357 26121 -3301
rect 26145 -3357 26201 -3301
rect 26225 -3357 26281 -3301
rect 26305 -3357 26361 -3301
rect 25905 -3442 25961 -3386
rect 25985 -3442 26041 -3386
rect 26065 -3442 26121 -3386
rect 26145 -3442 26201 -3386
rect 26225 -3442 26281 -3386
rect 26305 -3442 26361 -3386
rect 25905 -3527 25961 -3471
rect 25985 -3527 26041 -3471
rect 26065 -3527 26121 -3471
rect 26145 -3527 26201 -3471
rect 26225 -3527 26281 -3471
rect 26305 -3527 26361 -3471
rect 25905 -3612 25961 -3556
rect 25985 -3612 26041 -3556
rect 26065 -3612 26121 -3556
rect 26145 -3612 26201 -3556
rect 26225 -3612 26281 -3556
rect 26305 -3612 26361 -3556
rect 25905 -3697 25961 -3641
rect 25985 -3697 26041 -3641
rect 26065 -3697 26121 -3641
rect 26145 -3697 26201 -3641
rect 26225 -3697 26281 -3641
rect 26305 -3697 26361 -3641
rect 21547 -4287 21603 -4231
rect 21627 -4287 21683 -4231
rect 21707 -4287 21763 -4231
rect 21787 -4287 21843 -4231
rect 21867 -4287 21923 -4231
rect 21947 -4287 22003 -4231
rect 22027 -4287 22083 -4231
rect 21547 -4377 21603 -4321
rect 21627 -4377 21683 -4321
rect 21707 -4377 21763 -4321
rect 21787 -4377 21843 -4321
rect 21867 -4377 21923 -4321
rect 21947 -4377 22003 -4321
rect 22027 -4377 22083 -4321
rect 21547 -4467 21603 -4411
rect 21627 -4467 21683 -4411
rect 21707 -4467 21763 -4411
rect 21787 -4467 21843 -4411
rect 21867 -4467 21923 -4411
rect 21947 -4467 22003 -4411
rect 22027 -4467 22083 -4411
rect 21547 -4558 21603 -4502
rect 21627 -4558 21683 -4502
rect 21707 -4558 21763 -4502
rect 21787 -4558 21843 -4502
rect 21867 -4558 21923 -4502
rect 21947 -4558 22003 -4502
rect 22027 -4558 22083 -4502
rect 21547 -4649 21603 -4593
rect 21627 -4649 21683 -4593
rect 21707 -4649 21763 -4593
rect 21787 -4649 21843 -4593
rect 21867 -4649 21923 -4593
rect 21947 -4649 22003 -4593
rect 22027 -4649 22083 -4593
rect 21547 -4740 21603 -4684
rect 21627 -4740 21683 -4684
rect 21707 -4740 21763 -4684
rect 21787 -4740 21843 -4684
rect 21867 -4740 21923 -4684
rect 21947 -4740 22003 -4684
rect 22027 -4740 22083 -4684
rect 21547 -4831 21603 -4775
rect 21627 -4831 21683 -4775
rect 21707 -4831 21763 -4775
rect 21787 -4831 21843 -4775
rect 21867 -4831 21923 -4775
rect 21947 -4831 22003 -4775
rect 22027 -4831 22083 -4775
rect 27606 -459 27662 -403
rect 27686 -459 27742 -403
rect 27766 -459 27822 -403
rect 27846 -459 27902 -403
rect 27926 -459 27982 -403
rect 28345 4629 28401 4685
rect 28425 4629 28481 4685
rect 28505 4629 28561 4685
rect 28585 4629 28641 4685
rect 28345 4547 28401 4603
rect 28425 4547 28481 4603
rect 28505 4547 28561 4603
rect 28585 4547 28641 4603
rect 28345 4465 28401 4521
rect 28425 4465 28481 4521
rect 28505 4465 28561 4521
rect 28585 4465 28641 4521
rect 28345 4383 28401 4439
rect 28425 4383 28481 4439
rect 28505 4383 28561 4439
rect 28585 4383 28641 4439
rect 28345 4301 28401 4357
rect 28425 4301 28481 4357
rect 28505 4301 28561 4357
rect 28585 4301 28641 4357
rect 28345 4219 28401 4275
rect 28425 4219 28481 4275
rect 28505 4219 28561 4275
rect 28585 4219 28641 4275
rect 28345 4137 28401 4193
rect 28425 4137 28481 4193
rect 28505 4137 28561 4193
rect 28585 4137 28641 4193
rect 28345 4055 28401 4111
rect 28425 4055 28481 4111
rect 28505 4055 28561 4111
rect 28585 4055 28641 4111
rect 28345 3972 28401 4028
rect 28425 3972 28481 4028
rect 28505 3972 28561 4028
rect 28585 3972 28641 4028
rect 28345 3889 28401 3945
rect 28425 3889 28481 3945
rect 28505 3889 28561 3945
rect 28585 3889 28641 3945
rect 28345 3806 28401 3862
rect 28425 3806 28481 3862
rect 28505 3806 28561 3862
rect 28585 3806 28641 3862
rect 28345 3723 28401 3779
rect 28425 3723 28481 3779
rect 28505 3723 28561 3779
rect 28585 3723 28641 3779
rect 28345 270 28641 806
rect 28345 189 28401 245
rect 28425 189 28481 245
rect 28505 189 28561 245
rect 28585 189 28641 245
rect 28345 108 28401 164
rect 28425 108 28481 164
rect 28505 108 28561 164
rect 28585 108 28641 164
rect 28345 27 28401 83
rect 28425 27 28481 83
rect 28505 27 28561 83
rect 28585 27 28641 83
rect 28345 -54 28401 2
rect 28425 -54 28481 2
rect 28505 -54 28561 2
rect 28585 -54 28641 2
rect 28345 -135 28401 -79
rect 28425 -135 28481 -79
rect 28505 -135 28561 -79
rect 28585 -135 28641 -79
rect 28345 -216 28401 -160
rect 28425 -216 28481 -160
rect 28505 -216 28561 -160
rect 28585 -216 28641 -160
rect 28345 -297 28401 -241
rect 28425 -297 28481 -241
rect 28505 -297 28561 -241
rect 28585 -297 28641 -241
rect 28345 -378 28401 -322
rect 28425 -378 28481 -322
rect 28505 -378 28561 -322
rect 28585 -378 28641 -322
rect 28345 -459 28401 -403
rect 28425 -459 28481 -403
rect 28505 -459 28561 -403
rect 28585 -459 28641 -403
<< metal3 >>
rect 19258 22257 19883 22262
rect 19258 22201 19263 22257
rect 19319 22201 19357 22257
rect 19413 22201 19450 22257
rect 19506 22201 19543 22257
rect 19599 22201 19636 22257
rect 19692 22201 19729 22257
rect 19785 22201 19822 22257
rect 19878 22201 19883 22257
rect 19258 22177 19883 22201
rect 19258 22121 19263 22177
rect 19319 22121 19357 22177
rect 19413 22121 19450 22177
rect 19506 22121 19543 22177
rect 19599 22121 19636 22177
rect 19692 22121 19729 22177
rect 19785 22121 19822 22177
rect 19878 22121 19883 22177
rect 19258 22116 19883 22121
rect 21006 22258 21870 22271
rect 21006 22202 21011 22258
rect 21067 22202 21100 22258
rect 21156 22202 21189 22258
rect 21245 22202 21278 22258
rect 21334 22202 21367 22258
rect 21423 22202 21456 22258
rect 21512 22202 21545 22258
rect 21601 22202 21633 22258
rect 21689 22202 21721 22258
rect 21777 22202 21809 22258
rect 21865 22202 21870 22258
rect 21006 22178 21870 22202
rect 21006 22122 21011 22178
rect 21067 22122 21100 22178
rect 21156 22122 21189 22178
rect 21245 22122 21278 22178
rect 21334 22122 21367 22178
rect 21423 22122 21456 22178
rect 21512 22122 21545 22178
rect 21601 22122 21633 22178
rect 21689 22122 21721 22178
rect 21777 22122 21809 22178
rect 21865 22122 21870 22178
rect 21006 22109 21870 22122
rect 14144 21085 14370 21561
rect 1135 19652 1354 19866
rect 19198 18807 31448 18818
rect 19198 18751 19217 18807
rect 19273 18751 19298 18807
rect 19354 18751 19379 18807
rect 19435 18751 19460 18807
rect 19516 18751 19541 18807
rect 19597 18751 19622 18807
rect 19678 18751 19703 18807
rect 19759 18751 19784 18807
rect 19840 18751 19865 18807
rect 19198 18727 19865 18751
rect 19198 18671 19217 18727
rect 19273 18671 19298 18727
rect 19354 18671 19379 18727
rect 19435 18671 19460 18727
rect 19516 18671 19541 18727
rect 19597 18671 19622 18727
rect 19678 18671 19703 18727
rect 19759 18671 19784 18727
rect 19840 18671 19865 18727
rect 19198 18647 19865 18671
rect 19198 18591 19217 18647
rect 19273 18591 19298 18647
rect 19354 18591 19379 18647
rect 19435 18591 19460 18647
rect 19516 18591 19541 18647
rect 19597 18591 19622 18647
rect 19678 18591 19703 18647
rect 19759 18591 19784 18647
rect 19840 18591 19865 18647
rect 19198 18567 19865 18591
rect 19198 18511 19217 18567
rect 19273 18511 19298 18567
rect 19354 18511 19379 18567
rect 19435 18511 19460 18567
rect 19516 18511 19541 18567
rect 19597 18511 19622 18567
rect 19678 18511 19703 18567
rect 19759 18511 19784 18567
rect 19840 18511 19865 18567
rect 20561 18751 21048 18807
rect 21104 18751 21136 18807
rect 21192 18751 21224 18807
rect 21280 18751 21311 18807
rect 21367 18751 21398 18807
rect 21454 18751 21485 18807
rect 21541 18751 21572 18807
rect 21628 18751 21659 18807
rect 21715 18804 31448 18807
rect 21715 18802 31022 18804
rect 21715 18751 24092 18802
rect 20561 18746 24092 18751
rect 24148 18746 24172 18802
rect 24228 18746 24252 18802
rect 24308 18791 31022 18802
rect 24308 18746 29488 18791
rect 20561 18735 29488 18746
rect 29544 18735 29568 18791
rect 29624 18735 29648 18791
rect 29704 18735 29728 18791
rect 29784 18748 31022 18791
rect 31078 18748 31102 18804
rect 31158 18748 31182 18804
rect 31238 18748 31262 18804
rect 31318 18748 31342 18804
rect 31398 18748 31448 18804
rect 29784 18735 31448 18748
rect 20561 18727 31448 18735
rect 20561 18671 21048 18727
rect 21104 18671 21136 18727
rect 21192 18671 21224 18727
rect 21280 18671 21311 18727
rect 21367 18671 21398 18727
rect 21454 18671 21485 18727
rect 21541 18671 21572 18727
rect 21628 18671 21659 18727
rect 21715 18723 31448 18727
rect 21715 18705 31022 18723
rect 21715 18689 29488 18705
rect 21715 18671 24092 18689
rect 20561 18647 24092 18671
rect 20561 18591 21048 18647
rect 21104 18591 21136 18647
rect 21192 18591 21224 18647
rect 21280 18591 21311 18647
rect 21367 18591 21398 18647
rect 21454 18591 21485 18647
rect 21541 18591 21572 18647
rect 21628 18591 21659 18647
rect 21715 18633 24092 18647
rect 24148 18633 24172 18689
rect 24228 18633 24252 18689
rect 24308 18649 29488 18689
rect 29544 18649 29568 18705
rect 29624 18649 29648 18705
rect 29704 18649 29728 18705
rect 29784 18667 31022 18705
rect 31078 18667 31102 18723
rect 31158 18667 31182 18723
rect 31238 18667 31262 18723
rect 31318 18667 31342 18723
rect 31398 18667 31448 18723
rect 29784 18649 31448 18667
rect 24308 18642 31448 18649
rect 24308 18633 31022 18642
rect 21715 18618 31022 18633
rect 21715 18591 29488 18618
rect 20561 18575 29488 18591
rect 20561 18567 24092 18575
rect 20561 18511 21048 18567
rect 21104 18511 21136 18567
rect 21192 18511 21224 18567
rect 21280 18511 21311 18567
rect 21367 18511 21398 18567
rect 21454 18511 21485 18567
rect 21541 18511 21572 18567
rect 21628 18511 21659 18567
rect 21715 18519 24092 18567
rect 24148 18519 24172 18575
rect 24228 18519 24252 18575
rect 24308 18562 29488 18575
rect 29544 18562 29568 18618
rect 29624 18562 29648 18618
rect 29704 18562 29728 18618
rect 29784 18586 31022 18618
rect 31078 18586 31102 18642
rect 31158 18586 31182 18642
rect 31238 18586 31262 18642
rect 31318 18586 31342 18642
rect 31398 18586 31448 18642
rect 29784 18562 31448 18586
rect 24308 18561 31448 18562
rect 24308 18531 31022 18561
rect 24308 18519 29488 18531
rect 21715 18511 29488 18519
rect 19198 18475 29488 18511
rect 29544 18475 29568 18531
rect 29624 18475 29648 18531
rect 29704 18475 29728 18531
rect 29784 18505 31022 18531
rect 31078 18505 31102 18561
rect 31158 18505 31182 18561
rect 31238 18505 31262 18561
rect 31318 18505 31342 18561
rect 31398 18505 31448 18561
rect 29784 18480 31448 18505
rect 29784 18475 31022 18480
rect 19198 18444 31022 18475
rect 19198 18388 29488 18444
rect 29544 18388 29568 18444
rect 29624 18388 29648 18444
rect 29704 18388 29728 18444
rect 29784 18424 31022 18444
rect 31078 18424 31102 18480
rect 31158 18424 31182 18480
rect 31238 18424 31262 18480
rect 31318 18424 31342 18480
rect 31398 18424 31448 18480
rect 29784 18398 31448 18424
rect 29784 18388 31022 18398
rect 19198 18357 31022 18388
rect 19198 18301 29488 18357
rect 29544 18301 29568 18357
rect 29624 18301 29648 18357
rect 29704 18301 29728 18357
rect 29784 18342 31022 18357
rect 31078 18342 31102 18398
rect 31158 18342 31182 18398
rect 31238 18342 31262 18398
rect 31318 18342 31342 18398
rect 31398 18342 31448 18398
rect 29784 18316 31448 18342
rect 29784 18301 31022 18316
rect 19198 18270 31022 18301
rect 19198 18214 29488 18270
rect 29544 18214 29568 18270
rect 29624 18214 29648 18270
rect 29704 18214 29728 18270
rect 29784 18260 31022 18270
rect 31078 18260 31102 18316
rect 31158 18260 31182 18316
rect 31238 18260 31262 18316
rect 31318 18260 31342 18316
rect 31398 18260 31448 18316
rect 29784 18234 31448 18260
rect 29784 18214 31022 18234
rect 19198 18183 31022 18214
rect 19198 18127 29488 18183
rect 29544 18127 29568 18183
rect 29624 18127 29648 18183
rect 29704 18127 29728 18183
rect 29784 18178 31022 18183
rect 31078 18178 31102 18234
rect 31158 18178 31182 18234
rect 31238 18178 31262 18234
rect 31318 18178 31342 18234
rect 31398 18178 31448 18234
rect 29784 18152 31448 18178
rect 29784 18127 31022 18152
rect 19198 18096 31022 18127
rect 31078 18096 31102 18152
rect 31158 18096 31182 18152
rect 31238 18096 31262 18152
rect 31318 18096 31342 18152
rect 31398 18096 31448 18152
rect 19198 18040 29488 18096
rect 29544 18040 29568 18096
rect 29624 18040 29648 18096
rect 29704 18040 29728 18096
rect 29784 18070 31448 18096
rect 29784 18040 31022 18070
rect 19198 18014 31022 18040
rect 31078 18014 31102 18070
rect 31158 18014 31182 18070
rect 31238 18014 31262 18070
rect 31318 18014 31342 18070
rect 31398 18014 31448 18070
rect 19198 18009 31448 18014
rect 19198 17953 29488 18009
rect 29544 17953 29568 18009
rect 29624 17953 29648 18009
rect 29704 17953 29728 18009
rect 29784 17988 31448 18009
rect 29784 17953 31022 17988
rect 19198 17932 31022 17953
rect 31078 17932 31102 17988
rect 31158 17932 31182 17988
rect 31238 17932 31262 17988
rect 31318 17932 31342 17988
rect 31398 17932 31448 17988
rect 19198 17922 31448 17932
rect 19198 17914 29488 17922
rect 19198 17858 26328 17914
rect 26384 17858 26416 17914
rect 26472 17858 26504 17914
rect 26560 17866 29488 17914
rect 29544 17866 29568 17922
rect 29624 17866 29648 17922
rect 29704 17866 29728 17922
rect 29784 17906 31448 17922
rect 29784 17866 31022 17906
rect 26560 17858 31022 17866
rect 19198 17850 31022 17858
rect 31078 17850 31102 17906
rect 31158 17850 31182 17906
rect 31238 17850 31262 17906
rect 31318 17850 31342 17906
rect 31398 17850 31448 17906
rect 19198 17835 31448 17850
rect 19198 17834 29488 17835
rect 19198 17778 26328 17834
rect 26384 17778 26416 17834
rect 26472 17778 26504 17834
rect 26560 17779 29488 17834
rect 29544 17779 29568 17835
rect 29624 17779 29648 17835
rect 29704 17779 29728 17835
rect 29784 17824 31448 17835
rect 29784 17779 31022 17824
rect 26560 17778 31022 17779
rect 19198 17768 31022 17778
rect 31078 17768 31102 17824
rect 31158 17768 31182 17824
rect 31238 17768 31262 17824
rect 31318 17768 31342 17824
rect 31398 17768 31448 17824
rect 19198 17750 31448 17768
rect 19174 14803 22779 14817
rect 19174 14775 20888 14803
rect 19174 14719 19471 14775
rect 19527 14719 19551 14775
rect 19607 14719 19631 14775
rect 19687 14719 19711 14775
rect 19767 14719 19791 14775
rect 19847 14719 20888 14775
rect 19174 14694 20888 14719
rect 19174 14638 19471 14694
rect 19527 14638 19551 14694
rect 19607 14638 19631 14694
rect 19687 14638 19711 14694
rect 19767 14638 19791 14694
rect 19847 14638 20888 14694
rect 19174 14613 20888 14638
rect 19174 14557 19471 14613
rect 19527 14557 19551 14613
rect 19607 14557 19631 14613
rect 19687 14557 19711 14613
rect 19767 14557 19791 14613
rect 19847 14557 20888 14613
rect 19174 14532 20888 14557
rect 19174 14476 19471 14532
rect 19527 14476 19551 14532
rect 19607 14476 19631 14532
rect 19687 14476 19711 14532
rect 19767 14476 19791 14532
rect 19847 14476 20888 14532
rect 19174 14451 20888 14476
rect 19174 14395 19471 14451
rect 19527 14395 19551 14451
rect 19607 14395 19631 14451
rect 19687 14395 19711 14451
rect 19767 14395 19791 14451
rect 19847 14395 20888 14451
rect 19174 14370 20888 14395
rect 19174 14314 19471 14370
rect 19527 14314 19551 14370
rect 19607 14314 19631 14370
rect 19687 14314 19711 14370
rect 19767 14314 19791 14370
rect 19847 14314 20888 14370
rect 19174 14289 20888 14314
rect 19174 14233 19471 14289
rect 19527 14233 19551 14289
rect 19607 14233 19631 14289
rect 19687 14233 19711 14289
rect 19767 14233 19791 14289
rect 19847 14233 20888 14289
rect 19174 14208 20888 14233
rect 19174 14152 19471 14208
rect 19527 14152 19551 14208
rect 19607 14152 19631 14208
rect 19687 14152 19711 14208
rect 19767 14152 19791 14208
rect 19847 14152 20888 14208
rect 19174 14127 20888 14152
rect 19174 14071 19471 14127
rect 19527 14071 19551 14127
rect 19607 14071 19631 14127
rect 19687 14071 19711 14127
rect 19767 14071 19791 14127
rect 19847 14071 20888 14127
rect 19174 14046 20888 14071
rect 19174 13990 19471 14046
rect 19527 13990 19551 14046
rect 19607 13990 19631 14046
rect 19687 13990 19711 14046
rect 19767 13990 19791 14046
rect 19847 13990 20888 14046
rect 19174 13965 20888 13990
rect 19174 13909 19471 13965
rect 19527 13909 19551 13965
rect 19607 13909 19631 13965
rect 19687 13909 19711 13965
rect 19767 13909 19791 13965
rect 19847 13909 20888 13965
rect 19174 13884 20888 13909
rect 19174 13828 19471 13884
rect 19527 13828 19551 13884
rect 19607 13828 19631 13884
rect 19687 13828 19711 13884
rect 19767 13828 19791 13884
rect 19847 13828 20888 13884
rect 19174 13803 20888 13828
rect 19174 13747 19471 13803
rect 19527 13747 19551 13803
rect 19607 13747 19631 13803
rect 19687 13747 19711 13803
rect 19767 13747 19791 13803
rect 19847 13747 20888 13803
rect 19174 13722 20888 13747
rect 19174 13666 19471 13722
rect 19527 13666 19551 13722
rect 19607 13666 19631 13722
rect 19687 13666 19711 13722
rect 19767 13666 19791 13722
rect 19847 13666 20888 13722
rect 19174 13641 20888 13666
rect 19174 13585 19471 13641
rect 19527 13585 19551 13641
rect 19607 13585 19631 13641
rect 19687 13585 19711 13641
rect 19767 13585 19791 13641
rect 19847 13585 20888 13641
rect 19174 13560 20888 13585
rect 19174 13504 19471 13560
rect 19527 13504 19551 13560
rect 19607 13504 19631 13560
rect 19687 13504 19711 13560
rect 19767 13504 19791 13560
rect 19847 13504 20888 13560
rect 19174 13479 20888 13504
rect 19174 13423 19471 13479
rect 19527 13423 19551 13479
rect 19607 13423 19631 13479
rect 19687 13423 19711 13479
rect 19767 13423 19791 13479
rect 19847 13423 20888 13479
rect 19174 13398 20888 13423
rect 19174 13342 19471 13398
rect 19527 13342 19551 13398
rect 19607 13342 19631 13398
rect 19687 13342 19711 13398
rect 19767 13342 19791 13398
rect 19847 13342 20888 13398
rect 19174 13317 20888 13342
rect 19174 13261 19471 13317
rect 19527 13261 19551 13317
rect 19607 13261 19631 13317
rect 19687 13261 19711 13317
rect 19767 13261 19791 13317
rect 19847 13307 20888 13317
rect 21104 14801 22779 14803
rect 21104 13307 21641 14801
rect 19847 13282 21641 13307
rect 19847 13261 20888 13282
rect 19174 13236 20888 13261
rect 19174 13180 19471 13236
rect 19527 13180 19551 13236
rect 19607 13180 19631 13236
rect 19687 13180 19711 13236
rect 19767 13180 19791 13236
rect 19847 13226 20888 13236
rect 20944 13226 20968 13282
rect 21024 13226 21048 13282
rect 21104 13226 21641 13282
rect 19847 13201 21641 13226
rect 19847 13180 20888 13201
rect 19174 13155 20888 13180
rect 19174 13099 19471 13155
rect 19527 13099 19551 13155
rect 19607 13099 19631 13155
rect 19687 13099 19711 13155
rect 19767 13099 19791 13155
rect 19847 13145 20888 13155
rect 20944 13145 20968 13201
rect 21024 13145 21048 13201
rect 21104 13145 21641 13201
rect 19847 13120 21641 13145
rect 19847 13099 20888 13120
rect 19174 13074 20888 13099
rect 19174 13018 19471 13074
rect 19527 13018 19551 13074
rect 19607 13018 19631 13074
rect 19687 13018 19711 13074
rect 19767 13018 19791 13074
rect 19847 13064 20888 13074
rect 20944 13064 20968 13120
rect 21024 13064 21048 13120
rect 21104 13064 21641 13120
rect 19847 13039 21641 13064
rect 19847 13018 20888 13039
rect 19174 12993 20888 13018
rect 19174 12937 19471 12993
rect 19527 12937 19551 12993
rect 19607 12937 19631 12993
rect 19687 12937 19711 12993
rect 19767 12937 19791 12993
rect 19847 12983 20888 12993
rect 20944 12983 20968 13039
rect 21024 12983 21048 13039
rect 21104 12983 21641 13039
rect 19847 12958 21641 12983
rect 19847 12937 20888 12958
rect 19174 12912 20888 12937
rect 19174 12856 19471 12912
rect 19527 12856 19551 12912
rect 19607 12856 19631 12912
rect 19687 12856 19711 12912
rect 19767 12856 19791 12912
rect 19847 12902 20888 12912
rect 20944 12902 20968 12958
rect 21024 12902 21048 12958
rect 21104 12902 21641 12958
rect 19847 12877 21641 12902
rect 19847 12856 20888 12877
rect 19174 12831 20888 12856
rect 19174 12775 19471 12831
rect 19527 12775 19551 12831
rect 19607 12775 19631 12831
rect 19687 12775 19711 12831
rect 19767 12775 19791 12831
rect 19847 12821 20888 12831
rect 20944 12821 20968 12877
rect 21024 12821 21048 12877
rect 21104 12821 21641 12877
rect 19847 12796 21641 12821
rect 19847 12775 20888 12796
rect 19174 12750 20888 12775
rect 19174 12694 19471 12750
rect 19527 12694 19551 12750
rect 19607 12694 19631 12750
rect 19687 12694 19711 12750
rect 19767 12694 19791 12750
rect 19847 12740 20888 12750
rect 20944 12740 20968 12796
rect 21024 12740 21048 12796
rect 21104 12740 21641 12796
rect 19847 12715 21641 12740
rect 19847 12694 20888 12715
rect 19174 12669 20888 12694
rect 19174 12613 19471 12669
rect 19527 12613 19551 12669
rect 19607 12613 19631 12669
rect 19687 12613 19711 12669
rect 19767 12613 19791 12669
rect 19847 12659 20888 12669
rect 20944 12659 20968 12715
rect 21024 12659 21048 12715
rect 21104 12659 21641 12715
rect 19847 12634 21641 12659
rect 19847 12613 20888 12634
rect 19174 12588 20888 12613
rect 19174 12532 19471 12588
rect 19527 12532 19551 12588
rect 19607 12532 19631 12588
rect 19687 12532 19711 12588
rect 19767 12532 19791 12588
rect 19847 12578 20888 12588
rect 20944 12578 20968 12634
rect 21024 12578 21048 12634
rect 21104 12578 21641 12634
rect 19847 12553 21641 12578
rect 19847 12532 20888 12553
rect 19174 12507 20888 12532
rect 19174 12451 19471 12507
rect 19527 12451 19551 12507
rect 19607 12451 19631 12507
rect 19687 12451 19711 12507
rect 19767 12451 19791 12507
rect 19847 12497 20888 12507
rect 20944 12497 20968 12553
rect 21024 12497 21048 12553
rect 21104 12497 21641 12553
rect 19847 12472 21641 12497
rect 19847 12451 20888 12472
rect 19174 12426 20888 12451
rect 19174 12370 19471 12426
rect 19527 12370 19551 12426
rect 19607 12370 19631 12426
rect 19687 12370 19711 12426
rect 19767 12370 19791 12426
rect 19847 12416 20888 12426
rect 20944 12416 20968 12472
rect 21024 12416 21048 12472
rect 21104 12416 21641 12472
rect 19847 12391 21641 12416
rect 19847 12370 20888 12391
rect 19174 12345 20888 12370
rect 19174 12289 19471 12345
rect 19527 12289 19551 12345
rect 19607 12289 19631 12345
rect 19687 12289 19711 12345
rect 19767 12289 19791 12345
rect 19847 12335 20888 12345
rect 20944 12335 20968 12391
rect 21024 12335 21048 12391
rect 21104 12335 21641 12391
rect 19847 12310 21641 12335
rect 19847 12289 20888 12310
rect 19174 12264 20888 12289
rect 19174 12208 19471 12264
rect 19527 12208 19551 12264
rect 19607 12208 19631 12264
rect 19687 12208 19711 12264
rect 19767 12208 19791 12264
rect 19847 12254 20888 12264
rect 20944 12254 20968 12310
rect 21024 12254 21048 12310
rect 21104 12254 21641 12310
rect 19847 12229 21641 12254
rect 19847 12208 20888 12229
rect 19174 12183 20888 12208
rect 19174 12127 19471 12183
rect 19527 12127 19551 12183
rect 19607 12127 19631 12183
rect 19687 12127 19711 12183
rect 19767 12127 19791 12183
rect 19847 12173 20888 12183
rect 20944 12173 20968 12229
rect 21024 12173 21048 12229
rect 21104 12173 21641 12229
rect 19847 12148 21641 12173
rect 19847 12127 20888 12148
rect 19174 12102 20888 12127
rect 19174 12046 19471 12102
rect 19527 12046 19551 12102
rect 19607 12046 19631 12102
rect 19687 12046 19711 12102
rect 19767 12046 19791 12102
rect 19847 12092 20888 12102
rect 20944 12092 20968 12148
rect 21024 12092 21048 12148
rect 21104 12092 21641 12148
rect 19847 12067 21641 12092
rect 19847 12046 20888 12067
rect 19174 12021 20888 12046
rect 19174 11965 19471 12021
rect 19527 11965 19551 12021
rect 19607 11965 19631 12021
rect 19687 11965 19711 12021
rect 19767 11965 19791 12021
rect 19847 12011 20888 12021
rect 20944 12011 20968 12067
rect 21024 12011 21048 12067
rect 21104 12011 21641 12067
rect 19847 11986 21641 12011
rect 19847 11965 20888 11986
rect 19174 11939 20888 11965
rect 19174 11883 19471 11939
rect 19527 11883 19551 11939
rect 19607 11883 19631 11939
rect 19687 11883 19711 11939
rect 19767 11883 19791 11939
rect 19847 11930 20888 11939
rect 20944 11930 20968 11986
rect 21024 11930 21048 11986
rect 21104 11930 21641 11986
rect 19847 11905 21641 11930
rect 19847 11883 20888 11905
rect 19174 11857 20888 11883
rect 19174 11801 19471 11857
rect 19527 11801 19551 11857
rect 19607 11801 19631 11857
rect 19687 11801 19711 11857
rect 19767 11801 19791 11857
rect 19847 11849 20888 11857
rect 20944 11849 20968 11905
rect 21024 11849 21048 11905
rect 21104 11849 21641 11905
rect 19847 11824 21641 11849
rect 19847 11801 20888 11824
rect 19174 11775 20888 11801
rect 19174 11719 19471 11775
rect 19527 11719 19551 11775
rect 19607 11719 19631 11775
rect 19687 11719 19711 11775
rect 19767 11719 19791 11775
rect 19847 11768 20888 11775
rect 20944 11768 20968 11824
rect 21024 11768 21048 11824
rect 21104 11768 21641 11824
rect 19847 11743 21641 11768
rect 19847 11719 20888 11743
rect 19174 11693 20888 11719
rect 19174 11637 19471 11693
rect 19527 11637 19551 11693
rect 19607 11637 19631 11693
rect 19687 11637 19711 11693
rect 19767 11637 19791 11693
rect 19847 11687 20888 11693
rect 20944 11687 20968 11743
rect 21024 11687 21048 11743
rect 21104 11687 21641 11743
rect 19847 11662 21641 11687
rect 19847 11637 20888 11662
rect 19174 11611 20888 11637
rect 19174 11555 19471 11611
rect 19527 11555 19551 11611
rect 19607 11555 19631 11611
rect 19687 11555 19711 11611
rect 19767 11555 19791 11611
rect 19847 11606 20888 11611
rect 20944 11606 20968 11662
rect 21024 11606 21048 11662
rect 21104 11606 21641 11662
rect 19847 11581 21641 11606
rect 19847 11555 20888 11581
rect 19174 11529 20888 11555
rect 19174 11473 19471 11529
rect 19527 11473 19551 11529
rect 19607 11473 19631 11529
rect 19687 11473 19711 11529
rect 19767 11473 19791 11529
rect 19847 11525 20888 11529
rect 20944 11525 20968 11581
rect 21024 11525 21048 11581
rect 21104 11525 21641 11581
rect 19847 11500 21641 11525
rect 19847 11473 20888 11500
rect 19174 11447 20888 11473
rect 19174 11391 19471 11447
rect 19527 11391 19551 11447
rect 19607 11391 19631 11447
rect 19687 11391 19711 11447
rect 19767 11391 19791 11447
rect 19847 11444 20888 11447
rect 20944 11444 20968 11500
rect 21024 11444 21048 11500
rect 21104 11444 21641 11500
rect 19847 11419 21641 11444
rect 19847 11391 20888 11419
rect 19174 11363 20888 11391
rect 20944 11363 20968 11419
rect 21024 11363 21048 11419
rect 21104 11363 21641 11419
rect 19174 11338 21641 11363
rect 19174 11336 20888 11338
rect 19174 11280 19462 11336
rect 19518 11333 20888 11336
rect 19518 11280 19720 11333
rect 19174 11277 19720 11280
rect 19776 11277 19800 11333
rect 19856 11282 20888 11333
rect 20944 11282 20968 11338
rect 21024 11282 21048 11338
rect 21104 11282 21641 11338
rect 19856 11277 21641 11282
rect 19174 11257 21641 11277
rect 19174 11256 20888 11257
rect 19174 11200 19462 11256
rect 19518 11252 20888 11256
rect 19518 11200 19720 11252
rect 19174 11196 19720 11200
rect 19776 11196 19800 11252
rect 19856 11201 20888 11252
rect 20944 11201 20968 11257
rect 21024 11201 21048 11257
rect 21104 11201 21641 11257
rect 19856 11196 21641 11201
rect 19174 11176 21641 11196
rect 19174 11120 19462 11176
rect 19518 11171 20888 11176
rect 19518 11120 19720 11171
rect 19174 11115 19720 11120
rect 19776 11115 19800 11171
rect 19856 11120 20888 11171
rect 20944 11120 20968 11176
rect 21024 11120 21048 11176
rect 21104 11120 21641 11176
rect 19856 11115 21641 11120
rect 19174 11096 21641 11115
rect 19174 11040 19462 11096
rect 19518 11095 21641 11096
rect 19518 11090 20888 11095
rect 19518 11040 19720 11090
rect 19174 11034 19720 11040
rect 19776 11034 19800 11090
rect 19856 11039 20888 11090
rect 20944 11039 20968 11095
rect 21024 11039 21048 11095
rect 21104 11039 21641 11095
rect 19856 11034 21641 11039
rect 19174 11015 21641 11034
rect 19174 10959 19462 11015
rect 19518 11014 21641 11015
rect 19518 11009 20888 11014
rect 19518 10959 19720 11009
rect 19174 10953 19720 10959
rect 19776 10953 19800 11009
rect 19856 10958 20888 11009
rect 20944 10958 20968 11014
rect 21024 10958 21048 11014
rect 21104 10958 21641 11014
rect 19856 10953 21641 10958
rect 19174 10934 21641 10953
rect 19174 10878 19462 10934
rect 19518 10933 21641 10934
rect 19518 10928 20888 10933
rect 19518 10878 19720 10928
rect 19174 10872 19720 10878
rect 19776 10872 19800 10928
rect 19856 10877 20888 10928
rect 20944 10877 20968 10933
rect 21024 10877 21048 10933
rect 21104 10877 21641 10933
rect 19856 10872 21641 10877
rect 19174 10853 21641 10872
rect 19174 10797 19462 10853
rect 19518 10852 21641 10853
rect 19518 10847 20888 10852
rect 19518 10797 19720 10847
rect 19174 10791 19720 10797
rect 19776 10791 19800 10847
rect 19856 10796 20888 10847
rect 20944 10796 20968 10852
rect 21024 10796 21048 10852
rect 21104 10796 21641 10852
rect 19856 10791 21641 10796
rect 19174 10772 21641 10791
rect 19174 10716 19462 10772
rect 19518 10771 21641 10772
rect 19518 10766 20888 10771
rect 19518 10716 19720 10766
rect 19174 10710 19720 10716
rect 19776 10710 19800 10766
rect 19856 10715 20888 10766
rect 20944 10715 20968 10771
rect 21024 10715 21048 10771
rect 21104 10715 21641 10771
rect 19856 10710 21641 10715
rect 19174 10691 21641 10710
rect 19174 10635 19462 10691
rect 19518 10690 21641 10691
rect 19518 10685 20888 10690
rect 19518 10635 19720 10685
rect 19174 10629 19720 10635
rect 19776 10629 19800 10685
rect 19856 10634 20888 10685
rect 20944 10634 20968 10690
rect 21024 10634 21048 10690
rect 21104 10634 21641 10690
rect 19856 10629 21641 10634
rect 19174 10610 21641 10629
rect 19174 10554 19462 10610
rect 19518 10609 21641 10610
rect 19518 10604 20888 10609
rect 19518 10554 19720 10604
rect 19174 10548 19720 10554
rect 19776 10548 19800 10604
rect 19856 10553 20888 10604
rect 20944 10553 20968 10609
rect 21024 10553 21048 10609
rect 21104 10553 21641 10609
rect 19856 10548 21641 10553
rect 19174 10529 21641 10548
rect 19174 10473 19462 10529
rect 19518 10528 21641 10529
rect 19518 10523 20888 10528
rect 19518 10473 19720 10523
rect 19174 10467 19720 10473
rect 19776 10467 19800 10523
rect 19856 10472 20888 10523
rect 20944 10472 20968 10528
rect 21024 10472 21048 10528
rect 21104 10472 21641 10528
rect 19856 10467 21641 10472
rect 19174 10448 21641 10467
rect 19174 10392 19462 10448
rect 19518 10447 21641 10448
rect 19518 10442 20888 10447
rect 19518 10392 19720 10442
rect 19174 10386 19720 10392
rect 19776 10386 19800 10442
rect 19856 10391 20888 10442
rect 20944 10391 20968 10447
rect 21024 10391 21048 10447
rect 21104 10391 21641 10447
rect 19856 10386 21641 10391
rect 19174 10367 21641 10386
rect 19174 10311 19462 10367
rect 19518 10366 21641 10367
rect 19518 10361 20888 10366
rect 19518 10311 19720 10361
rect 19174 10305 19720 10311
rect 19776 10305 19800 10361
rect 19856 10310 20888 10361
rect 20944 10310 20968 10366
rect 21024 10310 21048 10366
rect 21104 10310 21641 10366
rect 19856 10305 21641 10310
rect 19174 10286 21641 10305
rect 19174 10230 19462 10286
rect 19518 10285 21641 10286
rect 19518 10280 20888 10285
rect 19518 10230 19720 10280
rect 19174 10224 19720 10230
rect 19776 10224 19800 10280
rect 19856 10229 20888 10280
rect 20944 10229 20968 10285
rect 21024 10229 21048 10285
rect 21104 10229 21641 10285
rect 19856 10224 21641 10229
rect 19174 10205 21641 10224
rect 19174 10149 19462 10205
rect 19518 10204 21641 10205
rect 19518 10199 20888 10204
rect 19518 10149 19720 10199
rect 19174 10143 19720 10149
rect 19776 10143 19800 10199
rect 19856 10148 20888 10199
rect 20944 10148 20968 10204
rect 21024 10148 21048 10204
rect 21104 10148 21641 10204
rect 19856 10143 21641 10148
rect 19174 10124 21641 10143
rect 19174 10068 19462 10124
rect 19518 10123 21641 10124
rect 19518 10118 20888 10123
rect 19518 10068 19720 10118
rect 19174 10062 19720 10068
rect 19776 10062 19800 10118
rect 19856 10067 20888 10118
rect 20944 10067 20968 10123
rect 21024 10067 21048 10123
rect 21104 10067 21641 10123
rect 19856 10062 21641 10067
rect 19174 10043 21641 10062
rect 19174 9987 19462 10043
rect 19518 10042 21641 10043
rect 19518 10037 20888 10042
rect 19518 9987 19720 10037
rect 19174 9981 19720 9987
rect 19776 9981 19800 10037
rect 19856 9986 20888 10037
rect 20944 9986 20968 10042
rect 21024 9986 21048 10042
rect 21104 9986 21641 10042
rect 19856 9981 21641 9986
rect 19174 9962 21641 9981
rect 19174 9906 19462 9962
rect 19518 9961 21641 9962
rect 19518 9956 20888 9961
rect 19518 9906 19720 9956
rect 19174 9900 19720 9906
rect 19776 9900 19800 9956
rect 19856 9905 20888 9956
rect 20944 9905 20968 9961
rect 21024 9905 21048 9961
rect 21104 9905 21641 9961
rect 19856 9900 21641 9905
rect 19174 9881 21641 9900
rect 19174 9825 19462 9881
rect 19518 9880 21641 9881
rect 19518 9875 20888 9880
rect 19518 9825 19720 9875
rect 19174 9819 19720 9825
rect 19776 9819 19800 9875
rect 19856 9824 20888 9875
rect 20944 9824 20968 9880
rect 21024 9824 21048 9880
rect 21104 9824 21641 9880
rect 19856 9819 21641 9824
rect 19174 9800 21641 9819
rect 19174 9744 19462 9800
rect 19518 9799 21641 9800
rect 19518 9794 20888 9799
rect 19518 9744 19720 9794
rect 19174 9738 19720 9744
rect 19776 9738 19800 9794
rect 19856 9743 20888 9794
rect 20944 9743 20968 9799
rect 21024 9743 21048 9799
rect 21104 9743 21641 9799
rect 19856 9738 21641 9743
rect 19174 9719 21641 9738
rect 19174 9663 19462 9719
rect 19518 9718 21641 9719
rect 19518 9713 20888 9718
rect 19518 9663 19720 9713
rect 19174 9657 19720 9663
rect 19776 9657 19800 9713
rect 19856 9662 20888 9713
rect 20944 9662 20968 9718
rect 21024 9662 21048 9718
rect 21104 9662 21641 9718
rect 19856 9657 21641 9662
rect 19174 9638 21641 9657
rect 19174 9582 19462 9638
rect 19518 9637 21641 9638
rect 19518 9631 20888 9637
rect 19518 9582 19720 9631
rect 19174 9575 19720 9582
rect 19776 9575 19800 9631
rect 19856 9581 20888 9631
rect 20944 9581 20968 9637
rect 21024 9581 21048 9637
rect 21104 9581 21641 9637
rect 19856 9575 21641 9581
rect 19174 9557 21641 9575
rect 19174 9501 19462 9557
rect 19518 9556 21641 9557
rect 19518 9549 20888 9556
rect 19518 9501 19720 9549
rect 19174 9493 19720 9501
rect 19776 9493 19800 9549
rect 19856 9500 20888 9549
rect 20944 9500 20968 9556
rect 21024 9500 21048 9556
rect 21104 9500 21641 9556
rect 19856 9493 21641 9500
rect 19174 9476 21641 9493
rect 19174 9420 19462 9476
rect 19518 9475 21641 9476
rect 19518 9467 20888 9475
rect 19518 9420 19720 9467
rect 19174 9411 19720 9420
rect 19776 9411 19800 9467
rect 19856 9419 20888 9467
rect 20944 9419 20968 9475
rect 21024 9419 21048 9475
rect 21104 9419 21641 9475
rect 19856 9411 21641 9419
rect 19174 9395 21641 9411
rect 19174 9339 19462 9395
rect 19518 9394 21641 9395
rect 19518 9385 20888 9394
rect 19518 9339 19720 9385
rect 19174 9329 19720 9339
rect 19776 9329 19800 9385
rect 19856 9338 20888 9385
rect 20944 9338 20968 9394
rect 21024 9338 21048 9394
rect 21104 9338 21641 9394
rect 19856 9329 21641 9338
rect 19174 9314 21641 9329
rect 19174 9258 19462 9314
rect 19518 9313 21641 9314
rect 19518 9303 20888 9313
rect 19518 9258 19720 9303
rect 19174 9247 19720 9258
rect 19776 9247 19800 9303
rect 19856 9257 20888 9303
rect 20944 9257 20968 9313
rect 21024 9257 21048 9313
rect 21104 9257 21641 9313
rect 19856 9247 21641 9257
rect 19174 9233 21641 9247
rect 19174 9177 19462 9233
rect 19518 9232 21641 9233
rect 19518 9221 20888 9232
rect 19518 9177 19720 9221
rect 19174 9165 19720 9177
rect 19776 9165 19800 9221
rect 19856 9176 20888 9221
rect 20944 9176 20968 9232
rect 21024 9176 21048 9232
rect 21104 9176 21641 9232
rect 19856 9165 21641 9176
rect 19174 9152 21641 9165
rect 19174 9096 19462 9152
rect 19518 9151 21641 9152
rect 19518 9139 20888 9151
rect 19518 9096 19720 9139
rect 19174 9083 19720 9096
rect 19776 9083 19800 9139
rect 19856 9095 20888 9139
rect 20944 9095 20968 9151
rect 21024 9095 21048 9151
rect 21104 9095 21641 9151
rect 19856 9083 21641 9095
rect 19174 9071 21641 9083
rect 19174 9015 19462 9071
rect 19518 9070 21641 9071
rect 19518 9057 20888 9070
rect 19518 9015 19720 9057
rect 19174 9001 19720 9015
rect 19776 9001 19800 9057
rect 19856 9014 20888 9057
rect 20944 9014 20968 9070
rect 21024 9014 21048 9070
rect 21104 9014 21641 9070
rect 19856 9001 21641 9014
rect 19174 8990 21641 9001
rect 19174 8934 19462 8990
rect 19518 8989 21641 8990
rect 19518 8975 20888 8989
rect 19518 8934 19720 8975
rect 19174 8919 19720 8934
rect 19776 8919 19800 8975
rect 19856 8933 20888 8975
rect 20944 8933 20968 8989
rect 21024 8933 21048 8989
rect 21104 8933 21641 8989
rect 19856 8919 21641 8933
rect 19174 8909 21641 8919
rect 19174 8853 19462 8909
rect 19518 8908 21641 8909
rect 19518 8893 20888 8908
rect 19518 8853 19720 8893
rect 19174 8837 19720 8853
rect 19776 8837 19800 8893
rect 19856 8852 20888 8893
rect 20944 8852 20968 8908
rect 21024 8852 21048 8908
rect 21104 8852 21641 8908
rect 19856 8837 21641 8852
rect 19174 8828 21641 8837
rect 19174 8772 19462 8828
rect 19518 8827 21641 8828
rect 19518 8811 20888 8827
rect 19518 8772 19720 8811
rect 19174 8755 19720 8772
rect 19776 8755 19800 8811
rect 19856 8771 20888 8811
rect 20944 8771 20968 8827
rect 21024 8771 21048 8827
rect 21104 8771 21641 8827
rect 19856 8755 21641 8771
rect 19174 8746 21641 8755
rect 19174 8690 20888 8746
rect 20944 8690 20968 8746
rect 21024 8690 21048 8746
rect 21104 8690 21641 8746
rect 19174 8669 21641 8690
rect 19174 8613 19482 8669
rect 19538 8613 19562 8669
rect 19618 8613 19642 8669
rect 19698 8613 19722 8669
rect 19778 8613 19802 8669
rect 19858 8665 21641 8669
rect 19858 8613 20888 8665
rect 19174 8609 20888 8613
rect 20944 8609 20968 8665
rect 21024 8609 21048 8665
rect 21104 8609 21641 8665
rect 19174 8584 21641 8609
rect 19174 8528 19482 8584
rect 19538 8528 19562 8584
rect 19618 8528 19642 8584
rect 19698 8528 19722 8584
rect 19778 8528 19802 8584
rect 19858 8528 20888 8584
rect 20944 8528 20968 8584
rect 21024 8528 21048 8584
rect 21104 8528 21641 8584
rect 19174 8503 21641 8528
rect 19174 8498 20888 8503
rect 19174 8442 19482 8498
rect 19538 8442 19562 8498
rect 19618 8442 19642 8498
rect 19698 8442 19722 8498
rect 19778 8442 19802 8498
rect 19858 8447 20888 8498
rect 20944 8447 20968 8503
rect 21024 8447 21048 8503
rect 21104 8447 21641 8503
rect 19858 8442 21641 8447
rect 19174 8425 21641 8442
rect 21937 8425 22779 14801
rect 19174 8422 22779 8425
rect 19174 8412 20888 8422
rect 19174 8356 19482 8412
rect 19538 8356 19562 8412
rect 19618 8356 19642 8412
rect 19698 8356 19722 8412
rect 19778 8356 19802 8412
rect 19858 8366 20888 8412
rect 20944 8366 20968 8422
rect 21024 8366 21048 8422
rect 21104 8400 22779 8422
rect 21104 8366 21641 8400
rect 19858 8356 21641 8366
rect 19174 8344 21641 8356
rect 21697 8344 21721 8400
rect 21777 8344 21801 8400
rect 21857 8344 21881 8400
rect 21937 8344 22779 8400
rect 19174 8341 22779 8344
rect 19174 8326 20888 8341
rect 19174 8270 19482 8326
rect 19538 8270 19562 8326
rect 19618 8270 19642 8326
rect 19698 8270 19722 8326
rect 19778 8270 19802 8326
rect 19858 8285 20888 8326
rect 20944 8285 20968 8341
rect 21024 8285 21048 8341
rect 21104 8319 22779 8341
rect 21104 8285 21641 8319
rect 19858 8270 21641 8285
rect 19174 8263 21641 8270
rect 21697 8263 21721 8319
rect 21777 8263 21801 8319
rect 21857 8263 21881 8319
rect 21937 8263 22779 8319
rect 19174 8260 22779 8263
rect 19174 8240 20888 8260
rect 19174 8184 19482 8240
rect 19538 8184 19562 8240
rect 19618 8184 19642 8240
rect 19698 8184 19722 8240
rect 19778 8184 19802 8240
rect 19858 8204 20888 8240
rect 20944 8204 20968 8260
rect 21024 8204 21048 8260
rect 21104 8238 22779 8260
rect 21104 8204 21641 8238
rect 19858 8184 21641 8204
rect 19174 8182 21641 8184
rect 21697 8182 21721 8238
rect 21777 8182 21801 8238
rect 21857 8182 21881 8238
rect 21937 8182 22779 8238
rect 19174 8179 22779 8182
rect 19174 8154 20888 8179
rect 19174 8098 19482 8154
rect 19538 8098 19562 8154
rect 19618 8098 19642 8154
rect 19698 8098 19722 8154
rect 19778 8098 19802 8154
rect 19858 8123 20888 8154
rect 20944 8123 20968 8179
rect 21024 8123 21048 8179
rect 21104 8157 22779 8179
rect 21104 8123 21641 8157
rect 19858 8101 21641 8123
rect 21697 8101 21721 8157
rect 21777 8101 21801 8157
rect 21857 8101 21881 8157
rect 21937 8101 22779 8157
rect 19858 8098 22779 8101
rect 19174 8068 20888 8098
rect 19174 8012 19482 8068
rect 19538 8012 19562 8068
rect 19618 8012 19642 8068
rect 19698 8012 19722 8068
rect 19778 8012 19802 8068
rect 19858 8042 20888 8068
rect 20944 8042 20968 8098
rect 21024 8042 21048 8098
rect 21104 8095 22779 8098
rect 21104 8076 22231 8095
rect 21104 8042 21641 8076
rect 19858 8020 21641 8042
rect 21697 8020 21721 8076
rect 21777 8020 21801 8076
rect 21857 8020 21881 8076
rect 21937 8039 22231 8076
rect 22287 8039 22316 8095
rect 22372 8039 22400 8095
rect 22456 8039 22484 8095
rect 22540 8039 22568 8095
rect 22624 8039 22652 8095
rect 22708 8039 22779 8095
rect 21937 8020 22779 8039
rect 19858 8017 22779 8020
rect 19858 8012 20888 8017
rect 19174 7982 20888 8012
rect 19174 7926 19482 7982
rect 19538 7926 19562 7982
rect 19618 7926 19642 7982
rect 19698 7926 19722 7982
rect 19778 7926 19802 7982
rect 19858 7961 20888 7982
rect 20944 7961 20968 8017
rect 21024 7961 21048 8017
rect 21104 8015 22779 8017
rect 21104 7995 22231 8015
rect 21104 7961 21641 7995
rect 19858 7939 21641 7961
rect 21697 7939 21721 7995
rect 21777 7939 21801 7995
rect 21857 7939 21881 7995
rect 21937 7959 22231 7995
rect 22287 7959 22316 8015
rect 22372 7959 22400 8015
rect 22456 7959 22484 8015
rect 22540 7959 22568 8015
rect 22624 7959 22652 8015
rect 22708 7959 22779 8015
rect 21937 7939 22779 7959
rect 19858 7936 22779 7939
rect 19858 7926 20888 7936
rect 19174 7880 20888 7926
rect 20944 7880 20968 7936
rect 21024 7880 21048 7936
rect 21104 7935 22779 7936
rect 21104 7914 22231 7935
rect 21104 7880 21641 7914
rect 19174 7858 21641 7880
rect 21697 7858 21721 7914
rect 21777 7858 21801 7914
rect 21857 7858 21881 7914
rect 21937 7879 22231 7914
rect 22287 7879 22316 7935
rect 22372 7879 22400 7935
rect 22456 7879 22484 7935
rect 22540 7879 22568 7935
rect 22624 7879 22652 7935
rect 22708 7879 22779 7935
rect 21937 7858 22779 7879
rect 19174 7837 22779 7858
rect 167 5555 2016 7452
rect 3016 5558 15125 7452
rect -1959 5550 -1413 5555
rect -1959 5094 -1954 5550
rect -1418 5094 -1413 5550
rect -1959 5069 -1413 5094
rect -1959 5013 -1954 5069
rect -1898 5013 -1874 5069
rect -1818 5013 -1794 5069
rect -1738 5013 -1714 5069
rect -1658 5013 -1634 5069
rect -1578 5013 -1554 5069
rect -1498 5013 -1474 5069
rect -1418 5013 -1413 5069
rect -1959 4988 -1413 5013
rect -1959 4932 -1954 4988
rect -1898 4932 -1874 4988
rect -1818 4932 -1794 4988
rect -1738 4932 -1714 4988
rect -1658 4932 -1634 4988
rect -1578 4932 -1554 4988
rect -1498 4932 -1474 4988
rect -1418 4932 -1413 4988
rect -1959 4907 -1413 4932
rect -1959 4851 -1954 4907
rect -1898 4851 -1874 4907
rect -1818 4851 -1794 4907
rect -1738 4851 -1714 4907
rect -1658 4851 -1634 4907
rect -1578 4851 -1554 4907
rect -1498 4851 -1474 4907
rect -1418 4851 -1413 4907
rect -1959 4826 -1413 4851
rect -1959 4770 -1954 4826
rect -1898 4770 -1874 4826
rect -1818 4770 -1794 4826
rect -1738 4770 -1714 4826
rect -1658 4770 -1634 4826
rect -1578 4770 -1554 4826
rect -1498 4770 -1474 4826
rect -1418 4770 -1413 4826
rect -1959 4745 -1413 4770
rect -1959 4689 -1954 4745
rect -1898 4689 -1874 4745
rect -1818 4689 -1794 4745
rect -1738 4689 -1714 4745
rect -1658 4689 -1634 4745
rect -1578 4689 -1554 4745
rect -1498 4689 -1474 4745
rect -1418 4689 -1413 4745
rect -1959 4664 -1413 4689
rect -1959 4608 -1954 4664
rect -1898 4608 -1874 4664
rect -1818 4608 -1794 4664
rect -1738 4608 -1714 4664
rect -1658 4608 -1634 4664
rect -1578 4608 -1554 4664
rect -1498 4608 -1474 4664
rect -1418 4608 -1413 4664
rect -1959 4583 -1413 4608
rect -1959 4527 -1954 4583
rect -1898 4527 -1874 4583
rect -1818 4527 -1794 4583
rect -1738 4527 -1714 4583
rect -1658 4527 -1634 4583
rect -1578 4527 -1554 4583
rect -1498 4527 -1474 4583
rect -1418 4527 -1413 4583
rect -1959 4502 -1413 4527
rect -1959 4446 -1954 4502
rect -1898 4446 -1874 4502
rect -1818 4446 -1794 4502
rect -1738 4446 -1714 4502
rect -1658 4446 -1634 4502
rect -1578 4446 -1554 4502
rect -1498 4446 -1474 4502
rect -1418 4446 -1413 4502
rect -1959 4441 -1413 4446
rect -168 5550 2198 5555
rect -168 5094 -163 5550
rect 373 5094 1657 5550
rect 2193 5094 2198 5550
rect -168 5069 2198 5094
rect -168 5013 -163 5069
rect -107 5013 -83 5069
rect -27 5013 -3 5069
rect 53 5013 77 5069
rect 133 5013 157 5069
rect 213 5013 237 5069
rect 293 5013 317 5069
rect 373 5013 1657 5069
rect 1713 5013 1737 5069
rect 1793 5013 1817 5069
rect 1873 5013 1897 5069
rect 1953 5013 1977 5069
rect 2033 5013 2057 5069
rect 2113 5013 2137 5069
rect 2193 5013 2198 5069
rect -168 4988 2198 5013
rect -168 4932 -163 4988
rect -107 4932 -83 4988
rect -27 4932 -3 4988
rect 53 4932 77 4988
rect 133 4932 157 4988
rect 213 4932 237 4988
rect 293 4932 317 4988
rect 373 4932 1657 4988
rect 1713 4932 1737 4988
rect 1793 4932 1817 4988
rect 1873 4932 1897 4988
rect 1953 4932 1977 4988
rect 2033 4932 2057 4988
rect 2113 4932 2137 4988
rect 2193 4932 2198 4988
rect -168 4907 2198 4932
rect -168 4851 -163 4907
rect -107 4851 -83 4907
rect -27 4851 -3 4907
rect 53 4851 77 4907
rect 133 4851 157 4907
rect 213 4851 237 4907
rect 293 4851 317 4907
rect 373 4851 1657 4907
rect 1713 4851 1737 4907
rect 1793 4851 1817 4907
rect 1873 4851 1897 4907
rect 1953 4851 1977 4907
rect 2033 4851 2057 4907
rect 2113 4851 2137 4907
rect 2193 4851 2198 4907
rect -168 4826 2198 4851
rect -168 4770 -163 4826
rect -107 4770 -83 4826
rect -27 4770 -3 4826
rect 53 4770 77 4826
rect 133 4770 157 4826
rect 213 4770 237 4826
rect 293 4770 317 4826
rect 373 4770 1657 4826
rect 1713 4770 1737 4826
rect 1793 4770 1817 4826
rect 1873 4770 1897 4826
rect 1953 4770 1977 4826
rect 2033 4770 2057 4826
rect 2113 4770 2137 4826
rect 2193 4770 2198 4826
rect -168 4745 2198 4770
rect -168 4689 -163 4745
rect -107 4689 -83 4745
rect -27 4689 -3 4745
rect 53 4689 77 4745
rect 133 4689 157 4745
rect 213 4689 237 4745
rect 293 4689 317 4745
rect 373 4689 1657 4745
rect 1713 4689 1737 4745
rect 1793 4689 1817 4745
rect 1873 4689 1897 4745
rect 1953 4689 1977 4745
rect 2033 4689 2057 4745
rect 2113 4689 2137 4745
rect 2193 4689 2198 4745
rect -168 4664 2198 4689
rect -168 4608 -163 4664
rect -107 4608 -83 4664
rect -27 4608 -3 4664
rect 53 4608 77 4664
rect 133 4608 157 4664
rect 213 4608 237 4664
rect 293 4608 317 4664
rect 373 4608 1657 4664
rect 1713 4608 1737 4664
rect 1793 4608 1817 4664
rect 1873 4608 1897 4664
rect 1953 4608 1977 4664
rect 2033 4608 2057 4664
rect 2113 4608 2137 4664
rect 2193 4608 2198 4664
rect -168 4583 2198 4608
rect -168 4527 -163 4583
rect -107 4527 -83 4583
rect -27 4527 -3 4583
rect 53 4527 77 4583
rect 133 4527 157 4583
rect 213 4527 237 4583
rect 293 4527 317 4583
rect 373 4527 1657 4583
rect 1713 4527 1737 4583
rect 1793 4527 1817 4583
rect 1873 4527 1897 4583
rect 1953 4527 1977 4583
rect 2033 4527 2057 4583
rect 2113 4527 2137 4583
rect 2193 4527 2198 4583
rect -168 4502 2198 4527
rect -168 4446 -163 4502
rect -107 4446 -83 4502
rect -27 4446 -3 4502
rect 53 4446 77 4502
rect 133 4446 157 4502
rect 213 4446 237 4502
rect 293 4446 317 4502
rect 373 4446 1657 4502
rect 1713 4446 1737 4502
rect 1793 4446 1817 4502
rect 1873 4446 1897 4502
rect 1953 4446 1977 4502
rect 2033 4446 2057 4502
rect 2113 4446 2137 4502
rect 2193 4446 2198 4502
rect -168 4441 2198 4446
rect 3016 5550 10660 5558
rect 3016 5094 3458 5550
rect 3994 5094 5266 5550
rect 5802 5494 7061 5550
rect 7117 5494 7141 5550
rect 7197 5494 7221 5550
rect 7277 5494 7301 5550
rect 7357 5494 7381 5550
rect 7437 5494 7461 5550
rect 7517 5494 7541 5550
rect 7597 5530 10660 5550
rect 7597 5494 8872 5530
rect 5802 5474 8872 5494
rect 8928 5474 8952 5530
rect 9008 5474 9032 5530
rect 9088 5474 9112 5530
rect 9168 5474 9192 5530
rect 9248 5474 9272 5530
rect 9328 5474 9352 5530
rect 9408 5502 10660 5530
rect 10716 5502 10740 5558
rect 10796 5502 10820 5558
rect 10876 5502 10900 5558
rect 10956 5502 10980 5558
rect 11036 5502 11060 5558
rect 11116 5502 11140 5558
rect 11196 5502 12465 5558
rect 12521 5502 12545 5558
rect 12601 5502 12625 5558
rect 12681 5502 12705 5558
rect 12761 5502 12785 5558
rect 12841 5502 12865 5558
rect 12921 5502 12945 5558
rect 13001 5502 14278 5558
rect 14334 5502 14358 5558
rect 14414 5502 14438 5558
rect 14494 5502 14518 5558
rect 14574 5502 14598 5558
rect 14654 5502 14678 5558
rect 14734 5502 14758 5558
rect 14814 5502 15125 5558
rect 9408 5476 15125 5502
rect 9408 5474 10660 5476
rect 5802 5467 10660 5474
rect 5802 5411 7061 5467
rect 7117 5411 7141 5467
rect 7197 5411 7221 5467
rect 7277 5411 7301 5467
rect 7357 5411 7381 5467
rect 7437 5411 7461 5467
rect 7517 5411 7541 5467
rect 7597 5449 10660 5467
rect 7597 5411 8872 5449
rect 5802 5393 8872 5411
rect 8928 5393 8952 5449
rect 9008 5393 9032 5449
rect 9088 5393 9112 5449
rect 9168 5393 9192 5449
rect 9248 5393 9272 5449
rect 9328 5393 9352 5449
rect 9408 5420 10660 5449
rect 10716 5420 10740 5476
rect 10796 5420 10820 5476
rect 10876 5420 10900 5476
rect 10956 5420 10980 5476
rect 11036 5420 11060 5476
rect 11116 5420 11140 5476
rect 11196 5420 12465 5476
rect 12521 5420 12545 5476
rect 12601 5420 12625 5476
rect 12681 5420 12705 5476
rect 12761 5420 12785 5476
rect 12841 5420 12865 5476
rect 12921 5420 12945 5476
rect 13001 5420 14278 5476
rect 14334 5420 14358 5476
rect 14414 5420 14438 5476
rect 14494 5420 14518 5476
rect 14574 5420 14598 5476
rect 14654 5420 14678 5476
rect 14734 5420 14758 5476
rect 14814 5420 15125 5476
rect 9408 5393 15125 5420
rect 5802 5384 10660 5393
rect 5802 5328 7061 5384
rect 7117 5328 7141 5384
rect 7197 5328 7221 5384
rect 7277 5328 7301 5384
rect 7357 5328 7381 5384
rect 7437 5328 7461 5384
rect 7517 5328 7541 5384
rect 7597 5368 10660 5384
rect 7597 5328 8872 5368
rect 5802 5312 8872 5328
rect 8928 5312 8952 5368
rect 9008 5312 9032 5368
rect 9088 5312 9112 5368
rect 9168 5312 9192 5368
rect 9248 5312 9272 5368
rect 9328 5312 9352 5368
rect 9408 5337 10660 5368
rect 10716 5337 10740 5393
rect 10796 5337 10820 5393
rect 10876 5337 10900 5393
rect 10956 5337 10980 5393
rect 11036 5337 11060 5393
rect 11116 5337 11140 5393
rect 11196 5337 12465 5393
rect 12521 5337 12545 5393
rect 12601 5337 12625 5393
rect 12681 5337 12705 5393
rect 12761 5337 12785 5393
rect 12841 5337 12865 5393
rect 12921 5337 12945 5393
rect 13001 5337 14278 5393
rect 14334 5337 14358 5393
rect 14414 5337 14438 5393
rect 14494 5337 14518 5393
rect 14574 5337 14598 5393
rect 14654 5337 14678 5393
rect 14734 5337 14758 5393
rect 14814 5337 15125 5393
rect 9408 5312 15125 5337
rect 5802 5310 15125 5312
rect 5802 5301 10660 5310
rect 5802 5245 7061 5301
rect 7117 5245 7141 5301
rect 7197 5245 7221 5301
rect 7277 5245 7301 5301
rect 7357 5245 7381 5301
rect 7437 5245 7461 5301
rect 7517 5245 7541 5301
rect 7597 5287 10660 5301
rect 7597 5245 8872 5287
rect 5802 5231 8872 5245
rect 8928 5231 8952 5287
rect 9008 5231 9032 5287
rect 9088 5231 9112 5287
rect 9168 5231 9192 5287
rect 9248 5231 9272 5287
rect 9328 5231 9352 5287
rect 9408 5254 10660 5287
rect 10716 5254 10740 5310
rect 10796 5254 10820 5310
rect 10876 5254 10900 5310
rect 10956 5254 10980 5310
rect 11036 5254 11060 5310
rect 11116 5254 11140 5310
rect 11196 5254 12465 5310
rect 12521 5254 12545 5310
rect 12601 5254 12625 5310
rect 12681 5254 12705 5310
rect 12761 5254 12785 5310
rect 12841 5254 12865 5310
rect 12921 5254 12945 5310
rect 13001 5254 14278 5310
rect 14334 5254 14358 5310
rect 14414 5254 14438 5310
rect 14494 5254 14518 5310
rect 14574 5254 14598 5310
rect 14654 5254 14678 5310
rect 14734 5254 14758 5310
rect 14814 5254 15125 5310
rect 9408 5231 15125 5254
rect 5802 5227 15125 5231
rect 5802 5218 10660 5227
rect 5802 5162 7061 5218
rect 7117 5162 7141 5218
rect 7197 5162 7221 5218
rect 7277 5162 7301 5218
rect 7357 5162 7381 5218
rect 7437 5162 7461 5218
rect 7517 5162 7541 5218
rect 7597 5206 10660 5218
rect 7597 5162 8872 5206
rect 5802 5150 8872 5162
rect 8928 5150 8952 5206
rect 9008 5150 9032 5206
rect 9088 5150 9112 5206
rect 9168 5150 9192 5206
rect 9248 5150 9272 5206
rect 9328 5150 9352 5206
rect 9408 5171 10660 5206
rect 10716 5171 10740 5227
rect 10796 5171 10820 5227
rect 10876 5171 10900 5227
rect 10956 5171 10980 5227
rect 11036 5171 11060 5227
rect 11116 5171 11140 5227
rect 11196 5171 12465 5227
rect 12521 5171 12545 5227
rect 12601 5171 12625 5227
rect 12681 5171 12705 5227
rect 12761 5171 12785 5227
rect 12841 5171 12865 5227
rect 12921 5171 12945 5227
rect 13001 5171 14278 5227
rect 14334 5171 14358 5227
rect 14414 5171 14438 5227
rect 14494 5171 14518 5227
rect 14574 5171 14598 5227
rect 14654 5171 14678 5227
rect 14734 5171 14758 5227
rect 14814 5171 15125 5227
rect 9408 5150 15125 5171
rect 5802 5144 15125 5150
rect 5802 5134 10660 5144
rect 5802 5094 7061 5134
rect 3016 5078 7061 5094
rect 7117 5078 7141 5134
rect 7197 5078 7221 5134
rect 7277 5078 7301 5134
rect 7357 5078 7381 5134
rect 7437 5078 7461 5134
rect 7517 5078 7541 5134
rect 7597 5125 10660 5134
rect 7597 5078 8872 5125
rect 3016 5069 8872 5078
rect 8928 5069 8952 5125
rect 9008 5069 9032 5125
rect 9088 5069 9112 5125
rect 9168 5069 9192 5125
rect 9248 5069 9272 5125
rect 9328 5069 9352 5125
rect 9408 5088 10660 5125
rect 10716 5088 10740 5144
rect 10796 5088 10820 5144
rect 10876 5088 10900 5144
rect 10956 5088 10980 5144
rect 11036 5088 11060 5144
rect 11116 5088 11140 5144
rect 11196 5088 12465 5144
rect 12521 5088 12545 5144
rect 12601 5088 12625 5144
rect 12681 5088 12705 5144
rect 12761 5088 12785 5144
rect 12841 5088 12865 5144
rect 12921 5088 12945 5144
rect 13001 5088 14278 5144
rect 14334 5088 14358 5144
rect 14414 5088 14438 5144
rect 14494 5088 14518 5144
rect 14574 5088 14598 5144
rect 14654 5088 14678 5144
rect 14734 5088 14758 5144
rect 14814 5088 15125 5144
rect 9408 5069 15125 5088
rect 3016 5013 3458 5069
rect 3514 5013 3538 5069
rect 3594 5013 3618 5069
rect 3674 5013 3698 5069
rect 3754 5013 3778 5069
rect 3834 5013 3858 5069
rect 3914 5013 3938 5069
rect 3994 5013 5266 5069
rect 5322 5013 5346 5069
rect 5402 5013 5426 5069
rect 5482 5013 5506 5069
rect 5562 5013 5586 5069
rect 5642 5013 5666 5069
rect 5722 5013 5746 5069
rect 5802 5061 15125 5069
rect 5802 5050 10660 5061
rect 5802 5013 7061 5050
rect 3016 4994 7061 5013
rect 7117 4994 7141 5050
rect 7197 4994 7221 5050
rect 7277 4994 7301 5050
rect 7357 4994 7381 5050
rect 7437 4994 7461 5050
rect 7517 4994 7541 5050
rect 7597 5044 10660 5050
rect 7597 4994 8872 5044
rect 3016 4988 8872 4994
rect 8928 4988 8952 5044
rect 9008 4988 9032 5044
rect 9088 4988 9112 5044
rect 9168 4988 9192 5044
rect 9248 4988 9272 5044
rect 9328 4988 9352 5044
rect 9408 5005 10660 5044
rect 10716 5005 10740 5061
rect 10796 5005 10820 5061
rect 10876 5005 10900 5061
rect 10956 5005 10980 5061
rect 11036 5005 11060 5061
rect 11116 5005 11140 5061
rect 11196 5005 12465 5061
rect 12521 5005 12545 5061
rect 12601 5005 12625 5061
rect 12681 5005 12705 5061
rect 12761 5005 12785 5061
rect 12841 5005 12865 5061
rect 12921 5005 12945 5061
rect 13001 5005 14278 5061
rect 14334 5005 14358 5061
rect 14414 5005 14438 5061
rect 14494 5005 14518 5061
rect 14574 5005 14598 5061
rect 14654 5005 14678 5061
rect 14734 5005 14758 5061
rect 14814 5005 15125 5061
rect 9408 4988 15125 5005
rect 3016 4932 3458 4988
rect 3514 4932 3538 4988
rect 3594 4932 3618 4988
rect 3674 4932 3698 4988
rect 3754 4932 3778 4988
rect 3834 4932 3858 4988
rect 3914 4932 3938 4988
rect 3994 4932 5266 4988
rect 5322 4932 5346 4988
rect 5402 4932 5426 4988
rect 5482 4932 5506 4988
rect 5562 4932 5586 4988
rect 5642 4932 5666 4988
rect 5722 4932 5746 4988
rect 5802 4978 15125 4988
rect 5802 4966 10660 4978
rect 5802 4932 7061 4966
rect 3016 4910 7061 4932
rect 7117 4910 7141 4966
rect 7197 4910 7221 4966
rect 7277 4910 7301 4966
rect 7357 4910 7381 4966
rect 7437 4910 7461 4966
rect 7517 4910 7541 4966
rect 7597 4963 10660 4966
rect 7597 4910 8872 4963
rect 3016 4907 8872 4910
rect 8928 4907 8952 4963
rect 9008 4907 9032 4963
rect 9088 4907 9112 4963
rect 9168 4907 9192 4963
rect 9248 4907 9272 4963
rect 9328 4907 9352 4963
rect 9408 4922 10660 4963
rect 10716 4922 10740 4978
rect 10796 4922 10820 4978
rect 10876 4922 10900 4978
rect 10956 4922 10980 4978
rect 11036 4922 11060 4978
rect 11116 4922 11140 4978
rect 11196 4922 12465 4978
rect 12521 4922 12545 4978
rect 12601 4922 12625 4978
rect 12681 4922 12705 4978
rect 12761 4922 12785 4978
rect 12841 4922 12865 4978
rect 12921 4922 12945 4978
rect 13001 4922 14278 4978
rect 14334 4922 14358 4978
rect 14414 4922 14438 4978
rect 14494 4922 14518 4978
rect 14574 4922 14598 4978
rect 14654 4922 14678 4978
rect 14734 4922 14758 4978
rect 14814 4922 15125 4978
rect 9408 4907 15125 4922
rect 3016 4851 3458 4907
rect 3514 4851 3538 4907
rect 3594 4851 3618 4907
rect 3674 4851 3698 4907
rect 3754 4851 3778 4907
rect 3834 4851 3858 4907
rect 3914 4851 3938 4907
rect 3994 4851 5266 4907
rect 5322 4851 5346 4907
rect 5402 4851 5426 4907
rect 5482 4851 5506 4907
rect 5562 4851 5586 4907
rect 5642 4851 5666 4907
rect 5722 4851 5746 4907
rect 5802 4895 15125 4907
rect 5802 4882 10660 4895
rect 5802 4851 7061 4882
rect 3016 4826 7061 4851
rect 7117 4826 7141 4882
rect 7197 4826 7221 4882
rect 7277 4826 7301 4882
rect 7357 4826 7381 4882
rect 7437 4826 7461 4882
rect 7517 4826 7541 4882
rect 7597 4881 10660 4882
rect 7597 4826 8872 4881
rect 3016 4770 3458 4826
rect 3514 4770 3538 4826
rect 3594 4770 3618 4826
rect 3674 4770 3698 4826
rect 3754 4770 3778 4826
rect 3834 4770 3858 4826
rect 3914 4770 3938 4826
rect 3994 4770 5266 4826
rect 5322 4770 5346 4826
rect 5402 4770 5426 4826
rect 5482 4770 5506 4826
rect 5562 4770 5586 4826
rect 5642 4770 5666 4826
rect 5722 4770 5746 4826
rect 5802 4825 8872 4826
rect 8928 4825 8952 4881
rect 9008 4825 9032 4881
rect 9088 4825 9112 4881
rect 9168 4825 9192 4881
rect 9248 4825 9272 4881
rect 9328 4825 9352 4881
rect 9408 4839 10660 4881
rect 10716 4839 10740 4895
rect 10796 4839 10820 4895
rect 10876 4839 10900 4895
rect 10956 4839 10980 4895
rect 11036 4839 11060 4895
rect 11116 4839 11140 4895
rect 11196 4839 12465 4895
rect 12521 4839 12545 4895
rect 12601 4839 12625 4895
rect 12681 4839 12705 4895
rect 12761 4839 12785 4895
rect 12841 4839 12865 4895
rect 12921 4839 12945 4895
rect 13001 4839 14278 4895
rect 14334 4839 14358 4895
rect 14414 4839 14438 4895
rect 14494 4839 14518 4895
rect 14574 4839 14598 4895
rect 14654 4839 14678 4895
rect 14734 4839 14758 4895
rect 14814 4839 15125 4895
rect 9408 4825 15125 4839
rect 5802 4812 15125 4825
rect 5802 4799 10660 4812
rect 5802 4798 8872 4799
rect 5802 4770 7061 4798
rect 3016 4745 7061 4770
rect 3016 4689 3458 4745
rect 3514 4689 3538 4745
rect 3594 4689 3618 4745
rect 3674 4689 3698 4745
rect 3754 4689 3778 4745
rect 3834 4689 3858 4745
rect 3914 4689 3938 4745
rect 3994 4689 5266 4745
rect 5322 4689 5346 4745
rect 5402 4689 5426 4745
rect 5482 4689 5506 4745
rect 5562 4689 5586 4745
rect 5642 4689 5666 4745
rect 5722 4689 5746 4745
rect 5802 4742 7061 4745
rect 7117 4742 7141 4798
rect 7197 4742 7221 4798
rect 7277 4742 7301 4798
rect 7357 4742 7381 4798
rect 7437 4742 7461 4798
rect 7517 4742 7541 4798
rect 7597 4743 8872 4798
rect 8928 4743 8952 4799
rect 9008 4743 9032 4799
rect 9088 4743 9112 4799
rect 9168 4743 9192 4799
rect 9248 4743 9272 4799
rect 9328 4743 9352 4799
rect 9408 4756 10660 4799
rect 10716 4756 10740 4812
rect 10796 4756 10820 4812
rect 10876 4756 10900 4812
rect 10956 4756 10980 4812
rect 11036 4756 11060 4812
rect 11116 4756 11140 4812
rect 11196 4756 12465 4812
rect 12521 4756 12545 4812
rect 12601 4756 12625 4812
rect 12681 4756 12705 4812
rect 12761 4756 12785 4812
rect 12841 4756 12865 4812
rect 12921 4756 12945 4812
rect 13001 4756 14278 4812
rect 14334 4756 14358 4812
rect 14414 4756 14438 4812
rect 14494 4756 14518 4812
rect 14574 4756 14598 4812
rect 14654 4756 14678 4812
rect 14734 4756 14758 4812
rect 14814 4756 15125 4812
rect 9408 4743 15125 4756
rect 7597 4742 15125 4743
rect 5802 4729 15125 4742
rect 5802 4717 10660 4729
rect 5802 4689 8872 4717
rect 3016 4664 8872 4689
rect 3016 4608 3458 4664
rect 3514 4608 3538 4664
rect 3594 4608 3618 4664
rect 3674 4608 3698 4664
rect 3754 4608 3778 4664
rect 3834 4608 3858 4664
rect 3914 4608 3938 4664
rect 3994 4608 5266 4664
rect 5322 4608 5346 4664
rect 5402 4608 5426 4664
rect 5482 4608 5506 4664
rect 5562 4608 5586 4664
rect 5642 4608 5666 4664
rect 5722 4608 5746 4664
rect 5802 4661 8872 4664
rect 8928 4661 8952 4717
rect 9008 4661 9032 4717
rect 9088 4661 9112 4717
rect 9168 4661 9192 4717
rect 9248 4661 9272 4717
rect 9328 4661 9352 4717
rect 9408 4673 10660 4717
rect 10716 4673 10740 4729
rect 10796 4673 10820 4729
rect 10876 4673 10900 4729
rect 10956 4673 10980 4729
rect 11036 4673 11060 4729
rect 11116 4673 11140 4729
rect 11196 4673 12465 4729
rect 12521 4673 12545 4729
rect 12601 4673 12625 4729
rect 12681 4673 12705 4729
rect 12761 4673 12785 4729
rect 12841 4673 12865 4729
rect 12921 4673 12945 4729
rect 13001 4673 14278 4729
rect 14334 4673 14358 4729
rect 14414 4673 14438 4729
rect 14494 4673 14518 4729
rect 14574 4673 14598 4729
rect 14654 4673 14678 4729
rect 14734 4673 14758 4729
rect 14814 4673 15125 4729
rect 9408 4661 15125 4673
rect 5802 4646 15125 4661
rect 5802 4635 10660 4646
rect 5802 4608 8872 4635
rect 3016 4583 8872 4608
rect 3016 4527 3458 4583
rect 3514 4527 3538 4583
rect 3594 4527 3618 4583
rect 3674 4527 3698 4583
rect 3754 4527 3778 4583
rect 3834 4527 3858 4583
rect 3914 4527 3938 4583
rect 3994 4527 5266 4583
rect 5322 4527 5346 4583
rect 5402 4527 5426 4583
rect 5482 4527 5506 4583
rect 5562 4527 5586 4583
rect 5642 4527 5666 4583
rect 5722 4527 5746 4583
rect 5802 4579 8872 4583
rect 8928 4579 8952 4635
rect 9008 4579 9032 4635
rect 9088 4579 9112 4635
rect 9168 4579 9192 4635
rect 9248 4579 9272 4635
rect 9328 4579 9352 4635
rect 9408 4590 10660 4635
rect 10716 4590 10740 4646
rect 10796 4590 10820 4646
rect 10876 4590 10900 4646
rect 10956 4590 10980 4646
rect 11036 4590 11060 4646
rect 11116 4590 11140 4646
rect 11196 4590 12465 4646
rect 12521 4590 12545 4646
rect 12601 4590 12625 4646
rect 12681 4590 12705 4646
rect 12761 4590 12785 4646
rect 12841 4590 12865 4646
rect 12921 4590 12945 4646
rect 13001 4590 14278 4646
rect 14334 4590 14358 4646
rect 14414 4590 14438 4646
rect 14494 4590 14518 4646
rect 14574 4590 14598 4646
rect 14654 4590 14678 4646
rect 14734 4590 14758 4646
rect 14814 4590 15125 4646
rect 9408 4579 15125 4590
rect 5802 4563 15125 4579
rect 5802 4553 10660 4563
rect 5802 4527 8872 4553
rect 3016 4502 8872 4527
rect 3016 4446 3458 4502
rect 3514 4446 3538 4502
rect 3594 4446 3618 4502
rect 3674 4446 3698 4502
rect 3754 4446 3778 4502
rect 3834 4446 3858 4502
rect 3914 4446 3938 4502
rect 3994 4446 5266 4502
rect 5322 4446 5346 4502
rect 5402 4446 5426 4502
rect 5482 4446 5506 4502
rect 5562 4446 5586 4502
rect 5642 4446 5666 4502
rect 5722 4446 5746 4502
rect 5802 4497 8872 4502
rect 8928 4497 8952 4553
rect 9008 4497 9032 4553
rect 9088 4497 9112 4553
rect 9168 4497 9192 4553
rect 9248 4497 9272 4553
rect 9328 4497 9352 4553
rect 9408 4507 10660 4553
rect 10716 4507 10740 4563
rect 10796 4507 10820 4563
rect 10876 4507 10900 4563
rect 10956 4507 10980 4563
rect 11036 4507 11060 4563
rect 11116 4507 11140 4563
rect 11196 4507 12465 4563
rect 12521 4507 12545 4563
rect 12601 4507 12625 4563
rect 12681 4507 12705 4563
rect 12761 4507 12785 4563
rect 12841 4507 12865 4563
rect 12921 4507 12945 4563
rect 13001 4507 14278 4563
rect 14334 4507 14358 4563
rect 14414 4507 14438 4563
rect 14494 4507 14518 4563
rect 14574 4507 14598 4563
rect 14654 4507 14678 4563
rect 14734 4507 14758 4563
rect 14814 4507 15125 4563
rect 9408 4497 15125 4507
rect 5802 4446 15125 4497
rect 167 4284 2016 4441
rect 167 4228 865 4284
rect 921 4228 945 4284
rect 1001 4228 1025 4284
rect 1081 4228 2016 4284
rect 167 4200 2016 4228
rect 167 4144 865 4200
rect 921 4144 945 4200
rect 1001 4144 1025 4200
rect 1081 4144 2016 4200
rect 167 4116 2016 4144
rect 167 4060 865 4116
rect 921 4060 945 4116
rect 1001 4060 1025 4116
rect 1081 4060 2016 4116
rect 167 4031 2016 4060
rect 167 3975 865 4031
rect 921 3975 945 4031
rect 1001 3975 1025 4031
rect 1081 3975 2016 4031
rect 167 3946 2016 3975
rect 167 3890 865 3946
rect 921 3890 945 3946
rect 1001 3890 1025 3946
rect 1081 3890 2016 3946
rect 167 3861 2016 3890
rect 167 3805 865 3861
rect 921 3805 945 3861
rect 1001 3805 1025 3861
rect 1081 3805 2016 3861
rect 167 3776 2016 3805
rect 167 3720 865 3776
rect 921 3720 945 3776
rect 1001 3720 1025 3776
rect 1081 3720 2016 3776
rect 167 3704 2016 3720
rect 3016 4340 15125 4446
rect 3016 4132 10609 4340
rect 3016 4076 8675 4132
rect 8731 4076 8755 4132
rect 8811 4076 8835 4132
rect 8891 4076 8915 4132
rect 8971 4076 8995 4132
rect 9051 4076 10609 4132
rect 3016 4048 10609 4076
rect 3016 3992 8675 4048
rect 8731 3992 8755 4048
rect 8811 3992 8835 4048
rect 8891 3992 8915 4048
rect 8971 3992 8995 4048
rect 9051 3992 10609 4048
rect 3016 3964 10609 3992
rect 10825 4100 15125 4340
rect 10825 4044 13307 4100
rect 13363 4044 13392 4100
rect 13448 4044 13476 4100
rect 13532 4044 13560 4100
rect 13616 4044 13644 4100
rect 13700 4044 13728 4100
rect 13784 4044 13812 4100
rect 13868 4044 15125 4100
rect 10825 4020 15125 4044
rect 10825 3964 13307 4020
rect 13363 3964 13392 4020
rect 13448 3964 13476 4020
rect 13532 3964 13560 4020
rect 13616 3964 13644 4020
rect 13700 3964 13728 4020
rect 13784 3964 13812 4020
rect 13868 3964 15125 4020
rect 3016 3908 8675 3964
rect 8731 3908 8755 3964
rect 8811 3908 8835 3964
rect 8891 3908 8915 3964
rect 8971 3908 8995 3964
rect 9051 3940 15125 3964
rect 9051 3939 13307 3940
rect 9051 3908 10609 3939
rect 3016 3883 10609 3908
rect 10665 3883 10689 3939
rect 10745 3883 10769 3939
rect 10825 3884 13307 3939
rect 13363 3884 13392 3940
rect 13448 3884 13476 3940
rect 13532 3884 13560 3940
rect 13616 3884 13644 3940
rect 13700 3884 13728 3940
rect 13784 3884 13812 3940
rect 13868 3884 15125 3940
rect 10825 3883 15125 3884
rect 3016 3880 15125 3883
rect 3016 3824 8675 3880
rect 8731 3824 8755 3880
rect 8811 3824 8835 3880
rect 8891 3824 8915 3880
rect 8971 3824 8995 3880
rect 9051 3860 15125 3880
rect 9051 3858 13307 3860
rect 9051 3824 10609 3858
rect 3016 3802 10609 3824
rect 10665 3802 10689 3858
rect 10745 3802 10769 3858
rect 10825 3804 13307 3858
rect 13363 3804 13392 3860
rect 13448 3804 13476 3860
rect 13532 3804 13560 3860
rect 13616 3804 13644 3860
rect 13700 3804 13728 3860
rect 13784 3804 13812 3860
rect 13868 3804 15125 3860
rect 10825 3802 15125 3804
rect 3016 3795 15125 3802
rect 3016 3739 8675 3795
rect 8731 3739 8755 3795
rect 8811 3739 8835 3795
rect 8891 3739 8915 3795
rect 8971 3739 8995 3795
rect 9051 3780 15125 3795
rect 9051 3777 13307 3780
rect 9051 3739 10609 3777
rect 3016 3721 10609 3739
rect 10665 3721 10689 3777
rect 10745 3721 10769 3777
rect 10825 3724 13307 3777
rect 13363 3724 13392 3780
rect 13448 3724 13476 3780
rect 13532 3724 13560 3780
rect 13616 3724 13644 3780
rect 13700 3724 13728 3780
rect 13784 3724 13812 3780
rect 13868 3724 15125 3780
rect 10825 3721 15125 3724
rect 3016 3704 15125 3721
rect 16016 5556 16632 7452
rect 16016 5500 16064 5556
rect 16120 5500 16144 5556
rect 16200 5500 16224 5556
rect 16280 5500 16304 5556
rect 16360 5500 16384 5556
rect 16440 5500 16464 5556
rect 16520 5500 16632 5556
rect 16016 5474 16632 5500
rect 16016 5418 16064 5474
rect 16120 5418 16144 5474
rect 16200 5418 16224 5474
rect 16280 5418 16304 5474
rect 16360 5418 16384 5474
rect 16440 5418 16464 5474
rect 16520 5418 16632 5474
rect 16016 5392 16632 5418
rect 16016 5336 16064 5392
rect 16120 5336 16144 5392
rect 16200 5336 16224 5392
rect 16280 5336 16304 5392
rect 16360 5336 16384 5392
rect 16440 5336 16464 5392
rect 16520 5336 16632 5392
rect 16016 5310 16632 5336
rect 16016 5254 16064 5310
rect 16120 5254 16144 5310
rect 16200 5254 16224 5310
rect 16280 5254 16304 5310
rect 16360 5254 16384 5310
rect 16440 5254 16464 5310
rect 16520 5254 16632 5310
rect 16016 5228 16632 5254
rect 16016 5172 16064 5228
rect 16120 5172 16144 5228
rect 16200 5172 16224 5228
rect 16280 5172 16304 5228
rect 16360 5172 16384 5228
rect 16440 5172 16464 5228
rect 16520 5172 16632 5228
rect 16016 5146 16632 5172
rect 16016 5090 16064 5146
rect 16120 5090 16144 5146
rect 16200 5090 16224 5146
rect 16280 5090 16304 5146
rect 16360 5090 16384 5146
rect 16440 5090 16464 5146
rect 16520 5090 16632 5146
rect 16016 5064 16632 5090
rect 16016 5008 16064 5064
rect 16120 5008 16144 5064
rect 16200 5008 16224 5064
rect 16280 5008 16304 5064
rect 16360 5008 16384 5064
rect 16440 5008 16464 5064
rect 16520 5008 16632 5064
rect 16016 4982 16632 5008
rect 16016 4926 16064 4982
rect 16120 4926 16144 4982
rect 16200 4926 16224 4982
rect 16280 4926 16304 4982
rect 16360 4926 16384 4982
rect 16440 4926 16464 4982
rect 16520 4926 16632 4982
rect 16016 4900 16632 4926
rect 16016 4844 16064 4900
rect 16120 4844 16144 4900
rect 16200 4844 16224 4900
rect 16280 4844 16304 4900
rect 16360 4844 16384 4900
rect 16440 4844 16464 4900
rect 16520 4844 16632 4900
rect 16016 4818 16632 4844
rect 16016 4762 16064 4818
rect 16120 4762 16144 4818
rect 16200 4762 16224 4818
rect 16280 4762 16304 4818
rect 16360 4762 16384 4818
rect 16440 4762 16464 4818
rect 16520 4762 16632 4818
rect 16016 4735 16632 4762
rect 16016 4679 16064 4735
rect 16120 4679 16144 4735
rect 16200 4679 16224 4735
rect 16280 4679 16304 4735
rect 16360 4679 16384 4735
rect 16440 4679 16464 4735
rect 16520 4679 16632 4735
rect 28321 4685 28665 4690
rect 16016 4652 16632 4679
rect 16016 4596 16064 4652
rect 16120 4596 16144 4652
rect 16200 4596 16224 4652
rect 16280 4596 16304 4652
rect 16360 4596 16384 4652
rect 16440 4596 16464 4652
rect 16520 4596 16632 4652
rect 16016 4569 16632 4596
rect 16016 4513 16064 4569
rect 16120 4513 16144 4569
rect 16200 4513 16224 4569
rect 16280 4513 16304 4569
rect 16360 4513 16384 4569
rect 16440 4513 16464 4569
rect 16520 4513 16632 4569
rect 16016 3704 16632 4513
rect 27594 4679 27994 4684
rect 27594 4623 27606 4679
rect 27662 4623 27686 4679
rect 27742 4623 27766 4679
rect 27822 4623 27846 4679
rect 27902 4623 27926 4679
rect 27982 4623 27994 4679
rect 27594 4598 27994 4623
rect 27594 4542 27606 4598
rect 27662 4542 27686 4598
rect 27742 4542 27766 4598
rect 27822 4542 27846 4598
rect 27902 4542 27926 4598
rect 27982 4542 27994 4598
rect 27594 4517 27994 4542
rect 27594 4461 27606 4517
rect 27662 4461 27686 4517
rect 27742 4461 27766 4517
rect 27822 4461 27846 4517
rect 27902 4461 27926 4517
rect 27982 4461 27994 4517
rect 27594 4435 27994 4461
rect 27594 4379 27606 4435
rect 27662 4379 27686 4435
rect 27742 4379 27766 4435
rect 27822 4379 27846 4435
rect 27902 4379 27926 4435
rect 27982 4379 27994 4435
rect 27594 4353 27994 4379
rect 27594 4297 27606 4353
rect 27662 4297 27686 4353
rect 27742 4297 27766 4353
rect 27822 4297 27846 4353
rect 27902 4297 27926 4353
rect 27982 4297 27994 4353
rect 27594 4271 27994 4297
rect 27594 4215 27606 4271
rect 27662 4215 27686 4271
rect 27742 4215 27766 4271
rect 27822 4215 27846 4271
rect 27902 4215 27926 4271
rect 27982 4215 27994 4271
rect 27594 4189 27994 4215
rect 27594 4133 27606 4189
rect 27662 4133 27686 4189
rect 27742 4133 27766 4189
rect 27822 4133 27846 4189
rect 27902 4133 27926 4189
rect 27982 4133 27994 4189
rect 27594 4107 27994 4133
rect 27594 4051 27606 4107
rect 27662 4051 27686 4107
rect 27742 4051 27766 4107
rect 27822 4051 27846 4107
rect 27902 4051 27926 4107
rect 27982 4051 27994 4107
rect 27594 4025 27994 4051
rect 27594 3969 27606 4025
rect 27662 3969 27686 4025
rect 27742 3969 27766 4025
rect 27822 3969 27846 4025
rect 27902 3969 27926 4025
rect 27982 3969 27994 4025
rect 27594 3943 27994 3969
rect 27594 3887 27606 3943
rect 27662 3887 27686 3943
rect 27742 3887 27766 3943
rect 27822 3887 27846 3943
rect 27902 3887 27926 3943
rect 27982 3887 27994 3943
rect 27594 3861 27994 3887
rect 27594 3805 27606 3861
rect 27662 3805 27686 3861
rect 27742 3805 27766 3861
rect 27822 3805 27846 3861
rect 27902 3805 27926 3861
rect 27982 3805 27994 3861
rect 27594 3779 27994 3805
rect 27594 3723 27606 3779
rect 27662 3723 27686 3779
rect 27742 3723 27766 3779
rect 27822 3723 27846 3779
rect 27902 3723 27926 3779
rect 27982 3723 27994 3779
rect 27594 3718 27994 3723
rect 28321 4629 28345 4685
rect 28401 4629 28425 4685
rect 28481 4629 28505 4685
rect 28561 4629 28585 4685
rect 28641 4629 28665 4685
rect 28321 4603 28665 4629
rect 28321 4547 28345 4603
rect 28401 4547 28425 4603
rect 28481 4547 28505 4603
rect 28561 4547 28585 4603
rect 28641 4547 28665 4603
rect 28321 4521 28665 4547
rect 28321 4465 28345 4521
rect 28401 4465 28425 4521
rect 28481 4465 28505 4521
rect 28561 4465 28585 4521
rect 28641 4465 28665 4521
rect 28321 4439 28665 4465
rect 28321 4383 28345 4439
rect 28401 4383 28425 4439
rect 28481 4383 28505 4439
rect 28561 4383 28585 4439
rect 28641 4383 28665 4439
rect 28321 4357 28665 4383
rect 28321 4301 28345 4357
rect 28401 4301 28425 4357
rect 28481 4301 28505 4357
rect 28561 4301 28585 4357
rect 28641 4301 28665 4357
rect 28321 4275 28665 4301
rect 28321 4219 28345 4275
rect 28401 4219 28425 4275
rect 28481 4219 28505 4275
rect 28561 4219 28585 4275
rect 28641 4219 28665 4275
rect 28321 4193 28665 4219
rect 28321 4137 28345 4193
rect 28401 4137 28425 4193
rect 28481 4137 28505 4193
rect 28561 4137 28585 4193
rect 28641 4137 28665 4193
rect 28321 4111 28665 4137
rect 28321 4055 28345 4111
rect 28401 4055 28425 4111
rect 28481 4055 28505 4111
rect 28561 4055 28585 4111
rect 28641 4055 28665 4111
rect 28321 4028 28665 4055
rect 28321 3972 28345 4028
rect 28401 3972 28425 4028
rect 28481 3972 28505 4028
rect 28561 3972 28585 4028
rect 28641 3972 28665 4028
rect 28321 3945 28665 3972
rect 28321 3889 28345 3945
rect 28401 3889 28425 3945
rect 28481 3889 28505 3945
rect 28561 3889 28585 3945
rect 28641 3889 28665 3945
rect 28321 3862 28665 3889
rect 28321 3806 28345 3862
rect 28401 3806 28425 3862
rect 28481 3806 28505 3862
rect 28561 3806 28585 3862
rect 28641 3806 28665 3862
rect 28321 3779 28665 3806
rect 28321 3723 28345 3779
rect 28401 3723 28425 3779
rect 28481 3723 28505 3779
rect 28561 3723 28585 3779
rect 28641 3723 28665 3779
rect 28321 3718 28665 3723
rect 167 3188 5228 3204
rect 123 3183 5228 3188
rect 123 1447 167 3183
rect 623 3127 2288 3183
rect 2344 3127 2368 3183
rect 2424 3127 2448 3183
rect 2504 3127 2528 3183
rect 2584 3127 2608 3183
rect 2664 3127 2688 3183
rect 2744 3138 5228 3183
rect 2744 3127 4228 3138
rect 623 3093 4228 3127
rect 623 3037 2288 3093
rect 2344 3037 2368 3093
rect 2424 3037 2448 3093
rect 2504 3037 2528 3093
rect 2584 3037 2608 3093
rect 2664 3037 2688 3093
rect 2744 3082 4228 3093
rect 4284 3082 4308 3138
rect 4364 3082 4388 3138
rect 4444 3082 4468 3138
rect 4524 3082 4548 3138
rect 4604 3082 4628 3138
rect 4684 3082 4708 3138
rect 4764 3082 4788 3138
rect 4844 3082 4868 3138
rect 4924 3082 4948 3138
rect 5004 3082 5028 3138
rect 5084 3082 5228 3138
rect 2744 3057 5228 3082
rect 2744 3037 4228 3057
rect 623 3003 4228 3037
rect 623 2947 2288 3003
rect 2344 2947 2368 3003
rect 2424 2947 2448 3003
rect 2504 2947 2528 3003
rect 2584 2947 2608 3003
rect 2664 2947 2688 3003
rect 2744 3001 4228 3003
rect 4284 3001 4308 3057
rect 4364 3001 4388 3057
rect 4444 3001 4468 3057
rect 4524 3001 4548 3057
rect 4604 3001 4628 3057
rect 4684 3001 4708 3057
rect 4764 3001 4788 3057
rect 4844 3001 4868 3057
rect 4924 3001 4948 3057
rect 5004 3001 5028 3057
rect 5084 3001 5228 3057
rect 2744 2976 5228 3001
rect 2744 2947 4228 2976
rect 623 2920 4228 2947
rect 4284 2920 4308 2976
rect 4364 2920 4388 2976
rect 4444 2920 4468 2976
rect 4524 2920 4548 2976
rect 4604 2920 4628 2976
rect 4684 2920 4708 2976
rect 4764 2920 4788 2976
rect 4844 2920 4868 2976
rect 4924 2920 4948 2976
rect 5004 2920 5028 2976
rect 5084 2920 5228 2976
rect 623 2913 5228 2920
rect 623 2857 2288 2913
rect 2344 2857 2368 2913
rect 2424 2857 2448 2913
rect 2504 2857 2528 2913
rect 2584 2857 2608 2913
rect 2664 2857 2688 2913
rect 2744 2895 5228 2913
rect 2744 2857 4228 2895
rect 623 2839 4228 2857
rect 4284 2839 4308 2895
rect 4364 2839 4388 2895
rect 4444 2839 4468 2895
rect 4524 2839 4548 2895
rect 4604 2839 4628 2895
rect 4684 2839 4708 2895
rect 4764 2839 4788 2895
rect 4844 2839 4868 2895
rect 4924 2839 4948 2895
rect 5004 2839 5028 2895
rect 5084 2839 5228 2895
rect 623 2823 5228 2839
rect 623 2767 2288 2823
rect 2344 2767 2368 2823
rect 2424 2767 2448 2823
rect 2504 2767 2528 2823
rect 2584 2767 2608 2823
rect 2664 2767 2688 2823
rect 2744 2814 5228 2823
rect 2744 2767 4228 2814
rect 623 2758 4228 2767
rect 4284 2758 4308 2814
rect 4364 2758 4388 2814
rect 4444 2758 4468 2814
rect 4524 2758 4548 2814
rect 4604 2758 4628 2814
rect 4684 2758 4708 2814
rect 4764 2758 4788 2814
rect 4844 2758 4868 2814
rect 4924 2758 4948 2814
rect 5004 2758 5028 2814
rect 5084 2758 5228 2814
rect 623 2733 5228 2758
rect 623 2677 2288 2733
rect 2344 2677 2368 2733
rect 2424 2677 2448 2733
rect 2504 2677 2528 2733
rect 2584 2677 2608 2733
rect 2664 2677 2688 2733
rect 2744 2677 4228 2733
rect 4284 2677 4308 2733
rect 4364 2677 4388 2733
rect 4444 2677 4468 2733
rect 4524 2677 4548 2733
rect 4604 2677 4628 2733
rect 4684 2677 4708 2733
rect 4764 2677 4788 2733
rect 4844 2677 4868 2733
rect 4924 2677 4948 2733
rect 5004 2677 5028 2733
rect 5084 2677 5228 2733
rect 623 2652 5228 2677
rect 623 2642 4228 2652
rect 623 2586 2288 2642
rect 2344 2586 2368 2642
rect 2424 2586 2448 2642
rect 2504 2586 2528 2642
rect 2584 2586 2608 2642
rect 2664 2586 2688 2642
rect 2744 2596 4228 2642
rect 4284 2596 4308 2652
rect 4364 2596 4388 2652
rect 4444 2596 4468 2652
rect 4524 2596 4548 2652
rect 4604 2596 4628 2652
rect 4684 2596 4708 2652
rect 4764 2596 4788 2652
rect 4844 2596 4868 2652
rect 4924 2596 4948 2652
rect 5004 2596 5028 2652
rect 5084 2596 5228 2652
rect 2744 2586 5228 2596
rect 623 2571 5228 2586
rect 623 2551 4228 2571
rect 623 2495 2288 2551
rect 2344 2495 2368 2551
rect 2424 2495 2448 2551
rect 2504 2495 2528 2551
rect 2584 2495 2608 2551
rect 2664 2495 2688 2551
rect 2744 2515 4228 2551
rect 4284 2515 4308 2571
rect 4364 2515 4388 2571
rect 4444 2515 4468 2571
rect 4524 2515 4548 2571
rect 4604 2515 4628 2571
rect 4684 2515 4708 2571
rect 4764 2515 4788 2571
rect 4844 2515 4868 2571
rect 4924 2515 4948 2571
rect 5004 2515 5028 2571
rect 5084 2515 5228 2571
rect 2744 2495 5228 2515
rect 623 2490 5228 2495
rect 623 2434 4228 2490
rect 4284 2434 4308 2490
rect 4364 2434 4388 2490
rect 4444 2434 4468 2490
rect 4524 2434 4548 2490
rect 4604 2434 4628 2490
rect 4684 2434 4708 2490
rect 4764 2434 4788 2490
rect 4844 2434 4868 2490
rect 4924 2434 4948 2490
rect 5004 2434 5028 2490
rect 5084 2434 5228 2490
rect 623 2408 5228 2434
rect 623 2352 4228 2408
rect 4284 2352 4308 2408
rect 4364 2352 4388 2408
rect 4444 2352 4468 2408
rect 4524 2352 4548 2408
rect 4604 2352 4628 2408
rect 4684 2352 4708 2408
rect 4764 2352 4788 2408
rect 4844 2352 4868 2408
rect 4924 2352 4948 2408
rect 5004 2352 5028 2408
rect 5084 2352 5228 2408
rect 623 2326 5228 2352
rect 623 2270 4228 2326
rect 4284 2270 4308 2326
rect 4364 2270 4388 2326
rect 4444 2270 4468 2326
rect 4524 2270 4548 2326
rect 4604 2270 4628 2326
rect 4684 2270 4708 2326
rect 4764 2270 4788 2326
rect 4844 2270 4868 2326
rect 4924 2270 4948 2326
rect 5004 2270 5028 2326
rect 5084 2270 5228 2326
rect 623 2244 5228 2270
rect 623 2188 4228 2244
rect 4284 2188 4308 2244
rect 4364 2188 4388 2244
rect 4444 2188 4468 2244
rect 4524 2188 4548 2244
rect 4604 2188 4628 2244
rect 4684 2188 4708 2244
rect 4764 2188 4788 2244
rect 4844 2188 4868 2244
rect 4924 2188 4948 2244
rect 5004 2188 5028 2244
rect 5084 2188 5228 2244
rect 623 2162 5228 2188
rect 623 2106 4228 2162
rect 4284 2106 4308 2162
rect 4364 2106 4388 2162
rect 4444 2106 4468 2162
rect 4524 2106 4548 2162
rect 4604 2106 4628 2162
rect 4684 2106 4708 2162
rect 4764 2106 4788 2162
rect 4844 2106 4868 2162
rect 4924 2106 4948 2162
rect 5004 2106 5028 2162
rect 5084 2106 5228 2162
rect 623 2080 5228 2106
rect 623 2024 4228 2080
rect 4284 2024 4308 2080
rect 4364 2024 4388 2080
rect 4444 2024 4468 2080
rect 4524 2024 4548 2080
rect 4604 2024 4628 2080
rect 4684 2024 4708 2080
rect 4764 2024 4788 2080
rect 4844 2024 4868 2080
rect 4924 2024 4948 2080
rect 5004 2024 5028 2080
rect 5084 2024 5228 2080
rect 623 2018 5228 2024
rect 623 1962 1594 2018
rect 1650 1962 1674 2018
rect 1730 1962 1754 2018
rect 1810 1962 1834 2018
rect 1890 1962 2415 2018
rect 2471 1962 2495 2018
rect 2551 1962 2575 2018
rect 2631 1962 2655 2018
rect 2711 1998 5228 2018
rect 2711 1962 4228 1998
rect 623 1942 4228 1962
rect 4284 1942 4308 1998
rect 4364 1942 4388 1998
rect 4444 1942 4468 1998
rect 4524 1942 4548 1998
rect 4604 1942 4628 1998
rect 4684 1942 4708 1998
rect 4764 1942 4788 1998
rect 4844 1942 4868 1998
rect 4924 1942 4948 1998
rect 5004 1942 5028 1998
rect 5084 1942 5228 1998
rect 623 1932 5228 1942
rect 623 1876 1594 1932
rect 1650 1876 1674 1932
rect 1730 1876 1754 1932
rect 1810 1876 1834 1932
rect 1890 1876 2415 1932
rect 2471 1876 2495 1932
rect 2551 1876 2575 1932
rect 2631 1876 2655 1932
rect 2711 1916 5228 1932
rect 2711 1876 4228 1916
rect 623 1860 4228 1876
rect 4284 1860 4308 1916
rect 4364 1860 4388 1916
rect 4444 1860 4468 1916
rect 4524 1860 4548 1916
rect 4604 1860 4628 1916
rect 4684 1860 4708 1916
rect 4764 1860 4788 1916
rect 4844 1860 4868 1916
rect 4924 1860 4948 1916
rect 5004 1860 5028 1916
rect 5084 1860 5228 1916
rect 623 1846 5228 1860
rect 623 1790 1594 1846
rect 1650 1790 1674 1846
rect 1730 1790 1754 1846
rect 1810 1790 1834 1846
rect 1890 1790 2415 1846
rect 2471 1790 2495 1846
rect 2551 1790 2575 1846
rect 2631 1790 2655 1846
rect 2711 1790 5228 1846
rect 623 1760 5228 1790
rect 623 1704 1594 1760
rect 1650 1704 1674 1760
rect 1730 1704 1754 1760
rect 1810 1704 1834 1760
rect 1890 1704 2415 1760
rect 2471 1704 2495 1760
rect 2551 1704 2575 1760
rect 2631 1704 2655 1760
rect 2711 1704 5228 1760
rect 623 1693 5228 1704
rect 623 1674 3161 1693
rect 623 1618 1594 1674
rect 1650 1618 1674 1674
rect 1730 1618 1754 1674
rect 1810 1618 1834 1674
rect 1890 1618 2415 1674
rect 2471 1618 2495 1674
rect 2551 1618 2575 1674
rect 2631 1618 2655 1674
rect 2711 1637 3161 1674
rect 3217 1637 3241 1693
rect 3297 1637 5228 1693
rect 2711 1618 5228 1637
rect 623 1601 5228 1618
rect 623 1587 3161 1601
rect 623 1531 1594 1587
rect 1650 1531 1674 1587
rect 1730 1531 1754 1587
rect 1810 1531 1834 1587
rect 1890 1531 2415 1587
rect 2471 1531 2495 1587
rect 2551 1531 2575 1587
rect 2631 1531 2655 1587
rect 2711 1545 3161 1587
rect 3217 1545 3241 1601
rect 3297 1545 5228 1601
rect 2711 1531 5228 1545
rect 623 1530 5228 1531
rect 623 1508 3321 1530
rect 623 1500 3161 1508
rect 623 1447 1594 1500
rect 123 1444 1594 1447
rect 1650 1444 1674 1500
rect 1730 1444 1754 1500
rect 1810 1444 1834 1500
rect 1890 1444 2415 1500
rect 2471 1444 2495 1500
rect 2551 1444 2575 1500
rect 2631 1444 2655 1500
rect 2711 1452 3161 1500
rect 3217 1452 3241 1508
rect 3297 1474 3321 1508
rect 3377 1474 3401 1530
rect 3457 1474 5228 1530
rect 3297 1452 5228 1474
rect 2711 1444 5228 1452
rect 123 1422 5228 1444
rect 123 1366 167 1422
rect 223 1366 247 1422
rect 303 1366 327 1422
rect 383 1366 407 1422
rect 463 1366 487 1422
rect 543 1366 567 1422
rect 623 1418 5228 1422
rect 623 1415 3321 1418
rect 623 1413 3161 1415
rect 623 1366 1594 1413
rect 123 1361 1594 1366
rect 167 1357 1594 1361
rect 1650 1357 1674 1413
rect 1730 1357 1754 1413
rect 1810 1357 1834 1413
rect 1890 1357 2415 1413
rect 2471 1357 2495 1413
rect 2551 1357 2575 1413
rect 2631 1357 2655 1413
rect 2711 1359 3161 1413
rect 3217 1359 3241 1415
rect 3297 1362 3321 1415
rect 3377 1362 3401 1418
rect 3457 1362 5228 1418
rect 3297 1359 5228 1362
rect 2711 1357 5228 1359
rect 167 1344 5228 1357
rect 6497 3149 8275 3204
rect 6497 3093 6798 3149
rect 6854 3093 6884 3149
rect 6940 3093 6970 3149
rect 7026 3093 7056 3149
rect 7112 3093 7142 3149
rect 7198 3093 7228 3149
rect 7284 3093 7314 3149
rect 7370 3093 7400 3149
rect 7456 3093 7486 3149
rect 7542 3093 7572 3149
rect 7628 3093 7657 3149
rect 7713 3093 8275 3149
rect 6497 3069 8275 3093
rect 6497 3013 6798 3069
rect 6854 3013 6884 3069
rect 6940 3013 6970 3069
rect 7026 3013 7056 3069
rect 7112 3013 7142 3069
rect 7198 3013 7228 3069
rect 7284 3013 7314 3069
rect 7370 3013 7400 3069
rect 7456 3013 7486 3069
rect 7542 3013 7572 3069
rect 7628 3013 7657 3069
rect 7713 3013 8275 3069
rect 6497 2989 8275 3013
rect 6497 2933 6798 2989
rect 6854 2933 6884 2989
rect 6940 2933 6970 2989
rect 7026 2933 7056 2989
rect 7112 2933 7142 2989
rect 7198 2933 7228 2989
rect 7284 2933 7314 2989
rect 7370 2933 7400 2989
rect 7456 2933 7486 2989
rect 7542 2933 7572 2989
rect 7628 2933 7657 2989
rect 7713 2933 8275 2989
rect 6497 2909 8275 2933
rect 6497 2853 6798 2909
rect 6854 2853 6884 2909
rect 6940 2853 6970 2909
rect 7026 2853 7056 2909
rect 7112 2853 7142 2909
rect 7198 2853 7228 2909
rect 7284 2853 7314 2909
rect 7370 2853 7400 2909
rect 7456 2853 7486 2909
rect 7542 2853 7572 2909
rect 7628 2853 7657 2909
rect 7713 2853 8275 2909
rect 6497 2829 8275 2853
rect 6497 2773 6798 2829
rect 6854 2773 6884 2829
rect 6940 2773 6970 2829
rect 7026 2773 7056 2829
rect 7112 2773 7142 2829
rect 7198 2773 7228 2829
rect 7284 2773 7314 2829
rect 7370 2773 7400 2829
rect 7456 2773 7486 2829
rect 7542 2773 7572 2829
rect 7628 2773 7657 2829
rect 7713 2773 8275 2829
rect 6497 2749 8275 2773
rect 6497 2693 6798 2749
rect 6854 2693 6884 2749
rect 6940 2693 6970 2749
rect 7026 2693 7056 2749
rect 7112 2693 7142 2749
rect 7198 2693 7228 2749
rect 7284 2693 7314 2749
rect 7370 2693 7400 2749
rect 7456 2693 7486 2749
rect 7542 2693 7572 2749
rect 7628 2693 7657 2749
rect 7713 2693 8275 2749
rect 6497 2669 8275 2693
rect 6497 2613 6798 2669
rect 6854 2613 6884 2669
rect 6940 2613 6970 2669
rect 7026 2613 7056 2669
rect 7112 2613 7142 2669
rect 7198 2613 7228 2669
rect 7284 2613 7314 2669
rect 7370 2613 7400 2669
rect 7456 2613 7486 2669
rect 7542 2613 7572 2669
rect 7628 2613 7657 2669
rect 7713 2613 8275 2669
rect 6497 2589 8275 2613
rect 6497 2533 6798 2589
rect 6854 2533 6884 2589
rect 6940 2533 6970 2589
rect 7026 2533 7056 2589
rect 7112 2533 7142 2589
rect 7198 2533 7228 2589
rect 7284 2533 7314 2589
rect 7370 2533 7400 2589
rect 7456 2533 7486 2589
rect 7542 2533 7572 2589
rect 7628 2533 7657 2589
rect 7713 2533 8275 2589
rect 6497 1831 8275 2533
rect 6497 1775 7794 1831
rect 7850 1775 7874 1831
rect 7930 1775 7954 1831
rect 8010 1775 8034 1831
rect 8090 1775 8114 1831
rect 8170 1775 8194 1831
rect 8250 1775 8275 1831
rect 6497 1748 8275 1775
rect 6497 1692 7794 1748
rect 7850 1692 7874 1748
rect 7930 1692 7954 1748
rect 8010 1692 8034 1748
rect 8090 1692 8114 1748
rect 8170 1692 8194 1748
rect 8250 1692 8275 1748
rect 6497 1665 8275 1692
rect 6497 1609 7794 1665
rect 7850 1609 7874 1665
rect 7930 1609 7954 1665
rect 8010 1609 8034 1665
rect 8090 1609 8114 1665
rect 8170 1609 8194 1665
rect 8250 1609 8275 1665
rect 6497 1582 8275 1609
rect 6497 1526 7794 1582
rect 7850 1526 7874 1582
rect 7930 1526 7954 1582
rect 8010 1526 8034 1582
rect 8090 1526 8114 1582
rect 8170 1526 8194 1582
rect 8250 1526 8275 1582
rect 6497 1498 8275 1526
rect 6497 1442 7794 1498
rect 7850 1442 7874 1498
rect 7930 1442 7954 1498
rect 8010 1442 8034 1498
rect 8090 1442 8114 1498
rect 8170 1442 8194 1498
rect 8250 1442 8275 1498
rect 6497 1414 8275 1442
rect 6497 1358 7794 1414
rect 7850 1358 7874 1414
rect 7930 1358 7954 1414
rect 8010 1358 8034 1414
rect 8090 1358 8114 1414
rect 8170 1358 8194 1414
rect 8250 1358 8275 1414
rect 6497 1344 8275 1358
rect 9475 3145 10916 3204
rect 9475 3089 9602 3145
rect 9658 3089 9682 3145
rect 9738 3089 9762 3145
rect 9818 3089 9842 3145
rect 9898 3089 9922 3145
rect 9978 3089 10002 3145
rect 10058 3089 10082 3145
rect 10138 3089 10162 3145
rect 10218 3089 10242 3145
rect 10298 3089 10916 3145
rect 9475 3058 10916 3089
rect 9475 3002 9602 3058
rect 9658 3002 9682 3058
rect 9738 3002 9762 3058
rect 9818 3002 9842 3058
rect 9898 3002 9922 3058
rect 9978 3002 10002 3058
rect 10058 3002 10082 3058
rect 10138 3002 10162 3058
rect 10218 3002 10242 3058
rect 10298 3002 10916 3058
rect 9475 2971 10916 3002
rect 9475 2915 9602 2971
rect 9658 2915 9682 2971
rect 9738 2915 9762 2971
rect 9818 2915 9842 2971
rect 9898 2915 9922 2971
rect 9978 2915 10002 2971
rect 10058 2915 10082 2971
rect 10138 2915 10162 2971
rect 10218 2915 10242 2971
rect 10298 2915 10916 2971
rect 9475 2884 10916 2915
rect 9475 2828 9602 2884
rect 9658 2828 9682 2884
rect 9738 2828 9762 2884
rect 9818 2828 9842 2884
rect 9898 2828 9922 2884
rect 9978 2828 10002 2884
rect 10058 2828 10082 2884
rect 10138 2828 10162 2884
rect 10218 2828 10242 2884
rect 10298 2828 10916 2884
rect 9475 2797 10916 2828
rect 9475 2741 9602 2797
rect 9658 2741 9682 2797
rect 9738 2741 9762 2797
rect 9818 2741 9842 2797
rect 9898 2741 9922 2797
rect 9978 2741 10002 2797
rect 10058 2741 10082 2797
rect 10138 2741 10162 2797
rect 10218 2741 10242 2797
rect 10298 2741 10916 2797
rect 9475 2710 10916 2741
rect 9475 2654 9602 2710
rect 9658 2654 9682 2710
rect 9738 2654 9762 2710
rect 9818 2654 9842 2710
rect 9898 2654 9922 2710
rect 9978 2654 10002 2710
rect 10058 2654 10082 2710
rect 10138 2654 10162 2710
rect 10218 2654 10242 2710
rect 10298 2654 10916 2710
rect 9475 2623 10916 2654
rect 9475 2567 9602 2623
rect 9658 2567 9682 2623
rect 9738 2567 9762 2623
rect 9818 2567 9842 2623
rect 9898 2567 9922 2623
rect 9978 2567 10002 2623
rect 10058 2567 10082 2623
rect 10138 2567 10162 2623
rect 10218 2567 10242 2623
rect 10298 2567 10916 2623
rect 9475 2536 10916 2567
rect 9475 2480 9602 2536
rect 9658 2480 9682 2536
rect 9738 2480 9762 2536
rect 9818 2480 9842 2536
rect 9898 2480 9922 2536
rect 9978 2480 10002 2536
rect 10058 2480 10082 2536
rect 10138 2480 10162 2536
rect 10218 2480 10242 2536
rect 10298 2480 10916 2536
rect 9475 2448 10916 2480
rect 9475 2392 9602 2448
rect 9658 2392 9682 2448
rect 9738 2392 9762 2448
rect 9818 2392 9842 2448
rect 9898 2392 9922 2448
rect 9978 2392 10002 2448
rect 10058 2392 10082 2448
rect 10138 2392 10162 2448
rect 10218 2392 10242 2448
rect 10298 2392 10916 2448
rect 9475 2360 10916 2392
rect 9475 2304 9602 2360
rect 9658 2304 9682 2360
rect 9738 2304 9762 2360
rect 9818 2304 9842 2360
rect 9898 2304 9922 2360
rect 9978 2304 10002 2360
rect 10058 2304 10082 2360
rect 10138 2304 10162 2360
rect 10218 2304 10242 2360
rect 10298 2304 10916 2360
rect 9475 2272 10916 2304
rect 9475 2216 9602 2272
rect 9658 2216 9682 2272
rect 9738 2216 9762 2272
rect 9818 2216 9842 2272
rect 9898 2216 9922 2272
rect 9978 2216 10002 2272
rect 10058 2216 10082 2272
rect 10138 2216 10162 2272
rect 10218 2216 10242 2272
rect 10298 2216 10916 2272
rect 9475 2049 10916 2216
rect 9475 1993 9735 2049
rect 9791 1993 9815 2049
rect 9871 1993 9895 2049
rect 9951 1993 10916 2049
rect 9475 1959 10916 1993
rect 9475 1903 9735 1959
rect 9791 1903 9815 1959
rect 9871 1903 9895 1959
rect 9951 1903 10916 1959
rect 9475 1869 10916 1903
rect 9475 1813 9735 1869
rect 9791 1813 9815 1869
rect 9871 1813 9895 1869
rect 9951 1813 10916 1869
rect 9475 1779 10916 1813
rect 9475 1723 9735 1779
rect 9791 1723 9815 1779
rect 9871 1723 9895 1779
rect 9951 1723 10916 1779
rect 9475 1689 10916 1723
rect 9475 1633 9735 1689
rect 9791 1633 9815 1689
rect 9871 1633 9895 1689
rect 9951 1633 10916 1689
rect 9475 1599 10916 1633
rect 9475 1543 9735 1599
rect 9791 1543 9815 1599
rect 9871 1543 9895 1599
rect 9951 1543 10916 1599
rect 9475 1509 10916 1543
rect 9475 1453 9735 1509
rect 9791 1453 9815 1509
rect 9871 1453 9895 1509
rect 9951 1453 10916 1509
rect 9475 1418 10916 1453
rect 9475 1362 9735 1418
rect 9791 1362 9815 1418
rect 9871 1362 9895 1418
rect 9951 1362 10916 1418
rect 9475 1344 10916 1362
rect 12116 3190 15234 3204
rect 12116 2494 12194 3190
rect 12650 3159 15234 3190
rect 12650 3103 13972 3159
rect 14028 3103 14063 3159
rect 14119 3103 14154 3159
rect 14210 3103 14244 3159
rect 14300 3103 14334 3159
rect 14390 3103 14424 3159
rect 14480 3103 14514 3159
rect 14570 3145 15234 3159
rect 14570 3103 14630 3145
rect 12650 3089 14630 3103
rect 14686 3089 14718 3145
rect 14774 3089 14806 3145
rect 14862 3089 14894 3145
rect 14950 3089 14982 3145
rect 15038 3089 15070 3145
rect 15126 3089 15158 3145
rect 15214 3089 15234 3145
rect 12650 3079 15234 3089
rect 12650 3023 13972 3079
rect 14028 3023 14063 3079
rect 14119 3023 14154 3079
rect 14210 3023 14244 3079
rect 14300 3023 14334 3079
rect 14390 3023 14424 3079
rect 14480 3023 14514 3079
rect 14570 3065 15234 3079
rect 23413 3189 23623 3194
rect 14570 3023 14630 3065
rect 12650 3009 14630 3023
rect 14686 3009 14718 3065
rect 14774 3009 14806 3065
rect 14862 3009 14894 3065
rect 14950 3009 14982 3065
rect 15038 3009 15070 3065
rect 15126 3009 15158 3065
rect 15214 3009 15234 3065
rect 12650 2999 15234 3009
rect 12650 2943 13972 2999
rect 14028 2943 14063 2999
rect 14119 2943 14154 2999
rect 14210 2943 14244 2999
rect 14300 2943 14334 2999
rect 14390 2943 14424 2999
rect 14480 2943 14514 2999
rect 14570 2985 15234 2999
rect 14570 2943 14630 2985
rect 12650 2929 14630 2943
rect 14686 2929 14718 2985
rect 14774 2929 14806 2985
rect 14862 2929 14894 2985
rect 14950 2929 14982 2985
rect 15038 2929 15070 2985
rect 15126 2929 15158 2985
rect 15214 2929 15234 2985
rect 12650 2919 15234 2929
rect 12650 2863 13972 2919
rect 14028 2863 14063 2919
rect 14119 2863 14154 2919
rect 14210 2863 14244 2919
rect 14300 2863 14334 2919
rect 14390 2863 14424 2919
rect 14480 2863 14514 2919
rect 14570 2905 15234 2919
rect 14570 2863 14630 2905
rect 12650 2849 14630 2863
rect 14686 2849 14718 2905
rect 14774 2849 14806 2905
rect 14862 2849 14894 2905
rect 14950 2849 14982 2905
rect 15038 2849 15070 2905
rect 15126 2849 15158 2905
rect 15214 2849 15234 2905
rect 12650 2839 15234 2849
rect 12650 2783 13972 2839
rect 14028 2783 14063 2839
rect 14119 2783 14154 2839
rect 14210 2783 14244 2839
rect 14300 2783 14334 2839
rect 14390 2783 14424 2839
rect 14480 2783 14514 2839
rect 14570 2789 15234 2839
rect 14570 2783 14641 2789
rect 12650 2759 14641 2783
rect 12650 2703 13972 2759
rect 14028 2703 14063 2759
rect 14119 2703 14154 2759
rect 14210 2703 14244 2759
rect 14300 2703 14334 2759
rect 14390 2703 14424 2759
rect 14480 2703 14514 2759
rect 14570 2733 14641 2759
rect 14697 2733 14721 2789
rect 14777 2733 14801 2789
rect 14857 2733 15234 2789
rect 14570 2703 15234 2733
rect 12650 2679 15234 2703
rect 12650 2623 13972 2679
rect 14028 2623 14063 2679
rect 14119 2623 14154 2679
rect 14210 2623 14244 2679
rect 14300 2623 14334 2679
rect 14390 2623 14424 2679
rect 14480 2623 14514 2679
rect 14570 2677 15234 2679
rect 14570 2623 14641 2677
rect 12650 2621 14641 2623
rect 14697 2621 14721 2677
rect 14777 2621 14801 2677
rect 14857 2621 15234 2677
rect 12650 2599 15234 2621
rect 12650 2543 13972 2599
rect 14028 2543 14063 2599
rect 14119 2543 14154 2599
rect 14210 2543 14244 2599
rect 14300 2543 14334 2599
rect 14390 2543 14424 2599
rect 14480 2543 14514 2599
rect 14570 2564 15234 2599
rect 14570 2543 14641 2564
rect 12650 2519 14641 2543
rect 12650 2494 13972 2519
rect 12116 2469 13972 2494
rect 12116 2413 12194 2469
rect 12250 2413 12274 2469
rect 12330 2413 12354 2469
rect 12410 2413 12434 2469
rect 12490 2413 12514 2469
rect 12570 2413 12594 2469
rect 12650 2463 13972 2469
rect 14028 2463 14063 2519
rect 14119 2463 14154 2519
rect 14210 2463 14244 2519
rect 14300 2463 14334 2519
rect 14390 2463 14424 2519
rect 14480 2463 14514 2519
rect 14570 2508 14641 2519
rect 14697 2508 14721 2564
rect 14777 2508 14801 2564
rect 14857 2508 15234 2564
rect 14570 2463 15234 2508
rect 12650 2439 15234 2463
rect 12650 2413 13972 2439
rect 12116 2388 13972 2413
rect 12116 2332 12194 2388
rect 12250 2332 12274 2388
rect 12330 2332 12354 2388
rect 12410 2332 12434 2388
rect 12490 2332 12514 2388
rect 12570 2332 12594 2388
rect 12650 2383 13972 2388
rect 14028 2383 14063 2439
rect 14119 2383 14154 2439
rect 14210 2383 14244 2439
rect 14300 2383 14334 2439
rect 14390 2383 14424 2439
rect 14480 2383 14514 2439
rect 14570 2383 15234 2439
rect 12650 2359 15234 2383
rect 12650 2332 13972 2359
rect 12116 2307 13972 2332
rect 12116 2251 12194 2307
rect 12250 2251 12274 2307
rect 12330 2251 12354 2307
rect 12410 2251 12434 2307
rect 12490 2251 12514 2307
rect 12570 2251 12594 2307
rect 12650 2303 13972 2307
rect 14028 2303 14063 2359
rect 14119 2303 14154 2359
rect 14210 2303 14244 2359
rect 14300 2303 14334 2359
rect 14390 2303 14424 2359
rect 14480 2303 14514 2359
rect 14570 2303 15234 2359
rect 12650 2279 15234 2303
rect 12650 2251 13972 2279
rect 12116 2226 13972 2251
rect 12116 2170 12194 2226
rect 12250 2170 12274 2226
rect 12330 2170 12354 2226
rect 12410 2170 12434 2226
rect 12490 2170 12514 2226
rect 12570 2170 12594 2226
rect 12650 2223 13972 2226
rect 14028 2223 14063 2279
rect 14119 2223 14154 2279
rect 14210 2223 14244 2279
rect 14300 2223 14334 2279
rect 14390 2223 14424 2279
rect 14480 2223 14514 2279
rect 14570 2223 15234 2279
rect 12650 2170 15234 2223
rect 12116 2145 15234 2170
rect 12116 2089 12194 2145
rect 12250 2089 12274 2145
rect 12330 2089 12354 2145
rect 12410 2089 12434 2145
rect 12490 2089 12514 2145
rect 12570 2089 12594 2145
rect 12650 2089 15234 2145
rect 12116 2064 15234 2089
rect 12116 2008 12194 2064
rect 12250 2008 12274 2064
rect 12330 2008 12354 2064
rect 12410 2008 12434 2064
rect 12490 2008 12514 2064
rect 12570 2008 12594 2064
rect 12650 2008 15234 2064
rect 12116 1983 15234 2008
rect 12116 1927 12194 1983
rect 12250 1927 12274 1983
rect 12330 1927 12354 1983
rect 12410 1927 12434 1983
rect 12490 1927 12514 1983
rect 12570 1927 12594 1983
rect 12650 1927 15234 1983
rect 12116 1902 15234 1927
rect 12116 1846 12194 1902
rect 12250 1846 12274 1902
rect 12330 1846 12354 1902
rect 12410 1846 12434 1902
rect 12490 1846 12514 1902
rect 12570 1846 12594 1902
rect 12650 1846 15234 1902
rect 22085 3063 22151 3068
rect 22085 3007 22090 3063
rect 22146 3007 22151 3063
rect 22085 2983 22151 3007
rect 22085 2927 22090 2983
rect 22146 2927 22151 2983
rect 22085 2903 22151 2927
rect 22085 2847 22090 2903
rect 22146 2847 22151 2903
rect 22085 2823 22151 2847
rect 22085 2767 22090 2823
rect 22146 2767 22151 2823
rect 22085 2743 22151 2767
rect 22085 2687 22090 2743
rect 22146 2687 22151 2743
rect 22085 2663 22151 2687
rect 22085 2607 22090 2663
rect 22146 2607 22151 2663
rect 22085 2583 22151 2607
rect 22085 2527 22090 2583
rect 22146 2527 22151 2583
rect 22085 2503 22151 2527
rect 22085 2447 22090 2503
rect 22146 2447 22151 2503
rect 22085 2423 22151 2447
rect 22085 2367 22090 2423
rect 22146 2367 22151 2423
rect 22085 2343 22151 2367
rect 22085 2287 22090 2343
rect 22146 2287 22151 2343
rect 22085 2263 22151 2287
rect 22085 2207 22090 2263
rect 22146 2207 22151 2263
rect 22085 2183 22151 2207
rect 22085 2127 22090 2183
rect 22146 2127 22151 2183
rect 22085 2103 22151 2127
rect 22085 2047 22090 2103
rect 22146 2047 22151 2103
rect 22085 2023 22151 2047
rect 22085 1967 22090 2023
rect 22146 1967 22151 2023
rect 22085 1943 22151 1967
rect 12116 1821 15234 1846
rect 12116 1765 12194 1821
rect 12250 1765 12274 1821
rect 12330 1765 12354 1821
rect 12410 1765 12434 1821
rect 12490 1765 12514 1821
rect 12570 1765 12594 1821
rect 12650 1765 15234 1821
rect 12116 1740 15234 1765
rect 12116 1684 12194 1740
rect 12250 1684 12274 1740
rect 12330 1684 12354 1740
rect 12410 1684 12434 1740
rect 12490 1684 12514 1740
rect 12570 1684 12594 1740
rect 12650 1684 15234 1740
rect 12116 1659 15234 1684
rect 12116 1603 12194 1659
rect 12250 1603 12274 1659
rect 12330 1603 12354 1659
rect 12410 1603 12434 1659
rect 12490 1603 12514 1659
rect 12570 1603 12594 1659
rect 12650 1603 15234 1659
rect 15619 1895 15977 1900
rect 12116 1578 15234 1603
rect 12116 1522 12194 1578
rect 12250 1522 12274 1578
rect 12330 1522 12354 1578
rect 12410 1522 12434 1578
rect 12490 1522 12514 1578
rect 12570 1522 12594 1578
rect 12650 1522 15234 1578
rect 12116 1497 15234 1522
rect 12116 1441 12194 1497
rect 12250 1441 12274 1497
rect 12330 1441 12354 1497
rect 12410 1441 12434 1497
rect 12490 1441 12514 1497
rect 12570 1441 12594 1497
rect 12650 1441 15234 1497
rect 12116 1416 15234 1441
rect 12116 1360 12194 1416
rect 12250 1360 12274 1416
rect 12330 1360 12354 1416
rect 12410 1360 12434 1416
rect 12490 1360 12514 1416
rect 12570 1360 12594 1416
rect 12650 1360 15234 1416
rect 15375 1638 15601 1643
rect 15375 1582 15380 1638
rect 15436 1582 15460 1638
rect 15516 1582 15540 1638
rect 15596 1582 15601 1638
rect 15375 1530 15601 1582
rect 15375 1474 15380 1530
rect 15436 1474 15460 1530
rect 15516 1474 15540 1530
rect 15596 1474 15601 1530
rect 15375 1421 15601 1474
rect 15375 1365 15380 1421
rect 15436 1365 15460 1421
rect 15516 1365 15540 1421
rect 15596 1365 15601 1421
rect 15375 1360 15601 1365
rect 12116 1344 15234 1360
rect 15619 1359 15650 1895
rect 15946 1359 15977 1895
rect 22085 1887 22090 1943
rect 22146 1887 22151 1943
rect 22085 1863 22151 1887
rect 22085 1807 22090 1863
rect 22146 1807 22151 1863
rect 22085 1782 22151 1807
rect 22085 1726 22090 1782
rect 22146 1726 22151 1782
rect 22085 1701 22151 1726
rect 22085 1645 22090 1701
rect 22146 1645 22151 1701
rect 22085 1620 22151 1645
rect 22085 1564 22090 1620
rect 22146 1564 22151 1620
rect 22085 1539 22151 1564
rect 22085 1483 22090 1539
rect 22146 1483 22151 1539
rect 22085 1478 22151 1483
rect 23413 2493 23450 3189
rect 23586 2493 23623 3189
rect 23413 2468 23623 2493
rect 23413 2412 23450 2468
rect 23506 2412 23530 2468
rect 23586 2412 23623 2468
rect 23413 2387 23623 2412
rect 23413 2331 23450 2387
rect 23506 2331 23530 2387
rect 23586 2331 23623 2387
rect 23413 2306 23623 2331
rect 23413 2250 23450 2306
rect 23506 2250 23530 2306
rect 23586 2250 23623 2306
rect 23413 2225 23623 2250
rect 23413 2169 23450 2225
rect 23506 2169 23530 2225
rect 23586 2169 23623 2225
rect 23413 2144 23623 2169
rect 23413 2088 23450 2144
rect 23506 2088 23530 2144
rect 23586 2088 23623 2144
rect 23413 2063 23623 2088
rect 23413 2007 23450 2063
rect 23506 2007 23530 2063
rect 23586 2007 23623 2063
rect 23413 1982 23623 2007
rect 23413 1926 23450 1982
rect 23506 1926 23530 1982
rect 23586 1926 23623 1982
rect 23413 1901 23623 1926
rect 23413 1845 23450 1901
rect 23506 1845 23530 1901
rect 23586 1845 23623 1901
rect 23413 1820 23623 1845
rect 23413 1764 23450 1820
rect 23506 1764 23530 1820
rect 23586 1764 23623 1820
rect 23413 1739 23623 1764
rect 23413 1683 23450 1739
rect 23506 1683 23530 1739
rect 23586 1683 23623 1739
rect 23413 1658 23623 1683
rect 23413 1602 23450 1658
rect 23506 1602 23530 1658
rect 23586 1602 23623 1658
rect 23413 1577 23623 1602
rect 23413 1521 23450 1577
rect 23506 1521 23530 1577
rect 23586 1521 23623 1577
rect 23413 1496 23623 1521
rect 15619 1354 15977 1359
rect 23413 1440 23450 1496
rect 23506 1440 23530 1496
rect 23586 1440 23623 1496
rect 23413 1415 23623 1440
rect 23413 1359 23450 1415
rect 23506 1359 23530 1415
rect 23586 1359 23623 1415
rect 23413 1354 23623 1359
rect 24152 3190 24428 3195
rect 24152 2734 24182 3190
rect 24398 2734 24428 3190
rect 24152 2709 24428 2734
rect 24152 2653 24182 2709
rect 24238 2653 24262 2709
rect 24318 2653 24342 2709
rect 24398 2653 24428 2709
rect 24152 2628 24428 2653
rect 24152 2572 24182 2628
rect 24238 2572 24262 2628
rect 24318 2572 24342 2628
rect 24398 2572 24428 2628
rect 24152 2547 24428 2572
rect 24152 2491 24182 2547
rect 24238 2491 24262 2547
rect 24318 2491 24342 2547
rect 24398 2491 24428 2547
rect 24152 2466 24428 2491
rect 24152 2410 24182 2466
rect 24238 2410 24262 2466
rect 24318 2410 24342 2466
rect 24398 2410 24428 2466
rect 24152 2385 24428 2410
rect 24152 2329 24182 2385
rect 24238 2329 24262 2385
rect 24318 2329 24342 2385
rect 24398 2329 24428 2385
rect 24152 2304 24428 2329
rect 24152 2248 24182 2304
rect 24238 2248 24262 2304
rect 24318 2248 24342 2304
rect 24398 2248 24428 2304
rect 24152 2223 24428 2248
rect 24152 2167 24182 2223
rect 24238 2167 24262 2223
rect 24318 2167 24342 2223
rect 24398 2167 24428 2223
rect 24152 2142 24428 2167
rect 24152 2086 24182 2142
rect 24238 2086 24262 2142
rect 24318 2086 24342 2142
rect 24398 2086 24428 2142
rect 24152 2061 24428 2086
rect 24152 2005 24182 2061
rect 24238 2005 24262 2061
rect 24318 2005 24342 2061
rect 24398 2005 24428 2061
rect 24152 1980 24428 2005
rect 24152 1924 24182 1980
rect 24238 1924 24262 1980
rect 24318 1924 24342 1980
rect 24398 1924 24428 1980
rect 24152 1899 24428 1924
rect 24152 1843 24182 1899
rect 24238 1843 24262 1899
rect 24318 1843 24342 1899
rect 24398 1843 24428 1899
rect 24152 1818 24428 1843
rect 24152 1762 24182 1818
rect 24238 1762 24262 1818
rect 24318 1762 24342 1818
rect 24398 1762 24428 1818
rect 24152 1737 24428 1762
rect 24152 1681 24182 1737
rect 24238 1681 24262 1737
rect 24318 1681 24342 1737
rect 24398 1681 24428 1737
rect 24152 1656 24428 1681
rect 24152 1600 24182 1656
rect 24238 1600 24262 1656
rect 24318 1600 24342 1656
rect 24398 1600 24428 1656
rect 24152 1575 24428 1600
rect 24152 1519 24182 1575
rect 24238 1519 24262 1575
rect 24318 1519 24342 1575
rect 24398 1519 24428 1575
rect 24152 1494 24428 1519
rect 24152 1438 24182 1494
rect 24238 1438 24262 1494
rect 24318 1438 24342 1494
rect 24398 1438 24428 1494
rect 24152 1413 24428 1438
rect 24152 1357 24182 1413
rect 24238 1357 24262 1413
rect 24318 1357 24342 1413
rect 24398 1357 24428 1413
rect 25888 2436 26382 2441
rect 25888 2380 25907 2436
rect 25963 2380 25987 2436
rect 26043 2380 26067 2436
rect 26123 2380 26147 2436
rect 26203 2380 26227 2436
rect 26283 2380 26307 2436
rect 26363 2380 26382 2436
rect 25888 2353 26382 2380
rect 25888 2297 25907 2353
rect 25963 2297 25987 2353
rect 26043 2297 26067 2353
rect 26123 2297 26147 2353
rect 26203 2297 26227 2353
rect 26283 2297 26307 2353
rect 26363 2297 26382 2353
rect 25888 2270 26382 2297
rect 25888 2214 25907 2270
rect 25963 2214 25987 2270
rect 26043 2214 26067 2270
rect 26123 2214 26147 2270
rect 26203 2214 26227 2270
rect 26283 2214 26307 2270
rect 26363 2214 26382 2270
rect 25888 2187 26382 2214
rect 25888 2131 25907 2187
rect 25963 2131 25987 2187
rect 26043 2131 26067 2187
rect 26123 2131 26147 2187
rect 26203 2131 26227 2187
rect 26283 2131 26307 2187
rect 26363 2131 26382 2187
rect 25888 2104 26382 2131
rect 25888 2048 25907 2104
rect 25963 2048 25987 2104
rect 26043 2048 26067 2104
rect 26123 2048 26147 2104
rect 26203 2048 26227 2104
rect 26283 2048 26307 2104
rect 26363 2048 26382 2104
rect 25888 2021 26382 2048
rect 25888 1965 25907 2021
rect 25963 1965 25987 2021
rect 26043 1965 26067 2021
rect 26123 1965 26147 2021
rect 26203 1965 26227 2021
rect 26283 1965 26307 2021
rect 26363 1965 26382 2021
rect 25888 1938 26382 1965
rect 25888 1882 25907 1938
rect 25963 1882 25987 1938
rect 26043 1882 26067 1938
rect 26123 1882 26147 1938
rect 26203 1882 26227 1938
rect 26283 1882 26307 1938
rect 26363 1882 26382 1938
rect 25888 1855 26382 1882
rect 25888 1799 25907 1855
rect 25963 1799 25987 1855
rect 26043 1799 26067 1855
rect 26123 1799 26147 1855
rect 26203 1799 26227 1855
rect 26283 1799 26307 1855
rect 26363 1799 26382 1855
rect 25888 1771 26382 1799
rect 25888 1715 25907 1771
rect 25963 1715 25987 1771
rect 26043 1715 26067 1771
rect 26123 1715 26147 1771
rect 26203 1715 26227 1771
rect 26283 1715 26307 1771
rect 26363 1715 26382 1771
rect 25888 1687 26382 1715
rect 25888 1631 25907 1687
rect 25963 1631 25987 1687
rect 26043 1631 26067 1687
rect 26123 1631 26147 1687
rect 26203 1631 26227 1687
rect 26283 1631 26307 1687
rect 26363 1631 26382 1687
rect 25888 1603 26382 1631
rect 25888 1547 25907 1603
rect 25963 1547 25987 1603
rect 26043 1547 26067 1603
rect 26123 1547 26147 1603
rect 26203 1547 26227 1603
rect 26283 1547 26307 1603
rect 26363 1547 26382 1603
rect 25888 1519 26382 1547
rect 25888 1463 25907 1519
rect 25963 1463 25987 1519
rect 26043 1463 26067 1519
rect 26123 1463 26147 1519
rect 26203 1463 26227 1519
rect 26283 1463 26307 1519
rect 26363 1463 26382 1519
rect 25888 1435 26382 1463
rect 25888 1379 25907 1435
rect 25963 1379 25987 1435
rect 26043 1379 26067 1435
rect 26123 1379 26147 1435
rect 26203 1379 26227 1435
rect 26283 1379 26307 1435
rect 26363 1379 26382 1435
rect 25888 1374 26382 1379
rect 24152 1352 24428 1357
rect 13296 832 13541 837
rect 2751 824 3039 829
rect 2751 -752 2787 824
rect 3003 -752 3039 824
rect 10381 827 10847 832
rect 10381 771 10386 827
rect 10442 771 10466 827
rect 10522 771 10546 827
rect 10602 771 10626 827
rect 10682 771 10706 827
rect 10762 771 10786 827
rect 10842 771 10847 827
rect 10381 740 10847 771
rect 10381 684 10386 740
rect 10442 684 10466 740
rect 10522 684 10546 740
rect 10602 684 10626 740
rect 10682 684 10706 740
rect 10762 684 10786 740
rect 10842 684 10847 740
rect 10381 652 10847 684
rect 10381 596 10386 652
rect 10442 596 10466 652
rect 10522 596 10546 652
rect 10602 596 10626 652
rect 10682 596 10706 652
rect 10762 596 10786 652
rect 10842 596 10847 652
rect 10381 564 10847 596
rect 10381 508 10386 564
rect 10442 508 10466 564
rect 10522 508 10546 564
rect 10602 508 10626 564
rect 10682 508 10706 564
rect 10762 508 10786 564
rect 10842 508 10847 564
rect 10381 476 10847 508
rect 10381 420 10386 476
rect 10442 420 10466 476
rect 10522 420 10546 476
rect 10602 420 10626 476
rect 10682 420 10706 476
rect 10762 420 10786 476
rect 10842 420 10847 476
rect 13296 776 13320 832
rect 13376 776 13400 832
rect 13456 776 13480 832
rect 13536 776 13541 832
rect 13296 746 13541 776
rect 13296 690 13320 746
rect 13376 690 13400 746
rect 13456 737 13541 746
rect 13456 690 13480 737
rect 13296 681 13480 690
rect 13536 681 13541 737
rect 13296 660 13541 681
rect 13296 604 13320 660
rect 13376 604 13400 660
rect 13456 641 13541 660
rect 13456 604 13480 641
rect 13296 585 13480 604
rect 13536 585 13541 641
rect 13296 574 13541 585
rect 13296 518 13320 574
rect 13376 518 13400 574
rect 13456 545 13541 574
rect 13555 832 13621 837
rect 13555 776 13560 832
rect 13616 776 13621 832
rect 13555 730 13621 776
rect 13555 674 13560 730
rect 13616 674 13621 730
rect 13555 628 13621 674
rect 13635 832 13701 837
rect 13635 776 13640 832
rect 13696 776 13701 832
rect 13635 706 13701 776
rect 13715 794 13781 837
rect 13715 738 13720 794
rect 13776 738 13781 794
rect 13715 733 13781 738
rect 27594 822 27994 827
rect 27594 766 27606 822
rect 27662 766 27686 822
rect 27742 766 27766 822
rect 27822 766 27846 822
rect 27902 766 27926 822
rect 27982 766 27994 822
rect 27594 741 27994 766
rect 13635 650 13640 706
rect 13696 650 13701 706
rect 13635 645 13701 650
rect 27594 685 27606 741
rect 27662 685 27686 741
rect 27742 685 27766 741
rect 27822 685 27846 741
rect 27902 685 27926 741
rect 27982 685 27994 741
rect 27594 660 27994 685
rect 13555 572 13560 628
rect 13616 572 13621 628
rect 13555 567 13621 572
rect 27594 604 27606 660
rect 27662 604 27686 660
rect 27742 604 27766 660
rect 27822 604 27846 660
rect 27902 604 27926 660
rect 27982 604 27994 660
rect 27594 579 27994 604
rect 13456 518 13480 545
rect 13296 489 13480 518
rect 13536 489 13541 545
rect 13296 487 13541 489
rect 13296 431 13320 487
rect 13376 431 13400 487
rect 13456 484 13541 487
rect 27594 523 27606 579
rect 27662 523 27686 579
rect 27742 523 27766 579
rect 27822 523 27846 579
rect 27902 523 27926 579
rect 27982 523 27994 579
rect 27594 498 27994 523
rect 13456 431 13480 484
rect 13296 426 13480 431
rect 27594 442 27606 498
rect 27662 442 27686 498
rect 27742 442 27766 498
rect 27822 442 27846 498
rect 27902 442 27926 498
rect 27982 442 27994 498
rect 10381 388 10847 420
rect 10381 332 10386 388
rect 10442 332 10466 388
rect 10522 332 10546 388
rect 10602 332 10626 388
rect 10682 332 10706 388
rect 10762 332 10786 388
rect 10842 332 10847 388
rect 10381 300 10847 332
rect 10381 244 10386 300
rect 10442 244 10466 300
rect 10522 244 10546 300
rect 10602 244 10626 300
rect 10682 244 10706 300
rect 10762 244 10786 300
rect 10842 244 10847 300
rect 10381 239 10847 244
rect 27594 417 27994 442
rect 27594 361 27606 417
rect 27662 361 27686 417
rect 27742 361 27766 417
rect 27822 361 27846 417
rect 27902 361 27926 417
rect 27982 361 27994 417
rect 27594 335 27994 361
rect 27594 279 27606 335
rect 27662 279 27686 335
rect 27742 279 27766 335
rect 27822 279 27846 335
rect 27902 279 27926 335
rect 27982 279 27994 335
rect 27594 253 27994 279
rect 27594 197 27606 253
rect 27662 197 27686 253
rect 27742 197 27766 253
rect 27822 197 27846 253
rect 27902 197 27926 253
rect 27982 197 27994 253
rect 27594 171 27994 197
rect 27594 115 27606 171
rect 27662 115 27686 171
rect 27742 115 27766 171
rect 27822 115 27846 171
rect 27902 115 27926 171
rect 27982 115 27994 171
rect 27594 89 27994 115
rect 27594 33 27606 89
rect 27662 33 27686 89
rect 27742 33 27766 89
rect 27822 33 27846 89
rect 27902 33 27926 89
rect 27982 33 27994 89
rect 27594 7 27994 33
rect 27594 -49 27606 7
rect 27662 -49 27686 7
rect 27742 -49 27766 7
rect 27822 -49 27846 7
rect 27902 -49 27926 7
rect 27982 -49 27994 7
rect 27594 -75 27994 -49
rect 27594 -131 27606 -75
rect 27662 -131 27686 -75
rect 27742 -131 27766 -75
rect 27822 -131 27846 -75
rect 27902 -131 27926 -75
rect 27982 -131 27994 -75
rect 27594 -157 27994 -131
rect 27594 -213 27606 -157
rect 27662 -213 27686 -157
rect 27742 -213 27766 -157
rect 27822 -213 27846 -157
rect 27902 -213 27926 -157
rect 27982 -213 27994 -157
rect 27594 -239 27994 -213
rect 27594 -295 27606 -239
rect 27662 -295 27686 -239
rect 27742 -295 27766 -239
rect 27822 -295 27846 -239
rect 27902 -295 27926 -239
rect 27982 -295 27994 -239
rect 27594 -321 27994 -295
rect 27594 -377 27606 -321
rect 27662 -377 27686 -321
rect 27742 -377 27766 -321
rect 27822 -377 27846 -321
rect 27902 -377 27926 -321
rect 27982 -377 27994 -321
rect 27594 -403 27994 -377
rect 27594 -459 27606 -403
rect 27662 -459 27686 -403
rect 27742 -459 27766 -403
rect 27822 -459 27846 -403
rect 27902 -459 27926 -403
rect 27982 -459 27994 -403
rect 27594 -464 27994 -459
rect 28321 806 28665 811
rect 28321 270 28345 806
rect 28641 270 28665 806
rect 28321 245 28665 270
rect 28321 189 28345 245
rect 28401 189 28425 245
rect 28481 189 28505 245
rect 28561 189 28585 245
rect 28641 189 28665 245
rect 28321 164 28665 189
rect 28321 108 28345 164
rect 28401 108 28425 164
rect 28481 108 28505 164
rect 28561 108 28585 164
rect 28641 108 28665 164
rect 28321 83 28665 108
rect 28321 27 28345 83
rect 28401 27 28425 83
rect 28481 27 28505 83
rect 28561 27 28585 83
rect 28641 27 28665 83
rect 28321 2 28665 27
rect 28321 -54 28345 2
rect 28401 -54 28425 2
rect 28481 -54 28505 2
rect 28561 -54 28585 2
rect 28641 -54 28665 2
rect 28321 -79 28665 -54
rect 28321 -135 28345 -79
rect 28401 -135 28425 -79
rect 28481 -135 28505 -79
rect 28561 -135 28585 -79
rect 28641 -135 28665 -79
rect 28321 -160 28665 -135
rect 28321 -216 28345 -160
rect 28401 -216 28425 -160
rect 28481 -216 28505 -160
rect 28561 -216 28585 -160
rect 28641 -216 28665 -160
rect 28321 -241 28665 -216
rect 28321 -297 28345 -241
rect 28401 -297 28425 -241
rect 28481 -297 28505 -241
rect 28561 -297 28585 -241
rect 28641 -297 28665 -241
rect 28321 -322 28665 -297
rect 28321 -378 28345 -322
rect 28401 -378 28425 -322
rect 28481 -378 28505 -322
rect 28561 -378 28585 -322
rect 28641 -378 28665 -322
rect 28321 -403 28665 -378
rect 28321 -459 28345 -403
rect 28401 -459 28425 -403
rect 28481 -459 28505 -403
rect 28561 -459 28585 -403
rect 28641 -459 28665 -403
rect 28321 -464 28665 -459
rect 2751 -777 3039 -752
rect 2751 -833 2787 -777
rect 2843 -833 2867 -777
rect 2923 -833 2947 -777
rect 3003 -833 3039 -777
rect 2751 -858 3039 -833
rect 2751 -914 2787 -858
rect 2843 -914 2867 -858
rect 2923 -914 2947 -858
rect 3003 -914 3039 -858
rect 2751 -939 3039 -914
rect 2751 -995 2787 -939
rect 2843 -995 2867 -939
rect 2923 -995 2947 -939
rect 3003 -995 3039 -939
rect 2751 -1020 3039 -995
rect 2751 -1076 2787 -1020
rect 2843 -1076 2867 -1020
rect 2923 -1076 2947 -1020
rect 3003 -1076 3039 -1020
rect 2751 -1101 3039 -1076
rect 2751 -1157 2787 -1101
rect 2843 -1157 2867 -1101
rect 2923 -1157 2947 -1101
rect 3003 -1157 3039 -1101
rect 2751 -1182 3039 -1157
rect 2751 -1238 2787 -1182
rect 2843 -1238 2867 -1182
rect 2923 -1238 2947 -1182
rect 3003 -1238 3039 -1182
rect 2751 -1263 3039 -1238
rect 2751 -1319 2787 -1263
rect 2843 -1319 2867 -1263
rect 2923 -1319 2947 -1263
rect 3003 -1319 3039 -1263
rect 2751 -1344 3039 -1319
rect 2751 -1400 2787 -1344
rect 2843 -1400 2867 -1344
rect 2923 -1400 2947 -1344
rect 3003 -1400 3039 -1344
rect 2751 -1425 3039 -1400
rect 2751 -1481 2787 -1425
rect 2843 -1481 2867 -1425
rect 2923 -1481 2947 -1425
rect 3003 -1481 3039 -1425
rect 2751 -1506 3039 -1481
rect 2751 -1562 2787 -1506
rect 2843 -1562 2867 -1506
rect 2923 -1562 2947 -1506
rect 3003 -1562 3039 -1506
rect 2751 -1587 3039 -1562
rect 2751 -1643 2787 -1587
rect 2843 -1643 2867 -1587
rect 2923 -1643 2947 -1587
rect 3003 -1643 3039 -1587
rect 2751 -1668 3039 -1643
rect 2751 -1724 2787 -1668
rect 2843 -1724 2867 -1668
rect 2923 -1724 2947 -1668
rect 3003 -1724 3039 -1668
rect 2751 -1749 3039 -1724
rect 2751 -1805 2787 -1749
rect 2843 -1805 2867 -1749
rect 2923 -1805 2947 -1749
rect 3003 -1805 3039 -1749
rect 2751 -1830 3039 -1805
rect 2751 -1886 2787 -1830
rect 2843 -1886 2867 -1830
rect 2923 -1886 2947 -1830
rect 3003 -1886 3039 -1830
rect 2751 -1911 3039 -1886
rect 2751 -1967 2787 -1911
rect 2843 -1967 2867 -1911
rect 2923 -1967 2947 -1911
rect 3003 -1967 3039 -1911
rect 2751 -1972 3039 -1967
tri 341 -1990 343 -1988 ne
tri 9056 -1990 9058 -1988 nw
rect 9723 -2871 9949 -2866
rect 9723 -2927 9728 -2871
rect 9784 -2927 9808 -2871
rect 9864 -2927 9888 -2871
rect 9944 -2927 9949 -2871
rect 23413 -2873 23621 -2868
rect 9723 -2955 9949 -2927
rect 9723 -3011 9728 -2955
rect 9784 -3011 9808 -2955
rect 9864 -3011 9888 -2955
rect 9944 -3011 9949 -2955
rect 9723 -3039 9949 -3011
rect 9723 -3095 9728 -3039
rect 9784 -3095 9808 -3039
rect 9864 -3095 9888 -3039
rect 9944 -3095 9949 -3039
rect 9723 -3123 9949 -3095
rect 9723 -3179 9728 -3123
rect 9784 -3179 9808 -3123
rect 9864 -3179 9888 -3123
rect 9944 -3179 9949 -3123
rect 9723 -3207 9949 -3179
rect 9723 -3263 9728 -3207
rect 9784 -3263 9808 -3207
rect 9864 -3263 9888 -3207
rect 9944 -3263 9949 -3207
rect 9723 -3291 9949 -3263
rect 9723 -3347 9728 -3291
rect 9784 -3347 9808 -3291
rect 9864 -3347 9888 -3291
rect 9944 -3347 9949 -3291
rect 9723 -3375 9949 -3347
rect 9723 -3431 9728 -3375
rect 9784 -3431 9808 -3375
rect 9864 -3431 9888 -3375
rect 9944 -3431 9949 -3375
rect 9723 -3459 9949 -3431
rect 9723 -3515 9728 -3459
rect 9784 -3515 9808 -3459
rect 9864 -3515 9888 -3459
rect 9944 -3515 9949 -3459
rect 9723 -3543 9949 -3515
rect 9723 -3599 9728 -3543
rect 9784 -3599 9808 -3543
rect 9864 -3599 9888 -3543
rect 9944 -3599 9949 -3543
rect 9723 -3628 9949 -3599
rect 9723 -3684 9728 -3628
rect 9784 -3684 9808 -3628
rect 9864 -3684 9888 -3628
rect 9944 -3684 9949 -3628
rect 9723 -3689 9949 -3684
rect 15210 -2881 15978 -2876
rect 15210 -2937 15246 -2881
rect 15302 -2937 15326 -2881
rect 15382 -2937 15406 -2881
rect 15462 -2937 15486 -2881
rect 15542 -2937 15566 -2881
rect 15622 -2937 15646 -2881
rect 15702 -2937 15726 -2881
rect 15782 -2937 15806 -2881
rect 15862 -2937 15886 -2881
rect 15942 -2937 15978 -2881
rect 15210 -2964 15978 -2937
rect 15210 -3020 15246 -2964
rect 15302 -3020 15326 -2964
rect 15382 -3020 15406 -2964
rect 15462 -3020 15486 -2964
rect 15542 -3020 15566 -2964
rect 15622 -3020 15646 -2964
rect 15702 -3020 15726 -2964
rect 15782 -3020 15806 -2964
rect 15862 -3020 15886 -2964
rect 15942 -3020 15978 -2964
rect 15210 -3047 15978 -3020
rect 15210 -3103 15246 -3047
rect 15302 -3103 15326 -3047
rect 15382 -3103 15406 -3047
rect 15462 -3103 15486 -3047
rect 15542 -3103 15566 -3047
rect 15622 -3103 15646 -3047
rect 15702 -3103 15726 -3047
rect 15782 -3103 15806 -3047
rect 15862 -3103 15886 -3047
rect 15942 -3103 15978 -3047
rect 15210 -3131 15978 -3103
rect 15210 -3187 15246 -3131
rect 15302 -3187 15326 -3131
rect 15382 -3187 15406 -3131
rect 15462 -3187 15486 -3131
rect 15542 -3187 15566 -3131
rect 15622 -3187 15646 -3131
rect 15702 -3187 15726 -3131
rect 15782 -3187 15806 -3131
rect 15862 -3187 15886 -3131
rect 15942 -3187 15978 -3131
rect 15210 -3215 15978 -3187
rect 15210 -3271 15246 -3215
rect 15302 -3271 15326 -3215
rect 15382 -3271 15406 -3215
rect 15462 -3271 15486 -3215
rect 15542 -3271 15566 -3215
rect 15622 -3271 15646 -3215
rect 15702 -3271 15726 -3215
rect 15782 -3271 15806 -3215
rect 15862 -3271 15886 -3215
rect 15942 -3271 15978 -3215
rect 15210 -3299 15978 -3271
rect 15210 -3355 15246 -3299
rect 15302 -3355 15326 -3299
rect 15382 -3355 15406 -3299
rect 15462 -3355 15486 -3299
rect 15542 -3355 15566 -3299
rect 15622 -3355 15646 -3299
rect 15702 -3355 15726 -3299
rect 15782 -3355 15806 -3299
rect 15862 -3355 15886 -3299
rect 15942 -3355 15978 -3299
rect 15210 -3383 15978 -3355
rect 15210 -3439 15246 -3383
rect 15302 -3439 15326 -3383
rect 15382 -3439 15406 -3383
rect 15462 -3439 15486 -3383
rect 15542 -3439 15566 -3383
rect 15622 -3439 15646 -3383
rect 15702 -3439 15726 -3383
rect 15782 -3439 15806 -3383
rect 15862 -3439 15886 -3383
rect 15942 -3439 15978 -3383
rect 15210 -3467 15978 -3439
rect 15210 -3523 15246 -3467
rect 15302 -3523 15326 -3467
rect 15382 -3523 15406 -3467
rect 15462 -3523 15486 -3467
rect 15542 -3523 15566 -3467
rect 15622 -3523 15646 -3467
rect 15702 -3523 15726 -3467
rect 15782 -3523 15806 -3467
rect 15862 -3523 15886 -3467
rect 15942 -3523 15978 -3467
rect 15210 -3551 15978 -3523
rect 15210 -3607 15246 -3551
rect 15302 -3607 15326 -3551
rect 15382 -3607 15406 -3551
rect 15462 -3607 15486 -3551
rect 15542 -3607 15566 -3551
rect 15622 -3607 15646 -3551
rect 15702 -3607 15726 -3551
rect 15782 -3607 15806 -3551
rect 15862 -3607 15886 -3551
rect 15942 -3607 15978 -3551
rect 15210 -3635 15978 -3607
rect 15210 -3691 15246 -3635
rect 15302 -3691 15326 -3635
rect 15382 -3691 15406 -3635
rect 15462 -3691 15486 -3635
rect 15542 -3691 15566 -3635
rect 15622 -3691 15646 -3635
rect 15702 -3691 15726 -3635
rect 15782 -3691 15806 -3635
rect 15862 -3691 15886 -3635
rect 15942 -3691 15978 -3635
rect 15210 -3696 15978 -3691
rect 23413 -2929 23449 -2873
rect 23505 -2929 23529 -2873
rect 23585 -2929 23621 -2873
rect 23413 -2958 23621 -2929
rect 23413 -3014 23449 -2958
rect 23505 -3014 23529 -2958
rect 23585 -3014 23621 -2958
rect 23413 -3043 23621 -3014
rect 23413 -3099 23449 -3043
rect 23505 -3099 23529 -3043
rect 23585 -3099 23621 -3043
rect 23413 -3128 23621 -3099
rect 23413 -3184 23449 -3128
rect 23505 -3184 23529 -3128
rect 23585 -3184 23621 -3128
rect 23413 -3214 23621 -3184
rect 23413 -3270 23449 -3214
rect 23505 -3270 23529 -3214
rect 23585 -3270 23621 -3214
rect 23413 -3300 23621 -3270
rect 23413 -3356 23449 -3300
rect 23505 -3356 23529 -3300
rect 23585 -3356 23621 -3300
rect 23413 -3386 23621 -3356
rect 23413 -3442 23449 -3386
rect 23505 -3442 23529 -3386
rect 23585 -3442 23621 -3386
rect 23413 -3472 23621 -3442
rect 23413 -3528 23449 -3472
rect 23505 -3528 23529 -3472
rect 23585 -3528 23621 -3472
rect 23413 -3558 23621 -3528
rect 23413 -3614 23449 -3558
rect 23505 -3614 23529 -3558
rect 23585 -3614 23621 -3558
rect 23413 -3644 23621 -3614
rect 23413 -3700 23449 -3644
rect 23505 -3700 23529 -3644
rect 23585 -3700 23621 -3644
rect 23413 -3705 23621 -3700
rect 24155 -2871 24427 -2866
rect 24155 -2927 24183 -2871
rect 24239 -2927 24263 -2871
rect 24319 -2927 24343 -2871
rect 24399 -2927 24427 -2871
rect 24155 -2957 24427 -2927
rect 24155 -3013 24183 -2957
rect 24239 -3013 24263 -2957
rect 24319 -3013 24343 -2957
rect 24399 -3013 24427 -2957
rect 24155 -3043 24427 -3013
rect 24155 -3099 24183 -3043
rect 24239 -3099 24263 -3043
rect 24319 -3099 24343 -3043
rect 24399 -3099 24427 -3043
rect 24155 -3129 24427 -3099
rect 24155 -3185 24183 -3129
rect 24239 -3185 24263 -3129
rect 24319 -3185 24343 -3129
rect 24399 -3185 24427 -3129
rect 24155 -3215 24427 -3185
rect 24155 -3271 24183 -3215
rect 24239 -3271 24263 -3215
rect 24319 -3271 24343 -3215
rect 24399 -3271 24427 -3215
rect 24155 -3301 24427 -3271
rect 24155 -3357 24183 -3301
rect 24239 -3357 24263 -3301
rect 24319 -3357 24343 -3301
rect 24399 -3357 24427 -3301
rect 24155 -3387 24427 -3357
rect 24155 -3443 24183 -3387
rect 24239 -3443 24263 -3387
rect 24319 -3443 24343 -3387
rect 24399 -3443 24427 -3387
rect 24155 -3473 24427 -3443
rect 24155 -3529 24183 -3473
rect 24239 -3529 24263 -3473
rect 24319 -3529 24343 -3473
rect 24399 -3529 24427 -3473
rect 24155 -3559 24427 -3529
rect 24155 -3615 24183 -3559
rect 24239 -3615 24263 -3559
rect 24319 -3615 24343 -3559
rect 24399 -3615 24427 -3559
rect 24155 -3646 24427 -3615
rect 24155 -3702 24183 -3646
rect 24239 -3702 24263 -3646
rect 24319 -3702 24343 -3646
rect 24399 -3702 24427 -3646
rect 25877 -2878 26389 -2873
rect 25877 -2934 25905 -2878
rect 25961 -2934 25985 -2878
rect 26041 -2934 26065 -2878
rect 26121 -2934 26145 -2878
rect 26201 -2934 26225 -2878
rect 26281 -2934 26305 -2878
rect 26361 -2934 26389 -2878
rect 25877 -2962 26389 -2934
rect 25877 -3018 25905 -2962
rect 25961 -3018 25985 -2962
rect 26041 -3018 26065 -2962
rect 26121 -3018 26145 -2962
rect 26201 -3018 26225 -2962
rect 26281 -3018 26305 -2962
rect 26361 -3018 26389 -2962
rect 25877 -3046 26389 -3018
rect 25877 -3102 25905 -3046
rect 25961 -3102 25985 -3046
rect 26041 -3102 26065 -3046
rect 26121 -3102 26145 -3046
rect 26201 -3102 26225 -3046
rect 26281 -3102 26305 -3046
rect 26361 -3102 26389 -3046
rect 25877 -3131 26389 -3102
rect 25877 -3187 25905 -3131
rect 25961 -3187 25985 -3131
rect 26041 -3187 26065 -3131
rect 26121 -3187 26145 -3131
rect 26201 -3187 26225 -3131
rect 26281 -3187 26305 -3131
rect 26361 -3187 26389 -3131
rect 25877 -3216 26389 -3187
rect 25877 -3272 25905 -3216
rect 25961 -3272 25985 -3216
rect 26041 -3272 26065 -3216
rect 26121 -3272 26145 -3216
rect 26201 -3272 26225 -3216
rect 26281 -3272 26305 -3216
rect 26361 -3272 26389 -3216
rect 25877 -3301 26389 -3272
rect 25877 -3357 25905 -3301
rect 25961 -3357 25985 -3301
rect 26041 -3357 26065 -3301
rect 26121 -3357 26145 -3301
rect 26201 -3357 26225 -3301
rect 26281 -3357 26305 -3301
rect 26361 -3357 26389 -3301
rect 25877 -3386 26389 -3357
rect 25877 -3442 25905 -3386
rect 25961 -3442 25985 -3386
rect 26041 -3442 26065 -3386
rect 26121 -3442 26145 -3386
rect 26201 -3442 26225 -3386
rect 26281 -3442 26305 -3386
rect 26361 -3442 26389 -3386
rect 25877 -3471 26389 -3442
rect 25877 -3527 25905 -3471
rect 25961 -3527 25985 -3471
rect 26041 -3527 26065 -3471
rect 26121 -3527 26145 -3471
rect 26201 -3527 26225 -3471
rect 26281 -3527 26305 -3471
rect 26361 -3527 26389 -3471
rect 25877 -3556 26389 -3527
rect 25877 -3612 25905 -3556
rect 25961 -3612 25985 -3556
rect 26041 -3612 26065 -3556
rect 26121 -3612 26145 -3556
rect 26201 -3612 26225 -3556
rect 26281 -3612 26305 -3556
rect 26361 -3612 26389 -3556
rect 25877 -3641 26389 -3612
rect 25877 -3697 25905 -3641
rect 25961 -3697 25985 -3641
rect 26041 -3697 26065 -3641
rect 26121 -3697 26145 -3641
rect 26201 -3697 26225 -3641
rect 26281 -3697 26305 -3641
rect 26361 -3697 26389 -3641
rect 25877 -3702 26389 -3697
rect 24155 -3707 24427 -3702
rect 21539 -4231 22091 -4226
rect 21539 -4287 21547 -4231
rect 21603 -4287 21627 -4231
rect 21683 -4287 21707 -4231
rect 21763 -4287 21787 -4231
rect 21843 -4287 21867 -4231
rect 21923 -4287 21947 -4231
rect 22003 -4287 22027 -4231
rect 22083 -4287 22091 -4231
rect 21539 -4321 22091 -4287
rect 21539 -4377 21547 -4321
rect 21603 -4377 21627 -4321
rect 21683 -4377 21707 -4321
rect 21763 -4377 21787 -4321
rect 21843 -4377 21867 -4321
rect 21923 -4377 21947 -4321
rect 22003 -4377 22027 -4321
rect 22083 -4377 22091 -4321
rect 21539 -4411 22091 -4377
rect 21539 -4467 21547 -4411
rect 21603 -4467 21627 -4411
rect 21683 -4467 21707 -4411
rect 21763 -4467 21787 -4411
rect 21843 -4467 21867 -4411
rect 21923 -4467 21947 -4411
rect 22003 -4467 22027 -4411
rect 22083 -4467 22091 -4411
rect 21539 -4502 22091 -4467
rect 21539 -4558 21547 -4502
rect 21603 -4558 21627 -4502
rect 21683 -4558 21707 -4502
rect 21763 -4558 21787 -4502
rect 21843 -4558 21867 -4502
rect 21923 -4558 21947 -4502
rect 22003 -4558 22027 -4502
rect 22083 -4558 22091 -4502
rect 21539 -4593 22091 -4558
rect 21539 -4649 21547 -4593
rect 21603 -4649 21627 -4593
rect 21683 -4649 21707 -4593
rect 21763 -4649 21787 -4593
rect 21843 -4649 21867 -4593
rect 21923 -4649 21947 -4593
rect 22003 -4649 22027 -4593
rect 22083 -4649 22091 -4593
rect 21539 -4684 22091 -4649
rect 21539 -4740 21547 -4684
rect 21603 -4740 21627 -4684
rect 21683 -4740 21707 -4684
rect 21763 -4740 21787 -4684
rect 21843 -4740 21867 -4684
rect 21923 -4740 21947 -4684
rect 22003 -4740 22027 -4684
rect 22083 -4740 22091 -4684
rect 21539 -4775 22091 -4740
rect 21539 -4831 21547 -4775
rect 21603 -4831 21627 -4775
rect 21683 -4831 21707 -4775
rect 21763 -4831 21787 -4775
rect 21843 -4831 21867 -4775
rect 21923 -4831 21947 -4775
rect 22003 -4831 22027 -4775
rect 22083 -4831 22091 -4775
rect 21539 -4836 22091 -4831
<< metal4 >>
rect 8792 23111 9011 23325
rect 13675 15116 14100 15987
rect 8358 8037 8761 8394
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1701704242
transform -1 0 102 0 -1 4031
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1701704242
transform 0 -1 79 1 0 3302
box 0 0 1 1
use L1M1_CDNS_524688791851241  L1M1_CDNS_524688791851241_0
timestamp 1701704242
transform -1 0 17218 0 -1 1613
box -12 -6 262 400
use L1M1_CDNS_524688791851441  L1M1_CDNS_524688791851441_0
timestamp 1701704242
transform 1 0 16636 0 1 179
box -12 -6 406 616
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_0
timestamp 1701704242
transform 0 1 25486 -1 0 -2862
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_1
timestamp 1701704242
transform -1 0 8362 0 1 3523
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_2
timestamp 1701704242
transform -1 0 7551 0 1 508
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_3
timestamp 1701704242
transform -1 0 114 0 -1 4043
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_4
timestamp 1701704242
transform -1 0 17560 0 -1 -2992
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_5
timestamp 1701704242
transform 0 -1 91 1 0 3288
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_6
timestamp 1701704242
transform 0 -1 -2837 1 0 4430
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_7
timestamp 1701704242
transform 0 -1 -2757 1 0 4430
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_8
timestamp 1701704242
transform 0 -1 -3157 1 0 4438
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_9
timestamp 1701704242
transform 0 -1 -2677 1 0 4417
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_10
timestamp 1701704242
transform 0 -1 -2517 1 0 4417
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_11
timestamp 1701704242
transform 1 0 9386 0 1 3609
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_12
timestamp 1701704242
transform 1 0 8402 0 1 4083
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_13
timestamp 1701704242
transform 1 0 9169 0 1 428
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_14
timestamp 1701704242
transform 1 0 9189 0 1 3121
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_15
timestamp 1701704242
transform 1 0 10434 0 1 3438
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_16
timestamp 1701704242
transform 1 0 6324 0 1 3358
box 0 0 1 1
use M1M2_CDNS_52468879185197  M1M2_CDNS_52468879185197_0
timestamp 1701704242
transform -1 0 20935 0 1 18164
box 0 0 256 116
use M1M2_CDNS_52468879185197  M1M2_CDNS_52468879185197_1
timestamp 1701704242
transform 1 0 2023 0 1 1941
box 0 0 256 116
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_0
timestamp 1701704242
transform 1 0 22460 0 1 6184
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_1
timestamp 1701704242
transform 1 0 19341 0 1 21961
box 0 0 1 1
use M1M2_CDNS_52468879185201  M1M2_CDNS_52468879185201_0
timestamp 1701704242
transform 1 0 29204 0 1 28354
box 0 0 320 116
use M1M2_CDNS_52468879185209  M1M2_CDNS_52468879185209_0
timestamp 1701704242
transform 0 1 23423 1 0 24141
box 0 0 128 244
use M1M2_CDNS_52468879185209  M1M2_CDNS_52468879185209_1
timestamp 1701704242
transform 0 1 23423 1 0 23878
box 0 0 128 244
use M1M2_CDNS_52468879185209  M1M2_CDNS_52468879185209_2
timestamp 1701704242
transform 0 1 23423 1 0 23613
box 0 0 128 244
use M1M2_CDNS_52468879185209  M1M2_CDNS_52468879185209_3
timestamp 1701704242
transform 0 1 23423 1 0 23349
box 0 0 128 244
use M1M2_CDNS_52468879185209  M1M2_CDNS_52468879185209_4
timestamp 1701704242
transform 0 1 23423 1 0 23089
box 0 0 128 244
use M1M2_CDNS_52468879185209  M1M2_CDNS_52468879185209_5
timestamp 1701704242
transform 0 1 23423 1 0 22825
box 0 0 128 244
use M1M2_CDNS_524688791851077  M1M2_CDNS_524688791851077_0
timestamp 1701704242
transform 1 0 29204 0 1 27561
box 0 0 320 180
use M1M2_CDNS_524688791851175  M1M2_CDNS_524688791851175_0
timestamp 1701704242
transform 0 1 20658 1 0 24145
box 0 0 128 308
use M1M2_CDNS_524688791851175  M1M2_CDNS_524688791851175_1
timestamp 1701704242
transform 0 1 20658 1 0 23878
box 0 0 128 308
use M1M2_CDNS_524688791851175  M1M2_CDNS_524688791851175_2
timestamp 1701704242
transform 0 1 20658 1 0 23613
box 0 0 128 308
use M1M2_CDNS_524688791851175  M1M2_CDNS_524688791851175_3
timestamp 1701704242
transform 0 1 20658 1 0 23349
box 0 0 128 308
use M1M2_CDNS_524688791851175  M1M2_CDNS_524688791851175_4
timestamp 1701704242
transform 0 1 20658 1 0 23089
box 0 0 128 308
use M1M2_CDNS_524688791851175  M1M2_CDNS_524688791851175_5
timestamp 1701704242
transform 0 1 20658 1 0 22825
box 0 0 128 308
use M1M2_CDNS_524688791851175  M1M2_CDNS_524688791851175_6
timestamp 1701704242
transform 0 1 17017 1 0 1931
box 0 0 128 308
use M1M2_CDNS_524688791851432  M1M2_CDNS_524688791851432_0
timestamp 1701704242
transform 1 0 11237 0 1 2977
box 0 0 832 1012
use M1M2_CDNS_524688791851433  M1M2_CDNS_524688791851433_0
timestamp 1701704242
transform 1 0 12730 0 1 2977
box 0 0 512 1140
use M1M2_CDNS_524688791851434  M1M2_CDNS_524688791851434_0
timestamp 1701704242
transform 1 0 16121 0 1 1420
box 0 0 512 372
use M1M2_CDNS_524688791851434  M1M2_CDNS_524688791851434_1
timestamp 1701704242
transform 1 0 16121 0 1 249
box 0 0 512 372
use M1M2_CDNS_524688791851435  M1M2_CDNS_524688791851435_0
timestamp 1701704242
transform 1 0 12730 0 -1 2709
box 0 0 512 564
use M1M2_CDNS_524688791851436  M1M2_CDNS_524688791851436_0
timestamp 1701704242
transform 1 0 10975 0 -1 2709
box 0 0 1088 564
use M1M2_CDNS_524688791851437  M1M2_CDNS_524688791851437_0
timestamp 1701704242
transform 1 0 10975 0 1 1218
box 0 0 1088 628
use M1M2_CDNS_524688791851438  M1M2_CDNS_524688791851438_0
timestamp 1701704242
transform 1 0 12730 0 1 1218
box 0 0 512 628
use M1M2_CDNS_524688791851439  M1M2_CDNS_524688791851439_0
timestamp 1701704242
transform 1 0 3602 0 1 21706
box 0 0 1920 116
use M1M2_CDNS_524688791851440  M1M2_CDNS_524688791851440_0
timestamp 1701704242
transform -1 0 6562 0 1 22492
box 0 0 1536 116
use M3M4_CDNS_524688791851431  M3M4_CDNS_524688791851431_0
timestamp 1701704242
transform 1 0 14145 0 1 21085
box -1 0 225 476
use nfet_CDNS_524688791851442  nfet_CDNS_524688791851442_0
timestamp 1701704242
transform 1 0 10748 0 1 751
box -79 -26 4079 110
use nfet_CDNS_524688791851442  nfet_CDNS_524688791851442_1
timestamp 1701704242
transform 1 0 10748 0 1 543
box -79 -26 4079 110
use nfet_CDNS_524688791851442  nfet_CDNS_524688791851442_2
timestamp 1701704242
transform 1 0 6567 0 1 543
box -79 -26 4079 110
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_0
timestamp 1701704242
transform 0 -1 95 -1 0 3356
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_1
timestamp 1701704242
transform 0 -1 95 1 0 4060
box 0 0 1 1
use PYres_CDNS_524688791851665  PYres_CDNS_524688791851665_0
timestamp 1701704242
transform 0 -1 112 1 0 3408
box -50 0 650 100
use sky130_fd_io__sio_hotswap  sky130_fd_io__sio_hotswap_0
timestamp 1701704242
transform 1 0 2449 0 1 17331
box -232 -2471 30116 15428
use sky130_fd_io__sio_odrvr_nonreg  sky130_fd_io__sio_odrvr_nonreg_0
timestamp 1701704242
transform 1 0 221 0 1 1066
box -3430 -3054 19072 25952
use sky130_fd_io__sio_pudrvr_reg  sky130_fd_io__sio_pudrvr_reg_0
timestamp 1701704242
transform 1 0 17264 0 1 -2889
box -16995 -5965 16495 36653
<< labels >>
flabel comment s 13078 3478 13078 3478 0 FreeSans 500 0 0 0 vnb
flabel comment s 11470 3411 11470 3411 0 FreeSans 500 0 0 0 vnb
flabel comment s 395 2932 395 2932 0 FreeSans 500 0 0 0 vcc_io
flabel comment s 2505 2938 2505 2938 0 FreeSans 500 0 0 0 vcc_io
flabel comment s 4696 2952 4696 2952 0 FreeSans 500 0 0 0 vcc_io
flabel comment s 7423 3133 7423 3133 0 FreeSans 500 0 0 0 vcc_io
flabel comment s 9916 3240 9916 3240 0 FreeSans 500 0 0 0 vcc_io
flabel comment s 8830 3113 8830 3113 0 FreeSans 500 0 0 0 vgnd_io
flabel comment s 5728 2905 5728 2905 0 FreeSans 500 0 0 0 vgnd_io
flabel comment s 3457 2871 3457 2871 0 FreeSans 500 0 0 0 vgnd_io
flabel comment s 5304 31872 5304 31872 0 FreeSans 300 90 0 0 1250ohm
flabel comment s 7781 888 7781 888 0 FreeSans 440 0 0 0 condiode
flabel metal1 s 17162 -2301 17229 -2249 3 FreeSans 200 0 0 0 slow_h_n
port 4 nsew
flabel metal1 s 17162 -2393 17231 -2341 3 FreeSans 200 0 0 0 vreg_en_h
port 5 nsew
flabel metal1 s 17162 -2533 17259 -2481 3 FreeSans 200 0 0 0 puen_reg_h
port 6 nsew
flabel metal1 s 15813 5198 15868 5252 7 FreeSans 400 0 0 0 pd_h<4>
port 3 nsew
flabel metal1 s 17162 -2613 17259 -2561 3 FreeSans 200 0 0 0 drvhi_h
port 7 nsew
flabel metal1 s 16911 21955 16938 22007 0 FreeSans 600 270 0 0 p2g
port 2 nsew
flabel metal4 s 13675 15116 14100 15987 0 FreeSans 200 0 0 0 pad
port 8 nsew
flabel metal4 s 8792 23111 9011 23325 0 FreeSans 200 0 0 0 pad
port 8 nsew
flabel metal4 s 8358 8037 8761 8394 0 FreeSans 200 0 0 0 pad
port 8 nsew
flabel metal3 s 1135 19652 1354 19866 0 FreeSans 200 0 0 0 pad
port 8 nsew
flabel metal2 s -2569 4464 -2517 4498 3 FreeSans 200 90 0 0 pu_h_n<2>
port 9 nsew
flabel metal2 s 16633 4464 16691 4521 3 FreeSans 200 90 0 0 pd_h<3>
port 10 nsew
flabel metal2 s 6327 4088 6379 4122 3 FreeSans 200 90 0 0 pd_h<1>
port 11 nsew
flabel metal2 s 8450 4092 8502 4126 3 FreeSans 200 90 0 0 pd_h<0>
port 12 nsew
flabel metal2 s 16786 4464 16844 4522 3 FreeSans 200 90 0 0 tie_lo_esd
port 13 nsew
flabel metal2 s 31290 14732 31434 14867 0 FreeSans 200 0 0 0 vpwr_ka
port 14 nsew
flabel metal2 s 15306 4464 15488 4538 0 FreeSans 400 0 0 0 vcc_io
port 15 nsew
flabel metal2 s 11737 4464 11919 4538 0 FreeSans 400 0 0 0 vcc_io
port 15 nsew
flabel metal2 s 9700 4464 9882 4538 0 FreeSans 400 0 0 0 vcc_io
port 15 nsew
flabel metal2 s 6330 4464 6512 4538 0 FreeSans 400 0 0 0 vcc_io
port 15 nsew
flabel metal2 s 4584 4464 4766 4538 0 FreeSans 400 0 0 0 vcc_io
port 15 nsew
flabel metal2 s 2409 4464 2591 4538 0 FreeSans 400 0 0 0 vcc_io
port 15 nsew
flabel metal2 s 17782 21612 18092 21652 0 FreeSans 200 0 0 0 vcc_io
port 15 nsew
flabel metal2 s 5416 4464 5638 4538 0 FreeSans 400 0 0 0 vgnd_io
port 16 nsew
flabel metal2 s 9024 4464 9246 4538 0 FreeSans 400 0 0 0 vgnd_io
port 16 nsew
flabel metal2 s 11022 4464 11243 4538 0 FreeSans 400 0 0 0 vgnd_io
port 16 nsew
flabel metal2 s 14436 4464 14658 4538 0 FreeSans 400 0 0 0 vgnd_io
port 16 nsew
flabel metal2 s 16190 4464 16412 4538 0 FreeSans 400 0 0 0 vgnd_io
port 16 nsew
flabel metal2 s 3612 4464 3834 4538 0 FreeSans 400 0 0 0 vgnd_io
port 16 nsew
flabel metal2 s 17012 4464 17332 4529 0 FreeSans 200 0 0 0 pad
port 8 nsew
flabel metal2 s 860 18818 860 18818 0 FreeSans 200 90 0 0 pghs_h
flabel metal2 s 775 20359 775 20359 0 FreeSans 200 90 0 0 pug_h<0>
flabel metal2 s 1262 20297 1262 20297 0 FreeSans 200 90 0 0 pug_h<1>
flabel metal2 s 1418 21055 1418 21055 0 FreeSans 200 90 0 0 pug_h<2>
flabel metal2 s 1576 21402 1576 21402 0 FreeSans 200 90 0 0 pug_h<3>
flabel metal2 s 24986 26640 24986 26640 0 FreeSans 200 180 0 0 pug_h<4>
flabel metal2 s 24981 26557 24981 26557 0 FreeSans 200 0 0 0 pug_h<5>
flabel metal2 s 836 6549 836 6549 0 FreeSans 200 90 0 0 tie_hi
flabel metal2 s 19373 26060 19373 26060 0 FreeSans 200 90 0 0 vpb_drvr
flabel metal2 s 22527 5384 22527 5384 0 FreeSans 200 90 0 0 vref_int
flabel metal2 s 20284 14889 20506 14963 0 FreeSans 400 0 0 0 vgnd_io
port 16 nsew
flabel metal2 s 15853 4464 15911 4521 3 FreeSans 200 90 0 0 pd_h<2>
port 17 nsew
flabel metal2 s -2409 4464 -2357 4498 3 FreeSans 200 90 0 0 pu_h_n<3>
port 18 nsew
flabel metal2 s -2729 4464 -2677 4498 3 FreeSans 200 90 0 0 pu_h_n<1>
port 19 nsew
flabel metal2 s 31700 14727 31828 14867 7 FreeSans 200 90 0 0 refleak_bias
port 20 nsew
flabel metal2 s 31514 14727 31642 14867 7 FreeSans 200 90 0 0 voutref
port 21 nsew
flabel metal2 s -3209 4464 -3157 4498 3 FreeSans 200 90 0 0 pu_h_n<0>
port 22 nsew
<< properties >>
string GDS_END 100306206
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 98937186
string path 545.375 -120.900 545.375 -105.650 
<< end >>
