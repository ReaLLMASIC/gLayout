magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< pwell >>
rect -79 -26 4079 110
<< mvnmos >>
rect 0 0 4000 84
<< mvndiff >>
rect -53 46 0 84
rect -53 12 -45 46
rect -11 12 0 46
rect -53 0 0 12
rect 4000 46 4053 84
rect 4000 12 4011 46
rect 4045 12 4053 46
rect 4000 0 4053 12
<< mvndiffc >>
rect -45 12 -11 46
rect 4011 12 4045 46
<< poly >>
rect 0 84 4000 110
rect 0 -26 4000 0
<< locali >>
rect -45 46 -11 62
rect -45 -4 -11 12
rect 4011 46 4045 62
<< viali >>
rect 4011 12 4045 30
rect 4011 -4 4045 12
<< metal1 >>
rect 4005 30 4051 42
rect 4005 -4 4011 30
rect 4045 -4 4051 30
rect 4005 -16 4051 -4
use hvDFL1sd_CDNS_52468879185349  hvDFL1sd_CDNS_52468879185349_0
timestamp 1701704242
transform -1 0 0 0 1 0
box 0 0 1 1
use hvDFM1sd_CDNS_52468879185145  hvDFM1sd_CDNS_52468879185145_0
timestamp 1701704242
transform 1 0 4000 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s -28 29 -28 29 0 FreeSans 300 0 0 0 S
flabel comment s 4028 13 4028 13 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 85979046
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85978156
<< end >>
