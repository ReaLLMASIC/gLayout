magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -38 261 1602 582
<< pwell >>
rect 1 21 1545 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 247 47 277 177
rect 331 47 361 177
rect 519 47 549 177
rect 603 47 633 177
rect 691 47 721 177
rect 775 47 805 177
rect 859 47 889 177
rect 943 47 973 177
rect 1031 47 1061 177
rect 1183 47 1213 177
rect 1307 47 1337 177
rect 1391 47 1421 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 247 297 277 497
rect 331 297 361 497
rect 415 297 445 497
rect 503 297 533 497
rect 691 297 721 497
rect 775 297 805 497
rect 859 297 889 497
rect 943 297 973 497
rect 1139 297 1169 497
rect 1223 297 1253 497
rect 1307 297 1337 497
rect 1391 297 1421 497
<< ndiff >>
rect 27 93 79 177
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 161 163 177
rect 109 127 119 161
rect 153 127 163 161
rect 109 93 163 127
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 93 247 177
rect 193 59 203 93
rect 237 59 247 93
rect 193 47 247 59
rect 277 161 331 177
rect 277 127 287 161
rect 321 127 331 161
rect 277 93 331 127
rect 277 59 287 93
rect 321 59 331 93
rect 277 47 331 59
rect 361 161 413 177
rect 361 127 371 161
rect 405 127 413 161
rect 361 93 413 127
rect 361 59 371 93
rect 405 59 413 93
rect 361 47 413 59
rect 467 93 519 177
rect 467 59 475 93
rect 509 59 519 93
rect 467 47 519 59
rect 549 161 603 177
rect 549 127 559 161
rect 593 127 603 161
rect 549 47 603 127
rect 633 161 691 177
rect 633 127 647 161
rect 681 127 691 161
rect 633 93 691 127
rect 633 59 647 93
rect 681 59 691 93
rect 633 47 691 59
rect 721 93 775 177
rect 721 59 731 93
rect 765 59 775 93
rect 721 47 775 59
rect 805 169 859 177
rect 805 135 815 169
rect 849 135 859 169
rect 805 101 859 135
rect 805 67 815 101
rect 849 67 859 101
rect 805 47 859 67
rect 889 93 943 177
rect 889 59 899 93
rect 933 59 943 93
rect 889 47 943 59
rect 973 169 1031 177
rect 973 135 983 169
rect 1017 135 1031 169
rect 973 101 1031 135
rect 973 67 983 101
rect 1017 67 1031 101
rect 973 47 1031 67
rect 1061 93 1183 177
rect 1061 59 1071 93
rect 1105 59 1139 93
rect 1173 59 1183 93
rect 1061 47 1183 59
rect 1213 169 1307 177
rect 1213 135 1248 169
rect 1282 135 1307 169
rect 1213 101 1307 135
rect 1213 67 1248 101
rect 1282 67 1307 101
rect 1213 47 1307 67
rect 1337 93 1391 177
rect 1337 59 1347 93
rect 1381 59 1391 93
rect 1337 47 1391 59
rect 1421 169 1519 177
rect 1421 135 1469 169
rect 1503 135 1519 169
rect 1421 101 1519 135
rect 1421 67 1469 101
rect 1503 67 1519 101
rect 1421 47 1519 67
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 417 79 451
rect 27 383 35 417
rect 69 383 79 417
rect 27 297 79 383
rect 109 485 163 497
rect 109 451 119 485
rect 153 451 163 485
rect 109 417 163 451
rect 109 383 119 417
rect 153 383 163 417
rect 109 349 163 383
rect 109 315 119 349
rect 153 315 163 349
rect 109 297 163 315
rect 193 485 247 497
rect 193 451 203 485
rect 237 451 247 485
rect 193 417 247 451
rect 193 383 203 417
rect 237 383 247 417
rect 193 297 247 383
rect 277 485 331 497
rect 277 451 287 485
rect 321 451 331 485
rect 277 417 331 451
rect 277 383 287 417
rect 321 383 331 417
rect 277 349 331 383
rect 277 315 287 349
rect 321 315 331 349
rect 277 297 331 315
rect 361 485 415 497
rect 361 451 371 485
rect 405 451 415 485
rect 361 417 415 451
rect 361 383 371 417
rect 405 383 415 417
rect 361 349 415 383
rect 361 315 371 349
rect 405 315 415 349
rect 361 297 415 315
rect 445 485 503 497
rect 445 451 459 485
rect 493 451 503 485
rect 445 417 503 451
rect 445 383 459 417
rect 493 383 503 417
rect 445 349 503 383
rect 445 315 459 349
rect 493 315 503 349
rect 445 297 503 315
rect 533 485 585 497
rect 533 451 543 485
rect 577 451 585 485
rect 533 417 585 451
rect 533 383 543 417
rect 577 383 585 417
rect 533 297 585 383
rect 639 485 691 497
rect 639 451 647 485
rect 681 451 691 485
rect 639 417 691 451
rect 639 383 647 417
rect 681 383 691 417
rect 639 297 691 383
rect 721 407 775 497
rect 721 373 731 407
rect 765 373 775 407
rect 721 339 775 373
rect 721 305 731 339
rect 765 305 775 339
rect 721 297 775 305
rect 805 475 859 497
rect 805 441 815 475
rect 849 441 859 475
rect 805 407 859 441
rect 805 373 815 407
rect 849 373 859 407
rect 805 339 859 373
rect 805 305 815 339
rect 849 305 859 339
rect 805 297 859 305
rect 889 475 943 497
rect 889 441 899 475
rect 933 441 943 475
rect 889 407 943 441
rect 889 373 899 407
rect 933 373 943 407
rect 889 297 943 373
rect 973 407 1029 497
rect 973 373 983 407
rect 1017 373 1029 407
rect 973 339 1029 373
rect 973 305 983 339
rect 1017 305 1029 339
rect 973 297 1029 305
rect 1083 407 1139 497
rect 1083 373 1095 407
rect 1129 373 1139 407
rect 1083 339 1139 373
rect 1083 305 1095 339
rect 1129 305 1139 339
rect 1083 297 1139 305
rect 1169 475 1223 497
rect 1169 441 1179 475
rect 1213 441 1223 475
rect 1169 407 1223 441
rect 1169 373 1179 407
rect 1213 373 1223 407
rect 1169 297 1223 373
rect 1253 475 1307 497
rect 1253 441 1263 475
rect 1297 441 1307 475
rect 1253 407 1307 441
rect 1253 373 1263 407
rect 1297 373 1307 407
rect 1253 339 1307 373
rect 1253 305 1263 339
rect 1297 305 1307 339
rect 1253 297 1307 305
rect 1337 475 1391 497
rect 1337 441 1347 475
rect 1381 441 1391 475
rect 1337 407 1391 441
rect 1337 373 1347 407
rect 1381 373 1391 407
rect 1337 297 1391 373
rect 1421 475 1519 497
rect 1421 441 1469 475
rect 1503 441 1519 475
rect 1421 407 1519 441
rect 1421 373 1469 407
rect 1503 373 1519 407
rect 1421 339 1519 373
rect 1421 305 1469 339
rect 1503 305 1519 339
rect 1421 297 1519 305
<< ndiffc >>
rect 35 59 69 93
rect 119 127 153 161
rect 119 59 153 93
rect 203 59 237 93
rect 287 127 321 161
rect 287 59 321 93
rect 371 127 405 161
rect 371 59 405 93
rect 475 59 509 93
rect 559 127 593 161
rect 647 127 681 161
rect 647 59 681 93
rect 731 59 765 93
rect 815 135 849 169
rect 815 67 849 101
rect 899 59 933 93
rect 983 135 1017 169
rect 983 67 1017 101
rect 1071 59 1105 93
rect 1139 59 1173 93
rect 1248 135 1282 169
rect 1248 67 1282 101
rect 1347 59 1381 93
rect 1469 135 1503 169
rect 1469 67 1503 101
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 119 451 153 485
rect 119 383 153 417
rect 119 315 153 349
rect 203 451 237 485
rect 203 383 237 417
rect 287 451 321 485
rect 287 383 321 417
rect 287 315 321 349
rect 371 451 405 485
rect 371 383 405 417
rect 371 315 405 349
rect 459 451 493 485
rect 459 383 493 417
rect 459 315 493 349
rect 543 451 577 485
rect 543 383 577 417
rect 647 451 681 485
rect 647 383 681 417
rect 731 373 765 407
rect 731 305 765 339
rect 815 441 849 475
rect 815 373 849 407
rect 815 305 849 339
rect 899 441 933 475
rect 899 373 933 407
rect 983 373 1017 407
rect 983 305 1017 339
rect 1095 373 1129 407
rect 1095 305 1129 339
rect 1179 441 1213 475
rect 1179 373 1213 407
rect 1263 441 1297 475
rect 1263 373 1297 407
rect 1263 305 1297 339
rect 1347 441 1381 475
rect 1347 373 1381 407
rect 1469 441 1503 475
rect 1469 373 1503 407
rect 1469 305 1503 339
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 247 497 277 523
rect 331 497 361 523
rect 415 497 445 523
rect 503 497 533 523
rect 691 497 721 523
rect 775 497 805 523
rect 859 497 889 523
rect 943 497 973 523
rect 1139 497 1169 523
rect 1223 497 1253 523
rect 1307 497 1337 523
rect 1391 497 1421 523
rect 79 259 109 297
rect 163 259 193 297
rect 247 259 277 297
rect 331 259 361 297
rect 79 249 361 259
rect 79 215 119 249
rect 153 215 203 249
rect 237 215 288 249
rect 322 215 361 249
rect 79 205 361 215
rect 415 259 445 297
rect 503 259 533 297
rect 691 259 721 297
rect 775 259 805 297
rect 415 249 633 259
rect 415 215 583 249
rect 617 215 633 249
rect 415 205 633 215
rect 79 177 109 205
rect 163 177 193 205
rect 247 177 277 205
rect 331 177 361 205
rect 519 177 549 205
rect 603 177 633 205
rect 691 249 805 259
rect 691 215 731 249
rect 765 215 805 249
rect 691 205 805 215
rect 691 177 721 205
rect 775 177 805 205
rect 859 259 889 297
rect 943 259 973 297
rect 1139 259 1169 297
rect 1223 259 1253 297
rect 1307 259 1337 297
rect 1391 259 1421 297
rect 859 249 973 259
rect 859 215 899 249
rect 933 215 973 249
rect 859 205 973 215
rect 1030 249 1262 259
rect 1030 215 1046 249
rect 1080 215 1133 249
rect 1167 215 1212 249
rect 1246 215 1262 249
rect 1030 205 1262 215
rect 1307 249 1496 259
rect 1307 215 1350 249
rect 1384 215 1446 249
rect 1480 215 1496 249
rect 1307 205 1496 215
rect 859 177 889 205
rect 943 177 973 205
rect 1031 177 1061 205
rect 1183 177 1213 205
rect 1307 177 1337 205
rect 1391 177 1421 205
rect 79 21 109 47
rect 163 21 193 47
rect 247 21 277 47
rect 331 21 361 47
rect 519 21 549 47
rect 603 21 633 47
rect 691 21 721 47
rect 775 21 805 47
rect 859 21 889 47
rect 943 21 973 47
rect 1031 21 1061 47
rect 1183 21 1213 47
rect 1307 21 1337 47
rect 1391 21 1421 47
<< polycont >>
rect 119 215 153 249
rect 203 215 237 249
rect 288 215 322 249
rect 583 215 617 249
rect 731 215 765 249
rect 899 215 933 249
rect 1046 215 1080 249
rect 1133 215 1167 249
rect 1212 215 1246 249
rect 1350 215 1384 249
rect 1446 215 1480 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 17 485 69 527
rect 17 451 35 485
rect 17 417 69 451
rect 17 383 35 417
rect 17 367 69 383
rect 103 485 169 493
rect 103 451 119 485
rect 153 451 169 485
rect 103 417 169 451
rect 103 383 119 417
rect 153 383 169 417
rect 103 349 169 383
rect 203 485 237 527
rect 203 417 237 451
rect 203 367 237 383
rect 271 485 337 493
rect 271 451 287 485
rect 321 451 337 485
rect 271 417 337 451
rect 271 383 287 417
rect 321 383 337 417
rect 103 333 119 349
rect 17 315 119 333
rect 153 333 169 349
rect 271 349 337 383
rect 271 333 287 349
rect 153 315 287 333
rect 321 315 337 349
rect 17 293 337 315
rect 371 485 405 527
rect 371 417 405 451
rect 371 349 405 383
rect 371 293 405 315
rect 439 485 509 493
rect 439 451 459 485
rect 493 451 509 485
rect 439 417 509 451
rect 439 383 459 417
rect 493 383 509 417
rect 439 349 509 383
rect 543 485 593 527
rect 577 451 593 485
rect 543 417 593 451
rect 577 383 593 417
rect 543 367 593 383
rect 627 485 865 493
rect 627 451 647 485
rect 681 475 865 485
rect 681 459 815 475
rect 627 417 681 451
rect 799 441 815 459
rect 849 441 865 475
rect 627 383 647 417
rect 627 367 681 383
rect 715 407 765 425
rect 715 373 731 407
rect 439 315 459 349
rect 493 323 509 349
rect 715 339 765 373
rect 715 323 731 339
rect 493 315 731 323
rect 439 305 731 315
rect 17 181 69 293
rect 439 289 765 305
rect 799 407 865 441
rect 799 373 815 407
rect 849 373 865 407
rect 799 339 865 373
rect 899 475 1229 493
rect 933 459 1179 475
rect 899 407 933 441
rect 1163 441 1179 459
rect 1213 441 1229 475
rect 899 357 933 373
rect 967 407 1033 423
rect 967 373 983 407
rect 1017 373 1033 407
rect 799 305 815 339
rect 849 323 865 339
rect 967 339 1033 373
rect 967 323 983 339
rect 849 305 983 323
rect 1017 305 1033 339
rect 799 289 1033 305
rect 1079 407 1129 423
rect 1079 373 1095 407
rect 1079 339 1129 373
rect 1163 407 1229 441
rect 1163 373 1179 407
rect 1213 373 1229 407
rect 1163 357 1229 373
rect 1263 475 1297 491
rect 1263 407 1297 441
rect 1079 305 1095 339
rect 1263 339 1297 373
rect 1331 475 1397 527
rect 1331 441 1347 475
rect 1381 441 1397 475
rect 1331 407 1397 441
rect 1331 373 1347 407
rect 1381 373 1397 407
rect 1331 357 1397 373
rect 1453 475 1519 493
rect 1453 441 1469 475
rect 1503 441 1519 475
rect 1453 407 1519 441
rect 1453 373 1469 407
rect 1503 373 1519 407
rect 1129 305 1263 323
rect 1453 339 1519 373
rect 1453 323 1469 339
rect 1297 305 1469 323
rect 1503 305 1519 339
rect 1079 289 1519 305
rect 439 259 509 289
rect 103 249 509 259
rect 567 249 633 255
rect 103 215 119 249
rect 153 215 203 249
rect 237 215 288 249
rect 322 215 533 249
rect 567 215 583 249
rect 617 215 633 249
rect 682 249 808 255
rect 682 215 731 249
rect 765 215 808 249
rect 866 249 992 255
rect 866 215 899 249
rect 933 215 992 249
rect 1030 249 1272 255
rect 1030 215 1046 249
rect 1080 215 1133 249
rect 1167 215 1212 249
rect 1246 215 1272 249
rect 1330 249 1547 255
rect 1330 215 1350 249
rect 1384 215 1446 249
rect 1480 215 1547 249
rect 459 181 533 215
rect 17 161 337 181
rect 17 143 119 161
rect 103 127 119 143
rect 153 143 287 161
rect 153 127 169 143
rect 17 93 69 109
rect 17 59 35 93
rect 17 17 69 59
rect 103 93 169 127
rect 271 127 287 143
rect 321 127 337 161
rect 103 59 119 93
rect 153 59 169 93
rect 103 51 169 59
rect 203 93 237 109
rect 203 17 237 59
rect 271 93 337 127
rect 271 59 287 93
rect 321 59 337 93
rect 271 51 337 59
rect 371 161 421 177
rect 405 127 421 161
rect 459 161 609 181
rect 459 127 559 161
rect 593 127 609 161
rect 647 169 1519 181
rect 647 161 815 169
rect 681 147 815 161
rect 681 127 697 147
rect 371 93 421 127
rect 647 93 697 127
rect 849 147 983 169
rect 405 59 421 93
rect 371 17 421 59
rect 459 59 475 93
rect 509 59 647 93
rect 681 59 697 93
rect 459 51 697 59
rect 731 93 775 109
rect 765 59 775 93
rect 731 17 775 59
rect 815 101 849 135
rect 1017 147 1248 169
rect 815 51 849 67
rect 889 93 943 109
rect 889 59 899 93
rect 933 59 943 93
rect 889 17 943 59
rect 983 101 1017 135
rect 1282 147 1469 169
rect 983 51 1017 67
rect 1061 93 1183 109
rect 1061 59 1071 93
rect 1105 59 1139 93
rect 1173 59 1183 93
rect 1061 17 1183 59
rect 1248 101 1282 135
rect 1453 135 1469 147
rect 1503 135 1519 169
rect 1248 51 1282 67
rect 1337 93 1391 109
rect 1337 59 1347 93
rect 1381 59 1391 93
rect 1337 17 1391 59
rect 1453 101 1519 135
rect 1453 67 1469 101
rect 1503 67 1519 101
rect 1453 51 1519 67
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
<< metal1 >>
rect 0 561 1564 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 0 496 1564 527
rect 0 17 1564 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
rect 0 -48 1564 -17
<< labels >>
flabel locali s 1510 221 1544 255 0 FreeSans 250 0 0 0 A1
port 1 nsew signal input
flabel locali s 1422 221 1456 255 0 FreeSans 250 0 0 0 A1
port 1 nsew signal input
flabel locali s 1330 221 1364 255 0 FreeSans 250 0 0 0 A1
port 1 nsew signal input
flabel locali s 1238 221 1272 255 0 FreeSans 250 0 0 0 A2
port 2 nsew signal input
flabel locali s 1146 221 1180 255 0 FreeSans 250 0 0 0 A2
port 2 nsew signal input
flabel locali s 1054 221 1088 255 0 FreeSans 250 0 0 0 A2
port 2 nsew signal input
flabel locali s 958 221 992 255 0 FreeSans 250 0 0 0 A3
port 3 nsew signal input
flabel locali s 866 221 900 255 0 FreeSans 250 0 0 0 A3
port 3 nsew signal input
flabel locali s 774 221 808 255 0 FreeSans 250 0 0 0 A4
port 4 nsew signal input
flabel locali s 682 221 716 255 0 FreeSans 250 0 0 0 A4
port 4 nsew signal input
flabel locali s 586 221 620 255 0 FreeSans 250 0 0 0 B1
port 5 nsew signal input
flabel locali s 30 289 64 323 0 FreeSans 250 0 0 0 X
port 10 nsew signal output
flabel locali s 30 221 64 255 0 FreeSans 250 0 0 0 X
port 10 nsew signal output
flabel locali s 30 153 64 187 0 FreeSans 250 0 0 0 X
port 10 nsew signal output
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 o41a_4
rlabel metal1 s 0 -48 1564 48 1 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1564 592 1 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1564 544
string GDS_END 712108
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 699004
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 7.820 0.000 
<< end >>
