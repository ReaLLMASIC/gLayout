magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< poly >>
rect -50 50 0 66
rect -50 16 -34 50
rect -50 0 0 16
rect 9412 50 9462 66
rect 9446 16 9462 50
rect 9412 0 9462 16
<< polycont >>
rect -34 16 0 50
rect 9412 16 9446 50
<< npolyres >>
rect 0 0 9412 66
<< locali >>
rect -34 50 0 66
rect -34 0 0 16
rect 9412 50 9446 66
rect 9412 0 9446 16
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_0
timestamp 1701704242
transform 1 0 9396 0 1 0
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_1
timestamp 1701704242
transform 1 0 -50 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 98008728
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 98008248
<< end >>
