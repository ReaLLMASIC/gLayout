magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -92 -36 125 636
<< pmos >>
rect 0 0 36 600
<< pdiff >>
rect -50 0 0 600
rect 36 0 86 600
<< poly >>
rect 0 600 36 626
rect 0 -26 36 0
<< locali >>
rect -45 -4 -11 538
rect 47 -4 81 538
use DFL1sd2_CDNS_5246887918535  DFL1sd2_CDNS_5246887918535_0
timestamp 1701704242
transform -1 0 0 0 1 0
box -36 -36 92 636
use DFL1sd_CDNS_5246887918534  DFL1sd_CDNS_5246887918534_0
timestamp 1701704242
transform 1 0 36 0 1 0
box -36 -36 89 636
<< labels >>
flabel comment s -28 267 -28 267 0 FreeSans 300 0 0 0 S
flabel comment s 64 267 64 267 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 79607820
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 79606934
<< end >>
