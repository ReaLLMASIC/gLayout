magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< pwell >>
rect -76 -26 256 2026
<< mvnnmos >>
rect 0 0 180 2000
<< mvndiff >>
rect -50 0 0 2000
rect 180 0 230 2000
<< poly >>
rect 0 2000 180 2052
rect 0 -52 180 0
<< locali >>
rect -45 -4 -11 1966
rect 191 -4 225 1966
use hvDFL1sd2_CDNS_52468879185991  hvDFL1sd2_CDNS_52468879185991_0
timestamp 1701704242
transform -1 0 0 0 1 0
box -26 -26 82 2026
use hvDFL1sd2_CDNS_52468879185991  hvDFL1sd2_CDNS_52468879185991_1
timestamp 1701704242
transform 1 0 180 0 1 0
box -26 -26 82 2026
<< labels >>
flabel comment s -28 981 -28 981 0 FreeSans 300 0 0 0 S
flabel comment s 208 981 208 981 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 86888270
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86887312
<< end >>
