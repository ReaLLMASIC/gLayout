magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< pwell >>
rect -76 -26 256 2026
<< mvnnmos >>
rect 0 0 180 2000
<< mvndiff >>
rect -50 0 0 2000
rect 180 0 230 2000
<< poly >>
rect 0 2000 180 2026
rect 0 -26 180 0
<< metal1 >>
rect -51 -16 -5 1986
rect 185 -16 231 1986
use DFM1sd_CDNS_524688791851117  DFM1sd_CDNS_524688791851117_0
timestamp 1701704242
transform -1 0 0 0 1 0
box -26 -26 79 2026
use DFM1sd_CDNS_524688791851117  DFM1sd_CDNS_524688791851117_1
timestamp 1701704242
transform 1 0 180 0 1 0
box -26 -26 79 2026
<< labels >>
flabel comment s -28 985 -28 985 0 FreeSans 300 0 0 0 S
flabel comment s 208 985 208 985 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 86364604
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86363650
<< end >>
