magic
tech sky130A
timestamp 1701704242
<< properties >>
string GDS_END 4737978
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_START 4737654
<< end >>
