magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 39 21 582 157
rect 39 17 63 21
rect 29 -17 63 17
<< locali >>
rect 72 365 157 493
rect 17 146 87 331
rect 121 177 157 365
rect 191 211 265 472
rect 299 211 369 347
rect 471 280 525 347
rect 407 214 525 280
rect 121 127 408 177
rect 471 132 525 214
rect 559 130 627 347
rect 157 123 408 127
rect 157 51 208 123
rect 342 56 408 123
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 308 417 374 493
rect 408 451 474 527
rect 508 417 574 493
rect 308 381 574 417
rect 57 17 123 93
rect 242 17 308 89
rect 494 17 560 96
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
rlabel locali s 471 132 525 214 6 A1
port 1 nsew signal input
rlabel locali s 407 214 525 280 6 A1
port 1 nsew signal input
rlabel locali s 471 280 525 347 6 A1
port 1 nsew signal input
rlabel locali s 559 130 627 347 6 A2
port 2 nsew signal input
rlabel locali s 299 211 369 347 6 B1
port 3 nsew signal input
rlabel locali s 191 211 265 472 6 C1
port 4 nsew signal input
rlabel locali s 17 146 87 331 6 D1
port 5 nsew signal input
rlabel metal1 s 0 -48 644 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 17 8 VNB
port 7 nsew ground bidirectional
rlabel pwell s 39 17 63 21 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 39 21 582 157 6 VNB
port 7 nsew ground bidirectional
rlabel nwell s -38 261 682 582 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 496 644 592 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 342 56 408 123 6 Y
port 10 nsew signal output
rlabel locali s 157 51 208 123 6 Y
port 10 nsew signal output
rlabel locali s 157 123 408 127 6 Y
port 10 nsew signal output
rlabel locali s 121 127 408 177 6 Y
port 10 nsew signal output
rlabel locali s 121 177 157 365 6 Y
port 10 nsew signal output
rlabel locali s 72 365 157 493 6 Y
port 10 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 644 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 3771120
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3763656
<< end >>
