magic
tech sky130B
timestamp 1701704242
<< metal1 >>
rect 0 0 3 3098
rect 285 0 288 3098
<< via1 >>
rect 3 0 285 3098
<< metal2 >>
rect 0 0 3 3098
rect 285 0 288 3098
<< properties >>
string GDS_END 93774886
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 93718882
<< end >>
