magic
tech sky130B
timestamp 1701704242
<< metal1 >>
rect 0 0 3 186
rect 125 0 128 186
<< via1 >>
rect 3 0 125 186
<< metal2 >>
rect 0 0 3 186
rect 125 0 128 186
<< properties >>
string GDS_END 88148752
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 88147084
<< end >>
