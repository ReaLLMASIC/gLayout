magic
tech sky130B
timestamp 1701704242
<< metal1 >>
rect 0 0 3 26
rect 29 0 35 26
rect 61 0 67 26
rect 93 0 99 26
rect 125 0 131 26
rect 157 0 163 26
rect 189 0 195 26
rect 221 0 227 26
rect 253 0 259 26
rect 285 0 291 26
rect 317 0 323 26
rect 349 0 355 26
rect 381 0 387 26
rect 413 0 419 26
rect 445 0 451 26
rect 477 0 483 26
rect 509 0 515 26
rect 541 0 547 26
rect 573 0 579 26
rect 605 0 611 26
rect 637 0 643 26
rect 669 0 675 26
rect 701 0 707 26
rect 733 0 739 26
rect 765 0 771 26
rect 797 0 803 26
rect 829 0 835 26
rect 861 0 867 26
rect 893 0 899 26
rect 925 0 931 26
rect 957 0 963 26
rect 989 0 995 26
rect 1021 0 1027 26
rect 1053 0 1059 26
rect 1085 0 1091 26
rect 1117 0 1123 26
rect 1149 0 1155 26
rect 1181 0 1187 26
rect 1213 0 1219 26
rect 1245 0 1251 26
rect 1277 0 1283 26
rect 1309 0 1315 26
rect 1341 0 1347 26
rect 1373 0 1379 26
rect 1405 0 1411 26
rect 1437 0 1443 26
rect 1469 0 1475 26
rect 1501 0 1507 26
rect 1533 0 1539 26
rect 1565 0 1571 26
rect 1597 0 1603 26
rect 1629 0 1635 26
rect 1661 0 1667 26
rect 1693 0 1699 26
rect 1725 0 1731 26
rect 1757 0 1763 26
rect 1789 0 1795 26
rect 1821 0 1827 26
rect 1853 0 1859 26
rect 1885 0 1891 26
rect 1917 0 1923 26
rect 1949 0 1955 26
rect 1981 0 1987 26
rect 2013 0 2019 26
rect 2045 0 2051 26
rect 2077 0 2083 26
rect 2109 0 2115 26
rect 2141 0 2147 26
rect 2173 0 2179 26
rect 2205 0 2211 26
rect 2237 0 2243 26
rect 2269 0 2275 26
rect 2301 0 2307 26
rect 2333 0 2339 26
rect 2365 0 2371 26
rect 2397 0 2403 26
rect 2429 0 2435 26
rect 2461 0 2467 26
rect 2493 0 2499 26
rect 2525 0 2531 26
rect 2557 0 2563 26
rect 2589 0 2595 26
rect 2621 0 2627 26
rect 2653 0 2659 26
rect 2685 0 2691 26
rect 2717 0 2723 26
rect 2749 0 2755 26
rect 2781 0 2787 26
rect 2813 0 2819 26
rect 2845 0 2851 26
rect 2877 0 2883 26
rect 2909 0 2915 26
rect 2941 0 2947 26
rect 2973 0 2979 26
rect 3005 0 3011 26
rect 3037 0 3043 26
rect 3069 0 3075 26
rect 3101 0 3107 26
rect 3133 0 3139 26
rect 3165 0 3171 26
rect 3197 0 3203 26
rect 3229 0 3235 26
rect 3261 0 3267 26
rect 3293 0 3299 26
rect 3325 0 3331 26
rect 3357 0 3363 26
rect 3389 0 3395 26
rect 3421 0 3427 26
rect 3453 0 3459 26
rect 3485 0 3491 26
rect 3517 0 3523 26
rect 3549 0 3555 26
rect 3581 0 3587 26
rect 3613 0 3619 26
rect 3645 0 3651 26
rect 3677 0 3683 26
rect 3709 0 3715 26
rect 3741 0 3747 26
rect 3773 0 3779 26
rect 3805 0 3811 26
rect 3837 0 3843 26
rect 3869 0 3875 26
rect 3901 0 3907 26
rect 3933 0 3939 26
rect 3965 0 3971 26
rect 3997 0 4003 26
rect 4029 0 4035 26
rect 4061 0 4067 26
rect 4093 0 4099 26
rect 4125 0 4131 26
rect 4157 0 4163 26
rect 4189 0 4195 26
rect 4221 0 4227 26
rect 4253 0 4259 26
rect 4285 0 4291 26
rect 4317 0 4323 26
rect 4349 0 4355 26
rect 4381 0 4387 26
rect 4413 0 4419 26
rect 4445 0 4451 26
rect 4477 0 4483 26
rect 4509 0 4515 26
rect 4541 0 4547 26
rect 4573 0 4579 26
rect 4605 0 4611 26
rect 4637 0 4643 26
rect 4669 0 4675 26
rect 4701 0 4707 26
rect 4733 0 4739 26
rect 4765 0 4771 26
rect 4797 0 4803 26
rect 4829 0 4835 26
rect 4861 0 4867 26
rect 4893 0 4899 26
rect 4925 0 4931 26
rect 4957 0 4963 26
rect 4989 0 4995 26
rect 5021 0 5027 26
rect 5053 0 5059 26
rect 5085 0 5091 26
rect 5117 0 5123 26
rect 5149 0 5155 26
rect 5181 0 5187 26
rect 5213 0 5219 26
rect 5245 0 5251 26
rect 5277 0 5283 26
rect 5309 0 5315 26
rect 5341 0 5347 26
rect 5373 0 5379 26
rect 5405 0 5411 26
rect 5437 0 5443 26
rect 5469 0 5475 26
rect 5501 0 5507 26
rect 5533 0 5539 26
rect 5565 0 5571 26
rect 5597 0 5603 26
rect 5629 0 5635 26
rect 5661 0 5667 26
rect 5693 0 5699 26
rect 5725 0 5731 26
rect 5757 0 5763 26
rect 5789 0 5795 26
rect 5821 0 5827 26
rect 5853 0 5856 26
<< via1 >>
rect 3 0 29 26
rect 35 0 61 26
rect 67 0 93 26
rect 99 0 125 26
rect 131 0 157 26
rect 163 0 189 26
rect 195 0 221 26
rect 227 0 253 26
rect 259 0 285 26
rect 291 0 317 26
rect 323 0 349 26
rect 355 0 381 26
rect 387 0 413 26
rect 419 0 445 26
rect 451 0 477 26
rect 483 0 509 26
rect 515 0 541 26
rect 547 0 573 26
rect 579 0 605 26
rect 611 0 637 26
rect 643 0 669 26
rect 675 0 701 26
rect 707 0 733 26
rect 739 0 765 26
rect 771 0 797 26
rect 803 0 829 26
rect 835 0 861 26
rect 867 0 893 26
rect 899 0 925 26
rect 931 0 957 26
rect 963 0 989 26
rect 995 0 1021 26
rect 1027 0 1053 26
rect 1059 0 1085 26
rect 1091 0 1117 26
rect 1123 0 1149 26
rect 1155 0 1181 26
rect 1187 0 1213 26
rect 1219 0 1245 26
rect 1251 0 1277 26
rect 1283 0 1309 26
rect 1315 0 1341 26
rect 1347 0 1373 26
rect 1379 0 1405 26
rect 1411 0 1437 26
rect 1443 0 1469 26
rect 1475 0 1501 26
rect 1507 0 1533 26
rect 1539 0 1565 26
rect 1571 0 1597 26
rect 1603 0 1629 26
rect 1635 0 1661 26
rect 1667 0 1693 26
rect 1699 0 1725 26
rect 1731 0 1757 26
rect 1763 0 1789 26
rect 1795 0 1821 26
rect 1827 0 1853 26
rect 1859 0 1885 26
rect 1891 0 1917 26
rect 1923 0 1949 26
rect 1955 0 1981 26
rect 1987 0 2013 26
rect 2019 0 2045 26
rect 2051 0 2077 26
rect 2083 0 2109 26
rect 2115 0 2141 26
rect 2147 0 2173 26
rect 2179 0 2205 26
rect 2211 0 2237 26
rect 2243 0 2269 26
rect 2275 0 2301 26
rect 2307 0 2333 26
rect 2339 0 2365 26
rect 2371 0 2397 26
rect 2403 0 2429 26
rect 2435 0 2461 26
rect 2467 0 2493 26
rect 2499 0 2525 26
rect 2531 0 2557 26
rect 2563 0 2589 26
rect 2595 0 2621 26
rect 2627 0 2653 26
rect 2659 0 2685 26
rect 2691 0 2717 26
rect 2723 0 2749 26
rect 2755 0 2781 26
rect 2787 0 2813 26
rect 2819 0 2845 26
rect 2851 0 2877 26
rect 2883 0 2909 26
rect 2915 0 2941 26
rect 2947 0 2973 26
rect 2979 0 3005 26
rect 3011 0 3037 26
rect 3043 0 3069 26
rect 3075 0 3101 26
rect 3107 0 3133 26
rect 3139 0 3165 26
rect 3171 0 3197 26
rect 3203 0 3229 26
rect 3235 0 3261 26
rect 3267 0 3293 26
rect 3299 0 3325 26
rect 3331 0 3357 26
rect 3363 0 3389 26
rect 3395 0 3421 26
rect 3427 0 3453 26
rect 3459 0 3485 26
rect 3491 0 3517 26
rect 3523 0 3549 26
rect 3555 0 3581 26
rect 3587 0 3613 26
rect 3619 0 3645 26
rect 3651 0 3677 26
rect 3683 0 3709 26
rect 3715 0 3741 26
rect 3747 0 3773 26
rect 3779 0 3805 26
rect 3811 0 3837 26
rect 3843 0 3869 26
rect 3875 0 3901 26
rect 3907 0 3933 26
rect 3939 0 3965 26
rect 3971 0 3997 26
rect 4003 0 4029 26
rect 4035 0 4061 26
rect 4067 0 4093 26
rect 4099 0 4125 26
rect 4131 0 4157 26
rect 4163 0 4189 26
rect 4195 0 4221 26
rect 4227 0 4253 26
rect 4259 0 4285 26
rect 4291 0 4317 26
rect 4323 0 4349 26
rect 4355 0 4381 26
rect 4387 0 4413 26
rect 4419 0 4445 26
rect 4451 0 4477 26
rect 4483 0 4509 26
rect 4515 0 4541 26
rect 4547 0 4573 26
rect 4579 0 4605 26
rect 4611 0 4637 26
rect 4643 0 4669 26
rect 4675 0 4701 26
rect 4707 0 4733 26
rect 4739 0 4765 26
rect 4771 0 4797 26
rect 4803 0 4829 26
rect 4835 0 4861 26
rect 4867 0 4893 26
rect 4899 0 4925 26
rect 4931 0 4957 26
rect 4963 0 4989 26
rect 4995 0 5021 26
rect 5027 0 5053 26
rect 5059 0 5085 26
rect 5091 0 5117 26
rect 5123 0 5149 26
rect 5155 0 5181 26
rect 5187 0 5213 26
rect 5219 0 5245 26
rect 5251 0 5277 26
rect 5283 0 5309 26
rect 5315 0 5341 26
rect 5347 0 5373 26
rect 5379 0 5405 26
rect 5411 0 5437 26
rect 5443 0 5469 26
rect 5475 0 5501 26
rect 5507 0 5533 26
rect 5539 0 5565 26
rect 5571 0 5597 26
rect 5603 0 5629 26
rect 5635 0 5661 26
rect 5667 0 5693 26
rect 5699 0 5725 26
rect 5731 0 5757 26
rect 5763 0 5789 26
rect 5795 0 5821 26
rect 5827 0 5853 26
<< metal2 >>
rect 0 0 3 26
rect 29 0 35 26
rect 61 0 67 26
rect 93 0 99 26
rect 125 0 131 26
rect 157 0 163 26
rect 189 0 195 26
rect 221 0 227 26
rect 253 0 259 26
rect 285 0 291 26
rect 317 0 323 26
rect 349 0 355 26
rect 381 0 387 26
rect 413 0 419 26
rect 445 0 451 26
rect 477 0 483 26
rect 509 0 515 26
rect 541 0 547 26
rect 573 0 579 26
rect 605 0 611 26
rect 637 0 643 26
rect 669 0 675 26
rect 701 0 707 26
rect 733 0 739 26
rect 765 0 771 26
rect 797 0 803 26
rect 829 0 835 26
rect 861 0 867 26
rect 893 0 899 26
rect 925 0 931 26
rect 957 0 963 26
rect 989 0 995 26
rect 1021 0 1027 26
rect 1053 0 1059 26
rect 1085 0 1091 26
rect 1117 0 1123 26
rect 1149 0 1155 26
rect 1181 0 1187 26
rect 1213 0 1219 26
rect 1245 0 1251 26
rect 1277 0 1283 26
rect 1309 0 1315 26
rect 1341 0 1347 26
rect 1373 0 1379 26
rect 1405 0 1411 26
rect 1437 0 1443 26
rect 1469 0 1475 26
rect 1501 0 1507 26
rect 1533 0 1539 26
rect 1565 0 1571 26
rect 1597 0 1603 26
rect 1629 0 1635 26
rect 1661 0 1667 26
rect 1693 0 1699 26
rect 1725 0 1731 26
rect 1757 0 1763 26
rect 1789 0 1795 26
rect 1821 0 1827 26
rect 1853 0 1859 26
rect 1885 0 1891 26
rect 1917 0 1923 26
rect 1949 0 1955 26
rect 1981 0 1987 26
rect 2013 0 2019 26
rect 2045 0 2051 26
rect 2077 0 2083 26
rect 2109 0 2115 26
rect 2141 0 2147 26
rect 2173 0 2179 26
rect 2205 0 2211 26
rect 2237 0 2243 26
rect 2269 0 2275 26
rect 2301 0 2307 26
rect 2333 0 2339 26
rect 2365 0 2371 26
rect 2397 0 2403 26
rect 2429 0 2435 26
rect 2461 0 2467 26
rect 2493 0 2499 26
rect 2525 0 2531 26
rect 2557 0 2563 26
rect 2589 0 2595 26
rect 2621 0 2627 26
rect 2653 0 2659 26
rect 2685 0 2691 26
rect 2717 0 2723 26
rect 2749 0 2755 26
rect 2781 0 2787 26
rect 2813 0 2819 26
rect 2845 0 2851 26
rect 2877 0 2883 26
rect 2909 0 2915 26
rect 2941 0 2947 26
rect 2973 0 2979 26
rect 3005 0 3011 26
rect 3037 0 3043 26
rect 3069 0 3075 26
rect 3101 0 3107 26
rect 3133 0 3139 26
rect 3165 0 3171 26
rect 3197 0 3203 26
rect 3229 0 3235 26
rect 3261 0 3267 26
rect 3293 0 3299 26
rect 3325 0 3331 26
rect 3357 0 3363 26
rect 3389 0 3395 26
rect 3421 0 3427 26
rect 3453 0 3459 26
rect 3485 0 3491 26
rect 3517 0 3523 26
rect 3549 0 3555 26
rect 3581 0 3587 26
rect 3613 0 3619 26
rect 3645 0 3651 26
rect 3677 0 3683 26
rect 3709 0 3715 26
rect 3741 0 3747 26
rect 3773 0 3779 26
rect 3805 0 3811 26
rect 3837 0 3843 26
rect 3869 0 3875 26
rect 3901 0 3907 26
rect 3933 0 3939 26
rect 3965 0 3971 26
rect 3997 0 4003 26
rect 4029 0 4035 26
rect 4061 0 4067 26
rect 4093 0 4099 26
rect 4125 0 4131 26
rect 4157 0 4163 26
rect 4189 0 4195 26
rect 4221 0 4227 26
rect 4253 0 4259 26
rect 4285 0 4291 26
rect 4317 0 4323 26
rect 4349 0 4355 26
rect 4381 0 4387 26
rect 4413 0 4419 26
rect 4445 0 4451 26
rect 4477 0 4483 26
rect 4509 0 4515 26
rect 4541 0 4547 26
rect 4573 0 4579 26
rect 4605 0 4611 26
rect 4637 0 4643 26
rect 4669 0 4675 26
rect 4701 0 4707 26
rect 4733 0 4739 26
rect 4765 0 4771 26
rect 4797 0 4803 26
rect 4829 0 4835 26
rect 4861 0 4867 26
rect 4893 0 4899 26
rect 4925 0 4931 26
rect 4957 0 4963 26
rect 4989 0 4995 26
rect 5021 0 5027 26
rect 5053 0 5059 26
rect 5085 0 5091 26
rect 5117 0 5123 26
rect 5149 0 5155 26
rect 5181 0 5187 26
rect 5213 0 5219 26
rect 5245 0 5251 26
rect 5277 0 5283 26
rect 5309 0 5315 26
rect 5341 0 5347 26
rect 5373 0 5379 26
rect 5405 0 5411 26
rect 5437 0 5443 26
rect 5469 0 5475 26
rect 5501 0 5507 26
rect 5533 0 5539 26
rect 5565 0 5571 26
rect 5597 0 5603 26
rect 5629 0 5635 26
rect 5661 0 5667 26
rect 5693 0 5699 26
rect 5725 0 5731 26
rect 5757 0 5763 26
rect 5789 0 5795 26
rect 5821 0 5827 26
rect 5853 0 5856 26
<< properties >>
string GDS_END 78988224
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 78976380
<< end >>
