magic
tech sky130B
timestamp 1701704242
<< metal1 >>
rect 0 0 3 122
rect 253 0 256 122
<< via1 >>
rect 3 0 253 122
<< metal2 >>
rect 0 0 3 122
rect 253 0 256 122
<< properties >>
string GDS_END 88147026
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 88144846
<< end >>
