magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -119 -66 531 1466
<< mvpmos >>
rect 0 0 100 1400
rect 156 0 256 1400
rect 312 0 412 1400
<< mvpdiff >>
rect -50 0 0 1400
rect 412 0 462 1400
<< poly >>
rect 0 1400 100 1452
rect 0 -52 100 0
rect 156 1400 256 1452
rect 156 -52 256 0
rect 312 1400 412 1452
rect 312 -52 412 0
<< locali >>
rect -45 -4 -11 1354
rect 111 -4 145 1354
rect 267 -4 301 1354
rect 423 -4 457 1354
use DFL1sd_CDNS_52468879185620  DFL1sd_CDNS_52468879185620_0
timestamp 1701704242
transform 1 0 412 0 1 0
box -36 -36 89 1436
use hvDFL1sd2_CDNS_5246887918575  hvDFL1sd2_CDNS_5246887918575_0
timestamp 1701704242
transform 1 0 256 0 1 0
box -36 -36 92 1436
use hvDFL1sd2_CDNS_5246887918575  hvDFL1sd2_CDNS_5246887918575_1
timestamp 1701704242
transform 1 0 100 0 1 0
box -36 -36 92 1436
use hvDFL1sd_CDNS_5246887918573  hvDFL1sd_CDNS_5246887918573_0
timestamp 1701704242
transform -1 0 0 0 1 0
box -36 -36 89 1436
<< labels >>
flabel comment s -28 675 -28 675 0 FreeSans 300 0 0 0 S
flabel comment s 128 675 128 675 0 FreeSans 300 0 0 0 D
flabel comment s 284 675 284 675 0 FreeSans 300 0 0 0 S
flabel comment s 440 675 440 675 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 80258120
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 80256108
<< end >>
