magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< pwell >>
rect -79 -26 370 226
<< nmoslvt >>
rect 0 0 30 200
rect 86 0 116 200
rect 172 0 202 200
rect 258 0 288 200
<< ndiff >>
rect -53 182 0 200
rect -53 148 -45 182
rect -11 148 0 182
rect -53 114 0 148
rect -53 80 -45 114
rect -11 80 0 114
rect -53 46 0 80
rect -53 12 -45 46
rect -11 12 0 46
rect -53 0 0 12
rect 30 182 86 200
rect 30 148 41 182
rect 75 148 86 182
rect 30 114 86 148
rect 30 80 41 114
rect 75 80 86 114
rect 30 46 86 80
rect 30 12 41 46
rect 75 12 86 46
rect 30 0 86 12
rect 116 182 172 200
rect 116 148 127 182
rect 161 148 172 182
rect 116 114 172 148
rect 116 80 127 114
rect 161 80 172 114
rect 116 46 172 80
rect 116 12 127 46
rect 161 12 172 46
rect 116 0 172 12
rect 202 182 258 200
rect 202 148 213 182
rect 247 148 258 182
rect 202 114 258 148
rect 202 80 213 114
rect 247 80 258 114
rect 202 46 258 80
rect 202 12 213 46
rect 247 12 258 46
rect 202 0 258 12
rect 288 182 344 200
rect 288 148 299 182
rect 333 148 344 182
rect 288 114 344 148
rect 288 80 299 114
rect 333 80 344 114
rect 288 46 344 80
rect 288 12 299 46
rect 333 12 344 46
rect 288 0 344 12
<< ndiffc >>
rect -45 148 -11 182
rect -45 80 -11 114
rect -45 12 -11 46
rect 41 148 75 182
rect 41 80 75 114
rect 41 12 75 46
rect 127 148 161 182
rect 127 80 161 114
rect 127 12 161 46
rect 213 148 247 182
rect 213 80 247 114
rect 213 12 247 46
rect 299 148 333 182
rect 299 80 333 114
rect 299 12 333 46
<< poly >>
rect 0 200 30 226
rect 86 200 116 226
rect 172 200 202 226
rect 258 200 288 226
rect 0 -26 30 0
rect 86 -26 116 0
rect 172 -26 202 0
rect 258 -26 288 0
<< locali >>
rect -45 182 -11 198
rect -45 114 -11 148
rect -45 46 -11 80
rect -45 -4 -11 12
rect 41 182 75 198
rect 41 114 75 148
rect 41 46 75 80
rect 41 -4 75 12
rect 127 182 161 198
rect 127 114 161 148
rect 127 46 161 80
rect 127 -4 161 12
rect 213 182 247 198
rect 213 114 247 148
rect 213 46 247 80
rect 213 -4 247 12
rect 299 182 333 198
rect 299 114 333 148
rect 299 46 333 80
rect 299 -4 333 12
use hvDFL1sd2_CDNS_52468879185133  hvDFL1sd2_CDNS_52468879185133_0
timestamp 1701704242
transform 1 0 288 0 1 0
box 0 0 1 1
use hvDFL1sd2_CDNS_52468879185133  hvDFL1sd2_CDNS_52468879185133_1
timestamp 1701704242
transform 1 0 202 0 1 0
box 0 0 1 1
use hvDFL1sd2_CDNS_52468879185133  hvDFL1sd2_CDNS_52468879185133_2
timestamp 1701704242
transform 1 0 116 0 1 0
box 0 0 1 1
use hvDFL1sd2_CDNS_52468879185133  hvDFL1sd2_CDNS_52468879185133_3
timestamp 1701704242
transform 1 0 30 0 1 0
box 0 0 1 1
use hvDFL1sd_CDNS_52468879185132  hvDFL1sd_CDNS_52468879185132_0
timestamp 1701704242
transform -1 0 0 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s -28 97 -28 97 0 FreeSans 300 0 0 0 D
flabel comment s 58 97 58 97 0 FreeSans 300 0 0 0 S
flabel comment s 144 97 144 97 0 FreeSans 300 0 0 0 D
flabel comment s 230 97 230 97 0 FreeSans 300 0 0 0 S
flabel comment s 316 97 316 97 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 21572278
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 21569886
<< end >>
