magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 2 67 813 203
rect 29 21 813 67
rect 29 -17 63 21
<< locali >>
rect 17 199 105 265
rect 217 323 251 493
rect 481 323 530 425
rect 217 289 530 323
rect 305 181 356 289
rect 390 215 618 255
rect 652 215 811 255
rect 305 129 371 181
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 36 333 70 383
rect 117 375 183 527
rect 36 299 173 333
rect 139 249 173 299
rect 294 359 344 527
rect 391 459 607 493
rect 391 359 447 459
rect 573 333 607 459
rect 641 367 707 527
rect 741 333 796 493
rect 573 291 796 333
rect 139 215 267 249
rect 139 165 173 215
rect 36 17 70 165
rect 120 89 173 165
rect 215 95 271 181
rect 405 145 796 181
rect 405 95 455 145
rect 215 51 455 95
rect 489 17 523 111
rect 557 51 623 145
rect 657 17 691 111
rect 725 53 796 145
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
rlabel locali s 652 215 811 255 6 A1
port 1 nsew signal input
rlabel locali s 390 215 618 255 6 A2
port 2 nsew signal input
rlabel locali s 17 199 105 265 6 B1_N
port 3 nsew signal input
rlabel metal1 s 0 -48 828 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 29 21 813 67 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 2 67 813 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 866 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 828 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 305 129 371 181 6 Y
port 8 nsew signal output
rlabel locali s 305 181 356 289 6 Y
port 8 nsew signal output
rlabel locali s 217 289 530 323 6 Y
port 8 nsew signal output
rlabel locali s 481 323 530 425 6 Y
port 8 nsew signal output
rlabel locali s 217 323 251 493 6 Y
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 828 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1322534
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1315478
<< end >>
