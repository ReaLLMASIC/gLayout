magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< nwell >>
rect 6329 1414 6495 2173
<< pwell >>
rect 2477 1941 3819 2231
rect 6314 888 6400 1283
rect 2477 77 3819 367
rect 5983 289 6400 888
rect 5521 73 5733 159
rect 5521 -206 5607 73
<< pdiff >>
rect 9652 262 9689 781
<< psubdiff >>
rect 2503 2171 2721 2205
rect 2755 2171 2790 2205
rect 2824 2171 2859 2205
rect 2893 2171 2928 2205
rect 2962 2171 2997 2205
rect 2503 2137 2997 2171
rect 2503 2103 2721 2137
rect 2755 2103 2790 2137
rect 2824 2103 2859 2137
rect 2893 2103 2928 2137
rect 2962 2103 2997 2137
rect 2503 2069 2997 2103
rect 2503 2035 2721 2069
rect 2755 2035 2790 2069
rect 2824 2035 2859 2069
rect 2893 2035 2928 2069
rect 2962 2035 2997 2069
rect 2503 2001 2997 2035
rect 2503 1967 2721 2001
rect 2755 1967 2790 2001
rect 2824 1967 2859 2001
rect 2893 1967 2928 2001
rect 2962 1967 2997 2001
rect 3575 1967 3793 2205
rect 6009 838 6374 862
rect 6009 804 6136 838
rect 6170 804 6204 838
rect 6238 804 6272 838
rect 6306 804 6340 838
rect 6009 760 6374 804
rect 6009 726 6136 760
rect 6170 726 6204 760
rect 6238 726 6272 760
rect 6306 726 6340 760
rect 6009 682 6374 726
rect 6009 648 6136 682
rect 6170 648 6204 682
rect 6238 648 6272 682
rect 6306 648 6340 682
rect 6009 604 6374 648
rect 6009 570 6136 604
rect 6170 570 6204 604
rect 6238 570 6272 604
rect 6306 570 6340 604
rect 6009 527 6374 570
rect 6009 493 6136 527
rect 6170 493 6204 527
rect 6238 493 6272 527
rect 6306 493 6340 527
rect 6009 450 6374 493
rect 6009 416 6136 450
rect 6170 416 6204 450
rect 6238 416 6272 450
rect 6306 416 6340 450
rect 6009 373 6374 416
rect 2503 307 2595 341
rect 2629 307 2678 341
rect 2712 307 2760 341
rect 2794 307 2842 341
rect 2876 307 3026 341
rect 3060 307 3096 341
rect 3130 307 3166 341
rect 3200 307 3236 341
rect 3270 307 3420 341
rect 3454 307 3503 341
rect 3537 307 3585 341
rect 3619 307 3667 341
rect 3701 307 3793 341
rect 6009 339 6136 373
rect 6170 339 6204 373
rect 6238 339 6272 373
rect 6306 339 6340 373
rect 6009 315 6374 339
rect 2503 273 3793 307
rect 2503 239 2595 273
rect 2629 239 2678 273
rect 2712 239 2760 273
rect 2794 239 2842 273
rect 2876 239 3026 273
rect 3060 239 3096 273
rect 3130 239 3166 273
rect 3200 239 3236 273
rect 3270 239 3420 273
rect 3454 239 3503 273
rect 3537 239 3585 273
rect 3619 239 3667 273
rect 3701 239 3793 273
rect 2503 205 3793 239
rect 2503 171 2595 205
rect 2629 171 2678 205
rect 2712 171 2760 205
rect 2794 171 2842 205
rect 2876 171 3026 205
rect 3060 171 3096 205
rect 3130 171 3166 205
rect 3200 171 3236 205
rect 3270 171 3420 205
rect 3454 171 3503 205
rect 3537 171 3585 205
rect 3619 171 3667 205
rect 3701 171 3793 205
rect 2503 137 3793 171
rect 2503 103 2595 137
rect 2629 103 2678 137
rect 2712 103 2760 137
rect 2794 103 2842 137
rect 2876 103 3026 137
rect 3060 103 3096 137
rect 3130 103 3166 137
rect 3200 103 3236 137
rect 3270 103 3420 137
rect 3454 103 3503 137
rect 3537 103 3585 137
rect 3619 103 3667 137
rect 3701 103 3793 137
rect 5547 109 5649 133
rect 5581 99 5649 109
rect 5683 99 5707 133
rect 5547 32 5581 75
rect 5547 -45 5581 -2
rect 5547 -122 5581 -79
rect 5547 -180 5581 -156
<< mvpsubdiff >>
rect 6340 1233 6374 1257
rect 6340 1115 6374 1199
rect 6340 1057 6374 1081
<< mvnsubdiff >>
rect 6395 2083 6429 2107
rect 6395 2014 6429 2049
rect 6395 1946 6429 1980
rect 6395 1878 6429 1912
rect 6395 1810 6429 1844
rect 6395 1742 6429 1776
rect 6395 1674 6429 1708
rect 6395 1606 6429 1640
rect 6395 1538 6429 1572
rect 6395 1480 6429 1504
<< psubdiffcont >>
rect 2721 2171 2755 2205
rect 2790 2171 2824 2205
rect 2859 2171 2893 2205
rect 2928 2171 2962 2205
rect 2721 2103 2755 2137
rect 2790 2103 2824 2137
rect 2859 2103 2893 2137
rect 2928 2103 2962 2137
rect 2721 2035 2755 2069
rect 2790 2035 2824 2069
rect 2859 2035 2893 2069
rect 2928 2035 2962 2069
rect 2721 1967 2755 2001
rect 2790 1967 2824 2001
rect 2859 1967 2893 2001
rect 2928 1967 2962 2001
rect 2997 1967 3575 2205
rect 6136 804 6170 838
rect 6204 804 6238 838
rect 6272 804 6306 838
rect 6340 804 6374 838
rect 6136 726 6170 760
rect 6204 726 6238 760
rect 6272 726 6306 760
rect 6340 726 6374 760
rect 6136 648 6170 682
rect 6204 648 6238 682
rect 6272 648 6306 682
rect 6340 648 6374 682
rect 6136 570 6170 604
rect 6204 570 6238 604
rect 6272 570 6306 604
rect 6340 570 6374 604
rect 6136 493 6170 527
rect 6204 493 6238 527
rect 6272 493 6306 527
rect 6340 493 6374 527
rect 6136 416 6170 450
rect 6204 416 6238 450
rect 6272 416 6306 450
rect 6340 416 6374 450
rect 2595 307 2629 341
rect 2678 307 2712 341
rect 2760 307 2794 341
rect 2842 307 2876 341
rect 3026 307 3060 341
rect 3096 307 3130 341
rect 3166 307 3200 341
rect 3236 307 3270 341
rect 3420 307 3454 341
rect 3503 307 3537 341
rect 3585 307 3619 341
rect 3667 307 3701 341
rect 6136 339 6170 373
rect 6204 339 6238 373
rect 6272 339 6306 373
rect 6340 339 6374 373
rect 2595 239 2629 273
rect 2678 239 2712 273
rect 2760 239 2794 273
rect 2842 239 2876 273
rect 3026 239 3060 273
rect 3096 239 3130 273
rect 3166 239 3200 273
rect 3236 239 3270 273
rect 3420 239 3454 273
rect 3503 239 3537 273
rect 3585 239 3619 273
rect 3667 239 3701 273
rect 2595 171 2629 205
rect 2678 171 2712 205
rect 2760 171 2794 205
rect 2842 171 2876 205
rect 3026 171 3060 205
rect 3096 171 3130 205
rect 3166 171 3200 205
rect 3236 171 3270 205
rect 3420 171 3454 205
rect 3503 171 3537 205
rect 3585 171 3619 205
rect 3667 171 3701 205
rect 2595 103 2629 137
rect 2678 103 2712 137
rect 2760 103 2794 137
rect 2842 103 2876 137
rect 3026 103 3060 137
rect 3096 103 3130 137
rect 3166 103 3200 137
rect 3236 103 3270 137
rect 3420 103 3454 137
rect 3503 103 3537 137
rect 3585 103 3619 137
rect 3667 103 3701 137
rect 5547 75 5581 109
rect 5649 99 5683 133
rect 5547 -2 5581 32
rect 5547 -79 5581 -45
rect 5547 -156 5581 -122
<< mvpsubdiffcont >>
rect 6340 1199 6374 1233
rect 6340 1081 6374 1115
<< mvnsubdiffcont >>
rect 6395 2049 6429 2083
rect 6395 1980 6429 2014
rect 6395 1912 6429 1946
rect 6395 1844 6429 1878
rect 6395 1776 6429 1810
rect 6395 1708 6429 1742
rect 6395 1640 6429 1674
rect 6395 1572 6429 1606
rect 6395 1504 6429 1538
<< poly >>
rect 852 991 918 1007
rect 852 957 868 991
rect 902 957 918 991
rect 852 941 918 957
rect 5375 991 5441 1007
rect 5375 957 5391 991
rect 5425 957 5441 991
rect 5375 941 5441 957
<< polycont >>
rect 868 957 902 991
rect 5391 957 5425 991
<< locali >>
rect 2697 2171 2721 2205
rect 2755 2171 2790 2205
rect 2824 2171 2859 2205
rect 2893 2171 2928 2205
rect 2962 2171 2997 2205
rect 2697 2137 2997 2171
rect 2697 2103 2721 2137
rect 2755 2103 2790 2137
rect 2824 2103 2859 2137
rect 2893 2103 2928 2137
rect 2962 2103 2997 2137
rect 2697 2069 2997 2103
rect 2697 2035 2721 2069
rect 2755 2035 2790 2069
rect 2824 2035 2859 2069
rect 2893 2035 2928 2069
rect 2962 2035 2997 2069
rect 2697 2001 2997 2035
rect 2697 1967 2721 2001
rect 2755 1967 2790 2001
rect 2824 1967 2859 2001
rect 2893 1967 2928 2001
rect 2962 1967 2997 2001
rect 3575 1967 3599 2205
rect 6395 2151 6429 2189
rect 6395 2083 6429 2117
rect 6395 2014 6429 2045
rect 6395 1946 6429 1980
rect 6395 1878 6429 1912
rect 6395 1810 6429 1844
rect 6395 1742 6429 1776
rect 6395 1674 6429 1708
rect 6395 1606 6429 1640
rect 522 1549 560 1583
rect 6395 1538 6429 1572
rect 6395 1480 6429 1504
rect 6340 1233 6374 1257
rect 413 1157 448 1203
rect 5831 1123 5869 1157
rect 6340 1115 6374 1199
rect 15114 1120 15171 1154
rect 15205 1120 15262 1154
rect 15296 1120 15352 1154
rect 852 991 918 1007
rect 852 957 868 991
rect 902 975 918 991
rect 852 941 884 957
rect 5375 991 5441 1007
rect 5375 957 5391 991
rect 5425 975 5441 991
rect 5375 941 5407 957
rect 6340 862 6374 1081
rect 6009 838 6374 862
rect 6009 804 6136 838
rect 6170 804 6204 838
rect 6238 804 6272 838
rect 6306 804 6340 838
rect 6009 760 6374 804
rect 6009 726 6136 760
rect 6170 726 6204 760
rect 6238 726 6272 760
rect 6306 726 6340 760
rect 15381 778 15415 816
rect 6009 682 6374 726
rect 6009 648 6136 682
rect 6170 648 6204 682
rect 6238 648 6272 682
rect 6306 648 6340 682
rect 6009 604 6374 648
rect 6009 570 6136 604
rect 6170 570 6204 604
rect 6238 570 6272 604
rect 6306 570 6340 604
rect 6009 527 6374 570
rect 6009 493 6136 527
rect 6170 493 6204 527
rect 6238 493 6272 527
rect 6306 493 6340 527
rect 6009 450 6374 493
rect 6009 416 6136 450
rect 6170 416 6204 450
rect 6238 416 6272 450
rect 6306 416 6340 450
rect 6009 373 6374 416
rect 2503 307 2595 341
rect 2629 307 2678 341
rect 2712 307 2760 341
rect 2794 307 2842 341
rect 2876 307 2900 341
rect 2503 273 2900 307
rect 2503 239 2595 273
rect 2629 239 2678 273
rect 2712 239 2760 273
rect 2794 239 2842 273
rect 2876 239 2900 273
rect 2503 211 2900 239
rect 3002 307 3026 341
rect 3060 307 3096 341
rect 3130 307 3166 341
rect 3200 307 3236 341
rect 3270 307 3294 341
rect 3002 273 3294 307
rect 3002 239 3026 273
rect 3060 239 3096 273
rect 3130 239 3166 273
rect 3200 239 3236 273
rect 3270 239 3294 273
rect 3002 211 3294 239
rect 3396 307 3420 341
rect 3454 307 3503 341
rect 3537 307 3585 341
rect 3619 307 3667 341
rect 3701 307 3793 341
rect 6009 339 6136 373
rect 6170 339 6204 373
rect 6238 339 6272 373
rect 6306 339 6340 373
rect 6009 315 6374 339
rect 3396 273 3793 307
rect 3396 239 3420 273
rect 3454 239 3503 273
rect 3537 239 3585 273
rect 3619 239 3667 273
rect 3701 239 3793 273
rect 3396 211 3793 239
rect 2503 205 3793 211
rect 2503 171 2595 205
rect 2629 171 2678 205
rect 2712 171 2760 205
rect 2794 171 2842 205
rect 2876 171 3026 205
rect 3060 171 3096 205
rect 3130 171 3166 205
rect 3200 171 3236 205
rect 3270 171 3420 205
rect 3454 171 3503 205
rect 3537 171 3585 205
rect 3619 171 3667 205
rect 3701 171 3793 205
rect 2503 137 3793 171
rect 2503 103 2595 137
rect 2629 103 2678 137
rect 2712 103 2760 137
rect 2794 103 2842 137
rect 2876 103 3026 137
rect 3060 103 3096 137
rect 3130 103 3166 137
rect 3200 103 3236 137
rect 3270 103 3420 137
rect 3454 103 3503 137
rect 3537 103 3585 137
rect 3619 103 3667 137
rect 3701 103 3793 137
rect 5547 109 5649 133
rect 1719 61 1889 95
rect 5581 99 5649 109
rect 5683 99 5707 133
rect 1096 -40 1136 6
rect 1783 -15 1889 61
rect 1817 -49 1855 -15
rect 4665 -21 4771 61
rect 5547 32 5581 75
rect 4699 -55 4737 -21
rect 5160 -40 5200 6
rect 4665 -60 4771 -55
rect 5547 -45 5581 -2
rect 5547 -122 5581 -79
rect 5547 -180 5581 -156
rect 9919 -637 9973 276
rect 10395 223 10433 257
rect 15156 158 15204 192
rect 15238 158 15286 192
rect 15320 158 15367 192
rect 15401 158 15448 192
rect 15482 158 15529 192
rect 15563 158 15610 192
rect 9919 -671 9929 -637
rect 9963 -671 9973 -637
rect 9919 -709 9973 -671
rect 9919 -743 9929 -709
rect 9963 -743 9973 -709
<< viali >>
rect 6395 2189 6429 2223
rect 6395 2117 6429 2151
rect 6395 2049 6429 2079
rect 6395 2045 6429 2049
rect 488 1549 522 1583
rect 560 1549 594 1583
rect 5797 1123 5831 1157
rect 5869 1123 5903 1157
rect 15080 1120 15114 1154
rect 15171 1120 15205 1154
rect 15262 1120 15296 1154
rect 15352 1120 15386 1154
rect 884 957 902 975
rect 902 957 918 975
rect 884 941 918 957
rect 5407 957 5425 975
rect 5425 957 5441 975
rect 5407 941 5441 957
rect 15381 816 15415 850
rect 15381 744 15415 778
rect 1783 -49 1817 -15
rect 1855 -49 1889 -15
rect 4665 -55 4699 -21
rect 4737 -55 4771 -21
rect 10361 223 10395 257
rect 10433 223 10467 257
rect 15122 158 15156 192
rect 15204 158 15238 192
rect 15286 158 15320 192
rect 15367 158 15401 192
rect 15448 158 15482 192
rect 15529 158 15563 192
rect 15610 158 15644 192
rect 9929 -671 9963 -637
rect 9929 -743 9963 -709
<< metal1 >>
rect -179 2033 -139 2235
rect 6389 2223 6435 2235
rect 6389 2189 6395 2223
rect 6429 2189 6435 2223
rect 6389 2151 6435 2189
rect 6389 2117 6395 2151
rect 6429 2117 6435 2151
rect 6389 2079 6435 2117
rect 6389 2045 6395 2079
rect 6429 2045 6435 2079
rect 6389 2033 6435 2045
rect -179 1875 -139 2005
rect 104 1998 220 2004
rect 104 1876 220 1882
rect 6475 1998 9656 2005
rect 6475 1882 9534 1998
rect 9650 1882 9656 1998
rect 6475 1875 9656 1882
rect 476 1583 6608 1589
rect 476 1549 488 1583
rect 522 1549 560 1583
rect 594 1549 6556 1583
rect 476 1543 6556 1549
tri 6531 1518 6556 1543 ne
rect 6556 1519 6608 1531
rect 6556 1461 6608 1467
rect 6267 1235 6642 1287
rect 6694 1235 6706 1287
rect 6758 1235 6764 1287
rect 5785 1157 6731 1166
rect 5785 1123 5797 1157
rect 5831 1123 5869 1157
rect 5903 1123 6731 1157
rect 5785 1114 6731 1123
rect 6783 1114 6795 1166
rect 6847 1114 6853 1166
rect 15068 1154 15512 1160
rect 15068 1120 15080 1154
rect 15114 1120 15171 1154
rect 15205 1120 15262 1154
rect 15296 1120 15352 1154
rect 15386 1120 15512 1154
rect 15068 1114 15512 1120
tri 15459 1089 15484 1114 ne
rect -179 884 -96 1086
rect 2949 991 2955 1043
rect 3007 991 3013 1043
rect 872 975 930 987
rect 872 941 884 975
rect 918 941 930 975
rect 872 929 930 941
rect 2949 979 3013 991
rect 2949 927 2955 979
rect 3007 927 3013 979
rect 5395 975 5453 987
rect 5395 941 5407 975
rect 5441 941 5453 975
rect 5395 929 5453 941
rect 9625 884 9665 1086
rect 6049 881 6682 884
tri 6682 881 6685 884 nw
rect 6049 856 6657 881
tri 6657 856 6682 881 nw
tri 15459 856 15484 881 se
rect 15484 856 15512 1114
rect 6049 850 6651 856
tri 6651 850 6657 856 nw
tri 13246 850 13252 856 se
rect 13252 850 15512 856
rect 6049 824 6617 850
rect -120 478 247 752
rect 2994 695 3304 696
rect 2949 643 2955 695
rect 3007 643 3304 695
rect 2949 631 3304 643
rect 2949 579 2955 631
rect 3007 579 3304 631
rect 2994 576 3304 579
rect 6049 478 6111 824
rect 6463 816 6617 824
tri 6617 816 6651 850 nw
tri 13237 841 13246 850 se
rect 13246 841 15381 850
rect 6463 778 6579 816
tri 6579 778 6617 816 nw
rect 6463 744 6545 778
tri 6545 744 6579 778 nw
rect 6463 738 6539 744
tri 6539 738 6545 744 nw
rect 6463 695 6496 738
tri 6496 695 6539 738 nw
rect 9733 708 9935 841
tri 13212 816 13237 841 se
rect 13237 816 15381 841
rect 15415 816 15512 850
tri 13174 778 13212 816 se
rect 13212 778 15512 816
tri 13140 744 13174 778 se
rect 13174 744 15381 778
rect 15415 744 15512 778
tri 13134 738 13140 744 se
rect 13140 738 15512 744
tri 13129 733 13134 738 se
rect 13134 733 13270 738
tri 9935 708 9960 733 sw
tri 13104 708 13129 733 se
rect 13129 708 13270 733
tri 13270 708 13300 738 nw
tri 6463 662 6496 695 nw
rect 9733 590 13152 708
tri 13152 590 13270 708 nw
rect 9733 469 9935 590
tri 9935 565 9960 590 nw
rect 10 93 45 441
tri 9973 257 9979 263 se
rect 9979 257 10479 263
tri 9939 223 9973 257 se
rect 9973 223 10361 257
rect 10395 223 10433 257
rect 10467 223 10479 257
tri 9933 217 9939 223 se
rect 9939 217 10479 223
tri 9914 198 9933 217 se
rect 9933 198 9980 217
tri 9980 198 9999 217 nw
tri 9913 197 9914 198 se
rect 9914 197 9979 198
tri 9979 197 9980 198 nw
tri 9908 192 9913 197 se
rect 9913 192 9974 197
tri 9974 192 9979 197 nw
rect 15110 192 15656 198
tri 9874 158 9908 192 se
rect 9908 158 9940 192
tri 9940 158 9974 192 nw
rect 15110 158 15122 192
rect 15156 158 15204 192
rect 15238 158 15286 192
rect 15320 158 15367 192
rect 15401 158 15448 192
rect 15482 158 15529 192
rect 15563 158 15610 192
rect 15644 158 15656 192
tri 9847 131 9874 158 se
rect 9874 131 9913 158
tri 9913 131 9940 158 nw
tri 9809 93 9847 131 se
tri 9781 65 9809 93 se
rect 9809 65 9847 93
tri 9847 65 9913 131 nw
tri 15070 65 15110 105 se
rect 15110 65 15656 158
rect 2690 19 2736 65
rect 3560 19 3606 65
rect 6636 55 6688 61
rect 6725 13 6731 65
rect 6783 13 6795 65
rect 6847 41 9823 65
tri 9823 41 9847 65 nw
tri 15046 41 15070 65 se
rect 15070 53 15656 65
rect 15070 41 15644 53
tri 15644 41 15656 53 nw
rect 6847 25 9807 41
tri 9807 25 9823 41 nw
tri 9847 25 9863 41 se
rect 9863 25 15592 41
rect 6847 13 9795 25
tri 9795 13 9807 25 nw
tri 9835 13 9847 25 se
rect 9847 13 15592 25
tri 9832 10 9835 13 se
rect 9835 10 15592 13
rect 6636 -9 6688 3
rect 1771 -15 2117 -9
rect 1771 -49 1783 -15
rect 1817 -49 1855 -15
rect 1889 -49 2117 -15
rect 1771 -55 2117 -49
tri 2104 -61 2110 -55 ne
rect 2110 -61 2117 -55
rect 2169 -61 2181 -9
rect 2233 -61 2239 -9
rect 4379 -61 4385 -9
rect 4437 -61 4449 -9
rect 4501 -15 4507 -9
tri 4507 -15 4513 -9 sw
rect 4501 -21 4783 -15
rect 4501 -55 4665 -21
rect 4699 -55 4737 -21
rect 4771 -55 4783 -21
rect 4501 -61 4783 -55
tri 6688 -15 6713 10 sw
tri 9807 -15 9832 10 se
rect 9832 -11 15592 10
tri 15592 -11 15644 41 nw
rect 9832 -15 9881 -11
tri 9881 -15 9885 -11 nw
rect 6688 -61 9829 -15
rect 6636 -67 9829 -61
tri 9829 -67 9881 -15 nw
rect 11133 -193 11183 -141
rect 10810 -353 10862 -301
rect 9729 -583 9769 -381
rect 6480 -683 6486 -631
rect 6538 -683 6550 -631
rect 6602 -637 9975 -631
rect 6602 -671 9929 -637
rect 9963 -671 9975 -637
rect 6602 -683 9975 -671
tri 9892 -708 9917 -683 ne
rect 9917 -709 9975 -683
rect 9917 -743 9929 -709
rect 9963 -743 9975 -709
rect 9917 -749 9975 -743
<< via1 >>
rect 104 1882 220 1998
rect 9534 1882 9650 1998
rect 6556 1531 6608 1583
rect 6556 1467 6608 1519
rect 6642 1235 6694 1287
rect 6706 1235 6758 1287
rect 6731 1114 6783 1166
rect 6795 1114 6847 1166
rect 2955 991 3007 1043
rect 2955 927 3007 979
rect 2955 643 3007 695
rect 2955 579 3007 631
rect 6636 3 6688 55
rect 6731 13 6783 65
rect 6795 13 6847 65
rect 2117 -61 2169 -9
rect 2181 -61 2233 -9
rect 4385 -61 4437 -9
rect 4449 -61 4501 -9
rect 6636 -61 6688 -9
rect 6486 -683 6538 -631
rect 6550 -683 6602 -631
<< metal2 >>
rect 104 1998 220 2004
tri 2891 1926 2938 1973 se
rect 2938 1933 3994 1973
rect 2938 1926 2949 1933
tri 2949 1926 2956 1933 nw
tri 3976 1926 3983 1933 ne
rect 3983 1926 3994 1933
tri 3994 1926 4041 1973 sw
tri 2880 1915 2891 1926 se
rect 2891 1915 2938 1926
tri 2938 1915 2949 1926 nw
tri 3983 1915 3994 1926 ne
rect 3994 1915 4041 1926
rect 104 745 220 1882
tri 2871 1906 2880 1915 se
rect 2880 1906 2929 1915
tri 2929 1906 2938 1915 nw
tri 3994 1908 4001 1915 ne
tri 2835 1043 2871 1079 se
rect 2871 1061 2911 1906
tri 2911 1888 2929 1906 nw
rect 2871 1043 2893 1061
tri 2893 1043 2911 1061 nw
tri 2813 1021 2835 1043 se
rect 2835 1021 2871 1043
tri 2871 1021 2893 1043 nw
tri 2809 1017 2813 1021 se
rect 2813 1017 2867 1021
tri 2867 1017 2871 1021 nw
tri 2265 991 2291 1017 se
rect 2291 991 2841 1017
tri 2841 991 2867 1017 nw
rect 2949 991 2955 1043
rect 3007 991 3013 1043
tri 2253 979 2265 991 se
rect 2265 979 2829 991
tri 2829 979 2841 991 nw
rect 2949 979 3013 991
tri 2233 959 2253 979 se
rect 2253 977 2827 979
tri 2827 977 2829 979 nw
rect 2253 959 2291 977
tri 2291 959 2309 977 nw
tri 2201 927 2233 959 se
rect 2233 927 2259 959
tri 2259 927 2291 959 nw
rect 2949 927 2955 979
rect 3007 927 3013 979
tri 2199 925 2201 927 se
rect 2201 925 2257 927
tri 2257 925 2259 927 nw
tri 2177 3 2199 25 se
rect 2199 3 2239 925
tri 2239 907 2257 925 nw
rect 2949 695 3013 927
rect 2949 643 2955 695
rect 3007 643 3013 695
rect 2949 631 3013 643
rect 2949 579 2955 631
rect 3007 579 3013 631
rect 4001 579 4041 1915
rect 9528 1882 9534 1998
rect 9650 1882 9656 1998
rect 6556 1583 6608 1589
rect 6556 1519 6608 1531
tri 4041 579 4047 585 sw
rect 4001 567 4047 579
tri 4001 533 4035 567 ne
rect 4035 533 4047 567
tri 4047 533 4093 579 sw
tri 4035 527 4041 533 ne
rect 4041 527 4390 533
tri 4041 493 4075 527 ne
rect 4075 493 4390 527
tri 4372 475 4390 493 ne
tri 4390 475 4448 533 sw
tri 4390 457 4408 475 ne
tri 4391 3 4408 20 se
rect 4408 3 4448 475
tri 4448 3 4495 50 sw
tri 2165 -9 2177 3 se
rect 2177 -9 2239 3
rect 2110 -61 2117 -9
rect 2169 -61 2181 -9
rect 2233 -61 2239 -9
tri 4379 -9 4391 3 se
rect 4391 -9 4495 3
tri 4495 -9 4507 3 sw
rect 4379 -61 4385 -9
rect 4437 -61 4449 -9
rect 4501 -61 4507 -9
rect 6128 -123 6448 816
tri 6531 -631 6556 -606 se
rect 6556 -631 6608 1467
rect 6636 1235 6642 1287
rect 6694 1235 6706 1287
rect 6758 1235 6764 1287
rect 6636 55 6688 1235
tri 6688 1210 6713 1235 nw
rect 6725 1114 6731 1166
rect 6783 1114 6795 1166
rect 6847 1114 6853 1166
rect 6725 65 6777 1114
tri 6777 1089 6802 1114 nw
rect 9528 469 9656 1882
rect 11136 579 11946 1247
tri 11136 534 11181 579 ne
tri 6777 65 6802 90 sw
rect 6725 13 6731 65
rect 6783 13 6795 65
rect 6847 13 6853 65
rect 6636 -9 6688 3
rect 6636 -67 6688 -61
rect 11181 -583 11946 579
rect 6480 -683 6486 -631
rect 6538 -683 6550 -631
rect 6602 -683 6608 -631
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_0
timestamp 1701704242
transform 1 0 9929 0 -1 -637
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_1
timestamp 1701704242
transform 1 0 15381 0 -1 850
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1701704242
transform -1 0 1889 0 1 -49
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1701704242
transform -1 0 5903 0 1 1123
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1701704242
transform -1 0 4771 0 1 -55
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_3
timestamp 1701704242
transform 1 0 488 0 1 1549
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_4
timestamp 1701704242
transform 1 0 10361 0 1 223
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_0
timestamp 1701704242
transform 0 -1 6429 1 0 2045
box 0 0 1 1
use L1M1_CDNS_52468879185191  L1M1_CDNS_52468879185191_0
timestamp 1701704242
transform -1 0 3570 0 1 1965
box -12 -6 838 40
use L1M1_CDNS_524688791851423  L1M1_CDNS_524688791851423_0
timestamp 1701704242
transform 0 1 6117 -1 0 812
box -12 -6 334 256
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_0
timestamp 1701704242
transform 0 -1 6608 -1 0 1589
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_1
timestamp 1701704242
transform 0 -1 6688 1 0 -67
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_2
timestamp 1701704242
transform 1 0 6480 0 1 -683
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_3
timestamp 1701704242
transform 1 0 6725 0 1 1114
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_4
timestamp 1701704242
transform 1 0 6636 0 1 1235
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_5
timestamp 1701704242
transform 1 0 6725 0 1 13
box 0 0 1 1
use M1M2_CDNS_52468879185197  M1M2_CDNS_52468879185197_0
timestamp 1701704242
transform 0 -1 220 1 0 489
box 0 0 256 116
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_0
timestamp 1701704242
transform 0 -1 220 -1 0 2004
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_1
timestamp 1701704242
transform 1 0 9528 0 1 1882
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_0
timestamp 1701704242
transform -1 0 3013 0 1 927
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_1
timestamp 1701704242
transform -1 0 3013 0 -1 695
box 0 0 1 1
use M1M2_CDNS_524688791851246  M1M2_CDNS_524688791851246_0
timestamp 1701704242
transform 1 0 6128 0 -1 803
box 0 0 320 308
use M1M2_CDNS_524688791851424  M1M2_CDNS_524688791851424_0
timestamp 1701704242
transform 0 1 11181 -1 0 -386
box 0 0 192 756
use PYM1_CDNS_524688791851422  PYM1_CDNS_524688791851422_0
timestamp 1701704242
transform 0 -1 918 1 0 941
box 0 0 1 1
use PYM1_CDNS_524688791851422  PYM1_CDNS_524688791851422_1
timestamp 1701704242
transform 0 -1 5441 1 0 941
box 0 0 1 1
use sky130_fd_io__sio_cclat  sky130_fd_io__sio_cclat_0
timestamp 1701704242
transform 1 0 9647 0 -1 1303
box -124 145 6234 2367
use sky130_fd_io__sio_com_dat_ls  sky130_fd_io__sio_com_dat_ls_0
timestamp 1701704242
transform -1 0 6296 0 -1 2339
box -179 14 3312 2420
use sky130_fd_io__sio_com_dat_ls  sky130_fd_io__sio_com_dat_ls_1
timestamp 1701704242
transform 1 0 0 0 -1 2339
box -179 14 3312 2420
<< labels >>
flabel comment s 9690 44 9690 44 0 FreeSans 300 0 0 0 pu_dis_h
flabel comment s 9687 -31 9687 -31 0 FreeSans 300 0 0 0 pd_dis_h
flabel comment s 6318 1571 6318 1571 0 FreeSans 300 0 0 0 oe_h_n
flabel comment s 6224 1264 6224 1264 0 FreeSans 300 0 0 0 pd_dis_h
flabel comment s 6228 1145 6228 1145 0 FreeSans 300 0 0 0 pu_dis_h
flabel metal1 s 9729 -583 9769 -381 3 FreeSans 300 0 0 0 vcc_io
port 2 nsew
flabel metal1 s 9625 884 9665 1086 3 FreeSans 300 0 0 0 vgnd
port 3 nsew
flabel metal1 s 2690 19 2736 65 7 FreeSans 300 0 0 0 oe_n
port 4 nsew
flabel metal1 s 3560 19 3606 65 3 FreeSans 300 0 0 0 din
port 5 nsew
flabel metal1 s 10 93 45 441 3 FreeSans 300 180 0 0 vpwr_ka
port 6 nsew
flabel metal1 s -179 884 -139 1086 3 FreeSans 300 180 0 0 vgnd
port 3 nsew
flabel metal1 s -179 2033 -139 2235 3 FreeSans 300 180 0 0 vcc_io
port 2 nsew
flabel metal1 s -179 1875 -139 2005 3 FreeSans 300 180 0 0 vgnd
port 3 nsew
flabel metal1 s 10810 -353 10862 -301 3 FreeSans 300 0 0 0 drvlo_h_n
port 7 nsew
flabel metal1 s 11133 -193 11183 -141 3 FreeSans 300 0 0 0 drvhi_h
port 8 nsew
flabel locali s 1096 -40 1136 6 7 FreeSans 300 180 0 0 od_h
port 9 nsew
flabel locali s 5160 -40 5200 6 3 FreeSans 300 180 0 0 od_h
port 9 nsew
flabel locali s 413 1157 448 1203 3 FreeSans 300 0 0 0 oe_h
port 10 nsew
flabel locali s 1816 -40 1856 6 7 FreeSans 300 180 0 0 hld_i_ovr_h
port 11 nsew
flabel metal2 s 6129 -122 6447 -90 0 FreeSans 200 0 0 0 vgnd
port 3 nsew
<< properties >>
string GDS_END 87654658
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 87633720
string path 55.975 -0.875 52.750 -0.875 
<< end >>
