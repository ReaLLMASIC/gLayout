magic
tech sky130B
timestamp 1701704242
<< properties >>
string GDS_END 16744910
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 16744458
<< end >>
