magic
tech sky130A
timestamp 1701704242
<< metal1 >>
rect 0 0 3 314
rect 541 0 544 314
<< via1 >>
rect 3 0 541 314
<< metal2 >>
rect 0 0 3 314
rect 541 0 544 314
<< properties >>
string GDS_END 88455536
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 88444524
<< end >>
