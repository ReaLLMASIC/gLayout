magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< pwell >>
rect -76 -26 4988 1426
<< nmos >>
rect 0 0 1600 1400
rect 1656 0 3256 1400
rect 3312 0 4912 1400
<< ndiff >>
rect -50 0 0 1400
rect 4912 0 4962 1400
<< poly >>
rect 0 1400 1600 1432
rect 0 -32 1600 0
rect 1656 1400 3256 1432
rect 1656 -32 3256 0
rect 3312 1400 4912 1432
rect 3312 -32 4912 0
<< locali >>
rect -45 -4 -11 1354
rect 1611 -4 1645 1354
rect 3267 -4 3301 1354
rect 4923 -4 4957 1354
use hvDFL1sd2_CDNS_55959141808559  hvDFL1sd2_CDNS_55959141808559_0
timestamp 1701704242
transform 1 0 1600 0 1 0
box -26 -26 82 1426
use hvDFL1sd2_CDNS_55959141808559  hvDFL1sd2_CDNS_55959141808559_1
timestamp 1701704242
transform 1 0 3256 0 1 0
box -26 -26 82 1426
use hvDFL1sd_CDNS_55959141808700  hvDFL1sd_CDNS_55959141808700_0
timestamp 1701704242
transform -1 0 0 0 1 0
box -26 -26 79 1426
use hvDFL1sd_CDNS_55959141808700  hvDFL1sd_CDNS_55959141808700_1
timestamp 1701704242
transform 1 0 4912 0 1 0
box -26 -26 79 1426
<< labels >>
flabel comment s 4940 675 4940 675 0 FreeSans 300 0 0 0 D
flabel comment s 3284 675 3284 675 0 FreeSans 300 0 0 0 S
flabel comment s 1628 675 1628 675 0 FreeSans 300 0 0 0 D
flabel comment s -28 675 -28 675 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 2737958
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 2736132
<< end >>
