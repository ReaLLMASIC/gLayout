magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -53 1526 529 2316
rect 3675 1526 4733 2312
rect 7879 1526 8937 2312
<< pwell >>
rect -43 97 43 1056
rect 4161 97 4247 749
rect 8365 97 8451 749
rect 12516 97 12602 749
rect 14957 97 15043 1056
<< nsubdiff >>
rect -17 2276 493 2280
rect -17 2252 93 2276
rect 17 2242 93 2252
rect 127 2242 201 2276
rect 235 2242 493 2276
rect 3945 2242 3969 2276
rect 4003 2242 4042 2276
rect 4076 2242 4115 2276
rect 4149 2242 4188 2276
rect 4222 2242 4261 2276
rect 4295 2242 4333 2276
rect 4367 2242 4405 2276
rect 4439 2242 4463 2276
rect 8149 2242 8173 2276
rect 8207 2242 8246 2276
rect 8280 2242 8319 2276
rect 8353 2242 8392 2276
rect 8426 2242 8465 2276
rect 8499 2242 8537 2276
rect 8571 2242 8609 2276
rect 8643 2242 8667 2276
rect -17 2182 17 2218
rect -17 2112 17 2148
rect -17 2042 17 2078
rect -17 1972 17 2008
rect -17 1902 17 1938
rect -17 1832 17 1868
rect -17 1762 17 1798
rect -17 1691 17 1728
rect -17 1620 17 1657
rect -17 1562 17 1586
rect 4187 2166 4221 2242
rect 4187 2097 4221 2132
rect 4187 2028 4221 2063
rect 4187 1960 4221 1994
rect 4187 1892 4221 1926
rect 4187 1824 4221 1858
rect 4187 1756 4221 1790
rect 4187 1688 4221 1722
rect 4187 1620 4221 1654
rect 4187 1562 4221 1586
rect 8391 2166 8425 2242
rect 8391 2097 8425 2132
rect 8391 2028 8425 2063
rect 8391 1960 8425 1994
rect 8391 1892 8425 1926
rect 8391 1824 8425 1858
rect 8391 1756 8425 1790
rect 8391 1688 8425 1722
rect 8391 1620 8425 1654
rect 8391 1562 8425 1586
<< mvpsubdiff >>
rect -17 1006 17 1030
rect -17 937 17 972
rect -17 868 17 903
rect -17 799 17 834
rect -17 730 17 765
rect 14983 1006 15017 1030
rect 14983 937 15017 972
rect 14983 868 15017 903
rect 14983 799 15017 834
rect 14983 730 15017 765
rect -17 661 17 696
rect -17 592 17 627
rect -17 523 17 558
rect -17 454 17 489
rect -17 385 17 420
rect -17 317 17 351
rect -17 249 17 283
rect -17 181 17 215
rect -17 123 17 147
rect 4187 699 4221 723
rect 4187 625 4221 665
rect 4187 551 4221 591
rect 4187 477 4221 517
rect 4187 403 4221 443
rect 4187 329 4221 369
rect 4187 255 4221 295
rect 4187 181 4221 221
rect 4187 123 4221 147
rect 8391 699 8425 723
rect 8391 625 8425 665
rect 8391 551 8425 591
rect 8391 477 8425 517
rect 8391 403 8425 443
rect 8391 329 8425 369
rect 8391 255 8425 295
rect 8391 181 8425 221
rect 8391 123 8425 147
rect 12542 699 12576 723
rect 12542 625 12576 665
rect 12542 551 12576 591
rect 12542 477 12576 517
rect 12542 403 12576 443
rect 12542 329 12576 369
rect 12542 255 12576 295
rect 12542 181 12576 221
rect 12542 123 12576 147
rect 14983 661 15017 696
rect 14983 592 15017 627
rect 14983 523 15017 558
rect 14983 454 15017 489
rect 14983 385 15017 420
rect 14983 317 15017 351
rect 14983 249 15017 283
rect 14983 181 15017 215
rect 14983 123 15017 147
<< nsubdiffcont >>
rect -17 2218 17 2252
rect 93 2242 127 2276
rect 201 2242 235 2276
rect 3969 2242 4003 2276
rect 4042 2242 4076 2276
rect 4115 2242 4149 2276
rect 4188 2242 4222 2276
rect 4261 2242 4295 2276
rect 4333 2242 4367 2276
rect 4405 2242 4439 2276
rect 8173 2242 8207 2276
rect 8246 2242 8280 2276
rect 8319 2242 8353 2276
rect 8392 2242 8426 2276
rect 8465 2242 8499 2276
rect 8537 2242 8571 2276
rect 8609 2242 8643 2276
rect -17 2148 17 2182
rect -17 2078 17 2112
rect -17 2008 17 2042
rect -17 1938 17 1972
rect -17 1868 17 1902
rect -17 1798 17 1832
rect -17 1728 17 1762
rect -17 1657 17 1691
rect -17 1586 17 1620
rect 4187 2132 4221 2166
rect 4187 2063 4221 2097
rect 4187 1994 4221 2028
rect 4187 1926 4221 1960
rect 4187 1858 4221 1892
rect 4187 1790 4221 1824
rect 4187 1722 4221 1756
rect 4187 1654 4221 1688
rect 4187 1586 4221 1620
rect 8391 2132 8425 2166
rect 8391 2063 8425 2097
rect 8391 1994 8425 2028
rect 8391 1926 8425 1960
rect 8391 1858 8425 1892
rect 8391 1790 8425 1824
rect 8391 1722 8425 1756
rect 8391 1654 8425 1688
rect 8391 1586 8425 1620
<< mvpsubdiffcont >>
rect -17 972 17 1006
rect -17 903 17 937
rect -17 834 17 868
rect -17 765 17 799
rect -17 696 17 730
rect 14983 972 15017 1006
rect 14983 903 15017 937
rect 14983 834 15017 868
rect 14983 765 15017 799
rect -17 627 17 661
rect -17 558 17 592
rect -17 489 17 523
rect -17 420 17 454
rect -17 351 17 385
rect -17 283 17 317
rect -17 215 17 249
rect -17 147 17 181
rect 4187 665 4221 699
rect 4187 591 4221 625
rect 4187 517 4221 551
rect 4187 443 4221 477
rect 4187 369 4221 403
rect 4187 295 4221 329
rect 4187 221 4221 255
rect 4187 147 4221 181
rect 8391 665 8425 699
rect 8391 591 8425 625
rect 8391 517 8425 551
rect 8391 443 8425 477
rect 8391 369 8425 403
rect 8391 295 8425 329
rect 8391 221 8425 255
rect 8391 147 8425 181
rect 12542 665 12576 699
rect 12542 591 12576 625
rect 12542 517 12576 551
rect 12542 443 12576 477
rect 12542 369 12576 403
rect 12542 295 12576 329
rect 12542 221 12576 255
rect 12542 147 12576 181
rect 14983 696 15017 730
rect 14983 627 15017 661
rect 14983 558 15017 592
rect 14983 489 15017 523
rect 14983 420 15017 454
rect 14983 351 15017 385
rect 14983 283 15017 317
rect 14983 215 15017 249
rect 14983 147 15017 181
<< locali >>
rect -17 2276 74 2280
rect 259 2276 493 2280
rect -17 2252 93 2276
rect 17 2246 93 2252
rect 69 2242 93 2246
rect 127 2242 201 2276
rect 235 2248 493 2276
rect 235 2242 259 2248
rect 3945 2242 3969 2276
rect 4003 2242 4042 2276
rect 4076 2242 4115 2276
rect 4149 2242 4188 2276
rect 4222 2242 4261 2276
rect 4295 2242 4333 2276
rect 4367 2242 4405 2276
rect 4439 2242 4463 2276
rect 8149 2242 8173 2276
rect 8207 2242 8246 2276
rect 8280 2242 8319 2276
rect 8353 2242 8392 2276
rect 8426 2242 8465 2276
rect 8499 2242 8537 2276
rect 8571 2242 8609 2276
rect 8643 2242 8667 2276
rect -17 2182 17 2218
rect -17 2112 17 2148
rect -17 2042 17 2078
rect -17 1972 17 2008
rect -17 1902 17 1938
rect -17 1832 17 1868
rect -17 1762 17 1798
rect -17 1691 17 1728
rect -17 1620 17 1657
rect -17 1562 17 1586
rect 2563 1205 2669 2227
rect 4187 2166 4221 2190
rect 4187 2097 4221 2132
rect 4187 2028 4221 2063
rect 4187 1960 4221 1994
rect 4187 1892 4221 1926
rect 4187 1824 4221 1858
rect 4187 1756 4221 1790
rect 4187 1688 4221 1722
rect 4187 1620 4221 1654
rect 4187 1562 4221 1586
rect 5739 1205 5845 2227
rect 6767 1205 6873 2227
rect 8391 2166 8425 2190
rect 8391 2097 8425 2132
rect 8391 2028 8425 2063
rect 8391 1960 8425 1994
rect 8391 1892 8425 1926
rect 8391 1824 8425 1858
rect 8391 1756 8425 1790
rect 8391 1688 8425 1722
rect 8391 1620 8425 1654
rect 8391 1562 8425 1586
rect 9943 1205 10049 2227
rect 10971 1205 11077 2227
rect -17 1006 17 1030
rect -17 937 17 972
rect -17 868 17 903
rect 14983 1006 15017 1030
rect 14983 937 15017 972
rect 14983 868 15017 903
rect -17 799 17 834
rect -17 730 17 765
rect -17 661 17 696
rect -17 592 17 627
rect -17 523 17 558
rect -17 454 17 489
rect -17 385 17 404
rect -17 317 17 332
rect -17 249 17 283
rect -17 181 17 215
rect -17 123 17 147
rect 4187 699 4221 856
rect 4187 625 4221 665
rect 4187 551 4221 591
rect 4187 477 4221 517
rect 4187 438 4221 443
rect 4187 403 4221 404
rect 4187 366 4221 369
rect 4187 329 4221 332
rect 4187 255 4221 295
rect 4187 181 4221 221
rect 4187 123 4221 147
rect 8391 699 8425 856
rect 12595 723 12629 823
rect 8391 625 8425 665
rect 8391 551 8425 591
rect 12542 699 12629 723
rect 12576 665 12629 699
rect 12542 625 12629 665
rect 12576 591 12629 625
rect 12542 551 12629 591
rect 8391 477 8425 517
rect 12212 484 12250 518
rect 12576 517 12629 551
rect 8391 438 8425 443
rect 8391 403 8425 404
rect 8391 366 8425 369
rect 8391 329 8425 332
rect 8391 255 8425 295
rect 8391 181 8425 221
rect 8391 123 8425 147
rect 12542 477 12629 517
rect 12576 443 12629 477
rect 12542 438 12629 443
rect 12542 404 12563 438
rect 12597 404 12629 438
rect 12542 403 12629 404
rect 12576 369 12629 403
rect 12542 366 12629 369
rect 12542 332 12563 366
rect 12597 332 12629 366
rect 12542 329 12629 332
rect 12576 295 12629 329
rect 12542 255 12629 295
rect 12576 221 12629 255
rect 12542 181 12629 221
rect 12576 147 12629 181
rect 12542 123 12629 147
rect 14983 799 15017 834
rect 14983 730 15017 765
rect 14983 661 15017 696
rect 14983 592 15017 627
rect 14983 523 15017 558
rect 14983 454 15017 489
rect 14983 385 15017 404
rect 14983 317 15017 332
rect 14983 249 15017 283
rect 14983 181 15017 215
rect 14983 123 15017 147
rect 245 16 283 50
rect 598 16 636 50
rect 670 16 708 50
rect 742 16 780 50
rect 814 16 852 50
rect 3294 16 3332 50
rect 3366 16 3404 50
rect 3438 16 3476 50
rect 3510 16 3548 50
rect 3582 16 3620 50
rect 3757 16 3795 50
rect 3947 16 3985 50
rect 4449 16 4487 50
rect 4787 16 4825 50
rect 4859 16 4897 50
rect 4931 16 4969 50
rect 5003 16 5041 50
rect 5075 16 5113 50
rect 7571 16 7609 50
rect 7643 16 7681 50
rect 7715 16 7753 50
rect 7787 16 7825 50
rect 7961 16 7999 50
rect 8151 16 8189 50
rect 8653 16 8691 50
rect 8823 16 8861 50
rect 8991 16 9029 50
rect 9063 16 9101 50
rect 9135 16 9173 50
rect 9207 16 9245 50
rect 9279 16 9317 50
rect 455 -22 489 16
rect 4659 -22 4693 16
rect 11657 -8 12063 50
rect 12165 16 12203 50
rect 11657 -42 11669 -8
rect 11703 -42 11741 -8
rect 11775 -42 11813 -8
rect 11847 -42 11885 -8
rect 11919 -42 11957 -8
rect 11991 -42 12029 -8
rect 12315 -21 12349 17
<< viali >>
rect -17 420 17 438
rect -17 404 17 420
rect -17 351 17 366
rect -17 332 17 351
rect 4187 404 4221 438
rect 4187 332 4221 366
rect 12178 484 12212 518
rect 12250 484 12284 518
rect 8391 404 8425 438
rect 8391 332 8425 366
rect 12563 404 12597 438
rect 12563 332 12597 366
rect 14983 420 15017 438
rect 14983 404 15017 420
rect 14983 351 15017 366
rect 14983 332 15017 351
rect 211 16 245 50
rect 283 16 317 50
rect 455 16 489 50
rect 564 16 598 50
rect 636 16 670 50
rect 708 16 742 50
rect 780 16 814 50
rect 852 16 886 50
rect 3260 16 3294 50
rect 3332 16 3366 50
rect 3404 16 3438 50
rect 3476 16 3510 50
rect 3548 16 3582 50
rect 3620 16 3654 50
rect 3723 16 3757 50
rect 3795 16 3829 50
rect 3913 16 3947 50
rect 3985 16 4019 50
rect 4415 16 4449 50
rect 4487 16 4521 50
rect 4659 16 4693 50
rect 4753 16 4787 50
rect 4825 16 4859 50
rect 4897 16 4931 50
rect 4969 16 5003 50
rect 5041 16 5075 50
rect 5113 16 5147 50
rect 7537 16 7571 50
rect 7609 16 7643 50
rect 7681 16 7715 50
rect 7753 16 7787 50
rect 7825 16 7859 50
rect 7927 16 7961 50
rect 7999 16 8033 50
rect 8117 16 8151 50
rect 8189 16 8223 50
rect 8619 16 8653 50
rect 8691 16 8725 50
rect 8789 16 8823 50
rect 8861 16 8895 50
rect 8957 16 8991 50
rect 9029 16 9063 50
rect 9101 16 9135 50
rect 9173 16 9207 50
rect 9245 16 9279 50
rect 9317 16 9351 50
rect 455 -56 489 -22
rect 4659 -56 4693 -22
rect 12131 16 12165 50
rect 12203 16 12237 50
rect 12315 17 12349 51
rect 11669 -42 11703 -8
rect 11741 -42 11775 -8
rect 11813 -42 11847 -8
rect 11885 -42 11919 -8
rect 11957 -42 11991 -8
rect 12029 -42 12063 -8
rect 12315 -55 12349 -21
<< metal1 >>
rect 846 2382 898 2388
tri 821 2312 846 2337 se
rect 846 2318 898 2330
rect 757 2266 846 2312
tri 898 2312 923 2337 sw
rect 898 2266 3323 2312
rect 757 2260 3323 2266
rect 3375 2260 3387 2312
rect 3439 2260 4980 2312
rect 5032 2260 5044 2312
rect 5096 2260 7760 2312
rect 7812 2260 7824 2312
rect 7876 2260 9184 2312
rect 9236 2260 9248 2312
rect 9300 2260 11866 2312
rect 11868 2311 11904 2312
rect 11867 2261 11905 2311
rect 11868 2260 11904 2261
rect 11906 2260 11964 2312
rect 12016 2260 12028 2312
rect 12080 2260 12086 2312
rect 12581 2114 12912 2232
rect 185 2086 12912 2114
rect 185 1884 219 2086
rect 4019 1884 4389 2086
rect 8223 1884 8593 2086
rect 12427 1884 12931 2086
tri 4072 1521 4091 1540 sw
tri 4317 1521 4336 1540 se
tri 1997 1515 2003 1521 se
rect 2003 1515 2760 1521
tri 2760 1515 2766 1521 sw
rect 4072 1515 4091 1521
tri 4091 1515 4097 1521 sw
tri 4311 1515 4317 1521 se
rect 4317 1515 4336 1521
tri 8276 1515 8301 1540 sw
tri 8515 1515 8540 1540 se
tri 12480 1515 12505 1540 sw
rect 1990 1469 2766 1515
rect 4050 1469 12594 1515
rect 12693 1469 13043 1515
rect -14 1239 12874 1441
rect 12495 1159 12898 1211
tri 12635 1134 12660 1159 nw
rect 54 1089 119 1097
rect 54 1043 175 1089
rect 4071 1049 4105 1083
rect 4303 1049 4337 1083
rect 8275 1049 8309 1083
rect 8507 1049 8541 1083
rect 12479 1049 12513 1083
rect 54 1039 119 1043
rect 12474 889 12784 941
tri 12635 864 12660 889 nw
rect 109 735 186 787
rect 188 786 224 787
rect 187 736 225 786
rect 226 781 303 787
rect 188 735 224 736
rect 226 735 251 781
rect 109 627 161 735
tri 161 710 186 735 nw
tri 226 710 251 735 ne
rect 251 717 303 729
rect 251 659 303 665
rect 304 660 305 786
rect 341 660 342 786
rect 343 659 401 787
rect 403 786 439 787
rect 402 660 440 786
rect 441 781 518 787
rect 493 735 518 781
rect 519 736 520 786
rect 556 736 557 786
rect 558 735 635 787
rect 441 717 493 729
tri 493 710 518 735 nw
tri 558 710 583 735 ne
rect 403 659 439 660
rect 441 659 493 665
tri 161 627 186 652 sw
tri 558 627 583 652 se
rect 583 627 635 735
rect 3569 735 3646 787
rect 3647 736 3648 786
rect 3684 736 3685 786
rect 3686 781 3763 787
rect 3765 786 3801 787
rect 3686 735 3711 781
rect 1747 663 1781 697
rect 2423 663 2457 697
tri 635 627 660 652 sw
tri 3544 627 3569 652 se
rect 3569 627 3621 735
tri 3621 710 3646 735 nw
tri 3686 710 3711 735 ne
rect 3711 717 3763 729
rect 3711 659 3763 665
rect 3764 660 3802 786
rect 3765 659 3801 660
rect 3803 659 3861 787
rect 3862 660 3863 786
rect 3899 660 3900 786
rect 3901 781 3978 787
rect 3980 786 4016 787
rect 3953 735 3978 781
rect 3979 736 4017 786
rect 3980 735 4016 736
rect 4018 735 4095 787
rect 3901 717 3953 729
tri 3953 710 3978 735 nw
tri 4018 710 4043 735 ne
rect 3901 659 3953 665
tri 3621 627 3646 652 sw
tri 4018 627 4043 652 se
rect 4043 627 4095 735
rect 4313 735 4390 787
rect 4392 786 4428 787
rect 4391 736 4429 786
rect 4430 781 4507 787
rect 4392 735 4428 736
rect 4430 735 4455 781
tri 4095 627 4120 652 sw
rect 4313 627 4365 735
tri 4365 710 4390 735 nw
tri 4430 710 4455 735 ne
rect 4455 717 4507 729
rect 4455 659 4507 665
rect 4508 660 4509 786
rect 4545 660 4546 786
rect 4547 659 4605 787
rect 4607 786 4643 787
rect 4606 660 4644 786
rect 4645 781 4722 787
rect 4697 735 4722 781
rect 4723 736 4724 786
rect 4760 736 4761 786
rect 4762 735 4839 787
rect 4645 717 4697 729
tri 4697 710 4722 735 nw
tri 4762 710 4787 735 ne
rect 4607 659 4643 660
rect 4645 659 4697 665
tri 4365 627 4390 652 sw
tri 4762 627 4787 652 se
rect 4787 627 4839 735
rect 7773 735 7850 787
rect 7851 736 7852 786
rect 7888 736 7889 786
rect 7890 781 7967 787
rect 7969 786 8005 787
rect 7890 735 7915 781
rect 5951 663 5985 697
rect 6627 663 6660 697
tri 4839 627 4864 652 sw
tri 7748 627 7773 652 se
rect 7773 627 7825 735
tri 7825 710 7850 735 nw
tri 7890 710 7915 735 ne
rect 7915 717 7967 729
rect 7915 659 7967 665
rect 7968 660 8006 786
rect 7969 659 8005 660
rect 8007 659 8065 787
rect 8066 660 8067 786
rect 8103 660 8104 786
rect 8105 781 8182 787
rect 8184 786 8220 787
rect 8157 735 8182 781
rect 8183 736 8221 786
rect 8184 735 8220 736
rect 8222 735 8299 787
rect 8105 717 8157 729
tri 8157 710 8182 735 nw
tri 8222 710 8247 735 ne
rect 8105 659 8157 665
tri 7825 627 7850 652 sw
tri 8222 627 8247 652 se
rect 8247 627 8299 735
rect 8517 735 8594 787
rect 8596 786 8632 787
rect 8595 736 8633 786
rect 8634 781 8711 787
rect 8596 735 8632 736
rect 8634 735 8659 781
tri 8299 627 8324 652 sw
tri 8492 627 8517 652 se
rect 8517 627 8569 735
tri 8569 710 8594 735 nw
tri 8634 710 8659 735 ne
rect 8659 717 8711 729
rect 8659 659 8711 665
rect 8712 660 8713 786
rect 8749 660 8750 786
rect 8751 659 8809 787
rect 8811 786 8847 787
rect 8810 660 8848 786
rect 8849 781 8926 787
rect 8901 735 8926 781
rect 8927 736 8928 786
rect 8964 736 8965 786
rect 8966 735 9043 787
rect 8849 717 8901 729
tri 8901 710 8926 735 nw
tri 8966 710 8991 735 ne
rect 8811 659 8847 660
rect 8849 659 8901 665
tri 8569 627 8594 652 sw
tri 8966 627 8991 652 se
rect 8991 627 9043 735
rect 11977 735 12054 787
rect 12055 736 12056 786
rect 12092 736 12093 786
rect 12094 781 12171 787
rect 12173 786 12209 787
rect 12094 735 12119 781
rect 10155 663 10189 697
rect 10831 663 10865 697
tri 9043 627 9068 652 sw
tri 11952 627 11977 652 se
rect 11977 627 12029 735
tri 12029 710 12054 735 nw
tri 12094 710 12119 735 ne
rect 12119 717 12171 729
rect 12119 659 12171 665
rect 12172 660 12210 786
rect 12173 659 12209 660
rect 12211 659 12269 787
rect 12270 660 12271 786
rect 12307 660 12308 786
rect 12309 781 12386 787
rect 12388 786 12424 787
rect 12361 735 12386 781
rect 12387 736 12425 786
rect 12388 735 12424 736
rect 12426 735 12503 787
rect 12309 717 12361 729
tri 12361 710 12386 735 nw
tri 12426 710 12451 735 ne
rect 12309 659 12361 665
tri 12029 627 12054 652 sw
tri 12426 627 12451 652 se
rect 12451 627 12503 735
tri 12503 627 12528 652 sw
rect 109 581 12697 627
rect 12166 536 12266 542
rect 12166 518 12214 536
tri 12266 524 12284 542 sw
rect 12266 518 12683 524
rect 12166 484 12178 518
rect 12212 484 12214 518
rect 12284 484 12683 518
rect 12166 478 12683 484
rect -23 438 34 450
rect -23 404 -17 438
rect 17 404 34 438
rect -23 366 34 404
rect -23 332 -17 366
rect 17 332 34 366
rect -23 320 34 332
rect 4181 438 4227 450
rect 4181 404 4187 438
rect 4221 404 4227 438
rect 4181 366 4227 404
rect 4181 332 4187 366
rect 4221 332 4227 366
rect 4181 320 4227 332
rect 8385 438 8431 450
rect 8385 404 8391 438
rect 8425 404 8431 438
rect 8385 366 8431 404
rect 8385 332 8391 366
rect 8425 332 8431 366
rect 8385 320 8431 332
rect 12557 438 15023 450
rect 12557 404 12563 438
rect 12597 404 14983 438
rect 15017 404 15023 438
rect 12557 366 15023 404
rect 12557 332 12563 366
rect 12597 332 14983 366
rect 15017 332 15023 366
rect 12557 320 15023 332
rect 0 90 34 292
tri 12009 65 12034 90 ne
rect 12034 65 12086 117
rect 12536 90 12885 292
tri 12086 65 12111 90 nw
rect 12035 63 12085 64
rect 199 56 329 62
rect 199 50 251 56
rect 303 50 329 56
rect 199 16 211 50
rect 245 16 251 50
rect 317 16 329 50
rect 199 10 251 16
tri 226 -8 244 10 ne
rect 244 4 251 10
rect 303 10 329 16
rect 441 56 495 62
rect 303 4 310 10
rect 244 -8 310 4
tri 310 -8 328 10 nw
rect 493 4 495 56
rect 552 56 898 62
rect 3317 56 3369 62
rect 3901 56 4031 62
rect 552 50 846 56
rect 552 16 564 50
rect 598 16 636 50
rect 670 16 708 50
rect 742 16 780 50
rect 814 16 846 50
rect 552 10 846 16
rect 441 -8 495 4
tri 821 -8 839 10 ne
rect 839 4 846 10
rect 3248 50 3317 56
rect 3369 50 3666 56
rect 3248 16 3260 50
rect 3294 16 3317 50
rect 3369 16 3404 50
rect 3438 16 3476 50
rect 3510 16 3548 50
rect 3582 16 3620 50
rect 3654 16 3666 50
rect 3248 10 3317 16
rect 839 -8 898 4
tri 3292 -8 3310 10 ne
rect 3310 4 3317 10
rect 3369 10 3666 16
rect 3711 50 3841 56
rect 3763 16 3795 50
rect 3829 16 3841 50
rect 3369 4 3376 10
rect 3310 -8 3376 4
tri 3376 -8 3394 10 nw
rect 3763 10 3841 16
rect 3953 50 4031 56
rect 3953 16 3985 50
rect 4019 16 4031 50
rect 3763 -2 3770 10
rect 3711 -8 3770 -2
tri 3770 -8 3788 10 nw
rect 3953 10 4031 16
rect 4403 56 4533 62
rect 4403 50 4455 56
rect 4507 50 4533 56
rect 4403 16 4415 50
rect 4449 16 4455 50
rect 4521 16 4533 50
rect 4403 10 4455 16
rect 3953 4 3972 10
rect 3901 -8 3972 4
tri 3972 -8 3990 10 nw
tri 4430 -8 4448 10 ne
rect 4448 4 4455 10
rect 4507 10 4533 16
rect 4645 56 4699 62
rect 4507 4 4514 10
rect 4448 -8 4514 4
tri 4514 -8 4532 10 nw
rect 4697 4 4699 56
rect 4741 56 5160 62
rect 4741 50 5050 56
rect 5102 50 5160 56
rect 4741 16 4753 50
rect 4787 16 4825 50
rect 4859 16 4897 50
rect 4931 16 4969 50
rect 5003 16 5041 50
rect 5102 16 5113 50
rect 5147 16 5160 50
rect 4741 10 5050 16
rect 4645 -8 4699 4
tri 5025 -8 5043 10 ne
rect 5043 4 5050 10
rect 5102 10 5160 16
rect 7525 56 7882 62
rect 7525 50 7830 56
rect 7525 16 7537 50
rect 7571 16 7609 50
rect 7643 16 7681 50
rect 7715 16 7753 50
rect 7787 16 7825 50
rect 7525 10 7830 16
rect 5102 4 5109 10
rect 5043 -8 5109 4
tri 5109 -8 5127 10 nw
tri 7805 -8 7823 10 ne
rect 7823 4 7830 10
rect 7915 10 7921 62
rect 7973 10 7985 62
rect 8037 10 8045 62
rect 8105 10 8111 62
rect 8163 10 8175 62
rect 8227 10 8235 62
rect 8607 56 8737 62
rect 8607 50 8659 56
rect 8711 50 8737 56
rect 8607 16 8619 50
rect 8653 16 8659 50
rect 8725 16 8737 50
rect 8607 10 8659 16
rect 7823 -8 7882 4
tri 8634 -8 8652 10 ne
rect 8652 4 8659 10
rect 8711 10 8737 16
rect 8783 56 8901 62
rect 8783 50 8849 56
rect 8783 16 8789 50
rect 8823 16 8849 50
rect 8711 4 8730 10
tri 8730 4 8736 10 nw
rect 8783 4 8849 16
rect 8945 56 9363 62
tri 12122 56 12128 62 se
rect 12128 56 12249 62
rect 8945 50 9254 56
rect 9306 50 9363 56
rect 8945 16 8957 50
rect 8991 16 9029 50
rect 9063 16 9101 50
rect 9135 16 9173 50
rect 9207 16 9245 50
rect 9306 16 9317 50
rect 9351 16 9363 50
rect 12035 26 12085 27
tri 12025 16 12034 25 se
rect 12034 16 12086 25
rect 8945 10 9254 16
rect 8652 -8 8718 4
tri 8718 -8 8730 4 nw
rect 8783 -8 8901 4
tri 9229 -8 9247 10 ne
rect 9247 4 9254 10
rect 9306 10 9363 16
tri 12019 10 12025 16 se
rect 12025 10 12086 16
rect 9306 4 9321 10
rect 9247 0 9321 4
tri 9321 0 9331 10 nw
tri 12009 0 12019 10 se
rect 12019 0 12086 10
rect 12119 10 12128 56
rect 12180 50 12249 56
rect 12180 16 12203 50
rect 12237 16 12249 50
tri 12119 1 12128 10 ne
rect 12180 4 12249 16
rect 9247 -2 9319 0
tri 9319 -2 9321 0 nw
rect 9247 -8 9313 -2
tri 9313 -8 9319 -2 nw
rect 11657 -8 11964 0
tri 244 -15 251 -8 ne
tri 303 -15 310 -8 nw
rect 251 -66 303 -60
rect 493 -60 495 -8
tri 839 -15 846 -8 ne
rect 441 -68 495 -60
tri 3310 -15 3317 -8 ne
rect 846 -66 898 -60
tri 3369 -15 3376 -8 nw
rect 3711 -14 3763 -8
rect 3317 -66 3369 -60
tri 3763 -15 3770 -8 nw
rect 3953 -15 3965 -8
tri 3965 -15 3972 -8 nw
tri 4448 -15 4455 -8 ne
rect 3953 -22 3958 -15
tri 3958 -22 3965 -15 nw
tri 3953 -27 3958 -22 nw
rect 3901 -66 3953 -60
tri 4507 -15 4514 -8 nw
rect 4455 -66 4507 -60
rect 4697 -60 4699 -8
tri 5043 -15 5050 -8 ne
rect 3711 -72 3763 -66
rect 4645 -68 4699 -60
tri 5102 -15 5109 -8 nw
tri 7823 -15 7830 -8 ne
rect 5050 -66 5102 -60
tri 8652 -15 8659 -8 ne
rect 7830 -66 7882 -60
tri 8711 -15 8718 -8 nw
rect 8659 -66 8711 -60
rect 8783 -60 8849 -8
tri 9247 -15 9254 -8 ne
rect 8783 -66 8901 -60
tri 9306 -15 9313 -8 nw
rect 11657 -42 11669 -8
rect 11703 -42 11741 -8
rect 11775 -42 11813 -8
rect 11847 -42 11885 -8
rect 11919 -42 11957 -8
rect 11657 -52 11964 -42
rect 12016 -52 12028 0
rect 12080 -52 12086 0
rect 12128 -8 12249 4
rect 9254 -66 9306 -60
rect 12180 -60 12249 -8
rect 12128 -66 12249 -60
rect 12303 56 12361 62
rect 12303 4 12309 56
rect 12303 -8 12361 4
rect 12303 -60 12309 -8
rect 12303 -66 12361 -60
<< rmetal1 >>
rect 11866 2311 11868 2312
rect 11904 2311 11906 2312
rect 11866 2261 11867 2311
rect 11905 2261 11906 2311
rect 11866 2260 11868 2261
rect 11904 2260 11906 2261
rect 186 786 188 787
rect 224 786 226 787
rect 186 736 187 786
rect 225 736 226 786
rect 303 786 305 787
rect 186 735 188 736
rect 224 735 226 736
rect 303 660 304 786
rect 303 659 305 660
rect 341 786 343 787
rect 342 660 343 786
rect 341 659 343 660
rect 401 786 403 787
rect 439 786 441 787
rect 401 660 402 786
rect 440 660 441 786
rect 518 786 520 787
rect 518 736 519 786
rect 518 735 520 736
rect 556 786 558 787
rect 557 736 558 786
rect 556 735 558 736
rect 401 659 403 660
rect 439 659 441 660
rect 3646 786 3648 787
rect 3646 736 3647 786
rect 3646 735 3648 736
rect 3684 786 3686 787
rect 3685 736 3686 786
rect 3763 786 3765 787
rect 3801 786 3803 787
rect 3684 735 3686 736
rect 3763 660 3764 786
rect 3802 660 3803 786
rect 3763 659 3765 660
rect 3801 659 3803 660
rect 3861 786 3863 787
rect 3861 660 3862 786
rect 3861 659 3863 660
rect 3899 786 3901 787
rect 3900 660 3901 786
rect 3978 786 3980 787
rect 4016 786 4018 787
rect 3978 736 3979 786
rect 4017 736 4018 786
rect 3978 735 3980 736
rect 4016 735 4018 736
rect 3899 659 3901 660
rect 4390 786 4392 787
rect 4428 786 4430 787
rect 4390 736 4391 786
rect 4429 736 4430 786
rect 4507 786 4509 787
rect 4390 735 4392 736
rect 4428 735 4430 736
rect 4507 660 4508 786
rect 4507 659 4509 660
rect 4545 786 4547 787
rect 4546 660 4547 786
rect 4545 659 4547 660
rect 4605 786 4607 787
rect 4643 786 4645 787
rect 4605 660 4606 786
rect 4644 660 4645 786
rect 4722 786 4724 787
rect 4722 736 4723 786
rect 4722 735 4724 736
rect 4760 786 4762 787
rect 4761 736 4762 786
rect 4760 735 4762 736
rect 4605 659 4607 660
rect 4643 659 4645 660
rect 7850 786 7852 787
rect 7850 736 7851 786
rect 7850 735 7852 736
rect 7888 786 7890 787
rect 7889 736 7890 786
rect 7967 786 7969 787
rect 8005 786 8007 787
rect 7888 735 7890 736
rect 7967 660 7968 786
rect 8006 660 8007 786
rect 7967 659 7969 660
rect 8005 659 8007 660
rect 8065 786 8067 787
rect 8065 660 8066 786
rect 8065 659 8067 660
rect 8103 786 8105 787
rect 8104 660 8105 786
rect 8182 786 8184 787
rect 8220 786 8222 787
rect 8182 736 8183 786
rect 8221 736 8222 786
rect 8182 735 8184 736
rect 8220 735 8222 736
rect 8103 659 8105 660
rect 8594 786 8596 787
rect 8632 786 8634 787
rect 8594 736 8595 786
rect 8633 736 8634 786
rect 8711 786 8713 787
rect 8594 735 8596 736
rect 8632 735 8634 736
rect 8711 660 8712 786
rect 8711 659 8713 660
rect 8749 786 8751 787
rect 8750 660 8751 786
rect 8749 659 8751 660
rect 8809 786 8811 787
rect 8847 786 8849 787
rect 8809 660 8810 786
rect 8848 660 8849 786
rect 8926 786 8928 787
rect 8926 736 8927 786
rect 8926 735 8928 736
rect 8964 786 8966 787
rect 8965 736 8966 786
rect 8964 735 8966 736
rect 8809 659 8811 660
rect 8847 659 8849 660
rect 12054 786 12056 787
rect 12054 736 12055 786
rect 12054 735 12056 736
rect 12092 786 12094 787
rect 12093 736 12094 786
rect 12171 786 12173 787
rect 12209 786 12211 787
rect 12092 735 12094 736
rect 12171 660 12172 786
rect 12210 660 12211 786
rect 12171 659 12173 660
rect 12209 659 12211 660
rect 12269 786 12271 787
rect 12269 660 12270 786
rect 12269 659 12271 660
rect 12307 786 12309 787
rect 12308 660 12309 786
rect 12386 786 12388 787
rect 12424 786 12426 787
rect 12386 736 12387 786
rect 12425 736 12426 786
rect 12386 735 12388 736
rect 12424 735 12426 736
rect 12307 659 12309 660
rect 12034 64 12086 65
rect 12034 63 12035 64
rect 12085 63 12086 64
rect 12034 26 12035 27
rect 12085 26 12086 27
rect 12034 25 12086 26
<< via1 >>
rect 846 2330 898 2382
rect 846 2266 898 2318
rect 3323 2260 3375 2312
rect 3387 2260 3439 2312
rect 4980 2260 5032 2312
rect 5044 2260 5096 2312
rect 7760 2260 7812 2312
rect 7824 2260 7876 2312
rect 9184 2260 9236 2312
rect 9248 2260 9300 2312
rect 11964 2260 12016 2312
rect 12028 2260 12080 2312
rect 251 729 303 781
rect 251 665 303 717
rect 441 729 493 781
rect 441 665 493 717
rect 3711 729 3763 781
rect 3711 665 3763 717
rect 3901 729 3953 781
rect 3901 665 3953 717
rect 4455 729 4507 781
rect 4455 665 4507 717
rect 4645 729 4697 781
rect 4645 665 4697 717
rect 7915 729 7967 781
rect 7915 665 7967 717
rect 8105 729 8157 781
rect 8105 665 8157 717
rect 8659 729 8711 781
rect 8659 665 8711 717
rect 8849 729 8901 781
rect 8849 665 8901 717
rect 12119 729 12171 781
rect 12119 665 12171 717
rect 12309 729 12361 781
rect 12309 665 12361 717
rect 12214 518 12266 536
rect 12214 484 12250 518
rect 12250 484 12266 518
rect 251 50 303 56
rect 251 16 283 50
rect 283 16 303 50
rect 251 4 303 16
rect 441 50 493 56
rect 441 16 455 50
rect 455 16 489 50
rect 489 16 493 50
rect 441 4 493 16
rect 846 50 898 56
rect 846 16 852 50
rect 852 16 886 50
rect 886 16 898 50
rect 846 4 898 16
rect 3317 50 3369 56
rect 3317 16 3332 50
rect 3332 16 3366 50
rect 3366 16 3369 50
rect 3317 4 3369 16
rect 3711 16 3723 50
rect 3723 16 3757 50
rect 3757 16 3763 50
rect 3711 -2 3763 16
rect 3901 50 3953 56
rect 3901 16 3913 50
rect 3913 16 3947 50
rect 3947 16 3953 50
rect 3901 4 3953 16
rect 4455 50 4507 56
rect 4455 16 4487 50
rect 4487 16 4507 50
rect 4455 4 4507 16
rect 4645 50 4697 56
rect 4645 16 4659 50
rect 4659 16 4693 50
rect 4693 16 4697 50
rect 4645 4 4697 16
rect 5050 50 5102 56
rect 5050 16 5075 50
rect 5075 16 5102 50
rect 5050 4 5102 16
rect 7830 50 7882 56
rect 7830 16 7859 50
rect 7859 16 7882 50
rect 7830 4 7882 16
rect 7921 50 7973 62
rect 7921 16 7927 50
rect 7927 16 7961 50
rect 7961 16 7973 50
rect 7921 10 7973 16
rect 7985 50 8037 62
rect 7985 16 7999 50
rect 7999 16 8033 50
rect 8033 16 8037 50
rect 7985 10 8037 16
rect 8111 50 8163 62
rect 8111 16 8117 50
rect 8117 16 8151 50
rect 8151 16 8163 50
rect 8111 10 8163 16
rect 8175 50 8227 62
rect 8175 16 8189 50
rect 8189 16 8223 50
rect 8223 16 8227 50
rect 8175 10 8227 16
rect 8659 50 8711 56
rect 8659 16 8691 50
rect 8691 16 8711 50
rect 8659 4 8711 16
rect 8849 50 8901 56
rect 8849 16 8861 50
rect 8861 16 8895 50
rect 8895 16 8901 50
rect 8849 4 8901 16
rect 9254 50 9306 56
rect 9254 16 9279 50
rect 9279 16 9306 50
rect 9254 4 9306 16
rect 12128 50 12180 56
rect 12128 16 12131 50
rect 12131 16 12165 50
rect 12165 16 12180 50
rect 12128 4 12180 16
rect 11964 -8 12016 0
rect 251 -60 303 -8
rect 441 -22 493 -8
rect 441 -56 455 -22
rect 455 -56 489 -22
rect 489 -56 493 -22
rect 441 -60 493 -56
rect 846 -60 898 -8
rect 3317 -60 3369 -8
rect 3711 -66 3763 -14
rect 3901 -60 3953 -8
rect 4455 -60 4507 -8
rect 4645 -22 4697 -8
rect 4645 -56 4659 -22
rect 4659 -56 4693 -22
rect 4693 -56 4697 -22
rect 4645 -60 4697 -56
rect 5050 -60 5102 -8
rect 7830 -60 7882 -8
rect 8659 -60 8711 -8
rect 8849 -60 8901 -8
rect 9254 -60 9306 -8
rect 11964 -42 11991 -8
rect 11991 -42 12016 -8
rect 11964 -52 12016 -42
rect 12028 -8 12080 0
rect 12028 -42 12029 -8
rect 12029 -42 12063 -8
rect 12063 -42 12080 -8
rect 12028 -52 12080 -42
rect 12128 -60 12180 -8
rect 12309 51 12361 56
rect 12309 17 12315 51
rect 12315 17 12349 51
rect 12349 17 12361 51
rect 12309 4 12361 17
rect 12309 -21 12361 -8
rect 12309 -55 12315 -21
rect 12315 -55 12349 -21
rect 12349 -55 12361 -21
rect 12309 -60 12361 -55
<< metal2 >>
rect 846 2382 898 2388
rect 846 2318 898 2330
rect 251 781 303 787
rect 251 717 303 729
rect 251 56 303 665
rect 251 -8 303 4
rect 251 -66 303 -60
rect 441 781 493 787
rect 441 717 493 729
rect 441 56 493 665
rect 441 -8 493 4
rect 441 -66 493 -60
rect 846 56 898 2266
rect 3317 2260 3323 2312
rect 3375 2260 3387 2312
rect 3439 2260 3445 2312
rect 4974 2260 4980 2312
rect 5032 2260 5044 2312
rect 5096 2260 5102 2312
rect 7754 2260 7760 2312
rect 7812 2260 7824 2312
rect 7876 2260 7882 2312
rect 9178 2260 9184 2312
rect 9236 2260 9248 2312
rect 9300 2260 9306 2312
rect 11958 2260 11964 2312
rect 12016 2260 12028 2312
rect 12080 2260 12086 2312
tri 3312 1950 3317 1955 se
rect 3317 1950 3369 2260
tri 3369 2235 3394 2260 nw
tri 5025 2235 5050 2260 ne
tri 3303 1941 3312 1950 se
rect 3312 1941 3355 1950
rect 1461 1049 1491 1079
rect 2713 1049 2743 1079
rect 3303 613 3355 1941
tri 3355 1936 3369 1950 nw
rect 3711 781 3763 787
rect 3711 717 3763 729
tri 3303 606 3310 613 ne
rect 3310 606 3355 613
tri 3355 606 3369 620 sw
tri 3310 599 3317 606 ne
rect 846 -8 898 4
rect 846 -66 898 -60
rect 3317 56 3369 606
rect 3317 -8 3369 4
rect 3317 -66 3369 -60
rect 3711 50 3763 665
rect 3711 -14 3763 -2
rect 3901 781 3953 787
rect 3901 717 3953 729
rect 3901 56 3953 665
rect 3901 -8 3953 4
rect 3901 -66 3953 -60
rect 4455 781 4507 787
rect 4455 717 4507 729
rect 4455 56 4507 665
rect 4455 -8 4507 4
rect 4455 -66 4507 -60
rect 4645 781 4697 787
rect 4645 717 4697 729
rect 4645 56 4697 665
rect 4645 -8 4697 4
rect 4645 -66 4697 -60
rect 5050 56 5102 2260
tri 7805 2235 7830 2260 ne
rect 5665 1049 5694 1079
rect 6917 1049 6947 1079
rect 5050 -8 5102 4
rect 5050 -66 5102 -60
rect 7830 56 7882 2260
tri 9229 2235 9254 2260 ne
rect 7915 781 7967 787
rect 7915 717 7967 729
rect 7915 62 7967 665
rect 8105 781 8157 787
rect 8105 717 8157 729
tri 7967 62 7992 87 sw
rect 8105 62 8157 665
rect 8659 781 8711 787
rect 8659 717 8711 729
tri 8157 62 8182 87 sw
rect 7915 10 7921 62
rect 7973 10 7985 62
rect 8037 10 8043 62
rect 8105 10 8111 62
rect 8163 10 8175 62
rect 8227 10 8233 62
rect 8659 56 8711 665
rect 7830 -8 7882 4
rect 7830 -66 7882 -60
rect 8659 -8 8711 4
rect 8659 -66 8711 -60
rect 8849 781 8901 787
rect 8849 717 8901 729
rect 8849 56 8901 665
rect 8849 -8 8901 4
rect 8849 -66 8901 -60
rect 9254 56 9306 2260
tri 12009 2235 12034 2260 ne
rect 9869 1049 9899 1079
rect 11121 1049 11151 1079
rect 9254 -8 9306 4
rect 12034 0 12086 2260
rect 12119 781 12171 787
rect 12119 717 12171 729
rect 12119 62 12171 665
rect 12309 781 12361 787
rect 12309 717 12361 729
rect 12214 536 12266 659
rect 12214 478 12266 484
tri 12171 62 12180 71 sw
rect 12119 56 12180 62
rect 12119 10 12128 56
tri 12119 4 12125 10 ne
rect 12125 4 12128 10
tri 12125 1 12128 4 ne
rect 11958 -52 11964 0
rect 12016 -52 12028 0
rect 12080 -52 12086 0
rect 12128 -8 12180 4
rect 9254 -66 9306 -60
rect 12128 -66 12180 -60
rect 12309 56 12361 665
rect 12309 -8 12361 4
rect 12309 -66 12361 -60
rect 3711 -72 3763 -66
<< comment >>
rect 12807 -10 12996 2319
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_0
timestamp 1701704242
transform 0 -1 8895 -1 0 50
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_1
timestamp 1701704242
transform 1 0 12315 0 -1 51
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1701704242
transform 0 -1 489 -1 0 50
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1701704242
transform 0 -1 4693 -1 0 50
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1701704242
transform -1 0 12284 0 1 484
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_3
timestamp 1701704242
transform -1 0 8725 0 1 16
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_4
timestamp 1701704242
transform -1 0 4521 0 1 16
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_5
timestamp 1701704242
transform -1 0 317 0 1 16
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_6
timestamp 1701704242
transform 0 1 12563 1 0 332
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_7
timestamp 1701704242
transform 0 -1 8425 1 0 332
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_8
timestamp 1701704242
transform 0 -1 4221 1 0 332
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_9
timestamp 1701704242
transform 0 -1 17 1 0 332
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_10
timestamp 1701704242
transform 0 -1 15017 1 0 332
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_11
timestamp 1701704242
transform 1 0 12131 0 -1 50
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_12
timestamp 1701704242
transform 1 0 8117 0 1 16
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_13
timestamp 1701704242
transform 1 0 7927 0 1 16
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_14
timestamp 1701704242
transform 1 0 3723 0 1 16
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_15
timestamp 1701704242
transform 1 0 3913 0 1 16
box 0 0 1 1
use L1M1_CDNS_52468879185193  L1M1_CDNS_52468879185193_0
timestamp 1701704242
transform -1 0 7859 0 1 16
box 0 0 1 1
use L1M1_CDNS_52468879185193  L1M1_CDNS_52468879185193_1
timestamp 1701704242
transform 1 0 564 0 -1 50
box 0 0 1 1
use L1M1_CDNS_52468879185308  L1M1_CDNS_52468879185308_0
timestamp 1701704242
transform -1 0 12063 0 1 -42
box 0 0 1 1
use L1M1_CDNS_52468879185308  L1M1_CDNS_52468879185308_1
timestamp 1701704242
transform -1 0 5147 0 1 16
box 0 0 1 1
use L1M1_CDNS_52468879185308  L1M1_CDNS_52468879185308_2
timestamp 1701704242
transform -1 0 9351 0 1 16
box 0 0 1 1
use L1M1_CDNS_52468879185308  L1M1_CDNS_52468879185308_3
timestamp 1701704242
transform 1 0 3260 0 1 16
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_0
timestamp 1701704242
transform 0 -1 3953 -1 0 787
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_1
timestamp 1701704242
transform 0 -1 303 -1 0 787
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_2
timestamp 1701704242
transform 0 -1 493 -1 0 787
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_3
timestamp 1701704242
transform 0 -1 3763 -1 0 56
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_4
timestamp 1701704242
transform 0 -1 7967 -1 0 787
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_5
timestamp 1701704242
transform 0 -1 8157 -1 0 787
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_6
timestamp 1701704242
transform 0 -1 4697 -1 0 787
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_7
timestamp 1701704242
transform 0 -1 8901 -1 0 787
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_8
timestamp 1701704242
transform 0 -1 8711 -1 0 787
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_9
timestamp 1701704242
transform 0 -1 12171 -1 0 787
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_10
timestamp 1701704242
transform 0 -1 12361 -1 0 787
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_11
timestamp 1701704242
transform 0 -1 4507 -1 0 787
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_12
timestamp 1701704242
transform 0 -1 3953 -1 0 62
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_13
timestamp 1701704242
transform 0 -1 3763 -1 0 787
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_14
timestamp 1701704242
transform -1 0 8233 0 1 10
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_15
timestamp 1701704242
transform -1 0 8043 0 1 10
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_16
timestamp 1701704242
transform -1 0 5102 0 -1 2312
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_17
timestamp 1701704242
transform -1 0 7882 0 -1 2312
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_18
timestamp 1701704242
transform -1 0 9306 0 -1 2312
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_19
timestamp 1701704242
transform -1 0 12086 0 -1 2312
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_20
timestamp 1701704242
transform 0 1 12309 1 0 -66
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_21
timestamp 1701704242
transform 0 1 12128 1 0 -66
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_22
timestamp 1701704242
transform 0 1 846 1 0 2260
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_23
timestamp 1701704242
transform 0 1 5050 1 0 -66
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_24
timestamp 1701704242
transform 0 1 9254 1 0 -66
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_25
timestamp 1701704242
transform 0 -1 3369 1 0 -66
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_26
timestamp 1701704242
transform 0 -1 493 1 0 -66
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_27
timestamp 1701704242
transform 0 -1 8711 1 0 -66
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_28
timestamp 1701704242
transform 0 -1 8901 1 0 -66
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_29
timestamp 1701704242
transform 0 -1 4507 1 0 -66
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_30
timestamp 1701704242
transform 0 -1 4697 1 0 -66
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_31
timestamp 1701704242
transform 0 -1 898 1 0 -66
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_32
timestamp 1701704242
transform 0 -1 303 1 0 -66
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_33
timestamp 1701704242
transform 0 -1 7882 1 0 -66
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_34
timestamp 1701704242
transform 1 0 11958 0 -1 0
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_35
timestamp 1701704242
transform 1 0 3317 0 -1 2312
box 0 0 1 1
use M1M2_CDNS_52468879185970  M1M2_CDNS_52468879185970_0
timestamp 1701704242
transform 0 -1 12266 -1 0 542
box 0 0 1 1
use sky130_fd_io__sio_com_ctl_ls  sky130_fd_io__sio_com_ctl_ls_0
timestamp 1701704242
transform -1 0 6306 0 1 0
box -91 0 2150 2319
use sky130_fd_io__sio_com_ctl_ls  sky130_fd_io__sio_com_ctl_ls_1
timestamp 1701704242
transform -1 0 2102 0 1 0
box -91 0 2150 2319
use sky130_fd_io__sio_com_ctl_ls  sky130_fd_io__sio_com_ctl_ls_2
timestamp 1701704242
transform -1 0 10510 0 1 0
box -91 0 2150 2319
use sky130_fd_io__sio_com_ctl_ls  sky130_fd_io__sio_com_ctl_ls_3
timestamp 1701704242
transform 1 0 2102 0 1 0
box -91 0 2150 2319
use sky130_fd_io__sio_com_ctl_ls  sky130_fd_io__sio_com_ctl_ls_4
timestamp 1701704242
transform 1 0 6306 0 1 0
box -91 0 2150 2319
use sky130_fd_io__sio_com_ctl_ls  sky130_fd_io__sio_com_ctl_ls_5
timestamp 1701704242
transform 1 0 10510 0 1 0
box -91 0 2150 2319
use sky130_fd_io__tk_em1o_CDNS_52468879185315  sky130_fd_io__tk_em1o_CDNS_52468879185315_0
timestamp 1701704242
transform 0 1 12034 -1 0 117
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185315  sky130_fd_io__tk_em1o_CDNS_52468879185315_1
timestamp 1701704242
transform -1 0 9018 0 1 735
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185315  sky130_fd_io__tk_em1o_CDNS_52468879185315_2
timestamp 1701704242
transform -1 0 4814 0 1 735
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185315  sky130_fd_io__tk_em1o_CDNS_52468879185315_3
timestamp 1701704242
transform -1 0 610 0 1 735
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185315  sky130_fd_io__tk_em1o_CDNS_52468879185315_4
timestamp 1701704242
transform 1 0 12002 0 1 735
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185315  sky130_fd_io__tk_em1o_CDNS_52468879185315_5
timestamp 1701704242
transform 1 0 7798 0 1 735
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185315  sky130_fd_io__tk_em1o_CDNS_52468879185315_6
timestamp 1701704242
transform 1 0 3594 0 1 735
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185338  sky130_fd_io__tk_em1o_CDNS_52468879185338_0
timestamp 1701704242
transform -1 0 8803 0 1 659
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185338  sky130_fd_io__tk_em1o_CDNS_52468879185338_1
timestamp 1701704242
transform -1 0 4599 0 1 659
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185338  sky130_fd_io__tk_em1o_CDNS_52468879185338_2
timestamp 1701704242
transform -1 0 395 0 1 659
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185338  sky130_fd_io__tk_em1o_CDNS_52468879185338_3
timestamp 1701704242
transform 1 0 8013 0 1 659
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185338  sky130_fd_io__tk_em1o_CDNS_52468879185338_4
timestamp 1701704242
transform 1 0 12217 0 1 659
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185338  sky130_fd_io__tk_em1o_CDNS_52468879185338_5
timestamp 1701704242
transform 1 0 3809 0 1 659
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185314  sky130_fd_io__tk_em1s_CDNS_52468879185314_0
timestamp 1701704242
transform -1 0 278 0 1 735
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185314  sky130_fd_io__tk_em1s_CDNS_52468879185314_1
timestamp 1701704242
transform -1 0 8686 0 1 735
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185314  sky130_fd_io__tk_em1s_CDNS_52468879185314_2
timestamp 1701704242
transform -1 0 4482 0 1 735
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185314  sky130_fd_io__tk_em1s_CDNS_52468879185314_3
timestamp 1701704242
transform -1 0 11958 0 -1 2312
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185314  sky130_fd_io__tk_em1s_CDNS_52468879185314_4
timestamp 1701704242
transform 1 0 8130 0 1 735
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185314  sky130_fd_io__tk_em1s_CDNS_52468879185314_5
timestamp 1701704242
transform 1 0 12334 0 1 735
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185314  sky130_fd_io__tk_em1s_CDNS_52468879185314_6
timestamp 1701704242
transform 1 0 3926 0 1 735
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_524688791851189  sky130_fd_io__tk_em1s_CDNS_524688791851189_0
timestamp 1701704242
transform -1 0 493 0 1 659
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_524688791851189  sky130_fd_io__tk_em1s_CDNS_524688791851189_1
timestamp 1701704242
transform -1 0 8901 0 1 659
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_524688791851189  sky130_fd_io__tk_em1s_CDNS_524688791851189_2
timestamp 1701704242
transform -1 0 4697 0 1 659
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_524688791851189  sky130_fd_io__tk_em1s_CDNS_524688791851189_3
timestamp 1701704242
transform 1 0 7915 0 1 659
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_524688791851189  sky130_fd_io__tk_em1s_CDNS_524688791851189_4
timestamp 1701704242
transform 1 0 12119 0 1 659
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_524688791851189  sky130_fd_io__tk_em1s_CDNS_524688791851189_5
timestamp 1701704242
transform 1 0 3711 0 1 659
box 0 0 1 1
<< labels >>
flabel comment s 464 125 464 125 0 FreeSans 200 90 0 0 dm_st_h<0>
flabel comment s 265 27 265 27 0 FreeSans 200 180 0 0 dm_rst_h<0>
flabel comment s 12337 607 12337 607 0 FreeSans 400 180 0 0 od_i_h
flabel comment s 5098 608 5098 608 0 FreeSans 400 180 0 0 od_i_h
flabel comment s 3766 33 3766 33 0 FreeSans 200 0 0 0 dm_st_h<1>
flabel comment s 968 604 968 604 0 FreeSans 400 180 0 0 od_i_h
flabel comment s 10964 2288 10964 2288 0 FreeSans 400 180 0 0 hld_i_h_n
flabel comment s 7337 530 7337 530 0 FreeSans 200 0 0 0 dm_st_h<0>
flabel comment s 7384 -96 7384 -96 0 FreeSans 200 0 0 0 dm_rst_h<0>
flabel comment s 115 1066 115 1066 0 FreeSans 400 180 0 0 dm<0>
flabel comment s 4088 1066 4088 1066 0 FreeSans 400 180 0 0 dm<1>
flabel comment s 4320 1066 4320 1066 0 FreeSans 400 180 0 0 dm<2>
flabel comment s 8292 1066 8292 1066 0 FreeSans 400 180 0 0 ibuf_sel
flabel comment s 8524 1066 8524 1066 0 FreeSans 400 180 0 0 vtrip_sel
flabel comment s 12496 1066 12496 1066 0 FreeSans 400 180 0 0 sio_diff_hyst_en
flabel comment s 11094 1072 11094 1072 0 FreeSans 200 180 0 0 sio_diff_hyst_sel_h
flabel comment s 10848 680 10848 680 0 FreeSans 400 180 0 0 sio_diff_hyst_sel_h_n
flabel comment s 10046 1064 10046 1064 0 FreeSans 400 180 0 0 vtrip_sel_h
flabel comment s 10172 680 10172 680 0 FreeSans 400 180 0 0 vtrip_sel_h_n
flabel comment s 6644 680 6644 680 0 FreeSans 400 180 0 0 ibuf_sel_h_n
flabel comment s 6735 1075 6735 1075 0 FreeSans 400 180 0 0 ibuf_sel_h
flabel comment s 5679 1064 5679 1064 0 FreeSans 400 180 0 0 dm_h<2>
flabel comment s 5968 680 5968 680 0 FreeSans 400 180 0 0 dm_h_n<2>
flabel comment s 2440 680 2440 680 0 FreeSans 400 180 0 0 dm_h_n<1>
flabel comment s 2728 1064 2728 1064 0 FreeSans 400 180 0 0 dm_h<1>
flabel comment s 1476 1064 1476 1064 0 FreeSans 400 180 0 0 dm_h<0>
flabel comment s 1764 680 1764 680 0 FreeSans 400 180 0 0 dm_h_n<0>
flabel metal1 s 12553 1469 12594 1515 3 FreeSans 520 0 0 0 hld_i_vpwr
port 2 nsew
flabel metal1 s 12479 1049 12513 1083 0 FreeSans 400 0 0 0 inp_dis
port 8 nsew
flabel metal1 s 0 320 34 450 3 FreeSans 400 0 0 0 vgnd
port 3 nsew
flabel metal1 s 10155 663 10189 697 0 FreeSans 400 0 0 0 vtrip_sel_h_n
port 4 nsew
flabel metal1 s 8507 1049 8541 1083 0 FreeSans 400 0 0 0 vtrip_sel
port 5 nsew
flabel metal1 s 185 1884 219 2086 3 FreeSans 400 0 0 0 vpwr
port 6 nsew
flabel metal1 s 0 1239 34 1441 3 FreeSans 400 0 0 0 vgnd
port 3 nsew
flabel metal1 s 0 90 34 292 3 FreeSans 400 0 0 0 vcc_io
port 7 nsew
flabel metal1 s 11828 585 11862 619 0 FreeSans 400 0 0 0 od_i_h
port 9 nsew
flabel metal1 s 10831 663 10865 697 0 FreeSans 400 0 0 0 inp_dis_h_n
port 10 nsew
flabel metal1 s 6627 663 6660 697 0 FreeSans 400 0 0 0 ibuf_sel_h_n
port 11 nsew
flabel metal1 s 8275 1049 8309 1083 0 FreeSans 400 0 0 0 ibuf_sel
port 12 nsew
flabel metal1 s 803 2266 841 2300 0 FreeSans 400 0 0 0 hld_i_h_n
port 13 nsew
flabel metal1 s 5951 663 5985 697 0 FreeSans 400 0 0 0 dm_h_n<2>
port 14 nsew
flabel metal1 s 2423 663 2457 697 0 FreeSans 400 0 0 0 dm_h_n<1>
port 15 nsew
flabel metal1 s 1747 663 1781 697 0 FreeSans 400 0 0 0 dm_h_n<0>
port 16 nsew
flabel metal1 s 4303 1049 4337 1083 0 FreeSans 400 0 0 0 dm<2>
port 17 nsew
flabel metal1 s 4071 1049 4105 1083 0 FreeSans 400 0 0 0 dm<1>
port 18 nsew
flabel metal1 s 98 1049 132 1083 0 FreeSans 400 0 0 0 dm<0>
port 19 nsew
flabel metal1 s 14966 320 15000 450 3 FreeSans 400 180 0 0 vgnd
port 3 nsew
flabel metal2 s 8871 179 8871 179 0 FreeSans 200 90 0 0 trip_sel_st_h
flabel metal2 s 8683 181 8683 181 0 FreeSans 200 90 0 0 trip_sel_rst_h
flabel metal2 s 12136 195 12136 195 0 FreeSans 200 90 0 0 sio_diff_hyst_en_st_h
flabel metal2 s 12335 195 12335 195 0 FreeSans 200 90 0 0 sio_diff_hyst_en_rst_h
flabel metal2 s 9869 1049 9899 1079 3 FreeSans 400 0 0 0 vtrip_sel_h
port 20 nsew
flabel metal2 s 11121 1049 11151 1079 0 FreeSans 400 0 0 0 inp_dis_h
port 21 nsew
flabel metal2 s 6917 1049 6947 1079 0 FreeSans 400 0 0 0 ibuf_sel_h
port 22 nsew
flabel metal2 s 5665 1049 5694 1079 0 FreeSans 400 0 0 0 dm_h<2>
port 23 nsew
flabel metal2 s 2713 1049 2743 1079 0 FreeSans 400 0 0 0 dm_h<1>
port 24 nsew
flabel metal2 s 1461 1049 1491 1079 0 FreeSans 400 0 0 0 dm_h<0>
port 25 nsew
<< properties >>
string GDS_END 85304966
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85272974
string path 105.100 55.400 105.100 38.400 
<< end >>
