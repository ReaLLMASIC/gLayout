magic
tech sky130A
timestamp 1701704242
<< properties >>
string GDS_END 30606002
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 30602734
<< end >>
