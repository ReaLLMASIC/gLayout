magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -823 2514 -323 3754
rect 91 3611 3610 3754
rect 91 3588 3619 3611
rect 91 2514 1322 3588
rect 1341 3548 2287 3588
rect 2683 3548 3619 3588
rect 1341 3332 3619 3548
rect 1341 2514 2287 3332
rect 2683 2879 3619 3332
rect 1634 2479 2287 2514
rect 4058 2188 4630 3720
rect 5030 2188 5652 3720
rect 6123 3391 6824 3433
rect 6123 2515 6832 3391
<< pwell >>
rect -32378 -9661 -27010 4370
rect 3912 3780 5798 3866
rect 207 1927 551 2263
rect 3912 2128 3998 3780
rect 4696 2128 4968 3780
rect 5712 3351 5798 3780
rect 5712 2596 6018 3351
rect 5712 2128 5798 2596
rect 3912 2042 5798 2128
rect 2663 1927 3389 1933
rect -258 875 1925 1927
rect 2663 1912 3673 1927
rect 2097 1275 3673 1912
rect 3912 1885 4196 2042
rect 3852 1633 4196 1885
rect 2097 1260 3389 1275
rect 117 853 1925 875
rect 2663 853 3389 1260
rect 117 767 3420 853
rect 117 4 2169 767
rect 2663 453 3236 767
<< mvnmos >>
rect 5852 3152 5992 3272
rect 5852 2976 5992 3096
rect 5852 2675 5992 2795
rect -176 901 -16 1901
rect 171 901 331 1901
rect 387 901 547 1901
rect 603 901 763 1901
rect 819 901 979 1901
rect 1035 901 1195 1901
rect 1251 901 1411 1901
rect 1467 901 1627 1901
rect 1683 901 1843 1901
rect 2176 1286 2276 1886
rect 2459 1286 2559 1886
rect 2742 907 2842 1907
rect 2898 907 2998 1907
rect 3054 907 3154 1907
rect 3210 907 3310 1907
rect 3491 1301 3591 1901
rect 2742 479 2842 679
rect 2898 479 2998 679
rect 3054 479 3154 679
<< mvpmos >>
rect -701 2580 -601 3580
rect -545 2580 -445 3580
rect 213 2580 313 3580
rect 369 2580 469 3580
rect 661 2580 761 3580
rect 817 2580 917 3580
rect 1100 2580 1200 3580
rect 1460 2580 1560 3580
rect 1753 2545 1853 3545
rect 1909 2545 2009 3545
rect 2065 2545 2165 3545
rect 2356 3398 2456 3482
rect 2512 3398 2612 3482
rect 2802 2945 2902 3545
rect 3085 2945 3185 3545
rect 3241 2945 3341 3545
rect 3397 2945 3497 3545
rect 4289 2545 4389 3545
rect 5261 3288 5421 3488
rect 5261 2782 5421 2982
rect 6190 3152 6390 3272
rect 6458 3152 6658 3272
rect 6190 2976 6390 3096
rect 6458 2976 6658 3096
rect 6190 2675 6390 2795
rect 6458 2675 6658 2795
<< mvnnmos >>
rect 289 2037 469 2237
rect 3934 1659 4114 1859
rect 143 449 2143 629
rect 143 86 2143 266
<< mvndiff >>
rect -31524 -8719 -31512 -8685
rect -31478 -8719 -31466 -8685
rect -31524 -8739 -31466 -8719
rect -29280 -8731 -29268 -8697
rect -29234 -8731 -29222 -8697
rect -29280 -8739 -29222 -8731
rect 233 2225 289 2237
rect 233 2191 244 2225
rect 278 2191 289 2225
rect 233 2157 289 2191
rect 233 2123 244 2157
rect 278 2123 289 2157
rect 233 2089 289 2123
rect 233 2055 244 2089
rect 278 2055 289 2089
rect 233 2037 289 2055
rect 469 2225 525 2237
rect 469 2191 480 2225
rect 514 2191 525 2225
rect 469 2157 525 2191
rect 469 2123 480 2157
rect 514 2123 525 2157
rect 469 2089 525 2123
rect 469 2055 480 2089
rect 514 2055 525 2089
rect 5852 3317 5992 3325
rect 5852 3283 5878 3317
rect 5912 3283 5946 3317
rect 5980 3283 5992 3317
rect 5852 3272 5992 3283
rect 5852 3096 5992 3152
rect 5852 2965 5992 2976
rect 5852 2931 5878 2965
rect 5912 2931 5946 2965
rect 5980 2931 5992 2965
rect 5852 2923 5992 2931
rect 5852 2840 5992 2848
rect 5852 2806 5878 2840
rect 5912 2806 5946 2840
rect 5980 2806 5992 2840
rect 5852 2795 5992 2806
rect 5852 2664 5992 2675
rect 5852 2630 5878 2664
rect 5912 2630 5946 2664
rect 5980 2630 5992 2664
rect 5852 2622 5992 2630
rect 469 2037 525 2055
rect -232 1831 -176 1901
rect -232 1797 -221 1831
rect -187 1797 -176 1831
rect -232 1763 -176 1797
rect -232 1729 -221 1763
rect -187 1729 -176 1763
rect -232 1695 -176 1729
rect -232 1661 -221 1695
rect -187 1661 -176 1695
rect -232 1627 -176 1661
rect -232 1593 -221 1627
rect -187 1593 -176 1627
rect -232 1559 -176 1593
rect -232 1525 -221 1559
rect -187 1525 -176 1559
rect -232 1491 -176 1525
rect -232 1457 -221 1491
rect -187 1457 -176 1491
rect -232 1423 -176 1457
rect -232 1389 -221 1423
rect -187 1389 -176 1423
rect -232 1355 -176 1389
rect -232 1321 -221 1355
rect -187 1321 -176 1355
rect -232 1287 -176 1321
rect -232 1253 -221 1287
rect -187 1253 -176 1287
rect -232 1219 -176 1253
rect -232 1185 -221 1219
rect -187 1185 -176 1219
rect -232 1151 -176 1185
rect -232 1117 -221 1151
rect -187 1117 -176 1151
rect -232 1083 -176 1117
rect -232 1049 -221 1083
rect -187 1049 -176 1083
rect -232 1015 -176 1049
rect -232 981 -221 1015
rect -187 981 -176 1015
rect -232 947 -176 981
rect -232 913 -221 947
rect -187 913 -176 947
rect -232 901 -176 913
rect -16 1831 40 1901
rect -16 1797 -5 1831
rect 29 1797 40 1831
rect -16 1763 40 1797
rect -16 1729 -5 1763
rect 29 1729 40 1763
rect -16 1695 40 1729
rect -16 1661 -5 1695
rect 29 1661 40 1695
rect -16 1627 40 1661
rect -16 1593 -5 1627
rect 29 1593 40 1627
rect -16 1559 40 1593
rect -16 1525 -5 1559
rect 29 1525 40 1559
rect -16 1491 40 1525
rect -16 1457 -5 1491
rect 29 1457 40 1491
rect -16 1423 40 1457
rect -16 1389 -5 1423
rect 29 1389 40 1423
rect -16 1355 40 1389
rect -16 1321 -5 1355
rect 29 1321 40 1355
rect -16 1287 40 1321
rect -16 1253 -5 1287
rect 29 1253 40 1287
rect -16 1219 40 1253
rect -16 1185 -5 1219
rect 29 1185 40 1219
rect -16 1151 40 1185
rect -16 1117 -5 1151
rect 29 1117 40 1151
rect -16 1083 40 1117
rect -16 1049 -5 1083
rect 29 1049 40 1083
rect -16 1015 40 1049
rect -16 981 -5 1015
rect 29 981 40 1015
rect -16 947 40 981
rect -16 913 -5 947
rect 29 913 40 947
rect -16 901 40 913
rect 115 1831 171 1901
rect 115 1797 126 1831
rect 160 1797 171 1831
rect 115 1763 171 1797
rect 115 1729 126 1763
rect 160 1729 171 1763
rect 115 1695 171 1729
rect 115 1661 126 1695
rect 160 1661 171 1695
rect 115 1627 171 1661
rect 115 1593 126 1627
rect 160 1593 171 1627
rect 115 1559 171 1593
rect 115 1525 126 1559
rect 160 1525 171 1559
rect 115 1491 171 1525
rect 115 1457 126 1491
rect 160 1457 171 1491
rect 115 1423 171 1457
rect 115 1389 126 1423
rect 160 1389 171 1423
rect 115 1355 171 1389
rect 115 1321 126 1355
rect 160 1321 171 1355
rect 115 1287 171 1321
rect 115 1253 126 1287
rect 160 1253 171 1287
rect 115 1219 171 1253
rect 115 1185 126 1219
rect 160 1185 171 1219
rect 115 1151 171 1185
rect 115 1117 126 1151
rect 160 1117 171 1151
rect 115 1083 171 1117
rect 115 1049 126 1083
rect 160 1049 171 1083
rect 115 1015 171 1049
rect 115 981 126 1015
rect 160 981 171 1015
rect 115 947 171 981
rect 115 913 126 947
rect 160 913 171 947
rect 115 901 171 913
rect 331 1831 387 1901
rect 331 1797 342 1831
rect 376 1797 387 1831
rect 331 1763 387 1797
rect 331 1729 342 1763
rect 376 1729 387 1763
rect 331 1695 387 1729
rect 331 1661 342 1695
rect 376 1661 387 1695
rect 331 1627 387 1661
rect 331 1593 342 1627
rect 376 1593 387 1627
rect 331 1559 387 1593
rect 331 1525 342 1559
rect 376 1525 387 1559
rect 331 1491 387 1525
rect 331 1457 342 1491
rect 376 1457 387 1491
rect 331 1423 387 1457
rect 331 1389 342 1423
rect 376 1389 387 1423
rect 331 1355 387 1389
rect 331 1321 342 1355
rect 376 1321 387 1355
rect 331 1287 387 1321
rect 331 1253 342 1287
rect 376 1253 387 1287
rect 331 1219 387 1253
rect 331 1185 342 1219
rect 376 1185 387 1219
rect 331 1151 387 1185
rect 331 1117 342 1151
rect 376 1117 387 1151
rect 331 1083 387 1117
rect 331 1049 342 1083
rect 376 1049 387 1083
rect 331 1015 387 1049
rect 331 981 342 1015
rect 376 981 387 1015
rect 331 947 387 981
rect 331 913 342 947
rect 376 913 387 947
rect 331 901 387 913
rect 547 1831 603 1901
rect 547 1797 558 1831
rect 592 1797 603 1831
rect 547 1763 603 1797
rect 547 1729 558 1763
rect 592 1729 603 1763
rect 547 1695 603 1729
rect 547 1661 558 1695
rect 592 1661 603 1695
rect 547 1627 603 1661
rect 547 1593 558 1627
rect 592 1593 603 1627
rect 547 1559 603 1593
rect 547 1525 558 1559
rect 592 1525 603 1559
rect 547 1491 603 1525
rect 547 1457 558 1491
rect 592 1457 603 1491
rect 547 1423 603 1457
rect 547 1389 558 1423
rect 592 1389 603 1423
rect 547 1355 603 1389
rect 547 1321 558 1355
rect 592 1321 603 1355
rect 547 1287 603 1321
rect 547 1253 558 1287
rect 592 1253 603 1287
rect 547 1219 603 1253
rect 547 1185 558 1219
rect 592 1185 603 1219
rect 547 1151 603 1185
rect 547 1117 558 1151
rect 592 1117 603 1151
rect 547 1083 603 1117
rect 547 1049 558 1083
rect 592 1049 603 1083
rect 547 1015 603 1049
rect 547 981 558 1015
rect 592 981 603 1015
rect 547 947 603 981
rect 547 913 558 947
rect 592 913 603 947
rect 547 901 603 913
rect 763 1831 819 1901
rect 763 1797 774 1831
rect 808 1797 819 1831
rect 763 1763 819 1797
rect 763 1729 774 1763
rect 808 1729 819 1763
rect 763 1695 819 1729
rect 763 1661 774 1695
rect 808 1661 819 1695
rect 763 1627 819 1661
rect 763 1593 774 1627
rect 808 1593 819 1627
rect 763 1559 819 1593
rect 763 1525 774 1559
rect 808 1525 819 1559
rect 763 1491 819 1525
rect 763 1457 774 1491
rect 808 1457 819 1491
rect 763 1423 819 1457
rect 763 1389 774 1423
rect 808 1389 819 1423
rect 763 1355 819 1389
rect 763 1321 774 1355
rect 808 1321 819 1355
rect 763 1287 819 1321
rect 763 1253 774 1287
rect 808 1253 819 1287
rect 763 1219 819 1253
rect 763 1185 774 1219
rect 808 1185 819 1219
rect 763 1151 819 1185
rect 763 1117 774 1151
rect 808 1117 819 1151
rect 763 1083 819 1117
rect 763 1049 774 1083
rect 808 1049 819 1083
rect 763 1015 819 1049
rect 763 981 774 1015
rect 808 981 819 1015
rect 763 947 819 981
rect 763 913 774 947
rect 808 913 819 947
rect 763 901 819 913
rect 979 1831 1035 1901
rect 979 1797 990 1831
rect 1024 1797 1035 1831
rect 979 1763 1035 1797
rect 979 1729 990 1763
rect 1024 1729 1035 1763
rect 979 1695 1035 1729
rect 979 1661 990 1695
rect 1024 1661 1035 1695
rect 979 1627 1035 1661
rect 979 1593 990 1627
rect 1024 1593 1035 1627
rect 979 1559 1035 1593
rect 979 1525 990 1559
rect 1024 1525 1035 1559
rect 979 1491 1035 1525
rect 979 1457 990 1491
rect 1024 1457 1035 1491
rect 979 1423 1035 1457
rect 979 1389 990 1423
rect 1024 1389 1035 1423
rect 979 1355 1035 1389
rect 979 1321 990 1355
rect 1024 1321 1035 1355
rect 979 1287 1035 1321
rect 979 1253 990 1287
rect 1024 1253 1035 1287
rect 979 1219 1035 1253
rect 979 1185 990 1219
rect 1024 1185 1035 1219
rect 979 1151 1035 1185
rect 979 1117 990 1151
rect 1024 1117 1035 1151
rect 979 1083 1035 1117
rect 979 1049 990 1083
rect 1024 1049 1035 1083
rect 979 1015 1035 1049
rect 979 981 990 1015
rect 1024 981 1035 1015
rect 979 947 1035 981
rect 979 913 990 947
rect 1024 913 1035 947
rect 979 901 1035 913
rect 1195 1831 1251 1901
rect 1195 1797 1206 1831
rect 1240 1797 1251 1831
rect 1195 1763 1251 1797
rect 1195 1729 1206 1763
rect 1240 1729 1251 1763
rect 1195 1695 1251 1729
rect 1195 1661 1206 1695
rect 1240 1661 1251 1695
rect 1195 1627 1251 1661
rect 1195 1593 1206 1627
rect 1240 1593 1251 1627
rect 1195 1559 1251 1593
rect 1195 1525 1206 1559
rect 1240 1525 1251 1559
rect 1195 1491 1251 1525
rect 1195 1457 1206 1491
rect 1240 1457 1251 1491
rect 1195 1423 1251 1457
rect 1195 1389 1206 1423
rect 1240 1389 1251 1423
rect 1195 1355 1251 1389
rect 1195 1321 1206 1355
rect 1240 1321 1251 1355
rect 1195 1287 1251 1321
rect 1195 1253 1206 1287
rect 1240 1253 1251 1287
rect 1195 1219 1251 1253
rect 1195 1185 1206 1219
rect 1240 1185 1251 1219
rect 1195 1151 1251 1185
rect 1195 1117 1206 1151
rect 1240 1117 1251 1151
rect 1195 1083 1251 1117
rect 1195 1049 1206 1083
rect 1240 1049 1251 1083
rect 1195 1015 1251 1049
rect 1195 981 1206 1015
rect 1240 981 1251 1015
rect 1195 947 1251 981
rect 1195 913 1206 947
rect 1240 913 1251 947
rect 1195 901 1251 913
rect 1411 1831 1467 1901
rect 1411 1797 1422 1831
rect 1456 1797 1467 1831
rect 1411 1763 1467 1797
rect 1411 1729 1422 1763
rect 1456 1729 1467 1763
rect 1411 1695 1467 1729
rect 1411 1661 1422 1695
rect 1456 1661 1467 1695
rect 1411 1627 1467 1661
rect 1411 1593 1422 1627
rect 1456 1593 1467 1627
rect 1411 1559 1467 1593
rect 1411 1525 1422 1559
rect 1456 1525 1467 1559
rect 1411 1491 1467 1525
rect 1411 1457 1422 1491
rect 1456 1457 1467 1491
rect 1411 1423 1467 1457
rect 1411 1389 1422 1423
rect 1456 1389 1467 1423
rect 1411 1355 1467 1389
rect 1411 1321 1422 1355
rect 1456 1321 1467 1355
rect 1411 1287 1467 1321
rect 1411 1253 1422 1287
rect 1456 1253 1467 1287
rect 1411 1219 1467 1253
rect 1411 1185 1422 1219
rect 1456 1185 1467 1219
rect 1411 1151 1467 1185
rect 1411 1117 1422 1151
rect 1456 1117 1467 1151
rect 1411 1083 1467 1117
rect 1411 1049 1422 1083
rect 1456 1049 1467 1083
rect 1411 1015 1467 1049
rect 1411 981 1422 1015
rect 1456 981 1467 1015
rect 1411 947 1467 981
rect 1411 913 1422 947
rect 1456 913 1467 947
rect 1411 901 1467 913
rect 1627 1831 1683 1901
rect 1627 1797 1638 1831
rect 1672 1797 1683 1831
rect 1627 1763 1683 1797
rect 1627 1729 1638 1763
rect 1672 1729 1683 1763
rect 1627 1695 1683 1729
rect 1627 1661 1638 1695
rect 1672 1661 1683 1695
rect 1627 1627 1683 1661
rect 1627 1593 1638 1627
rect 1672 1593 1683 1627
rect 1627 1559 1683 1593
rect 1627 1525 1638 1559
rect 1672 1525 1683 1559
rect 1627 1491 1683 1525
rect 1627 1457 1638 1491
rect 1672 1457 1683 1491
rect 1627 1423 1683 1457
rect 1627 1389 1638 1423
rect 1672 1389 1683 1423
rect 1627 1355 1683 1389
rect 1627 1321 1638 1355
rect 1672 1321 1683 1355
rect 1627 1287 1683 1321
rect 1627 1253 1638 1287
rect 1672 1253 1683 1287
rect 1627 1219 1683 1253
rect 1627 1185 1638 1219
rect 1672 1185 1683 1219
rect 1627 1151 1683 1185
rect 1627 1117 1638 1151
rect 1672 1117 1683 1151
rect 1627 1083 1683 1117
rect 1627 1049 1638 1083
rect 1672 1049 1683 1083
rect 1627 1015 1683 1049
rect 1627 981 1638 1015
rect 1672 981 1683 1015
rect 1627 947 1683 981
rect 1627 913 1638 947
rect 1672 913 1683 947
rect 1627 901 1683 913
rect 1843 1831 1899 1901
rect 1843 1797 1854 1831
rect 1888 1797 1899 1831
rect 1843 1763 1899 1797
rect 1843 1729 1854 1763
rect 1888 1729 1899 1763
rect 1843 1695 1899 1729
rect 1843 1661 1854 1695
rect 1888 1661 1899 1695
rect 1843 1627 1899 1661
rect 1843 1593 1854 1627
rect 1888 1593 1899 1627
rect 1843 1559 1899 1593
rect 1843 1525 1854 1559
rect 1888 1525 1899 1559
rect 1843 1491 1899 1525
rect 1843 1457 1854 1491
rect 1888 1457 1899 1491
rect 1843 1423 1899 1457
rect 1843 1389 1854 1423
rect 1888 1389 1899 1423
rect 1843 1355 1899 1389
rect 1843 1321 1854 1355
rect 1888 1321 1899 1355
rect 1843 1287 1899 1321
rect 1843 1253 1854 1287
rect 1888 1253 1899 1287
rect 2123 1808 2176 1886
rect 2123 1774 2131 1808
rect 2165 1774 2176 1808
rect 2123 1740 2176 1774
rect 2123 1706 2131 1740
rect 2165 1706 2176 1740
rect 2123 1672 2176 1706
rect 2123 1638 2131 1672
rect 2165 1638 2176 1672
rect 2123 1604 2176 1638
rect 2123 1570 2131 1604
rect 2165 1570 2176 1604
rect 2123 1536 2176 1570
rect 2123 1502 2131 1536
rect 2165 1502 2176 1536
rect 2123 1468 2176 1502
rect 2123 1434 2131 1468
rect 2165 1434 2176 1468
rect 2123 1400 2176 1434
rect 2123 1366 2131 1400
rect 2165 1366 2176 1400
rect 2123 1332 2176 1366
rect 2123 1298 2131 1332
rect 2165 1298 2176 1332
rect 2123 1286 2176 1298
rect 2276 1808 2332 1886
rect 2276 1774 2287 1808
rect 2321 1774 2332 1808
rect 2276 1740 2332 1774
rect 2276 1706 2287 1740
rect 2321 1706 2332 1740
rect 2276 1672 2332 1706
rect 2276 1638 2287 1672
rect 2321 1638 2332 1672
rect 2276 1604 2332 1638
rect 2276 1570 2287 1604
rect 2321 1570 2332 1604
rect 2276 1536 2332 1570
rect 2276 1502 2287 1536
rect 2321 1502 2332 1536
rect 2276 1468 2332 1502
rect 2276 1434 2287 1468
rect 2321 1434 2332 1468
rect 2276 1400 2332 1434
rect 2276 1366 2287 1400
rect 2321 1366 2332 1400
rect 2276 1332 2332 1366
rect 2276 1298 2287 1332
rect 2321 1298 2332 1332
rect 2276 1286 2332 1298
rect 2406 1808 2459 1886
rect 2406 1774 2414 1808
rect 2448 1774 2459 1808
rect 2406 1740 2459 1774
rect 2406 1706 2414 1740
rect 2448 1706 2459 1740
rect 2406 1672 2459 1706
rect 2406 1638 2414 1672
rect 2448 1638 2459 1672
rect 2406 1604 2459 1638
rect 2406 1570 2414 1604
rect 2448 1570 2459 1604
rect 2406 1536 2459 1570
rect 2406 1502 2414 1536
rect 2448 1502 2459 1536
rect 2406 1468 2459 1502
rect 2406 1434 2414 1468
rect 2448 1434 2459 1468
rect 2406 1400 2459 1434
rect 2406 1366 2414 1400
rect 2448 1366 2459 1400
rect 2406 1332 2459 1366
rect 2406 1298 2414 1332
rect 2448 1298 2459 1332
rect 2406 1286 2459 1298
rect 2559 1808 2615 1886
rect 2559 1774 2570 1808
rect 2604 1774 2615 1808
rect 2559 1740 2615 1774
rect 2559 1706 2570 1740
rect 2604 1706 2615 1740
rect 2559 1672 2615 1706
rect 2559 1638 2570 1672
rect 2604 1638 2615 1672
rect 2559 1604 2615 1638
rect 2559 1570 2570 1604
rect 2604 1570 2615 1604
rect 2559 1536 2615 1570
rect 2559 1502 2570 1536
rect 2604 1502 2615 1536
rect 2559 1468 2615 1502
rect 2559 1434 2570 1468
rect 2604 1434 2615 1468
rect 2559 1400 2615 1434
rect 2559 1366 2570 1400
rect 2604 1366 2615 1400
rect 2559 1332 2615 1366
rect 2559 1298 2570 1332
rect 2604 1298 2615 1332
rect 2559 1286 2615 1298
rect 2689 1837 2742 1907
rect 2689 1803 2697 1837
rect 2731 1803 2742 1837
rect 2689 1769 2742 1803
rect 2689 1735 2697 1769
rect 2731 1735 2742 1769
rect 2689 1701 2742 1735
rect 2689 1667 2697 1701
rect 2731 1667 2742 1701
rect 2689 1633 2742 1667
rect 2689 1599 2697 1633
rect 2731 1599 2742 1633
rect 2689 1565 2742 1599
rect 2689 1531 2697 1565
rect 2731 1531 2742 1565
rect 2689 1497 2742 1531
rect 2689 1463 2697 1497
rect 2731 1463 2742 1497
rect 2689 1429 2742 1463
rect 2689 1395 2697 1429
rect 2731 1395 2742 1429
rect 2689 1361 2742 1395
rect 2689 1327 2697 1361
rect 2731 1327 2742 1361
rect 2689 1293 2742 1327
rect 2689 1259 2697 1293
rect 2731 1259 2742 1293
rect 1843 1219 1899 1253
rect 1843 1185 1854 1219
rect 1888 1185 1899 1219
rect 1843 1151 1899 1185
rect 1843 1117 1854 1151
rect 1888 1117 1899 1151
rect 1843 1083 1899 1117
rect 1843 1049 1854 1083
rect 1888 1049 1899 1083
rect 1843 1015 1899 1049
rect 1843 981 1854 1015
rect 1888 981 1899 1015
rect 1843 947 1899 981
rect 1843 913 1854 947
rect 1888 913 1899 947
rect 1843 901 1899 913
rect 2689 1225 2742 1259
rect 2689 1191 2697 1225
rect 2731 1191 2742 1225
rect 2689 1157 2742 1191
rect 2689 1123 2697 1157
rect 2731 1123 2742 1157
rect 2689 1089 2742 1123
rect 2689 1055 2697 1089
rect 2731 1055 2742 1089
rect 2689 1021 2742 1055
rect 2689 987 2697 1021
rect 2731 987 2742 1021
rect 2689 953 2742 987
rect 2689 919 2697 953
rect 2731 919 2742 953
rect 2689 907 2742 919
rect 2842 1837 2898 1907
rect 2842 1803 2853 1837
rect 2887 1803 2898 1837
rect 2842 1769 2898 1803
rect 2842 1735 2853 1769
rect 2887 1735 2898 1769
rect 2842 1701 2898 1735
rect 2842 1667 2853 1701
rect 2887 1667 2898 1701
rect 2842 1633 2898 1667
rect 2842 1599 2853 1633
rect 2887 1599 2898 1633
rect 2842 1565 2898 1599
rect 2842 1531 2853 1565
rect 2887 1531 2898 1565
rect 2842 1497 2898 1531
rect 2842 1463 2853 1497
rect 2887 1463 2898 1497
rect 2842 1429 2898 1463
rect 2842 1395 2853 1429
rect 2887 1395 2898 1429
rect 2842 1361 2898 1395
rect 2842 1327 2853 1361
rect 2887 1327 2898 1361
rect 2842 1293 2898 1327
rect 2842 1259 2853 1293
rect 2887 1259 2898 1293
rect 2842 1225 2898 1259
rect 2842 1191 2853 1225
rect 2887 1191 2898 1225
rect 2842 1157 2898 1191
rect 2842 1123 2853 1157
rect 2887 1123 2898 1157
rect 2842 1089 2898 1123
rect 2842 1055 2853 1089
rect 2887 1055 2898 1089
rect 2842 1021 2898 1055
rect 2842 987 2853 1021
rect 2887 987 2898 1021
rect 2842 953 2898 987
rect 2842 919 2853 953
rect 2887 919 2898 953
rect 2842 907 2898 919
rect 2998 1837 3054 1907
rect 2998 1803 3009 1837
rect 3043 1803 3054 1837
rect 2998 1769 3054 1803
rect 2998 1735 3009 1769
rect 3043 1735 3054 1769
rect 2998 1701 3054 1735
rect 2998 1667 3009 1701
rect 3043 1667 3054 1701
rect 2998 1633 3054 1667
rect 2998 1599 3009 1633
rect 3043 1599 3054 1633
rect 2998 1565 3054 1599
rect 2998 1531 3009 1565
rect 3043 1531 3054 1565
rect 2998 1497 3054 1531
rect 2998 1463 3009 1497
rect 3043 1463 3054 1497
rect 2998 1429 3054 1463
rect 2998 1395 3009 1429
rect 3043 1395 3054 1429
rect 2998 1361 3054 1395
rect 2998 1327 3009 1361
rect 3043 1327 3054 1361
rect 2998 1293 3054 1327
rect 2998 1259 3009 1293
rect 3043 1259 3054 1293
rect 2998 1225 3054 1259
rect 2998 1191 3009 1225
rect 3043 1191 3054 1225
rect 2998 1157 3054 1191
rect 2998 1123 3009 1157
rect 3043 1123 3054 1157
rect 2998 1089 3054 1123
rect 2998 1055 3009 1089
rect 3043 1055 3054 1089
rect 2998 1021 3054 1055
rect 2998 987 3009 1021
rect 3043 987 3054 1021
rect 2998 953 3054 987
rect 2998 919 3009 953
rect 3043 919 3054 953
rect 2998 907 3054 919
rect 3154 1837 3210 1907
rect 3154 1803 3165 1837
rect 3199 1803 3210 1837
rect 3154 1769 3210 1803
rect 3154 1735 3165 1769
rect 3199 1735 3210 1769
rect 3154 1701 3210 1735
rect 3154 1667 3165 1701
rect 3199 1667 3210 1701
rect 3154 1633 3210 1667
rect 3154 1599 3165 1633
rect 3199 1599 3210 1633
rect 3154 1565 3210 1599
rect 3154 1531 3165 1565
rect 3199 1531 3210 1565
rect 3154 1497 3210 1531
rect 3154 1463 3165 1497
rect 3199 1463 3210 1497
rect 3154 1429 3210 1463
rect 3154 1395 3165 1429
rect 3199 1395 3210 1429
rect 3154 1361 3210 1395
rect 3154 1327 3165 1361
rect 3199 1327 3210 1361
rect 3154 1293 3210 1327
rect 3154 1259 3165 1293
rect 3199 1259 3210 1293
rect 3154 1225 3210 1259
rect 3154 1191 3165 1225
rect 3199 1191 3210 1225
rect 3154 1157 3210 1191
rect 3154 1123 3165 1157
rect 3199 1123 3210 1157
rect 3154 1089 3210 1123
rect 3154 1055 3165 1089
rect 3199 1055 3210 1089
rect 3154 1021 3210 1055
rect 3154 987 3165 1021
rect 3199 987 3210 1021
rect 3154 953 3210 987
rect 3154 919 3165 953
rect 3199 919 3210 953
rect 3154 907 3210 919
rect 3310 1837 3363 1907
rect 3310 1803 3321 1837
rect 3355 1803 3363 1837
rect 3310 1769 3363 1803
rect 3310 1735 3321 1769
rect 3355 1735 3363 1769
rect 3310 1701 3363 1735
rect 3310 1667 3321 1701
rect 3355 1667 3363 1701
rect 3310 1633 3363 1667
rect 3310 1599 3321 1633
rect 3355 1599 3363 1633
rect 3310 1565 3363 1599
rect 3310 1531 3321 1565
rect 3355 1531 3363 1565
rect 3310 1497 3363 1531
rect 3310 1463 3321 1497
rect 3355 1463 3363 1497
rect 3310 1429 3363 1463
rect 3310 1395 3321 1429
rect 3355 1395 3363 1429
rect 3310 1361 3363 1395
rect 3310 1327 3321 1361
rect 3355 1327 3363 1361
rect 3310 1293 3363 1327
rect 3438 1823 3491 1901
rect 3438 1789 3446 1823
rect 3480 1789 3491 1823
rect 3438 1755 3491 1789
rect 3438 1721 3446 1755
rect 3480 1721 3491 1755
rect 3438 1687 3491 1721
rect 3438 1653 3446 1687
rect 3480 1653 3491 1687
rect 3438 1619 3491 1653
rect 3438 1585 3446 1619
rect 3480 1585 3491 1619
rect 3438 1551 3491 1585
rect 3438 1517 3446 1551
rect 3480 1517 3491 1551
rect 3438 1483 3491 1517
rect 3438 1449 3446 1483
rect 3480 1449 3491 1483
rect 3438 1415 3491 1449
rect 3438 1381 3446 1415
rect 3480 1381 3491 1415
rect 3438 1347 3491 1381
rect 3438 1313 3446 1347
rect 3480 1313 3491 1347
rect 3438 1301 3491 1313
rect 3591 1823 3647 1901
rect 3591 1789 3602 1823
rect 3636 1789 3647 1823
rect 3591 1755 3647 1789
rect 3591 1721 3602 1755
rect 3636 1721 3647 1755
rect 3591 1687 3647 1721
rect 3591 1653 3602 1687
rect 3636 1653 3647 1687
rect 3878 1841 3934 1859
rect 3878 1807 3889 1841
rect 3923 1807 3934 1841
rect 3878 1773 3934 1807
rect 3878 1739 3889 1773
rect 3923 1739 3934 1773
rect 3878 1705 3934 1739
rect 3878 1671 3889 1705
rect 3923 1671 3934 1705
rect 3878 1659 3934 1671
rect 4114 1841 4170 1859
rect 4114 1807 4125 1841
rect 4159 1807 4170 1841
rect 4114 1773 4170 1807
rect 4114 1739 4125 1773
rect 4159 1739 4170 1773
rect 4114 1705 4170 1739
rect 4114 1671 4125 1705
rect 4159 1671 4170 1705
rect 4114 1659 4170 1671
rect 3591 1619 3647 1653
rect 3591 1585 3602 1619
rect 3636 1585 3647 1619
rect 3591 1551 3647 1585
rect 3591 1517 3602 1551
rect 3636 1517 3647 1551
rect 3591 1483 3647 1517
rect 3591 1449 3602 1483
rect 3636 1449 3647 1483
rect 3591 1415 3647 1449
rect 3591 1381 3602 1415
rect 3636 1381 3647 1415
rect 3591 1347 3647 1381
rect 3591 1313 3602 1347
rect 3636 1313 3647 1347
rect 3591 1301 3647 1313
rect 3310 1259 3321 1293
rect 3355 1259 3363 1293
rect 3310 1225 3363 1259
rect 3310 1191 3321 1225
rect 3355 1191 3363 1225
rect 3310 1157 3363 1191
rect 3310 1123 3321 1157
rect 3355 1123 3363 1157
rect 3310 1089 3363 1123
rect 3310 1055 3321 1089
rect 3355 1055 3363 1089
rect 3310 1021 3363 1055
rect 3310 987 3321 1021
rect 3355 987 3363 1021
rect 3310 953 3363 987
rect 3310 919 3321 953
rect 3355 919 3363 953
rect 3310 907 3363 919
rect 143 674 2143 685
rect 143 640 193 674
rect 227 640 261 674
rect 295 640 329 674
rect 363 640 397 674
rect 431 640 465 674
rect 499 640 533 674
rect 567 640 601 674
rect 635 640 669 674
rect 703 640 737 674
rect 771 640 805 674
rect 839 640 873 674
rect 907 640 941 674
rect 975 640 1009 674
rect 1043 640 1077 674
rect 1111 640 1145 674
rect 1179 640 1213 674
rect 1247 640 1281 674
rect 1315 640 1349 674
rect 1383 640 1417 674
rect 1451 640 1485 674
rect 1519 640 1553 674
rect 1587 640 1621 674
rect 1655 640 1689 674
rect 1723 640 1757 674
rect 1791 640 1825 674
rect 1859 640 1893 674
rect 1927 640 1961 674
rect 1995 640 2029 674
rect 2063 640 2097 674
rect 2131 640 2143 674
rect 143 629 2143 640
rect 2689 667 2742 679
rect 2689 633 2697 667
rect 2731 633 2742 667
rect 2689 599 2742 633
rect 2689 565 2697 599
rect 2731 565 2742 599
rect 2689 531 2742 565
rect 2689 497 2697 531
rect 2731 497 2742 531
rect 2689 479 2742 497
rect 2842 667 2898 679
rect 2842 633 2853 667
rect 2887 633 2898 667
rect 2842 599 2898 633
rect 2842 565 2853 599
rect 2887 565 2898 599
rect 2842 531 2898 565
rect 2842 497 2853 531
rect 2887 497 2898 531
rect 2842 479 2898 497
rect 2998 667 3054 679
rect 2998 633 3009 667
rect 3043 633 3054 667
rect 2998 599 3054 633
rect 2998 565 3009 599
rect 3043 565 3054 599
rect 2998 531 3054 565
rect 2998 497 3009 531
rect 3043 497 3054 531
rect 2998 479 3054 497
rect 3154 667 3210 679
rect 3154 633 3165 667
rect 3199 633 3210 667
rect 3154 599 3210 633
rect 3154 565 3165 599
rect 3199 565 3210 599
rect 3154 531 3210 565
rect 3154 497 3165 531
rect 3199 497 3210 531
rect 3154 479 3210 497
rect 143 438 2143 449
rect 143 404 193 438
rect 227 404 261 438
rect 295 404 329 438
rect 363 404 397 438
rect 431 404 465 438
rect 499 404 533 438
rect 567 404 601 438
rect 635 404 669 438
rect 703 404 737 438
rect 771 404 805 438
rect 839 404 873 438
rect 907 404 941 438
rect 975 404 1009 438
rect 1043 404 1077 438
rect 1111 404 1145 438
rect 1179 404 1213 438
rect 1247 404 1281 438
rect 1315 404 1349 438
rect 1383 404 1417 438
rect 1451 404 1485 438
rect 1519 404 1553 438
rect 1587 404 1621 438
rect 1655 404 1689 438
rect 1723 404 1757 438
rect 1791 404 1825 438
rect 1859 404 1893 438
rect 1927 404 1961 438
rect 1995 404 2029 438
rect 2063 404 2097 438
rect 2131 404 2143 438
rect 143 393 2143 404
rect 143 311 2143 319
rect 143 277 193 311
rect 227 277 261 311
rect 295 277 329 311
rect 363 277 397 311
rect 431 277 465 311
rect 499 277 533 311
rect 567 277 601 311
rect 635 277 669 311
rect 703 277 737 311
rect 771 277 805 311
rect 839 277 873 311
rect 907 277 941 311
rect 975 277 1009 311
rect 1043 277 1077 311
rect 1111 277 1145 311
rect 1179 277 1213 311
rect 1247 277 1281 311
rect 1315 277 1349 311
rect 1383 277 1417 311
rect 1451 277 1485 311
rect 1519 277 1553 311
rect 1587 277 1621 311
rect 1655 277 1689 311
rect 1723 277 1757 311
rect 1791 277 1825 311
rect 1859 277 1893 311
rect 1927 277 1961 311
rect 1995 277 2029 311
rect 2063 277 2097 311
rect 2131 277 2143 311
rect 143 266 2143 277
rect 143 75 2143 86
rect 143 41 193 75
rect 227 41 261 75
rect 295 41 329 75
rect 363 41 397 75
rect 431 41 465 75
rect 499 41 533 75
rect 567 41 601 75
rect 635 41 669 75
rect 703 41 737 75
rect 771 41 805 75
rect 839 41 873 75
rect 907 41 941 75
rect 975 41 1009 75
rect 1043 41 1077 75
rect 1111 41 1145 75
rect 1179 41 1213 75
rect 1247 41 1281 75
rect 1315 41 1349 75
rect 1383 41 1417 75
rect 1451 41 1485 75
rect 1519 41 1553 75
rect 1587 41 1621 75
rect 1655 41 1689 75
rect 1723 41 1757 75
rect 1791 41 1825 75
rect 1859 41 1893 75
rect 1927 41 1961 75
rect 1995 41 2029 75
rect 2063 41 2097 75
rect 2131 41 2143 75
rect 143 30 2143 41
<< mvpdiff >>
rect -757 3510 -701 3580
rect -757 3476 -746 3510
rect -712 3476 -701 3510
rect -757 3442 -701 3476
rect -757 3408 -746 3442
rect -712 3408 -701 3442
rect -757 3374 -701 3408
rect -757 3340 -746 3374
rect -712 3340 -701 3374
rect -757 3306 -701 3340
rect -757 3272 -746 3306
rect -712 3272 -701 3306
rect -757 3238 -701 3272
rect -757 3204 -746 3238
rect -712 3204 -701 3238
rect -757 3170 -701 3204
rect -757 3136 -746 3170
rect -712 3136 -701 3170
rect -757 3102 -701 3136
rect -757 3068 -746 3102
rect -712 3068 -701 3102
rect -757 3034 -701 3068
rect -757 3000 -746 3034
rect -712 3000 -701 3034
rect -757 2966 -701 3000
rect -757 2932 -746 2966
rect -712 2932 -701 2966
rect -757 2898 -701 2932
rect -757 2864 -746 2898
rect -712 2864 -701 2898
rect -757 2830 -701 2864
rect -757 2796 -746 2830
rect -712 2796 -701 2830
rect -757 2762 -701 2796
rect -757 2728 -746 2762
rect -712 2728 -701 2762
rect -757 2694 -701 2728
rect -757 2660 -746 2694
rect -712 2660 -701 2694
rect -757 2626 -701 2660
rect -757 2592 -746 2626
rect -712 2592 -701 2626
rect -757 2580 -701 2592
rect -601 3510 -545 3580
rect -601 3476 -590 3510
rect -556 3476 -545 3510
rect -601 3442 -545 3476
rect -601 3408 -590 3442
rect -556 3408 -545 3442
rect -601 3374 -545 3408
rect -601 3340 -590 3374
rect -556 3340 -545 3374
rect -601 3306 -545 3340
rect -601 3272 -590 3306
rect -556 3272 -545 3306
rect -601 3238 -545 3272
rect -601 3204 -590 3238
rect -556 3204 -545 3238
rect -601 3170 -545 3204
rect -601 3136 -590 3170
rect -556 3136 -545 3170
rect -601 3102 -545 3136
rect -601 3068 -590 3102
rect -556 3068 -545 3102
rect -601 3034 -545 3068
rect -601 3000 -590 3034
rect -556 3000 -545 3034
rect -601 2966 -545 3000
rect -601 2932 -590 2966
rect -556 2932 -545 2966
rect -601 2898 -545 2932
rect -601 2864 -590 2898
rect -556 2864 -545 2898
rect -601 2830 -545 2864
rect -601 2796 -590 2830
rect -556 2796 -545 2830
rect -601 2762 -545 2796
rect -601 2728 -590 2762
rect -556 2728 -545 2762
rect -601 2694 -545 2728
rect -601 2660 -590 2694
rect -556 2660 -545 2694
rect -601 2626 -545 2660
rect -601 2592 -590 2626
rect -556 2592 -545 2626
rect -601 2580 -545 2592
rect -445 3510 -389 3580
rect -445 3476 -434 3510
rect -400 3476 -389 3510
rect -445 3442 -389 3476
rect -445 3408 -434 3442
rect -400 3408 -389 3442
rect -445 3374 -389 3408
rect -445 3340 -434 3374
rect -400 3340 -389 3374
rect -445 3306 -389 3340
rect -445 3272 -434 3306
rect -400 3272 -389 3306
rect -445 3238 -389 3272
rect -445 3204 -434 3238
rect -400 3204 -389 3238
rect -445 3170 -389 3204
rect -445 3136 -434 3170
rect -400 3136 -389 3170
rect -445 3102 -389 3136
rect -445 3068 -434 3102
rect -400 3068 -389 3102
rect -445 3034 -389 3068
rect -445 3000 -434 3034
rect -400 3000 -389 3034
rect -445 2966 -389 3000
rect -445 2932 -434 2966
rect -400 2932 -389 2966
rect -445 2898 -389 2932
rect -445 2864 -434 2898
rect -400 2864 -389 2898
rect -445 2830 -389 2864
rect -445 2796 -434 2830
rect -400 2796 -389 2830
rect -445 2762 -389 2796
rect -445 2728 -434 2762
rect -400 2728 -389 2762
rect -445 2694 -389 2728
rect -445 2660 -434 2694
rect -400 2660 -389 2694
rect -445 2626 -389 2660
rect -445 2592 -434 2626
rect -400 2592 -389 2626
rect -445 2580 -389 2592
rect 157 3510 213 3580
rect 157 3476 168 3510
rect 202 3476 213 3510
rect 157 3442 213 3476
rect 157 3408 168 3442
rect 202 3408 213 3442
rect 157 3374 213 3408
rect 157 3340 168 3374
rect 202 3340 213 3374
rect 157 3306 213 3340
rect 157 3272 168 3306
rect 202 3272 213 3306
rect 157 3238 213 3272
rect 157 3204 168 3238
rect 202 3204 213 3238
rect 157 3170 213 3204
rect 157 3136 168 3170
rect 202 3136 213 3170
rect 157 3102 213 3136
rect 157 3068 168 3102
rect 202 3068 213 3102
rect 157 3034 213 3068
rect 157 3000 168 3034
rect 202 3000 213 3034
rect 157 2966 213 3000
rect 157 2932 168 2966
rect 202 2932 213 2966
rect 157 2898 213 2932
rect 157 2864 168 2898
rect 202 2864 213 2898
rect 157 2830 213 2864
rect 157 2796 168 2830
rect 202 2796 213 2830
rect 157 2762 213 2796
rect 157 2728 168 2762
rect 202 2728 213 2762
rect 157 2694 213 2728
rect 157 2660 168 2694
rect 202 2660 213 2694
rect 157 2626 213 2660
rect 157 2592 168 2626
rect 202 2592 213 2626
rect 157 2580 213 2592
rect 313 3510 369 3580
rect 313 3476 324 3510
rect 358 3476 369 3510
rect 313 3442 369 3476
rect 313 3408 324 3442
rect 358 3408 369 3442
rect 313 3374 369 3408
rect 313 3340 324 3374
rect 358 3340 369 3374
rect 313 3306 369 3340
rect 313 3272 324 3306
rect 358 3272 369 3306
rect 313 3238 369 3272
rect 313 3204 324 3238
rect 358 3204 369 3238
rect 313 3170 369 3204
rect 313 3136 324 3170
rect 358 3136 369 3170
rect 313 3102 369 3136
rect 313 3068 324 3102
rect 358 3068 369 3102
rect 313 3034 369 3068
rect 313 3000 324 3034
rect 358 3000 369 3034
rect 313 2966 369 3000
rect 313 2932 324 2966
rect 358 2932 369 2966
rect 313 2898 369 2932
rect 313 2864 324 2898
rect 358 2864 369 2898
rect 313 2830 369 2864
rect 313 2796 324 2830
rect 358 2796 369 2830
rect 313 2762 369 2796
rect 313 2728 324 2762
rect 358 2728 369 2762
rect 313 2694 369 2728
rect 313 2660 324 2694
rect 358 2660 369 2694
rect 313 2626 369 2660
rect 313 2592 324 2626
rect 358 2592 369 2626
rect 313 2580 369 2592
rect 469 3510 525 3580
rect 469 3476 480 3510
rect 514 3476 525 3510
rect 469 3442 525 3476
rect 469 3408 480 3442
rect 514 3408 525 3442
rect 469 3374 525 3408
rect 469 3340 480 3374
rect 514 3340 525 3374
rect 469 3306 525 3340
rect 469 3272 480 3306
rect 514 3272 525 3306
rect 469 3238 525 3272
rect 469 3204 480 3238
rect 514 3204 525 3238
rect 469 3170 525 3204
rect 469 3136 480 3170
rect 514 3136 525 3170
rect 469 3102 525 3136
rect 469 3068 480 3102
rect 514 3068 525 3102
rect 469 3034 525 3068
rect 469 3000 480 3034
rect 514 3000 525 3034
rect 469 2966 525 3000
rect 469 2932 480 2966
rect 514 2932 525 2966
rect 469 2898 525 2932
rect 469 2864 480 2898
rect 514 2864 525 2898
rect 469 2830 525 2864
rect 469 2796 480 2830
rect 514 2796 525 2830
rect 469 2762 525 2796
rect 469 2728 480 2762
rect 514 2728 525 2762
rect 469 2694 525 2728
rect 469 2660 480 2694
rect 514 2660 525 2694
rect 469 2626 525 2660
rect 469 2592 480 2626
rect 514 2592 525 2626
rect 469 2580 525 2592
rect 605 3510 661 3580
rect 605 3476 616 3510
rect 650 3476 661 3510
rect 605 3442 661 3476
rect 605 3408 616 3442
rect 650 3408 661 3442
rect 605 3374 661 3408
rect 605 3340 616 3374
rect 650 3340 661 3374
rect 605 3306 661 3340
rect 605 3272 616 3306
rect 650 3272 661 3306
rect 605 3238 661 3272
rect 605 3204 616 3238
rect 650 3204 661 3238
rect 605 3170 661 3204
rect 605 3136 616 3170
rect 650 3136 661 3170
rect 605 3102 661 3136
rect 605 3068 616 3102
rect 650 3068 661 3102
rect 605 3034 661 3068
rect 605 3000 616 3034
rect 650 3000 661 3034
rect 605 2966 661 3000
rect 605 2932 616 2966
rect 650 2932 661 2966
rect 605 2898 661 2932
rect 605 2864 616 2898
rect 650 2864 661 2898
rect 605 2830 661 2864
rect 605 2796 616 2830
rect 650 2796 661 2830
rect 605 2762 661 2796
rect 605 2728 616 2762
rect 650 2728 661 2762
rect 605 2694 661 2728
rect 605 2660 616 2694
rect 650 2660 661 2694
rect 605 2626 661 2660
rect 605 2592 616 2626
rect 650 2592 661 2626
rect 605 2580 661 2592
rect 761 3510 817 3580
rect 761 3476 772 3510
rect 806 3476 817 3510
rect 761 3442 817 3476
rect 761 3408 772 3442
rect 806 3408 817 3442
rect 761 3374 817 3408
rect 761 3340 772 3374
rect 806 3340 817 3374
rect 761 3306 817 3340
rect 761 3272 772 3306
rect 806 3272 817 3306
rect 761 3238 817 3272
rect 761 3204 772 3238
rect 806 3204 817 3238
rect 761 3170 817 3204
rect 761 3136 772 3170
rect 806 3136 817 3170
rect 761 3102 817 3136
rect 761 3068 772 3102
rect 806 3068 817 3102
rect 761 3034 817 3068
rect 761 3000 772 3034
rect 806 3000 817 3034
rect 761 2966 817 3000
rect 761 2932 772 2966
rect 806 2932 817 2966
rect 761 2898 817 2932
rect 761 2864 772 2898
rect 806 2864 817 2898
rect 761 2830 817 2864
rect 761 2796 772 2830
rect 806 2796 817 2830
rect 761 2762 817 2796
rect 761 2728 772 2762
rect 806 2728 817 2762
rect 761 2694 817 2728
rect 761 2660 772 2694
rect 806 2660 817 2694
rect 761 2626 817 2660
rect 761 2592 772 2626
rect 806 2592 817 2626
rect 761 2580 817 2592
rect 917 3510 970 3580
rect 917 3476 928 3510
rect 962 3476 970 3510
rect 917 3442 970 3476
rect 917 3408 928 3442
rect 962 3408 970 3442
rect 917 3374 970 3408
rect 917 3340 928 3374
rect 962 3340 970 3374
rect 917 3306 970 3340
rect 917 3272 928 3306
rect 962 3272 970 3306
rect 917 3238 970 3272
rect 917 3204 928 3238
rect 962 3204 970 3238
rect 917 3170 970 3204
rect 917 3136 928 3170
rect 962 3136 970 3170
rect 917 3102 970 3136
rect 917 3068 928 3102
rect 962 3068 970 3102
rect 917 3034 970 3068
rect 917 3000 928 3034
rect 962 3000 970 3034
rect 917 2966 970 3000
rect 917 2932 928 2966
rect 962 2932 970 2966
rect 917 2898 970 2932
rect 917 2864 928 2898
rect 962 2864 970 2898
rect 917 2830 970 2864
rect 917 2796 928 2830
rect 962 2796 970 2830
rect 917 2762 970 2796
rect 917 2728 928 2762
rect 962 2728 970 2762
rect 917 2694 970 2728
rect 917 2660 928 2694
rect 962 2660 970 2694
rect 917 2626 970 2660
rect 917 2592 928 2626
rect 962 2592 970 2626
rect 917 2580 970 2592
rect 1044 3510 1100 3580
rect 1044 3476 1055 3510
rect 1089 3476 1100 3510
rect 1044 3442 1100 3476
rect 1044 3408 1055 3442
rect 1089 3408 1100 3442
rect 1044 3374 1100 3408
rect 1044 3340 1055 3374
rect 1089 3340 1100 3374
rect 1044 3306 1100 3340
rect 1044 3272 1055 3306
rect 1089 3272 1100 3306
rect 1044 3238 1100 3272
rect 1044 3204 1055 3238
rect 1089 3204 1100 3238
rect 1044 3170 1100 3204
rect 1044 3136 1055 3170
rect 1089 3136 1100 3170
rect 1044 3102 1100 3136
rect 1044 3068 1055 3102
rect 1089 3068 1100 3102
rect 1044 3034 1100 3068
rect 1044 3000 1055 3034
rect 1089 3000 1100 3034
rect 1044 2966 1100 3000
rect 1044 2932 1055 2966
rect 1089 2932 1100 2966
rect 1044 2898 1100 2932
rect 1044 2864 1055 2898
rect 1089 2864 1100 2898
rect 1044 2830 1100 2864
rect 1044 2796 1055 2830
rect 1089 2796 1100 2830
rect 1044 2762 1100 2796
rect 1044 2728 1055 2762
rect 1089 2728 1100 2762
rect 1044 2694 1100 2728
rect 1044 2660 1055 2694
rect 1089 2660 1100 2694
rect 1044 2626 1100 2660
rect 1044 2592 1055 2626
rect 1089 2592 1100 2626
rect 1044 2580 1100 2592
rect 1200 3510 1256 3580
rect 1200 3476 1211 3510
rect 1245 3476 1256 3510
rect 1200 3442 1256 3476
rect 1200 3408 1211 3442
rect 1245 3408 1256 3442
rect 1200 3374 1256 3408
rect 1200 3340 1211 3374
rect 1245 3340 1256 3374
rect 1200 3306 1256 3340
rect 1200 3272 1211 3306
rect 1245 3272 1256 3306
rect 1200 3238 1256 3272
rect 1200 3204 1211 3238
rect 1245 3204 1256 3238
rect 1200 3170 1256 3204
rect 1200 3136 1211 3170
rect 1245 3136 1256 3170
rect 1200 3102 1256 3136
rect 1200 3068 1211 3102
rect 1245 3068 1256 3102
rect 1200 3034 1256 3068
rect 1200 3000 1211 3034
rect 1245 3000 1256 3034
rect 1200 2966 1256 3000
rect 1200 2932 1211 2966
rect 1245 2932 1256 2966
rect 1200 2898 1256 2932
rect 1200 2864 1211 2898
rect 1245 2864 1256 2898
rect 1200 2830 1256 2864
rect 1200 2796 1211 2830
rect 1245 2796 1256 2830
rect 1200 2762 1256 2796
rect 1200 2728 1211 2762
rect 1245 2728 1256 2762
rect 1200 2694 1256 2728
rect 1200 2660 1211 2694
rect 1245 2660 1256 2694
rect 1200 2626 1256 2660
rect 1200 2592 1211 2626
rect 1245 2592 1256 2626
rect 1200 2580 1256 2592
rect 1407 3510 1460 3580
rect 1407 3476 1415 3510
rect 1449 3476 1460 3510
rect 1407 3442 1460 3476
rect 1407 3408 1415 3442
rect 1449 3408 1460 3442
rect 1407 3374 1460 3408
rect 1407 3340 1415 3374
rect 1449 3340 1460 3374
rect 1407 3306 1460 3340
rect 1407 3272 1415 3306
rect 1449 3272 1460 3306
rect 1407 3238 1460 3272
rect 1407 3204 1415 3238
rect 1449 3204 1460 3238
rect 1407 3170 1460 3204
rect 1407 3136 1415 3170
rect 1449 3136 1460 3170
rect 1407 3102 1460 3136
rect 1407 3068 1415 3102
rect 1449 3068 1460 3102
rect 1407 3034 1460 3068
rect 1407 3000 1415 3034
rect 1449 3000 1460 3034
rect 1407 2966 1460 3000
rect 1407 2932 1415 2966
rect 1449 2932 1460 2966
rect 1407 2898 1460 2932
rect 1407 2864 1415 2898
rect 1449 2864 1460 2898
rect 1407 2830 1460 2864
rect 1407 2796 1415 2830
rect 1449 2796 1460 2830
rect 1407 2762 1460 2796
rect 1407 2728 1415 2762
rect 1449 2728 1460 2762
rect 1407 2694 1460 2728
rect 1407 2660 1415 2694
rect 1449 2660 1460 2694
rect 1407 2626 1460 2660
rect 1407 2592 1415 2626
rect 1449 2592 1460 2626
rect 1407 2580 1460 2592
rect 1560 3510 1616 3580
rect 1560 3476 1571 3510
rect 1605 3476 1616 3510
rect 1560 3442 1616 3476
rect 1560 3408 1571 3442
rect 1605 3408 1616 3442
rect 1560 3374 1616 3408
rect 1560 3340 1571 3374
rect 1605 3340 1616 3374
rect 1560 3306 1616 3340
rect 1560 3272 1571 3306
rect 1605 3272 1616 3306
rect 1560 3238 1616 3272
rect 1560 3204 1571 3238
rect 1605 3204 1616 3238
rect 1560 3170 1616 3204
rect 1560 3136 1571 3170
rect 1605 3136 1616 3170
rect 1560 3102 1616 3136
rect 1560 3068 1571 3102
rect 1605 3068 1616 3102
rect 1560 3034 1616 3068
rect 1560 3000 1571 3034
rect 1605 3000 1616 3034
rect 1560 2966 1616 3000
rect 1560 2932 1571 2966
rect 1605 2932 1616 2966
rect 1560 2898 1616 2932
rect 1560 2864 1571 2898
rect 1605 2864 1616 2898
rect 1560 2830 1616 2864
rect 1560 2796 1571 2830
rect 1605 2796 1616 2830
rect 1560 2762 1616 2796
rect 1560 2728 1571 2762
rect 1605 2728 1616 2762
rect 1560 2694 1616 2728
rect 1560 2660 1571 2694
rect 1605 2660 1616 2694
rect 1560 2626 1616 2660
rect 1560 2592 1571 2626
rect 1605 2592 1616 2626
rect 1560 2580 1616 2592
rect 1700 3475 1753 3545
rect 1700 3441 1708 3475
rect 1742 3441 1753 3475
rect 1700 3407 1753 3441
rect 1700 3373 1708 3407
rect 1742 3373 1753 3407
rect 1700 3339 1753 3373
rect 1700 3305 1708 3339
rect 1742 3305 1753 3339
rect 1700 3271 1753 3305
rect 1700 3237 1708 3271
rect 1742 3237 1753 3271
rect 1700 3203 1753 3237
rect 1700 3169 1708 3203
rect 1742 3169 1753 3203
rect 1700 3135 1753 3169
rect 1700 3101 1708 3135
rect 1742 3101 1753 3135
rect 1700 3067 1753 3101
rect 1700 3033 1708 3067
rect 1742 3033 1753 3067
rect 1700 2999 1753 3033
rect 1700 2965 1708 2999
rect 1742 2965 1753 2999
rect 1700 2931 1753 2965
rect 1700 2897 1708 2931
rect 1742 2897 1753 2931
rect 1700 2863 1753 2897
rect 1700 2829 1708 2863
rect 1742 2829 1753 2863
rect 1700 2795 1753 2829
rect 1700 2761 1708 2795
rect 1742 2761 1753 2795
rect 1700 2727 1753 2761
rect 1700 2693 1708 2727
rect 1742 2693 1753 2727
rect 1700 2659 1753 2693
rect 1700 2625 1708 2659
rect 1742 2625 1753 2659
rect 1700 2591 1753 2625
rect 1700 2557 1708 2591
rect 1742 2557 1753 2591
rect 1700 2545 1753 2557
rect 1853 3475 1909 3545
rect 1853 3441 1864 3475
rect 1898 3441 1909 3475
rect 1853 3407 1909 3441
rect 1853 3373 1864 3407
rect 1898 3373 1909 3407
rect 1853 3339 1909 3373
rect 1853 3305 1864 3339
rect 1898 3305 1909 3339
rect 1853 3271 1909 3305
rect 1853 3237 1864 3271
rect 1898 3237 1909 3271
rect 1853 3203 1909 3237
rect 1853 3169 1864 3203
rect 1898 3169 1909 3203
rect 1853 3135 1909 3169
rect 1853 3101 1864 3135
rect 1898 3101 1909 3135
rect 1853 3067 1909 3101
rect 1853 3033 1864 3067
rect 1898 3033 1909 3067
rect 1853 2999 1909 3033
rect 1853 2965 1864 2999
rect 1898 2965 1909 2999
rect 1853 2931 1909 2965
rect 1853 2897 1864 2931
rect 1898 2897 1909 2931
rect 1853 2863 1909 2897
rect 1853 2829 1864 2863
rect 1898 2829 1909 2863
rect 1853 2795 1909 2829
rect 1853 2761 1864 2795
rect 1898 2761 1909 2795
rect 1853 2727 1909 2761
rect 1853 2693 1864 2727
rect 1898 2693 1909 2727
rect 1853 2659 1909 2693
rect 1853 2625 1864 2659
rect 1898 2625 1909 2659
rect 1853 2591 1909 2625
rect 1853 2557 1864 2591
rect 1898 2557 1909 2591
rect 1853 2545 1909 2557
rect 2009 3475 2065 3545
rect 2009 3441 2020 3475
rect 2054 3441 2065 3475
rect 2009 3407 2065 3441
rect 2009 3373 2020 3407
rect 2054 3373 2065 3407
rect 2009 3339 2065 3373
rect 2009 3305 2020 3339
rect 2054 3305 2065 3339
rect 2009 3271 2065 3305
rect 2009 3237 2020 3271
rect 2054 3237 2065 3271
rect 2009 3203 2065 3237
rect 2009 3169 2020 3203
rect 2054 3169 2065 3203
rect 2009 3135 2065 3169
rect 2009 3101 2020 3135
rect 2054 3101 2065 3135
rect 2009 3067 2065 3101
rect 2009 3033 2020 3067
rect 2054 3033 2065 3067
rect 2009 2999 2065 3033
rect 2009 2965 2020 2999
rect 2054 2965 2065 2999
rect 2009 2931 2065 2965
rect 2009 2897 2020 2931
rect 2054 2897 2065 2931
rect 2009 2863 2065 2897
rect 2009 2829 2020 2863
rect 2054 2829 2065 2863
rect 2009 2795 2065 2829
rect 2009 2761 2020 2795
rect 2054 2761 2065 2795
rect 2009 2727 2065 2761
rect 2009 2693 2020 2727
rect 2054 2693 2065 2727
rect 2009 2659 2065 2693
rect 2009 2625 2020 2659
rect 2054 2625 2065 2659
rect 2009 2591 2065 2625
rect 2009 2557 2020 2591
rect 2054 2557 2065 2591
rect 2009 2545 2065 2557
rect 2165 3475 2221 3545
rect 2749 3533 2802 3545
rect 2749 3499 2757 3533
rect 2791 3499 2802 3533
rect 2165 3441 2176 3475
rect 2210 3441 2221 3475
rect 2165 3407 2221 3441
rect 2165 3373 2176 3407
rect 2210 3373 2221 3407
rect 2300 3470 2356 3482
rect 2300 3436 2311 3470
rect 2345 3436 2356 3470
rect 2300 3398 2356 3436
rect 2456 3470 2512 3482
rect 2456 3436 2467 3470
rect 2501 3436 2512 3470
rect 2456 3398 2512 3436
rect 2612 3470 2668 3482
rect 2612 3436 2623 3470
rect 2657 3436 2668 3470
rect 2612 3398 2668 3436
rect 2749 3465 2802 3499
rect 2749 3431 2757 3465
rect 2791 3431 2802 3465
rect 2165 3339 2221 3373
rect 2165 3305 2176 3339
rect 2210 3305 2221 3339
rect 2165 3271 2221 3305
rect 2165 3237 2176 3271
rect 2210 3237 2221 3271
rect 2165 3203 2221 3237
rect 2165 3169 2176 3203
rect 2210 3169 2221 3203
rect 2165 3135 2221 3169
rect 2165 3101 2176 3135
rect 2210 3101 2221 3135
rect 2749 3397 2802 3431
rect 2749 3363 2757 3397
rect 2791 3363 2802 3397
rect 2749 3329 2802 3363
rect 2749 3295 2757 3329
rect 2791 3295 2802 3329
rect 2749 3261 2802 3295
rect 2749 3227 2757 3261
rect 2791 3227 2802 3261
rect 2749 3193 2802 3227
rect 2749 3159 2757 3193
rect 2791 3159 2802 3193
rect 2749 3125 2802 3159
rect 2165 3067 2221 3101
rect 2165 3033 2176 3067
rect 2210 3033 2221 3067
rect 2165 2999 2221 3033
rect 2165 2965 2176 2999
rect 2210 2965 2221 2999
rect 2165 2931 2221 2965
rect 2749 3091 2757 3125
rect 2791 3091 2802 3125
rect 2749 3057 2802 3091
rect 2749 3023 2757 3057
rect 2791 3023 2802 3057
rect 2749 2945 2802 3023
rect 2902 3533 2958 3545
rect 2902 3499 2913 3533
rect 2947 3499 2958 3533
rect 2902 3465 2958 3499
rect 2902 3431 2913 3465
rect 2947 3431 2958 3465
rect 2902 3397 2958 3431
rect 2902 3363 2913 3397
rect 2947 3363 2958 3397
rect 2902 3329 2958 3363
rect 2902 3295 2913 3329
rect 2947 3295 2958 3329
rect 2902 3261 2958 3295
rect 2902 3227 2913 3261
rect 2947 3227 2958 3261
rect 2902 3193 2958 3227
rect 2902 3159 2913 3193
rect 2947 3159 2958 3193
rect 2902 3125 2958 3159
rect 2902 3091 2913 3125
rect 2947 3091 2958 3125
rect 2902 3057 2958 3091
rect 2902 3023 2913 3057
rect 2947 3023 2958 3057
rect 2902 2945 2958 3023
rect 3032 3533 3085 3545
rect 3032 3499 3040 3533
rect 3074 3499 3085 3533
rect 3032 3465 3085 3499
rect 3032 3431 3040 3465
rect 3074 3431 3085 3465
rect 3032 3397 3085 3431
rect 3032 3363 3040 3397
rect 3074 3363 3085 3397
rect 3032 3329 3085 3363
rect 3032 3295 3040 3329
rect 3074 3295 3085 3329
rect 3032 3261 3085 3295
rect 3032 3227 3040 3261
rect 3074 3227 3085 3261
rect 3032 3193 3085 3227
rect 3032 3159 3040 3193
rect 3074 3159 3085 3193
rect 3032 3125 3085 3159
rect 3032 3091 3040 3125
rect 3074 3091 3085 3125
rect 3032 3057 3085 3091
rect 3032 3023 3040 3057
rect 3074 3023 3085 3057
rect 3032 2945 3085 3023
rect 3185 3533 3241 3545
rect 3185 3499 3196 3533
rect 3230 3499 3241 3533
rect 3185 3465 3241 3499
rect 3185 3431 3196 3465
rect 3230 3431 3241 3465
rect 3185 3397 3241 3431
rect 3185 3363 3196 3397
rect 3230 3363 3241 3397
rect 3185 3329 3241 3363
rect 3185 3295 3196 3329
rect 3230 3295 3241 3329
rect 3185 3261 3241 3295
rect 3185 3227 3196 3261
rect 3230 3227 3241 3261
rect 3185 3193 3241 3227
rect 3185 3159 3196 3193
rect 3230 3159 3241 3193
rect 3185 3125 3241 3159
rect 3185 3091 3196 3125
rect 3230 3091 3241 3125
rect 3185 3057 3241 3091
rect 3185 3023 3196 3057
rect 3230 3023 3241 3057
rect 3185 2945 3241 3023
rect 3341 3533 3397 3545
rect 3341 3499 3352 3533
rect 3386 3499 3397 3533
rect 3341 3465 3397 3499
rect 3341 3431 3352 3465
rect 3386 3431 3397 3465
rect 3341 3397 3397 3431
rect 3341 3363 3352 3397
rect 3386 3363 3397 3397
rect 3341 3329 3397 3363
rect 3341 3295 3352 3329
rect 3386 3295 3397 3329
rect 3341 3261 3397 3295
rect 3341 3227 3352 3261
rect 3386 3227 3397 3261
rect 3341 3193 3397 3227
rect 3341 3159 3352 3193
rect 3386 3159 3397 3193
rect 3341 3125 3397 3159
rect 3341 3091 3352 3125
rect 3386 3091 3397 3125
rect 3341 3057 3397 3091
rect 3341 3023 3352 3057
rect 3386 3023 3397 3057
rect 3341 2945 3397 3023
rect 3497 3533 3553 3545
rect 3497 3499 3508 3533
rect 3542 3499 3553 3533
rect 3497 3465 3553 3499
rect 3497 3431 3508 3465
rect 3542 3431 3553 3465
rect 3497 3397 3553 3431
rect 3497 3363 3508 3397
rect 3542 3363 3553 3397
rect 3497 3329 3553 3363
rect 3497 3295 3508 3329
rect 3542 3295 3553 3329
rect 3497 3261 3553 3295
rect 3497 3227 3508 3261
rect 3542 3227 3553 3261
rect 3497 3193 3553 3227
rect 3497 3159 3508 3193
rect 3542 3159 3553 3193
rect 3497 3125 3553 3159
rect 3497 3091 3508 3125
rect 3542 3091 3553 3125
rect 3497 3057 3553 3091
rect 3497 3023 3508 3057
rect 3542 3023 3553 3057
rect 3497 2945 3553 3023
rect 2165 2897 2176 2931
rect 2210 2897 2221 2931
rect 2165 2863 2221 2897
rect 2165 2829 2176 2863
rect 2210 2829 2221 2863
rect 2165 2795 2221 2829
rect 2165 2761 2176 2795
rect 2210 2761 2221 2795
rect 2165 2727 2221 2761
rect 2165 2693 2176 2727
rect 2210 2693 2221 2727
rect 2165 2659 2221 2693
rect 2165 2625 2176 2659
rect 2210 2625 2221 2659
rect 2165 2591 2221 2625
rect 2165 2557 2176 2591
rect 2210 2557 2221 2591
rect 2165 2545 2221 2557
rect 4233 3533 4289 3545
rect 4233 3499 4244 3533
rect 4278 3499 4289 3533
rect 4233 3465 4289 3499
rect 4233 3431 4244 3465
rect 4278 3431 4289 3465
rect 4233 3397 4289 3431
rect 4233 3363 4244 3397
rect 4278 3363 4289 3397
rect 4233 3329 4289 3363
rect 4233 3295 4244 3329
rect 4278 3295 4289 3329
rect 4233 3261 4289 3295
rect 4233 3227 4244 3261
rect 4278 3227 4289 3261
rect 4233 3193 4289 3227
rect 4233 3159 4244 3193
rect 4278 3159 4289 3193
rect 4233 3125 4289 3159
rect 4233 3091 4244 3125
rect 4278 3091 4289 3125
rect 4233 3057 4289 3091
rect 4233 3023 4244 3057
rect 4278 3023 4289 3057
rect 4233 2989 4289 3023
rect 4233 2955 4244 2989
rect 4278 2955 4289 2989
rect 4233 2921 4289 2955
rect 4233 2887 4244 2921
rect 4278 2887 4289 2921
rect 4233 2853 4289 2887
rect 4233 2819 4244 2853
rect 4278 2819 4289 2853
rect 4233 2785 4289 2819
rect 4233 2751 4244 2785
rect 4278 2751 4289 2785
rect 4233 2717 4289 2751
rect 4233 2683 4244 2717
rect 4278 2683 4289 2717
rect 4233 2649 4289 2683
rect 4233 2615 4244 2649
rect 4278 2615 4289 2649
rect 4233 2545 4289 2615
rect 4389 3533 4445 3545
rect 4389 3499 4400 3533
rect 4434 3499 4445 3533
rect 4389 3465 4445 3499
rect 4389 3431 4400 3465
rect 4434 3431 4445 3465
rect 4389 3397 4445 3431
rect 4389 3363 4400 3397
rect 4434 3363 4445 3397
rect 4389 3329 4445 3363
rect 4389 3295 4400 3329
rect 4434 3295 4445 3329
rect 4389 3261 4445 3295
rect 4389 3227 4400 3261
rect 4434 3227 4445 3261
rect 4389 3193 4445 3227
rect 4389 3159 4400 3193
rect 4434 3159 4445 3193
rect 4389 3125 4445 3159
rect 4389 3091 4400 3125
rect 4434 3091 4445 3125
rect 4389 3057 4445 3091
rect 4389 3023 4400 3057
rect 4434 3023 4445 3057
rect 4389 2989 4445 3023
rect 4389 2955 4400 2989
rect 4434 2955 4445 2989
rect 4389 2921 4445 2955
rect 4389 2887 4400 2921
rect 4434 2887 4445 2921
rect 4389 2853 4445 2887
rect 4389 2819 4400 2853
rect 4434 2819 4445 2853
rect 4389 2785 4445 2819
rect 4389 2751 4400 2785
rect 4434 2751 4445 2785
rect 4389 2717 4445 2751
rect 4389 2683 4400 2717
rect 4434 2683 4445 2717
rect 4389 2649 4445 2683
rect 4389 2615 4400 2649
rect 4434 2615 4445 2649
rect 4389 2545 4445 2615
rect 5205 3470 5261 3488
rect 5205 3436 5216 3470
rect 5250 3436 5261 3470
rect 5205 3402 5261 3436
rect 5205 3368 5216 3402
rect 5250 3368 5261 3402
rect 5205 3334 5261 3368
rect 5205 3300 5216 3334
rect 5250 3300 5261 3334
rect 5205 3288 5261 3300
rect 5421 3470 5477 3488
rect 5421 3436 5432 3470
rect 5466 3436 5477 3470
rect 5421 3402 5477 3436
rect 5421 3368 5432 3402
rect 5466 3368 5477 3402
rect 5421 3334 5477 3368
rect 5421 3300 5432 3334
rect 5466 3300 5477 3334
rect 5421 3288 5477 3300
rect 5205 2964 5261 2982
rect 5205 2930 5216 2964
rect 5250 2930 5261 2964
rect 5205 2896 5261 2930
rect 5205 2862 5216 2896
rect 5250 2862 5261 2896
rect 5205 2828 5261 2862
rect 5205 2794 5216 2828
rect 5250 2794 5261 2828
rect 5205 2782 5261 2794
rect 5421 2964 5477 2982
rect 5421 2930 5432 2964
rect 5466 2930 5477 2964
rect 5421 2896 5477 2930
rect 5421 2862 5432 2896
rect 5466 2862 5477 2896
rect 5421 2828 5477 2862
rect 5421 2794 5432 2828
rect 5466 2794 5477 2828
rect 5421 2782 5477 2794
rect 6190 3317 6390 3325
rect 6190 3283 6208 3317
rect 6242 3283 6276 3317
rect 6310 3283 6344 3317
rect 6378 3283 6390 3317
rect 6190 3272 6390 3283
rect 6458 3317 6658 3325
rect 6458 3283 6470 3317
rect 6504 3283 6538 3317
rect 6572 3283 6606 3317
rect 6640 3283 6658 3317
rect 6458 3272 6658 3283
rect 6190 3141 6390 3152
rect 6190 3107 6208 3141
rect 6242 3107 6276 3141
rect 6310 3107 6344 3141
rect 6378 3107 6390 3141
rect 6190 3096 6390 3107
rect 6458 3141 6658 3152
rect 6458 3107 6470 3141
rect 6504 3107 6538 3141
rect 6572 3107 6606 3141
rect 6640 3107 6658 3141
rect 6458 3096 6658 3107
rect 6190 2965 6390 2976
rect 6190 2931 6208 2965
rect 6242 2931 6276 2965
rect 6310 2931 6344 2965
rect 6378 2931 6390 2965
rect 6190 2923 6390 2931
rect 6458 2965 6658 2976
rect 6458 2931 6470 2965
rect 6504 2931 6538 2965
rect 6572 2931 6606 2965
rect 6640 2931 6658 2965
rect 6458 2923 6658 2931
rect 6190 2840 6390 2848
rect 6190 2806 6208 2840
rect 6242 2806 6276 2840
rect 6310 2806 6344 2840
rect 6378 2806 6390 2840
rect 6190 2795 6390 2806
rect 6458 2840 6658 2848
rect 6458 2806 6470 2840
rect 6504 2806 6538 2840
rect 6572 2806 6606 2840
rect 6640 2806 6658 2840
rect 6458 2795 6658 2806
rect 6190 2664 6390 2675
rect 6190 2630 6208 2664
rect 6242 2630 6276 2664
rect 6310 2630 6344 2664
rect 6378 2630 6390 2664
rect 6190 2622 6390 2630
rect 6458 2664 6658 2675
rect 6458 2630 6470 2664
rect 6504 2630 6538 2664
rect 6572 2630 6606 2664
rect 6640 2630 6658 2664
rect 6458 2622 6658 2630
<< mvndiffc >>
rect -31512 -8719 -31478 -8685
rect -29268 -8731 -29234 -8697
rect 244 2191 278 2225
rect 244 2123 278 2157
rect 244 2055 278 2089
rect 480 2191 514 2225
rect 480 2123 514 2157
rect 480 2055 514 2089
rect 5878 3283 5912 3317
rect 5946 3283 5980 3317
rect 5878 2931 5912 2965
rect 5946 2931 5980 2965
rect 5878 2806 5912 2840
rect 5946 2806 5980 2840
rect 5878 2630 5912 2664
rect 5946 2630 5980 2664
rect -221 1797 -187 1831
rect -221 1729 -187 1763
rect -221 1661 -187 1695
rect -221 1593 -187 1627
rect -221 1525 -187 1559
rect -221 1457 -187 1491
rect -221 1389 -187 1423
rect -221 1321 -187 1355
rect -221 1253 -187 1287
rect -221 1185 -187 1219
rect -221 1117 -187 1151
rect -221 1049 -187 1083
rect -221 981 -187 1015
rect -221 913 -187 947
rect -5 1797 29 1831
rect -5 1729 29 1763
rect -5 1661 29 1695
rect -5 1593 29 1627
rect -5 1525 29 1559
rect -5 1457 29 1491
rect -5 1389 29 1423
rect -5 1321 29 1355
rect -5 1253 29 1287
rect -5 1185 29 1219
rect -5 1117 29 1151
rect -5 1049 29 1083
rect -5 981 29 1015
rect -5 913 29 947
rect 126 1797 160 1831
rect 126 1729 160 1763
rect 126 1661 160 1695
rect 126 1593 160 1627
rect 126 1525 160 1559
rect 126 1457 160 1491
rect 126 1389 160 1423
rect 126 1321 160 1355
rect 126 1253 160 1287
rect 126 1185 160 1219
rect 126 1117 160 1151
rect 126 1049 160 1083
rect 126 981 160 1015
rect 126 913 160 947
rect 342 1797 376 1831
rect 342 1729 376 1763
rect 342 1661 376 1695
rect 342 1593 376 1627
rect 342 1525 376 1559
rect 342 1457 376 1491
rect 342 1389 376 1423
rect 342 1321 376 1355
rect 342 1253 376 1287
rect 342 1185 376 1219
rect 342 1117 376 1151
rect 342 1049 376 1083
rect 342 981 376 1015
rect 342 913 376 947
rect 558 1797 592 1831
rect 558 1729 592 1763
rect 558 1661 592 1695
rect 558 1593 592 1627
rect 558 1525 592 1559
rect 558 1457 592 1491
rect 558 1389 592 1423
rect 558 1321 592 1355
rect 558 1253 592 1287
rect 558 1185 592 1219
rect 558 1117 592 1151
rect 558 1049 592 1083
rect 558 981 592 1015
rect 558 913 592 947
rect 774 1797 808 1831
rect 774 1729 808 1763
rect 774 1661 808 1695
rect 774 1593 808 1627
rect 774 1525 808 1559
rect 774 1457 808 1491
rect 774 1389 808 1423
rect 774 1321 808 1355
rect 774 1253 808 1287
rect 774 1185 808 1219
rect 774 1117 808 1151
rect 774 1049 808 1083
rect 774 981 808 1015
rect 774 913 808 947
rect 990 1797 1024 1831
rect 990 1729 1024 1763
rect 990 1661 1024 1695
rect 990 1593 1024 1627
rect 990 1525 1024 1559
rect 990 1457 1024 1491
rect 990 1389 1024 1423
rect 990 1321 1024 1355
rect 990 1253 1024 1287
rect 990 1185 1024 1219
rect 990 1117 1024 1151
rect 990 1049 1024 1083
rect 990 981 1024 1015
rect 990 913 1024 947
rect 1206 1797 1240 1831
rect 1206 1729 1240 1763
rect 1206 1661 1240 1695
rect 1206 1593 1240 1627
rect 1206 1525 1240 1559
rect 1206 1457 1240 1491
rect 1206 1389 1240 1423
rect 1206 1321 1240 1355
rect 1206 1253 1240 1287
rect 1206 1185 1240 1219
rect 1206 1117 1240 1151
rect 1206 1049 1240 1083
rect 1206 981 1240 1015
rect 1206 913 1240 947
rect 1422 1797 1456 1831
rect 1422 1729 1456 1763
rect 1422 1661 1456 1695
rect 1422 1593 1456 1627
rect 1422 1525 1456 1559
rect 1422 1457 1456 1491
rect 1422 1389 1456 1423
rect 1422 1321 1456 1355
rect 1422 1253 1456 1287
rect 1422 1185 1456 1219
rect 1422 1117 1456 1151
rect 1422 1049 1456 1083
rect 1422 981 1456 1015
rect 1422 913 1456 947
rect 1638 1797 1672 1831
rect 1638 1729 1672 1763
rect 1638 1661 1672 1695
rect 1638 1593 1672 1627
rect 1638 1525 1672 1559
rect 1638 1457 1672 1491
rect 1638 1389 1672 1423
rect 1638 1321 1672 1355
rect 1638 1253 1672 1287
rect 1638 1185 1672 1219
rect 1638 1117 1672 1151
rect 1638 1049 1672 1083
rect 1638 981 1672 1015
rect 1638 913 1672 947
rect 1854 1797 1888 1831
rect 1854 1729 1888 1763
rect 1854 1661 1888 1695
rect 1854 1593 1888 1627
rect 1854 1525 1888 1559
rect 1854 1457 1888 1491
rect 1854 1389 1888 1423
rect 1854 1321 1888 1355
rect 1854 1253 1888 1287
rect 2131 1774 2165 1808
rect 2131 1706 2165 1740
rect 2131 1638 2165 1672
rect 2131 1570 2165 1604
rect 2131 1502 2165 1536
rect 2131 1434 2165 1468
rect 2131 1366 2165 1400
rect 2131 1298 2165 1332
rect 2287 1774 2321 1808
rect 2287 1706 2321 1740
rect 2287 1638 2321 1672
rect 2287 1570 2321 1604
rect 2287 1502 2321 1536
rect 2287 1434 2321 1468
rect 2287 1366 2321 1400
rect 2287 1298 2321 1332
rect 2414 1774 2448 1808
rect 2414 1706 2448 1740
rect 2414 1638 2448 1672
rect 2414 1570 2448 1604
rect 2414 1502 2448 1536
rect 2414 1434 2448 1468
rect 2414 1366 2448 1400
rect 2414 1298 2448 1332
rect 2570 1774 2604 1808
rect 2570 1706 2604 1740
rect 2570 1638 2604 1672
rect 2570 1570 2604 1604
rect 2570 1502 2604 1536
rect 2570 1434 2604 1468
rect 2570 1366 2604 1400
rect 2570 1298 2604 1332
rect 2697 1803 2731 1837
rect 2697 1735 2731 1769
rect 2697 1667 2731 1701
rect 2697 1599 2731 1633
rect 2697 1531 2731 1565
rect 2697 1463 2731 1497
rect 2697 1395 2731 1429
rect 2697 1327 2731 1361
rect 2697 1259 2731 1293
rect 1854 1185 1888 1219
rect 1854 1117 1888 1151
rect 1854 1049 1888 1083
rect 1854 981 1888 1015
rect 1854 913 1888 947
rect 2697 1191 2731 1225
rect 2697 1123 2731 1157
rect 2697 1055 2731 1089
rect 2697 987 2731 1021
rect 2697 919 2731 953
rect 2853 1803 2887 1837
rect 2853 1735 2887 1769
rect 2853 1667 2887 1701
rect 2853 1599 2887 1633
rect 2853 1531 2887 1565
rect 2853 1463 2887 1497
rect 2853 1395 2887 1429
rect 2853 1327 2887 1361
rect 2853 1259 2887 1293
rect 2853 1191 2887 1225
rect 2853 1123 2887 1157
rect 2853 1055 2887 1089
rect 2853 987 2887 1021
rect 2853 919 2887 953
rect 3009 1803 3043 1837
rect 3009 1735 3043 1769
rect 3009 1667 3043 1701
rect 3009 1599 3043 1633
rect 3009 1531 3043 1565
rect 3009 1463 3043 1497
rect 3009 1395 3043 1429
rect 3009 1327 3043 1361
rect 3009 1259 3043 1293
rect 3009 1191 3043 1225
rect 3009 1123 3043 1157
rect 3009 1055 3043 1089
rect 3009 987 3043 1021
rect 3009 919 3043 953
rect 3165 1803 3199 1837
rect 3165 1735 3199 1769
rect 3165 1667 3199 1701
rect 3165 1599 3199 1633
rect 3165 1531 3199 1565
rect 3165 1463 3199 1497
rect 3165 1395 3199 1429
rect 3165 1327 3199 1361
rect 3165 1259 3199 1293
rect 3165 1191 3199 1225
rect 3165 1123 3199 1157
rect 3165 1055 3199 1089
rect 3165 987 3199 1021
rect 3165 919 3199 953
rect 3321 1803 3355 1837
rect 3321 1735 3355 1769
rect 3321 1667 3355 1701
rect 3321 1599 3355 1633
rect 3321 1531 3355 1565
rect 3321 1463 3355 1497
rect 3321 1395 3355 1429
rect 3321 1327 3355 1361
rect 3446 1789 3480 1823
rect 3446 1721 3480 1755
rect 3446 1653 3480 1687
rect 3446 1585 3480 1619
rect 3446 1517 3480 1551
rect 3446 1449 3480 1483
rect 3446 1381 3480 1415
rect 3446 1313 3480 1347
rect 3602 1789 3636 1823
rect 3602 1721 3636 1755
rect 3602 1653 3636 1687
rect 3889 1807 3923 1841
rect 3889 1739 3923 1773
rect 3889 1671 3923 1705
rect 4125 1807 4159 1841
rect 4125 1739 4159 1773
rect 4125 1671 4159 1705
rect 3602 1585 3636 1619
rect 3602 1517 3636 1551
rect 3602 1449 3636 1483
rect 3602 1381 3636 1415
rect 3602 1313 3636 1347
rect 3321 1259 3355 1293
rect 3321 1191 3355 1225
rect 3321 1123 3355 1157
rect 3321 1055 3355 1089
rect 3321 987 3355 1021
rect 3321 919 3355 953
rect 193 640 227 674
rect 261 640 295 674
rect 329 640 363 674
rect 397 640 431 674
rect 465 640 499 674
rect 533 640 567 674
rect 601 640 635 674
rect 669 640 703 674
rect 737 640 771 674
rect 805 640 839 674
rect 873 640 907 674
rect 941 640 975 674
rect 1009 640 1043 674
rect 1077 640 1111 674
rect 1145 640 1179 674
rect 1213 640 1247 674
rect 1281 640 1315 674
rect 1349 640 1383 674
rect 1417 640 1451 674
rect 1485 640 1519 674
rect 1553 640 1587 674
rect 1621 640 1655 674
rect 1689 640 1723 674
rect 1757 640 1791 674
rect 1825 640 1859 674
rect 1893 640 1927 674
rect 1961 640 1995 674
rect 2029 640 2063 674
rect 2097 640 2131 674
rect 2697 633 2731 667
rect 2697 565 2731 599
rect 2697 497 2731 531
rect 2853 633 2887 667
rect 2853 565 2887 599
rect 2853 497 2887 531
rect 3009 633 3043 667
rect 3009 565 3043 599
rect 3009 497 3043 531
rect 3165 633 3199 667
rect 3165 565 3199 599
rect 3165 497 3199 531
rect 193 404 227 438
rect 261 404 295 438
rect 329 404 363 438
rect 397 404 431 438
rect 465 404 499 438
rect 533 404 567 438
rect 601 404 635 438
rect 669 404 703 438
rect 737 404 771 438
rect 805 404 839 438
rect 873 404 907 438
rect 941 404 975 438
rect 1009 404 1043 438
rect 1077 404 1111 438
rect 1145 404 1179 438
rect 1213 404 1247 438
rect 1281 404 1315 438
rect 1349 404 1383 438
rect 1417 404 1451 438
rect 1485 404 1519 438
rect 1553 404 1587 438
rect 1621 404 1655 438
rect 1689 404 1723 438
rect 1757 404 1791 438
rect 1825 404 1859 438
rect 1893 404 1927 438
rect 1961 404 1995 438
rect 2029 404 2063 438
rect 2097 404 2131 438
rect 193 277 227 311
rect 261 277 295 311
rect 329 277 363 311
rect 397 277 431 311
rect 465 277 499 311
rect 533 277 567 311
rect 601 277 635 311
rect 669 277 703 311
rect 737 277 771 311
rect 805 277 839 311
rect 873 277 907 311
rect 941 277 975 311
rect 1009 277 1043 311
rect 1077 277 1111 311
rect 1145 277 1179 311
rect 1213 277 1247 311
rect 1281 277 1315 311
rect 1349 277 1383 311
rect 1417 277 1451 311
rect 1485 277 1519 311
rect 1553 277 1587 311
rect 1621 277 1655 311
rect 1689 277 1723 311
rect 1757 277 1791 311
rect 1825 277 1859 311
rect 1893 277 1927 311
rect 1961 277 1995 311
rect 2029 277 2063 311
rect 2097 277 2131 311
rect 193 41 227 75
rect 261 41 295 75
rect 329 41 363 75
rect 397 41 431 75
rect 465 41 499 75
rect 533 41 567 75
rect 601 41 635 75
rect 669 41 703 75
rect 737 41 771 75
rect 805 41 839 75
rect 873 41 907 75
rect 941 41 975 75
rect 1009 41 1043 75
rect 1077 41 1111 75
rect 1145 41 1179 75
rect 1213 41 1247 75
rect 1281 41 1315 75
rect 1349 41 1383 75
rect 1417 41 1451 75
rect 1485 41 1519 75
rect 1553 41 1587 75
rect 1621 41 1655 75
rect 1689 41 1723 75
rect 1757 41 1791 75
rect 1825 41 1859 75
rect 1893 41 1927 75
rect 1961 41 1995 75
rect 2029 41 2063 75
rect 2097 41 2131 75
<< mvpdiffc >>
rect -746 3476 -712 3510
rect -746 3408 -712 3442
rect -746 3340 -712 3374
rect -746 3272 -712 3306
rect -746 3204 -712 3238
rect -746 3136 -712 3170
rect -746 3068 -712 3102
rect -746 3000 -712 3034
rect -746 2932 -712 2966
rect -746 2864 -712 2898
rect -746 2796 -712 2830
rect -746 2728 -712 2762
rect -746 2660 -712 2694
rect -746 2592 -712 2626
rect -590 3476 -556 3510
rect -590 3408 -556 3442
rect -590 3340 -556 3374
rect -590 3272 -556 3306
rect -590 3204 -556 3238
rect -590 3136 -556 3170
rect -590 3068 -556 3102
rect -590 3000 -556 3034
rect -590 2932 -556 2966
rect -590 2864 -556 2898
rect -590 2796 -556 2830
rect -590 2728 -556 2762
rect -590 2660 -556 2694
rect -590 2592 -556 2626
rect -434 3476 -400 3510
rect -434 3408 -400 3442
rect -434 3340 -400 3374
rect -434 3272 -400 3306
rect -434 3204 -400 3238
rect -434 3136 -400 3170
rect -434 3068 -400 3102
rect -434 3000 -400 3034
rect -434 2932 -400 2966
rect -434 2864 -400 2898
rect -434 2796 -400 2830
rect -434 2728 -400 2762
rect -434 2660 -400 2694
rect -434 2592 -400 2626
rect 168 3476 202 3510
rect 168 3408 202 3442
rect 168 3340 202 3374
rect 168 3272 202 3306
rect 168 3204 202 3238
rect 168 3136 202 3170
rect 168 3068 202 3102
rect 168 3000 202 3034
rect 168 2932 202 2966
rect 168 2864 202 2898
rect 168 2796 202 2830
rect 168 2728 202 2762
rect 168 2660 202 2694
rect 168 2592 202 2626
rect 324 3476 358 3510
rect 324 3408 358 3442
rect 324 3340 358 3374
rect 324 3272 358 3306
rect 324 3204 358 3238
rect 324 3136 358 3170
rect 324 3068 358 3102
rect 324 3000 358 3034
rect 324 2932 358 2966
rect 324 2864 358 2898
rect 324 2796 358 2830
rect 324 2728 358 2762
rect 324 2660 358 2694
rect 324 2592 358 2626
rect 480 3476 514 3510
rect 480 3408 514 3442
rect 480 3340 514 3374
rect 480 3272 514 3306
rect 480 3204 514 3238
rect 480 3136 514 3170
rect 480 3068 514 3102
rect 480 3000 514 3034
rect 480 2932 514 2966
rect 480 2864 514 2898
rect 480 2796 514 2830
rect 480 2728 514 2762
rect 480 2660 514 2694
rect 480 2592 514 2626
rect 616 3476 650 3510
rect 616 3408 650 3442
rect 616 3340 650 3374
rect 616 3272 650 3306
rect 616 3204 650 3238
rect 616 3136 650 3170
rect 616 3068 650 3102
rect 616 3000 650 3034
rect 616 2932 650 2966
rect 616 2864 650 2898
rect 616 2796 650 2830
rect 616 2728 650 2762
rect 616 2660 650 2694
rect 616 2592 650 2626
rect 772 3476 806 3510
rect 772 3408 806 3442
rect 772 3340 806 3374
rect 772 3272 806 3306
rect 772 3204 806 3238
rect 772 3136 806 3170
rect 772 3068 806 3102
rect 772 3000 806 3034
rect 772 2932 806 2966
rect 772 2864 806 2898
rect 772 2796 806 2830
rect 772 2728 806 2762
rect 772 2660 806 2694
rect 772 2592 806 2626
rect 928 3476 962 3510
rect 928 3408 962 3442
rect 928 3340 962 3374
rect 928 3272 962 3306
rect 928 3204 962 3238
rect 928 3136 962 3170
rect 928 3068 962 3102
rect 928 3000 962 3034
rect 928 2932 962 2966
rect 928 2864 962 2898
rect 928 2796 962 2830
rect 928 2728 962 2762
rect 928 2660 962 2694
rect 928 2592 962 2626
rect 1055 3476 1089 3510
rect 1055 3408 1089 3442
rect 1055 3340 1089 3374
rect 1055 3272 1089 3306
rect 1055 3204 1089 3238
rect 1055 3136 1089 3170
rect 1055 3068 1089 3102
rect 1055 3000 1089 3034
rect 1055 2932 1089 2966
rect 1055 2864 1089 2898
rect 1055 2796 1089 2830
rect 1055 2728 1089 2762
rect 1055 2660 1089 2694
rect 1055 2592 1089 2626
rect 1211 3476 1245 3510
rect 1211 3408 1245 3442
rect 1211 3340 1245 3374
rect 1211 3272 1245 3306
rect 1211 3204 1245 3238
rect 1211 3136 1245 3170
rect 1211 3068 1245 3102
rect 1211 3000 1245 3034
rect 1211 2932 1245 2966
rect 1211 2864 1245 2898
rect 1211 2796 1245 2830
rect 1211 2728 1245 2762
rect 1211 2660 1245 2694
rect 1211 2592 1245 2626
rect 1415 3476 1449 3510
rect 1415 3408 1449 3442
rect 1415 3340 1449 3374
rect 1415 3272 1449 3306
rect 1415 3204 1449 3238
rect 1415 3136 1449 3170
rect 1415 3068 1449 3102
rect 1415 3000 1449 3034
rect 1415 2932 1449 2966
rect 1415 2864 1449 2898
rect 1415 2796 1449 2830
rect 1415 2728 1449 2762
rect 1415 2660 1449 2694
rect 1415 2592 1449 2626
rect 1571 3476 1605 3510
rect 1571 3408 1605 3442
rect 1571 3340 1605 3374
rect 1571 3272 1605 3306
rect 1571 3204 1605 3238
rect 1571 3136 1605 3170
rect 1571 3068 1605 3102
rect 1571 3000 1605 3034
rect 1571 2932 1605 2966
rect 1571 2864 1605 2898
rect 1571 2796 1605 2830
rect 1571 2728 1605 2762
rect 1571 2660 1605 2694
rect 1571 2592 1605 2626
rect 1708 3441 1742 3475
rect 1708 3373 1742 3407
rect 1708 3305 1742 3339
rect 1708 3237 1742 3271
rect 1708 3169 1742 3203
rect 1708 3101 1742 3135
rect 1708 3033 1742 3067
rect 1708 2965 1742 2999
rect 1708 2897 1742 2931
rect 1708 2829 1742 2863
rect 1708 2761 1742 2795
rect 1708 2693 1742 2727
rect 1708 2625 1742 2659
rect 1708 2557 1742 2591
rect 1864 3441 1898 3475
rect 1864 3373 1898 3407
rect 1864 3305 1898 3339
rect 1864 3237 1898 3271
rect 1864 3169 1898 3203
rect 1864 3101 1898 3135
rect 1864 3033 1898 3067
rect 1864 2965 1898 2999
rect 1864 2897 1898 2931
rect 1864 2829 1898 2863
rect 1864 2761 1898 2795
rect 1864 2693 1898 2727
rect 1864 2625 1898 2659
rect 1864 2557 1898 2591
rect 2020 3441 2054 3475
rect 2020 3373 2054 3407
rect 2020 3305 2054 3339
rect 2020 3237 2054 3271
rect 2020 3169 2054 3203
rect 2020 3101 2054 3135
rect 2020 3033 2054 3067
rect 2020 2965 2054 2999
rect 2020 2897 2054 2931
rect 2020 2829 2054 2863
rect 2020 2761 2054 2795
rect 2020 2693 2054 2727
rect 2020 2625 2054 2659
rect 2020 2557 2054 2591
rect 2757 3499 2791 3533
rect 2176 3441 2210 3475
rect 2176 3373 2210 3407
rect 2311 3436 2345 3470
rect 2467 3436 2501 3470
rect 2623 3436 2657 3470
rect 2757 3431 2791 3465
rect 2176 3305 2210 3339
rect 2176 3237 2210 3271
rect 2176 3169 2210 3203
rect 2176 3101 2210 3135
rect 2757 3363 2791 3397
rect 2757 3295 2791 3329
rect 2757 3227 2791 3261
rect 2757 3159 2791 3193
rect 2176 3033 2210 3067
rect 2176 2965 2210 2999
rect 2757 3091 2791 3125
rect 2757 3023 2791 3057
rect 2913 3499 2947 3533
rect 2913 3431 2947 3465
rect 2913 3363 2947 3397
rect 2913 3295 2947 3329
rect 2913 3227 2947 3261
rect 2913 3159 2947 3193
rect 2913 3091 2947 3125
rect 2913 3023 2947 3057
rect 3040 3499 3074 3533
rect 3040 3431 3074 3465
rect 3040 3363 3074 3397
rect 3040 3295 3074 3329
rect 3040 3227 3074 3261
rect 3040 3159 3074 3193
rect 3040 3091 3074 3125
rect 3040 3023 3074 3057
rect 3196 3499 3230 3533
rect 3196 3431 3230 3465
rect 3196 3363 3230 3397
rect 3196 3295 3230 3329
rect 3196 3227 3230 3261
rect 3196 3159 3230 3193
rect 3196 3091 3230 3125
rect 3196 3023 3230 3057
rect 3352 3499 3386 3533
rect 3352 3431 3386 3465
rect 3352 3363 3386 3397
rect 3352 3295 3386 3329
rect 3352 3227 3386 3261
rect 3352 3159 3386 3193
rect 3352 3091 3386 3125
rect 3352 3023 3386 3057
rect 3508 3499 3542 3533
rect 3508 3431 3542 3465
rect 3508 3363 3542 3397
rect 3508 3295 3542 3329
rect 3508 3227 3542 3261
rect 3508 3159 3542 3193
rect 3508 3091 3542 3125
rect 3508 3023 3542 3057
rect 2176 2897 2210 2931
rect 2176 2829 2210 2863
rect 2176 2761 2210 2795
rect 2176 2693 2210 2727
rect 2176 2625 2210 2659
rect 2176 2557 2210 2591
rect 4244 3499 4278 3533
rect 4244 3431 4278 3465
rect 4244 3363 4278 3397
rect 4244 3295 4278 3329
rect 4244 3227 4278 3261
rect 4244 3159 4278 3193
rect 4244 3091 4278 3125
rect 4244 3023 4278 3057
rect 4244 2955 4278 2989
rect 4244 2887 4278 2921
rect 4244 2819 4278 2853
rect 4244 2751 4278 2785
rect 4244 2683 4278 2717
rect 4244 2615 4278 2649
rect 4400 3499 4434 3533
rect 4400 3431 4434 3465
rect 4400 3363 4434 3397
rect 4400 3295 4434 3329
rect 4400 3227 4434 3261
rect 4400 3159 4434 3193
rect 4400 3091 4434 3125
rect 4400 3023 4434 3057
rect 4400 2955 4434 2989
rect 4400 2887 4434 2921
rect 4400 2819 4434 2853
rect 4400 2751 4434 2785
rect 4400 2683 4434 2717
rect 4400 2615 4434 2649
rect 5216 3436 5250 3470
rect 5216 3368 5250 3402
rect 5216 3300 5250 3334
rect 5432 3436 5466 3470
rect 5432 3368 5466 3402
rect 5432 3300 5466 3334
rect 5216 2930 5250 2964
rect 5216 2862 5250 2896
rect 5216 2794 5250 2828
rect 5432 2930 5466 2964
rect 5432 2862 5466 2896
rect 5432 2794 5466 2828
rect 6208 3283 6242 3317
rect 6276 3283 6310 3317
rect 6344 3283 6378 3317
rect 6470 3283 6504 3317
rect 6538 3283 6572 3317
rect 6606 3283 6640 3317
rect 6208 3107 6242 3141
rect 6276 3107 6310 3141
rect 6344 3107 6378 3141
rect 6470 3107 6504 3141
rect 6538 3107 6572 3141
rect 6606 3107 6640 3141
rect 6208 2931 6242 2965
rect 6276 2931 6310 2965
rect 6344 2931 6378 2965
rect 6470 2931 6504 2965
rect 6538 2931 6572 2965
rect 6606 2931 6640 2965
rect 6208 2806 6242 2840
rect 6276 2806 6310 2840
rect 6344 2806 6378 2840
rect 6470 2806 6504 2840
rect 6538 2806 6572 2840
rect 6606 2806 6640 2840
rect 6208 2630 6242 2664
rect 6276 2630 6310 2664
rect 6344 2630 6378 2664
rect 6470 2630 6504 2664
rect 6538 2630 6572 2664
rect 6606 2630 6640 2664
<< psubdiff >>
rect 3938 3806 4106 3840
rect 4140 3806 4174 3840
rect 4208 3806 4242 3840
rect 4276 3806 4310 3840
rect 4344 3806 4378 3840
rect 4412 3806 4446 3840
rect 4480 3806 4514 3840
rect 4548 3806 4582 3840
rect 4616 3806 4650 3840
rect 4684 3806 4718 3840
rect 4752 3806 4786 3840
rect 4820 3806 4854 3840
rect 4888 3806 4922 3840
rect 4956 3806 4990 3840
rect 5024 3806 5058 3840
rect 5092 3806 5126 3840
rect 5160 3806 5194 3840
rect 5228 3806 5262 3840
rect 5296 3806 5330 3840
rect 5364 3806 5398 3840
rect 5432 3806 5466 3840
rect 5500 3806 5534 3840
rect 5568 3806 5602 3840
rect 5636 3806 5670 3840
rect 5704 3806 5772 3840
rect 3938 3734 3972 3806
rect 3938 3666 3972 3700
rect 4722 3772 4942 3806
rect 4722 3738 4723 3772
rect 4757 3738 4815 3772
rect 4849 3738 4907 3772
rect 4941 3738 4942 3772
rect 4722 3703 4942 3738
rect 4722 3669 4723 3703
rect 4757 3669 4815 3703
rect 4849 3669 4907 3703
rect 4941 3669 4942 3703
rect 3938 3598 3972 3632
rect 3938 3530 3972 3564
rect 3938 3462 3972 3496
rect 3938 3394 3972 3428
rect 3938 3326 3972 3360
rect 3938 3258 3972 3292
rect 3938 3190 3972 3224
rect 3938 3122 3972 3156
rect 3938 3054 3972 3088
rect 3938 2986 3972 3020
rect 3938 2918 3972 2952
rect 3938 2850 3972 2884
rect 3938 2782 3972 2816
rect 3938 2714 3972 2748
rect 3938 2646 3972 2680
rect 3938 2578 3972 2612
rect 3938 2510 3972 2544
rect 3938 2442 3972 2476
rect 3938 2374 3972 2408
rect 3938 2306 3972 2340
rect 3938 2238 3972 2272
rect 4722 3634 4942 3669
rect 5738 3772 5772 3806
rect 5738 3704 5772 3738
rect 4722 3600 4723 3634
rect 4757 3600 4815 3634
rect 4849 3600 4907 3634
rect 4941 3600 4942 3634
rect 4722 3565 4942 3600
rect 4722 3531 4723 3565
rect 4757 3531 4815 3565
rect 4849 3531 4907 3565
rect 4941 3531 4942 3565
rect 4722 3496 4942 3531
rect 4722 3462 4723 3496
rect 4757 3462 4815 3496
rect 4849 3462 4907 3496
rect 4941 3462 4942 3496
rect 4722 3427 4942 3462
rect 4722 3393 4723 3427
rect 4757 3393 4815 3427
rect 4849 3393 4907 3427
rect 4941 3393 4942 3427
rect 4722 3358 4942 3393
rect 4722 3324 4723 3358
rect 4757 3324 4815 3358
rect 4849 3324 4907 3358
rect 4941 3324 4942 3358
rect 4722 3289 4942 3324
rect 4722 3255 4723 3289
rect 4757 3255 4815 3289
rect 4849 3255 4907 3289
rect 4941 3255 4942 3289
rect 4722 3220 4942 3255
rect 4722 3186 4723 3220
rect 4757 3186 4815 3220
rect 4849 3186 4907 3220
rect 4941 3186 4942 3220
rect 4722 3150 4942 3186
rect 4722 3116 4723 3150
rect 4757 3116 4815 3150
rect 4849 3116 4907 3150
rect 4941 3116 4942 3150
rect 4722 3080 4942 3116
rect 4722 3046 4723 3080
rect 4757 3046 4815 3080
rect 4849 3046 4907 3080
rect 4941 3046 4942 3080
rect 4722 3010 4942 3046
rect 4722 2976 4723 3010
rect 4757 2976 4815 3010
rect 4849 2976 4907 3010
rect 4941 2976 4942 3010
rect 4722 2940 4942 2976
rect 4722 2906 4723 2940
rect 4757 2906 4815 2940
rect 4849 2906 4907 2940
rect 4941 2906 4942 2940
rect 4722 2870 4942 2906
rect 4722 2836 4723 2870
rect 4757 2836 4815 2870
rect 4849 2836 4907 2870
rect 4941 2836 4942 2870
rect 4722 2800 4942 2836
rect 4722 2766 4723 2800
rect 4757 2766 4815 2800
rect 4849 2766 4907 2800
rect 4941 2766 4942 2800
rect 4722 2730 4942 2766
rect 4722 2696 4723 2730
rect 4757 2696 4815 2730
rect 4849 2696 4907 2730
rect 4941 2696 4942 2730
rect 4722 2660 4942 2696
rect 4722 2626 4723 2660
rect 4757 2626 4815 2660
rect 4849 2626 4907 2660
rect 4941 2626 4942 2660
rect 4722 2590 4942 2626
rect 4722 2556 4723 2590
rect 4757 2556 4815 2590
rect 4849 2556 4907 2590
rect 4941 2556 4942 2590
rect 4722 2520 4942 2556
rect 4722 2486 4723 2520
rect 4757 2486 4815 2520
rect 4849 2486 4907 2520
rect 4941 2486 4942 2520
rect 4722 2450 4942 2486
rect 4722 2416 4723 2450
rect 4757 2416 4815 2450
rect 4849 2416 4907 2450
rect 4941 2416 4942 2450
rect 4722 2380 4942 2416
rect 4722 2346 4723 2380
rect 4757 2346 4815 2380
rect 4849 2346 4907 2380
rect 4941 2346 4942 2380
rect 4722 2310 4942 2346
rect 4722 2276 4723 2310
rect 4757 2276 4815 2310
rect 4849 2276 4907 2310
rect 4941 2276 4942 2310
rect 3938 2170 3972 2204
rect 3938 2102 3972 2136
rect 4722 2240 4942 2276
rect 5738 3636 5772 3670
rect 5738 3568 5772 3602
rect 5738 3500 5772 3534
rect 5738 3433 5772 3466
rect 4722 2206 4723 2240
rect 4757 2206 4815 2240
rect 4849 2206 4907 2240
rect 4941 2206 4942 2240
rect 4722 2170 4942 2206
rect 4722 2136 4723 2170
rect 4757 2136 4815 2170
rect 4849 2136 4907 2170
rect 4941 2136 4942 2170
rect 4722 2102 4942 2136
rect 5738 2102 5772 2509
rect 3938 2068 4038 2102
rect 4072 2068 4106 2102
rect 4140 2068 4174 2102
rect 4208 2068 4242 2102
rect 4276 2068 4310 2102
rect 4344 2068 4378 2102
rect 4412 2068 4446 2102
rect 4480 2068 4514 2102
rect 4548 2068 4582 2102
rect 4616 2068 4650 2102
rect 4684 2068 4718 2102
rect 4752 2068 4786 2102
rect 4820 2068 4854 2102
rect 4888 2068 4922 2102
rect 4956 2068 4990 2102
rect 5024 2068 5058 2102
rect 5092 2068 5126 2102
rect 5160 2068 5194 2102
rect 5228 2068 5262 2102
rect 5296 2068 5330 2102
rect 5364 2068 5398 2102
rect 5432 2068 5466 2102
rect 5500 2068 5534 2102
rect 5568 2068 5602 2102
rect 5636 2068 5670 2102
rect 5704 2068 5772 2102
rect 144 793 168 827
rect 202 793 237 827
rect 271 793 306 827
rect 340 793 375 827
rect 409 793 444 827
rect 478 793 513 827
rect 547 793 582 827
rect 616 793 651 827
rect 685 793 720 827
rect 754 793 789 827
rect 823 793 858 827
rect 892 793 927 827
rect 961 793 996 827
rect 1030 793 1065 827
rect 1099 793 1134 827
rect 1168 793 1203 827
rect 1237 793 1272 827
rect 1306 793 1341 827
rect 1375 793 1410 827
rect 1444 793 1479 827
rect 1513 793 1548 827
rect 1582 793 1617 827
rect 1651 793 1686 827
rect 1720 793 1755 827
rect 1789 793 1824 827
rect 1858 793 1893 827
rect 1927 793 1962 827
rect 1996 793 2031 827
rect 2065 793 2100 827
rect 2134 793 2169 827
rect 2203 793 2238 827
rect 2272 793 2307 827
rect 2341 793 2376 827
rect 2410 793 2445 827
rect 2479 793 2514 827
rect 2548 793 2583 827
rect 2617 793 2652 827
rect 2686 793 2721 827
rect 2755 793 2790 827
rect 2824 793 2859 827
rect 2893 793 2928 827
rect 2962 793 2996 827
rect 3030 793 3064 827
rect 3098 793 3132 827
rect 3166 793 3200 827
rect 3234 793 3268 827
rect 3302 793 3336 827
rect 3370 793 3394 827
<< nsubdiff >>
rect 4125 3619 4293 3653
rect 4327 3619 4361 3653
rect 4395 3619 4429 3653
rect 4463 3619 4563 3653
rect 4125 3581 4159 3619
rect 4529 3585 4563 3619
rect 4125 3513 4159 3547
rect 4125 3445 4159 3479
rect 4125 3377 4159 3411
rect 4125 3309 4159 3343
rect 4125 3241 4159 3275
rect 4125 3173 4159 3207
rect 4125 3105 4159 3139
rect 4125 3037 4159 3071
rect 4125 2969 4159 3003
rect 4125 2901 4159 2935
rect 4125 2833 4159 2867
rect 4125 2765 4159 2799
rect 4125 2697 4159 2731
rect 4125 2629 4159 2663
rect 4125 2561 4159 2595
rect 4529 3517 4563 3551
rect 4529 3449 4563 3483
rect 4529 3381 4563 3415
rect 4529 3313 4563 3347
rect 4529 3245 4563 3279
rect 4529 3177 4563 3211
rect 4529 3109 4563 3143
rect 4529 3041 4563 3075
rect 4529 2973 4563 3007
rect 4529 2905 4563 2939
rect 4529 2837 4563 2871
rect 4529 2769 4563 2803
rect 4529 2701 4563 2735
rect 4529 2633 4563 2667
rect 4529 2565 4563 2599
rect 4125 2493 4159 2527
rect 4125 2425 4159 2459
rect 4125 2357 4159 2391
rect 4529 2497 4563 2531
rect 4529 2429 4563 2463
rect 4125 2289 4159 2323
rect 4529 2361 4563 2395
rect 4529 2289 4563 2327
rect 4125 2255 4257 2289
rect 4291 2255 4325 2289
rect 4359 2255 4393 2289
rect 4427 2255 4461 2289
rect 4495 2255 4563 2289
rect 5097 3619 5197 3653
rect 5231 3619 5265 3653
rect 5299 3619 5333 3653
rect 5367 3619 5483 3653
rect 5517 3619 5585 3653
rect 5097 3585 5131 3619
rect 5097 3517 5131 3551
rect 5551 3581 5585 3619
rect 5551 3513 5585 3547
rect 5097 3449 5131 3483
rect 5097 3381 5131 3415
rect 5097 3313 5131 3347
rect 5551 3445 5585 3479
rect 5551 3377 5585 3411
rect 5551 3309 5585 3343
rect 5097 3245 5131 3279
rect 5097 3177 5131 3211
rect 5097 3109 5131 3143
rect 5551 3241 5585 3275
rect 5551 3173 5585 3207
rect 5551 3105 5585 3139
rect 5097 3041 5131 3075
rect 5551 3037 5585 3071
rect 5097 2973 5131 3007
rect 5097 2905 5131 2939
rect 5097 2837 5131 2871
rect 5097 2769 5131 2803
rect 5551 2969 5585 3003
rect 5551 2901 5585 2935
rect 5551 2833 5585 2867
rect 5097 2701 5131 2735
rect 5097 2633 5131 2667
rect 5097 2565 5131 2599
rect 5551 2765 5585 2799
rect 5551 2697 5585 2731
rect 5551 2629 5585 2663
rect 5097 2497 5131 2531
rect 5097 2429 5131 2463
rect 5097 2361 5131 2395
rect 5097 2289 5131 2327
rect 5551 2561 5585 2595
rect 5551 2493 5585 2527
rect 5551 2425 5585 2459
rect 5551 2357 5585 2391
rect 5551 2289 5585 2323
rect 5097 2255 5165 2289
rect 5199 2255 5233 2289
rect 5267 2255 5301 2289
rect 5335 2255 5369 2289
rect 5403 2255 5437 2289
rect 5471 2255 5585 2289
<< mvpsubdiff >>
rect -32352 4310 -32315 4344
rect -32281 4310 -32247 4344
rect -32213 4310 -32179 4344
rect -32145 4310 -32111 4344
rect -32077 4310 -32043 4344
rect -32009 4310 -31975 4344
rect -31941 4310 -31907 4344
rect -31873 4310 -31839 4344
rect -31805 4310 -31771 4344
rect -31737 4310 -31703 4344
rect -31669 4310 -29078 4344
rect -29044 4310 -29010 4344
rect -28976 4310 -28942 4344
rect -28908 4310 -28874 4344
rect -28840 4310 -28806 4344
rect -28772 4310 -28738 4344
rect -28704 4310 -28670 4344
rect -28636 4310 -28602 4344
rect -28568 4310 -28534 4344
rect -28500 4310 -28466 4344
rect -28432 4310 -28398 4344
rect -28364 4310 -28330 4344
rect -28296 4310 -28262 4344
rect -28228 4310 -28194 4344
rect -28160 4310 -28126 4344
rect -28092 4310 -28058 4344
rect -28024 4310 -27990 4344
rect -27956 4310 -27922 4344
rect -27888 4310 -27854 4344
rect -27820 4310 -27786 4344
rect -27752 4310 -27718 4344
rect -27684 4310 -27650 4344
rect -27616 4310 -27582 4344
rect -27548 4310 -27514 4344
rect -27480 4310 -27446 4344
rect -27412 4310 -27378 4344
rect -27344 4310 -27310 4344
rect -27276 4310 -27242 4344
rect -27208 4310 -27174 4344
rect -27140 4310 -27106 4344
rect -27072 4310 -27036 4344
rect -32352 4276 -27036 4310
rect -32352 4275 -31632 4276
rect -32352 4241 -32315 4275
rect -32281 4241 -32247 4275
rect -32213 4241 -32179 4275
rect -32145 4241 -32111 4275
rect -32077 4241 -32043 4275
rect -32009 4241 -31975 4275
rect -31941 4241 -31907 4275
rect -31873 4241 -31839 4275
rect -31805 4241 -31771 4275
rect -31737 4241 -31703 4275
rect -31669 4242 -31632 4275
rect -31598 4242 -31563 4276
rect -31529 4242 -31494 4276
rect -31460 4242 -31425 4276
rect -31391 4242 -31356 4276
rect -31322 4242 -31287 4276
rect -31253 4242 -31218 4276
rect -31184 4242 -31149 4276
rect -31115 4242 -31080 4276
rect -31046 4242 -31011 4276
rect -30977 4242 -30942 4276
rect -30908 4242 -30873 4276
rect -30839 4242 -30804 4276
rect -30770 4242 -30735 4276
rect -30701 4242 -30666 4276
rect -30632 4242 -30597 4276
rect -30563 4242 -30528 4276
rect -30494 4242 -30459 4276
rect -30425 4242 -30390 4276
rect -30356 4242 -30321 4276
rect -30287 4242 -30252 4276
rect -30218 4242 -30183 4276
rect -30149 4242 -30114 4276
rect -30080 4242 -30045 4276
rect -30011 4242 -29976 4276
rect -29942 4242 -29907 4276
rect -29873 4242 -29838 4276
rect -29804 4242 -29769 4276
rect -29735 4242 -29700 4276
rect -29666 4242 -29631 4276
rect -29597 4242 -29562 4276
rect -29528 4242 -29493 4276
rect -29459 4242 -29424 4276
rect -29390 4242 -29355 4276
rect -29321 4242 -29286 4276
rect -29252 4242 -29217 4276
rect -29183 4242 -29148 4276
rect -29114 4275 -27036 4276
rect -29114 4242 -29078 4275
rect -31669 4241 -29078 4242
rect -29044 4241 -29010 4275
rect -28976 4241 -28942 4275
rect -28908 4241 -28874 4275
rect -28840 4241 -28806 4275
rect -28772 4241 -28738 4275
rect -28704 4241 -28670 4275
rect -28636 4241 -28602 4275
rect -28568 4241 -28534 4275
rect -28500 4241 -28466 4275
rect -28432 4241 -28398 4275
rect -28364 4241 -28330 4275
rect -28296 4241 -28262 4275
rect -28228 4241 -28194 4275
rect -28160 4241 -28126 4275
rect -28092 4241 -28058 4275
rect -28024 4241 -27990 4275
rect -27956 4241 -27922 4275
rect -27888 4241 -27854 4275
rect -27820 4241 -27786 4275
rect -27752 4241 -27718 4275
rect -27684 4241 -27650 4275
rect -27616 4241 -27582 4275
rect -27548 4241 -27514 4275
rect -27480 4241 -27446 4275
rect -27412 4241 -27378 4275
rect -27344 4241 -27310 4275
rect -27276 4241 -27242 4275
rect -27208 4241 -27174 4275
rect -27140 4241 -27106 4275
rect -27072 4241 -27036 4275
rect -32352 4206 -27036 4241
rect -32352 4172 -32315 4206
rect -32281 4172 -32247 4206
rect -32213 4172 -32179 4206
rect -32145 4172 -32111 4206
rect -32077 4172 -32043 4206
rect -32009 4172 -31975 4206
rect -31941 4172 -31907 4206
rect -31873 4172 -31839 4206
rect -31805 4172 -31771 4206
rect -31737 4172 -31703 4206
rect -31669 4172 -31632 4206
rect -31598 4172 -31563 4206
rect -31529 4172 -31494 4206
rect -31460 4172 -31425 4206
rect -31391 4172 -31356 4206
rect -31322 4172 -31287 4206
rect -31253 4172 -31218 4206
rect -31184 4172 -31149 4206
rect -31115 4172 -31080 4206
rect -31046 4172 -31011 4206
rect -30977 4172 -30942 4206
rect -30908 4172 -30873 4206
rect -30839 4172 -30804 4206
rect -30770 4172 -30735 4206
rect -30701 4172 -30666 4206
rect -30632 4172 -30597 4206
rect -30563 4172 -30528 4206
rect -30494 4172 -30459 4206
rect -30425 4172 -30390 4206
rect -30356 4172 -30321 4206
rect -30287 4172 -30252 4206
rect -30218 4172 -30183 4206
rect -30149 4172 -30114 4206
rect -30080 4172 -30045 4206
rect -30011 4172 -29976 4206
rect -29942 4172 -29907 4206
rect -29873 4172 -29838 4206
rect -29804 4172 -29769 4206
rect -29735 4172 -29700 4206
rect -29666 4172 -29631 4206
rect -29597 4172 -29562 4206
rect -29528 4172 -29493 4206
rect -29459 4172 -29424 4206
rect -29390 4172 -29355 4206
rect -29321 4172 -29286 4206
rect -29252 4172 -29217 4206
rect -29183 4172 -29148 4206
rect -29114 4172 -29078 4206
rect -29044 4172 -29010 4206
rect -28976 4172 -28942 4206
rect -28908 4172 -28874 4206
rect -28840 4172 -28806 4206
rect -28772 4172 -28738 4206
rect -28704 4172 -28670 4206
rect -28636 4172 -28602 4206
rect -28568 4172 -28534 4206
rect -28500 4172 -28466 4206
rect -28432 4172 -28398 4206
rect -28364 4172 -28330 4206
rect -28296 4172 -28262 4206
rect -28228 4172 -28194 4206
rect -28160 4172 -28126 4206
rect -28092 4172 -28058 4206
rect -28024 4172 -27990 4206
rect -27956 4172 -27922 4206
rect -27888 4172 -27854 4206
rect -27820 4172 -27786 4206
rect -27752 4172 -27718 4206
rect -27684 4172 -27650 4206
rect -27616 4172 -27582 4206
rect -27548 4172 -27514 4206
rect -27480 4172 -27446 4206
rect -27412 4172 -27378 4206
rect -27344 4172 -27310 4206
rect -27276 4172 -27242 4206
rect -27208 4172 -27174 4206
rect -27140 4172 -27106 4206
rect -27072 4172 -27036 4206
rect -32352 4137 -27036 4172
rect -32352 4103 -32315 4137
rect -32281 4103 -32247 4137
rect -32213 4103 -32179 4137
rect -32145 4103 -32111 4137
rect -32077 4103 -32043 4137
rect -32009 4103 -31975 4137
rect -31941 4103 -31907 4137
rect -31873 4103 -31839 4137
rect -31805 4103 -31771 4137
rect -31737 4103 -31703 4137
rect -31669 4136 -29078 4137
rect -31669 4103 -31632 4136
rect -32352 4102 -31632 4103
rect -31598 4102 -31563 4136
rect -31529 4102 -31494 4136
rect -31460 4102 -31425 4136
rect -31391 4102 -31356 4136
rect -31322 4102 -31287 4136
rect -31253 4102 -31218 4136
rect -31184 4102 -31149 4136
rect -31115 4102 -31080 4136
rect -31046 4102 -31011 4136
rect -30977 4102 -30942 4136
rect -30908 4102 -30873 4136
rect -30839 4102 -30804 4136
rect -30770 4102 -30735 4136
rect -30701 4102 -30666 4136
rect -30632 4102 -30597 4136
rect -30563 4102 -30528 4136
rect -30494 4102 -30459 4136
rect -30425 4102 -30390 4136
rect -30356 4102 -30321 4136
rect -30287 4102 -30252 4136
rect -30218 4102 -30183 4136
rect -30149 4102 -30114 4136
rect -30080 4102 -30045 4136
rect -30011 4102 -29976 4136
rect -29942 4102 -29907 4136
rect -29873 4102 -29838 4136
rect -29804 4102 -29769 4136
rect -29735 4102 -29700 4136
rect -29666 4102 -29631 4136
rect -29597 4102 -29562 4136
rect -29528 4102 -29493 4136
rect -29459 4102 -29424 4136
rect -29390 4102 -29355 4136
rect -29321 4102 -29286 4136
rect -29252 4102 -29217 4136
rect -29183 4102 -29148 4136
rect -29114 4103 -29078 4136
rect -29044 4103 -29010 4137
rect -28976 4103 -28942 4137
rect -28908 4103 -28874 4137
rect -28840 4103 -28806 4137
rect -28772 4103 -28738 4137
rect -28704 4103 -28670 4137
rect -28636 4103 -28602 4137
rect -28568 4103 -28534 4137
rect -28500 4103 -28466 4137
rect -28432 4103 -28398 4137
rect -28364 4103 -28330 4137
rect -28296 4103 -28262 4137
rect -28228 4103 -28194 4137
rect -28160 4103 -28126 4137
rect -28092 4103 -28058 4137
rect -28024 4103 -27990 4137
rect -27956 4103 -27922 4137
rect -27888 4103 -27854 4137
rect -27820 4103 -27786 4137
rect -27752 4103 -27718 4137
rect -27684 4103 -27650 4137
rect -27616 4103 -27582 4137
rect -27548 4103 -27514 4137
rect -27480 4103 -27446 4137
rect -27412 4103 -27378 4137
rect -27344 4103 -27310 4137
rect -27276 4103 -27242 4137
rect -27208 4103 -27174 4137
rect -27140 4103 -27106 4137
rect -27072 4103 -27036 4137
rect -29114 4102 -27036 4103
rect -32352 4068 -27036 4102
rect -32352 4034 -32315 4068
rect -32281 4034 -32247 4068
rect -32213 4034 -32179 4068
rect -32145 4034 -32111 4068
rect -32077 4034 -32043 4068
rect -32009 4034 -31975 4068
rect -31941 4034 -31907 4068
rect -31873 4034 -31839 4068
rect -31805 4034 -31771 4068
rect -31737 4034 -31703 4068
rect -31669 4066 -29078 4068
rect -31669 4034 -31632 4066
rect -32352 4032 -31632 4034
rect -31598 4032 -31563 4066
rect -31529 4032 -31494 4066
rect -31460 4032 -31425 4066
rect -31391 4032 -31356 4066
rect -31322 4032 -31287 4066
rect -31253 4032 -31218 4066
rect -31184 4032 -31149 4066
rect -31115 4032 -31080 4066
rect -31046 4032 -31011 4066
rect -30977 4032 -30942 4066
rect -30908 4032 -30873 4066
rect -30839 4032 -30804 4066
rect -30770 4032 -30735 4066
rect -30701 4032 -30666 4066
rect -30632 4032 -30597 4066
rect -30563 4032 -30528 4066
rect -30494 4032 -30459 4066
rect -30425 4032 -30390 4066
rect -30356 4032 -30321 4066
rect -30287 4032 -30252 4066
rect -30218 4032 -30183 4066
rect -30149 4032 -30114 4066
rect -30080 4032 -30045 4066
rect -30011 4032 -29976 4066
rect -29942 4032 -29907 4066
rect -29873 4032 -29838 4066
rect -29804 4032 -29769 4066
rect -29735 4032 -29700 4066
rect -29666 4032 -29631 4066
rect -29597 4032 -29562 4066
rect -29528 4032 -29493 4066
rect -29459 4032 -29424 4066
rect -29390 4032 -29355 4066
rect -29321 4032 -29286 4066
rect -29252 4032 -29217 4066
rect -29183 4032 -29148 4066
rect -29114 4034 -29078 4066
rect -29044 4034 -29010 4068
rect -28976 4034 -28942 4068
rect -28908 4034 -28874 4068
rect -28840 4034 -28806 4068
rect -28772 4034 -28738 4068
rect -28704 4034 -28670 4068
rect -28636 4034 -28602 4068
rect -28568 4034 -28534 4068
rect -28500 4034 -28466 4068
rect -28432 4034 -28398 4068
rect -28364 4034 -28330 4068
rect -28296 4034 -28262 4068
rect -28228 4034 -28194 4068
rect -28160 4034 -28126 4068
rect -28092 4034 -28058 4068
rect -28024 4034 -27990 4068
rect -27956 4034 -27922 4068
rect -27888 4034 -27854 4068
rect -27820 4034 -27786 4068
rect -27752 4034 -27718 4068
rect -27684 4034 -27650 4068
rect -27616 4034 -27582 4068
rect -27548 4034 -27514 4068
rect -27480 4034 -27446 4068
rect -27412 4034 -27378 4068
rect -27344 4034 -27310 4068
rect -27276 4034 -27242 4068
rect -27208 4034 -27174 4068
rect -27140 4034 -27106 4068
rect -27072 4034 -27036 4068
rect -29114 4032 -27036 4034
rect -32352 3999 -27036 4032
rect -32352 -9635 -32315 3999
rect -31669 3996 -29078 3999
rect -31669 3962 -31632 3996
rect -31598 3962 -31563 3996
rect -31529 3962 -31494 3996
rect -31460 3962 -31425 3996
rect -31391 3962 -31356 3996
rect -31322 3962 -31287 3996
rect -31253 3962 -31218 3996
rect -31184 3962 -31149 3996
rect -31115 3962 -31080 3996
rect -31046 3962 -31011 3996
rect -30977 3962 -30942 3996
rect -30908 3962 -30873 3996
rect -30839 3962 -30804 3996
rect -30770 3962 -30735 3996
rect -30701 3962 -30666 3996
rect -30632 3962 -30597 3996
rect -30563 3962 -30528 3996
rect -30494 3962 -30459 3996
rect -30425 3962 -30390 3996
rect -30356 3962 -30321 3996
rect -30287 3962 -30252 3996
rect -30218 3962 -30183 3996
rect -30149 3962 -30114 3996
rect -30080 3962 -30045 3996
rect -30011 3962 -29976 3996
rect -29942 3962 -29907 3996
rect -29873 3962 -29838 3996
rect -29804 3962 -29769 3996
rect -29735 3962 -29700 3996
rect -29666 3962 -29631 3996
rect -29597 3962 -29562 3996
rect -29528 3962 -29493 3996
rect -29459 3962 -29424 3996
rect -29390 3962 -29355 3996
rect -29321 3962 -29286 3996
rect -29252 3962 -29217 3996
rect -29183 3962 -29148 3996
rect -29114 3965 -29078 3996
rect -29044 3965 -29010 3999
rect -28976 3965 -28942 3999
rect -28908 3965 -28874 3999
rect -28840 3965 -28806 3999
rect -28772 3965 -28738 3999
rect -28704 3965 -28670 3999
rect -28636 3965 -28602 3999
rect -28568 3965 -28534 3999
rect -28500 3965 -28466 3999
rect -28432 3965 -28398 3999
rect -28364 3965 -28330 3999
rect -28296 3965 -28262 3999
rect -28228 3965 -28194 3999
rect -28160 3965 -28126 3999
rect -28092 3965 -28058 3999
rect -28024 3965 -27990 3999
rect -27956 3965 -27922 3999
rect -27888 3965 -27854 3999
rect -27820 3965 -27786 3999
rect -27752 3965 -27718 3999
rect -27684 3965 -27650 3999
rect -27616 3965 -27582 3999
rect -27548 3965 -27514 3999
rect -27480 3965 -27446 3999
rect -27412 3965 -27378 3999
rect -27344 3965 -27310 3999
rect -27276 3965 -27242 3999
rect -27208 3965 -27174 3999
rect -27140 3965 -27106 3999
rect -27072 3965 -27036 3999
rect -29114 3962 -27036 3965
rect -31669 3930 -27036 3962
rect -31669 3926 -29078 3930
rect -31669 3892 -31632 3926
rect -31598 3892 -31563 3926
rect -31529 3892 -31494 3926
rect -31460 3892 -31425 3926
rect -31391 3892 -31356 3926
rect -31322 3892 -31287 3926
rect -31253 3892 -31218 3926
rect -31184 3892 -31149 3926
rect -31115 3892 -31080 3926
rect -31046 3892 -31011 3926
rect -30977 3892 -30942 3926
rect -30908 3892 -30873 3926
rect -30839 3892 -30804 3926
rect -30770 3892 -30735 3926
rect -30701 3892 -30666 3926
rect -30632 3892 -30597 3926
rect -30563 3892 -30528 3926
rect -30494 3892 -30459 3926
rect -30425 3892 -30390 3926
rect -30356 3892 -30321 3926
rect -30287 3892 -30252 3926
rect -30218 3892 -30183 3926
rect -30149 3892 -30114 3926
rect -30080 3892 -30045 3926
rect -30011 3892 -29976 3926
rect -29942 3892 -29907 3926
rect -29873 3892 -29838 3926
rect -29804 3892 -29769 3926
rect -29735 3892 -29700 3926
rect -29666 3892 -29631 3926
rect -29597 3892 -29562 3926
rect -29528 3892 -29493 3926
rect -29459 3892 -29424 3926
rect -29390 3892 -29355 3926
rect -29321 3892 -29286 3926
rect -29252 3892 -29217 3926
rect -29183 3892 -29148 3926
rect -29114 3896 -29078 3926
rect -29044 3896 -29010 3930
rect -28976 3896 -28942 3930
rect -28908 3896 -28874 3930
rect -28840 3896 -28806 3930
rect -28772 3896 -28738 3930
rect -28704 3896 -28670 3930
rect -28636 3896 -28602 3930
rect -28568 3896 -28534 3930
rect -28500 3896 -28466 3930
rect -28432 3896 -28398 3930
rect -28364 3896 -28330 3930
rect -28296 3896 -28262 3930
rect -28228 3896 -28194 3930
rect -28160 3896 -28126 3930
rect -28092 3896 -28058 3930
rect -28024 3896 -27990 3930
rect -27956 3896 -27922 3930
rect -27888 3896 -27854 3930
rect -27820 3896 -27786 3930
rect -27752 3896 -27718 3930
rect -27684 3896 -27650 3930
rect -27616 3896 -27582 3930
rect -27548 3896 -27514 3930
rect -27480 3896 -27446 3930
rect -27412 3896 -27378 3930
rect -27344 3896 -27310 3930
rect -27276 3896 -27242 3930
rect -27208 3896 -27174 3930
rect -27140 3896 -27106 3930
rect -27072 3896 -27036 3930
rect -29114 3892 -27036 3896
rect -31669 3861 -27036 3892
rect -31669 3856 -29078 3861
rect -31669 3822 -31632 3856
rect -31598 3822 -31563 3856
rect -31529 3822 -31494 3856
rect -31460 3822 -31425 3856
rect -31391 3822 -31356 3856
rect -31322 3822 -31287 3856
rect -31253 3822 -31218 3856
rect -31184 3822 -31149 3856
rect -31115 3822 -31080 3856
rect -31046 3822 -31011 3856
rect -30977 3822 -30942 3856
rect -30908 3822 -30873 3856
rect -30839 3822 -30804 3856
rect -30770 3822 -30735 3856
rect -30701 3822 -30666 3856
rect -30632 3822 -30597 3856
rect -30563 3822 -30528 3856
rect -30494 3822 -30459 3856
rect -30425 3822 -30390 3856
rect -30356 3822 -30321 3856
rect -30287 3822 -30252 3856
rect -30218 3822 -30183 3856
rect -30149 3822 -30114 3856
rect -30080 3822 -30045 3856
rect -30011 3822 -29976 3856
rect -29942 3822 -29907 3856
rect -29873 3822 -29838 3856
rect -29804 3822 -29769 3856
rect -29735 3822 -29700 3856
rect -29666 3822 -29631 3856
rect -29597 3822 -29562 3856
rect -29528 3822 -29493 3856
rect -29459 3822 -29424 3856
rect -29390 3822 -29355 3856
rect -29321 3822 -29286 3856
rect -29252 3822 -29217 3856
rect -29183 3822 -29148 3856
rect -29114 3827 -29078 3856
rect -29044 3827 -29010 3861
rect -28976 3827 -28942 3861
rect -28908 3827 -28874 3861
rect -28840 3827 -28806 3861
rect -28772 3827 -28738 3861
rect -28704 3827 -28670 3861
rect -28636 3827 -28602 3861
rect -28568 3827 -28534 3861
rect -28500 3827 -28466 3861
rect -28432 3827 -28398 3861
rect -28364 3827 -28330 3861
rect -28296 3827 -28262 3861
rect -28228 3827 -28194 3861
rect -28160 3827 -28126 3861
rect -28092 3827 -28058 3861
rect -28024 3827 -27990 3861
rect -27956 3827 -27922 3861
rect -27888 3827 -27854 3861
rect -27820 3827 -27786 3861
rect -27752 3827 -27718 3861
rect -27684 3827 -27650 3861
rect -27616 3827 -27582 3861
rect -27548 3827 -27514 3861
rect -27480 3827 -27446 3861
rect -27412 3827 -27378 3861
rect -27344 3827 -27310 3861
rect -27276 3827 -27242 3861
rect -27208 3827 -27174 3861
rect -27140 3827 -27106 3861
rect -27072 3827 -27036 3861
rect -29114 3822 -27036 3827
rect -31669 3792 -27036 3822
rect -31669 3786 -29078 3792
rect -31669 3752 -31632 3786
rect -31598 3752 -31563 3786
rect -31529 3752 -31494 3786
rect -31460 3752 -31425 3786
rect -31391 3752 -31356 3786
rect -31322 3752 -31287 3786
rect -31253 3752 -31218 3786
rect -31184 3752 -31149 3786
rect -31115 3752 -31080 3786
rect -31046 3752 -31011 3786
rect -30977 3752 -30942 3786
rect -30908 3752 -30873 3786
rect -30839 3752 -30804 3786
rect -30770 3752 -30735 3786
rect -30701 3752 -30666 3786
rect -30632 3752 -30597 3786
rect -30563 3752 -30528 3786
rect -30494 3752 -30459 3786
rect -30425 3752 -30390 3786
rect -30356 3752 -30321 3786
rect -30287 3752 -30252 3786
rect -30218 3752 -30183 3786
rect -30149 3752 -30114 3786
rect -30080 3752 -30045 3786
rect -30011 3752 -29976 3786
rect -29942 3752 -29907 3786
rect -29873 3752 -29838 3786
rect -29804 3752 -29769 3786
rect -29735 3752 -29700 3786
rect -29666 3752 -29631 3786
rect -29597 3752 -29562 3786
rect -29528 3752 -29493 3786
rect -29459 3752 -29424 3786
rect -29390 3752 -29355 3786
rect -29321 3752 -29286 3786
rect -29252 3752 -29217 3786
rect -29183 3752 -29148 3786
rect -29114 3758 -29078 3786
rect -29044 3758 -29010 3792
rect -28976 3758 -28942 3792
rect -28908 3758 -28874 3792
rect -28840 3758 -28806 3792
rect -28772 3758 -28738 3792
rect -28704 3758 -28670 3792
rect -28636 3758 -28602 3792
rect -28568 3758 -28534 3792
rect -28500 3758 -28466 3792
rect -28432 3758 -28398 3792
rect -28364 3758 -28330 3792
rect -28296 3758 -28262 3792
rect -28228 3758 -28194 3792
rect -28160 3758 -28126 3792
rect -28092 3758 -28058 3792
rect -28024 3758 -27990 3792
rect -27956 3758 -27922 3792
rect -27888 3758 -27854 3792
rect -27820 3758 -27786 3792
rect -27752 3758 -27718 3792
rect -27684 3758 -27650 3792
rect -27616 3758 -27582 3792
rect -27548 3758 -27514 3792
rect -27480 3758 -27446 3792
rect -27412 3758 -27378 3792
rect -27344 3758 -27310 3792
rect -27276 3758 -27242 3792
rect -27208 3758 -27174 3792
rect -27140 3758 -27106 3792
rect -27072 3758 -27036 3792
rect -29114 3752 -27036 3758
rect -31669 3723 -27036 3752
rect -31669 3716 -29078 3723
rect -31669 3682 -31632 3716
rect -31598 3682 -31563 3716
rect -31529 3682 -31494 3716
rect -31460 3682 -31425 3716
rect -31391 3682 -31356 3716
rect -31322 3682 -31287 3716
rect -31253 3682 -31218 3716
rect -31184 3682 -31149 3716
rect -31115 3682 -31080 3716
rect -31046 3682 -31011 3716
rect -30977 3682 -30942 3716
rect -30908 3682 -30873 3716
rect -30839 3682 -30804 3716
rect -30770 3682 -30735 3716
rect -30701 3682 -30666 3716
rect -30632 3682 -30597 3716
rect -30563 3682 -30528 3716
rect -30494 3682 -30459 3716
rect -30425 3682 -30390 3716
rect -30356 3682 -30321 3716
rect -30287 3682 -30252 3716
rect -30218 3682 -30183 3716
rect -30149 3682 -30114 3716
rect -30080 3682 -30045 3716
rect -30011 3682 -29976 3716
rect -29942 3682 -29907 3716
rect -29873 3682 -29838 3716
rect -29804 3682 -29769 3716
rect -29735 3682 -29700 3716
rect -29666 3682 -29631 3716
rect -29597 3682 -29562 3716
rect -29528 3682 -29493 3716
rect -29459 3682 -29424 3716
rect -29390 3682 -29355 3716
rect -29321 3682 -29286 3716
rect -29252 3682 -29217 3716
rect -29183 3682 -29148 3716
rect -29114 3689 -29078 3716
rect -29044 3689 -29010 3723
rect -28976 3689 -28942 3723
rect -28908 3689 -28874 3723
rect -28840 3689 -28806 3723
rect -28772 3689 -28738 3723
rect -28704 3689 -28670 3723
rect -28636 3689 -28602 3723
rect -28568 3689 -28534 3723
rect -28500 3689 -28466 3723
rect -28432 3689 -28398 3723
rect -28364 3689 -28330 3723
rect -28296 3689 -28262 3723
rect -28228 3689 -28194 3723
rect -28160 3689 -28126 3723
rect -28092 3689 -28058 3723
rect -28024 3689 -27990 3723
rect -27956 3689 -27922 3723
rect -27888 3689 -27854 3723
rect -27820 3689 -27786 3723
rect -27752 3689 -27718 3723
rect -27684 3689 -27650 3723
rect -27616 3689 -27582 3723
rect -27548 3689 -27514 3723
rect -27480 3689 -27446 3723
rect -27412 3689 -27378 3723
rect -27344 3689 -27310 3723
rect -27276 3689 -27242 3723
rect -27208 3689 -27174 3723
rect -27140 3689 -27106 3723
rect -27072 3689 -27036 3723
rect -29114 3682 -27036 3689
rect -31669 3654 -27036 3682
rect -31669 3646 -29078 3654
rect -31669 3612 -31632 3646
rect -31598 3612 -31563 3646
rect -31529 3612 -31494 3646
rect -31460 3612 -31425 3646
rect -31391 3612 -31356 3646
rect -31322 3612 -31287 3646
rect -31253 3612 -31218 3646
rect -31184 3612 -31149 3646
rect -31115 3612 -31080 3646
rect -31046 3612 -31011 3646
rect -30977 3612 -30942 3646
rect -30908 3612 -30873 3646
rect -30839 3612 -30804 3646
rect -30770 3612 -30735 3646
rect -30701 3612 -30666 3646
rect -30632 3612 -30597 3646
rect -30563 3612 -30528 3646
rect -30494 3612 -30459 3646
rect -30425 3612 -30390 3646
rect -30356 3612 -30321 3646
rect -30287 3612 -30252 3646
rect -30218 3612 -30183 3646
rect -30149 3612 -30114 3646
rect -30080 3612 -30045 3646
rect -30011 3612 -29976 3646
rect -29942 3612 -29907 3646
rect -29873 3612 -29838 3646
rect -29804 3612 -29769 3646
rect -29735 3612 -29700 3646
rect -29666 3612 -29631 3646
rect -29597 3612 -29562 3646
rect -29528 3612 -29493 3646
rect -29459 3612 -29424 3646
rect -29390 3612 -29355 3646
rect -29321 3612 -29286 3646
rect -29252 3612 -29217 3646
rect -29183 3612 -29148 3646
rect -29114 3620 -29078 3646
rect -29044 3620 -29010 3654
rect -28976 3620 -28942 3654
rect -28908 3620 -28874 3654
rect -28840 3620 -28806 3654
rect -28772 3620 -28738 3654
rect -28704 3620 -28670 3654
rect -28636 3620 -28602 3654
rect -28568 3620 -28534 3654
rect -28500 3620 -28466 3654
rect -28432 3620 -28398 3654
rect -28364 3620 -28330 3654
rect -28296 3620 -28262 3654
rect -28228 3620 -28194 3654
rect -28160 3620 -28126 3654
rect -28092 3620 -28058 3654
rect -28024 3620 -27990 3654
rect -27956 3620 -27922 3654
rect -27888 3620 -27854 3654
rect -27820 3620 -27786 3654
rect -27752 3620 -27718 3654
rect -27684 3620 -27650 3654
rect -27616 3620 -27582 3654
rect -27548 3620 -27514 3654
rect -27480 3620 -27446 3654
rect -27412 3620 -27378 3654
rect -27344 3620 -27310 3654
rect -27276 3620 -27242 3654
rect -27208 3620 -27174 3654
rect -27140 3620 -27106 3654
rect -27072 3620 -27036 3654
rect -29114 3612 -27036 3620
rect -31669 3585 -27036 3612
rect -31669 3576 -29078 3585
rect -31669 3542 -31632 3576
rect -31598 3542 -31563 3576
rect -31529 3542 -31494 3576
rect -31460 3542 -31425 3576
rect -31391 3542 -31356 3576
rect -31322 3542 -31287 3576
rect -31253 3542 -31218 3576
rect -31184 3542 -31149 3576
rect -31115 3542 -31080 3576
rect -31046 3542 -31011 3576
rect -30977 3542 -30942 3576
rect -30908 3542 -30873 3576
rect -30839 3542 -30804 3576
rect -30770 3542 -30735 3576
rect -30701 3542 -30666 3576
rect -30632 3542 -30597 3576
rect -30563 3542 -30528 3576
rect -30494 3542 -30459 3576
rect -30425 3542 -30390 3576
rect -30356 3542 -30321 3576
rect -30287 3542 -30252 3576
rect -30218 3542 -30183 3576
rect -30149 3542 -30114 3576
rect -30080 3542 -30045 3576
rect -30011 3542 -29976 3576
rect -29942 3542 -29907 3576
rect -29873 3542 -29838 3576
rect -29804 3542 -29769 3576
rect -29735 3542 -29700 3576
rect -29666 3542 -29631 3576
rect -29597 3542 -29562 3576
rect -29528 3542 -29493 3576
rect -29459 3542 -29424 3576
rect -29390 3542 -29355 3576
rect -29321 3542 -29286 3576
rect -29252 3542 -29217 3576
rect -29183 3542 -29148 3576
rect -29114 3551 -29078 3576
rect -29044 3551 -29010 3585
rect -28976 3551 -28942 3585
rect -28908 3551 -28874 3585
rect -28840 3551 -28806 3585
rect -28772 3551 -28738 3585
rect -28704 3551 -28670 3585
rect -28636 3551 -28602 3585
rect -28568 3551 -28534 3585
rect -28500 3551 -28466 3585
rect -28432 3551 -28398 3585
rect -28364 3551 -28330 3585
rect -28296 3551 -28262 3585
rect -28228 3551 -28194 3585
rect -28160 3551 -28126 3585
rect -28092 3551 -28058 3585
rect -28024 3551 -27990 3585
rect -27956 3551 -27922 3585
rect -27888 3551 -27854 3585
rect -27820 3551 -27786 3585
rect -27752 3551 -27718 3585
rect -27684 3551 -27650 3585
rect -27616 3551 -27582 3585
rect -27548 3551 -27514 3585
rect -27480 3551 -27446 3585
rect -27412 3551 -27378 3585
rect -27344 3551 -27310 3585
rect -27276 3551 -27242 3585
rect -27208 3551 -27174 3585
rect -27140 3551 -27106 3585
rect -27072 3551 -27036 3585
rect -29114 3542 -27036 3551
rect -31669 3516 -27036 3542
rect -31669 3506 -29078 3516
rect -31669 3472 -31632 3506
rect -31598 3472 -31563 3506
rect -31529 3472 -31494 3506
rect -31460 3472 -31425 3506
rect -31391 3472 -31356 3506
rect -31322 3472 -31287 3506
rect -31253 3472 -31218 3506
rect -31184 3472 -31149 3506
rect -31115 3472 -31080 3506
rect -31046 3472 -31011 3506
rect -30977 3472 -30942 3506
rect -30908 3472 -30873 3506
rect -30839 3472 -30804 3506
rect -30770 3472 -30735 3506
rect -30701 3472 -30666 3506
rect -30632 3472 -30597 3506
rect -30563 3472 -30528 3506
rect -30494 3472 -30459 3506
rect -30425 3472 -30390 3506
rect -30356 3472 -30321 3506
rect -30287 3472 -30252 3506
rect -30218 3472 -30183 3506
rect -30149 3472 -30114 3506
rect -30080 3472 -30045 3506
rect -30011 3472 -29976 3506
rect -29942 3472 -29907 3506
rect -29873 3472 -29838 3506
rect -29804 3472 -29769 3506
rect -29735 3472 -29700 3506
rect -29666 3472 -29631 3506
rect -29597 3472 -29562 3506
rect -29528 3472 -29493 3506
rect -29459 3472 -29424 3506
rect -29390 3472 -29355 3506
rect -29321 3472 -29286 3506
rect -29252 3472 -29217 3506
rect -29183 3472 -29148 3506
rect -29114 3482 -29078 3506
rect -29044 3482 -29010 3516
rect -28976 3482 -28942 3516
rect -28908 3482 -28874 3516
rect -28840 3482 -28806 3516
rect -28772 3482 -28738 3516
rect -28704 3482 -28670 3516
rect -28636 3482 -28602 3516
rect -28568 3482 -28534 3516
rect -28500 3482 -28466 3516
rect -28432 3482 -28398 3516
rect -28364 3482 -28330 3516
rect -28296 3482 -28262 3516
rect -28228 3482 -28194 3516
rect -28160 3482 -28126 3516
rect -28092 3482 -28058 3516
rect -28024 3482 -27990 3516
rect -27956 3482 -27922 3516
rect -27888 3482 -27854 3516
rect -27820 3482 -27786 3516
rect -27752 3482 -27718 3516
rect -27684 3482 -27650 3516
rect -27616 3482 -27582 3516
rect -27548 3482 -27514 3516
rect -27480 3482 -27446 3516
rect -27412 3482 -27378 3516
rect -27344 3482 -27310 3516
rect -27276 3482 -27242 3516
rect -27208 3482 -27174 3516
rect -27140 3482 -27106 3516
rect -27072 3482 -27036 3516
rect -29114 3472 -27036 3482
rect -31669 3447 -27036 3472
rect -31669 3436 -29078 3447
rect -31669 3402 -31632 3436
rect -31598 3402 -31563 3436
rect -31529 3402 -31494 3436
rect -31460 3402 -31425 3436
rect -31391 3402 -31356 3436
rect -31322 3402 -31287 3436
rect -31253 3402 -31218 3436
rect -31184 3402 -31149 3436
rect -31115 3402 -31080 3436
rect -31046 3402 -31011 3436
rect -30977 3402 -30942 3436
rect -30908 3402 -30873 3436
rect -30839 3402 -30804 3436
rect -30770 3402 -30735 3436
rect -30701 3402 -30666 3436
rect -30632 3402 -30597 3436
rect -30563 3402 -30528 3436
rect -30494 3402 -30459 3436
rect -30425 3402 -30390 3436
rect -30356 3402 -30321 3436
rect -30287 3402 -30252 3436
rect -30218 3402 -30183 3436
rect -30149 3402 -30114 3436
rect -30080 3402 -30045 3436
rect -30011 3402 -29976 3436
rect -29942 3402 -29907 3436
rect -29873 3402 -29838 3436
rect -29804 3402 -29769 3436
rect -29735 3402 -29700 3436
rect -29666 3402 -29631 3436
rect -29597 3402 -29562 3436
rect -29528 3402 -29493 3436
rect -29459 3402 -29424 3436
rect -29390 3402 -29355 3436
rect -29321 3402 -29286 3436
rect -29252 3402 -29217 3436
rect -29183 3402 -29148 3436
rect -29114 3413 -29078 3436
rect -29044 3413 -29010 3447
rect -28976 3413 -28942 3447
rect -28908 3413 -28874 3447
rect -28840 3413 -28806 3447
rect -28772 3413 -28738 3447
rect -28704 3413 -28670 3447
rect -28636 3413 -28602 3447
rect -28568 3413 -28534 3447
rect -28500 3413 -28466 3447
rect -28432 3413 -28398 3447
rect -28364 3413 -28330 3447
rect -28296 3413 -28262 3447
rect -28228 3413 -28194 3447
rect -28160 3413 -28126 3447
rect -28092 3413 -28058 3447
rect -28024 3413 -27990 3447
rect -27956 3413 -27922 3447
rect -27888 3413 -27854 3447
rect -27820 3413 -27786 3447
rect -27752 3413 -27718 3447
rect -27684 3413 -27650 3447
rect -27616 3413 -27582 3447
rect -27548 3413 -27514 3447
rect -27480 3413 -27446 3447
rect -27412 3413 -27378 3447
rect -27344 3413 -27310 3447
rect -27276 3413 -27242 3447
rect -27208 3413 -27174 3447
rect -27140 3413 -27106 3447
rect -27072 3413 -27036 3447
rect -29114 3402 -27036 3413
rect -31669 3378 -27036 3402
rect -31669 3344 -29078 3378
rect -29044 3344 -29010 3378
rect -28976 3344 -28942 3378
rect -28908 3344 -28874 3378
rect -28840 3344 -28806 3378
rect -28772 3344 -28738 3378
rect -28704 3344 -28670 3378
rect -28636 3344 -28602 3378
rect -28568 3344 -28534 3378
rect -28500 3344 -28466 3378
rect -28432 3344 -28398 3378
rect -28364 3344 -28330 3378
rect -28296 3344 -28262 3378
rect -28228 3344 -28194 3378
rect -28160 3344 -28126 3378
rect -28092 3344 -28058 3378
rect -28024 3344 -27990 3378
rect -27956 3344 -27922 3378
rect -27888 3344 -27854 3378
rect -27820 3344 -27786 3378
rect -27752 3344 -27718 3378
rect -27684 3344 -27650 3378
rect -27616 3344 -27582 3378
rect -27548 3344 -27514 3378
rect -27480 3344 -27446 3378
rect -27412 3344 -27378 3378
rect -27344 3344 -27310 3378
rect -27276 3344 -27242 3378
rect -27208 3344 -27174 3378
rect -27140 3344 -27106 3378
rect -27072 3344 -27036 3378
rect -31669 3334 -27036 3344
rect -31669 3300 -31564 3334
rect -31530 3300 -31496 3334
rect -31462 3300 -31428 3334
rect -31394 3300 -31360 3334
rect -31326 3300 -31292 3334
rect -31258 3300 -31224 3334
rect -31190 3300 -31156 3334
rect -31122 3300 -31088 3334
rect -31054 3300 -31020 3334
rect -30986 3300 -30952 3334
rect -30918 3300 -30884 3334
rect -30850 3300 -30816 3334
rect -30782 3300 -30748 3334
rect -30714 3300 -30680 3334
rect -30646 3300 -30612 3334
rect -30578 3300 -30544 3334
rect -30510 3300 -30476 3334
rect -30442 3300 -30408 3334
rect -30374 3300 -30340 3334
rect -30306 3300 -30272 3334
rect -30238 3300 -30204 3334
rect -30170 3300 -30136 3334
rect -30102 3300 -30068 3334
rect -30034 3300 -30000 3334
rect -29966 3300 -29932 3334
rect -29898 3300 -29864 3334
rect -29830 3300 -29796 3334
rect -29762 3300 -29728 3334
rect -29694 3300 -29660 3334
rect -29626 3300 -29592 3334
rect -29558 3300 -29524 3334
rect -29490 3300 -29456 3334
rect -29422 3300 -29388 3334
rect -29354 3300 -29260 3334
rect -29226 3309 -27036 3334
rect -29226 3300 -29078 3309
rect -31669 3223 -31598 3300
rect -31669 3189 -31632 3223
rect -29148 3275 -29078 3300
rect -29044 3275 -29010 3309
rect -28976 3275 -28942 3309
rect -28908 3275 -28874 3309
rect -28840 3275 -28806 3309
rect -28772 3275 -28738 3309
rect -28704 3275 -28670 3309
rect -28636 3275 -28602 3309
rect -28568 3275 -28534 3309
rect -28500 3275 -28466 3309
rect -28432 3275 -28398 3309
rect -28364 3275 -28330 3309
rect -28296 3275 -28262 3309
rect -28228 3275 -28194 3309
rect -28160 3275 -28126 3309
rect -28092 3275 -28058 3309
rect -28024 3275 -27990 3309
rect -27956 3275 -27922 3309
rect -27888 3275 -27854 3309
rect -27820 3275 -27786 3309
rect -27752 3275 -27718 3309
rect -27684 3275 -27650 3309
rect -27616 3275 -27582 3309
rect -27548 3275 -27514 3309
rect -27480 3275 -27446 3309
rect -27412 3275 -27378 3309
rect -27344 3275 -27310 3309
rect -27276 3275 -27242 3309
rect -27208 3275 -27174 3309
rect -27140 3275 -27106 3309
rect -27072 3275 -27036 3309
rect -29148 3266 -27036 3275
rect -29114 3240 -27036 3266
rect -29114 3232 -29078 3240
rect -31669 3155 -31598 3189
rect -31669 3121 -31632 3155
rect -31669 3087 -31598 3121
rect -31669 3053 -31632 3087
rect -31669 3019 -31598 3053
rect -31669 2985 -31632 3019
rect -31669 2951 -31598 2985
rect -31669 2917 -31632 2951
rect -31669 2883 -31598 2917
rect -31669 2849 -31632 2883
rect -31669 2815 -31598 2849
rect -31669 2781 -31632 2815
rect -31669 2747 -31598 2781
rect -31669 2713 -31632 2747
rect -31669 2679 -31598 2713
rect -31669 2645 -31632 2679
rect -31669 2611 -31598 2645
rect -31669 2577 -31632 2611
rect -31669 2543 -31598 2577
rect -31669 2509 -31632 2543
rect -31669 2475 -31598 2509
rect -31669 2441 -31632 2475
rect -31669 2407 -31598 2441
rect -31669 2373 -31632 2407
rect -31669 2339 -31598 2373
rect -31669 2305 -31632 2339
rect -31669 2271 -31598 2305
rect -31669 2237 -31632 2271
rect -31669 2203 -31598 2237
rect -31669 2169 -31632 2203
rect -31669 2135 -31598 2169
rect -31669 2101 -31632 2135
rect -31669 2067 -31598 2101
rect -31669 2033 -31632 2067
rect -31669 1999 -31598 2033
rect -31669 1965 -31632 1999
rect -31669 1931 -31598 1965
rect -31669 1897 -31632 1931
rect -31669 1863 -31598 1897
rect -31669 1829 -31632 1863
rect -31669 1795 -31598 1829
rect -31669 1761 -31632 1795
rect -31669 1727 -31598 1761
rect -31669 1693 -31632 1727
rect -31669 1659 -31598 1693
rect -31669 1625 -31632 1659
rect -31669 1591 -31598 1625
rect -31669 1557 -31632 1591
rect -31669 1523 -31598 1557
rect -31669 1489 -31632 1523
rect -31669 1455 -31598 1489
rect -31669 1421 -31632 1455
rect -31669 1387 -31598 1421
rect -31669 1353 -31632 1387
rect -31669 1319 -31598 1353
rect -31669 1285 -31632 1319
rect -31669 1251 -31598 1285
rect -31669 1217 -31632 1251
rect -31669 1183 -31598 1217
rect -31669 1149 -31632 1183
rect -31669 1115 -31598 1149
rect -31669 1081 -31632 1115
rect -31669 1047 -31598 1081
rect -31669 1013 -31632 1047
rect -31669 979 -31598 1013
rect -31669 945 -31632 979
rect -31669 911 -31598 945
rect -31669 877 -31632 911
rect -31669 843 -31598 877
rect -31669 809 -31632 843
rect -31669 775 -31598 809
rect -31669 741 -31632 775
rect -31669 707 -31598 741
rect -31669 673 -31632 707
rect -31669 639 -31598 673
rect -31669 605 -31632 639
rect -31669 571 -31598 605
rect -31669 537 -31632 571
rect -31669 503 -31598 537
rect -31669 469 -31632 503
rect -31669 435 -31598 469
rect -31669 401 -31632 435
rect -31669 367 -31598 401
rect -31669 333 -31632 367
rect -31669 299 -31598 333
rect -31669 265 -31632 299
rect -31669 231 -31598 265
rect -31669 197 -31632 231
rect -31669 163 -31598 197
rect -31669 129 -31632 163
rect -31669 95 -31598 129
rect -31669 61 -31632 95
rect -31669 27 -31598 61
rect -31669 -7 -31632 27
rect -31669 -41 -31598 -7
rect -31669 -75 -31632 -41
rect -31669 -109 -31598 -75
rect -31669 -143 -31632 -109
rect -31669 -177 -31598 -143
rect -31669 -211 -31632 -177
rect -31669 -245 -31598 -211
rect -31669 -279 -31632 -245
rect -31669 -313 -31598 -279
rect -31669 -347 -31632 -313
rect -31669 -381 -31598 -347
rect -31669 -415 -31632 -381
rect -31669 -449 -31598 -415
rect -31669 -483 -31632 -449
rect -31669 -517 -31598 -483
rect -31669 -551 -31632 -517
rect -31669 -585 -31598 -551
rect -31669 -619 -31632 -585
rect -31669 -653 -31598 -619
rect -31669 -687 -31632 -653
rect -31669 -721 -31598 -687
rect -31669 -755 -31632 -721
rect -31669 -789 -31598 -755
rect -31669 -823 -31632 -789
rect -31669 -857 -31598 -823
rect -31669 -891 -31632 -857
rect -31669 -925 -31598 -891
rect -31669 -959 -31632 -925
rect -31669 -993 -31598 -959
rect -31669 -1027 -31632 -993
rect -31669 -1061 -31598 -1027
rect -31669 -1095 -31632 -1061
rect -31669 -1129 -31598 -1095
rect -31669 -1163 -31632 -1129
rect -31669 -1197 -31598 -1163
rect -31669 -1231 -31632 -1197
rect -31669 -1265 -31598 -1231
rect -31669 -1299 -31632 -1265
rect -31669 -1333 -31598 -1299
rect -31669 -1367 -31632 -1333
rect -31669 -1401 -31598 -1367
rect -31669 -1435 -31632 -1401
rect -31669 -1469 -31598 -1435
rect -31669 -1503 -31632 -1469
rect -31669 -1537 -31598 -1503
rect -31669 -1571 -31632 -1537
rect -31669 -1605 -31598 -1571
rect -31669 -1639 -31632 -1605
rect -31669 -1673 -31598 -1639
rect -31669 -1707 -31632 -1673
rect -31669 -1741 -31598 -1707
rect -31669 -1775 -31632 -1741
rect -31669 -1809 -31598 -1775
rect -31669 -1843 -31632 -1809
rect -31669 -1877 -31598 -1843
rect -31669 -1911 -31632 -1877
rect -31669 -1945 -31598 -1911
rect -31669 -1979 -31632 -1945
rect -31669 -2013 -31598 -1979
rect -31669 -2047 -31632 -2013
rect -31669 -2081 -31598 -2047
rect -31669 -2115 -31632 -2081
rect -31669 -2149 -31598 -2115
rect -31669 -2183 -31632 -2149
rect -31669 -2217 -31598 -2183
rect -31669 -2251 -31632 -2217
rect -31669 -2285 -31598 -2251
rect -31669 -2319 -31632 -2285
rect -31669 -2353 -31598 -2319
rect -31669 -2387 -31632 -2353
rect -31669 -2421 -31598 -2387
rect -31669 -2455 -31632 -2421
rect -31669 -2489 -31598 -2455
rect -31669 -2523 -31632 -2489
rect -31669 -2557 -31598 -2523
rect -31669 -2591 -31632 -2557
rect -31669 -2625 -31598 -2591
rect -31669 -2659 -31632 -2625
rect -31669 -2693 -31598 -2659
rect -31669 -2727 -31632 -2693
rect -31669 -2761 -31598 -2727
rect -31669 -2795 -31632 -2761
rect -31669 -2829 -31598 -2795
rect -31669 -2863 -31632 -2829
rect -31669 -2897 -31598 -2863
rect -31669 -2931 -31632 -2897
rect -31669 -2965 -31598 -2931
rect -31669 -2999 -31632 -2965
rect -31669 -3033 -31598 -2999
rect -31669 -3067 -31632 -3033
rect -31669 -3101 -31598 -3067
rect -31669 -3135 -31632 -3101
rect -31669 -3169 -31598 -3135
rect -31669 -3203 -31632 -3169
rect -31669 -3237 -31598 -3203
rect -31669 -3271 -31632 -3237
rect -31669 -3305 -31598 -3271
rect -31669 -3339 -31632 -3305
rect -31669 -3373 -31598 -3339
rect -31669 -3407 -31632 -3373
rect -31669 -3441 -31598 -3407
rect -31669 -3475 -31632 -3441
rect -31669 -3509 -31598 -3475
rect -31669 -3543 -31632 -3509
rect -31669 -3577 -31598 -3543
rect -31669 -3611 -31632 -3577
rect -31669 -3645 -31598 -3611
rect -31669 -3679 -31632 -3645
rect -31669 -3713 -31598 -3679
rect -31669 -3747 -31632 -3713
rect -31669 -3781 -31598 -3747
rect -31669 -3815 -31632 -3781
rect -31669 -3849 -31598 -3815
rect -31669 -3883 -31632 -3849
rect -31669 -3917 -31598 -3883
rect -31669 -3951 -31632 -3917
rect -31669 -3985 -31598 -3951
rect -31669 -4019 -31632 -3985
rect -31669 -4053 -31598 -4019
rect -31669 -4087 -31632 -4053
rect -31669 -4121 -31598 -4087
rect -31669 -4155 -31632 -4121
rect -31669 -4189 -31598 -4155
rect -31669 -4223 -31632 -4189
rect -31669 -4257 -31598 -4223
rect -31669 -4291 -31632 -4257
rect -31669 -4325 -31598 -4291
rect -31669 -4359 -31632 -4325
rect -31669 -4393 -31598 -4359
rect -31669 -4427 -31632 -4393
rect -31669 -4461 -31598 -4427
rect -31669 -4495 -31632 -4461
rect -31669 -4529 -31598 -4495
rect -31669 -4563 -31632 -4529
rect -31669 -4597 -31598 -4563
rect -31669 -4631 -31632 -4597
rect -31669 -4665 -31598 -4631
rect -31669 -4699 -31632 -4665
rect -31669 -4733 -31598 -4699
rect -31669 -4767 -31632 -4733
rect -31669 -4801 -31598 -4767
rect -31669 -4835 -31632 -4801
rect -31669 -4869 -31598 -4835
rect -31669 -4903 -31632 -4869
rect -31669 -4937 -31598 -4903
rect -31669 -4971 -31632 -4937
rect -31669 -5005 -31598 -4971
rect -31669 -5039 -31632 -5005
rect -31669 -5073 -31598 -5039
rect -31669 -5107 -31632 -5073
rect -31669 -5141 -31598 -5107
rect -31669 -5175 -31632 -5141
rect -31669 -5209 -31598 -5175
rect -31669 -5243 -31632 -5209
rect -31669 -5277 -31598 -5243
rect -31669 -5311 -31632 -5277
rect -31669 -5345 -31598 -5311
rect -31669 -5379 -31632 -5345
rect -31669 -5413 -31598 -5379
rect -31669 -5447 -31632 -5413
rect -31669 -5481 -31598 -5447
rect -31669 -5515 -31632 -5481
rect -31669 -5549 -31598 -5515
rect -31669 -5583 -31632 -5549
rect -31669 -5617 -31598 -5583
rect -31669 -5651 -31632 -5617
rect -31669 -5685 -31598 -5651
rect -31669 -5719 -31632 -5685
rect -31669 -5753 -31598 -5719
rect -31669 -5787 -31632 -5753
rect -31669 -5821 -31598 -5787
rect -31669 -5855 -31632 -5821
rect -31669 -5889 -31598 -5855
rect -31669 -5923 -31632 -5889
rect -31669 -5957 -31598 -5923
rect -31669 -5991 -31632 -5957
rect -31669 -6025 -31598 -5991
rect -31669 -6059 -31632 -6025
rect -31669 -6093 -31598 -6059
rect -31669 -6127 -31632 -6093
rect -31669 -6161 -31598 -6127
rect -31669 -6195 -31632 -6161
rect -31669 -6229 -31598 -6195
rect -31669 -6263 -31632 -6229
rect -31669 -6297 -31598 -6263
rect -31669 -6331 -31632 -6297
rect -31669 -6365 -31598 -6331
rect -31669 -6399 -31632 -6365
rect -31669 -6433 -31598 -6399
rect -31669 -6467 -31632 -6433
rect -31669 -6501 -31598 -6467
rect -31669 -6535 -31632 -6501
rect -31669 -6569 -31598 -6535
rect -31669 -6603 -31632 -6569
rect -31669 -6637 -31598 -6603
rect -31669 -6671 -31632 -6637
rect -31669 -6705 -31598 -6671
rect -31669 -6739 -31632 -6705
rect -31669 -6773 -31598 -6739
rect -31669 -6807 -31632 -6773
rect -31669 -6841 -31598 -6807
rect -31669 -6875 -31632 -6841
rect -31669 -6909 -31598 -6875
rect -31669 -6943 -31632 -6909
rect -31669 -6977 -31598 -6943
rect -31669 -7011 -31632 -6977
rect -31669 -7045 -31598 -7011
rect -31669 -7079 -31632 -7045
rect -31669 -7113 -31598 -7079
rect -31669 -7147 -31632 -7113
rect -31669 -7181 -31598 -7147
rect -31669 -7215 -31632 -7181
rect -31669 -7249 -31598 -7215
rect -31669 -7283 -31632 -7249
rect -31669 -7317 -31598 -7283
rect -31669 -7351 -31632 -7317
rect -31669 -7385 -31598 -7351
rect -31669 -7419 -31632 -7385
rect -31669 -7453 -31598 -7419
rect -31669 -7487 -31632 -7453
rect -31669 -7521 -31598 -7487
rect -31669 -7555 -31632 -7521
rect -31669 -7589 -31598 -7555
rect -31669 -7623 -31632 -7589
rect -31669 -7657 -31598 -7623
rect -31669 -7691 -31632 -7657
rect -31669 -7725 -31598 -7691
rect -31669 -7759 -31632 -7725
rect -31669 -7793 -31598 -7759
rect -31669 -7827 -31632 -7793
rect -31669 -7861 -31598 -7827
rect -31669 -7895 -31632 -7861
rect -31669 -7929 -31598 -7895
rect -31669 -7963 -31632 -7929
rect -31669 -7997 -31598 -7963
rect -31669 -8031 -31632 -7997
rect -31669 -8065 -31598 -8031
rect -31669 -8099 -31632 -8065
rect -31669 -8133 -31598 -8099
rect -31669 -8167 -31632 -8133
rect -31669 -8201 -31598 -8167
rect -31669 -8235 -31632 -8201
rect -31669 -8269 -31598 -8235
rect -31669 -8303 -31632 -8269
rect -31669 -8337 -31598 -8303
rect -31669 -8371 -31632 -8337
rect -31669 -8405 -31598 -8371
rect -31669 -8439 -31632 -8405
rect -31669 -8473 -31598 -8439
rect -31669 -8507 -31632 -8473
rect -31669 -8541 -31598 -8507
rect -31669 -8575 -31632 -8541
rect -31669 -8609 -31598 -8575
rect -31669 -8643 -31632 -8609
rect -31669 -8677 -31598 -8643
rect -31669 -8711 -31632 -8677
rect -31669 -8745 -31598 -8711
rect -29148 3206 -29078 3232
rect -29044 3206 -29010 3240
rect -28976 3206 -28942 3240
rect -28908 3206 -28874 3240
rect -28840 3206 -28806 3240
rect -28772 3206 -28738 3240
rect -28704 3206 -28670 3240
rect -28636 3206 -28602 3240
rect -28568 3206 -28534 3240
rect -28500 3206 -28466 3240
rect -28432 3206 -28398 3240
rect -28364 3206 -28330 3240
rect -28296 3206 -28262 3240
rect -28228 3206 -28194 3240
rect -28160 3206 -28126 3240
rect -28092 3206 -28058 3240
rect -28024 3206 -27990 3240
rect -27956 3206 -27922 3240
rect -27888 3206 -27854 3240
rect -27820 3206 -27786 3240
rect -27752 3206 -27718 3240
rect -27684 3206 -27650 3240
rect -27616 3206 -27582 3240
rect -27548 3206 -27514 3240
rect -27480 3206 -27446 3240
rect -27412 3206 -27378 3240
rect -27344 3206 -27310 3240
rect -27276 3206 -27242 3240
rect -27208 3206 -27174 3240
rect -27140 3206 -27106 3240
rect -27072 3206 -27036 3240
rect -29148 3198 -27036 3206
rect -29114 3171 -27036 3198
rect -29114 3164 -29078 3171
rect -29148 3137 -29078 3164
rect -29044 3137 -29010 3171
rect -28976 3137 -28942 3171
rect -28908 3137 -28874 3171
rect -28840 3137 -28806 3171
rect -28772 3137 -28738 3171
rect -28704 3137 -28670 3171
rect -28636 3137 -28602 3171
rect -28568 3137 -28534 3171
rect -28500 3137 -28466 3171
rect -28432 3137 -28398 3171
rect -28364 3137 -28330 3171
rect -28296 3137 -28262 3171
rect -28228 3137 -28194 3171
rect -28160 3137 -28126 3171
rect -28092 3137 -28058 3171
rect -28024 3137 -27990 3171
rect -27956 3137 -27922 3171
rect -27888 3137 -27854 3171
rect -27820 3137 -27786 3171
rect -27752 3137 -27718 3171
rect -27684 3137 -27650 3171
rect -27616 3137 -27582 3171
rect -27548 3137 -27514 3171
rect -27480 3137 -27446 3171
rect -27412 3137 -27378 3171
rect -27344 3137 -27310 3171
rect -27276 3137 -27242 3171
rect -27208 3137 -27174 3171
rect -27140 3137 -27106 3171
rect -27072 3137 -27036 3171
rect -29148 3130 -27036 3137
rect -29114 3102 -27036 3130
rect -29114 3096 -29078 3102
rect -29148 3068 -29078 3096
rect -29044 3068 -29010 3102
rect -28976 3068 -28942 3102
rect -28908 3068 -28874 3102
rect -28840 3068 -28806 3102
rect -28772 3068 -28738 3102
rect -28704 3068 -28670 3102
rect -28636 3068 -28602 3102
rect -28568 3068 -28534 3102
rect -28500 3068 -28466 3102
rect -28432 3068 -28398 3102
rect -28364 3068 -28330 3102
rect -28296 3068 -28262 3102
rect -28228 3068 -28194 3102
rect -28160 3068 -28126 3102
rect -28092 3068 -28058 3102
rect -28024 3068 -27990 3102
rect -27956 3068 -27922 3102
rect -27888 3068 -27854 3102
rect -27820 3068 -27786 3102
rect -27752 3068 -27718 3102
rect -27684 3068 -27650 3102
rect -27616 3068 -27582 3102
rect -27548 3068 -27514 3102
rect -27480 3068 -27446 3102
rect -27412 3068 -27378 3102
rect -27344 3068 -27310 3102
rect -27276 3068 -27242 3102
rect -27208 3068 -27174 3102
rect -27140 3068 -27106 3102
rect -27072 3068 -27036 3102
rect -29148 3062 -27036 3068
rect -29114 3033 -27036 3062
rect -29114 3028 -29078 3033
rect -29148 2999 -29078 3028
rect -29044 2999 -29010 3033
rect -28976 2999 -28942 3033
rect -28908 2999 -28874 3033
rect -28840 2999 -28806 3033
rect -28772 2999 -28738 3033
rect -28704 2999 -28670 3033
rect -28636 2999 -28602 3033
rect -28568 2999 -28534 3033
rect -28500 2999 -28466 3033
rect -28432 2999 -28398 3033
rect -28364 2999 -28330 3033
rect -28296 2999 -28262 3033
rect -28228 2999 -28194 3033
rect -28160 2999 -28126 3033
rect -28092 2999 -28058 3033
rect -28024 2999 -27990 3033
rect -27956 2999 -27922 3033
rect -27888 2999 -27854 3033
rect -27820 2999 -27786 3033
rect -27752 2999 -27718 3033
rect -27684 2999 -27650 3033
rect -27616 2999 -27582 3033
rect -27548 2999 -27514 3033
rect -27480 2999 -27446 3033
rect -27412 2999 -27378 3033
rect -27344 2999 -27310 3033
rect -27276 2999 -27242 3033
rect -27208 2999 -27174 3033
rect -27140 2999 -27106 3033
rect -27072 2999 -27036 3033
rect -29148 2994 -27036 2999
rect -29114 2964 -27036 2994
rect -29114 2960 -29078 2964
rect -29148 2930 -29078 2960
rect -29044 2930 -29010 2964
rect -28976 2930 -28942 2964
rect -28908 2930 -28874 2964
rect -28840 2930 -28806 2964
rect -28772 2930 -28738 2964
rect -28704 2930 -28670 2964
rect -28636 2930 -28602 2964
rect -28568 2930 -28534 2964
rect -28500 2930 -28466 2964
rect -28432 2930 -28398 2964
rect -28364 2930 -28330 2964
rect -28296 2930 -28262 2964
rect -28228 2930 -28194 2964
rect -28160 2930 -28126 2964
rect -28092 2930 -28058 2964
rect -28024 2930 -27990 2964
rect -27956 2930 -27922 2964
rect -27888 2930 -27854 2964
rect -27820 2930 -27786 2964
rect -27752 2930 -27718 2964
rect -27684 2930 -27650 2964
rect -27616 2930 -27582 2964
rect -27548 2930 -27514 2964
rect -27480 2930 -27446 2964
rect -27412 2930 -27378 2964
rect -27344 2930 -27310 2964
rect -27276 2930 -27242 2964
rect -27208 2930 -27174 2964
rect -27140 2930 -27106 2964
rect -27072 2930 -27036 2964
rect -29148 2926 -27036 2930
rect -29114 2895 -27036 2926
rect -29114 2892 -29078 2895
rect -29148 2861 -29078 2892
rect -29044 2861 -29010 2895
rect -28976 2861 -28942 2895
rect -28908 2861 -28874 2895
rect -28840 2861 -28806 2895
rect -28772 2861 -28738 2895
rect -28704 2861 -28670 2895
rect -28636 2861 -28602 2895
rect -28568 2861 -28534 2895
rect -28500 2861 -28466 2895
rect -28432 2861 -28398 2895
rect -28364 2861 -28330 2895
rect -28296 2861 -28262 2895
rect -28228 2861 -28194 2895
rect -28160 2861 -28126 2895
rect -28092 2861 -28058 2895
rect -28024 2861 -27990 2895
rect -27956 2861 -27922 2895
rect -27888 2861 -27854 2895
rect -27820 2861 -27786 2895
rect -27752 2861 -27718 2895
rect -27684 2861 -27650 2895
rect -27616 2861 -27582 2895
rect -27548 2861 -27514 2895
rect -27480 2861 -27446 2895
rect -27412 2861 -27378 2895
rect -27344 2861 -27310 2895
rect -27276 2861 -27242 2895
rect -27208 2861 -27174 2895
rect -27140 2861 -27106 2895
rect -27072 2861 -27036 2895
rect -29148 2858 -27036 2861
rect -29114 2826 -27036 2858
rect -29114 2824 -29078 2826
rect -29148 2792 -29078 2824
rect -29044 2792 -29010 2826
rect -28976 2792 -28942 2826
rect -28908 2792 -28874 2826
rect -28840 2792 -28806 2826
rect -28772 2792 -28738 2826
rect -28704 2792 -28670 2826
rect -28636 2792 -28602 2826
rect -28568 2792 -28534 2826
rect -28500 2792 -28466 2826
rect -28432 2792 -28398 2826
rect -28364 2792 -28330 2826
rect -28296 2792 -28262 2826
rect -28228 2792 -28194 2826
rect -28160 2792 -28126 2826
rect -28092 2792 -28058 2826
rect -28024 2792 -27990 2826
rect -27956 2792 -27922 2826
rect -27888 2792 -27854 2826
rect -27820 2792 -27786 2826
rect -27752 2792 -27718 2826
rect -27684 2792 -27650 2826
rect -27616 2792 -27582 2826
rect -27548 2792 -27514 2826
rect -27480 2792 -27446 2826
rect -27412 2792 -27378 2826
rect -27344 2792 -27310 2826
rect -27276 2792 -27242 2826
rect -27208 2792 -27174 2826
rect -27140 2792 -27106 2826
rect -27072 2792 -27036 2826
rect -29148 2790 -27036 2792
rect -29114 2757 -27036 2790
rect -29114 2756 -29078 2757
rect -29148 2723 -29078 2756
rect -29044 2723 -29010 2757
rect -28976 2723 -28942 2757
rect -28908 2723 -28874 2757
rect -28840 2723 -28806 2757
rect -28772 2723 -28738 2757
rect -28704 2723 -28670 2757
rect -28636 2723 -28602 2757
rect -28568 2723 -28534 2757
rect -28500 2723 -28466 2757
rect -28432 2723 -28398 2757
rect -28364 2723 -28330 2757
rect -28296 2723 -28262 2757
rect -28228 2723 -28194 2757
rect -28160 2723 -28126 2757
rect -28092 2723 -28058 2757
rect -28024 2723 -27990 2757
rect -27956 2723 -27922 2757
rect -27888 2723 -27854 2757
rect -27820 2723 -27786 2757
rect -27752 2723 -27718 2757
rect -27684 2723 -27650 2757
rect -27616 2723 -27582 2757
rect -27548 2723 -27514 2757
rect -27480 2723 -27446 2757
rect -27412 2723 -27378 2757
rect -27344 2723 -27310 2757
rect -27276 2723 -27242 2757
rect -27208 2723 -27174 2757
rect -27140 2723 -27106 2757
rect -27072 2723 -27036 2757
rect -29148 2722 -27036 2723
rect -29114 2688 -27036 2722
rect -29148 2654 -29078 2688
rect -29044 2654 -29010 2688
rect -28976 2654 -28942 2688
rect -28908 2654 -28874 2688
rect -28840 2654 -28806 2688
rect -28772 2654 -28738 2688
rect -28704 2654 -28670 2688
rect -28636 2654 -28602 2688
rect -28568 2654 -28534 2688
rect -28500 2654 -28466 2688
rect -28432 2654 -28398 2688
rect -28364 2654 -28330 2688
rect -28296 2654 -28262 2688
rect -28228 2654 -28194 2688
rect -28160 2654 -28126 2688
rect -28092 2654 -28058 2688
rect -28024 2654 -27990 2688
rect -27956 2654 -27922 2688
rect -27888 2654 -27854 2688
rect -27820 2654 -27786 2688
rect -27752 2654 -27718 2688
rect -27684 2654 -27650 2688
rect -27616 2654 -27582 2688
rect -27548 2654 -27514 2688
rect -27480 2654 -27446 2688
rect -27412 2654 -27378 2688
rect -27344 2654 -27310 2688
rect -27276 2654 -27242 2688
rect -27208 2654 -27174 2688
rect -27140 2654 -27106 2688
rect -27072 2654 -27036 2688
rect -29114 2620 -27036 2654
rect -29148 2619 -27036 2620
rect -29148 2586 -29078 2619
rect -29114 2585 -29078 2586
rect -29044 2585 -29010 2619
rect -28976 2585 -28942 2619
rect -28908 2585 -28874 2619
rect -28840 2585 -28806 2619
rect -28772 2585 -28738 2619
rect -28704 2585 -28670 2619
rect -28636 2585 -28602 2619
rect -28568 2585 -28534 2619
rect -28500 2585 -28466 2619
rect -28432 2585 -28398 2619
rect -28364 2585 -28330 2619
rect -28296 2585 -28262 2619
rect -28228 2585 -28194 2619
rect -28160 2585 -28126 2619
rect -28092 2585 -28058 2619
rect -28024 2585 -27990 2619
rect -27956 2585 -27922 2619
rect -27888 2585 -27854 2619
rect -27820 2585 -27786 2619
rect -27752 2585 -27718 2619
rect -27684 2585 -27650 2619
rect -27616 2585 -27582 2619
rect -27548 2585 -27514 2619
rect -27480 2585 -27446 2619
rect -27412 2585 -27378 2619
rect -27344 2585 -27310 2619
rect -27276 2585 -27242 2619
rect -27208 2585 -27174 2619
rect -27140 2585 -27106 2619
rect -27072 2585 -27036 2619
rect -29114 2552 -27036 2585
rect -29148 2550 -27036 2552
rect -29148 2518 -29078 2550
rect -29114 2516 -29078 2518
rect -29044 2516 -29010 2550
rect -28976 2516 -28942 2550
rect -28908 2516 -28874 2550
rect -28840 2516 -28806 2550
rect -28772 2516 -28738 2550
rect -28704 2516 -28670 2550
rect -28636 2516 -28602 2550
rect -28568 2516 -28534 2550
rect -28500 2516 -28466 2550
rect -28432 2516 -28398 2550
rect -28364 2516 -28330 2550
rect -28296 2516 -28262 2550
rect -28228 2516 -28194 2550
rect -28160 2516 -28126 2550
rect -28092 2516 -28058 2550
rect -28024 2516 -27990 2550
rect -27956 2516 -27922 2550
rect -27888 2516 -27854 2550
rect -27820 2516 -27786 2550
rect -27752 2516 -27718 2550
rect -27684 2516 -27650 2550
rect -27616 2516 -27582 2550
rect -27548 2516 -27514 2550
rect -27480 2516 -27446 2550
rect -27412 2516 -27378 2550
rect -27344 2516 -27310 2550
rect -27276 2516 -27242 2550
rect -27208 2516 -27174 2550
rect -27140 2516 -27106 2550
rect -27072 2516 -27036 2550
rect -29114 2484 -27036 2516
rect -29148 2481 -27036 2484
rect -29148 2450 -29078 2481
rect -29114 2447 -29078 2450
rect -29044 2447 -29010 2481
rect -28976 2447 -28942 2481
rect -28908 2447 -28874 2481
rect -28840 2447 -28806 2481
rect -28772 2447 -28738 2481
rect -28704 2447 -28670 2481
rect -28636 2447 -28602 2481
rect -28568 2447 -28534 2481
rect -28500 2447 -28466 2481
rect -28432 2447 -28398 2481
rect -28364 2447 -28330 2481
rect -28296 2447 -28262 2481
rect -28228 2447 -28194 2481
rect -28160 2447 -28126 2481
rect -28092 2447 -28058 2481
rect -28024 2447 -27990 2481
rect -27956 2447 -27922 2481
rect -27888 2447 -27854 2481
rect -27820 2447 -27786 2481
rect -27752 2447 -27718 2481
rect -27684 2447 -27650 2481
rect -27616 2447 -27582 2481
rect -27548 2447 -27514 2481
rect -27480 2447 -27446 2481
rect -27412 2447 -27378 2481
rect -27344 2447 -27310 2481
rect -27276 2447 -27242 2481
rect -27208 2447 -27174 2481
rect -27140 2447 -27106 2481
rect -27072 2447 -27036 2481
rect -29114 2416 -27036 2447
rect -29148 2412 -27036 2416
rect -29148 2382 -29078 2412
rect -29114 2378 -29078 2382
rect -29044 2378 -29010 2412
rect -28976 2378 -28942 2412
rect -28908 2378 -28874 2412
rect -28840 2378 -28806 2412
rect -28772 2378 -28738 2412
rect -28704 2378 -28670 2412
rect -28636 2378 -28602 2412
rect -28568 2378 -28534 2412
rect -28500 2378 -28466 2412
rect -28432 2378 -28398 2412
rect -28364 2378 -28330 2412
rect -28296 2378 -28262 2412
rect -28228 2378 -28194 2412
rect -28160 2378 -28126 2412
rect -28092 2378 -28058 2412
rect -28024 2378 -27990 2412
rect -27956 2378 -27922 2412
rect -27888 2378 -27854 2412
rect -27820 2378 -27786 2412
rect -27752 2378 -27718 2412
rect -27684 2378 -27650 2412
rect -27616 2378 -27582 2412
rect -27548 2378 -27514 2412
rect -27480 2378 -27446 2412
rect -27412 2378 -27378 2412
rect -27344 2378 -27310 2412
rect -27276 2378 -27242 2412
rect -27208 2378 -27174 2412
rect -27140 2378 -27106 2412
rect -27072 2378 -27036 2412
rect -29114 2348 -27036 2378
rect -29148 2343 -27036 2348
rect -29148 2314 -29078 2343
rect -29114 2309 -29078 2314
rect -29044 2309 -29010 2343
rect -28976 2309 -28942 2343
rect -28908 2309 -28874 2343
rect -28840 2309 -28806 2343
rect -28772 2309 -28738 2343
rect -28704 2309 -28670 2343
rect -28636 2309 -28602 2343
rect -28568 2309 -28534 2343
rect -28500 2309 -28466 2343
rect -28432 2309 -28398 2343
rect -28364 2309 -28330 2343
rect -28296 2309 -28262 2343
rect -28228 2309 -28194 2343
rect -28160 2309 -28126 2343
rect -28092 2309 -28058 2343
rect -28024 2309 -27990 2343
rect -27956 2309 -27922 2343
rect -27888 2309 -27854 2343
rect -27820 2309 -27786 2343
rect -27752 2309 -27718 2343
rect -27684 2309 -27650 2343
rect -27616 2309 -27582 2343
rect -27548 2309 -27514 2343
rect -27480 2309 -27446 2343
rect -27412 2309 -27378 2343
rect -27344 2309 -27310 2343
rect -27276 2309 -27242 2343
rect -27208 2309 -27174 2343
rect -27140 2309 -27106 2343
rect -27072 2309 -27036 2343
rect -29114 2280 -27036 2309
rect -29148 2274 -27036 2280
rect -29148 2246 -29078 2274
rect -29114 2240 -29078 2246
rect -29044 2240 -29010 2274
rect -28976 2240 -28942 2274
rect -28908 2240 -28874 2274
rect -28840 2240 -28806 2274
rect -28772 2240 -28738 2274
rect -28704 2240 -28670 2274
rect -28636 2240 -28602 2274
rect -28568 2240 -28534 2274
rect -28500 2240 -28466 2274
rect -28432 2240 -28398 2274
rect -28364 2240 -28330 2274
rect -28296 2240 -28262 2274
rect -28228 2240 -28194 2274
rect -28160 2240 -28126 2274
rect -28092 2240 -28058 2274
rect -28024 2240 -27990 2274
rect -27956 2240 -27922 2274
rect -27888 2240 -27854 2274
rect -27820 2240 -27786 2274
rect -27752 2240 -27718 2274
rect -27684 2240 -27650 2274
rect -27616 2240 -27582 2274
rect -27548 2240 -27514 2274
rect -27480 2240 -27446 2274
rect -27412 2240 -27378 2274
rect -27344 2240 -27310 2274
rect -27276 2240 -27242 2274
rect -27208 2240 -27174 2274
rect -27140 2240 -27106 2274
rect -27072 2240 -27036 2274
rect -29114 2212 -27036 2240
rect -29148 2205 -27036 2212
rect -29148 2178 -29078 2205
rect -29114 2171 -29078 2178
rect -29044 2171 -29010 2205
rect -28976 2171 -28942 2205
rect -28908 2171 -28874 2205
rect -28840 2171 -28806 2205
rect -28772 2171 -28738 2205
rect -28704 2171 -28670 2205
rect -28636 2171 -28602 2205
rect -28568 2171 -28534 2205
rect -28500 2171 -28466 2205
rect -28432 2171 -28398 2205
rect -28364 2171 -28330 2205
rect -28296 2171 -28262 2205
rect -28228 2171 -28194 2205
rect -28160 2171 -28126 2205
rect -28092 2171 -28058 2205
rect -28024 2171 -27990 2205
rect -27956 2171 -27922 2205
rect -27888 2171 -27854 2205
rect -27820 2171 -27786 2205
rect -27752 2171 -27718 2205
rect -27684 2171 -27650 2205
rect -27616 2171 -27582 2205
rect -27548 2171 -27514 2205
rect -27480 2171 -27446 2205
rect -27412 2171 -27378 2205
rect -27344 2171 -27310 2205
rect -27276 2171 -27242 2205
rect -27208 2171 -27174 2205
rect -27140 2171 -27106 2205
rect -27072 2171 -27036 2205
rect -29114 2144 -27036 2171
rect -29148 2136 -27036 2144
rect -29148 2110 -29078 2136
rect -29114 2102 -29078 2110
rect -29044 2102 -29010 2136
rect -28976 2102 -28942 2136
rect -28908 2102 -28874 2136
rect -28840 2102 -28806 2136
rect -28772 2102 -28738 2136
rect -28704 2102 -28670 2136
rect -28636 2102 -28602 2136
rect -28568 2102 -28534 2136
rect -28500 2102 -28466 2136
rect -28432 2102 -28398 2136
rect -28364 2102 -28330 2136
rect -28296 2102 -28262 2136
rect -28228 2102 -28194 2136
rect -28160 2102 -28126 2136
rect -28092 2102 -28058 2136
rect -28024 2102 -27990 2136
rect -27956 2102 -27922 2136
rect -27888 2102 -27854 2136
rect -27820 2102 -27786 2136
rect -27752 2102 -27718 2136
rect -27684 2102 -27650 2136
rect -27616 2102 -27582 2136
rect -27548 2102 -27514 2136
rect -27480 2102 -27446 2136
rect -27412 2102 -27378 2136
rect -27344 2102 -27310 2136
rect -27276 2102 -27242 2136
rect -27208 2102 -27174 2136
rect -27140 2102 -27106 2136
rect -27072 2102 -27036 2136
rect -29114 2076 -27036 2102
rect -29148 2067 -27036 2076
rect -29148 2042 -29078 2067
rect -29114 2008 -29078 2042
rect -29148 1974 -29078 2008
rect -29114 1940 -29078 1974
rect -29148 1906 -29078 1940
rect -29114 1872 -29078 1906
rect -29148 1838 -29078 1872
rect -29114 1804 -29078 1838
rect -29148 1770 -29078 1804
rect -29114 1736 -29078 1770
rect -29148 1702 -29078 1736
rect -29114 1668 -29078 1702
rect -29148 1634 -29078 1668
rect -29114 1600 -29078 1634
rect -29148 1566 -29078 1600
rect -29114 1532 -29078 1566
rect -29148 1498 -29078 1532
rect -29114 1464 -29078 1498
rect -29148 1430 -29078 1464
rect -29114 1396 -29078 1430
rect -29148 1362 -29078 1396
rect -29114 1328 -29078 1362
rect -29148 1294 -29078 1328
rect -29114 1260 -29078 1294
rect -29148 1226 -29078 1260
rect -29114 1192 -29078 1226
rect -29148 1158 -29078 1192
rect -29114 1124 -29078 1158
rect -29148 1090 -29078 1124
rect -29114 1056 -29078 1090
rect -29148 1022 -29078 1056
rect -29114 988 -29078 1022
rect -29148 954 -29078 988
rect -29114 920 -29078 954
rect -29148 886 -29078 920
rect -29114 852 -29078 886
rect -29148 818 -29078 852
rect -29114 784 -29078 818
rect -29148 750 -29078 784
rect -29114 716 -29078 750
rect -29148 682 -29078 716
rect -29114 648 -29078 682
rect -29148 614 -29078 648
rect -29114 580 -29078 614
rect -29148 546 -29078 580
rect -29114 512 -29078 546
rect -29148 478 -29078 512
rect -29114 444 -29078 478
rect -29148 410 -29078 444
rect -29114 376 -29078 410
rect -29148 342 -29078 376
rect -29114 308 -29078 342
rect -29148 274 -29078 308
rect -29114 240 -29078 274
rect -29148 206 -29078 240
rect -29114 172 -29078 206
rect -29148 138 -29078 172
rect -29114 104 -29078 138
rect -29148 70 -29078 104
rect -29114 36 -29078 70
rect -29148 2 -29078 36
rect -29114 -32 -29078 2
rect -29148 -66 -29078 -32
rect -29114 -100 -29078 -66
rect -29148 -134 -29078 -100
rect -29114 -168 -29078 -134
rect -29148 -202 -29078 -168
rect -29114 -236 -29078 -202
rect -29148 -270 -29078 -236
rect -29114 -304 -29078 -270
rect -29148 -338 -29078 -304
rect -29114 -372 -29078 -338
rect -29148 -406 -29078 -372
rect -29114 -440 -29078 -406
rect -29148 -474 -29078 -440
rect -29114 -508 -29078 -474
rect -29148 -542 -29078 -508
rect -29114 -576 -29078 -542
rect -29148 -610 -29078 -576
rect -29114 -644 -29078 -610
rect -29148 -678 -29078 -644
rect -29114 -712 -29078 -678
rect -29148 -746 -29078 -712
rect -29114 -780 -29078 -746
rect -29148 -814 -29078 -780
rect -29114 -848 -29078 -814
rect -29148 -882 -29078 -848
rect -29114 -916 -29078 -882
rect -29148 -950 -29078 -916
rect -29114 -984 -29078 -950
rect -29148 -1018 -29078 -984
rect -29114 -1052 -29078 -1018
rect -29148 -1086 -29078 -1052
rect -29114 -1120 -29078 -1086
rect -29148 -1154 -29078 -1120
rect -29114 -1188 -29078 -1154
rect -29148 -1222 -29078 -1188
rect -29114 -1256 -29078 -1222
rect -29148 -1290 -29078 -1256
rect -29114 -1324 -29078 -1290
rect -29148 -1358 -29078 -1324
rect -29114 -1392 -29078 -1358
rect -29148 -1426 -29078 -1392
rect -29114 -1460 -29078 -1426
rect -29148 -1494 -29078 -1460
rect -29114 -1528 -29078 -1494
rect -29148 -1562 -29078 -1528
rect -29114 -1596 -29078 -1562
rect -29148 -1630 -29078 -1596
rect -29114 -1664 -29078 -1630
rect -29148 -1698 -29078 -1664
rect -29114 -1732 -29078 -1698
rect -29148 -1766 -29078 -1732
rect -29114 -1800 -29078 -1766
rect -29148 -1834 -29078 -1800
rect -29114 -1868 -29078 -1834
rect -29148 -1902 -29078 -1868
rect -29114 -1936 -29078 -1902
rect -29148 -1970 -29078 -1936
rect -29114 -2004 -29078 -1970
rect -29148 -2038 -29078 -2004
rect -29114 -2072 -29078 -2038
rect -29148 -2106 -29078 -2072
rect -29114 -2140 -29078 -2106
rect -29148 -2174 -29078 -2140
rect -29114 -2208 -29078 -2174
rect -29148 -2242 -29078 -2208
rect -29114 -2276 -29078 -2242
rect -29148 -2310 -29078 -2276
rect -29114 -2344 -29078 -2310
rect -29148 -2378 -29078 -2344
rect -29114 -2412 -29078 -2378
rect -29148 -2446 -29078 -2412
rect -29114 -2480 -29078 -2446
rect -29148 -2514 -29078 -2480
rect -29114 -2548 -29078 -2514
rect -29148 -2582 -29078 -2548
rect -29114 -2616 -29078 -2582
rect -29148 -2650 -29078 -2616
rect -29114 -2684 -29078 -2650
rect -29148 -2718 -29078 -2684
rect -29114 -2752 -29078 -2718
rect -29148 -2786 -29078 -2752
rect -29114 -2820 -29078 -2786
rect -29148 -2854 -29078 -2820
rect -29114 -2888 -29078 -2854
rect -29148 -2922 -29078 -2888
rect -29114 -2956 -29078 -2922
rect -29148 -2990 -29078 -2956
rect -29114 -3024 -29078 -2990
rect -29148 -3058 -29078 -3024
rect -29114 -3092 -29078 -3058
rect -29148 -3126 -29078 -3092
rect -29114 -3160 -29078 -3126
rect -29148 -3194 -29078 -3160
rect -29114 -3228 -29078 -3194
rect -29148 -3262 -29078 -3228
rect -29114 -3296 -29078 -3262
rect -29148 -3330 -29078 -3296
rect -29114 -3364 -29078 -3330
rect -29148 -3398 -29078 -3364
rect -29114 -3432 -29078 -3398
rect -29148 -3466 -29078 -3432
rect -29114 -3500 -29078 -3466
rect -29148 -3534 -29078 -3500
rect -29114 -3568 -29078 -3534
rect -29148 -3602 -29078 -3568
rect -29114 -3636 -29078 -3602
rect -29148 -3670 -29078 -3636
rect -29114 -3704 -29078 -3670
rect -29148 -3738 -29078 -3704
rect -29114 -3772 -29078 -3738
rect -29148 -3806 -29078 -3772
rect -29114 -3840 -29078 -3806
rect -29148 -3874 -29078 -3840
rect -29114 -3908 -29078 -3874
rect -29148 -3942 -29078 -3908
rect -29114 -3976 -29078 -3942
rect -29148 -4010 -29078 -3976
rect -29114 -4044 -29078 -4010
rect -29148 -4078 -29078 -4044
rect -29114 -4112 -29078 -4078
rect -29148 -4146 -29078 -4112
rect -29114 -4180 -29078 -4146
rect -29148 -4214 -29078 -4180
rect -29114 -4248 -29078 -4214
rect -29148 -4282 -29078 -4248
rect -29114 -4316 -29078 -4282
rect -29148 -4350 -29078 -4316
rect -29114 -4384 -29078 -4350
rect -29148 -4418 -29078 -4384
rect -29114 -4452 -29078 -4418
rect -29148 -4486 -29078 -4452
rect -29114 -4520 -29078 -4486
rect -29148 -4554 -29078 -4520
rect -29114 -4588 -29078 -4554
rect -29148 -4622 -29078 -4588
rect -29114 -4656 -29078 -4622
rect -29148 -4690 -29078 -4656
rect -29114 -4724 -29078 -4690
rect -29148 -4758 -29078 -4724
rect -29114 -4792 -29078 -4758
rect -29148 -4826 -29078 -4792
rect -29114 -4860 -29078 -4826
rect -29148 -4894 -29078 -4860
rect -29114 -4928 -29078 -4894
rect -29148 -4962 -29078 -4928
rect -29114 -4996 -29078 -4962
rect -29148 -5030 -29078 -4996
rect -29114 -5064 -29078 -5030
rect -29148 -5098 -29078 -5064
rect -29114 -5132 -29078 -5098
rect -29148 -5166 -29078 -5132
rect -29114 -5200 -29078 -5166
rect -29148 -5234 -29078 -5200
rect -29114 -5268 -29078 -5234
rect -29148 -5302 -29078 -5268
rect -29114 -5336 -29078 -5302
rect -29148 -5370 -29078 -5336
rect -29114 -5404 -29078 -5370
rect -29148 -5438 -29078 -5404
rect -29114 -5472 -29078 -5438
rect -29148 -5506 -29078 -5472
rect -29114 -5540 -29078 -5506
rect -29148 -5574 -29078 -5540
rect -29114 -5608 -29078 -5574
rect -29148 -5642 -29078 -5608
rect -29114 -5676 -29078 -5642
rect -29148 -5710 -29078 -5676
rect -29114 -5744 -29078 -5710
rect -29148 -5778 -29078 -5744
rect -29114 -5812 -29078 -5778
rect -29148 -5846 -29078 -5812
rect -29114 -5880 -29078 -5846
rect -29148 -5914 -29078 -5880
rect -29114 -5948 -29078 -5914
rect -29148 -5982 -29078 -5948
rect -29114 -6016 -29078 -5982
rect -29148 -6050 -29078 -6016
rect -29114 -6084 -29078 -6050
rect -29148 -6118 -29078 -6084
rect -29114 -6152 -29078 -6118
rect -29148 -6186 -29078 -6152
rect -29114 -6220 -29078 -6186
rect -29148 -6254 -29078 -6220
rect -29114 -6288 -29078 -6254
rect -29148 -6322 -29078 -6288
rect -29114 -6356 -29078 -6322
rect -29148 -6390 -29078 -6356
rect -29114 -6424 -29078 -6390
rect -29148 -6458 -29078 -6424
rect -29114 -6492 -29078 -6458
rect -29148 -6526 -29078 -6492
rect -29114 -6560 -29078 -6526
rect -29148 -6594 -29078 -6560
rect -29114 -6628 -29078 -6594
rect -29148 -6662 -29078 -6628
rect -29114 -6696 -29078 -6662
rect -29148 -6730 -29078 -6696
rect -29114 -6764 -29078 -6730
rect -29148 -6798 -29078 -6764
rect -29114 -6832 -29078 -6798
rect -29148 -6866 -29078 -6832
rect -29114 -6900 -29078 -6866
rect -29148 -6934 -29078 -6900
rect -29114 -6968 -29078 -6934
rect -29148 -7002 -29078 -6968
rect -29114 -7036 -29078 -7002
rect -29148 -7070 -29078 -7036
rect -29114 -7104 -29078 -7070
rect -29148 -7138 -29078 -7104
rect -29114 -7172 -29078 -7138
rect -29148 -7206 -29078 -7172
rect -29114 -7240 -29078 -7206
rect -29148 -7274 -29078 -7240
rect -29114 -7308 -29078 -7274
rect -29148 -7342 -29078 -7308
rect -29114 -7376 -29078 -7342
rect -29148 -7410 -29078 -7376
rect -29114 -7444 -29078 -7410
rect -29148 -7478 -29078 -7444
rect -29114 -7512 -29078 -7478
rect -29148 -7546 -29078 -7512
rect -29114 -7580 -29078 -7546
rect -29148 -7614 -29078 -7580
rect -29114 -7648 -29078 -7614
rect -29148 -7682 -29078 -7648
rect -29114 -7716 -29078 -7682
rect -29148 -7750 -29078 -7716
rect -29114 -7784 -29078 -7750
rect -29148 -7818 -29078 -7784
rect -29114 -7852 -29078 -7818
rect -29148 -7886 -29078 -7852
rect -29114 -7920 -29078 -7886
rect -29148 -7954 -29078 -7920
rect -29114 -7988 -29078 -7954
rect -29148 -8022 -29078 -7988
rect -29114 -8056 -29078 -8022
rect -29148 -8090 -29078 -8056
rect -29114 -8124 -29078 -8090
rect -29148 -8158 -29078 -8124
rect -29114 -8192 -29078 -8158
rect -29148 -8226 -29078 -8192
rect -29114 -8260 -29078 -8226
rect -29148 -8294 -29078 -8260
rect -29114 -8328 -29078 -8294
rect -29148 -8362 -29078 -8328
rect -29114 -8396 -29078 -8362
rect -29148 -8430 -29078 -8396
rect -29114 -8464 -29078 -8430
rect -29148 -8498 -29078 -8464
rect -29114 -8532 -29078 -8498
rect -29148 -8566 -29078 -8532
rect -29114 -8600 -29078 -8566
rect -29148 -8634 -29078 -8600
rect -29114 -8668 -29078 -8634
rect -29148 -8702 -29078 -8668
rect -29114 -8736 -29078 -8702
rect -31669 -8779 -31632 -8745
rect -31669 -8813 -31598 -8779
rect -29148 -8813 -29078 -8736
rect -31669 -8847 -31528 -8813
rect -31494 -8847 -31460 -8813
rect -31426 -8847 -31392 -8813
rect -31358 -8847 -31324 -8813
rect -31290 -8847 -31256 -8813
rect -31222 -8847 -31188 -8813
rect -31154 -8847 -31120 -8813
rect -31086 -8847 -31052 -8813
rect -31018 -8847 -30984 -8813
rect -30950 -8847 -30916 -8813
rect -30882 -8847 -30848 -8813
rect -30814 -8847 -30780 -8813
rect -30746 -8847 -30712 -8813
rect -30678 -8847 -30644 -8813
rect -30610 -8847 -30576 -8813
rect -30542 -8847 -30508 -8813
rect -30474 -8847 -30440 -8813
rect -30406 -8847 -30372 -8813
rect -30338 -8847 -30304 -8813
rect -30270 -8847 -30236 -8813
rect -30202 -8847 -30168 -8813
rect -30134 -8847 -30100 -8813
rect -30066 -8847 -30032 -8813
rect -29998 -8847 -29964 -8813
rect -29930 -8847 -29896 -8813
rect -29862 -8847 -29828 -8813
rect -29794 -8847 -29760 -8813
rect -29726 -8847 -29692 -8813
rect -29658 -8847 -29624 -8813
rect -29590 -8847 -29556 -8813
rect -29522 -8847 -29488 -8813
rect -29454 -8847 -29420 -8813
rect -29386 -8847 -29352 -8813
rect -29318 -8847 -29284 -8813
rect -29250 -8847 -29216 -8813
rect -29182 -8847 -29078 -8813
rect -27072 -8847 -27036 2067
rect 5738 3432 5772 3433
rect 5738 3364 5772 3398
rect 5738 3296 5772 3330
rect 5738 3228 5772 3262
rect 5738 3160 5772 3194
rect 5738 3092 5772 3126
rect 5738 3024 5772 3058
rect 5738 2956 5772 2990
rect 5738 2888 5772 2922
rect 5738 2820 5772 2854
rect 5738 2752 5772 2786
rect 5738 2684 5772 2718
rect 5738 2616 5772 2650
rect 5738 2548 5772 2582
rect 5738 2509 5772 2514
rect -31669 -8884 -27036 -8847
rect -31669 -9598 -31632 -8884
rect -27450 -8918 -27415 -8884
rect -27381 -8918 -27346 -8884
rect -27312 -8918 -27277 -8884
rect -27243 -8918 -27208 -8884
rect -27174 -8918 -27139 -8884
rect -27105 -8918 -27070 -8884
rect -27450 -8952 -27036 -8918
rect -27450 -8986 -27415 -8952
rect -27381 -8986 -27346 -8952
rect -27312 -8986 -27277 -8952
rect -27243 -8986 -27208 -8952
rect -27174 -8986 -27139 -8952
rect -27105 -8986 -27070 -8952
rect -27450 -9020 -27036 -8986
rect -27450 -9054 -27415 -9020
rect -27381 -9054 -27346 -9020
rect -27312 -9054 -27277 -9020
rect -27243 -9054 -27208 -9020
rect -27174 -9054 -27139 -9020
rect -27105 -9054 -27070 -9020
rect -27450 -9088 -27036 -9054
rect -27450 -9122 -27415 -9088
rect -27381 -9122 -27346 -9088
rect -27312 -9122 -27277 -9088
rect -27243 -9122 -27208 -9088
rect -27174 -9122 -27139 -9088
rect -27105 -9122 -27070 -9088
rect -27450 -9156 -27036 -9122
rect -27450 -9190 -27415 -9156
rect -27381 -9190 -27346 -9156
rect -27312 -9190 -27277 -9156
rect -27243 -9190 -27208 -9156
rect -27174 -9190 -27139 -9156
rect -27105 -9190 -27070 -9156
rect -27450 -9224 -27036 -9190
rect -27450 -9258 -27415 -9224
rect -27381 -9258 -27346 -9224
rect -27312 -9258 -27277 -9224
rect -27243 -9258 -27208 -9224
rect -27174 -9258 -27139 -9224
rect -27105 -9258 -27070 -9224
rect -27450 -9292 -27036 -9258
rect -27450 -9326 -27415 -9292
rect -27381 -9326 -27346 -9292
rect -27312 -9326 -27277 -9292
rect -27243 -9326 -27208 -9292
rect -27174 -9326 -27139 -9292
rect -27105 -9326 -27070 -9292
rect -27450 -9360 -27036 -9326
rect -27450 -9394 -27415 -9360
rect -27381 -9394 -27346 -9360
rect -27312 -9394 -27277 -9360
rect -27243 -9394 -27208 -9360
rect -27174 -9394 -27139 -9360
rect -27105 -9394 -27070 -9360
rect -27450 -9428 -27036 -9394
rect -27450 -9462 -27415 -9428
rect -27381 -9462 -27346 -9428
rect -27312 -9462 -27277 -9428
rect -27243 -9462 -27208 -9428
rect -27174 -9462 -27139 -9428
rect -27105 -9462 -27070 -9428
rect -27450 -9496 -27036 -9462
rect -27450 -9530 -27415 -9496
rect -27381 -9530 -27346 -9496
rect -27312 -9530 -27277 -9496
rect -27243 -9530 -27208 -9496
rect -27174 -9530 -27139 -9496
rect -27105 -9530 -27070 -9496
rect -27450 -9564 -27036 -9530
rect -27450 -9598 -27415 -9564
rect -27381 -9598 -27346 -9564
rect -27312 -9598 -27277 -9564
rect -27243 -9598 -27208 -9564
rect -27174 -9598 -27139 -9564
rect -27105 -9598 -27070 -9564
rect -31669 -9635 -27036 -9598
<< mvnsubdiff >>
rect -757 3654 -733 3688
rect -699 3654 -662 3688
rect -628 3654 -591 3688
rect -557 3654 -519 3688
rect -485 3654 -447 3688
rect -413 3654 -389 3688
rect 157 3654 181 3688
rect 215 3654 250 3688
rect 284 3654 319 3688
rect 353 3654 388 3688
rect 422 3654 457 3688
rect 491 3654 526 3688
rect 560 3654 595 3688
rect 629 3654 664 3688
rect 698 3654 733 3688
rect 767 3654 802 3688
rect 836 3654 871 3688
rect 905 3654 940 3688
rect 974 3654 1009 3688
rect 1043 3654 1078 3688
rect 1112 3654 1147 3688
rect 1181 3654 1216 3688
rect 1250 3654 1285 3688
rect 1319 3654 1354 3688
rect 1388 3654 1423 3688
rect 1457 3654 1492 3688
rect 1526 3654 1561 3688
rect 1595 3654 1630 3688
rect 1664 3654 1699 3688
rect 1733 3654 1768 3688
rect 1802 3654 1837 3688
rect 1871 3654 1906 3688
rect 1940 3654 1975 3688
rect 2009 3654 2044 3688
rect 2078 3654 2113 3688
rect 2147 3654 2182 3688
rect 2216 3654 2251 3688
rect 2285 3654 2320 3688
rect 2354 3654 2389 3688
rect 2423 3654 2458 3688
rect 2492 3654 2527 3688
rect 2561 3654 2596 3688
rect 2630 3654 2665 3688
rect 2699 3654 2734 3688
rect 2768 3654 2803 3688
rect 2837 3654 2872 3688
rect 2906 3654 2941 3688
rect 2975 3654 3010 3688
rect 3044 3654 3078 3688
rect 3112 3654 3146 3688
rect 3180 3654 3214 3688
rect 3248 3654 3282 3688
rect 3316 3654 3350 3688
rect 3384 3654 3418 3688
rect 3452 3654 3486 3688
rect 3520 3654 3544 3688
rect 6732 3301 6766 3325
rect 6732 3227 6766 3267
rect 6732 3153 6766 3193
rect 6732 3079 6766 3119
rect 6732 3005 6766 3045
rect 6732 2931 6766 2971
rect 6732 2858 6766 2897
rect 6732 2785 6766 2824
rect 6732 2712 6766 2751
rect 6732 2639 6766 2678
rect 6732 2581 6766 2605
<< psubdiffcont >>
rect 4106 3806 4140 3840
rect 4174 3806 4208 3840
rect 4242 3806 4276 3840
rect 4310 3806 4344 3840
rect 4378 3806 4412 3840
rect 4446 3806 4480 3840
rect 4514 3806 4548 3840
rect 4582 3806 4616 3840
rect 4650 3806 4684 3840
rect 4718 3806 4752 3840
rect 4786 3806 4820 3840
rect 4854 3806 4888 3840
rect 4922 3806 4956 3840
rect 4990 3806 5024 3840
rect 5058 3806 5092 3840
rect 5126 3806 5160 3840
rect 5194 3806 5228 3840
rect 5262 3806 5296 3840
rect 5330 3806 5364 3840
rect 5398 3806 5432 3840
rect 5466 3806 5500 3840
rect 5534 3806 5568 3840
rect 5602 3806 5636 3840
rect 5670 3806 5704 3840
rect 3938 3700 3972 3734
rect 3938 3632 3972 3666
rect 4723 3738 4757 3772
rect 4815 3738 4849 3772
rect 4907 3738 4941 3772
rect 4723 3669 4757 3703
rect 4815 3669 4849 3703
rect 4907 3669 4941 3703
rect 3938 3564 3972 3598
rect 3938 3496 3972 3530
rect 3938 3428 3972 3462
rect 3938 3360 3972 3394
rect 3938 3292 3972 3326
rect 3938 3224 3972 3258
rect 3938 3156 3972 3190
rect 3938 3088 3972 3122
rect 3938 3020 3972 3054
rect 3938 2952 3972 2986
rect 3938 2884 3972 2918
rect 3938 2816 3972 2850
rect 3938 2748 3972 2782
rect 3938 2680 3972 2714
rect 3938 2612 3972 2646
rect 3938 2544 3972 2578
rect 3938 2476 3972 2510
rect 3938 2408 3972 2442
rect 3938 2340 3972 2374
rect 3938 2272 3972 2306
rect 5738 3738 5772 3772
rect 5738 3670 5772 3704
rect 4723 3600 4757 3634
rect 4815 3600 4849 3634
rect 4907 3600 4941 3634
rect 4723 3531 4757 3565
rect 4815 3531 4849 3565
rect 4907 3531 4941 3565
rect 4723 3462 4757 3496
rect 4815 3462 4849 3496
rect 4907 3462 4941 3496
rect 4723 3393 4757 3427
rect 4815 3393 4849 3427
rect 4907 3393 4941 3427
rect 4723 3324 4757 3358
rect 4815 3324 4849 3358
rect 4907 3324 4941 3358
rect 4723 3255 4757 3289
rect 4815 3255 4849 3289
rect 4907 3255 4941 3289
rect 4723 3186 4757 3220
rect 4815 3186 4849 3220
rect 4907 3186 4941 3220
rect 4723 3116 4757 3150
rect 4815 3116 4849 3150
rect 4907 3116 4941 3150
rect 4723 3046 4757 3080
rect 4815 3046 4849 3080
rect 4907 3046 4941 3080
rect 4723 2976 4757 3010
rect 4815 2976 4849 3010
rect 4907 2976 4941 3010
rect 4723 2906 4757 2940
rect 4815 2906 4849 2940
rect 4907 2906 4941 2940
rect 4723 2836 4757 2870
rect 4815 2836 4849 2870
rect 4907 2836 4941 2870
rect 4723 2766 4757 2800
rect 4815 2766 4849 2800
rect 4907 2766 4941 2800
rect 4723 2696 4757 2730
rect 4815 2696 4849 2730
rect 4907 2696 4941 2730
rect 4723 2626 4757 2660
rect 4815 2626 4849 2660
rect 4907 2626 4941 2660
rect 4723 2556 4757 2590
rect 4815 2556 4849 2590
rect 4907 2556 4941 2590
rect 4723 2486 4757 2520
rect 4815 2486 4849 2520
rect 4907 2486 4941 2520
rect 4723 2416 4757 2450
rect 4815 2416 4849 2450
rect 4907 2416 4941 2450
rect 4723 2346 4757 2380
rect 4815 2346 4849 2380
rect 4907 2346 4941 2380
rect 4723 2276 4757 2310
rect 4815 2276 4849 2310
rect 4907 2276 4941 2310
rect 3938 2204 3972 2238
rect 3938 2136 3972 2170
rect 5738 3602 5772 3636
rect 5738 3534 5772 3568
rect 5738 3466 5772 3500
rect 4723 2206 4757 2240
rect 4815 2206 4849 2240
rect 4907 2206 4941 2240
rect 4723 2136 4757 2170
rect 4815 2136 4849 2170
rect 4907 2136 4941 2170
rect 4038 2068 4072 2102
rect 4106 2068 4140 2102
rect 4174 2068 4208 2102
rect 4242 2068 4276 2102
rect 4310 2068 4344 2102
rect 4378 2068 4412 2102
rect 4446 2068 4480 2102
rect 4514 2068 4548 2102
rect 4582 2068 4616 2102
rect 4650 2068 4684 2102
rect 4718 2068 4752 2102
rect 4786 2068 4820 2102
rect 4854 2068 4888 2102
rect 4922 2068 4956 2102
rect 4990 2068 5024 2102
rect 5058 2068 5092 2102
rect 5126 2068 5160 2102
rect 5194 2068 5228 2102
rect 5262 2068 5296 2102
rect 5330 2068 5364 2102
rect 5398 2068 5432 2102
rect 5466 2068 5500 2102
rect 5534 2068 5568 2102
rect 5602 2068 5636 2102
rect 5670 2068 5704 2102
rect 168 793 202 827
rect 237 793 271 827
rect 306 793 340 827
rect 375 793 409 827
rect 444 793 478 827
rect 513 793 547 827
rect 582 793 616 827
rect 651 793 685 827
rect 720 793 754 827
rect 789 793 823 827
rect 858 793 892 827
rect 927 793 961 827
rect 996 793 1030 827
rect 1065 793 1099 827
rect 1134 793 1168 827
rect 1203 793 1237 827
rect 1272 793 1306 827
rect 1341 793 1375 827
rect 1410 793 1444 827
rect 1479 793 1513 827
rect 1548 793 1582 827
rect 1617 793 1651 827
rect 1686 793 1720 827
rect 1755 793 1789 827
rect 1824 793 1858 827
rect 1893 793 1927 827
rect 1962 793 1996 827
rect 2031 793 2065 827
rect 2100 793 2134 827
rect 2169 793 2203 827
rect 2238 793 2272 827
rect 2307 793 2341 827
rect 2376 793 2410 827
rect 2445 793 2479 827
rect 2514 793 2548 827
rect 2583 793 2617 827
rect 2652 793 2686 827
rect 2721 793 2755 827
rect 2790 793 2824 827
rect 2859 793 2893 827
rect 2928 793 2962 827
rect 2996 793 3030 827
rect 3064 793 3098 827
rect 3132 793 3166 827
rect 3200 793 3234 827
rect 3268 793 3302 827
rect 3336 793 3370 827
<< nsubdiffcont >>
rect 4293 3619 4327 3653
rect 4361 3619 4395 3653
rect 4429 3619 4463 3653
rect 4125 3547 4159 3581
rect 4529 3551 4563 3585
rect 4125 3479 4159 3513
rect 4125 3411 4159 3445
rect 4125 3343 4159 3377
rect 4125 3275 4159 3309
rect 4125 3207 4159 3241
rect 4125 3139 4159 3173
rect 4125 3071 4159 3105
rect 4125 3003 4159 3037
rect 4125 2935 4159 2969
rect 4125 2867 4159 2901
rect 4125 2799 4159 2833
rect 4125 2731 4159 2765
rect 4125 2663 4159 2697
rect 4125 2595 4159 2629
rect 4125 2527 4159 2561
rect 4529 3483 4563 3517
rect 4529 3415 4563 3449
rect 4529 3347 4563 3381
rect 4529 3279 4563 3313
rect 4529 3211 4563 3245
rect 4529 3143 4563 3177
rect 4529 3075 4563 3109
rect 4529 3007 4563 3041
rect 4529 2939 4563 2973
rect 4529 2871 4563 2905
rect 4529 2803 4563 2837
rect 4529 2735 4563 2769
rect 4529 2667 4563 2701
rect 4529 2599 4563 2633
rect 4125 2459 4159 2493
rect 4125 2391 4159 2425
rect 4529 2531 4563 2565
rect 4529 2463 4563 2497
rect 4529 2395 4563 2429
rect 4125 2323 4159 2357
rect 4529 2327 4563 2361
rect 4257 2255 4291 2289
rect 4325 2255 4359 2289
rect 4393 2255 4427 2289
rect 4461 2255 4495 2289
rect 5197 3619 5231 3653
rect 5265 3619 5299 3653
rect 5333 3619 5367 3653
rect 5483 3619 5517 3653
rect 5097 3551 5131 3585
rect 5551 3547 5585 3581
rect 5097 3483 5131 3517
rect 5097 3415 5131 3449
rect 5097 3347 5131 3381
rect 5097 3279 5131 3313
rect 5551 3479 5585 3513
rect 5551 3411 5585 3445
rect 5551 3343 5585 3377
rect 5097 3211 5131 3245
rect 5097 3143 5131 3177
rect 5097 3075 5131 3109
rect 5551 3275 5585 3309
rect 5551 3207 5585 3241
rect 5551 3139 5585 3173
rect 5097 3007 5131 3041
rect 5551 3071 5585 3105
rect 5551 3003 5585 3037
rect 5097 2939 5131 2973
rect 5097 2871 5131 2905
rect 5097 2803 5131 2837
rect 5551 2935 5585 2969
rect 5551 2867 5585 2901
rect 5551 2799 5585 2833
rect 5097 2735 5131 2769
rect 5097 2667 5131 2701
rect 5097 2599 5131 2633
rect 5551 2731 5585 2765
rect 5551 2663 5585 2697
rect 5551 2595 5585 2629
rect 5097 2531 5131 2565
rect 5097 2463 5131 2497
rect 5097 2395 5131 2429
rect 5097 2327 5131 2361
rect 5551 2527 5585 2561
rect 5551 2459 5585 2493
rect 5551 2391 5585 2425
rect 5551 2323 5585 2357
rect 5165 2255 5199 2289
rect 5233 2255 5267 2289
rect 5301 2255 5335 2289
rect 5369 2255 5403 2289
rect 5437 2255 5471 2289
<< mvpsubdiffcont >>
rect -32315 4310 -32281 4344
rect -32247 4310 -32213 4344
rect -32179 4310 -32145 4344
rect -32111 4310 -32077 4344
rect -32043 4310 -32009 4344
rect -31975 4310 -31941 4344
rect -31907 4310 -31873 4344
rect -31839 4310 -31805 4344
rect -31771 4310 -31737 4344
rect -31703 4310 -31669 4344
rect -29078 4310 -29044 4344
rect -29010 4310 -28976 4344
rect -28942 4310 -28908 4344
rect -28874 4310 -28840 4344
rect -28806 4310 -28772 4344
rect -28738 4310 -28704 4344
rect -28670 4310 -28636 4344
rect -28602 4310 -28568 4344
rect -28534 4310 -28500 4344
rect -28466 4310 -28432 4344
rect -28398 4310 -28364 4344
rect -28330 4310 -28296 4344
rect -28262 4310 -28228 4344
rect -28194 4310 -28160 4344
rect -28126 4310 -28092 4344
rect -28058 4310 -28024 4344
rect -27990 4310 -27956 4344
rect -27922 4310 -27888 4344
rect -27854 4310 -27820 4344
rect -27786 4310 -27752 4344
rect -27718 4310 -27684 4344
rect -27650 4310 -27616 4344
rect -27582 4310 -27548 4344
rect -27514 4310 -27480 4344
rect -27446 4310 -27412 4344
rect -27378 4310 -27344 4344
rect -27310 4310 -27276 4344
rect -27242 4310 -27208 4344
rect -27174 4310 -27140 4344
rect -27106 4310 -27072 4344
rect -32315 4241 -32281 4275
rect -32247 4241 -32213 4275
rect -32179 4241 -32145 4275
rect -32111 4241 -32077 4275
rect -32043 4241 -32009 4275
rect -31975 4241 -31941 4275
rect -31907 4241 -31873 4275
rect -31839 4241 -31805 4275
rect -31771 4241 -31737 4275
rect -31703 4241 -31669 4275
rect -31632 4242 -31598 4276
rect -31563 4242 -31529 4276
rect -31494 4242 -31460 4276
rect -31425 4242 -31391 4276
rect -31356 4242 -31322 4276
rect -31287 4242 -31253 4276
rect -31218 4242 -31184 4276
rect -31149 4242 -31115 4276
rect -31080 4242 -31046 4276
rect -31011 4242 -30977 4276
rect -30942 4242 -30908 4276
rect -30873 4242 -30839 4276
rect -30804 4242 -30770 4276
rect -30735 4242 -30701 4276
rect -30666 4242 -30632 4276
rect -30597 4242 -30563 4276
rect -30528 4242 -30494 4276
rect -30459 4242 -30425 4276
rect -30390 4242 -30356 4276
rect -30321 4242 -30287 4276
rect -30252 4242 -30218 4276
rect -30183 4242 -30149 4276
rect -30114 4242 -30080 4276
rect -30045 4242 -30011 4276
rect -29976 4242 -29942 4276
rect -29907 4242 -29873 4276
rect -29838 4242 -29804 4276
rect -29769 4242 -29735 4276
rect -29700 4242 -29666 4276
rect -29631 4242 -29597 4276
rect -29562 4242 -29528 4276
rect -29493 4242 -29459 4276
rect -29424 4242 -29390 4276
rect -29355 4242 -29321 4276
rect -29286 4242 -29252 4276
rect -29217 4242 -29183 4276
rect -29148 4242 -29114 4276
rect -29078 4241 -29044 4275
rect -29010 4241 -28976 4275
rect -28942 4241 -28908 4275
rect -28874 4241 -28840 4275
rect -28806 4241 -28772 4275
rect -28738 4241 -28704 4275
rect -28670 4241 -28636 4275
rect -28602 4241 -28568 4275
rect -28534 4241 -28500 4275
rect -28466 4241 -28432 4275
rect -28398 4241 -28364 4275
rect -28330 4241 -28296 4275
rect -28262 4241 -28228 4275
rect -28194 4241 -28160 4275
rect -28126 4241 -28092 4275
rect -28058 4241 -28024 4275
rect -27990 4241 -27956 4275
rect -27922 4241 -27888 4275
rect -27854 4241 -27820 4275
rect -27786 4241 -27752 4275
rect -27718 4241 -27684 4275
rect -27650 4241 -27616 4275
rect -27582 4241 -27548 4275
rect -27514 4241 -27480 4275
rect -27446 4241 -27412 4275
rect -27378 4241 -27344 4275
rect -27310 4241 -27276 4275
rect -27242 4241 -27208 4275
rect -27174 4241 -27140 4275
rect -27106 4241 -27072 4275
rect -32315 4172 -32281 4206
rect -32247 4172 -32213 4206
rect -32179 4172 -32145 4206
rect -32111 4172 -32077 4206
rect -32043 4172 -32009 4206
rect -31975 4172 -31941 4206
rect -31907 4172 -31873 4206
rect -31839 4172 -31805 4206
rect -31771 4172 -31737 4206
rect -31703 4172 -31669 4206
rect -31632 4172 -31598 4206
rect -31563 4172 -31529 4206
rect -31494 4172 -31460 4206
rect -31425 4172 -31391 4206
rect -31356 4172 -31322 4206
rect -31287 4172 -31253 4206
rect -31218 4172 -31184 4206
rect -31149 4172 -31115 4206
rect -31080 4172 -31046 4206
rect -31011 4172 -30977 4206
rect -30942 4172 -30908 4206
rect -30873 4172 -30839 4206
rect -30804 4172 -30770 4206
rect -30735 4172 -30701 4206
rect -30666 4172 -30632 4206
rect -30597 4172 -30563 4206
rect -30528 4172 -30494 4206
rect -30459 4172 -30425 4206
rect -30390 4172 -30356 4206
rect -30321 4172 -30287 4206
rect -30252 4172 -30218 4206
rect -30183 4172 -30149 4206
rect -30114 4172 -30080 4206
rect -30045 4172 -30011 4206
rect -29976 4172 -29942 4206
rect -29907 4172 -29873 4206
rect -29838 4172 -29804 4206
rect -29769 4172 -29735 4206
rect -29700 4172 -29666 4206
rect -29631 4172 -29597 4206
rect -29562 4172 -29528 4206
rect -29493 4172 -29459 4206
rect -29424 4172 -29390 4206
rect -29355 4172 -29321 4206
rect -29286 4172 -29252 4206
rect -29217 4172 -29183 4206
rect -29148 4172 -29114 4206
rect -29078 4172 -29044 4206
rect -29010 4172 -28976 4206
rect -28942 4172 -28908 4206
rect -28874 4172 -28840 4206
rect -28806 4172 -28772 4206
rect -28738 4172 -28704 4206
rect -28670 4172 -28636 4206
rect -28602 4172 -28568 4206
rect -28534 4172 -28500 4206
rect -28466 4172 -28432 4206
rect -28398 4172 -28364 4206
rect -28330 4172 -28296 4206
rect -28262 4172 -28228 4206
rect -28194 4172 -28160 4206
rect -28126 4172 -28092 4206
rect -28058 4172 -28024 4206
rect -27990 4172 -27956 4206
rect -27922 4172 -27888 4206
rect -27854 4172 -27820 4206
rect -27786 4172 -27752 4206
rect -27718 4172 -27684 4206
rect -27650 4172 -27616 4206
rect -27582 4172 -27548 4206
rect -27514 4172 -27480 4206
rect -27446 4172 -27412 4206
rect -27378 4172 -27344 4206
rect -27310 4172 -27276 4206
rect -27242 4172 -27208 4206
rect -27174 4172 -27140 4206
rect -27106 4172 -27072 4206
rect -32315 4103 -32281 4137
rect -32247 4103 -32213 4137
rect -32179 4103 -32145 4137
rect -32111 4103 -32077 4137
rect -32043 4103 -32009 4137
rect -31975 4103 -31941 4137
rect -31907 4103 -31873 4137
rect -31839 4103 -31805 4137
rect -31771 4103 -31737 4137
rect -31703 4103 -31669 4137
rect -31632 4102 -31598 4136
rect -31563 4102 -31529 4136
rect -31494 4102 -31460 4136
rect -31425 4102 -31391 4136
rect -31356 4102 -31322 4136
rect -31287 4102 -31253 4136
rect -31218 4102 -31184 4136
rect -31149 4102 -31115 4136
rect -31080 4102 -31046 4136
rect -31011 4102 -30977 4136
rect -30942 4102 -30908 4136
rect -30873 4102 -30839 4136
rect -30804 4102 -30770 4136
rect -30735 4102 -30701 4136
rect -30666 4102 -30632 4136
rect -30597 4102 -30563 4136
rect -30528 4102 -30494 4136
rect -30459 4102 -30425 4136
rect -30390 4102 -30356 4136
rect -30321 4102 -30287 4136
rect -30252 4102 -30218 4136
rect -30183 4102 -30149 4136
rect -30114 4102 -30080 4136
rect -30045 4102 -30011 4136
rect -29976 4102 -29942 4136
rect -29907 4102 -29873 4136
rect -29838 4102 -29804 4136
rect -29769 4102 -29735 4136
rect -29700 4102 -29666 4136
rect -29631 4102 -29597 4136
rect -29562 4102 -29528 4136
rect -29493 4102 -29459 4136
rect -29424 4102 -29390 4136
rect -29355 4102 -29321 4136
rect -29286 4102 -29252 4136
rect -29217 4102 -29183 4136
rect -29148 4102 -29114 4136
rect -29078 4103 -29044 4137
rect -29010 4103 -28976 4137
rect -28942 4103 -28908 4137
rect -28874 4103 -28840 4137
rect -28806 4103 -28772 4137
rect -28738 4103 -28704 4137
rect -28670 4103 -28636 4137
rect -28602 4103 -28568 4137
rect -28534 4103 -28500 4137
rect -28466 4103 -28432 4137
rect -28398 4103 -28364 4137
rect -28330 4103 -28296 4137
rect -28262 4103 -28228 4137
rect -28194 4103 -28160 4137
rect -28126 4103 -28092 4137
rect -28058 4103 -28024 4137
rect -27990 4103 -27956 4137
rect -27922 4103 -27888 4137
rect -27854 4103 -27820 4137
rect -27786 4103 -27752 4137
rect -27718 4103 -27684 4137
rect -27650 4103 -27616 4137
rect -27582 4103 -27548 4137
rect -27514 4103 -27480 4137
rect -27446 4103 -27412 4137
rect -27378 4103 -27344 4137
rect -27310 4103 -27276 4137
rect -27242 4103 -27208 4137
rect -27174 4103 -27140 4137
rect -27106 4103 -27072 4137
rect -32315 4034 -32281 4068
rect -32247 4034 -32213 4068
rect -32179 4034 -32145 4068
rect -32111 4034 -32077 4068
rect -32043 4034 -32009 4068
rect -31975 4034 -31941 4068
rect -31907 4034 -31873 4068
rect -31839 4034 -31805 4068
rect -31771 4034 -31737 4068
rect -31703 4034 -31669 4068
rect -31632 4032 -31598 4066
rect -31563 4032 -31529 4066
rect -31494 4032 -31460 4066
rect -31425 4032 -31391 4066
rect -31356 4032 -31322 4066
rect -31287 4032 -31253 4066
rect -31218 4032 -31184 4066
rect -31149 4032 -31115 4066
rect -31080 4032 -31046 4066
rect -31011 4032 -30977 4066
rect -30942 4032 -30908 4066
rect -30873 4032 -30839 4066
rect -30804 4032 -30770 4066
rect -30735 4032 -30701 4066
rect -30666 4032 -30632 4066
rect -30597 4032 -30563 4066
rect -30528 4032 -30494 4066
rect -30459 4032 -30425 4066
rect -30390 4032 -30356 4066
rect -30321 4032 -30287 4066
rect -30252 4032 -30218 4066
rect -30183 4032 -30149 4066
rect -30114 4032 -30080 4066
rect -30045 4032 -30011 4066
rect -29976 4032 -29942 4066
rect -29907 4032 -29873 4066
rect -29838 4032 -29804 4066
rect -29769 4032 -29735 4066
rect -29700 4032 -29666 4066
rect -29631 4032 -29597 4066
rect -29562 4032 -29528 4066
rect -29493 4032 -29459 4066
rect -29424 4032 -29390 4066
rect -29355 4032 -29321 4066
rect -29286 4032 -29252 4066
rect -29217 4032 -29183 4066
rect -29148 4032 -29114 4066
rect -29078 4034 -29044 4068
rect -29010 4034 -28976 4068
rect -28942 4034 -28908 4068
rect -28874 4034 -28840 4068
rect -28806 4034 -28772 4068
rect -28738 4034 -28704 4068
rect -28670 4034 -28636 4068
rect -28602 4034 -28568 4068
rect -28534 4034 -28500 4068
rect -28466 4034 -28432 4068
rect -28398 4034 -28364 4068
rect -28330 4034 -28296 4068
rect -28262 4034 -28228 4068
rect -28194 4034 -28160 4068
rect -28126 4034 -28092 4068
rect -28058 4034 -28024 4068
rect -27990 4034 -27956 4068
rect -27922 4034 -27888 4068
rect -27854 4034 -27820 4068
rect -27786 4034 -27752 4068
rect -27718 4034 -27684 4068
rect -27650 4034 -27616 4068
rect -27582 4034 -27548 4068
rect -27514 4034 -27480 4068
rect -27446 4034 -27412 4068
rect -27378 4034 -27344 4068
rect -27310 4034 -27276 4068
rect -27242 4034 -27208 4068
rect -27174 4034 -27140 4068
rect -27106 4034 -27072 4068
rect -32315 -9635 -31669 3999
rect -31632 3962 -31598 3996
rect -31563 3962 -31529 3996
rect -31494 3962 -31460 3996
rect -31425 3962 -31391 3996
rect -31356 3962 -31322 3996
rect -31287 3962 -31253 3996
rect -31218 3962 -31184 3996
rect -31149 3962 -31115 3996
rect -31080 3962 -31046 3996
rect -31011 3962 -30977 3996
rect -30942 3962 -30908 3996
rect -30873 3962 -30839 3996
rect -30804 3962 -30770 3996
rect -30735 3962 -30701 3996
rect -30666 3962 -30632 3996
rect -30597 3962 -30563 3996
rect -30528 3962 -30494 3996
rect -30459 3962 -30425 3996
rect -30390 3962 -30356 3996
rect -30321 3962 -30287 3996
rect -30252 3962 -30218 3996
rect -30183 3962 -30149 3996
rect -30114 3962 -30080 3996
rect -30045 3962 -30011 3996
rect -29976 3962 -29942 3996
rect -29907 3962 -29873 3996
rect -29838 3962 -29804 3996
rect -29769 3962 -29735 3996
rect -29700 3962 -29666 3996
rect -29631 3962 -29597 3996
rect -29562 3962 -29528 3996
rect -29493 3962 -29459 3996
rect -29424 3962 -29390 3996
rect -29355 3962 -29321 3996
rect -29286 3962 -29252 3996
rect -29217 3962 -29183 3996
rect -29148 3962 -29114 3996
rect -29078 3965 -29044 3999
rect -29010 3965 -28976 3999
rect -28942 3965 -28908 3999
rect -28874 3965 -28840 3999
rect -28806 3965 -28772 3999
rect -28738 3965 -28704 3999
rect -28670 3965 -28636 3999
rect -28602 3965 -28568 3999
rect -28534 3965 -28500 3999
rect -28466 3965 -28432 3999
rect -28398 3965 -28364 3999
rect -28330 3965 -28296 3999
rect -28262 3965 -28228 3999
rect -28194 3965 -28160 3999
rect -28126 3965 -28092 3999
rect -28058 3965 -28024 3999
rect -27990 3965 -27956 3999
rect -27922 3965 -27888 3999
rect -27854 3965 -27820 3999
rect -27786 3965 -27752 3999
rect -27718 3965 -27684 3999
rect -27650 3965 -27616 3999
rect -27582 3965 -27548 3999
rect -27514 3965 -27480 3999
rect -27446 3965 -27412 3999
rect -27378 3965 -27344 3999
rect -27310 3965 -27276 3999
rect -27242 3965 -27208 3999
rect -27174 3965 -27140 3999
rect -27106 3965 -27072 3999
rect -31632 3892 -31598 3926
rect -31563 3892 -31529 3926
rect -31494 3892 -31460 3926
rect -31425 3892 -31391 3926
rect -31356 3892 -31322 3926
rect -31287 3892 -31253 3926
rect -31218 3892 -31184 3926
rect -31149 3892 -31115 3926
rect -31080 3892 -31046 3926
rect -31011 3892 -30977 3926
rect -30942 3892 -30908 3926
rect -30873 3892 -30839 3926
rect -30804 3892 -30770 3926
rect -30735 3892 -30701 3926
rect -30666 3892 -30632 3926
rect -30597 3892 -30563 3926
rect -30528 3892 -30494 3926
rect -30459 3892 -30425 3926
rect -30390 3892 -30356 3926
rect -30321 3892 -30287 3926
rect -30252 3892 -30218 3926
rect -30183 3892 -30149 3926
rect -30114 3892 -30080 3926
rect -30045 3892 -30011 3926
rect -29976 3892 -29942 3926
rect -29907 3892 -29873 3926
rect -29838 3892 -29804 3926
rect -29769 3892 -29735 3926
rect -29700 3892 -29666 3926
rect -29631 3892 -29597 3926
rect -29562 3892 -29528 3926
rect -29493 3892 -29459 3926
rect -29424 3892 -29390 3926
rect -29355 3892 -29321 3926
rect -29286 3892 -29252 3926
rect -29217 3892 -29183 3926
rect -29148 3892 -29114 3926
rect -29078 3896 -29044 3930
rect -29010 3896 -28976 3930
rect -28942 3896 -28908 3930
rect -28874 3896 -28840 3930
rect -28806 3896 -28772 3930
rect -28738 3896 -28704 3930
rect -28670 3896 -28636 3930
rect -28602 3896 -28568 3930
rect -28534 3896 -28500 3930
rect -28466 3896 -28432 3930
rect -28398 3896 -28364 3930
rect -28330 3896 -28296 3930
rect -28262 3896 -28228 3930
rect -28194 3896 -28160 3930
rect -28126 3896 -28092 3930
rect -28058 3896 -28024 3930
rect -27990 3896 -27956 3930
rect -27922 3896 -27888 3930
rect -27854 3896 -27820 3930
rect -27786 3896 -27752 3930
rect -27718 3896 -27684 3930
rect -27650 3896 -27616 3930
rect -27582 3896 -27548 3930
rect -27514 3896 -27480 3930
rect -27446 3896 -27412 3930
rect -27378 3896 -27344 3930
rect -27310 3896 -27276 3930
rect -27242 3896 -27208 3930
rect -27174 3896 -27140 3930
rect -27106 3896 -27072 3930
rect -31632 3822 -31598 3856
rect -31563 3822 -31529 3856
rect -31494 3822 -31460 3856
rect -31425 3822 -31391 3856
rect -31356 3822 -31322 3856
rect -31287 3822 -31253 3856
rect -31218 3822 -31184 3856
rect -31149 3822 -31115 3856
rect -31080 3822 -31046 3856
rect -31011 3822 -30977 3856
rect -30942 3822 -30908 3856
rect -30873 3822 -30839 3856
rect -30804 3822 -30770 3856
rect -30735 3822 -30701 3856
rect -30666 3822 -30632 3856
rect -30597 3822 -30563 3856
rect -30528 3822 -30494 3856
rect -30459 3822 -30425 3856
rect -30390 3822 -30356 3856
rect -30321 3822 -30287 3856
rect -30252 3822 -30218 3856
rect -30183 3822 -30149 3856
rect -30114 3822 -30080 3856
rect -30045 3822 -30011 3856
rect -29976 3822 -29942 3856
rect -29907 3822 -29873 3856
rect -29838 3822 -29804 3856
rect -29769 3822 -29735 3856
rect -29700 3822 -29666 3856
rect -29631 3822 -29597 3856
rect -29562 3822 -29528 3856
rect -29493 3822 -29459 3856
rect -29424 3822 -29390 3856
rect -29355 3822 -29321 3856
rect -29286 3822 -29252 3856
rect -29217 3822 -29183 3856
rect -29148 3822 -29114 3856
rect -29078 3827 -29044 3861
rect -29010 3827 -28976 3861
rect -28942 3827 -28908 3861
rect -28874 3827 -28840 3861
rect -28806 3827 -28772 3861
rect -28738 3827 -28704 3861
rect -28670 3827 -28636 3861
rect -28602 3827 -28568 3861
rect -28534 3827 -28500 3861
rect -28466 3827 -28432 3861
rect -28398 3827 -28364 3861
rect -28330 3827 -28296 3861
rect -28262 3827 -28228 3861
rect -28194 3827 -28160 3861
rect -28126 3827 -28092 3861
rect -28058 3827 -28024 3861
rect -27990 3827 -27956 3861
rect -27922 3827 -27888 3861
rect -27854 3827 -27820 3861
rect -27786 3827 -27752 3861
rect -27718 3827 -27684 3861
rect -27650 3827 -27616 3861
rect -27582 3827 -27548 3861
rect -27514 3827 -27480 3861
rect -27446 3827 -27412 3861
rect -27378 3827 -27344 3861
rect -27310 3827 -27276 3861
rect -27242 3827 -27208 3861
rect -27174 3827 -27140 3861
rect -27106 3827 -27072 3861
rect -31632 3752 -31598 3786
rect -31563 3752 -31529 3786
rect -31494 3752 -31460 3786
rect -31425 3752 -31391 3786
rect -31356 3752 -31322 3786
rect -31287 3752 -31253 3786
rect -31218 3752 -31184 3786
rect -31149 3752 -31115 3786
rect -31080 3752 -31046 3786
rect -31011 3752 -30977 3786
rect -30942 3752 -30908 3786
rect -30873 3752 -30839 3786
rect -30804 3752 -30770 3786
rect -30735 3752 -30701 3786
rect -30666 3752 -30632 3786
rect -30597 3752 -30563 3786
rect -30528 3752 -30494 3786
rect -30459 3752 -30425 3786
rect -30390 3752 -30356 3786
rect -30321 3752 -30287 3786
rect -30252 3752 -30218 3786
rect -30183 3752 -30149 3786
rect -30114 3752 -30080 3786
rect -30045 3752 -30011 3786
rect -29976 3752 -29942 3786
rect -29907 3752 -29873 3786
rect -29838 3752 -29804 3786
rect -29769 3752 -29735 3786
rect -29700 3752 -29666 3786
rect -29631 3752 -29597 3786
rect -29562 3752 -29528 3786
rect -29493 3752 -29459 3786
rect -29424 3752 -29390 3786
rect -29355 3752 -29321 3786
rect -29286 3752 -29252 3786
rect -29217 3752 -29183 3786
rect -29148 3752 -29114 3786
rect -29078 3758 -29044 3792
rect -29010 3758 -28976 3792
rect -28942 3758 -28908 3792
rect -28874 3758 -28840 3792
rect -28806 3758 -28772 3792
rect -28738 3758 -28704 3792
rect -28670 3758 -28636 3792
rect -28602 3758 -28568 3792
rect -28534 3758 -28500 3792
rect -28466 3758 -28432 3792
rect -28398 3758 -28364 3792
rect -28330 3758 -28296 3792
rect -28262 3758 -28228 3792
rect -28194 3758 -28160 3792
rect -28126 3758 -28092 3792
rect -28058 3758 -28024 3792
rect -27990 3758 -27956 3792
rect -27922 3758 -27888 3792
rect -27854 3758 -27820 3792
rect -27786 3758 -27752 3792
rect -27718 3758 -27684 3792
rect -27650 3758 -27616 3792
rect -27582 3758 -27548 3792
rect -27514 3758 -27480 3792
rect -27446 3758 -27412 3792
rect -27378 3758 -27344 3792
rect -27310 3758 -27276 3792
rect -27242 3758 -27208 3792
rect -27174 3758 -27140 3792
rect -27106 3758 -27072 3792
rect -31632 3682 -31598 3716
rect -31563 3682 -31529 3716
rect -31494 3682 -31460 3716
rect -31425 3682 -31391 3716
rect -31356 3682 -31322 3716
rect -31287 3682 -31253 3716
rect -31218 3682 -31184 3716
rect -31149 3682 -31115 3716
rect -31080 3682 -31046 3716
rect -31011 3682 -30977 3716
rect -30942 3682 -30908 3716
rect -30873 3682 -30839 3716
rect -30804 3682 -30770 3716
rect -30735 3682 -30701 3716
rect -30666 3682 -30632 3716
rect -30597 3682 -30563 3716
rect -30528 3682 -30494 3716
rect -30459 3682 -30425 3716
rect -30390 3682 -30356 3716
rect -30321 3682 -30287 3716
rect -30252 3682 -30218 3716
rect -30183 3682 -30149 3716
rect -30114 3682 -30080 3716
rect -30045 3682 -30011 3716
rect -29976 3682 -29942 3716
rect -29907 3682 -29873 3716
rect -29838 3682 -29804 3716
rect -29769 3682 -29735 3716
rect -29700 3682 -29666 3716
rect -29631 3682 -29597 3716
rect -29562 3682 -29528 3716
rect -29493 3682 -29459 3716
rect -29424 3682 -29390 3716
rect -29355 3682 -29321 3716
rect -29286 3682 -29252 3716
rect -29217 3682 -29183 3716
rect -29148 3682 -29114 3716
rect -29078 3689 -29044 3723
rect -29010 3689 -28976 3723
rect -28942 3689 -28908 3723
rect -28874 3689 -28840 3723
rect -28806 3689 -28772 3723
rect -28738 3689 -28704 3723
rect -28670 3689 -28636 3723
rect -28602 3689 -28568 3723
rect -28534 3689 -28500 3723
rect -28466 3689 -28432 3723
rect -28398 3689 -28364 3723
rect -28330 3689 -28296 3723
rect -28262 3689 -28228 3723
rect -28194 3689 -28160 3723
rect -28126 3689 -28092 3723
rect -28058 3689 -28024 3723
rect -27990 3689 -27956 3723
rect -27922 3689 -27888 3723
rect -27854 3689 -27820 3723
rect -27786 3689 -27752 3723
rect -27718 3689 -27684 3723
rect -27650 3689 -27616 3723
rect -27582 3689 -27548 3723
rect -27514 3689 -27480 3723
rect -27446 3689 -27412 3723
rect -27378 3689 -27344 3723
rect -27310 3689 -27276 3723
rect -27242 3689 -27208 3723
rect -27174 3689 -27140 3723
rect -27106 3689 -27072 3723
rect -31632 3612 -31598 3646
rect -31563 3612 -31529 3646
rect -31494 3612 -31460 3646
rect -31425 3612 -31391 3646
rect -31356 3612 -31322 3646
rect -31287 3612 -31253 3646
rect -31218 3612 -31184 3646
rect -31149 3612 -31115 3646
rect -31080 3612 -31046 3646
rect -31011 3612 -30977 3646
rect -30942 3612 -30908 3646
rect -30873 3612 -30839 3646
rect -30804 3612 -30770 3646
rect -30735 3612 -30701 3646
rect -30666 3612 -30632 3646
rect -30597 3612 -30563 3646
rect -30528 3612 -30494 3646
rect -30459 3612 -30425 3646
rect -30390 3612 -30356 3646
rect -30321 3612 -30287 3646
rect -30252 3612 -30218 3646
rect -30183 3612 -30149 3646
rect -30114 3612 -30080 3646
rect -30045 3612 -30011 3646
rect -29976 3612 -29942 3646
rect -29907 3612 -29873 3646
rect -29838 3612 -29804 3646
rect -29769 3612 -29735 3646
rect -29700 3612 -29666 3646
rect -29631 3612 -29597 3646
rect -29562 3612 -29528 3646
rect -29493 3612 -29459 3646
rect -29424 3612 -29390 3646
rect -29355 3612 -29321 3646
rect -29286 3612 -29252 3646
rect -29217 3612 -29183 3646
rect -29148 3612 -29114 3646
rect -29078 3620 -29044 3654
rect -29010 3620 -28976 3654
rect -28942 3620 -28908 3654
rect -28874 3620 -28840 3654
rect -28806 3620 -28772 3654
rect -28738 3620 -28704 3654
rect -28670 3620 -28636 3654
rect -28602 3620 -28568 3654
rect -28534 3620 -28500 3654
rect -28466 3620 -28432 3654
rect -28398 3620 -28364 3654
rect -28330 3620 -28296 3654
rect -28262 3620 -28228 3654
rect -28194 3620 -28160 3654
rect -28126 3620 -28092 3654
rect -28058 3620 -28024 3654
rect -27990 3620 -27956 3654
rect -27922 3620 -27888 3654
rect -27854 3620 -27820 3654
rect -27786 3620 -27752 3654
rect -27718 3620 -27684 3654
rect -27650 3620 -27616 3654
rect -27582 3620 -27548 3654
rect -27514 3620 -27480 3654
rect -27446 3620 -27412 3654
rect -27378 3620 -27344 3654
rect -27310 3620 -27276 3654
rect -27242 3620 -27208 3654
rect -27174 3620 -27140 3654
rect -27106 3620 -27072 3654
rect -31632 3542 -31598 3576
rect -31563 3542 -31529 3576
rect -31494 3542 -31460 3576
rect -31425 3542 -31391 3576
rect -31356 3542 -31322 3576
rect -31287 3542 -31253 3576
rect -31218 3542 -31184 3576
rect -31149 3542 -31115 3576
rect -31080 3542 -31046 3576
rect -31011 3542 -30977 3576
rect -30942 3542 -30908 3576
rect -30873 3542 -30839 3576
rect -30804 3542 -30770 3576
rect -30735 3542 -30701 3576
rect -30666 3542 -30632 3576
rect -30597 3542 -30563 3576
rect -30528 3542 -30494 3576
rect -30459 3542 -30425 3576
rect -30390 3542 -30356 3576
rect -30321 3542 -30287 3576
rect -30252 3542 -30218 3576
rect -30183 3542 -30149 3576
rect -30114 3542 -30080 3576
rect -30045 3542 -30011 3576
rect -29976 3542 -29942 3576
rect -29907 3542 -29873 3576
rect -29838 3542 -29804 3576
rect -29769 3542 -29735 3576
rect -29700 3542 -29666 3576
rect -29631 3542 -29597 3576
rect -29562 3542 -29528 3576
rect -29493 3542 -29459 3576
rect -29424 3542 -29390 3576
rect -29355 3542 -29321 3576
rect -29286 3542 -29252 3576
rect -29217 3542 -29183 3576
rect -29148 3542 -29114 3576
rect -29078 3551 -29044 3585
rect -29010 3551 -28976 3585
rect -28942 3551 -28908 3585
rect -28874 3551 -28840 3585
rect -28806 3551 -28772 3585
rect -28738 3551 -28704 3585
rect -28670 3551 -28636 3585
rect -28602 3551 -28568 3585
rect -28534 3551 -28500 3585
rect -28466 3551 -28432 3585
rect -28398 3551 -28364 3585
rect -28330 3551 -28296 3585
rect -28262 3551 -28228 3585
rect -28194 3551 -28160 3585
rect -28126 3551 -28092 3585
rect -28058 3551 -28024 3585
rect -27990 3551 -27956 3585
rect -27922 3551 -27888 3585
rect -27854 3551 -27820 3585
rect -27786 3551 -27752 3585
rect -27718 3551 -27684 3585
rect -27650 3551 -27616 3585
rect -27582 3551 -27548 3585
rect -27514 3551 -27480 3585
rect -27446 3551 -27412 3585
rect -27378 3551 -27344 3585
rect -27310 3551 -27276 3585
rect -27242 3551 -27208 3585
rect -27174 3551 -27140 3585
rect -27106 3551 -27072 3585
rect -31632 3472 -31598 3506
rect -31563 3472 -31529 3506
rect -31494 3472 -31460 3506
rect -31425 3472 -31391 3506
rect -31356 3472 -31322 3506
rect -31287 3472 -31253 3506
rect -31218 3472 -31184 3506
rect -31149 3472 -31115 3506
rect -31080 3472 -31046 3506
rect -31011 3472 -30977 3506
rect -30942 3472 -30908 3506
rect -30873 3472 -30839 3506
rect -30804 3472 -30770 3506
rect -30735 3472 -30701 3506
rect -30666 3472 -30632 3506
rect -30597 3472 -30563 3506
rect -30528 3472 -30494 3506
rect -30459 3472 -30425 3506
rect -30390 3472 -30356 3506
rect -30321 3472 -30287 3506
rect -30252 3472 -30218 3506
rect -30183 3472 -30149 3506
rect -30114 3472 -30080 3506
rect -30045 3472 -30011 3506
rect -29976 3472 -29942 3506
rect -29907 3472 -29873 3506
rect -29838 3472 -29804 3506
rect -29769 3472 -29735 3506
rect -29700 3472 -29666 3506
rect -29631 3472 -29597 3506
rect -29562 3472 -29528 3506
rect -29493 3472 -29459 3506
rect -29424 3472 -29390 3506
rect -29355 3472 -29321 3506
rect -29286 3472 -29252 3506
rect -29217 3472 -29183 3506
rect -29148 3472 -29114 3506
rect -29078 3482 -29044 3516
rect -29010 3482 -28976 3516
rect -28942 3482 -28908 3516
rect -28874 3482 -28840 3516
rect -28806 3482 -28772 3516
rect -28738 3482 -28704 3516
rect -28670 3482 -28636 3516
rect -28602 3482 -28568 3516
rect -28534 3482 -28500 3516
rect -28466 3482 -28432 3516
rect -28398 3482 -28364 3516
rect -28330 3482 -28296 3516
rect -28262 3482 -28228 3516
rect -28194 3482 -28160 3516
rect -28126 3482 -28092 3516
rect -28058 3482 -28024 3516
rect -27990 3482 -27956 3516
rect -27922 3482 -27888 3516
rect -27854 3482 -27820 3516
rect -27786 3482 -27752 3516
rect -27718 3482 -27684 3516
rect -27650 3482 -27616 3516
rect -27582 3482 -27548 3516
rect -27514 3482 -27480 3516
rect -27446 3482 -27412 3516
rect -27378 3482 -27344 3516
rect -27310 3482 -27276 3516
rect -27242 3482 -27208 3516
rect -27174 3482 -27140 3516
rect -27106 3482 -27072 3516
rect -31632 3402 -31598 3436
rect -31563 3402 -31529 3436
rect -31494 3402 -31460 3436
rect -31425 3402 -31391 3436
rect -31356 3402 -31322 3436
rect -31287 3402 -31253 3436
rect -31218 3402 -31184 3436
rect -31149 3402 -31115 3436
rect -31080 3402 -31046 3436
rect -31011 3402 -30977 3436
rect -30942 3402 -30908 3436
rect -30873 3402 -30839 3436
rect -30804 3402 -30770 3436
rect -30735 3402 -30701 3436
rect -30666 3402 -30632 3436
rect -30597 3402 -30563 3436
rect -30528 3402 -30494 3436
rect -30459 3402 -30425 3436
rect -30390 3402 -30356 3436
rect -30321 3402 -30287 3436
rect -30252 3402 -30218 3436
rect -30183 3402 -30149 3436
rect -30114 3402 -30080 3436
rect -30045 3402 -30011 3436
rect -29976 3402 -29942 3436
rect -29907 3402 -29873 3436
rect -29838 3402 -29804 3436
rect -29769 3402 -29735 3436
rect -29700 3402 -29666 3436
rect -29631 3402 -29597 3436
rect -29562 3402 -29528 3436
rect -29493 3402 -29459 3436
rect -29424 3402 -29390 3436
rect -29355 3402 -29321 3436
rect -29286 3402 -29252 3436
rect -29217 3402 -29183 3436
rect -29148 3402 -29114 3436
rect -29078 3413 -29044 3447
rect -29010 3413 -28976 3447
rect -28942 3413 -28908 3447
rect -28874 3413 -28840 3447
rect -28806 3413 -28772 3447
rect -28738 3413 -28704 3447
rect -28670 3413 -28636 3447
rect -28602 3413 -28568 3447
rect -28534 3413 -28500 3447
rect -28466 3413 -28432 3447
rect -28398 3413 -28364 3447
rect -28330 3413 -28296 3447
rect -28262 3413 -28228 3447
rect -28194 3413 -28160 3447
rect -28126 3413 -28092 3447
rect -28058 3413 -28024 3447
rect -27990 3413 -27956 3447
rect -27922 3413 -27888 3447
rect -27854 3413 -27820 3447
rect -27786 3413 -27752 3447
rect -27718 3413 -27684 3447
rect -27650 3413 -27616 3447
rect -27582 3413 -27548 3447
rect -27514 3413 -27480 3447
rect -27446 3413 -27412 3447
rect -27378 3413 -27344 3447
rect -27310 3413 -27276 3447
rect -27242 3413 -27208 3447
rect -27174 3413 -27140 3447
rect -27106 3413 -27072 3447
rect -29078 3344 -29044 3378
rect -29010 3344 -28976 3378
rect -28942 3344 -28908 3378
rect -28874 3344 -28840 3378
rect -28806 3344 -28772 3378
rect -28738 3344 -28704 3378
rect -28670 3344 -28636 3378
rect -28602 3344 -28568 3378
rect -28534 3344 -28500 3378
rect -28466 3344 -28432 3378
rect -28398 3344 -28364 3378
rect -28330 3344 -28296 3378
rect -28262 3344 -28228 3378
rect -28194 3344 -28160 3378
rect -28126 3344 -28092 3378
rect -28058 3344 -28024 3378
rect -27990 3344 -27956 3378
rect -27922 3344 -27888 3378
rect -27854 3344 -27820 3378
rect -27786 3344 -27752 3378
rect -27718 3344 -27684 3378
rect -27650 3344 -27616 3378
rect -27582 3344 -27548 3378
rect -27514 3344 -27480 3378
rect -27446 3344 -27412 3378
rect -27378 3344 -27344 3378
rect -27310 3344 -27276 3378
rect -27242 3344 -27208 3378
rect -27174 3344 -27140 3378
rect -27106 3344 -27072 3378
rect -31564 3300 -31530 3334
rect -31496 3300 -31462 3334
rect -31428 3300 -31394 3334
rect -31360 3300 -31326 3334
rect -31292 3300 -31258 3334
rect -31224 3300 -31190 3334
rect -31156 3300 -31122 3334
rect -31088 3300 -31054 3334
rect -31020 3300 -30986 3334
rect -30952 3300 -30918 3334
rect -30884 3300 -30850 3334
rect -30816 3300 -30782 3334
rect -30748 3300 -30714 3334
rect -30680 3300 -30646 3334
rect -30612 3300 -30578 3334
rect -30544 3300 -30510 3334
rect -30476 3300 -30442 3334
rect -30408 3300 -30374 3334
rect -30340 3300 -30306 3334
rect -30272 3300 -30238 3334
rect -30204 3300 -30170 3334
rect -30136 3300 -30102 3334
rect -30068 3300 -30034 3334
rect -30000 3300 -29966 3334
rect -29932 3300 -29898 3334
rect -29864 3300 -29830 3334
rect -29796 3300 -29762 3334
rect -29728 3300 -29694 3334
rect -29660 3300 -29626 3334
rect -29592 3300 -29558 3334
rect -29524 3300 -29490 3334
rect -29456 3300 -29422 3334
rect -29388 3300 -29354 3334
rect -29260 3300 -29226 3334
rect -31632 3189 -31598 3223
rect -29078 3275 -29044 3309
rect -29010 3275 -28976 3309
rect -28942 3275 -28908 3309
rect -28874 3275 -28840 3309
rect -28806 3275 -28772 3309
rect -28738 3275 -28704 3309
rect -28670 3275 -28636 3309
rect -28602 3275 -28568 3309
rect -28534 3275 -28500 3309
rect -28466 3275 -28432 3309
rect -28398 3275 -28364 3309
rect -28330 3275 -28296 3309
rect -28262 3275 -28228 3309
rect -28194 3275 -28160 3309
rect -28126 3275 -28092 3309
rect -28058 3275 -28024 3309
rect -27990 3275 -27956 3309
rect -27922 3275 -27888 3309
rect -27854 3275 -27820 3309
rect -27786 3275 -27752 3309
rect -27718 3275 -27684 3309
rect -27650 3275 -27616 3309
rect -27582 3275 -27548 3309
rect -27514 3275 -27480 3309
rect -27446 3275 -27412 3309
rect -27378 3275 -27344 3309
rect -27310 3275 -27276 3309
rect -27242 3275 -27208 3309
rect -27174 3275 -27140 3309
rect -27106 3275 -27072 3309
rect -29148 3232 -29114 3266
rect -31632 3121 -31598 3155
rect -31632 3053 -31598 3087
rect -31632 2985 -31598 3019
rect -31632 2917 -31598 2951
rect -31632 2849 -31598 2883
rect -31632 2781 -31598 2815
rect -31632 2713 -31598 2747
rect -31632 2645 -31598 2679
rect -31632 2577 -31598 2611
rect -31632 2509 -31598 2543
rect -31632 2441 -31598 2475
rect -31632 2373 -31598 2407
rect -31632 2305 -31598 2339
rect -31632 2237 -31598 2271
rect -31632 2169 -31598 2203
rect -31632 2101 -31598 2135
rect -31632 2033 -31598 2067
rect -31632 1965 -31598 1999
rect -31632 1897 -31598 1931
rect -31632 1829 -31598 1863
rect -31632 1761 -31598 1795
rect -31632 1693 -31598 1727
rect -31632 1625 -31598 1659
rect -31632 1557 -31598 1591
rect -31632 1489 -31598 1523
rect -31632 1421 -31598 1455
rect -31632 1353 -31598 1387
rect -31632 1285 -31598 1319
rect -31632 1217 -31598 1251
rect -31632 1149 -31598 1183
rect -31632 1081 -31598 1115
rect -31632 1013 -31598 1047
rect -31632 945 -31598 979
rect -31632 877 -31598 911
rect -31632 809 -31598 843
rect -31632 741 -31598 775
rect -31632 673 -31598 707
rect -31632 605 -31598 639
rect -31632 537 -31598 571
rect -31632 469 -31598 503
rect -31632 401 -31598 435
rect -31632 333 -31598 367
rect -31632 265 -31598 299
rect -31632 197 -31598 231
rect -31632 129 -31598 163
rect -31632 61 -31598 95
rect -31632 -7 -31598 27
rect -31632 -75 -31598 -41
rect -31632 -143 -31598 -109
rect -31632 -211 -31598 -177
rect -31632 -279 -31598 -245
rect -31632 -347 -31598 -313
rect -31632 -415 -31598 -381
rect -31632 -483 -31598 -449
rect -31632 -551 -31598 -517
rect -31632 -619 -31598 -585
rect -31632 -687 -31598 -653
rect -31632 -755 -31598 -721
rect -31632 -823 -31598 -789
rect -31632 -891 -31598 -857
rect -31632 -959 -31598 -925
rect -31632 -1027 -31598 -993
rect -31632 -1095 -31598 -1061
rect -31632 -1163 -31598 -1129
rect -31632 -1231 -31598 -1197
rect -31632 -1299 -31598 -1265
rect -31632 -1367 -31598 -1333
rect -31632 -1435 -31598 -1401
rect -31632 -1503 -31598 -1469
rect -31632 -1571 -31598 -1537
rect -31632 -1639 -31598 -1605
rect -31632 -1707 -31598 -1673
rect -31632 -1775 -31598 -1741
rect -31632 -1843 -31598 -1809
rect -31632 -1911 -31598 -1877
rect -31632 -1979 -31598 -1945
rect -31632 -2047 -31598 -2013
rect -31632 -2115 -31598 -2081
rect -31632 -2183 -31598 -2149
rect -31632 -2251 -31598 -2217
rect -31632 -2319 -31598 -2285
rect -31632 -2387 -31598 -2353
rect -31632 -2455 -31598 -2421
rect -31632 -2523 -31598 -2489
rect -31632 -2591 -31598 -2557
rect -31632 -2659 -31598 -2625
rect -31632 -2727 -31598 -2693
rect -31632 -2795 -31598 -2761
rect -31632 -2863 -31598 -2829
rect -31632 -2931 -31598 -2897
rect -31632 -2999 -31598 -2965
rect -31632 -3067 -31598 -3033
rect -31632 -3135 -31598 -3101
rect -31632 -3203 -31598 -3169
rect -31632 -3271 -31598 -3237
rect -31632 -3339 -31598 -3305
rect -31632 -3407 -31598 -3373
rect -31632 -3475 -31598 -3441
rect -31632 -3543 -31598 -3509
rect -31632 -3611 -31598 -3577
rect -31632 -3679 -31598 -3645
rect -31632 -3747 -31598 -3713
rect -31632 -3815 -31598 -3781
rect -31632 -3883 -31598 -3849
rect -31632 -3951 -31598 -3917
rect -31632 -4019 -31598 -3985
rect -31632 -4087 -31598 -4053
rect -31632 -4155 -31598 -4121
rect -31632 -4223 -31598 -4189
rect -31632 -4291 -31598 -4257
rect -31632 -4359 -31598 -4325
rect -31632 -4427 -31598 -4393
rect -31632 -4495 -31598 -4461
rect -31632 -4563 -31598 -4529
rect -31632 -4631 -31598 -4597
rect -31632 -4699 -31598 -4665
rect -31632 -4767 -31598 -4733
rect -31632 -4835 -31598 -4801
rect -31632 -4903 -31598 -4869
rect -31632 -4971 -31598 -4937
rect -31632 -5039 -31598 -5005
rect -31632 -5107 -31598 -5073
rect -31632 -5175 -31598 -5141
rect -31632 -5243 -31598 -5209
rect -31632 -5311 -31598 -5277
rect -31632 -5379 -31598 -5345
rect -31632 -5447 -31598 -5413
rect -31632 -5515 -31598 -5481
rect -31632 -5583 -31598 -5549
rect -31632 -5651 -31598 -5617
rect -31632 -5719 -31598 -5685
rect -31632 -5787 -31598 -5753
rect -31632 -5855 -31598 -5821
rect -31632 -5923 -31598 -5889
rect -31632 -5991 -31598 -5957
rect -31632 -6059 -31598 -6025
rect -31632 -6127 -31598 -6093
rect -31632 -6195 -31598 -6161
rect -31632 -6263 -31598 -6229
rect -31632 -6331 -31598 -6297
rect -31632 -6399 -31598 -6365
rect -31632 -6467 -31598 -6433
rect -31632 -6535 -31598 -6501
rect -31632 -6603 -31598 -6569
rect -31632 -6671 -31598 -6637
rect -31632 -6739 -31598 -6705
rect -31632 -6807 -31598 -6773
rect -31632 -6875 -31598 -6841
rect -31632 -6943 -31598 -6909
rect -31632 -7011 -31598 -6977
rect -31632 -7079 -31598 -7045
rect -31632 -7147 -31598 -7113
rect -31632 -7215 -31598 -7181
rect -31632 -7283 -31598 -7249
rect -31632 -7351 -31598 -7317
rect -31632 -7419 -31598 -7385
rect -31632 -7487 -31598 -7453
rect -31632 -7555 -31598 -7521
rect -31632 -7623 -31598 -7589
rect -31632 -7691 -31598 -7657
rect -31632 -7759 -31598 -7725
rect -31632 -7827 -31598 -7793
rect -31632 -7895 -31598 -7861
rect -31632 -7963 -31598 -7929
rect -31632 -8031 -31598 -7997
rect -31632 -8099 -31598 -8065
rect -31632 -8167 -31598 -8133
rect -31632 -8235 -31598 -8201
rect -31632 -8303 -31598 -8269
rect -31632 -8371 -31598 -8337
rect -31632 -8439 -31598 -8405
rect -31632 -8507 -31598 -8473
rect -31632 -8575 -31598 -8541
rect -31632 -8643 -31598 -8609
rect -31632 -8711 -31598 -8677
rect -29078 3206 -29044 3240
rect -29010 3206 -28976 3240
rect -28942 3206 -28908 3240
rect -28874 3206 -28840 3240
rect -28806 3206 -28772 3240
rect -28738 3206 -28704 3240
rect -28670 3206 -28636 3240
rect -28602 3206 -28568 3240
rect -28534 3206 -28500 3240
rect -28466 3206 -28432 3240
rect -28398 3206 -28364 3240
rect -28330 3206 -28296 3240
rect -28262 3206 -28228 3240
rect -28194 3206 -28160 3240
rect -28126 3206 -28092 3240
rect -28058 3206 -28024 3240
rect -27990 3206 -27956 3240
rect -27922 3206 -27888 3240
rect -27854 3206 -27820 3240
rect -27786 3206 -27752 3240
rect -27718 3206 -27684 3240
rect -27650 3206 -27616 3240
rect -27582 3206 -27548 3240
rect -27514 3206 -27480 3240
rect -27446 3206 -27412 3240
rect -27378 3206 -27344 3240
rect -27310 3206 -27276 3240
rect -27242 3206 -27208 3240
rect -27174 3206 -27140 3240
rect -27106 3206 -27072 3240
rect -29148 3164 -29114 3198
rect -29078 3137 -29044 3171
rect -29010 3137 -28976 3171
rect -28942 3137 -28908 3171
rect -28874 3137 -28840 3171
rect -28806 3137 -28772 3171
rect -28738 3137 -28704 3171
rect -28670 3137 -28636 3171
rect -28602 3137 -28568 3171
rect -28534 3137 -28500 3171
rect -28466 3137 -28432 3171
rect -28398 3137 -28364 3171
rect -28330 3137 -28296 3171
rect -28262 3137 -28228 3171
rect -28194 3137 -28160 3171
rect -28126 3137 -28092 3171
rect -28058 3137 -28024 3171
rect -27990 3137 -27956 3171
rect -27922 3137 -27888 3171
rect -27854 3137 -27820 3171
rect -27786 3137 -27752 3171
rect -27718 3137 -27684 3171
rect -27650 3137 -27616 3171
rect -27582 3137 -27548 3171
rect -27514 3137 -27480 3171
rect -27446 3137 -27412 3171
rect -27378 3137 -27344 3171
rect -27310 3137 -27276 3171
rect -27242 3137 -27208 3171
rect -27174 3137 -27140 3171
rect -27106 3137 -27072 3171
rect -29148 3096 -29114 3130
rect -29078 3068 -29044 3102
rect -29010 3068 -28976 3102
rect -28942 3068 -28908 3102
rect -28874 3068 -28840 3102
rect -28806 3068 -28772 3102
rect -28738 3068 -28704 3102
rect -28670 3068 -28636 3102
rect -28602 3068 -28568 3102
rect -28534 3068 -28500 3102
rect -28466 3068 -28432 3102
rect -28398 3068 -28364 3102
rect -28330 3068 -28296 3102
rect -28262 3068 -28228 3102
rect -28194 3068 -28160 3102
rect -28126 3068 -28092 3102
rect -28058 3068 -28024 3102
rect -27990 3068 -27956 3102
rect -27922 3068 -27888 3102
rect -27854 3068 -27820 3102
rect -27786 3068 -27752 3102
rect -27718 3068 -27684 3102
rect -27650 3068 -27616 3102
rect -27582 3068 -27548 3102
rect -27514 3068 -27480 3102
rect -27446 3068 -27412 3102
rect -27378 3068 -27344 3102
rect -27310 3068 -27276 3102
rect -27242 3068 -27208 3102
rect -27174 3068 -27140 3102
rect -27106 3068 -27072 3102
rect -29148 3028 -29114 3062
rect -29078 2999 -29044 3033
rect -29010 2999 -28976 3033
rect -28942 2999 -28908 3033
rect -28874 2999 -28840 3033
rect -28806 2999 -28772 3033
rect -28738 2999 -28704 3033
rect -28670 2999 -28636 3033
rect -28602 2999 -28568 3033
rect -28534 2999 -28500 3033
rect -28466 2999 -28432 3033
rect -28398 2999 -28364 3033
rect -28330 2999 -28296 3033
rect -28262 2999 -28228 3033
rect -28194 2999 -28160 3033
rect -28126 2999 -28092 3033
rect -28058 2999 -28024 3033
rect -27990 2999 -27956 3033
rect -27922 2999 -27888 3033
rect -27854 2999 -27820 3033
rect -27786 2999 -27752 3033
rect -27718 2999 -27684 3033
rect -27650 2999 -27616 3033
rect -27582 2999 -27548 3033
rect -27514 2999 -27480 3033
rect -27446 2999 -27412 3033
rect -27378 2999 -27344 3033
rect -27310 2999 -27276 3033
rect -27242 2999 -27208 3033
rect -27174 2999 -27140 3033
rect -27106 2999 -27072 3033
rect -29148 2960 -29114 2994
rect -29078 2930 -29044 2964
rect -29010 2930 -28976 2964
rect -28942 2930 -28908 2964
rect -28874 2930 -28840 2964
rect -28806 2930 -28772 2964
rect -28738 2930 -28704 2964
rect -28670 2930 -28636 2964
rect -28602 2930 -28568 2964
rect -28534 2930 -28500 2964
rect -28466 2930 -28432 2964
rect -28398 2930 -28364 2964
rect -28330 2930 -28296 2964
rect -28262 2930 -28228 2964
rect -28194 2930 -28160 2964
rect -28126 2930 -28092 2964
rect -28058 2930 -28024 2964
rect -27990 2930 -27956 2964
rect -27922 2930 -27888 2964
rect -27854 2930 -27820 2964
rect -27786 2930 -27752 2964
rect -27718 2930 -27684 2964
rect -27650 2930 -27616 2964
rect -27582 2930 -27548 2964
rect -27514 2930 -27480 2964
rect -27446 2930 -27412 2964
rect -27378 2930 -27344 2964
rect -27310 2930 -27276 2964
rect -27242 2930 -27208 2964
rect -27174 2930 -27140 2964
rect -27106 2930 -27072 2964
rect -29148 2892 -29114 2926
rect -29078 2861 -29044 2895
rect -29010 2861 -28976 2895
rect -28942 2861 -28908 2895
rect -28874 2861 -28840 2895
rect -28806 2861 -28772 2895
rect -28738 2861 -28704 2895
rect -28670 2861 -28636 2895
rect -28602 2861 -28568 2895
rect -28534 2861 -28500 2895
rect -28466 2861 -28432 2895
rect -28398 2861 -28364 2895
rect -28330 2861 -28296 2895
rect -28262 2861 -28228 2895
rect -28194 2861 -28160 2895
rect -28126 2861 -28092 2895
rect -28058 2861 -28024 2895
rect -27990 2861 -27956 2895
rect -27922 2861 -27888 2895
rect -27854 2861 -27820 2895
rect -27786 2861 -27752 2895
rect -27718 2861 -27684 2895
rect -27650 2861 -27616 2895
rect -27582 2861 -27548 2895
rect -27514 2861 -27480 2895
rect -27446 2861 -27412 2895
rect -27378 2861 -27344 2895
rect -27310 2861 -27276 2895
rect -27242 2861 -27208 2895
rect -27174 2861 -27140 2895
rect -27106 2861 -27072 2895
rect -29148 2824 -29114 2858
rect -29078 2792 -29044 2826
rect -29010 2792 -28976 2826
rect -28942 2792 -28908 2826
rect -28874 2792 -28840 2826
rect -28806 2792 -28772 2826
rect -28738 2792 -28704 2826
rect -28670 2792 -28636 2826
rect -28602 2792 -28568 2826
rect -28534 2792 -28500 2826
rect -28466 2792 -28432 2826
rect -28398 2792 -28364 2826
rect -28330 2792 -28296 2826
rect -28262 2792 -28228 2826
rect -28194 2792 -28160 2826
rect -28126 2792 -28092 2826
rect -28058 2792 -28024 2826
rect -27990 2792 -27956 2826
rect -27922 2792 -27888 2826
rect -27854 2792 -27820 2826
rect -27786 2792 -27752 2826
rect -27718 2792 -27684 2826
rect -27650 2792 -27616 2826
rect -27582 2792 -27548 2826
rect -27514 2792 -27480 2826
rect -27446 2792 -27412 2826
rect -27378 2792 -27344 2826
rect -27310 2792 -27276 2826
rect -27242 2792 -27208 2826
rect -27174 2792 -27140 2826
rect -27106 2792 -27072 2826
rect -29148 2756 -29114 2790
rect -29078 2723 -29044 2757
rect -29010 2723 -28976 2757
rect -28942 2723 -28908 2757
rect -28874 2723 -28840 2757
rect -28806 2723 -28772 2757
rect -28738 2723 -28704 2757
rect -28670 2723 -28636 2757
rect -28602 2723 -28568 2757
rect -28534 2723 -28500 2757
rect -28466 2723 -28432 2757
rect -28398 2723 -28364 2757
rect -28330 2723 -28296 2757
rect -28262 2723 -28228 2757
rect -28194 2723 -28160 2757
rect -28126 2723 -28092 2757
rect -28058 2723 -28024 2757
rect -27990 2723 -27956 2757
rect -27922 2723 -27888 2757
rect -27854 2723 -27820 2757
rect -27786 2723 -27752 2757
rect -27718 2723 -27684 2757
rect -27650 2723 -27616 2757
rect -27582 2723 -27548 2757
rect -27514 2723 -27480 2757
rect -27446 2723 -27412 2757
rect -27378 2723 -27344 2757
rect -27310 2723 -27276 2757
rect -27242 2723 -27208 2757
rect -27174 2723 -27140 2757
rect -27106 2723 -27072 2757
rect -29148 2688 -29114 2722
rect -29078 2654 -29044 2688
rect -29010 2654 -28976 2688
rect -28942 2654 -28908 2688
rect -28874 2654 -28840 2688
rect -28806 2654 -28772 2688
rect -28738 2654 -28704 2688
rect -28670 2654 -28636 2688
rect -28602 2654 -28568 2688
rect -28534 2654 -28500 2688
rect -28466 2654 -28432 2688
rect -28398 2654 -28364 2688
rect -28330 2654 -28296 2688
rect -28262 2654 -28228 2688
rect -28194 2654 -28160 2688
rect -28126 2654 -28092 2688
rect -28058 2654 -28024 2688
rect -27990 2654 -27956 2688
rect -27922 2654 -27888 2688
rect -27854 2654 -27820 2688
rect -27786 2654 -27752 2688
rect -27718 2654 -27684 2688
rect -27650 2654 -27616 2688
rect -27582 2654 -27548 2688
rect -27514 2654 -27480 2688
rect -27446 2654 -27412 2688
rect -27378 2654 -27344 2688
rect -27310 2654 -27276 2688
rect -27242 2654 -27208 2688
rect -27174 2654 -27140 2688
rect -27106 2654 -27072 2688
rect -29148 2620 -29114 2654
rect -29148 2552 -29114 2586
rect -29078 2585 -29044 2619
rect -29010 2585 -28976 2619
rect -28942 2585 -28908 2619
rect -28874 2585 -28840 2619
rect -28806 2585 -28772 2619
rect -28738 2585 -28704 2619
rect -28670 2585 -28636 2619
rect -28602 2585 -28568 2619
rect -28534 2585 -28500 2619
rect -28466 2585 -28432 2619
rect -28398 2585 -28364 2619
rect -28330 2585 -28296 2619
rect -28262 2585 -28228 2619
rect -28194 2585 -28160 2619
rect -28126 2585 -28092 2619
rect -28058 2585 -28024 2619
rect -27990 2585 -27956 2619
rect -27922 2585 -27888 2619
rect -27854 2585 -27820 2619
rect -27786 2585 -27752 2619
rect -27718 2585 -27684 2619
rect -27650 2585 -27616 2619
rect -27582 2585 -27548 2619
rect -27514 2585 -27480 2619
rect -27446 2585 -27412 2619
rect -27378 2585 -27344 2619
rect -27310 2585 -27276 2619
rect -27242 2585 -27208 2619
rect -27174 2585 -27140 2619
rect -27106 2585 -27072 2619
rect -29148 2484 -29114 2518
rect -29078 2516 -29044 2550
rect -29010 2516 -28976 2550
rect -28942 2516 -28908 2550
rect -28874 2516 -28840 2550
rect -28806 2516 -28772 2550
rect -28738 2516 -28704 2550
rect -28670 2516 -28636 2550
rect -28602 2516 -28568 2550
rect -28534 2516 -28500 2550
rect -28466 2516 -28432 2550
rect -28398 2516 -28364 2550
rect -28330 2516 -28296 2550
rect -28262 2516 -28228 2550
rect -28194 2516 -28160 2550
rect -28126 2516 -28092 2550
rect -28058 2516 -28024 2550
rect -27990 2516 -27956 2550
rect -27922 2516 -27888 2550
rect -27854 2516 -27820 2550
rect -27786 2516 -27752 2550
rect -27718 2516 -27684 2550
rect -27650 2516 -27616 2550
rect -27582 2516 -27548 2550
rect -27514 2516 -27480 2550
rect -27446 2516 -27412 2550
rect -27378 2516 -27344 2550
rect -27310 2516 -27276 2550
rect -27242 2516 -27208 2550
rect -27174 2516 -27140 2550
rect -27106 2516 -27072 2550
rect -29148 2416 -29114 2450
rect -29078 2447 -29044 2481
rect -29010 2447 -28976 2481
rect -28942 2447 -28908 2481
rect -28874 2447 -28840 2481
rect -28806 2447 -28772 2481
rect -28738 2447 -28704 2481
rect -28670 2447 -28636 2481
rect -28602 2447 -28568 2481
rect -28534 2447 -28500 2481
rect -28466 2447 -28432 2481
rect -28398 2447 -28364 2481
rect -28330 2447 -28296 2481
rect -28262 2447 -28228 2481
rect -28194 2447 -28160 2481
rect -28126 2447 -28092 2481
rect -28058 2447 -28024 2481
rect -27990 2447 -27956 2481
rect -27922 2447 -27888 2481
rect -27854 2447 -27820 2481
rect -27786 2447 -27752 2481
rect -27718 2447 -27684 2481
rect -27650 2447 -27616 2481
rect -27582 2447 -27548 2481
rect -27514 2447 -27480 2481
rect -27446 2447 -27412 2481
rect -27378 2447 -27344 2481
rect -27310 2447 -27276 2481
rect -27242 2447 -27208 2481
rect -27174 2447 -27140 2481
rect -27106 2447 -27072 2481
rect -29148 2348 -29114 2382
rect -29078 2378 -29044 2412
rect -29010 2378 -28976 2412
rect -28942 2378 -28908 2412
rect -28874 2378 -28840 2412
rect -28806 2378 -28772 2412
rect -28738 2378 -28704 2412
rect -28670 2378 -28636 2412
rect -28602 2378 -28568 2412
rect -28534 2378 -28500 2412
rect -28466 2378 -28432 2412
rect -28398 2378 -28364 2412
rect -28330 2378 -28296 2412
rect -28262 2378 -28228 2412
rect -28194 2378 -28160 2412
rect -28126 2378 -28092 2412
rect -28058 2378 -28024 2412
rect -27990 2378 -27956 2412
rect -27922 2378 -27888 2412
rect -27854 2378 -27820 2412
rect -27786 2378 -27752 2412
rect -27718 2378 -27684 2412
rect -27650 2378 -27616 2412
rect -27582 2378 -27548 2412
rect -27514 2378 -27480 2412
rect -27446 2378 -27412 2412
rect -27378 2378 -27344 2412
rect -27310 2378 -27276 2412
rect -27242 2378 -27208 2412
rect -27174 2378 -27140 2412
rect -27106 2378 -27072 2412
rect -29148 2280 -29114 2314
rect -29078 2309 -29044 2343
rect -29010 2309 -28976 2343
rect -28942 2309 -28908 2343
rect -28874 2309 -28840 2343
rect -28806 2309 -28772 2343
rect -28738 2309 -28704 2343
rect -28670 2309 -28636 2343
rect -28602 2309 -28568 2343
rect -28534 2309 -28500 2343
rect -28466 2309 -28432 2343
rect -28398 2309 -28364 2343
rect -28330 2309 -28296 2343
rect -28262 2309 -28228 2343
rect -28194 2309 -28160 2343
rect -28126 2309 -28092 2343
rect -28058 2309 -28024 2343
rect -27990 2309 -27956 2343
rect -27922 2309 -27888 2343
rect -27854 2309 -27820 2343
rect -27786 2309 -27752 2343
rect -27718 2309 -27684 2343
rect -27650 2309 -27616 2343
rect -27582 2309 -27548 2343
rect -27514 2309 -27480 2343
rect -27446 2309 -27412 2343
rect -27378 2309 -27344 2343
rect -27310 2309 -27276 2343
rect -27242 2309 -27208 2343
rect -27174 2309 -27140 2343
rect -27106 2309 -27072 2343
rect -29148 2212 -29114 2246
rect -29078 2240 -29044 2274
rect -29010 2240 -28976 2274
rect -28942 2240 -28908 2274
rect -28874 2240 -28840 2274
rect -28806 2240 -28772 2274
rect -28738 2240 -28704 2274
rect -28670 2240 -28636 2274
rect -28602 2240 -28568 2274
rect -28534 2240 -28500 2274
rect -28466 2240 -28432 2274
rect -28398 2240 -28364 2274
rect -28330 2240 -28296 2274
rect -28262 2240 -28228 2274
rect -28194 2240 -28160 2274
rect -28126 2240 -28092 2274
rect -28058 2240 -28024 2274
rect -27990 2240 -27956 2274
rect -27922 2240 -27888 2274
rect -27854 2240 -27820 2274
rect -27786 2240 -27752 2274
rect -27718 2240 -27684 2274
rect -27650 2240 -27616 2274
rect -27582 2240 -27548 2274
rect -27514 2240 -27480 2274
rect -27446 2240 -27412 2274
rect -27378 2240 -27344 2274
rect -27310 2240 -27276 2274
rect -27242 2240 -27208 2274
rect -27174 2240 -27140 2274
rect -27106 2240 -27072 2274
rect -29148 2144 -29114 2178
rect -29078 2171 -29044 2205
rect -29010 2171 -28976 2205
rect -28942 2171 -28908 2205
rect -28874 2171 -28840 2205
rect -28806 2171 -28772 2205
rect -28738 2171 -28704 2205
rect -28670 2171 -28636 2205
rect -28602 2171 -28568 2205
rect -28534 2171 -28500 2205
rect -28466 2171 -28432 2205
rect -28398 2171 -28364 2205
rect -28330 2171 -28296 2205
rect -28262 2171 -28228 2205
rect -28194 2171 -28160 2205
rect -28126 2171 -28092 2205
rect -28058 2171 -28024 2205
rect -27990 2171 -27956 2205
rect -27922 2171 -27888 2205
rect -27854 2171 -27820 2205
rect -27786 2171 -27752 2205
rect -27718 2171 -27684 2205
rect -27650 2171 -27616 2205
rect -27582 2171 -27548 2205
rect -27514 2171 -27480 2205
rect -27446 2171 -27412 2205
rect -27378 2171 -27344 2205
rect -27310 2171 -27276 2205
rect -27242 2171 -27208 2205
rect -27174 2171 -27140 2205
rect -27106 2171 -27072 2205
rect -29148 2076 -29114 2110
rect -29078 2102 -29044 2136
rect -29010 2102 -28976 2136
rect -28942 2102 -28908 2136
rect -28874 2102 -28840 2136
rect -28806 2102 -28772 2136
rect -28738 2102 -28704 2136
rect -28670 2102 -28636 2136
rect -28602 2102 -28568 2136
rect -28534 2102 -28500 2136
rect -28466 2102 -28432 2136
rect -28398 2102 -28364 2136
rect -28330 2102 -28296 2136
rect -28262 2102 -28228 2136
rect -28194 2102 -28160 2136
rect -28126 2102 -28092 2136
rect -28058 2102 -28024 2136
rect -27990 2102 -27956 2136
rect -27922 2102 -27888 2136
rect -27854 2102 -27820 2136
rect -27786 2102 -27752 2136
rect -27718 2102 -27684 2136
rect -27650 2102 -27616 2136
rect -27582 2102 -27548 2136
rect -27514 2102 -27480 2136
rect -27446 2102 -27412 2136
rect -27378 2102 -27344 2136
rect -27310 2102 -27276 2136
rect -27242 2102 -27208 2136
rect -27174 2102 -27140 2136
rect -27106 2102 -27072 2136
rect -29148 2008 -29114 2042
rect -29148 1940 -29114 1974
rect -29148 1872 -29114 1906
rect -29148 1804 -29114 1838
rect -29148 1736 -29114 1770
rect -29148 1668 -29114 1702
rect -29148 1600 -29114 1634
rect -29148 1532 -29114 1566
rect -29148 1464 -29114 1498
rect -29148 1396 -29114 1430
rect -29148 1328 -29114 1362
rect -29148 1260 -29114 1294
rect -29148 1192 -29114 1226
rect -29148 1124 -29114 1158
rect -29148 1056 -29114 1090
rect -29148 988 -29114 1022
rect -29148 920 -29114 954
rect -29148 852 -29114 886
rect -29148 784 -29114 818
rect -29148 716 -29114 750
rect -29148 648 -29114 682
rect -29148 580 -29114 614
rect -29148 512 -29114 546
rect -29148 444 -29114 478
rect -29148 376 -29114 410
rect -29148 308 -29114 342
rect -29148 240 -29114 274
rect -29148 172 -29114 206
rect -29148 104 -29114 138
rect -29148 36 -29114 70
rect -29148 -32 -29114 2
rect -29148 -100 -29114 -66
rect -29148 -168 -29114 -134
rect -29148 -236 -29114 -202
rect -29148 -304 -29114 -270
rect -29148 -372 -29114 -338
rect -29148 -440 -29114 -406
rect -29148 -508 -29114 -474
rect -29148 -576 -29114 -542
rect -29148 -644 -29114 -610
rect -29148 -712 -29114 -678
rect -29148 -780 -29114 -746
rect -29148 -848 -29114 -814
rect -29148 -916 -29114 -882
rect -29148 -984 -29114 -950
rect -29148 -1052 -29114 -1018
rect -29148 -1120 -29114 -1086
rect -29148 -1188 -29114 -1154
rect -29148 -1256 -29114 -1222
rect -29148 -1324 -29114 -1290
rect -29148 -1392 -29114 -1358
rect -29148 -1460 -29114 -1426
rect -29148 -1528 -29114 -1494
rect -29148 -1596 -29114 -1562
rect -29148 -1664 -29114 -1630
rect -29148 -1732 -29114 -1698
rect -29148 -1800 -29114 -1766
rect -29148 -1868 -29114 -1834
rect -29148 -1936 -29114 -1902
rect -29148 -2004 -29114 -1970
rect -29148 -2072 -29114 -2038
rect -29148 -2140 -29114 -2106
rect -29148 -2208 -29114 -2174
rect -29148 -2276 -29114 -2242
rect -29148 -2344 -29114 -2310
rect -29148 -2412 -29114 -2378
rect -29148 -2480 -29114 -2446
rect -29148 -2548 -29114 -2514
rect -29148 -2616 -29114 -2582
rect -29148 -2684 -29114 -2650
rect -29148 -2752 -29114 -2718
rect -29148 -2820 -29114 -2786
rect -29148 -2888 -29114 -2854
rect -29148 -2956 -29114 -2922
rect -29148 -3024 -29114 -2990
rect -29148 -3092 -29114 -3058
rect -29148 -3160 -29114 -3126
rect -29148 -3228 -29114 -3194
rect -29148 -3296 -29114 -3262
rect -29148 -3364 -29114 -3330
rect -29148 -3432 -29114 -3398
rect -29148 -3500 -29114 -3466
rect -29148 -3568 -29114 -3534
rect -29148 -3636 -29114 -3602
rect -29148 -3704 -29114 -3670
rect -29148 -3772 -29114 -3738
rect -29148 -3840 -29114 -3806
rect -29148 -3908 -29114 -3874
rect -29148 -3976 -29114 -3942
rect -29148 -4044 -29114 -4010
rect -29148 -4112 -29114 -4078
rect -29148 -4180 -29114 -4146
rect -29148 -4248 -29114 -4214
rect -29148 -4316 -29114 -4282
rect -29148 -4384 -29114 -4350
rect -29148 -4452 -29114 -4418
rect -29148 -4520 -29114 -4486
rect -29148 -4588 -29114 -4554
rect -29148 -4656 -29114 -4622
rect -29148 -4724 -29114 -4690
rect -29148 -4792 -29114 -4758
rect -29148 -4860 -29114 -4826
rect -29148 -4928 -29114 -4894
rect -29148 -4996 -29114 -4962
rect -29148 -5064 -29114 -5030
rect -29148 -5132 -29114 -5098
rect -29148 -5200 -29114 -5166
rect -29148 -5268 -29114 -5234
rect -29148 -5336 -29114 -5302
rect -29148 -5404 -29114 -5370
rect -29148 -5472 -29114 -5438
rect -29148 -5540 -29114 -5506
rect -29148 -5608 -29114 -5574
rect -29148 -5676 -29114 -5642
rect -29148 -5744 -29114 -5710
rect -29148 -5812 -29114 -5778
rect -29148 -5880 -29114 -5846
rect -29148 -5948 -29114 -5914
rect -29148 -6016 -29114 -5982
rect -29148 -6084 -29114 -6050
rect -29148 -6152 -29114 -6118
rect -29148 -6220 -29114 -6186
rect -29148 -6288 -29114 -6254
rect -29148 -6356 -29114 -6322
rect -29148 -6424 -29114 -6390
rect -29148 -6492 -29114 -6458
rect -29148 -6560 -29114 -6526
rect -29148 -6628 -29114 -6594
rect -29148 -6696 -29114 -6662
rect -29148 -6764 -29114 -6730
rect -29148 -6832 -29114 -6798
rect -29148 -6900 -29114 -6866
rect -29148 -6968 -29114 -6934
rect -29148 -7036 -29114 -7002
rect -29148 -7104 -29114 -7070
rect -29148 -7172 -29114 -7138
rect -29148 -7240 -29114 -7206
rect -29148 -7308 -29114 -7274
rect -29148 -7376 -29114 -7342
rect -29148 -7444 -29114 -7410
rect -29148 -7512 -29114 -7478
rect -29148 -7580 -29114 -7546
rect -29148 -7648 -29114 -7614
rect -29148 -7716 -29114 -7682
rect -29148 -7784 -29114 -7750
rect -29148 -7852 -29114 -7818
rect -29148 -7920 -29114 -7886
rect -29148 -7988 -29114 -7954
rect -29148 -8056 -29114 -8022
rect -29148 -8124 -29114 -8090
rect -29148 -8192 -29114 -8158
rect -29148 -8260 -29114 -8226
rect -29148 -8328 -29114 -8294
rect -29148 -8396 -29114 -8362
rect -29148 -8464 -29114 -8430
rect -29148 -8532 -29114 -8498
rect -29148 -8600 -29114 -8566
rect -29148 -8668 -29114 -8634
rect -29148 -8736 -29114 -8702
rect -31632 -8779 -31598 -8745
rect -31528 -8847 -31494 -8813
rect -31460 -8847 -31426 -8813
rect -31392 -8847 -31358 -8813
rect -31324 -8847 -31290 -8813
rect -31256 -8847 -31222 -8813
rect -31188 -8847 -31154 -8813
rect -31120 -8847 -31086 -8813
rect -31052 -8847 -31018 -8813
rect -30984 -8847 -30950 -8813
rect -30916 -8847 -30882 -8813
rect -30848 -8847 -30814 -8813
rect -30780 -8847 -30746 -8813
rect -30712 -8847 -30678 -8813
rect -30644 -8847 -30610 -8813
rect -30576 -8847 -30542 -8813
rect -30508 -8847 -30474 -8813
rect -30440 -8847 -30406 -8813
rect -30372 -8847 -30338 -8813
rect -30304 -8847 -30270 -8813
rect -30236 -8847 -30202 -8813
rect -30168 -8847 -30134 -8813
rect -30100 -8847 -30066 -8813
rect -30032 -8847 -29998 -8813
rect -29964 -8847 -29930 -8813
rect -29896 -8847 -29862 -8813
rect -29828 -8847 -29794 -8813
rect -29760 -8847 -29726 -8813
rect -29692 -8847 -29658 -8813
rect -29624 -8847 -29590 -8813
rect -29556 -8847 -29522 -8813
rect -29488 -8847 -29454 -8813
rect -29420 -8847 -29386 -8813
rect -29352 -8847 -29318 -8813
rect -29284 -8847 -29250 -8813
rect -29216 -8847 -29182 -8813
rect -29078 -8847 -27072 2067
rect 5738 3398 5772 3432
rect 5738 3330 5772 3364
rect 5738 3262 5772 3296
rect 5738 3194 5772 3228
rect 5738 3126 5772 3160
rect 5738 3058 5772 3092
rect 5738 2990 5772 3024
rect 5738 2922 5772 2956
rect 5738 2854 5772 2888
rect 5738 2786 5772 2820
rect 5738 2718 5772 2752
rect 5738 2650 5772 2684
rect 5738 2582 5772 2616
rect 5738 2514 5772 2548
rect -31632 -9598 -27450 -8884
rect -27415 -8918 -27381 -8884
rect -27346 -8918 -27312 -8884
rect -27277 -8918 -27243 -8884
rect -27208 -8918 -27174 -8884
rect -27139 -8918 -27105 -8884
rect -27070 -8918 -27036 -8884
rect -27415 -8986 -27381 -8952
rect -27346 -8986 -27312 -8952
rect -27277 -8986 -27243 -8952
rect -27208 -8986 -27174 -8952
rect -27139 -8986 -27105 -8952
rect -27070 -8986 -27036 -8952
rect -27415 -9054 -27381 -9020
rect -27346 -9054 -27312 -9020
rect -27277 -9054 -27243 -9020
rect -27208 -9054 -27174 -9020
rect -27139 -9054 -27105 -9020
rect -27070 -9054 -27036 -9020
rect -27415 -9122 -27381 -9088
rect -27346 -9122 -27312 -9088
rect -27277 -9122 -27243 -9088
rect -27208 -9122 -27174 -9088
rect -27139 -9122 -27105 -9088
rect -27070 -9122 -27036 -9088
rect -27415 -9190 -27381 -9156
rect -27346 -9190 -27312 -9156
rect -27277 -9190 -27243 -9156
rect -27208 -9190 -27174 -9156
rect -27139 -9190 -27105 -9156
rect -27070 -9190 -27036 -9156
rect -27415 -9258 -27381 -9224
rect -27346 -9258 -27312 -9224
rect -27277 -9258 -27243 -9224
rect -27208 -9258 -27174 -9224
rect -27139 -9258 -27105 -9224
rect -27070 -9258 -27036 -9224
rect -27415 -9326 -27381 -9292
rect -27346 -9326 -27312 -9292
rect -27277 -9326 -27243 -9292
rect -27208 -9326 -27174 -9292
rect -27139 -9326 -27105 -9292
rect -27070 -9326 -27036 -9292
rect -27415 -9394 -27381 -9360
rect -27346 -9394 -27312 -9360
rect -27277 -9394 -27243 -9360
rect -27208 -9394 -27174 -9360
rect -27139 -9394 -27105 -9360
rect -27070 -9394 -27036 -9360
rect -27415 -9462 -27381 -9428
rect -27346 -9462 -27312 -9428
rect -27277 -9462 -27243 -9428
rect -27208 -9462 -27174 -9428
rect -27139 -9462 -27105 -9428
rect -27070 -9462 -27036 -9428
rect -27415 -9530 -27381 -9496
rect -27346 -9530 -27312 -9496
rect -27277 -9530 -27243 -9496
rect -27208 -9530 -27174 -9496
rect -27139 -9530 -27105 -9496
rect -27070 -9530 -27036 -9496
rect -27415 -9598 -27381 -9564
rect -27346 -9598 -27312 -9564
rect -27277 -9598 -27243 -9564
rect -27208 -9598 -27174 -9564
rect -27139 -9598 -27105 -9564
rect -27070 -9598 -27036 -9564
<< mvnsubdiffcont >>
rect -733 3654 -699 3688
rect -662 3654 -628 3688
rect -591 3654 -557 3688
rect -519 3654 -485 3688
rect -447 3654 -413 3688
rect 181 3654 215 3688
rect 250 3654 284 3688
rect 319 3654 353 3688
rect 388 3654 422 3688
rect 457 3654 491 3688
rect 526 3654 560 3688
rect 595 3654 629 3688
rect 664 3654 698 3688
rect 733 3654 767 3688
rect 802 3654 836 3688
rect 871 3654 905 3688
rect 940 3654 974 3688
rect 1009 3654 1043 3688
rect 1078 3654 1112 3688
rect 1147 3654 1181 3688
rect 1216 3654 1250 3688
rect 1285 3654 1319 3688
rect 1354 3654 1388 3688
rect 1423 3654 1457 3688
rect 1492 3654 1526 3688
rect 1561 3654 1595 3688
rect 1630 3654 1664 3688
rect 1699 3654 1733 3688
rect 1768 3654 1802 3688
rect 1837 3654 1871 3688
rect 1906 3654 1940 3688
rect 1975 3654 2009 3688
rect 2044 3654 2078 3688
rect 2113 3654 2147 3688
rect 2182 3654 2216 3688
rect 2251 3654 2285 3688
rect 2320 3654 2354 3688
rect 2389 3654 2423 3688
rect 2458 3654 2492 3688
rect 2527 3654 2561 3688
rect 2596 3654 2630 3688
rect 2665 3654 2699 3688
rect 2734 3654 2768 3688
rect 2803 3654 2837 3688
rect 2872 3654 2906 3688
rect 2941 3654 2975 3688
rect 3010 3654 3044 3688
rect 3078 3654 3112 3688
rect 3146 3654 3180 3688
rect 3214 3654 3248 3688
rect 3282 3654 3316 3688
rect 3350 3654 3384 3688
rect 3418 3654 3452 3688
rect 3486 3654 3520 3688
rect 6732 3267 6766 3301
rect 6732 3193 6766 3227
rect 6732 3119 6766 3153
rect 6732 3045 6766 3079
rect 6732 2971 6766 3005
rect 6732 2897 6766 2931
rect 6732 2824 6766 2858
rect 6732 2751 6766 2785
rect 6732 2678 6766 2712
rect 6732 2605 6766 2639
<< poly >>
rect -9813 4312 -9733 4328
rect -9813 4278 -9790 4312
rect -9756 4278 -9733 4312
rect -11573 -8693 -11550 -8659
rect -11516 -8693 -11493 -8659
rect -11573 -8727 -11493 -8693
rect -9813 4244 -9733 4278
rect -9813 4210 -9790 4244
rect -9756 4210 -9733 4244
rect -701 3580 -601 3612
rect -545 3580 -445 3612
rect 213 3580 313 3612
rect 369 3580 469 3612
rect 661 3580 761 3612
rect 817 3580 917 3612
rect 1100 3580 1200 3612
rect 1460 3580 1560 3612
rect 1753 3545 1853 3577
rect 1909 3545 2009 3577
rect 2065 3545 2165 3577
rect 2802 3545 2902 3577
rect 3085 3545 3185 3577
rect 3241 3545 3341 3577
rect 3397 3545 3497 3577
rect -701 2548 -601 2580
rect -545 2548 -445 2580
rect -701 2532 -445 2548
rect -701 2498 -685 2532
rect -651 2498 -590 2532
rect -556 2498 -495 2532
rect -461 2498 -445 2532
rect -701 2482 -445 2498
rect 213 2524 313 2580
rect 213 2490 248 2524
rect 282 2490 313 2524
rect 213 2456 313 2490
rect 213 2422 248 2456
rect 282 2422 313 2456
rect 213 2406 313 2422
rect 369 2524 469 2580
rect 369 2490 404 2524
rect 438 2490 469 2524
rect 369 2456 469 2490
rect 369 2422 404 2456
rect 438 2422 469 2456
rect 369 2406 469 2422
rect 661 2524 761 2580
rect 661 2490 696 2524
rect 730 2490 761 2524
rect 661 2456 761 2490
rect 661 2422 696 2456
rect 730 2422 761 2456
rect 661 2406 761 2422
rect 817 2524 917 2580
rect 817 2490 852 2524
rect 886 2490 917 2524
rect 817 2456 917 2490
rect 817 2422 852 2456
rect 886 2422 917 2456
rect 817 2406 917 2422
rect 1100 2524 1200 2580
rect 1100 2490 1135 2524
rect 1169 2490 1200 2524
rect 1100 2456 1200 2490
rect 1100 2422 1135 2456
rect 1169 2422 1200 2456
rect 1100 2406 1200 2422
rect 1460 2524 1560 2580
rect 2356 3482 2456 3514
rect 2512 3482 2612 3514
rect 2356 3233 2456 3398
rect 2356 3199 2394 3233
rect 2428 3199 2456 3233
rect 2356 3165 2456 3199
rect 2356 3131 2394 3165
rect 2428 3131 2456 3165
rect 2356 3115 2456 3131
rect 2512 3233 2612 3398
rect 2512 3199 2550 3233
rect 2584 3199 2612 3233
rect 2512 3165 2612 3199
rect 2512 3131 2550 3165
rect 2584 3131 2612 3165
rect 2512 3115 2612 3131
rect 2802 2884 2902 2945
rect 2802 2850 2822 2884
rect 2856 2850 2902 2884
rect 2802 2816 2902 2850
rect 3085 2913 3185 2945
rect 3241 2913 3341 2945
rect 3397 2913 3497 2945
rect 3085 2897 3497 2913
rect 3085 2863 3101 2897
rect 3135 2863 3171 2897
rect 3205 2863 3240 2897
rect 3274 2863 3309 2897
rect 3343 2863 3378 2897
rect 3412 2863 3447 2897
rect 3481 2863 3497 2897
rect 3085 2847 3497 2863
rect 2802 2782 2822 2816
rect 2856 2782 2902 2816
rect 2802 2752 2902 2782
rect 1460 2490 1495 2524
rect 1529 2490 1560 2524
rect 1460 2456 1560 2490
rect 1460 2422 1495 2456
rect 1529 2422 1560 2456
rect 1460 2406 1560 2422
rect 1753 2489 1853 2545
rect 1753 2455 1788 2489
rect 1822 2455 1853 2489
rect 1753 2421 1853 2455
rect 1753 2387 1788 2421
rect 1822 2387 1853 2421
rect 1753 2371 1853 2387
rect 1909 2489 2009 2545
rect 1909 2455 1944 2489
rect 1978 2455 2009 2489
rect 1909 2421 2009 2455
rect 1909 2387 1944 2421
rect 1978 2387 2009 2421
rect 1909 2371 2009 2387
rect 2065 2489 2165 2545
rect 2065 2455 2100 2489
rect 2134 2455 2165 2489
rect 2065 2421 2165 2455
rect 2065 2387 2100 2421
rect 2134 2387 2165 2421
rect 2065 2371 2165 2387
rect 289 2237 469 2269
rect 4289 3545 4389 3577
rect 4289 2489 4389 2545
rect 4289 2455 4324 2489
rect 4358 2455 4389 2489
rect 4289 2421 4389 2455
rect 4289 2387 4324 2421
rect 4358 2387 4389 2421
rect 4289 2371 4389 2387
rect 5261 3488 5421 3520
rect 5261 3216 5421 3288
rect 5261 3182 5326 3216
rect 5360 3182 5421 3216
rect 5261 3148 5421 3182
rect 5261 3114 5326 3148
rect 5360 3114 5421 3148
rect 5261 3078 5421 3114
rect 5261 2982 5421 3014
rect 5261 2710 5421 2782
rect 5261 2676 5326 2710
rect 5360 2676 5421 2710
rect 5261 2642 5421 2676
rect 5261 2608 5326 2642
rect 5360 2608 5421 2642
rect 5261 2572 5421 2608
rect 5826 3152 5852 3272
rect 5992 3226 6190 3272
rect 5992 3192 6040 3226
rect 6074 3192 6108 3226
rect 6142 3192 6190 3226
rect 5992 3152 6190 3192
rect 6390 3152 6458 3272
rect 6658 3152 6684 3272
rect 5826 2976 5852 3096
rect 5992 3055 6190 3096
rect 5992 3021 6040 3055
rect 6074 3021 6108 3055
rect 6142 3021 6190 3055
rect 5992 2976 6190 3021
rect 6390 2976 6458 3096
rect 6658 2976 6684 3096
rect 5826 2675 5852 2795
rect 5992 2751 6190 2795
rect 5992 2717 6040 2751
rect 6074 2717 6108 2751
rect 6142 2717 6190 2751
rect 5992 2675 6190 2717
rect 6390 2675 6458 2795
rect 6658 2675 6684 2795
rect 2176 2049 2276 2069
rect 3491 2065 3591 2081
rect 289 2005 469 2037
rect 2176 2015 2206 2049
rect 2240 2015 2276 2049
rect -176 1983 -16 1999
rect -176 1949 -160 1983
rect -126 1949 -66 1983
rect -32 1949 -16 1983
rect -176 1901 -16 1949
rect 171 1986 979 2005
rect 171 1952 187 1986
rect 221 1952 262 1986
rect 296 1952 337 1986
rect 371 1952 411 1986
rect 445 1952 485 1986
rect 519 1952 559 1986
rect 593 1952 633 1986
rect 667 1952 707 1986
rect 741 1952 781 1986
rect 815 1952 855 1986
rect 889 1952 929 1986
rect 963 1952 979 1986
rect 171 1933 979 1952
rect 171 1901 331 1933
rect 387 1901 547 1933
rect 603 1901 763 1933
rect 819 1901 979 1933
rect 1035 1983 1843 1999
rect 1035 1949 1051 1983
rect 1085 1949 1125 1983
rect 1159 1949 1199 1983
rect 1233 1949 1273 1983
rect 1307 1949 1347 1983
rect 1381 1949 1421 1983
rect 1455 1949 1495 1983
rect 1529 1949 1569 1983
rect 1603 1949 1643 1983
rect 1677 1949 1718 1983
rect 1752 1949 1793 1983
rect 1827 1949 1843 1983
rect 1035 1933 1843 1949
rect 1035 1901 1195 1933
rect 1251 1901 1411 1933
rect 1467 1901 1627 1933
rect 1683 1901 1843 1933
rect 2176 1981 2276 2015
rect 2176 1947 2206 1981
rect 2240 1947 2276 1981
rect 2176 1886 2276 1947
rect 2459 2049 2559 2065
rect 2459 2015 2489 2049
rect 2523 2015 2559 2049
rect 2459 1981 2559 2015
rect 3491 2031 3530 2065
rect 3564 2031 3591 2065
rect 2459 1947 2489 1981
rect 2523 1947 2559 1981
rect 2459 1886 2559 1947
rect 2742 1989 2998 2005
rect 2742 1955 2758 1989
rect 2792 1955 2853 1989
rect 2887 1955 2948 1989
rect 2982 1955 2998 1989
rect 2742 1939 2998 1955
rect 2742 1907 2842 1939
rect 2898 1907 2998 1939
rect 3054 1989 3310 2005
rect 3054 1955 3070 1989
rect 3104 1955 3165 1989
rect 3199 1955 3260 1989
rect 3294 1955 3310 1989
rect 3054 1939 3310 1955
rect 3054 1907 3154 1939
rect 3210 1907 3310 1939
rect 3491 1997 3591 2031
rect 3491 1963 3530 1997
rect 3564 1963 3591 1997
rect 2176 1254 2276 1286
rect 2459 1254 2559 1286
rect 3491 1901 3591 1963
rect 3934 1956 4114 1972
rect 3934 1922 3950 1956
rect 3984 1922 4064 1956
rect 4098 1922 4114 1956
rect 3934 1859 4114 1922
rect 3934 1627 4114 1659
rect 3491 1269 3591 1301
rect -176 869 -16 901
rect 171 869 331 901
rect 387 869 547 901
rect 603 869 763 901
rect 819 869 979 901
rect 1035 869 1195 901
rect 1251 869 1411 901
rect 1467 869 1627 901
rect 1683 869 1843 901
rect 2742 875 2842 907
rect 2898 875 2998 907
rect 3054 875 3154 907
rect 3210 875 3310 907
rect 2742 679 2842 711
rect 2898 679 2998 711
rect 3054 679 3154 711
rect 111 449 143 629
rect 2143 628 2175 629
rect 2143 612 2241 628
rect 2143 578 2191 612
rect 2225 578 2241 612
rect 2143 498 2241 578
rect 2143 464 2191 498
rect 2225 464 2241 498
rect 2143 449 2241 464
rect 2175 448 2241 449
rect 2742 447 2842 479
rect 2898 447 2998 479
rect 3054 447 3154 479
rect 2742 431 3154 447
rect 2742 397 2758 431
rect 2792 397 2828 431
rect 2862 397 2897 431
rect 2931 397 2966 431
rect 3000 397 3035 431
rect 3069 397 3104 431
rect 3138 397 3154 431
rect 2742 381 3154 397
rect 111 86 143 266
rect 2143 250 2241 266
rect 2143 216 2191 250
rect 2225 216 2241 250
rect 2143 136 2241 216
rect 2143 102 2191 136
rect 2225 102 2241 136
rect 2143 86 2241 102
rect -11573 -8761 -11550 -8727
rect -11516 -8761 -11493 -8727
rect -11573 -8777 -11493 -8761
<< polycont >>
rect -9790 4278 -9756 4312
rect -11550 -8693 -11516 -8659
rect -9790 4210 -9756 4244
rect -685 2498 -651 2532
rect -590 2498 -556 2532
rect -495 2498 -461 2532
rect 248 2490 282 2524
rect 248 2422 282 2456
rect 404 2490 438 2524
rect 404 2422 438 2456
rect 696 2490 730 2524
rect 696 2422 730 2456
rect 852 2490 886 2524
rect 852 2422 886 2456
rect 1135 2490 1169 2524
rect 1135 2422 1169 2456
rect 2394 3199 2428 3233
rect 2394 3131 2428 3165
rect 2550 3199 2584 3233
rect 2550 3131 2584 3165
rect 2822 2850 2856 2884
rect 3101 2863 3135 2897
rect 3171 2863 3205 2897
rect 3240 2863 3274 2897
rect 3309 2863 3343 2897
rect 3378 2863 3412 2897
rect 3447 2863 3481 2897
rect 2822 2782 2856 2816
rect 1495 2490 1529 2524
rect 1495 2422 1529 2456
rect 1788 2455 1822 2489
rect 1788 2387 1822 2421
rect 1944 2455 1978 2489
rect 1944 2387 1978 2421
rect 2100 2455 2134 2489
rect 2100 2387 2134 2421
rect 4324 2455 4358 2489
rect 4324 2387 4358 2421
rect 5326 3182 5360 3216
rect 5326 3114 5360 3148
rect 5326 2676 5360 2710
rect 5326 2608 5360 2642
rect 6040 3192 6074 3226
rect 6108 3192 6142 3226
rect 6040 3021 6074 3055
rect 6108 3021 6142 3055
rect 6040 2717 6074 2751
rect 6108 2717 6142 2751
rect 2206 2015 2240 2049
rect -160 1949 -126 1983
rect -66 1949 -32 1983
rect 187 1952 221 1986
rect 262 1952 296 1986
rect 337 1952 371 1986
rect 411 1952 445 1986
rect 485 1952 519 1986
rect 559 1952 593 1986
rect 633 1952 667 1986
rect 707 1952 741 1986
rect 781 1952 815 1986
rect 855 1952 889 1986
rect 929 1952 963 1986
rect 1051 1949 1085 1983
rect 1125 1949 1159 1983
rect 1199 1949 1233 1983
rect 1273 1949 1307 1983
rect 1347 1949 1381 1983
rect 1421 1949 1455 1983
rect 1495 1949 1529 1983
rect 1569 1949 1603 1983
rect 1643 1949 1677 1983
rect 1718 1949 1752 1983
rect 1793 1949 1827 1983
rect 2206 1947 2240 1981
rect 2489 2015 2523 2049
rect 3530 2031 3564 2065
rect 2489 1947 2523 1981
rect 2758 1955 2792 1989
rect 2853 1955 2887 1989
rect 2948 1955 2982 1989
rect 3070 1955 3104 1989
rect 3165 1955 3199 1989
rect 3260 1955 3294 1989
rect 3530 1963 3564 1997
rect 3950 1922 3984 1956
rect 4064 1922 4098 1956
rect 2191 578 2225 612
rect 2191 464 2225 498
rect 2758 397 2792 431
rect 2828 397 2862 431
rect 2897 397 2931 431
rect 2966 397 3000 431
rect 3035 397 3069 431
rect 3104 397 3138 431
rect 2191 216 2225 250
rect 2191 102 2225 136
rect -11550 -8761 -11516 -8727
<< npolyres >>
rect -11573 4180 -11317 4260
rect -11573 -8659 -11493 4180
rect -11397 -8631 -11317 4180
rect -11221 4180 -10965 4260
rect -11221 -8631 -11141 4180
rect -11397 -8711 -11141 -8631
rect -11045 -8631 -10965 4180
rect -10869 4180 -10613 4260
rect -10869 -8631 -10789 4180
rect -11045 -8711 -10789 -8631
rect -10693 -8631 -10613 4180
rect -10517 4180 -10261 4260
rect -10517 -8631 -10437 4180
rect -10693 -8711 -10437 -8631
rect -10341 -8631 -10261 4180
rect -10165 4180 -9909 4260
rect -10165 -8631 -10085 4180
rect -10341 -8711 -10085 -8631
rect -9989 -8631 -9909 4180
rect -9813 -8631 -9733 4210
rect -9989 -8711 -9733 -8631
<< mvndiffres >>
rect -31524 3162 -31334 3220
rect -31524 -8685 -31466 3162
rect -31392 -8681 -31334 3162
rect -31260 3162 -31070 3220
rect -31260 -8681 -31202 3162
rect -31392 -8739 -31202 -8681
rect -31128 -8681 -31070 3162
rect -30996 3162 -30806 3220
rect -30996 -8681 -30938 3162
rect -31128 -8739 -30938 -8681
rect -30864 -8681 -30806 3162
rect -30732 3162 -30542 3220
rect -30732 -8681 -30674 3162
rect -30864 -8739 -30674 -8681
rect -30600 -8681 -30542 3162
rect -30468 3162 -30278 3220
rect -30468 -8681 -30410 3162
rect -30600 -8739 -30410 -8681
rect -30336 -8681 -30278 3162
rect -30204 3162 -30014 3220
rect -30204 -8681 -30146 3162
rect -30336 -8739 -30146 -8681
rect -30072 -8681 -30014 3162
rect -29940 3162 -29750 3220
rect -29940 -8681 -29882 3162
rect -30072 -8739 -29882 -8681
rect -29808 -8681 -29750 3162
rect -29676 3162 -29486 3220
rect -29676 -8681 -29618 3162
rect -29808 -8739 -29618 -8681
rect -29544 -8681 -29486 3162
rect -29412 3162 -29222 3220
rect -29412 -8681 -29354 3162
rect -29544 -8739 -29354 -8681
rect -29280 -8697 -29222 3162
<< locali >>
rect -32352 4332 -32315 4344
rect -32281 4332 -32247 4344
rect -32213 4332 -32179 4344
rect -32352 4298 -32344 4332
rect -32281 4310 -32266 4332
rect -32213 4310 -32188 4332
rect -32145 4310 -32111 4344
rect -32077 4332 -32043 4344
rect -32009 4332 -31975 4344
rect -31941 4332 -31907 4344
rect -31873 4332 -31839 4344
rect -32076 4310 -32043 4332
rect -31998 4310 -31975 4332
rect -31920 4310 -31907 4332
rect -31842 4310 -31839 4332
rect -31805 4332 -31771 4344
rect -31737 4333 -31703 4344
rect -31669 4333 -29078 4344
rect -29044 4333 -29010 4344
rect -31805 4310 -31798 4332
rect -31737 4310 -31718 4333
rect -31669 4310 -31645 4333
rect -32310 4298 -32266 4310
rect -32232 4298 -32188 4310
rect -32154 4298 -32110 4310
rect -32076 4298 -32032 4310
rect -31998 4298 -31954 4310
rect -31920 4298 -31876 4310
rect -31842 4298 -31798 4310
rect -31764 4299 -31718 4310
rect -31684 4299 -31645 4310
rect -31611 4299 -31572 4333
rect -31538 4299 -31499 4333
rect -31465 4299 -31426 4333
rect -31392 4299 -31353 4333
rect -31319 4299 -31280 4333
rect -31246 4299 -31207 4333
rect -31173 4299 -31134 4333
rect -31100 4299 -31061 4333
rect -31027 4299 -30988 4333
rect -30954 4299 -30915 4333
rect -30881 4299 -30842 4333
rect -30808 4299 -30768 4333
rect -30734 4299 -30694 4333
rect -30660 4299 -30620 4333
rect -30586 4299 -30546 4333
rect -30512 4299 -30472 4333
rect -30438 4299 -30398 4333
rect -30364 4299 -30324 4333
rect -30290 4299 -30250 4333
rect -30216 4299 -30176 4333
rect -30142 4299 -30102 4333
rect -30068 4299 -30028 4333
rect -29994 4299 -29954 4333
rect -29920 4299 -29880 4333
rect -29846 4299 -29806 4333
rect -29772 4299 -29732 4333
rect -29698 4299 -29658 4333
rect -29624 4299 -29584 4333
rect -29550 4299 -29510 4333
rect -29476 4299 -29436 4333
rect -29402 4299 -29362 4333
rect -29328 4299 -29288 4333
rect -29254 4299 -29214 4333
rect -29180 4299 -29134 4333
rect -29100 4310 -29078 4333
rect -29012 4310 -29010 4333
rect -28976 4333 -28942 4344
rect -28976 4310 -28958 4333
rect -28908 4310 -28874 4344
rect -28840 4333 -28806 4344
rect -28836 4310 -28806 4333
rect -28772 4310 -28738 4344
rect -28704 4310 -28670 4344
rect -28636 4310 -28602 4344
rect -28568 4310 -28534 4344
rect -28500 4310 -28466 4344
rect -28432 4310 -28398 4344
rect -28364 4310 -28330 4344
rect -28296 4310 -28262 4344
rect -28228 4310 -28194 4344
rect -28160 4310 -28126 4344
rect -28092 4310 -28058 4344
rect -28024 4310 -27990 4344
rect -27956 4310 -27922 4344
rect -27888 4310 -27854 4344
rect -27820 4310 -27786 4344
rect -27752 4310 -27718 4344
rect -27684 4310 -27650 4344
rect -27616 4310 -27582 4344
rect -27548 4310 -27514 4344
rect -27480 4310 -27446 4344
rect -27412 4310 -27378 4344
rect -27344 4310 -27310 4344
rect -27276 4310 -27242 4344
rect -27208 4310 -27174 4344
rect -27140 4310 -27106 4344
rect -27072 4310 -27036 4344
rect -29100 4299 -29046 4310
rect -29012 4299 -28958 4310
rect -28924 4299 -28870 4310
rect -28836 4299 -27036 4310
rect -31764 4298 -27036 4299
rect -32352 4276 -27036 4298
rect -32352 4275 -31632 4276
rect -32352 4259 -32315 4275
rect -32281 4259 -32247 4275
rect -32213 4259 -32179 4275
rect -32352 4225 -32344 4259
rect -32281 4241 -32266 4259
rect -32213 4241 -32188 4259
rect -32145 4241 -32111 4275
rect -32077 4259 -32043 4275
rect -32009 4259 -31975 4275
rect -31941 4259 -31907 4275
rect -31873 4259 -31839 4275
rect -32076 4241 -32043 4259
rect -31998 4241 -31975 4259
rect -31920 4241 -31907 4259
rect -31842 4241 -31839 4259
rect -31805 4259 -31771 4275
rect -31737 4261 -31703 4275
rect -31669 4261 -31632 4275
rect -31598 4261 -31563 4276
rect -31529 4261 -31494 4276
rect -31460 4261 -31425 4276
rect -31805 4241 -31798 4259
rect -31737 4241 -31718 4261
rect -31669 4241 -31645 4261
rect -31598 4242 -31572 4261
rect -31529 4242 -31499 4261
rect -31460 4242 -31426 4261
rect -31391 4242 -31356 4276
rect -31322 4261 -31287 4276
rect -31253 4261 -31218 4276
rect -31184 4261 -31149 4276
rect -31115 4261 -31080 4276
rect -31046 4261 -31011 4276
rect -30977 4261 -30942 4276
rect -30908 4261 -30873 4276
rect -30839 4261 -30804 4276
rect -31319 4242 -31287 4261
rect -31246 4242 -31218 4261
rect -31173 4242 -31149 4261
rect -31100 4242 -31080 4261
rect -31027 4242 -31011 4261
rect -30954 4242 -30942 4261
rect -30881 4242 -30873 4261
rect -30808 4242 -30804 4261
rect -30770 4261 -30735 4276
rect -30701 4261 -30666 4276
rect -30632 4261 -30597 4276
rect -30563 4261 -30528 4276
rect -30494 4261 -30459 4276
rect -30425 4261 -30390 4276
rect -30356 4261 -30321 4276
rect -30770 4242 -30768 4261
rect -30701 4242 -30694 4261
rect -30632 4242 -30620 4261
rect -30563 4242 -30546 4261
rect -30494 4242 -30472 4261
rect -30425 4242 -30398 4261
rect -30356 4242 -30324 4261
rect -30287 4242 -30252 4276
rect -30218 4261 -30183 4276
rect -30149 4261 -30114 4276
rect -30080 4261 -30045 4276
rect -30011 4261 -29976 4276
rect -29942 4261 -29907 4276
rect -29873 4261 -29838 4276
rect -29804 4261 -29769 4276
rect -30216 4242 -30183 4261
rect -30142 4242 -30114 4261
rect -30068 4242 -30045 4261
rect -29994 4242 -29976 4261
rect -29920 4242 -29907 4261
rect -29846 4242 -29838 4261
rect -29772 4242 -29769 4261
rect -29735 4261 -29700 4276
rect -29666 4261 -29631 4276
rect -29597 4261 -29562 4276
rect -29528 4261 -29493 4276
rect -29459 4261 -29424 4276
rect -29390 4261 -29355 4276
rect -29321 4261 -29286 4276
rect -29735 4242 -29732 4261
rect -29666 4242 -29658 4261
rect -29597 4242 -29584 4261
rect -29528 4242 -29510 4261
rect -29459 4242 -29436 4261
rect -29390 4242 -29362 4261
rect -29321 4242 -29288 4261
rect -29252 4242 -29217 4276
rect -29183 4261 -29148 4276
rect -29180 4242 -29148 4261
rect -29114 4275 -27036 4276
rect -29114 4260 -29078 4275
rect -29044 4260 -29010 4275
rect -32310 4225 -32266 4241
rect -32232 4225 -32188 4241
rect -32154 4225 -32110 4241
rect -32076 4225 -32032 4241
rect -31998 4225 -31954 4241
rect -31920 4225 -31876 4241
rect -31842 4225 -31798 4241
rect -31764 4227 -31718 4241
rect -31684 4227 -31645 4241
rect -31611 4227 -31572 4242
rect -31538 4227 -31499 4242
rect -31465 4227 -31426 4242
rect -31392 4227 -31353 4242
rect -31319 4227 -31280 4242
rect -31246 4227 -31207 4242
rect -31173 4227 -31134 4242
rect -31100 4227 -31061 4242
rect -31027 4227 -30988 4242
rect -30954 4227 -30915 4242
rect -30881 4227 -30842 4242
rect -30808 4227 -30768 4242
rect -30734 4227 -30694 4242
rect -30660 4227 -30620 4242
rect -30586 4227 -30546 4242
rect -30512 4227 -30472 4242
rect -30438 4227 -30398 4242
rect -30364 4227 -30324 4242
rect -30290 4227 -30250 4242
rect -30216 4227 -30176 4242
rect -30142 4227 -30102 4242
rect -30068 4227 -30028 4242
rect -29994 4227 -29954 4242
rect -29920 4227 -29880 4242
rect -29846 4227 -29806 4242
rect -29772 4227 -29732 4242
rect -29698 4227 -29658 4242
rect -29624 4227 -29584 4242
rect -29550 4227 -29510 4242
rect -29476 4227 -29436 4242
rect -29402 4227 -29362 4242
rect -29328 4227 -29288 4242
rect -29254 4227 -29214 4242
rect -29180 4227 -29134 4242
rect -31764 4226 -29134 4227
rect -29100 4241 -29078 4260
rect -29012 4241 -29010 4260
rect -28976 4260 -28942 4275
rect -28976 4241 -28958 4260
rect -28908 4241 -28874 4275
rect -28840 4260 -28806 4275
rect -28836 4241 -28806 4260
rect -28772 4241 -28738 4275
rect -28704 4241 -28670 4275
rect -28636 4241 -28602 4275
rect -28568 4241 -28534 4275
rect -28500 4241 -28466 4275
rect -28432 4241 -28398 4275
rect -28364 4241 -28330 4275
rect -28296 4241 -28262 4275
rect -28228 4241 -28194 4275
rect -28160 4241 -28126 4275
rect -28092 4241 -28058 4275
rect -28024 4241 -27990 4275
rect -27956 4241 -27922 4275
rect -27888 4241 -27854 4275
rect -27820 4241 -27786 4275
rect -27752 4241 -27718 4275
rect -27684 4241 -27650 4275
rect -27616 4241 -27582 4275
rect -27548 4241 -27514 4275
rect -27480 4241 -27446 4275
rect -27412 4241 -27378 4275
rect -27344 4241 -27310 4275
rect -27276 4241 -27242 4275
rect -27208 4241 -27174 4275
rect -27140 4241 -27106 4275
rect -27072 4241 -27036 4275
rect -29100 4226 -29046 4241
rect -29012 4226 -28958 4241
rect -28924 4226 -28870 4241
rect -28836 4239 -27036 4241
rect -28836 4226 -28189 4239
rect -31764 4225 -28189 4226
rect -32352 4206 -28189 4225
rect -28155 4206 -28115 4239
rect -28081 4206 -28041 4239
rect -28007 4206 -27967 4239
rect -27933 4206 -27893 4239
rect -27859 4206 -27819 4239
rect -27785 4206 -27745 4239
rect -27711 4206 -27671 4239
rect -27637 4206 -27597 4239
rect -27563 4206 -27523 4239
rect -27489 4206 -27449 4239
rect -27415 4206 -27375 4239
rect -27341 4206 -27301 4239
rect -27267 4206 -27227 4239
rect -27193 4206 -27153 4239
rect -27119 4206 -27036 4239
rect -32352 4186 -32315 4206
rect -32281 4186 -32247 4206
rect -32213 4186 -32179 4206
rect -32352 4152 -32344 4186
rect -32281 4172 -32266 4186
rect -32213 4172 -32188 4186
rect -32145 4172 -32111 4206
rect -32077 4186 -32043 4206
rect -32009 4186 -31975 4206
rect -31941 4186 -31907 4206
rect -31873 4186 -31839 4206
rect -32076 4172 -32043 4186
rect -31998 4172 -31975 4186
rect -31920 4172 -31907 4186
rect -31842 4172 -31839 4186
rect -31805 4186 -31771 4206
rect -31737 4189 -31703 4206
rect -31669 4189 -31632 4206
rect -31598 4189 -31563 4206
rect -31529 4189 -31494 4206
rect -31460 4189 -31425 4206
rect -31805 4172 -31798 4186
rect -31737 4172 -31718 4189
rect -31669 4172 -31645 4189
rect -31598 4172 -31572 4189
rect -31529 4172 -31499 4189
rect -31460 4172 -31426 4189
rect -31391 4172 -31356 4206
rect -31322 4189 -31287 4206
rect -31253 4189 -31218 4206
rect -31184 4189 -31149 4206
rect -31115 4189 -31080 4206
rect -31046 4189 -31011 4206
rect -30977 4189 -30942 4206
rect -30908 4189 -30873 4206
rect -30839 4189 -30804 4206
rect -31319 4172 -31287 4189
rect -31246 4172 -31218 4189
rect -31173 4172 -31149 4189
rect -31100 4172 -31080 4189
rect -31027 4172 -31011 4189
rect -30954 4172 -30942 4189
rect -30881 4172 -30873 4189
rect -30808 4172 -30804 4189
rect -30770 4189 -30735 4206
rect -30701 4189 -30666 4206
rect -30632 4189 -30597 4206
rect -30563 4189 -30528 4206
rect -30494 4189 -30459 4206
rect -30425 4189 -30390 4206
rect -30356 4189 -30321 4206
rect -30770 4172 -30768 4189
rect -30701 4172 -30694 4189
rect -30632 4172 -30620 4189
rect -30563 4172 -30546 4189
rect -30494 4172 -30472 4189
rect -30425 4172 -30398 4189
rect -30356 4172 -30324 4189
rect -30287 4172 -30252 4206
rect -30218 4189 -30183 4206
rect -30149 4189 -30114 4206
rect -30080 4189 -30045 4206
rect -30011 4189 -29976 4206
rect -29942 4189 -29907 4206
rect -29873 4189 -29838 4206
rect -29804 4189 -29769 4206
rect -30216 4172 -30183 4189
rect -30142 4172 -30114 4189
rect -30068 4172 -30045 4189
rect -29994 4172 -29976 4189
rect -29920 4172 -29907 4189
rect -29846 4172 -29838 4189
rect -29772 4172 -29769 4189
rect -29735 4189 -29700 4206
rect -29666 4189 -29631 4206
rect -29597 4189 -29562 4206
rect -29528 4189 -29493 4206
rect -29459 4189 -29424 4206
rect -29390 4189 -29355 4206
rect -29321 4189 -29286 4206
rect -29735 4172 -29732 4189
rect -29666 4172 -29658 4189
rect -29597 4172 -29584 4189
rect -29528 4172 -29510 4189
rect -29459 4172 -29436 4189
rect -29390 4172 -29362 4189
rect -29321 4172 -29288 4189
rect -29252 4172 -29217 4206
rect -29183 4189 -29148 4206
rect -29180 4172 -29148 4189
rect -29114 4187 -29078 4206
rect -29044 4187 -29010 4206
rect -29100 4172 -29078 4187
rect -29012 4172 -29010 4187
rect -28976 4187 -28942 4206
rect -28976 4172 -28958 4187
rect -28908 4172 -28874 4206
rect -28840 4187 -28806 4206
rect -28836 4172 -28806 4187
rect -28772 4172 -28738 4206
rect -28704 4172 -28670 4206
rect -28636 4172 -28602 4206
rect -28568 4172 -28534 4206
rect -28500 4172 -28466 4206
rect -28432 4172 -28398 4206
rect -28364 4172 -28330 4206
rect -28296 4172 -28262 4206
rect -28228 4172 -28194 4206
rect -28155 4205 -28126 4206
rect -28081 4205 -28058 4206
rect -28007 4205 -27990 4206
rect -27933 4205 -27922 4206
rect -27859 4205 -27854 4206
rect -28160 4172 -28126 4205
rect -28092 4172 -28058 4205
rect -28024 4172 -27990 4205
rect -27956 4172 -27922 4205
rect -27888 4172 -27854 4205
rect -27820 4205 -27819 4206
rect -27752 4205 -27745 4206
rect -27684 4205 -27671 4206
rect -27616 4205 -27597 4206
rect -27548 4205 -27523 4206
rect -27480 4205 -27449 4206
rect -27820 4172 -27786 4205
rect -27752 4172 -27718 4205
rect -27684 4172 -27650 4205
rect -27616 4172 -27582 4205
rect -27548 4172 -27514 4205
rect -27480 4172 -27446 4205
rect -27412 4172 -27378 4206
rect -27341 4205 -27310 4206
rect -27267 4205 -27242 4206
rect -27193 4205 -27174 4206
rect -27119 4205 -27106 4206
rect -27344 4172 -27310 4205
rect -27276 4172 -27242 4205
rect -27208 4172 -27174 4205
rect -27140 4172 -27106 4205
rect -27072 4172 -27036 4206
rect -9806 4312 -9740 4328
rect -9806 4278 -9790 4312
rect -9756 4278 -9740 4312
rect -9806 4244 -9740 4278
rect -9806 4206 -9790 4244
rect -9756 4206 -9740 4244
rect -9806 4194 -9740 4206
rect -32310 4152 -32266 4172
rect -32232 4152 -32188 4172
rect -32154 4152 -32110 4172
rect -32076 4152 -32032 4172
rect -31998 4152 -31954 4172
rect -31920 4152 -31876 4172
rect -31842 4152 -31798 4172
rect -31764 4155 -31718 4172
rect -31684 4155 -31645 4172
rect -31611 4155 -31572 4172
rect -31538 4155 -31499 4172
rect -31465 4155 -31426 4172
rect -31392 4155 -31353 4172
rect -31319 4155 -31280 4172
rect -31246 4155 -31207 4172
rect -31173 4155 -31134 4172
rect -31100 4155 -31061 4172
rect -31027 4155 -30988 4172
rect -30954 4155 -30915 4172
rect -30881 4155 -30842 4172
rect -30808 4155 -30768 4172
rect -30734 4155 -30694 4172
rect -30660 4155 -30620 4172
rect -30586 4155 -30546 4172
rect -30512 4155 -30472 4172
rect -30438 4155 -30398 4172
rect -30364 4155 -30324 4172
rect -30290 4155 -30250 4172
rect -30216 4155 -30176 4172
rect -30142 4155 -30102 4172
rect -30068 4155 -30028 4172
rect -29994 4155 -29954 4172
rect -29920 4155 -29880 4172
rect -29846 4155 -29806 4172
rect -29772 4155 -29732 4172
rect -29698 4155 -29658 4172
rect -29624 4155 -29584 4172
rect -29550 4155 -29510 4172
rect -29476 4155 -29436 4172
rect -29402 4155 -29362 4172
rect -29328 4155 -29288 4172
rect -29254 4155 -29214 4172
rect -29180 4155 -29134 4172
rect -31764 4153 -29134 4155
rect -29100 4153 -29046 4172
rect -29012 4153 -28958 4172
rect -28924 4153 -28870 4172
rect -28836 4166 -27036 4172
rect -28836 4153 -28189 4166
rect -31764 4152 -28189 4153
rect -32352 4137 -28189 4152
rect -28155 4137 -28115 4166
rect -28081 4137 -28041 4166
rect -28007 4137 -27967 4166
rect -27933 4137 -27893 4166
rect -27859 4137 -27819 4166
rect -27785 4137 -27745 4166
rect -27711 4137 -27671 4166
rect -27637 4137 -27597 4166
rect -27563 4137 -27523 4166
rect -27489 4137 -27449 4166
rect -27415 4137 -27375 4166
rect -27341 4137 -27301 4166
rect -27267 4137 -27227 4166
rect -27193 4137 -27153 4166
rect -27119 4137 -27036 4166
rect -32352 4113 -32315 4137
rect -32281 4113 -32247 4137
rect -32213 4113 -32179 4137
rect -32352 4079 -32344 4113
rect -32281 4103 -32266 4113
rect -32213 4103 -32188 4113
rect -32145 4103 -32111 4137
rect -32077 4113 -32043 4137
rect -32009 4113 -31975 4137
rect -31941 4113 -31907 4137
rect -31873 4113 -31839 4137
rect -32076 4103 -32043 4113
rect -31998 4103 -31975 4113
rect -31920 4103 -31907 4113
rect -31842 4103 -31839 4113
rect -31805 4113 -31771 4137
rect -31737 4117 -31703 4137
rect -31669 4136 -29078 4137
rect -31669 4117 -31632 4136
rect -31598 4117 -31563 4136
rect -31529 4117 -31494 4136
rect -31460 4117 -31425 4136
rect -31805 4103 -31798 4113
rect -31737 4103 -31718 4117
rect -31669 4103 -31645 4117
rect -32310 4079 -32266 4103
rect -32232 4079 -32188 4103
rect -32154 4079 -32110 4103
rect -32076 4079 -32032 4103
rect -31998 4079 -31954 4103
rect -31920 4079 -31876 4103
rect -31842 4079 -31798 4103
rect -31764 4083 -31718 4103
rect -31684 4083 -31645 4103
rect -31598 4102 -31572 4117
rect -31529 4102 -31499 4117
rect -31460 4102 -31426 4117
rect -31391 4102 -31356 4136
rect -31322 4117 -31287 4136
rect -31253 4117 -31218 4136
rect -31184 4117 -31149 4136
rect -31115 4117 -31080 4136
rect -31046 4117 -31011 4136
rect -30977 4117 -30942 4136
rect -30908 4117 -30873 4136
rect -30839 4117 -30804 4136
rect -31319 4102 -31287 4117
rect -31246 4102 -31218 4117
rect -31173 4102 -31149 4117
rect -31100 4102 -31080 4117
rect -31027 4102 -31011 4117
rect -30954 4102 -30942 4117
rect -30881 4102 -30873 4117
rect -30808 4102 -30804 4117
rect -30770 4117 -30735 4136
rect -30701 4117 -30666 4136
rect -30632 4117 -30597 4136
rect -30563 4117 -30528 4136
rect -30494 4117 -30459 4136
rect -30425 4117 -30390 4136
rect -30356 4117 -30321 4136
rect -30770 4102 -30768 4117
rect -30701 4102 -30694 4117
rect -30632 4102 -30620 4117
rect -30563 4102 -30546 4117
rect -30494 4102 -30472 4117
rect -30425 4102 -30398 4117
rect -30356 4102 -30324 4117
rect -30287 4102 -30252 4136
rect -30218 4117 -30183 4136
rect -30149 4117 -30114 4136
rect -30080 4117 -30045 4136
rect -30011 4117 -29976 4136
rect -29942 4117 -29907 4136
rect -29873 4117 -29838 4136
rect -29804 4117 -29769 4136
rect -30216 4102 -30183 4117
rect -30142 4102 -30114 4117
rect -30068 4102 -30045 4117
rect -29994 4102 -29976 4117
rect -29920 4102 -29907 4117
rect -29846 4102 -29838 4117
rect -29772 4102 -29769 4117
rect -29735 4117 -29700 4136
rect -29666 4117 -29631 4136
rect -29597 4117 -29562 4136
rect -29528 4117 -29493 4136
rect -29459 4117 -29424 4136
rect -29390 4117 -29355 4136
rect -29321 4117 -29286 4136
rect -29735 4102 -29732 4117
rect -29666 4102 -29658 4117
rect -29597 4102 -29584 4117
rect -29528 4102 -29510 4117
rect -29459 4102 -29436 4117
rect -29390 4102 -29362 4117
rect -29321 4102 -29288 4117
rect -29252 4102 -29217 4136
rect -29183 4117 -29148 4136
rect -29180 4102 -29148 4117
rect -29114 4114 -29078 4136
rect -29044 4114 -29010 4137
rect -29100 4103 -29078 4114
rect -29012 4103 -29010 4114
rect -28976 4114 -28942 4137
rect -28976 4103 -28958 4114
rect -28908 4103 -28874 4137
rect -28840 4114 -28806 4137
rect -28836 4103 -28806 4114
rect -28772 4103 -28738 4137
rect -28704 4103 -28670 4137
rect -28636 4103 -28602 4137
rect -28568 4103 -28534 4137
rect -28500 4103 -28466 4137
rect -28432 4103 -28398 4137
rect -28364 4103 -28330 4137
rect -28296 4103 -28262 4137
rect -28228 4103 -28194 4137
rect -28155 4132 -28126 4137
rect -28081 4132 -28058 4137
rect -28007 4132 -27990 4137
rect -27933 4132 -27922 4137
rect -27859 4132 -27854 4137
rect -28160 4103 -28126 4132
rect -28092 4103 -28058 4132
rect -28024 4103 -27990 4132
rect -27956 4103 -27922 4132
rect -27888 4103 -27854 4132
rect -27820 4132 -27819 4137
rect -27752 4132 -27745 4137
rect -27684 4132 -27671 4137
rect -27616 4132 -27597 4137
rect -27548 4132 -27523 4137
rect -27480 4132 -27449 4137
rect -27820 4103 -27786 4132
rect -27752 4103 -27718 4132
rect -27684 4103 -27650 4132
rect -27616 4103 -27582 4132
rect -27548 4103 -27514 4132
rect -27480 4103 -27446 4132
rect -27412 4103 -27378 4137
rect -27341 4132 -27310 4137
rect -27267 4132 -27242 4137
rect -27193 4132 -27174 4137
rect -27119 4132 -27106 4137
rect -27344 4103 -27310 4132
rect -27276 4103 -27242 4132
rect -27208 4103 -27174 4132
rect -27140 4103 -27106 4132
rect -27072 4103 -27036 4137
rect -31611 4083 -31572 4102
rect -31538 4083 -31499 4102
rect -31465 4083 -31426 4102
rect -31392 4083 -31353 4102
rect -31319 4083 -31280 4102
rect -31246 4083 -31207 4102
rect -31173 4083 -31134 4102
rect -31100 4083 -31061 4102
rect -31027 4083 -30988 4102
rect -30954 4083 -30915 4102
rect -30881 4083 -30842 4102
rect -30808 4083 -30768 4102
rect -30734 4083 -30694 4102
rect -30660 4083 -30620 4102
rect -30586 4083 -30546 4102
rect -30512 4083 -30472 4102
rect -30438 4083 -30398 4102
rect -30364 4083 -30324 4102
rect -30290 4083 -30250 4102
rect -30216 4083 -30176 4102
rect -30142 4083 -30102 4102
rect -30068 4083 -30028 4102
rect -29994 4083 -29954 4102
rect -29920 4083 -29880 4102
rect -29846 4083 -29806 4102
rect -29772 4083 -29732 4102
rect -29698 4083 -29658 4102
rect -29624 4083 -29584 4102
rect -29550 4083 -29510 4102
rect -29476 4083 -29436 4102
rect -29402 4083 -29362 4102
rect -29328 4083 -29288 4102
rect -29254 4083 -29214 4102
rect -29180 4083 -29134 4102
rect -31764 4080 -29134 4083
rect -29100 4080 -29046 4103
rect -29012 4080 -28958 4103
rect -28924 4080 -28870 4103
rect -28836 4093 -27036 4103
rect -28836 4080 -28189 4093
rect -31764 4079 -28189 4080
rect -32352 4068 -28189 4079
rect -28155 4068 -28115 4093
rect -28081 4068 -28041 4093
rect -28007 4068 -27967 4093
rect -27933 4068 -27893 4093
rect -27859 4068 -27819 4093
rect -27785 4068 -27745 4093
rect -27711 4068 -27671 4093
rect -27637 4068 -27597 4093
rect -27563 4068 -27523 4093
rect -27489 4068 -27449 4093
rect -27415 4068 -27375 4093
rect -27341 4068 -27301 4093
rect -27267 4068 -27227 4093
rect -27193 4068 -27153 4093
rect -27119 4068 -27036 4093
rect -32352 4040 -32315 4068
rect -32281 4040 -32247 4068
rect -32213 4040 -32179 4068
rect -32352 4006 -32344 4040
rect -32281 4034 -32266 4040
rect -32213 4034 -32188 4040
rect -32145 4034 -32111 4068
rect -32077 4040 -32043 4068
rect -32009 4040 -31975 4068
rect -31941 4040 -31907 4068
rect -31873 4040 -31839 4068
rect -32076 4034 -32043 4040
rect -31998 4034 -31975 4040
rect -31920 4034 -31907 4040
rect -31842 4034 -31839 4040
rect -31805 4040 -31771 4068
rect -31737 4045 -31703 4068
rect -31669 4066 -29078 4068
rect -31669 4045 -31632 4066
rect -31598 4045 -31563 4066
rect -31529 4045 -31494 4066
rect -31460 4045 -31425 4066
rect -31805 4034 -31798 4040
rect -31737 4034 -31718 4045
rect -31669 4034 -31645 4045
rect -32310 4006 -32266 4034
rect -32232 4006 -32188 4034
rect -32154 4006 -32110 4034
rect -32076 4006 -32032 4034
rect -31998 4006 -31954 4034
rect -31920 4006 -31876 4034
rect -31842 4006 -31798 4034
rect -31764 4011 -31718 4034
rect -31684 4011 -31645 4034
rect -31598 4032 -31572 4045
rect -31529 4032 -31499 4045
rect -31460 4032 -31426 4045
rect -31391 4032 -31356 4066
rect -31322 4045 -31287 4066
rect -31253 4045 -31218 4066
rect -31184 4045 -31149 4066
rect -31115 4045 -31080 4066
rect -31046 4045 -31011 4066
rect -30977 4045 -30942 4066
rect -30908 4045 -30873 4066
rect -30839 4045 -30804 4066
rect -31319 4032 -31287 4045
rect -31246 4032 -31218 4045
rect -31173 4032 -31149 4045
rect -31100 4032 -31080 4045
rect -31027 4032 -31011 4045
rect -30954 4032 -30942 4045
rect -30881 4032 -30873 4045
rect -30808 4032 -30804 4045
rect -30770 4045 -30735 4066
rect -30701 4045 -30666 4066
rect -30632 4045 -30597 4066
rect -30563 4045 -30528 4066
rect -30494 4045 -30459 4066
rect -30425 4045 -30390 4066
rect -30356 4045 -30321 4066
rect -30770 4032 -30768 4045
rect -30701 4032 -30694 4045
rect -30632 4032 -30620 4045
rect -30563 4032 -30546 4045
rect -30494 4032 -30472 4045
rect -30425 4032 -30398 4045
rect -30356 4032 -30324 4045
rect -30287 4032 -30252 4066
rect -30218 4045 -30183 4066
rect -30149 4045 -30114 4066
rect -30080 4045 -30045 4066
rect -30011 4045 -29976 4066
rect -29942 4045 -29907 4066
rect -29873 4045 -29838 4066
rect -29804 4045 -29769 4066
rect -30216 4032 -30183 4045
rect -30142 4032 -30114 4045
rect -30068 4032 -30045 4045
rect -29994 4032 -29976 4045
rect -29920 4032 -29907 4045
rect -29846 4032 -29838 4045
rect -29772 4032 -29769 4045
rect -29735 4045 -29700 4066
rect -29666 4045 -29631 4066
rect -29597 4045 -29562 4066
rect -29528 4045 -29493 4066
rect -29459 4045 -29424 4066
rect -29390 4045 -29355 4066
rect -29321 4045 -29286 4066
rect -29735 4032 -29732 4045
rect -29666 4032 -29658 4045
rect -29597 4032 -29584 4045
rect -29528 4032 -29510 4045
rect -29459 4032 -29436 4045
rect -29390 4032 -29362 4045
rect -29321 4032 -29288 4045
rect -29252 4032 -29217 4066
rect -29183 4045 -29148 4066
rect -29180 4032 -29148 4045
rect -29114 4041 -29078 4066
rect -29044 4041 -29010 4068
rect -29100 4034 -29078 4041
rect -29012 4034 -29010 4041
rect -28976 4041 -28942 4068
rect -28976 4034 -28958 4041
rect -28908 4034 -28874 4068
rect -28840 4041 -28806 4068
rect -28836 4034 -28806 4041
rect -28772 4034 -28738 4068
rect -28704 4034 -28670 4068
rect -28636 4034 -28602 4068
rect -28568 4034 -28534 4068
rect -28500 4034 -28466 4068
rect -28432 4034 -28398 4068
rect -28364 4034 -28330 4068
rect -28296 4034 -28262 4068
rect -28228 4034 -28194 4068
rect -28155 4059 -28126 4068
rect -28081 4059 -28058 4068
rect -28007 4059 -27990 4068
rect -27933 4059 -27922 4068
rect -27859 4059 -27854 4068
rect -28160 4034 -28126 4059
rect -28092 4034 -28058 4059
rect -28024 4034 -27990 4059
rect -27956 4034 -27922 4059
rect -27888 4034 -27854 4059
rect -27820 4059 -27819 4068
rect -27752 4059 -27745 4068
rect -27684 4059 -27671 4068
rect -27616 4059 -27597 4068
rect -27548 4059 -27523 4068
rect -27480 4059 -27449 4068
rect -27820 4034 -27786 4059
rect -27752 4034 -27718 4059
rect -27684 4034 -27650 4059
rect -27616 4034 -27582 4059
rect -27548 4034 -27514 4059
rect -27480 4034 -27446 4059
rect -27412 4034 -27378 4068
rect -27341 4059 -27310 4068
rect -27267 4059 -27242 4068
rect -27193 4059 -27174 4068
rect -27119 4059 -27106 4068
rect -27344 4034 -27310 4059
rect -27276 4034 -27242 4059
rect -27208 4034 -27174 4059
rect -27140 4034 -27106 4059
rect -27072 4034 -27036 4068
rect -31611 4011 -31572 4032
rect -31538 4011 -31499 4032
rect -31465 4011 -31426 4032
rect -31392 4011 -31353 4032
rect -31319 4011 -31280 4032
rect -31246 4011 -31207 4032
rect -31173 4011 -31134 4032
rect -31100 4011 -31061 4032
rect -31027 4011 -30988 4032
rect -30954 4011 -30915 4032
rect -30881 4011 -30842 4032
rect -30808 4011 -30768 4032
rect -30734 4011 -30694 4032
rect -30660 4011 -30620 4032
rect -30586 4011 -30546 4032
rect -30512 4011 -30472 4032
rect -30438 4011 -30398 4032
rect -30364 4011 -30324 4032
rect -30290 4011 -30250 4032
rect -30216 4011 -30176 4032
rect -30142 4011 -30102 4032
rect -30068 4011 -30028 4032
rect -29994 4011 -29954 4032
rect -29920 4011 -29880 4032
rect -29846 4011 -29806 4032
rect -29772 4011 -29732 4032
rect -29698 4011 -29658 4032
rect -29624 4011 -29584 4032
rect -29550 4011 -29510 4032
rect -29476 4011 -29436 4032
rect -29402 4011 -29362 4032
rect -29328 4011 -29288 4032
rect -29254 4011 -29214 4032
rect -29180 4011 -29134 4032
rect -31764 4007 -29134 4011
rect -29100 4007 -29046 4034
rect -29012 4007 -28958 4034
rect -28924 4007 -28870 4034
rect -28836 4020 -27036 4034
rect -28836 4007 -28189 4020
rect -31764 4006 -28189 4007
rect -32352 3999 -28189 4006
rect -28155 3999 -28115 4020
rect -28081 3999 -28041 4020
rect -28007 3999 -27967 4020
rect -27933 3999 -27893 4020
rect -27859 3999 -27819 4020
rect -27785 3999 -27745 4020
rect -27711 3999 -27671 4020
rect -27637 3999 -27597 4020
rect -27563 3999 -27523 4020
rect -27489 3999 -27449 4020
rect -27415 3999 -27375 4020
rect -27341 3999 -27301 4020
rect -27267 3999 -27227 4020
rect -27193 3999 -27153 4020
rect -27119 3999 -27036 4020
rect -32352 3967 -32315 3999
rect -31669 3996 -29078 3999
rect -31669 3973 -31632 3996
rect -31598 3973 -31563 3996
rect -31529 3973 -31494 3996
rect -31460 3973 -31425 3996
rect -32352 3933 -32344 3967
rect -31669 3939 -31645 3973
rect -31598 3962 -31572 3973
rect -31529 3962 -31499 3973
rect -31460 3962 -31426 3973
rect -31391 3962 -31356 3996
rect -31322 3973 -31287 3996
rect -31253 3973 -31218 3996
rect -31184 3973 -31149 3996
rect -31115 3973 -31080 3996
rect -31046 3973 -31011 3996
rect -30977 3973 -30942 3996
rect -30908 3973 -30873 3996
rect -30839 3973 -30804 3996
rect -31319 3962 -31287 3973
rect -31246 3962 -31218 3973
rect -31173 3962 -31149 3973
rect -31100 3962 -31080 3973
rect -31027 3962 -31011 3973
rect -30954 3962 -30942 3973
rect -30881 3962 -30873 3973
rect -30808 3962 -30804 3973
rect -30770 3973 -30735 3996
rect -30701 3973 -30666 3996
rect -30632 3973 -30597 3996
rect -30563 3973 -30528 3996
rect -30494 3973 -30459 3996
rect -30425 3973 -30390 3996
rect -30356 3973 -30321 3996
rect -30770 3962 -30768 3973
rect -30701 3962 -30694 3973
rect -30632 3962 -30620 3973
rect -30563 3962 -30546 3973
rect -30494 3962 -30472 3973
rect -30425 3962 -30398 3973
rect -30356 3962 -30324 3973
rect -30287 3962 -30252 3996
rect -30218 3973 -30183 3996
rect -30149 3973 -30114 3996
rect -30080 3973 -30045 3996
rect -30011 3973 -29976 3996
rect -29942 3973 -29907 3996
rect -29873 3973 -29838 3996
rect -29804 3973 -29769 3996
rect -30216 3962 -30183 3973
rect -30142 3962 -30114 3973
rect -30068 3962 -30045 3973
rect -29994 3962 -29976 3973
rect -29920 3962 -29907 3973
rect -29846 3962 -29838 3973
rect -29772 3962 -29769 3973
rect -29735 3973 -29700 3996
rect -29666 3973 -29631 3996
rect -29597 3973 -29562 3996
rect -29528 3973 -29493 3996
rect -29459 3973 -29424 3996
rect -29390 3973 -29355 3996
rect -29321 3973 -29286 3996
rect -29735 3962 -29732 3973
rect -29666 3962 -29658 3973
rect -29597 3962 -29584 3973
rect -29528 3962 -29510 3973
rect -29459 3962 -29436 3973
rect -29390 3962 -29362 3973
rect -29321 3962 -29288 3973
rect -29252 3962 -29217 3996
rect -29183 3973 -29148 3996
rect -29180 3962 -29148 3973
rect -29114 3968 -29078 3996
rect -29044 3968 -29010 3999
rect -29100 3965 -29078 3968
rect -29012 3965 -29010 3968
rect -28976 3968 -28942 3999
rect -28976 3965 -28958 3968
rect -28908 3965 -28874 3999
rect -28840 3968 -28806 3999
rect -28836 3965 -28806 3968
rect -28772 3965 -28738 3999
rect -28704 3965 -28670 3999
rect -28636 3965 -28602 3999
rect -28568 3965 -28534 3999
rect -28500 3965 -28466 3999
rect -28432 3965 -28398 3999
rect -28364 3965 -28330 3999
rect -28296 3965 -28262 3999
rect -28228 3965 -28194 3999
rect -28155 3986 -28126 3999
rect -28081 3986 -28058 3999
rect -28007 3986 -27990 3999
rect -27933 3986 -27922 3999
rect -27859 3986 -27854 3999
rect -28160 3965 -28126 3986
rect -28092 3965 -28058 3986
rect -28024 3965 -27990 3986
rect -27956 3965 -27922 3986
rect -27888 3965 -27854 3986
rect -27820 3986 -27819 3999
rect -27752 3986 -27745 3999
rect -27684 3986 -27671 3999
rect -27616 3986 -27597 3999
rect -27548 3986 -27523 3999
rect -27480 3986 -27449 3999
rect -27820 3965 -27786 3986
rect -27752 3965 -27718 3986
rect -27684 3965 -27650 3986
rect -27616 3965 -27582 3986
rect -27548 3965 -27514 3986
rect -27480 3965 -27446 3986
rect -27412 3965 -27378 3999
rect -27341 3986 -27310 3999
rect -27267 3986 -27242 3999
rect -27193 3986 -27174 3999
rect -27119 3986 -27106 3999
rect -27344 3965 -27310 3986
rect -27276 3965 -27242 3986
rect -27208 3965 -27174 3986
rect -27140 3965 -27106 3986
rect -27072 3965 -27036 3999
rect -31611 3939 -31572 3962
rect -31538 3939 -31499 3962
rect -31465 3939 -31426 3962
rect -31392 3939 -31353 3962
rect -31319 3939 -31280 3962
rect -31246 3939 -31207 3962
rect -31173 3939 -31134 3962
rect -31100 3939 -31061 3962
rect -31027 3939 -30988 3962
rect -30954 3939 -30915 3962
rect -30881 3939 -30842 3962
rect -30808 3939 -30768 3962
rect -30734 3939 -30694 3962
rect -30660 3939 -30620 3962
rect -30586 3939 -30546 3962
rect -30512 3939 -30472 3962
rect -30438 3939 -30398 3962
rect -30364 3939 -30324 3962
rect -30290 3939 -30250 3962
rect -30216 3939 -30176 3962
rect -30142 3939 -30102 3962
rect -30068 3939 -30028 3962
rect -29994 3939 -29954 3962
rect -29920 3939 -29880 3962
rect -29846 3939 -29806 3962
rect -29772 3939 -29732 3962
rect -29698 3939 -29658 3962
rect -29624 3939 -29584 3962
rect -29550 3939 -29510 3962
rect -29476 3939 -29436 3962
rect -29402 3939 -29362 3962
rect -29328 3939 -29288 3962
rect -29254 3939 -29214 3962
rect -29180 3939 -29134 3962
rect -31669 3934 -29134 3939
rect -29100 3934 -29046 3965
rect -29012 3934 -28958 3965
rect -28924 3934 -28870 3965
rect -28836 3947 -27036 3965
rect -28836 3934 -28189 3947
rect -32352 3894 -32315 3933
rect -31669 3930 -28189 3934
rect -28155 3930 -28115 3947
rect -28081 3930 -28041 3947
rect -28007 3930 -27967 3947
rect -27933 3930 -27893 3947
rect -27859 3930 -27819 3947
rect -27785 3930 -27745 3947
rect -27711 3930 -27671 3947
rect -27637 3930 -27597 3947
rect -27563 3930 -27523 3947
rect -27489 3930 -27449 3947
rect -27415 3930 -27375 3947
rect -27341 3930 -27301 3947
rect -27267 3930 -27227 3947
rect -27193 3930 -27153 3947
rect -27119 3930 -27036 3947
rect -31669 3926 -29078 3930
rect -31669 3901 -31632 3926
rect -31598 3901 -31563 3926
rect -31529 3901 -31494 3926
rect -31460 3901 -31425 3926
rect -32352 3860 -32344 3894
rect -31669 3867 -31645 3901
rect -31598 3892 -31572 3901
rect -31529 3892 -31499 3901
rect -31460 3892 -31426 3901
rect -31391 3892 -31356 3926
rect -31322 3901 -31287 3926
rect -31253 3901 -31218 3926
rect -31184 3901 -31149 3926
rect -31115 3901 -31080 3926
rect -31046 3901 -31011 3926
rect -30977 3901 -30942 3926
rect -30908 3901 -30873 3926
rect -30839 3901 -30804 3926
rect -31319 3892 -31287 3901
rect -31246 3892 -31218 3901
rect -31173 3892 -31149 3901
rect -31100 3892 -31080 3901
rect -31027 3892 -31011 3901
rect -30954 3892 -30942 3901
rect -30881 3892 -30873 3901
rect -30808 3892 -30804 3901
rect -30770 3901 -30735 3926
rect -30701 3901 -30666 3926
rect -30632 3901 -30597 3926
rect -30563 3901 -30528 3926
rect -30494 3901 -30459 3926
rect -30425 3901 -30390 3926
rect -30356 3901 -30321 3926
rect -30770 3892 -30768 3901
rect -30701 3892 -30694 3901
rect -30632 3892 -30620 3901
rect -30563 3892 -30546 3901
rect -30494 3892 -30472 3901
rect -30425 3892 -30398 3901
rect -30356 3892 -30324 3901
rect -30287 3892 -30252 3926
rect -30218 3901 -30183 3926
rect -30149 3901 -30114 3926
rect -30080 3901 -30045 3926
rect -30011 3901 -29976 3926
rect -29942 3901 -29907 3926
rect -29873 3901 -29838 3926
rect -29804 3901 -29769 3926
rect -30216 3892 -30183 3901
rect -30142 3892 -30114 3901
rect -30068 3892 -30045 3901
rect -29994 3892 -29976 3901
rect -29920 3892 -29907 3901
rect -29846 3892 -29838 3901
rect -29772 3892 -29769 3901
rect -29735 3901 -29700 3926
rect -29666 3901 -29631 3926
rect -29597 3901 -29562 3926
rect -29528 3901 -29493 3926
rect -29459 3901 -29424 3926
rect -29390 3901 -29355 3926
rect -29321 3901 -29286 3926
rect -29735 3892 -29732 3901
rect -29666 3892 -29658 3901
rect -29597 3892 -29584 3901
rect -29528 3892 -29510 3901
rect -29459 3892 -29436 3901
rect -29390 3892 -29362 3901
rect -29321 3892 -29288 3901
rect -29252 3892 -29217 3926
rect -29183 3901 -29148 3926
rect -29180 3892 -29148 3901
rect -29114 3896 -29078 3926
rect -29044 3896 -29010 3930
rect -28976 3896 -28942 3930
rect -28908 3896 -28874 3930
rect -28840 3896 -28806 3930
rect -28772 3896 -28738 3930
rect -28704 3896 -28670 3930
rect -28636 3896 -28602 3930
rect -28568 3896 -28534 3930
rect -28500 3896 -28466 3930
rect -28432 3896 -28398 3930
rect -28364 3896 -28330 3930
rect -28296 3896 -28262 3930
rect -28228 3896 -28194 3930
rect -28155 3913 -28126 3930
rect -28081 3913 -28058 3930
rect -28007 3913 -27990 3930
rect -27933 3913 -27922 3930
rect -27859 3913 -27854 3930
rect -28160 3896 -28126 3913
rect -28092 3896 -28058 3913
rect -28024 3896 -27990 3913
rect -27956 3896 -27922 3913
rect -27888 3896 -27854 3913
rect -27820 3913 -27819 3930
rect -27752 3913 -27745 3930
rect -27684 3913 -27671 3930
rect -27616 3913 -27597 3930
rect -27548 3913 -27523 3930
rect -27480 3913 -27449 3930
rect -27820 3896 -27786 3913
rect -27752 3896 -27718 3913
rect -27684 3896 -27650 3913
rect -27616 3896 -27582 3913
rect -27548 3896 -27514 3913
rect -27480 3896 -27446 3913
rect -27412 3896 -27378 3930
rect -27341 3913 -27310 3930
rect -27267 3913 -27242 3930
rect -27193 3913 -27174 3930
rect -27119 3913 -27106 3930
rect -27344 3896 -27310 3913
rect -27276 3896 -27242 3913
rect -27208 3896 -27174 3913
rect -27140 3896 -27106 3913
rect -27072 3896 -27036 3930
rect -29114 3895 -27036 3896
rect -31611 3867 -31572 3892
rect -31538 3867 -31499 3892
rect -31465 3867 -31426 3892
rect -31392 3867 -31353 3892
rect -31319 3867 -31280 3892
rect -31246 3867 -31207 3892
rect -31173 3867 -31134 3892
rect -31100 3867 -31061 3892
rect -31027 3867 -30988 3892
rect -30954 3867 -30915 3892
rect -30881 3867 -30842 3892
rect -30808 3867 -30768 3892
rect -30734 3867 -30694 3892
rect -30660 3867 -30620 3892
rect -30586 3867 -30546 3892
rect -30512 3867 -30472 3892
rect -30438 3867 -30398 3892
rect -30364 3867 -30324 3892
rect -30290 3867 -30250 3892
rect -30216 3867 -30176 3892
rect -30142 3867 -30102 3892
rect -30068 3867 -30028 3892
rect -29994 3867 -29954 3892
rect -29920 3867 -29880 3892
rect -29846 3867 -29806 3892
rect -29772 3867 -29732 3892
rect -29698 3867 -29658 3892
rect -29624 3867 -29584 3892
rect -29550 3867 -29510 3892
rect -29476 3867 -29436 3892
rect -29402 3867 -29362 3892
rect -29328 3867 -29288 3892
rect -29254 3867 -29214 3892
rect -29180 3867 -29134 3892
rect -31669 3861 -29134 3867
rect -29100 3861 -29046 3895
rect -29012 3861 -28958 3895
rect -28924 3861 -28870 3895
rect -28836 3874 -27036 3895
rect -28836 3861 -28189 3874
rect -28155 3861 -28115 3874
rect -28081 3861 -28041 3874
rect -28007 3861 -27967 3874
rect -27933 3861 -27893 3874
rect -27859 3861 -27819 3874
rect -27785 3861 -27745 3874
rect -27711 3861 -27671 3874
rect -27637 3861 -27597 3874
rect -27563 3861 -27523 3874
rect -27489 3861 -27449 3874
rect -27415 3861 -27375 3874
rect -27341 3861 -27301 3874
rect -27267 3861 -27227 3874
rect -27193 3861 -27153 3874
rect -27119 3861 -27036 3874
rect -32352 3821 -32315 3860
rect -31669 3856 -29078 3861
rect -31669 3829 -31632 3856
rect -31598 3829 -31563 3856
rect -31529 3829 -31494 3856
rect -31460 3829 -31425 3856
rect -32352 3787 -32344 3821
rect -31669 3795 -31645 3829
rect -31598 3822 -31572 3829
rect -31529 3822 -31499 3829
rect -31460 3822 -31426 3829
rect -31391 3822 -31356 3856
rect -31322 3829 -31287 3856
rect -31253 3829 -31218 3856
rect -31184 3829 -31149 3856
rect -31115 3829 -31080 3856
rect -31046 3829 -31011 3856
rect -30977 3829 -30942 3856
rect -30908 3829 -30873 3856
rect -30839 3829 -30804 3856
rect -31319 3822 -31287 3829
rect -31246 3822 -31218 3829
rect -31173 3822 -31149 3829
rect -31100 3822 -31080 3829
rect -31027 3822 -31011 3829
rect -30954 3822 -30942 3829
rect -30881 3822 -30873 3829
rect -30808 3822 -30804 3829
rect -30770 3829 -30735 3856
rect -30701 3829 -30666 3856
rect -30632 3829 -30597 3856
rect -30563 3829 -30528 3856
rect -30494 3829 -30459 3856
rect -30425 3829 -30390 3856
rect -30356 3829 -30321 3856
rect -30770 3822 -30768 3829
rect -30701 3822 -30694 3829
rect -30632 3822 -30620 3829
rect -30563 3822 -30546 3829
rect -30494 3822 -30472 3829
rect -30425 3822 -30398 3829
rect -30356 3822 -30324 3829
rect -30287 3822 -30252 3856
rect -30218 3829 -30183 3856
rect -30149 3829 -30114 3856
rect -30080 3829 -30045 3856
rect -30011 3829 -29976 3856
rect -29942 3829 -29907 3856
rect -29873 3829 -29838 3856
rect -29804 3829 -29769 3856
rect -30216 3822 -30183 3829
rect -30142 3822 -30114 3829
rect -30068 3822 -30045 3829
rect -29994 3822 -29976 3829
rect -29920 3822 -29907 3829
rect -29846 3822 -29838 3829
rect -29772 3822 -29769 3829
rect -29735 3829 -29700 3856
rect -29666 3829 -29631 3856
rect -29597 3829 -29562 3856
rect -29528 3829 -29493 3856
rect -29459 3829 -29424 3856
rect -29390 3829 -29355 3856
rect -29321 3829 -29286 3856
rect -29735 3822 -29732 3829
rect -29666 3822 -29658 3829
rect -29597 3822 -29584 3829
rect -29528 3822 -29510 3829
rect -29459 3822 -29436 3829
rect -29390 3822 -29362 3829
rect -29321 3822 -29288 3829
rect -29252 3822 -29217 3856
rect -29183 3829 -29148 3856
rect -29180 3822 -29148 3829
rect -29114 3827 -29078 3856
rect -29044 3827 -29010 3861
rect -28976 3827 -28942 3861
rect -28908 3827 -28874 3861
rect -28840 3827 -28806 3861
rect -28772 3827 -28738 3861
rect -28704 3827 -28670 3861
rect -28636 3827 -28602 3861
rect -28568 3827 -28534 3861
rect -28500 3827 -28466 3861
rect -28432 3827 -28398 3861
rect -28364 3827 -28330 3861
rect -28296 3827 -28262 3861
rect -28228 3827 -28194 3861
rect -28155 3840 -28126 3861
rect -28081 3840 -28058 3861
rect -28007 3840 -27990 3861
rect -27933 3840 -27922 3861
rect -27859 3840 -27854 3861
rect -28160 3827 -28126 3840
rect -28092 3827 -28058 3840
rect -28024 3827 -27990 3840
rect -27956 3827 -27922 3840
rect -27888 3827 -27854 3840
rect -27820 3840 -27819 3861
rect -27752 3840 -27745 3861
rect -27684 3840 -27671 3861
rect -27616 3840 -27597 3861
rect -27548 3840 -27523 3861
rect -27480 3840 -27449 3861
rect -27820 3827 -27786 3840
rect -27752 3827 -27718 3840
rect -27684 3827 -27650 3840
rect -27616 3827 -27582 3840
rect -27548 3827 -27514 3840
rect -27480 3827 -27446 3840
rect -27412 3827 -27378 3861
rect -27341 3840 -27310 3861
rect -27267 3840 -27242 3861
rect -27193 3840 -27174 3861
rect -27119 3840 -27106 3861
rect -27344 3827 -27310 3840
rect -27276 3827 -27242 3840
rect -27208 3827 -27174 3840
rect -27140 3827 -27106 3840
rect -27072 3827 -27036 3861
rect -29114 3822 -27036 3827
rect -31611 3795 -31572 3822
rect -31538 3795 -31499 3822
rect -31465 3795 -31426 3822
rect -31392 3795 -31353 3822
rect -31319 3795 -31280 3822
rect -31246 3795 -31207 3822
rect -31173 3795 -31134 3822
rect -31100 3795 -31061 3822
rect -31027 3795 -30988 3822
rect -30954 3795 -30915 3822
rect -30881 3795 -30842 3822
rect -30808 3795 -30768 3822
rect -30734 3795 -30694 3822
rect -30660 3795 -30620 3822
rect -30586 3795 -30546 3822
rect -30512 3795 -30472 3822
rect -30438 3795 -30398 3822
rect -30364 3795 -30324 3822
rect -30290 3795 -30250 3822
rect -30216 3795 -30176 3822
rect -30142 3795 -30102 3822
rect -30068 3795 -30028 3822
rect -29994 3795 -29954 3822
rect -29920 3795 -29880 3822
rect -29846 3795 -29806 3822
rect -29772 3795 -29732 3822
rect -29698 3795 -29658 3822
rect -29624 3795 -29584 3822
rect -29550 3795 -29510 3822
rect -29476 3795 -29436 3822
rect -29402 3795 -29362 3822
rect -29328 3795 -29288 3822
rect -29254 3795 -29214 3822
rect -29180 3795 -29134 3822
rect -31669 3788 -29134 3795
rect -29100 3792 -29046 3822
rect -29012 3792 -28958 3822
rect -28924 3792 -28870 3822
rect -28836 3801 -27036 3822
rect -28836 3792 -28189 3801
rect -28155 3792 -28115 3801
rect -28081 3792 -28041 3801
rect -28007 3792 -27967 3801
rect -27933 3792 -27893 3801
rect -27859 3792 -27819 3801
rect -27785 3792 -27745 3801
rect -27711 3792 -27671 3801
rect -27637 3792 -27597 3801
rect -27563 3792 -27523 3801
rect -27489 3792 -27449 3801
rect -27415 3792 -27375 3801
rect -27341 3792 -27301 3801
rect -27267 3792 -27227 3801
rect -27193 3792 -27153 3801
rect -27119 3792 -27036 3801
rect -29100 3788 -29078 3792
rect -29012 3788 -29010 3792
rect -32352 3748 -32315 3787
rect -31669 3786 -29078 3788
rect -31669 3757 -31632 3786
rect -31598 3757 -31563 3786
rect -31529 3757 -31494 3786
rect -31460 3757 -31425 3786
rect -32352 3714 -32344 3748
rect -31669 3723 -31645 3757
rect -31598 3752 -31572 3757
rect -31529 3752 -31499 3757
rect -31460 3752 -31426 3757
rect -31391 3752 -31356 3786
rect -31322 3757 -31287 3786
rect -31253 3757 -31218 3786
rect -31184 3757 -31149 3786
rect -31115 3757 -31080 3786
rect -31046 3757 -31011 3786
rect -30977 3757 -30942 3786
rect -30908 3757 -30873 3786
rect -30839 3757 -30804 3786
rect -31319 3752 -31287 3757
rect -31246 3752 -31218 3757
rect -31173 3752 -31149 3757
rect -31100 3752 -31080 3757
rect -31027 3752 -31011 3757
rect -30954 3752 -30942 3757
rect -30881 3752 -30873 3757
rect -30808 3752 -30804 3757
rect -30770 3757 -30735 3786
rect -30701 3757 -30666 3786
rect -30632 3757 -30597 3786
rect -30563 3757 -30528 3786
rect -30494 3757 -30459 3786
rect -30425 3757 -30390 3786
rect -30356 3757 -30321 3786
rect -30770 3752 -30768 3757
rect -30701 3752 -30694 3757
rect -30632 3752 -30620 3757
rect -30563 3752 -30546 3757
rect -30494 3752 -30472 3757
rect -30425 3752 -30398 3757
rect -30356 3752 -30324 3757
rect -30287 3752 -30252 3786
rect -30218 3757 -30183 3786
rect -30149 3757 -30114 3786
rect -30080 3757 -30045 3786
rect -30011 3757 -29976 3786
rect -29942 3757 -29907 3786
rect -29873 3757 -29838 3786
rect -29804 3757 -29769 3786
rect -30216 3752 -30183 3757
rect -30142 3752 -30114 3757
rect -30068 3752 -30045 3757
rect -29994 3752 -29976 3757
rect -29920 3752 -29907 3757
rect -29846 3752 -29838 3757
rect -29772 3752 -29769 3757
rect -29735 3757 -29700 3786
rect -29666 3757 -29631 3786
rect -29597 3757 -29562 3786
rect -29528 3757 -29493 3786
rect -29459 3757 -29424 3786
rect -29390 3757 -29355 3786
rect -29321 3757 -29286 3786
rect -29735 3752 -29732 3757
rect -29666 3752 -29658 3757
rect -29597 3752 -29584 3757
rect -29528 3752 -29510 3757
rect -29459 3752 -29436 3757
rect -29390 3752 -29362 3757
rect -29321 3752 -29288 3757
rect -29252 3752 -29217 3786
rect -29183 3757 -29148 3786
rect -29180 3752 -29148 3757
rect -29114 3758 -29078 3786
rect -29044 3758 -29010 3788
rect -28976 3788 -28958 3792
rect -28976 3758 -28942 3788
rect -28908 3758 -28874 3792
rect -28836 3788 -28806 3792
rect -28840 3758 -28806 3788
rect -28772 3758 -28738 3792
rect -28704 3758 -28670 3792
rect -28636 3758 -28602 3792
rect -28568 3758 -28534 3792
rect -28500 3758 -28466 3792
rect -28432 3758 -28398 3792
rect -28364 3758 -28330 3792
rect -28296 3758 -28262 3792
rect -28228 3758 -28194 3792
rect -28155 3767 -28126 3792
rect -28081 3767 -28058 3792
rect -28007 3767 -27990 3792
rect -27933 3767 -27922 3792
rect -27859 3767 -27854 3792
rect -28160 3758 -28126 3767
rect -28092 3758 -28058 3767
rect -28024 3758 -27990 3767
rect -27956 3758 -27922 3767
rect -27888 3758 -27854 3767
rect -27820 3767 -27819 3792
rect -27752 3767 -27745 3792
rect -27684 3767 -27671 3792
rect -27616 3767 -27597 3792
rect -27548 3767 -27523 3792
rect -27480 3767 -27449 3792
rect -27820 3758 -27786 3767
rect -27752 3758 -27718 3767
rect -27684 3758 -27650 3767
rect -27616 3758 -27582 3767
rect -27548 3758 -27514 3767
rect -27480 3758 -27446 3767
rect -27412 3758 -27378 3792
rect -27341 3767 -27310 3792
rect -27267 3767 -27242 3792
rect -27193 3767 -27174 3792
rect -27119 3767 -27106 3792
rect -27344 3758 -27310 3767
rect -27276 3758 -27242 3767
rect -27208 3758 -27174 3767
rect -27140 3758 -27106 3767
rect -27072 3758 -27036 3792
rect -29114 3752 -27036 3758
rect -31611 3723 -31572 3752
rect -31538 3723 -31499 3752
rect -31465 3723 -31426 3752
rect -31392 3723 -31353 3752
rect -31319 3723 -31280 3752
rect -31246 3723 -31207 3752
rect -31173 3723 -31134 3752
rect -31100 3723 -31061 3752
rect -31027 3723 -30988 3752
rect -30954 3723 -30915 3752
rect -30881 3723 -30842 3752
rect -30808 3723 -30768 3752
rect -30734 3723 -30694 3752
rect -30660 3723 -30620 3752
rect -30586 3723 -30546 3752
rect -30512 3723 -30472 3752
rect -30438 3723 -30398 3752
rect -30364 3723 -30324 3752
rect -30290 3723 -30250 3752
rect -30216 3723 -30176 3752
rect -30142 3723 -30102 3752
rect -30068 3723 -30028 3752
rect -29994 3723 -29954 3752
rect -29920 3723 -29880 3752
rect -29846 3723 -29806 3752
rect -29772 3723 -29732 3752
rect -29698 3723 -29658 3752
rect -29624 3723 -29584 3752
rect -29550 3723 -29510 3752
rect -29476 3723 -29436 3752
rect -29402 3723 -29362 3752
rect -29328 3723 -29288 3752
rect -29254 3723 -29214 3752
rect -29180 3749 -27036 3752
rect -29180 3723 -29134 3749
rect -31669 3716 -29134 3723
rect -29100 3723 -29046 3749
rect -29012 3723 -28958 3749
rect -28924 3723 -28870 3749
rect -28836 3728 -27036 3749
rect -28836 3723 -28189 3728
rect -28155 3723 -28115 3728
rect -28081 3723 -28041 3728
rect -28007 3723 -27967 3728
rect -27933 3723 -27893 3728
rect -27859 3723 -27819 3728
rect -27785 3723 -27745 3728
rect -27711 3723 -27671 3728
rect -27637 3723 -27597 3728
rect -27563 3723 -27523 3728
rect -27489 3723 -27449 3728
rect -27415 3723 -27375 3728
rect -27341 3723 -27301 3728
rect -27267 3723 -27227 3728
rect -27193 3723 -27153 3728
rect -27119 3723 -27036 3728
rect -32352 3675 -32315 3714
rect -31669 3685 -31632 3716
rect -31598 3685 -31563 3716
rect -31529 3685 -31494 3716
rect -31460 3685 -31425 3716
rect -32352 3641 -32344 3675
rect -31669 3651 -31645 3685
rect -31598 3682 -31572 3685
rect -31529 3682 -31499 3685
rect -31460 3682 -31426 3685
rect -31391 3682 -31356 3716
rect -31322 3685 -31287 3716
rect -31253 3685 -31218 3716
rect -31184 3685 -31149 3716
rect -31115 3685 -31080 3716
rect -31046 3685 -31011 3716
rect -30977 3685 -30942 3716
rect -30908 3685 -30873 3716
rect -30839 3685 -30804 3716
rect -31319 3682 -31287 3685
rect -31246 3682 -31218 3685
rect -31173 3682 -31149 3685
rect -31100 3682 -31080 3685
rect -31027 3682 -31011 3685
rect -30954 3682 -30942 3685
rect -30881 3682 -30873 3685
rect -30808 3682 -30804 3685
rect -30770 3685 -30735 3716
rect -30701 3685 -30666 3716
rect -30632 3685 -30597 3716
rect -30563 3685 -30528 3716
rect -30494 3685 -30459 3716
rect -30425 3685 -30390 3716
rect -30356 3685 -30321 3716
rect -30770 3682 -30768 3685
rect -30701 3682 -30694 3685
rect -30632 3682 -30620 3685
rect -30563 3682 -30546 3685
rect -30494 3682 -30472 3685
rect -30425 3682 -30398 3685
rect -30356 3682 -30324 3685
rect -30287 3682 -30252 3716
rect -30218 3685 -30183 3716
rect -30149 3685 -30114 3716
rect -30080 3685 -30045 3716
rect -30011 3685 -29976 3716
rect -29942 3685 -29907 3716
rect -29873 3685 -29838 3716
rect -29804 3685 -29769 3716
rect -30216 3682 -30183 3685
rect -30142 3682 -30114 3685
rect -30068 3682 -30045 3685
rect -29994 3682 -29976 3685
rect -29920 3682 -29907 3685
rect -29846 3682 -29838 3685
rect -29772 3682 -29769 3685
rect -29735 3685 -29700 3716
rect -29666 3685 -29631 3716
rect -29597 3685 -29562 3716
rect -29528 3685 -29493 3716
rect -29459 3685 -29424 3716
rect -29390 3685 -29355 3716
rect -29321 3685 -29286 3716
rect -29735 3682 -29732 3685
rect -29666 3682 -29658 3685
rect -29597 3682 -29584 3685
rect -29528 3682 -29510 3685
rect -29459 3682 -29436 3685
rect -29390 3682 -29362 3685
rect -29321 3682 -29288 3685
rect -29252 3682 -29217 3716
rect -29183 3685 -29148 3716
rect -29100 3715 -29078 3723
rect -29012 3715 -29010 3723
rect -29180 3682 -29148 3685
rect -29114 3689 -29078 3715
rect -29044 3689 -29010 3715
rect -28976 3715 -28958 3723
rect -28976 3689 -28942 3715
rect -28908 3689 -28874 3723
rect -28836 3715 -28806 3723
rect -28840 3689 -28806 3715
rect -28772 3689 -28738 3723
rect -28704 3689 -28670 3723
rect -28636 3689 -28602 3723
rect -28568 3689 -28534 3723
rect -28500 3689 -28466 3723
rect -28432 3689 -28398 3723
rect -28364 3689 -28330 3723
rect -28296 3689 -28262 3723
rect -28228 3689 -28194 3723
rect -28155 3694 -28126 3723
rect -28081 3694 -28058 3723
rect -28007 3694 -27990 3723
rect -27933 3694 -27922 3723
rect -27859 3694 -27854 3723
rect -28160 3689 -28126 3694
rect -28092 3689 -28058 3694
rect -28024 3689 -27990 3694
rect -27956 3689 -27922 3694
rect -27888 3689 -27854 3694
rect -27820 3694 -27819 3723
rect -27752 3694 -27745 3723
rect -27684 3694 -27671 3723
rect -27616 3694 -27597 3723
rect -27548 3694 -27523 3723
rect -27480 3694 -27449 3723
rect -27820 3689 -27786 3694
rect -27752 3689 -27718 3694
rect -27684 3689 -27650 3694
rect -27616 3689 -27582 3694
rect -27548 3689 -27514 3694
rect -27480 3689 -27446 3694
rect -27412 3689 -27378 3723
rect -27341 3694 -27310 3723
rect -27267 3694 -27242 3723
rect -27193 3694 -27174 3723
rect -27119 3694 -27106 3723
rect -27344 3689 -27310 3694
rect -27276 3689 -27242 3694
rect -27208 3689 -27174 3694
rect -27140 3689 -27106 3694
rect -27072 3689 -27036 3723
rect -29114 3682 -27036 3689
rect 3938 3806 4010 3840
rect 4044 3806 4082 3840
rect 4140 3806 4154 3840
rect 4208 3806 4226 3840
rect 4276 3806 4298 3840
rect 4344 3806 4370 3840
rect 4412 3806 4442 3840
rect 4480 3806 4514 3840
rect 4548 3806 4582 3840
rect 4620 3806 4650 3840
rect 4692 3806 4718 3840
rect 4764 3806 4786 3840
rect 4836 3806 4854 3840
rect 4908 3806 4922 3840
rect 4980 3806 4990 3840
rect 5052 3806 5058 3840
rect 5124 3806 5126 3840
rect 5160 3806 5162 3840
rect 5228 3806 5234 3840
rect 5296 3806 5306 3840
rect 5364 3806 5378 3840
rect 5432 3806 5450 3840
rect 5500 3806 5522 3840
rect 5568 3806 5594 3840
rect 5636 3806 5666 3840
rect 5704 3806 5772 3840
rect 3938 3768 3972 3806
rect 4722 3772 4942 3806
rect 4722 3753 4723 3772
rect 4757 3753 4815 3772
rect 4849 3753 4907 3772
rect 3938 3692 3972 3700
rect -31611 3651 -31572 3682
rect -31538 3651 -31499 3682
rect -31465 3651 -31426 3682
rect -31392 3651 -31353 3682
rect -31319 3651 -31280 3682
rect -31246 3651 -31207 3682
rect -31173 3651 -31134 3682
rect -31100 3651 -31061 3682
rect -31027 3651 -30988 3682
rect -30954 3651 -30915 3682
rect -30881 3651 -30842 3682
rect -30808 3651 -30768 3682
rect -30734 3651 -30694 3682
rect -30660 3651 -30620 3682
rect -30586 3651 -30546 3682
rect -30512 3651 -30472 3682
rect -30438 3651 -30398 3682
rect -30364 3651 -30324 3682
rect -30290 3651 -30250 3682
rect -30216 3651 -30176 3682
rect -30142 3651 -30102 3682
rect -30068 3651 -30028 3682
rect -29994 3651 -29954 3682
rect -29920 3651 -29880 3682
rect -29846 3651 -29806 3682
rect -29772 3651 -29732 3682
rect -29698 3651 -29658 3682
rect -29624 3651 -29584 3682
rect -29550 3651 -29510 3682
rect -29476 3651 -29436 3682
rect -29402 3651 -29362 3682
rect -29328 3651 -29288 3682
rect -29254 3651 -29214 3682
rect -29180 3676 -27036 3682
rect -29180 3651 -29134 3676
rect -31669 3646 -29134 3651
rect -29100 3654 -29046 3676
rect -29012 3654 -28958 3676
rect -28924 3654 -28870 3676
rect -28836 3655 -27036 3676
rect -28836 3654 -28189 3655
rect -28155 3654 -28115 3655
rect -28081 3654 -28041 3655
rect -28007 3654 -27967 3655
rect -27933 3654 -27893 3655
rect -27859 3654 -27819 3655
rect -27785 3654 -27745 3655
rect -27711 3654 -27671 3655
rect -27637 3654 -27597 3655
rect -27563 3654 -27523 3655
rect -27489 3654 -27449 3655
rect -27415 3654 -27375 3655
rect -27341 3654 -27301 3655
rect -27267 3654 -27227 3655
rect -27193 3654 -27153 3655
rect -27119 3654 -27036 3655
rect -699 3654 -677 3688
rect -628 3654 -597 3688
rect -557 3654 -519 3688
rect -482 3654 -447 3688
rect -401 3654 -389 3688
rect 157 3654 171 3688
rect 215 3654 244 3688
rect 284 3654 317 3688
rect 353 3654 388 3688
rect 424 3654 457 3688
rect 497 3654 526 3688
rect 570 3654 595 3688
rect 643 3654 664 3688
rect 716 3654 733 3688
rect 789 3654 802 3688
rect 862 3654 871 3688
rect 935 3654 940 3688
rect 1008 3654 1009 3688
rect 1043 3654 1047 3688
rect 1112 3654 1120 3688
rect 1181 3654 1193 3688
rect 1250 3654 1266 3688
rect 1319 3654 1339 3688
rect 1388 3654 1412 3688
rect 1457 3654 1485 3688
rect 1526 3654 1558 3688
rect 1595 3654 1630 3688
rect 1665 3654 1699 3688
rect 1738 3654 1768 3688
rect 1811 3654 1837 3688
rect 1884 3654 1906 3688
rect 1957 3654 1975 3688
rect 2029 3654 2044 3688
rect 2101 3654 2113 3688
rect 2173 3654 2182 3688
rect 2245 3654 2251 3688
rect 2317 3654 2320 3688
rect 2354 3654 2355 3688
rect 2423 3654 2427 3688
rect 2492 3654 2499 3688
rect 2561 3654 2571 3688
rect 2630 3654 2643 3688
rect 2699 3654 2715 3688
rect 2768 3654 2787 3688
rect 2837 3654 2859 3688
rect 2906 3654 2931 3688
rect 2975 3654 3003 3688
rect 3044 3654 3075 3688
rect 3112 3654 3146 3688
rect 3181 3654 3214 3688
rect 3253 3654 3282 3688
rect 3325 3654 3350 3688
rect 3397 3654 3418 3688
rect 3469 3654 3486 3688
rect 3541 3654 3544 3688
rect -32352 3602 -32315 3641
rect -31669 3613 -31632 3646
rect -31598 3613 -31563 3646
rect -31529 3613 -31494 3646
rect -31460 3613 -31425 3646
rect -32352 3568 -32344 3602
rect -31669 3579 -31645 3613
rect -31598 3612 -31572 3613
rect -31529 3612 -31499 3613
rect -31460 3612 -31426 3613
rect -31391 3612 -31356 3646
rect -31322 3613 -31287 3646
rect -31253 3613 -31218 3646
rect -31184 3613 -31149 3646
rect -31115 3613 -31080 3646
rect -31046 3613 -31011 3646
rect -30977 3613 -30942 3646
rect -30908 3613 -30873 3646
rect -30839 3613 -30804 3646
rect -31319 3612 -31287 3613
rect -31246 3612 -31218 3613
rect -31173 3612 -31149 3613
rect -31100 3612 -31080 3613
rect -31027 3612 -31011 3613
rect -30954 3612 -30942 3613
rect -30881 3612 -30873 3613
rect -30808 3612 -30804 3613
rect -30770 3613 -30735 3646
rect -30701 3613 -30666 3646
rect -30632 3613 -30597 3646
rect -30563 3613 -30528 3646
rect -30494 3613 -30459 3646
rect -30425 3613 -30390 3646
rect -30356 3613 -30321 3646
rect -30770 3612 -30768 3613
rect -30701 3612 -30694 3613
rect -30632 3612 -30620 3613
rect -30563 3612 -30546 3613
rect -30494 3612 -30472 3613
rect -30425 3612 -30398 3613
rect -30356 3612 -30324 3613
rect -30287 3612 -30252 3646
rect -30218 3613 -30183 3646
rect -30149 3613 -30114 3646
rect -30080 3613 -30045 3646
rect -30011 3613 -29976 3646
rect -29942 3613 -29907 3646
rect -29873 3613 -29838 3646
rect -29804 3613 -29769 3646
rect -30216 3612 -30183 3613
rect -30142 3612 -30114 3613
rect -30068 3612 -30045 3613
rect -29994 3612 -29976 3613
rect -29920 3612 -29907 3613
rect -29846 3612 -29838 3613
rect -29772 3612 -29769 3613
rect -29735 3613 -29700 3646
rect -29666 3613 -29631 3646
rect -29597 3613 -29562 3646
rect -29528 3613 -29493 3646
rect -29459 3613 -29424 3646
rect -29390 3613 -29355 3646
rect -29321 3613 -29286 3646
rect -29735 3612 -29732 3613
rect -29666 3612 -29658 3613
rect -29597 3612 -29584 3613
rect -29528 3612 -29510 3613
rect -29459 3612 -29436 3613
rect -29390 3612 -29362 3613
rect -29321 3612 -29288 3613
rect -29252 3612 -29217 3646
rect -29183 3613 -29148 3646
rect -29100 3642 -29078 3654
rect -29012 3642 -29010 3654
rect -29180 3612 -29148 3613
rect -29114 3620 -29078 3642
rect -29044 3620 -29010 3642
rect -28976 3642 -28958 3654
rect -28976 3620 -28942 3642
rect -28908 3620 -28874 3654
rect -28836 3642 -28806 3654
rect -28840 3620 -28806 3642
rect -28772 3620 -28738 3654
rect -28704 3620 -28670 3654
rect -28636 3620 -28602 3654
rect -28568 3620 -28534 3654
rect -28500 3620 -28466 3654
rect -28432 3620 -28398 3654
rect -28364 3620 -28330 3654
rect -28296 3620 -28262 3654
rect -28228 3620 -28194 3654
rect -28155 3621 -28126 3654
rect -28081 3621 -28058 3654
rect -28007 3621 -27990 3654
rect -27933 3621 -27922 3654
rect -27859 3621 -27854 3654
rect -28160 3620 -28126 3621
rect -28092 3620 -28058 3621
rect -28024 3620 -27990 3621
rect -27956 3620 -27922 3621
rect -27888 3620 -27854 3621
rect -27820 3621 -27819 3654
rect -27752 3621 -27745 3654
rect -27684 3621 -27671 3654
rect -27616 3621 -27597 3654
rect -27548 3621 -27523 3654
rect -27480 3621 -27449 3654
rect -27820 3620 -27786 3621
rect -27752 3620 -27718 3621
rect -27684 3620 -27650 3621
rect -27616 3620 -27582 3621
rect -27548 3620 -27514 3621
rect -27480 3620 -27446 3621
rect -27412 3620 -27378 3654
rect -27341 3621 -27310 3654
rect -27267 3621 -27242 3654
rect -27193 3621 -27174 3654
rect -27119 3621 -27106 3654
rect -27344 3620 -27310 3621
rect -27276 3620 -27242 3621
rect -27208 3620 -27174 3621
rect -27140 3620 -27106 3621
rect -27072 3620 -27036 3654
rect -29114 3612 -27036 3620
rect -31611 3579 -31572 3612
rect -31538 3579 -31499 3612
rect -31465 3579 -31426 3612
rect -31392 3579 -31353 3612
rect -31319 3579 -31280 3612
rect -31246 3579 -31207 3612
rect -31173 3579 -31134 3612
rect -31100 3579 -31061 3612
rect -31027 3579 -30988 3612
rect -30954 3579 -30915 3612
rect -30881 3579 -30842 3612
rect -30808 3579 -30768 3612
rect -30734 3579 -30694 3612
rect -30660 3579 -30620 3612
rect -30586 3579 -30546 3612
rect -30512 3579 -30472 3612
rect -30438 3579 -30398 3612
rect -30364 3579 -30324 3612
rect -30290 3579 -30250 3612
rect -30216 3579 -30176 3612
rect -30142 3579 -30102 3612
rect -30068 3579 -30028 3612
rect -29994 3579 -29954 3612
rect -29920 3579 -29880 3612
rect -29846 3579 -29806 3612
rect -29772 3579 -29732 3612
rect -29698 3579 -29658 3612
rect -29624 3579 -29584 3612
rect -29550 3579 -29510 3612
rect -29476 3579 -29436 3612
rect -29402 3579 -29362 3612
rect -29328 3579 -29288 3612
rect -29254 3579 -29214 3612
rect -29180 3603 -27036 3612
rect -29180 3579 -29134 3603
rect -31669 3576 -29134 3579
rect -29100 3585 -29046 3603
rect -29012 3585 -28958 3603
rect -28924 3585 -28870 3603
rect -28836 3585 -27036 3603
rect -32352 3529 -32315 3568
rect -31669 3542 -31632 3576
rect -31598 3542 -31563 3576
rect -31529 3542 -31494 3576
rect -31460 3542 -31425 3576
rect -31391 3542 -31356 3576
rect -31322 3542 -31287 3576
rect -31253 3542 -31218 3576
rect -31184 3542 -31149 3576
rect -31115 3542 -31080 3576
rect -31046 3542 -31011 3576
rect -30977 3542 -30942 3576
rect -30908 3542 -30873 3576
rect -30839 3542 -30804 3576
rect -30770 3542 -30735 3576
rect -30701 3542 -30666 3576
rect -30632 3542 -30597 3576
rect -30563 3542 -30528 3576
rect -30494 3542 -30459 3576
rect -30425 3542 -30390 3576
rect -30356 3542 -30321 3576
rect -30287 3542 -30252 3576
rect -30218 3542 -30183 3576
rect -30149 3542 -30114 3576
rect -30080 3542 -30045 3576
rect -30011 3542 -29976 3576
rect -29942 3542 -29907 3576
rect -29873 3542 -29838 3576
rect -29804 3542 -29769 3576
rect -29735 3542 -29700 3576
rect -29666 3542 -29631 3576
rect -29597 3542 -29562 3576
rect -29528 3542 -29493 3576
rect -29459 3542 -29424 3576
rect -29390 3542 -29355 3576
rect -29321 3542 -29286 3576
rect -29252 3542 -29217 3576
rect -29183 3542 -29148 3576
rect -29100 3569 -29078 3585
rect -29012 3569 -29010 3585
rect -29114 3551 -29078 3569
rect -29044 3551 -29010 3569
rect -28976 3569 -28958 3585
rect -28976 3551 -28942 3569
rect -28908 3551 -28874 3585
rect -28836 3569 -28806 3585
rect -28840 3551 -28806 3569
rect -28772 3551 -28738 3585
rect -28704 3551 -28670 3585
rect -28636 3551 -28602 3585
rect -28568 3551 -28534 3585
rect -28500 3551 -28466 3585
rect -28432 3551 -28398 3585
rect -28364 3551 -28330 3585
rect -28296 3551 -28262 3585
rect -28228 3551 -28194 3585
rect -28160 3582 -28126 3585
rect -28092 3582 -28058 3585
rect -28024 3582 -27990 3585
rect -27956 3582 -27922 3585
rect -27888 3582 -27854 3585
rect -28155 3551 -28126 3582
rect -28081 3551 -28058 3582
rect -28007 3551 -27990 3582
rect -27933 3551 -27922 3582
rect -27859 3551 -27854 3582
rect -27820 3582 -27786 3585
rect -27752 3582 -27718 3585
rect -27684 3582 -27650 3585
rect -27616 3582 -27582 3585
rect -27548 3582 -27514 3585
rect -27480 3582 -27446 3585
rect -27820 3551 -27819 3582
rect -27752 3551 -27745 3582
rect -27684 3551 -27671 3582
rect -27616 3551 -27597 3582
rect -27548 3551 -27523 3582
rect -27480 3551 -27449 3582
rect -27412 3551 -27378 3585
rect -27344 3582 -27310 3585
rect -27276 3582 -27242 3585
rect -27208 3582 -27174 3585
rect -27140 3582 -27106 3585
rect -27341 3551 -27310 3582
rect -27267 3551 -27242 3582
rect -27193 3551 -27174 3582
rect -27119 3551 -27106 3582
rect -27072 3551 -27036 3585
rect 4757 3738 4802 3753
rect 4849 3738 4886 3753
rect 4941 3738 4942 3772
rect 4752 3719 4802 3738
rect 4836 3719 4886 3738
rect 4920 3719 4942 3738
rect 4718 3703 4942 3719
rect 4718 3678 4723 3703
rect 4757 3678 4815 3703
rect 4849 3678 4907 3703
rect 4757 3669 4802 3678
rect 4849 3669 4886 3678
rect 4941 3669 4942 3703
rect 3938 3616 3972 3632
rect -29114 3548 -28189 3551
rect -28155 3548 -28115 3551
rect -28081 3548 -28041 3551
rect -28007 3548 -27967 3551
rect -27933 3548 -27893 3551
rect -27859 3548 -27819 3551
rect -27785 3548 -27745 3551
rect -27711 3548 -27671 3551
rect -27637 3548 -27597 3551
rect -27563 3548 -27523 3551
rect -27489 3548 -27449 3551
rect -27415 3548 -27375 3551
rect -27341 3548 -27301 3551
rect -27267 3548 -27227 3551
rect -27193 3548 -27153 3551
rect -27119 3548 -27036 3551
rect -29114 3542 -27036 3548
rect -31669 3541 -27036 3542
rect -32352 3495 -32344 3529
rect -31669 3507 -31645 3541
rect -31611 3507 -31572 3541
rect -31538 3507 -31499 3541
rect -31465 3507 -31426 3541
rect -31392 3507 -31353 3541
rect -31319 3507 -31280 3541
rect -31246 3507 -31207 3541
rect -31173 3507 -31134 3541
rect -31100 3507 -31061 3541
rect -31027 3507 -30988 3541
rect -30954 3507 -30915 3541
rect -30881 3507 -30842 3541
rect -30808 3507 -30768 3541
rect -30734 3507 -30694 3541
rect -30660 3507 -30620 3541
rect -30586 3507 -30546 3541
rect -30512 3507 -30472 3541
rect -30438 3507 -30398 3541
rect -30364 3507 -30324 3541
rect -30290 3507 -30250 3541
rect -30216 3507 -30176 3541
rect -30142 3507 -30102 3541
rect -30068 3507 -30028 3541
rect -29994 3507 -29954 3541
rect -29920 3507 -29880 3541
rect -29846 3507 -29806 3541
rect -29772 3507 -29732 3541
rect -29698 3507 -29658 3541
rect -29624 3507 -29584 3541
rect -29550 3507 -29510 3541
rect -29476 3507 -29436 3541
rect -29402 3507 -29362 3541
rect -29328 3507 -29288 3541
rect -29254 3507 -29214 3541
rect -29180 3530 -27036 3541
rect -29180 3507 -29134 3530
rect -31669 3506 -29134 3507
rect -29100 3516 -29046 3530
rect -29012 3516 -28958 3530
rect -28924 3516 -28870 3530
rect -28836 3516 -27036 3530
rect -32352 3456 -32315 3495
rect -31669 3472 -31632 3506
rect -31598 3472 -31563 3506
rect -31529 3472 -31494 3506
rect -31460 3472 -31425 3506
rect -31391 3472 -31356 3506
rect -31322 3472 -31287 3506
rect -31253 3472 -31218 3506
rect -31184 3472 -31149 3506
rect -31115 3472 -31080 3506
rect -31046 3472 -31011 3506
rect -30977 3472 -30942 3506
rect -30908 3472 -30873 3506
rect -30839 3472 -30804 3506
rect -30770 3472 -30735 3506
rect -30701 3472 -30666 3506
rect -30632 3472 -30597 3506
rect -30563 3472 -30528 3506
rect -30494 3472 -30459 3506
rect -30425 3472 -30390 3506
rect -30356 3472 -30321 3506
rect -30287 3472 -30252 3506
rect -30218 3472 -30183 3506
rect -30149 3472 -30114 3506
rect -30080 3472 -30045 3506
rect -30011 3472 -29976 3506
rect -29942 3472 -29907 3506
rect -29873 3472 -29838 3506
rect -29804 3472 -29769 3506
rect -29735 3472 -29700 3506
rect -29666 3472 -29631 3506
rect -29597 3472 -29562 3506
rect -29528 3472 -29493 3506
rect -29459 3472 -29424 3506
rect -29390 3472 -29355 3506
rect -29321 3472 -29286 3506
rect -29252 3472 -29217 3506
rect -29183 3472 -29148 3506
rect -29100 3496 -29078 3516
rect -29012 3496 -29010 3516
rect -29114 3482 -29078 3496
rect -29044 3482 -29010 3496
rect -28976 3496 -28958 3516
rect -28976 3482 -28942 3496
rect -28908 3482 -28874 3516
rect -28836 3496 -28806 3516
rect -28840 3482 -28806 3496
rect -28772 3482 -28738 3516
rect -28704 3482 -28670 3516
rect -28636 3482 -28602 3516
rect -28568 3482 -28534 3516
rect -28500 3482 -28466 3516
rect -28432 3482 -28398 3516
rect -28364 3482 -28330 3516
rect -28296 3482 -28262 3516
rect -28228 3482 -28194 3516
rect -28160 3509 -28126 3516
rect -28092 3509 -28058 3516
rect -28024 3509 -27990 3516
rect -27956 3509 -27922 3516
rect -27888 3509 -27854 3516
rect -28155 3482 -28126 3509
rect -28081 3482 -28058 3509
rect -28007 3482 -27990 3509
rect -27933 3482 -27922 3509
rect -27859 3482 -27854 3509
rect -27820 3509 -27786 3516
rect -27752 3509 -27718 3516
rect -27684 3509 -27650 3516
rect -27616 3509 -27582 3516
rect -27548 3509 -27514 3516
rect -27480 3509 -27446 3516
rect -27820 3482 -27819 3509
rect -27752 3482 -27745 3509
rect -27684 3482 -27671 3509
rect -27616 3482 -27597 3509
rect -27548 3482 -27523 3509
rect -27480 3482 -27449 3509
rect -27412 3482 -27378 3516
rect -27344 3509 -27310 3516
rect -27276 3509 -27242 3516
rect -27208 3509 -27174 3516
rect -27140 3509 -27106 3516
rect -27341 3482 -27310 3509
rect -27267 3482 -27242 3509
rect -27193 3482 -27174 3509
rect -27119 3482 -27106 3509
rect -27072 3482 -27036 3516
rect -29114 3475 -28189 3482
rect -28155 3475 -28115 3482
rect -28081 3475 -28041 3482
rect -28007 3475 -27967 3482
rect -27933 3475 -27893 3482
rect -27859 3475 -27819 3482
rect -27785 3475 -27745 3482
rect -27711 3475 -27671 3482
rect -27637 3475 -27597 3482
rect -27563 3475 -27523 3482
rect -27489 3475 -27449 3482
rect -27415 3475 -27375 3482
rect -27341 3475 -27301 3482
rect -27267 3475 -27227 3482
rect -27193 3475 -27153 3482
rect -27119 3475 -27036 3482
rect -29114 3472 -27036 3475
rect -31669 3469 -27036 3472
rect -32352 3422 -32344 3456
rect -31669 3435 -31645 3469
rect -31611 3436 -31572 3469
rect -31538 3436 -31499 3469
rect -31465 3436 -31426 3469
rect -31392 3436 -31353 3469
rect -31319 3436 -31280 3469
rect -31246 3436 -31207 3469
rect -31173 3436 -31134 3469
rect -31100 3436 -31061 3469
rect -31027 3436 -30988 3469
rect -30954 3436 -30915 3469
rect -30881 3436 -30842 3469
rect -30808 3436 -30768 3469
rect -30734 3436 -30694 3469
rect -30660 3436 -30620 3469
rect -30586 3436 -30546 3469
rect -30512 3436 -30472 3469
rect -30438 3436 -30398 3469
rect -30364 3436 -30324 3469
rect -30290 3436 -30250 3469
rect -30216 3436 -30176 3469
rect -30142 3436 -30102 3469
rect -30068 3436 -30028 3469
rect -29994 3436 -29954 3469
rect -29920 3436 -29880 3469
rect -29846 3436 -29806 3469
rect -29772 3436 -29732 3469
rect -29698 3436 -29658 3469
rect -29624 3436 -29584 3469
rect -29550 3436 -29510 3469
rect -29476 3436 -29436 3469
rect -29402 3436 -29362 3469
rect -29328 3436 -29288 3469
rect -29254 3436 -29214 3469
rect -29180 3457 -27036 3469
rect -29180 3436 -29134 3457
rect -29100 3447 -29046 3457
rect -29012 3447 -28958 3457
rect -28924 3447 -28870 3457
rect -28836 3447 -27036 3457
rect -31598 3435 -31572 3436
rect -31529 3435 -31499 3436
rect -31460 3435 -31426 3436
rect -32352 3383 -32315 3422
rect -31669 3402 -31632 3435
rect -31598 3402 -31563 3435
rect -31529 3402 -31494 3435
rect -31460 3402 -31425 3435
rect -31391 3402 -31356 3436
rect -31319 3435 -31287 3436
rect -31246 3435 -31218 3436
rect -31173 3435 -31149 3436
rect -31100 3435 -31080 3436
rect -31027 3435 -31011 3436
rect -30954 3435 -30942 3436
rect -30881 3435 -30873 3436
rect -30808 3435 -30804 3436
rect -31322 3402 -31287 3435
rect -31253 3402 -31218 3435
rect -31184 3402 -31149 3435
rect -31115 3402 -31080 3435
rect -31046 3402 -31011 3435
rect -30977 3402 -30942 3435
rect -30908 3402 -30873 3435
rect -30839 3402 -30804 3435
rect -30770 3435 -30768 3436
rect -30701 3435 -30694 3436
rect -30632 3435 -30620 3436
rect -30563 3435 -30546 3436
rect -30494 3435 -30472 3436
rect -30425 3435 -30398 3436
rect -30356 3435 -30324 3436
rect -30770 3402 -30735 3435
rect -30701 3402 -30666 3435
rect -30632 3402 -30597 3435
rect -30563 3402 -30528 3435
rect -30494 3402 -30459 3435
rect -30425 3402 -30390 3435
rect -30356 3402 -30321 3435
rect -30287 3402 -30252 3436
rect -30216 3435 -30183 3436
rect -30142 3435 -30114 3436
rect -30068 3435 -30045 3436
rect -29994 3435 -29976 3436
rect -29920 3435 -29907 3436
rect -29846 3435 -29838 3436
rect -29772 3435 -29769 3436
rect -30218 3402 -30183 3435
rect -30149 3402 -30114 3435
rect -30080 3402 -30045 3435
rect -30011 3402 -29976 3435
rect -29942 3402 -29907 3435
rect -29873 3402 -29838 3435
rect -29804 3402 -29769 3435
rect -29735 3435 -29732 3436
rect -29666 3435 -29658 3436
rect -29597 3435 -29584 3436
rect -29528 3435 -29510 3436
rect -29459 3435 -29436 3436
rect -29390 3435 -29362 3436
rect -29321 3435 -29288 3436
rect -29735 3402 -29700 3435
rect -29666 3402 -29631 3435
rect -29597 3402 -29562 3435
rect -29528 3402 -29493 3435
rect -29459 3402 -29424 3435
rect -29390 3402 -29355 3435
rect -29321 3402 -29286 3435
rect -29252 3402 -29217 3436
rect -29180 3435 -29148 3436
rect -29183 3402 -29148 3435
rect -29100 3423 -29078 3447
rect -29012 3423 -29010 3447
rect -29114 3413 -29078 3423
rect -29044 3413 -29010 3423
rect -28976 3423 -28958 3447
rect -28976 3413 -28942 3423
rect -28908 3413 -28874 3447
rect -28836 3423 -28806 3447
rect -28840 3413 -28806 3423
rect -28772 3413 -28738 3447
rect -28704 3413 -28670 3447
rect -28636 3413 -28602 3447
rect -28568 3413 -28534 3447
rect -28500 3413 -28466 3447
rect -28432 3413 -28398 3447
rect -28364 3413 -28330 3447
rect -28296 3413 -28262 3447
rect -28228 3413 -28194 3447
rect -28160 3436 -28126 3447
rect -28092 3436 -28058 3447
rect -28024 3436 -27990 3447
rect -27956 3436 -27922 3447
rect -27888 3436 -27854 3447
rect -28155 3413 -28126 3436
rect -28081 3413 -28058 3436
rect -28007 3413 -27990 3436
rect -27933 3413 -27922 3436
rect -27859 3413 -27854 3436
rect -27820 3436 -27786 3447
rect -27752 3436 -27718 3447
rect -27684 3436 -27650 3447
rect -27616 3436 -27582 3447
rect -27548 3436 -27514 3447
rect -27480 3436 -27446 3447
rect -27820 3413 -27819 3436
rect -27752 3413 -27745 3436
rect -27684 3413 -27671 3436
rect -27616 3413 -27597 3436
rect -27548 3413 -27523 3436
rect -27480 3413 -27449 3436
rect -27412 3413 -27378 3447
rect -27344 3436 -27310 3447
rect -27276 3436 -27242 3447
rect -27208 3436 -27174 3447
rect -27140 3436 -27106 3447
rect -27341 3413 -27310 3436
rect -27267 3413 -27242 3436
rect -27193 3413 -27174 3436
rect -27119 3413 -27106 3436
rect -27072 3413 -27036 3447
rect -29114 3402 -28189 3413
rect -28155 3402 -28115 3413
rect -28081 3402 -28041 3413
rect -28007 3402 -27967 3413
rect -27933 3402 -27893 3413
rect -27859 3402 -27819 3413
rect -27785 3402 -27745 3413
rect -27711 3402 -27671 3413
rect -27637 3402 -27597 3413
rect -27563 3402 -27523 3413
rect -27489 3402 -27449 3413
rect -27415 3402 -27375 3413
rect -27341 3402 -27301 3413
rect -27267 3402 -27227 3413
rect -27193 3402 -27153 3413
rect -27119 3402 -27036 3413
rect -31669 3397 -27036 3402
rect -32352 3349 -32344 3383
rect -31669 3363 -31645 3397
rect -31611 3363 -31572 3397
rect -31538 3363 -31499 3397
rect -31465 3363 -31426 3397
rect -31392 3363 -31353 3397
rect -31319 3363 -31280 3397
rect -31246 3363 -31207 3397
rect -31173 3363 -31134 3397
rect -31100 3363 -31061 3397
rect -31027 3363 -30988 3397
rect -30954 3363 -30915 3397
rect -30881 3363 -30842 3397
rect -30808 3363 -30768 3397
rect -30734 3363 -30694 3397
rect -30660 3363 -30620 3397
rect -30586 3363 -30546 3397
rect -30512 3363 -30472 3397
rect -30438 3363 -30398 3397
rect -30364 3363 -30324 3397
rect -30290 3363 -30250 3397
rect -30216 3363 -30176 3397
rect -30142 3363 -30102 3397
rect -30068 3363 -30028 3397
rect -29994 3363 -29954 3397
rect -29920 3363 -29880 3397
rect -29846 3363 -29806 3397
rect -29772 3363 -29732 3397
rect -29698 3363 -29658 3397
rect -29624 3363 -29584 3397
rect -29550 3363 -29510 3397
rect -29476 3363 -29436 3397
rect -29402 3363 -29362 3397
rect -29328 3363 -29288 3397
rect -29254 3363 -29214 3397
rect -29180 3384 -27036 3397
rect -29180 3363 -29134 3384
rect -31669 3350 -29134 3363
rect -29100 3378 -29046 3384
rect -29012 3378 -28958 3384
rect -28924 3378 -28870 3384
rect -28836 3378 -27036 3384
rect -29100 3350 -29078 3378
rect -29012 3350 -29010 3378
rect -32352 3310 -32315 3349
rect -31669 3344 -29078 3350
rect -29044 3344 -29010 3350
rect -28976 3350 -28958 3378
rect -28976 3344 -28942 3350
rect -28908 3344 -28874 3378
rect -28836 3350 -28806 3378
rect -28840 3344 -28806 3350
rect -28772 3344 -28738 3378
rect -28704 3344 -28670 3378
rect -28636 3344 -28602 3378
rect -28568 3344 -28534 3378
rect -28500 3344 -28466 3378
rect -28432 3344 -28398 3378
rect -28364 3344 -28330 3378
rect -28296 3344 -28262 3378
rect -28228 3344 -28194 3378
rect -28160 3363 -28126 3378
rect -28092 3363 -28058 3378
rect -28024 3363 -27990 3378
rect -27956 3363 -27922 3378
rect -27888 3363 -27854 3378
rect -28155 3344 -28126 3363
rect -28081 3344 -28058 3363
rect -28007 3344 -27990 3363
rect -27933 3344 -27922 3363
rect -27859 3344 -27854 3363
rect -27820 3363 -27786 3378
rect -27752 3363 -27718 3378
rect -27684 3363 -27650 3378
rect -27616 3363 -27582 3378
rect -27548 3363 -27514 3378
rect -27480 3363 -27446 3378
rect -27820 3344 -27819 3363
rect -27752 3344 -27745 3363
rect -27684 3344 -27671 3363
rect -27616 3344 -27597 3363
rect -27548 3344 -27523 3363
rect -27480 3344 -27449 3363
rect -27412 3344 -27378 3378
rect -27344 3363 -27310 3378
rect -27276 3363 -27242 3378
rect -27208 3363 -27174 3378
rect -27140 3363 -27106 3378
rect -27341 3344 -27310 3363
rect -27267 3344 -27242 3363
rect -27193 3344 -27174 3363
rect -27119 3344 -27106 3363
rect -27072 3344 -27036 3378
rect -31669 3334 -28189 3344
rect -32352 3276 -32344 3310
rect -31669 3300 -31564 3334
rect -31530 3300 -31496 3334
rect -31462 3300 -31428 3334
rect -31394 3300 -31360 3334
rect -31326 3300 -31292 3334
rect -31258 3300 -31224 3334
rect -31190 3300 -31156 3334
rect -31122 3300 -31088 3334
rect -31054 3300 -31020 3334
rect -30986 3300 -30952 3334
rect -30918 3300 -30884 3334
rect -30850 3300 -30816 3334
rect -30782 3300 -30748 3334
rect -30714 3300 -30680 3334
rect -30646 3300 -30612 3334
rect -30578 3300 -30544 3334
rect -30510 3300 -30476 3334
rect -30442 3300 -30408 3334
rect -30374 3300 -30340 3334
rect -30306 3300 -30272 3334
rect -30238 3300 -30204 3334
rect -30170 3300 -30136 3334
rect -30102 3300 -30068 3334
rect -30034 3300 -30000 3334
rect -29966 3300 -29932 3334
rect -29898 3300 -29864 3334
rect -29830 3300 -29796 3334
rect -29762 3300 -29728 3334
rect -29694 3300 -29660 3334
rect -29626 3300 -29592 3334
rect -29558 3300 -29524 3334
rect -29490 3300 -29456 3334
rect -29422 3300 -29388 3334
rect -29354 3300 -29260 3334
rect -29226 3329 -28189 3334
rect -28155 3329 -28115 3344
rect -28081 3329 -28041 3344
rect -28007 3329 -27967 3344
rect -27933 3329 -27893 3344
rect -27859 3329 -27819 3344
rect -27785 3329 -27745 3344
rect -27711 3329 -27671 3344
rect -27637 3329 -27597 3344
rect -27563 3329 -27523 3344
rect -27489 3329 -27449 3344
rect -27415 3329 -27375 3344
rect -27341 3329 -27301 3344
rect -27267 3329 -27227 3344
rect -27193 3329 -27153 3344
rect -27119 3329 -27036 3344
rect -29226 3311 -27036 3329
rect -29226 3300 -29134 3311
rect -32352 3237 -32315 3276
rect -32352 3203 -32344 3237
rect -31669 3223 -31598 3300
rect -32352 3164 -32315 3203
rect -31669 3189 -31632 3223
rect -32352 3130 -32344 3164
rect -31669 3155 -31598 3189
rect -32352 3091 -32315 3130
rect -31669 3121 -31632 3155
rect -32352 3057 -32344 3091
rect -31669 3087 -31598 3121
rect -32352 3018 -32315 3057
rect -31669 3053 -31632 3087
rect -31669 3019 -31598 3053
rect -32352 2984 -32344 3018
rect -31669 2985 -31632 3019
rect -32352 2945 -32315 2984
rect -31669 2951 -31598 2985
rect -32352 2911 -32344 2945
rect -31669 2917 -31632 2951
rect -32352 2872 -32315 2911
rect -31669 2883 -31598 2917
rect -32352 2838 -32344 2872
rect -31669 2849 -31632 2883
rect -32352 2799 -32315 2838
rect -31669 2815 -31598 2849
rect -32352 2765 -32344 2799
rect -31669 2781 -31632 2815
rect -32352 2726 -32315 2765
rect -31669 2747 -31598 2781
rect -32352 2692 -32344 2726
rect -31669 2713 -31632 2747
rect -32352 2653 -32315 2692
rect -31669 2679 -31598 2713
rect -32352 2619 -32344 2653
rect -31669 2645 -31632 2679
rect -32352 2580 -32315 2619
rect -31669 2611 -31598 2645
rect -32352 2546 -32344 2580
rect -31669 2577 -31632 2611
rect -32352 2507 -32315 2546
rect -31669 2543 -31598 2577
rect -31669 2509 -31632 2543
rect -32352 2473 -32344 2507
rect -31669 2475 -31598 2509
rect -32352 2434 -32315 2473
rect -31669 2441 -31632 2475
rect -32352 2400 -32344 2434
rect -31669 2407 -31598 2441
rect -32352 2361 -32315 2400
rect -31669 2373 -31632 2407
rect -32352 2327 -32344 2361
rect -31669 2339 -31598 2373
rect -32352 2288 -32315 2327
rect -31669 2305 -31632 2339
rect -32352 2254 -32344 2288
rect -31669 2271 -31598 2305
rect -32352 2215 -32315 2254
rect -31669 2237 -31632 2271
rect -32352 2181 -32344 2215
rect -31669 2203 -31598 2237
rect -32352 2142 -32315 2181
rect -31669 2169 -31632 2203
rect -32352 2108 -32344 2142
rect -31669 2135 -31598 2169
rect -32352 2069 -32315 2108
rect -31669 2101 -31632 2135
rect -32352 2035 -32344 2069
rect -31669 2067 -31598 2101
rect -32352 1996 -32315 2035
rect -31669 2033 -31632 2067
rect -31669 1999 -31598 2033
rect -32352 1962 -32344 1996
rect -31669 1965 -31632 1999
rect -32352 1923 -32315 1962
rect -31669 1931 -31598 1965
rect -32352 1889 -32344 1923
rect -31669 1897 -31632 1931
rect -32352 1850 -32315 1889
rect -31669 1863 -31598 1897
rect -32352 1816 -32344 1850
rect -31669 1829 -31632 1863
rect -32352 1777 -32315 1816
rect -31669 1795 -31598 1829
rect -32352 1743 -32344 1777
rect -31669 1761 -31632 1795
rect -32352 1704 -32315 1743
rect -31669 1727 -31598 1761
rect -32352 1670 -32344 1704
rect -31669 1693 -31632 1727
rect -32352 1631 -32315 1670
rect -31669 1659 -31598 1693
rect -32352 1597 -32344 1631
rect -31669 1625 -31632 1659
rect -32352 1558 -32315 1597
rect -31669 1591 -31598 1625
rect -32352 1524 -32344 1558
rect -31669 1557 -31632 1591
rect -32352 1485 -32315 1524
rect -31669 1523 -31598 1557
rect -31669 1489 -31632 1523
rect -32352 1451 -32344 1485
rect -31669 1455 -31598 1489
rect -32352 1412 -32315 1451
rect -31669 1421 -31632 1455
rect -32352 1378 -32344 1412
rect -31669 1387 -31598 1421
rect -32352 1339 -32315 1378
rect -31669 1353 -31632 1387
rect -32352 1305 -32344 1339
rect -31669 1319 -31598 1353
rect -32352 1266 -32315 1305
rect -31669 1285 -31632 1319
rect -32352 1232 -32344 1266
rect -31669 1251 -31598 1285
rect -32352 1193 -32315 1232
rect -31669 1217 -31632 1251
rect -32352 1159 -32344 1193
rect -31669 1183 -31598 1217
rect -32352 1120 -32315 1159
rect -31669 1149 -31632 1183
rect -32352 1086 -32344 1120
rect -31669 1115 -31598 1149
rect -32352 1047 -32315 1086
rect -31669 1081 -31632 1115
rect -31669 1047 -31598 1081
rect -32352 1013 -32344 1047
rect -31669 1013 -31632 1047
rect -32352 974 -32315 1013
rect -31669 979 -31598 1013
rect -32352 940 -32344 974
rect -31669 945 -31632 979
rect -32352 901 -32315 940
rect -31669 911 -31598 945
rect -32352 867 -32344 901
rect -31669 877 -31632 911
rect -32352 828 -32315 867
rect -31669 843 -31598 877
rect -32352 794 -32344 828
rect -31669 809 -31632 843
rect -32352 755 -32315 794
rect -31669 775 -31598 809
rect -32352 721 -32344 755
rect -31669 741 -31632 775
rect -32352 682 -32315 721
rect -31669 707 -31598 741
rect -32352 648 -32344 682
rect -31669 673 -31632 707
rect -32352 610 -32315 648
rect -31669 639 -31598 673
rect -32352 576 -32344 610
rect -31669 605 -31632 639
rect -32352 538 -32315 576
rect -31669 571 -31598 605
rect -32352 504 -32344 538
rect -31669 537 -31632 571
rect -32352 466 -32315 504
rect -31669 503 -31598 537
rect -31669 469 -31632 503
rect -32352 432 -32344 466
rect -31669 435 -31598 469
rect -32352 394 -32315 432
rect -31669 401 -31632 435
rect -32352 360 -32344 394
rect -31669 367 -31598 401
rect -32352 322 -32315 360
rect -31669 333 -31632 367
rect -32352 288 -32344 322
rect -31669 299 -31598 333
rect -32352 250 -32315 288
rect -31669 265 -31632 299
rect -32352 216 -32344 250
rect -31669 231 -31598 265
rect -32352 178 -32315 216
rect -31669 197 -31632 231
rect -32352 144 -32344 178
rect -31669 163 -31598 197
rect -32352 106 -32315 144
rect -31669 129 -31632 163
rect -32352 72 -32344 106
rect -31669 95 -31598 129
rect -32352 34 -32315 72
rect -31669 61 -31632 95
rect -32352 0 -32344 34
rect -31669 27 -31598 61
rect -32352 -38 -32315 0
rect -31669 -7 -31632 27
rect -32352 -72 -32344 -38
rect -31669 -41 -31598 -7
rect -32352 -110 -32315 -72
rect -31669 -75 -31632 -41
rect -31669 -109 -31598 -75
rect -32352 -144 -32344 -110
rect -31669 -143 -31632 -109
rect -32352 -182 -32315 -144
rect -31669 -177 -31598 -143
rect -32352 -216 -32344 -182
rect -31669 -211 -31632 -177
rect -32352 -254 -32315 -216
rect -31669 -245 -31598 -211
rect -32352 -288 -32344 -254
rect -31669 -279 -31632 -245
rect -32352 -326 -32315 -288
rect -31669 -313 -31598 -279
rect -32352 -360 -32344 -326
rect -31669 -347 -31632 -313
rect -32352 -398 -32315 -360
rect -31669 -381 -31598 -347
rect -32352 -432 -32344 -398
rect -31669 -415 -31632 -381
rect -32352 -470 -32315 -432
rect -31669 -449 -31598 -415
rect -32352 -504 -32344 -470
rect -31669 -483 -31632 -449
rect -32352 -542 -32315 -504
rect -31669 -517 -31598 -483
rect -32352 -576 -32344 -542
rect -31669 -551 -31632 -517
rect -32352 -614 -32315 -576
rect -31669 -585 -31598 -551
rect -32352 -648 -32344 -614
rect -31669 -619 -31632 -585
rect -32352 -686 -32315 -648
rect -31669 -653 -31598 -619
rect -32352 -720 -32344 -686
rect -31669 -687 -31632 -653
rect -32352 -758 -32315 -720
rect -31669 -721 -31598 -687
rect -31669 -755 -31632 -721
rect -32352 -792 -32344 -758
rect -31669 -789 -31598 -755
rect -32352 -830 -32315 -792
rect -31669 -823 -31632 -789
rect -32352 -864 -32344 -830
rect -31669 -857 -31598 -823
rect -32352 -902 -32315 -864
rect -31669 -891 -31632 -857
rect -32352 -936 -32344 -902
rect -31669 -925 -31598 -891
rect -32352 -974 -32315 -936
rect -31669 -959 -31632 -925
rect -32352 -1008 -32344 -974
rect -31669 -993 -31598 -959
rect -32352 -1046 -32315 -1008
rect -31669 -1027 -31632 -993
rect -32352 -1080 -32344 -1046
rect -31669 -1061 -31598 -1027
rect -32352 -1118 -32315 -1080
rect -31669 -1095 -31632 -1061
rect -32352 -1152 -32344 -1118
rect -31669 -1129 -31598 -1095
rect -32352 -1190 -32315 -1152
rect -31669 -1163 -31632 -1129
rect -32352 -1224 -32344 -1190
rect -31669 -1197 -31598 -1163
rect -32352 -1262 -32315 -1224
rect -31669 -1231 -31632 -1197
rect -32352 -1296 -32344 -1262
rect -31669 -1265 -31598 -1231
rect -32352 -1334 -32315 -1296
rect -31669 -1299 -31632 -1265
rect -31669 -1333 -31598 -1299
rect -32352 -1368 -32344 -1334
rect -31669 -1367 -31632 -1333
rect -32352 -1406 -32315 -1368
rect -31669 -1401 -31598 -1367
rect -32352 -1440 -32344 -1406
rect -31669 -1435 -31632 -1401
rect -32352 -1478 -32315 -1440
rect -31669 -1469 -31598 -1435
rect -32352 -1512 -32344 -1478
rect -31669 -1503 -31632 -1469
rect -32352 -1550 -32315 -1512
rect -31669 -1537 -31598 -1503
rect -32352 -1584 -32344 -1550
rect -31669 -1571 -31632 -1537
rect -32352 -1622 -32315 -1584
rect -31669 -1605 -31598 -1571
rect -32352 -1656 -32344 -1622
rect -31669 -1639 -31632 -1605
rect -32352 -1694 -32315 -1656
rect -31669 -1673 -31598 -1639
rect -32352 -1728 -32344 -1694
rect -31669 -1707 -31632 -1673
rect -32352 -1766 -32315 -1728
rect -31669 -1741 -31598 -1707
rect -32352 -1800 -32344 -1766
rect -31669 -1775 -31632 -1741
rect -32352 -1838 -32315 -1800
rect -31669 -1809 -31598 -1775
rect -32352 -1872 -32344 -1838
rect -31669 -1843 -31632 -1809
rect -32352 -1910 -32315 -1872
rect -31669 -1877 -31598 -1843
rect -32352 -1944 -32344 -1910
rect -31669 -1911 -31632 -1877
rect -32352 -1982 -32315 -1944
rect -31669 -1945 -31598 -1911
rect -31669 -1979 -31632 -1945
rect -32352 -2016 -32344 -1982
rect -31669 -2013 -31598 -1979
rect -32352 -2054 -32315 -2016
rect -31669 -2047 -31632 -2013
rect -32352 -2088 -32344 -2054
rect -31669 -2081 -31598 -2047
rect -32352 -2126 -32315 -2088
rect -31669 -2115 -31632 -2081
rect -32352 -2160 -32344 -2126
rect -31669 -2149 -31598 -2115
rect -32352 -2198 -32315 -2160
rect -31669 -2183 -31632 -2149
rect -32352 -2232 -32344 -2198
rect -31669 -2217 -31598 -2183
rect -32352 -2270 -32315 -2232
rect -31669 -2251 -31632 -2217
rect -32352 -2304 -32344 -2270
rect -31669 -2285 -31598 -2251
rect -32352 -2342 -32315 -2304
rect -31669 -2319 -31632 -2285
rect -32352 -2376 -32344 -2342
rect -31669 -2353 -31598 -2319
rect -32352 -2414 -32315 -2376
rect -31669 -2387 -31632 -2353
rect -32352 -2448 -32344 -2414
rect -31669 -2421 -31598 -2387
rect -32352 -2486 -32315 -2448
rect -31669 -2455 -31632 -2421
rect -32352 -2520 -32344 -2486
rect -31669 -2489 -31598 -2455
rect -32352 -2558 -32315 -2520
rect -31669 -2523 -31632 -2489
rect -31669 -2557 -31598 -2523
rect -32352 -2592 -32344 -2558
rect -31669 -2591 -31632 -2557
rect -32352 -2630 -32315 -2592
rect -31669 -2625 -31598 -2591
rect -32352 -2664 -32344 -2630
rect -31669 -2659 -31632 -2625
rect -32352 -2702 -32315 -2664
rect -31669 -2693 -31598 -2659
rect -32352 -2736 -32344 -2702
rect -31669 -2727 -31632 -2693
rect -32352 -2774 -32315 -2736
rect -31669 -2761 -31598 -2727
rect -32352 -2808 -32344 -2774
rect -31669 -2795 -31632 -2761
rect -32352 -2846 -32315 -2808
rect -31669 -2829 -31598 -2795
rect -32352 -2880 -32344 -2846
rect -31669 -2863 -31632 -2829
rect -32352 -2918 -32315 -2880
rect -31669 -2897 -31598 -2863
rect -32352 -2952 -32344 -2918
rect -31669 -2931 -31632 -2897
rect -32352 -2990 -32315 -2952
rect -31669 -2965 -31598 -2931
rect -32352 -3024 -32344 -2990
rect -31669 -2999 -31632 -2965
rect -32352 -3062 -32315 -3024
rect -31669 -3033 -31598 -2999
rect -32352 -3096 -32344 -3062
rect -31669 -3067 -31632 -3033
rect -32352 -3134 -32315 -3096
rect -31669 -3101 -31598 -3067
rect -32352 -3168 -32344 -3134
rect -31669 -3135 -31632 -3101
rect -32352 -3206 -32315 -3168
rect -31669 -3169 -31598 -3135
rect -31669 -3203 -31632 -3169
rect -32352 -3240 -32344 -3206
rect -31669 -3237 -31598 -3203
rect -32352 -3278 -32315 -3240
rect -31669 -3271 -31632 -3237
rect -32352 -3312 -32344 -3278
rect -31669 -3305 -31598 -3271
rect -32352 -3350 -32315 -3312
rect -31669 -3339 -31632 -3305
rect -32352 -3384 -32344 -3350
rect -31669 -3373 -31598 -3339
rect -32352 -3422 -32315 -3384
rect -31669 -3407 -31632 -3373
rect -32352 -3456 -32344 -3422
rect -31669 -3441 -31598 -3407
rect -32352 -3494 -32315 -3456
rect -31669 -3475 -31632 -3441
rect -32352 -3528 -32344 -3494
rect -31669 -3509 -31598 -3475
rect -32352 -3566 -32315 -3528
rect -31669 -3543 -31632 -3509
rect -32352 -3600 -32344 -3566
rect -31669 -3577 -31598 -3543
rect -32352 -3638 -32315 -3600
rect -31669 -3611 -31632 -3577
rect -32352 -3672 -32344 -3638
rect -31669 -3645 -31598 -3611
rect -32352 -3710 -32315 -3672
rect -31669 -3679 -31632 -3645
rect -32352 -3744 -32344 -3710
rect -31669 -3713 -31598 -3679
rect -32352 -3782 -32315 -3744
rect -31669 -3747 -31632 -3713
rect -31669 -3781 -31598 -3747
rect -32352 -3816 -32344 -3782
rect -31669 -3815 -31632 -3781
rect -32352 -3854 -32315 -3816
rect -31669 -3849 -31598 -3815
rect -32352 -3888 -32344 -3854
rect -31669 -3883 -31632 -3849
rect -32352 -3926 -32315 -3888
rect -31669 -3917 -31598 -3883
rect -32352 -3960 -32344 -3926
rect -31669 -3951 -31632 -3917
rect -32352 -3998 -32315 -3960
rect -31669 -3985 -31598 -3951
rect -32352 -4032 -32344 -3998
rect -31669 -4019 -31632 -3985
rect -32352 -4070 -32315 -4032
rect -31669 -4053 -31598 -4019
rect -32352 -4104 -32344 -4070
rect -31669 -4087 -31632 -4053
rect -32352 -4142 -32315 -4104
rect -31669 -4121 -31598 -4087
rect -32352 -4176 -32344 -4142
rect -31669 -4155 -31632 -4121
rect -32352 -4214 -32315 -4176
rect -31669 -4189 -31598 -4155
rect -32352 -4248 -32344 -4214
rect -31669 -4223 -31632 -4189
rect -32352 -4286 -32315 -4248
rect -31669 -4257 -31598 -4223
rect -32352 -4320 -32344 -4286
rect -31669 -4291 -31632 -4257
rect -32352 -4358 -32315 -4320
rect -31669 -4325 -31598 -4291
rect -32352 -4392 -32344 -4358
rect -31669 -4359 -31632 -4325
rect -32352 -4430 -32315 -4392
rect -31669 -4393 -31598 -4359
rect -31669 -4427 -31632 -4393
rect -32352 -4464 -32344 -4430
rect -31669 -4461 -31598 -4427
rect -32352 -4502 -32315 -4464
rect -31669 -4495 -31632 -4461
rect -32352 -4536 -32344 -4502
rect -31669 -4529 -31598 -4495
rect -32352 -4574 -32315 -4536
rect -31669 -4563 -31632 -4529
rect -32352 -4608 -32344 -4574
rect -31669 -4597 -31598 -4563
rect -32352 -4646 -32315 -4608
rect -31669 -4631 -31632 -4597
rect -32352 -4680 -32344 -4646
rect -31669 -4665 -31598 -4631
rect -32352 -4718 -32315 -4680
rect -31669 -4699 -31632 -4665
rect -32352 -4752 -32344 -4718
rect -31669 -4733 -31598 -4699
rect -32352 -4790 -32315 -4752
rect -31669 -4767 -31632 -4733
rect -32352 -4824 -32344 -4790
rect -31669 -4801 -31598 -4767
rect -32352 -4862 -32315 -4824
rect -31669 -4835 -31632 -4801
rect -32352 -4896 -32344 -4862
rect -31669 -4869 -31598 -4835
rect -32352 -4934 -32315 -4896
rect -31669 -4903 -31632 -4869
rect -32352 -4968 -32344 -4934
rect -31669 -4937 -31598 -4903
rect -32352 -5006 -32315 -4968
rect -31669 -4971 -31632 -4937
rect -31669 -5005 -31598 -4971
rect -32352 -5040 -32344 -5006
rect -31669 -5039 -31632 -5005
rect -32352 -5078 -32315 -5040
rect -31669 -5073 -31598 -5039
rect -32352 -5112 -32344 -5078
rect -31669 -5107 -31632 -5073
rect -32352 -5150 -32315 -5112
rect -31669 -5141 -31598 -5107
rect -32352 -5184 -32344 -5150
rect -31669 -5175 -31632 -5141
rect -32352 -5222 -32315 -5184
rect -31669 -5209 -31598 -5175
rect -32352 -5256 -32344 -5222
rect -31669 -5243 -31632 -5209
rect -32352 -5294 -32315 -5256
rect -31669 -5277 -31598 -5243
rect -32352 -5328 -32344 -5294
rect -31669 -5311 -31632 -5277
rect -32352 -5366 -32315 -5328
rect -31669 -5345 -31598 -5311
rect -32352 -5400 -32344 -5366
rect -31669 -5379 -31632 -5345
rect -32352 -5438 -32315 -5400
rect -31669 -5413 -31598 -5379
rect -32352 -5472 -32344 -5438
rect -31669 -5447 -31632 -5413
rect -32352 -5510 -32315 -5472
rect -31669 -5481 -31598 -5447
rect -32352 -5544 -32344 -5510
rect -31669 -5515 -31632 -5481
rect -32352 -5582 -32315 -5544
rect -31669 -5549 -31598 -5515
rect -32352 -5616 -32344 -5582
rect -31669 -5583 -31632 -5549
rect -32352 -5654 -32315 -5616
rect -31669 -5617 -31598 -5583
rect -31669 -5651 -31632 -5617
rect -32352 -5688 -32344 -5654
rect -31669 -5685 -31598 -5651
rect -32352 -5726 -32315 -5688
rect -31669 -5719 -31632 -5685
rect -32352 -5760 -32344 -5726
rect -31669 -5753 -31598 -5719
rect -32352 -5798 -32315 -5760
rect -31669 -5787 -31632 -5753
rect -32352 -5832 -32344 -5798
rect -31669 -5821 -31598 -5787
rect -32352 -5870 -32315 -5832
rect -31669 -5855 -31632 -5821
rect -32352 -5904 -32344 -5870
rect -31669 -5889 -31598 -5855
rect -32352 -5942 -32315 -5904
rect -31669 -5923 -31632 -5889
rect -32352 -5976 -32344 -5942
rect -31669 -5957 -31598 -5923
rect -32352 -6014 -32315 -5976
rect -31669 -5991 -31632 -5957
rect -32352 -6048 -32344 -6014
rect -31669 -6025 -31598 -5991
rect -32352 -6086 -32315 -6048
rect -31669 -6059 -31632 -6025
rect -32352 -6120 -32344 -6086
rect -31669 -6093 -31598 -6059
rect -32352 -6158 -32315 -6120
rect -31669 -6127 -31632 -6093
rect -32352 -6192 -32344 -6158
rect -31669 -6161 -31598 -6127
rect -32352 -6230 -32315 -6192
rect -31669 -6195 -31632 -6161
rect -31669 -6229 -31598 -6195
rect -32352 -6264 -32344 -6230
rect -31669 -6263 -31632 -6229
rect -32352 -6302 -32315 -6264
rect -31669 -6297 -31598 -6263
rect -32352 -6336 -32344 -6302
rect -31669 -6331 -31632 -6297
rect -32352 -6374 -32315 -6336
rect -31669 -6365 -31598 -6331
rect -32352 -6408 -32344 -6374
rect -31669 -6399 -31632 -6365
rect -32352 -6446 -32315 -6408
rect -31669 -6433 -31598 -6399
rect -32352 -6480 -32344 -6446
rect -31669 -6467 -31632 -6433
rect -32352 -6518 -32315 -6480
rect -31669 -6501 -31598 -6467
rect -32352 -6552 -32344 -6518
rect -31669 -6535 -31632 -6501
rect -32352 -6590 -32315 -6552
rect -31669 -6569 -31598 -6535
rect -32352 -6624 -32344 -6590
rect -31669 -6603 -31632 -6569
rect -32352 -6662 -32315 -6624
rect -31669 -6637 -31598 -6603
rect -32352 -6696 -32344 -6662
rect -31669 -6671 -31632 -6637
rect -32352 -6734 -32315 -6696
rect -31669 -6705 -31598 -6671
rect -32352 -6768 -32344 -6734
rect -31669 -6739 -31632 -6705
rect -32352 -6806 -32315 -6768
rect -31669 -6773 -31598 -6739
rect -32352 -6840 -32344 -6806
rect -31669 -6807 -31632 -6773
rect -32352 -6878 -32315 -6840
rect -31669 -6841 -31598 -6807
rect -31669 -6875 -31632 -6841
rect -32352 -6912 -32344 -6878
rect -31669 -6909 -31598 -6875
rect -32352 -6950 -32315 -6912
rect -31669 -6943 -31632 -6909
rect -32352 -6984 -32344 -6950
rect -31669 -6977 -31598 -6943
rect -32352 -7022 -32315 -6984
rect -31669 -7011 -31632 -6977
rect -32352 -7056 -32344 -7022
rect -31669 -7045 -31598 -7011
rect -32352 -7094 -32315 -7056
rect -31669 -7079 -31632 -7045
rect -32352 -7128 -32344 -7094
rect -31669 -7113 -31598 -7079
rect -32352 -7166 -32315 -7128
rect -31669 -7147 -31632 -7113
rect -32352 -7200 -32344 -7166
rect -31669 -7181 -31598 -7147
rect -32352 -7238 -32315 -7200
rect -31669 -7215 -31632 -7181
rect -32352 -7272 -32344 -7238
rect -31669 -7249 -31598 -7215
rect -32352 -7310 -32315 -7272
rect -31669 -7283 -31632 -7249
rect -32352 -7344 -32344 -7310
rect -31669 -7317 -31598 -7283
rect -32352 -7382 -32315 -7344
rect -31669 -7351 -31632 -7317
rect -32352 -7416 -32344 -7382
rect -31669 -7385 -31598 -7351
rect -32352 -7454 -32315 -7416
rect -31669 -7419 -31632 -7385
rect -31669 -7453 -31598 -7419
rect -32352 -7488 -32344 -7454
rect -31669 -7487 -31632 -7453
rect -32352 -7526 -32315 -7488
rect -31669 -7521 -31598 -7487
rect -32352 -7560 -32344 -7526
rect -31669 -7555 -31632 -7521
rect -32352 -7598 -32315 -7560
rect -31669 -7589 -31598 -7555
rect -32352 -7632 -32344 -7598
rect -31669 -7623 -31632 -7589
rect -32352 -7670 -32315 -7632
rect -31669 -7657 -31598 -7623
rect -32352 -7704 -32344 -7670
rect -31669 -7691 -31632 -7657
rect -32352 -7742 -32315 -7704
rect -31669 -7725 -31598 -7691
rect -32352 -7776 -32344 -7742
rect -31669 -7759 -31632 -7725
rect -32352 -7814 -32315 -7776
rect -31669 -7793 -31598 -7759
rect -32352 -7848 -32344 -7814
rect -31669 -7827 -31632 -7793
rect -32352 -7886 -32315 -7848
rect -31669 -7861 -31598 -7827
rect -32352 -7920 -32344 -7886
rect -31669 -7895 -31632 -7861
rect -32352 -7958 -32315 -7920
rect -31669 -7929 -31598 -7895
rect -32352 -7992 -32344 -7958
rect -31669 -7963 -31632 -7929
rect -32352 -8030 -32315 -7992
rect -31669 -7997 -31598 -7963
rect -32352 -8064 -32344 -8030
rect -31669 -8031 -31632 -7997
rect -32352 -8102 -32315 -8064
rect -31669 -8065 -31598 -8031
rect -31669 -8099 -31632 -8065
rect -32352 -8136 -32344 -8102
rect -31669 -8133 -31598 -8099
rect -32352 -8174 -32315 -8136
rect -31669 -8167 -31632 -8133
rect -32352 -8208 -32344 -8174
rect -31669 -8201 -31598 -8167
rect -32352 -8246 -32315 -8208
rect -31669 -8235 -31632 -8201
rect -32352 -8280 -32344 -8246
rect -31669 -8269 -31598 -8235
rect -32352 -8318 -32315 -8280
rect -31669 -8303 -31632 -8269
rect -32352 -8352 -32344 -8318
rect -31669 -8337 -31598 -8303
rect -32352 -8390 -32315 -8352
rect -31669 -8371 -31632 -8337
rect -32352 -8424 -32344 -8390
rect -31669 -8405 -31598 -8371
rect -32352 -8462 -32315 -8424
rect -31669 -8439 -31632 -8405
rect -32352 -8496 -32344 -8462
rect -31669 -8473 -31598 -8439
rect -32352 -8534 -32315 -8496
rect -31669 -8507 -31632 -8473
rect -32352 -8568 -32344 -8534
rect -31669 -8541 -31598 -8507
rect -32352 -8606 -32315 -8568
rect -31669 -8575 -31632 -8541
rect -32352 -8640 -32344 -8606
rect -31669 -8609 -31598 -8575
rect -29148 3277 -29134 3300
rect -29100 3309 -29046 3311
rect -29012 3309 -28958 3311
rect -28924 3309 -28870 3311
rect -28836 3309 -27036 3311
rect -29100 3277 -29078 3309
rect -29012 3277 -29010 3309
rect -29148 3275 -29078 3277
rect -29044 3275 -29010 3277
rect -28976 3277 -28958 3309
rect -28976 3275 -28942 3277
rect -28908 3275 -28874 3309
rect -28836 3277 -28806 3309
rect -28840 3275 -28806 3277
rect -28772 3275 -28738 3309
rect -28704 3275 -28670 3309
rect -28636 3275 -28602 3309
rect -28568 3275 -28534 3309
rect -28500 3275 -28466 3309
rect -28432 3275 -28398 3309
rect -28364 3275 -28330 3309
rect -28296 3275 -28262 3309
rect -28228 3275 -28194 3309
rect -28160 3290 -28126 3309
rect -28092 3290 -28058 3309
rect -28024 3290 -27990 3309
rect -27956 3290 -27922 3309
rect -27888 3290 -27854 3309
rect -28155 3275 -28126 3290
rect -28081 3275 -28058 3290
rect -28007 3275 -27990 3290
rect -27933 3275 -27922 3290
rect -27859 3275 -27854 3290
rect -27820 3290 -27786 3309
rect -27752 3290 -27718 3309
rect -27684 3290 -27650 3309
rect -27616 3290 -27582 3309
rect -27548 3290 -27514 3309
rect -27480 3290 -27446 3309
rect -27820 3275 -27819 3290
rect -27752 3275 -27745 3290
rect -27684 3275 -27671 3290
rect -27616 3275 -27597 3290
rect -27548 3275 -27523 3290
rect -27480 3275 -27449 3290
rect -27412 3275 -27378 3309
rect -27344 3290 -27310 3309
rect -27276 3290 -27242 3309
rect -27208 3290 -27174 3309
rect -27140 3290 -27106 3309
rect -27341 3275 -27310 3290
rect -27267 3275 -27242 3290
rect -27193 3275 -27174 3290
rect -27119 3275 -27106 3290
rect -27072 3275 -27036 3309
rect -29148 3266 -28189 3275
rect -29114 3256 -28189 3266
rect -28155 3256 -28115 3275
rect -28081 3256 -28041 3275
rect -28007 3256 -27967 3275
rect -27933 3256 -27893 3275
rect -27859 3256 -27819 3275
rect -27785 3256 -27745 3275
rect -27711 3256 -27671 3275
rect -27637 3256 -27597 3275
rect -27563 3256 -27523 3275
rect -27489 3256 -27449 3275
rect -27415 3256 -27375 3275
rect -27341 3256 -27301 3275
rect -27267 3256 -27227 3275
rect -27193 3256 -27153 3275
rect -27119 3256 -27036 3275
rect -29114 3240 -27036 3256
rect -29114 3238 -29078 3240
rect -29044 3238 -29010 3240
rect -29148 3204 -29134 3232
rect -29100 3206 -29078 3238
rect -29012 3206 -29010 3238
rect -28976 3238 -28942 3240
rect -28976 3206 -28958 3238
rect -28908 3206 -28874 3240
rect -28840 3238 -28806 3240
rect -28836 3206 -28806 3238
rect -28772 3206 -28738 3240
rect -28704 3206 -28670 3240
rect -28636 3206 -28602 3240
rect -28568 3206 -28534 3240
rect -28500 3206 -28466 3240
rect -28432 3206 -28398 3240
rect -28364 3206 -28330 3240
rect -28296 3206 -28262 3240
rect -28228 3206 -28194 3240
rect -28160 3217 -28126 3240
rect -28092 3217 -28058 3240
rect -28024 3217 -27990 3240
rect -27956 3217 -27922 3240
rect -27888 3217 -27854 3240
rect -28155 3206 -28126 3217
rect -28081 3206 -28058 3217
rect -28007 3206 -27990 3217
rect -27933 3206 -27922 3217
rect -27859 3206 -27854 3217
rect -27820 3217 -27786 3240
rect -27752 3217 -27718 3240
rect -27684 3217 -27650 3240
rect -27616 3217 -27582 3240
rect -27548 3217 -27514 3240
rect -27480 3217 -27446 3240
rect -27820 3206 -27819 3217
rect -27752 3206 -27745 3217
rect -27684 3206 -27671 3217
rect -27616 3206 -27597 3217
rect -27548 3206 -27523 3217
rect -27480 3206 -27449 3217
rect -27412 3206 -27378 3240
rect -27344 3217 -27310 3240
rect -27276 3217 -27242 3240
rect -27208 3217 -27174 3240
rect -27140 3217 -27106 3240
rect -27341 3206 -27310 3217
rect -27267 3206 -27242 3217
rect -27193 3206 -27174 3217
rect -27119 3206 -27106 3217
rect -27072 3206 -27036 3240
rect -29100 3204 -29046 3206
rect -29012 3204 -28958 3206
rect -28924 3204 -28870 3206
rect -28836 3204 -28189 3206
rect -29148 3198 -28189 3204
rect -29114 3183 -28189 3198
rect -28155 3183 -28115 3206
rect -28081 3183 -28041 3206
rect -28007 3183 -27967 3206
rect -27933 3183 -27893 3206
rect -27859 3183 -27819 3206
rect -27785 3183 -27745 3206
rect -27711 3183 -27671 3206
rect -27637 3183 -27597 3206
rect -27563 3183 -27523 3206
rect -27489 3183 -27449 3206
rect -27415 3183 -27375 3206
rect -27341 3183 -27301 3206
rect -27267 3183 -27227 3206
rect -27193 3183 -27153 3206
rect -27119 3183 -27036 3206
rect -29114 3171 -27036 3183
rect -29114 3165 -29078 3171
rect -29044 3165 -29010 3171
rect -29148 3131 -29134 3164
rect -29100 3137 -29078 3165
rect -29012 3137 -29010 3165
rect -28976 3165 -28942 3171
rect -28976 3137 -28958 3165
rect -28908 3137 -28874 3171
rect -28840 3165 -28806 3171
rect -28836 3137 -28806 3165
rect -28772 3137 -28738 3171
rect -28704 3137 -28670 3171
rect -28636 3137 -28602 3171
rect -28568 3137 -28534 3171
rect -28500 3137 -28466 3171
rect -28432 3137 -28398 3171
rect -28364 3137 -28330 3171
rect -28296 3137 -28262 3171
rect -28228 3137 -28194 3171
rect -28160 3144 -28126 3171
rect -28092 3144 -28058 3171
rect -28024 3144 -27990 3171
rect -27956 3144 -27922 3171
rect -27888 3144 -27854 3171
rect -28155 3137 -28126 3144
rect -28081 3137 -28058 3144
rect -28007 3137 -27990 3144
rect -27933 3137 -27922 3144
rect -27859 3137 -27854 3144
rect -27820 3144 -27786 3171
rect -27752 3144 -27718 3171
rect -27684 3144 -27650 3171
rect -27616 3144 -27582 3171
rect -27548 3144 -27514 3171
rect -27480 3144 -27446 3171
rect -27820 3137 -27819 3144
rect -27752 3137 -27745 3144
rect -27684 3137 -27671 3144
rect -27616 3137 -27597 3144
rect -27548 3137 -27523 3144
rect -27480 3137 -27449 3144
rect -27412 3137 -27378 3171
rect -27344 3144 -27310 3171
rect -27276 3144 -27242 3171
rect -27208 3144 -27174 3171
rect -27140 3144 -27106 3171
rect -27341 3137 -27310 3144
rect -27267 3137 -27242 3144
rect -27193 3137 -27174 3144
rect -27119 3137 -27106 3144
rect -27072 3137 -27036 3171
rect -29100 3131 -29046 3137
rect -29012 3131 -28958 3137
rect -28924 3131 -28870 3137
rect -28836 3131 -28189 3137
rect -29148 3130 -28189 3131
rect -29114 3110 -28189 3130
rect -28155 3110 -28115 3137
rect -28081 3110 -28041 3137
rect -28007 3110 -27967 3137
rect -27933 3110 -27893 3137
rect -27859 3110 -27819 3137
rect -27785 3110 -27745 3137
rect -27711 3110 -27671 3137
rect -27637 3110 -27597 3137
rect -27563 3110 -27523 3137
rect -27489 3110 -27449 3137
rect -27415 3110 -27375 3137
rect -27341 3110 -27301 3137
rect -27267 3110 -27227 3137
rect -27193 3110 -27153 3137
rect -27119 3110 -27036 3137
rect -29114 3102 -27036 3110
rect -29114 3096 -29078 3102
rect -29148 3092 -29078 3096
rect -29044 3092 -29010 3102
rect -29148 3062 -29134 3092
rect -29100 3068 -29078 3092
rect -29012 3068 -29010 3092
rect -28976 3092 -28942 3102
rect -28976 3068 -28958 3092
rect -28908 3068 -28874 3102
rect -28840 3092 -28806 3102
rect -28836 3068 -28806 3092
rect -28772 3068 -28738 3102
rect -28704 3068 -28670 3102
rect -28636 3068 -28602 3102
rect -28568 3068 -28534 3102
rect -28500 3068 -28466 3102
rect -28432 3068 -28398 3102
rect -28364 3068 -28330 3102
rect -28296 3068 -28262 3102
rect -28228 3068 -28194 3102
rect -28160 3071 -28126 3102
rect -28092 3071 -28058 3102
rect -28024 3071 -27990 3102
rect -27956 3071 -27922 3102
rect -27888 3071 -27854 3102
rect -28155 3068 -28126 3071
rect -28081 3068 -28058 3071
rect -28007 3068 -27990 3071
rect -27933 3068 -27922 3071
rect -27859 3068 -27854 3071
rect -27820 3071 -27786 3102
rect -27752 3071 -27718 3102
rect -27684 3071 -27650 3102
rect -27616 3071 -27582 3102
rect -27548 3071 -27514 3102
rect -27480 3071 -27446 3102
rect -27820 3068 -27819 3071
rect -27752 3068 -27745 3071
rect -27684 3068 -27671 3071
rect -27616 3068 -27597 3071
rect -27548 3068 -27523 3071
rect -27480 3068 -27449 3071
rect -27412 3068 -27378 3102
rect -27344 3071 -27310 3102
rect -27276 3071 -27242 3102
rect -27208 3071 -27174 3102
rect -27140 3071 -27106 3102
rect -27341 3068 -27310 3071
rect -27267 3068 -27242 3071
rect -27193 3068 -27174 3071
rect -27119 3068 -27106 3071
rect -27072 3068 -27036 3102
rect -29100 3058 -29046 3068
rect -29012 3058 -28958 3068
rect -28924 3058 -28870 3068
rect -28836 3058 -28189 3068
rect -29114 3037 -28189 3058
rect -28155 3037 -28115 3068
rect -28081 3037 -28041 3068
rect -28007 3037 -27967 3068
rect -27933 3037 -27893 3068
rect -27859 3037 -27819 3068
rect -27785 3037 -27745 3068
rect -27711 3037 -27671 3068
rect -27637 3037 -27597 3068
rect -27563 3037 -27523 3068
rect -27489 3037 -27449 3068
rect -27415 3037 -27375 3068
rect -27341 3037 -27301 3068
rect -27267 3037 -27227 3068
rect -27193 3037 -27153 3068
rect -27119 3037 -27036 3068
rect -29114 3033 -27036 3037
rect -29114 3028 -29078 3033
rect -29148 3019 -29078 3028
rect -29044 3019 -29010 3033
rect -29148 2994 -29134 3019
rect -29100 2999 -29078 3019
rect -29012 2999 -29010 3019
rect -28976 3019 -28942 3033
rect -28976 2999 -28958 3019
rect -28908 2999 -28874 3033
rect -28840 3019 -28806 3033
rect -28836 2999 -28806 3019
rect -28772 2999 -28738 3033
rect -28704 2999 -28670 3033
rect -28636 2999 -28602 3033
rect -28568 2999 -28534 3033
rect -28500 2999 -28466 3033
rect -28432 2999 -28398 3033
rect -28364 2999 -28330 3033
rect -28296 2999 -28262 3033
rect -28228 2999 -28194 3033
rect -28160 2999 -28126 3033
rect -28092 2999 -28058 3033
rect -28024 2999 -27990 3033
rect -27956 2999 -27922 3033
rect -27888 2999 -27854 3033
rect -27820 2999 -27786 3033
rect -27752 2999 -27718 3033
rect -27684 2999 -27650 3033
rect -27616 2999 -27582 3033
rect -27548 2999 -27514 3033
rect -27480 2999 -27446 3033
rect -27412 2999 -27378 3033
rect -27344 2999 -27310 3033
rect -27276 2999 -27242 3033
rect -27208 2999 -27174 3033
rect -27140 2999 -27106 3033
rect -27072 2999 -27036 3033
rect -29100 2985 -29046 2999
rect -29012 2985 -28958 2999
rect -28924 2985 -28870 2999
rect -28836 2998 -27036 2999
rect -28836 2985 -28189 2998
rect -29114 2964 -28189 2985
rect -28155 2964 -28115 2998
rect -28081 2964 -28041 2998
rect -28007 2964 -27967 2998
rect -27933 2964 -27893 2998
rect -27859 2964 -27819 2998
rect -27785 2964 -27745 2998
rect -27711 2964 -27671 2998
rect -27637 2964 -27597 2998
rect -27563 2964 -27523 2998
rect -27489 2964 -27449 2998
rect -27415 2964 -27375 2998
rect -27341 2964 -27301 2998
rect -27267 2964 -27227 2998
rect -27193 2964 -27153 2998
rect -27119 2964 -27036 2998
rect -29114 2960 -29078 2964
rect -29148 2946 -29078 2960
rect -29044 2946 -29010 2964
rect -29148 2926 -29134 2946
rect -29100 2930 -29078 2946
rect -29012 2930 -29010 2946
rect -28976 2946 -28942 2964
rect -28976 2930 -28958 2946
rect -28908 2930 -28874 2964
rect -28840 2946 -28806 2964
rect -28836 2930 -28806 2946
rect -28772 2930 -28738 2964
rect -28704 2930 -28670 2964
rect -28636 2930 -28602 2964
rect -28568 2930 -28534 2964
rect -28500 2930 -28466 2964
rect -28432 2930 -28398 2964
rect -28364 2930 -28330 2964
rect -28296 2930 -28262 2964
rect -28228 2930 -28194 2964
rect -28160 2930 -28126 2964
rect -28092 2930 -28058 2964
rect -28024 2930 -27990 2964
rect -27956 2930 -27922 2964
rect -27888 2930 -27854 2964
rect -27820 2930 -27786 2964
rect -27752 2930 -27718 2964
rect -27684 2930 -27650 2964
rect -27616 2930 -27582 2964
rect -27548 2930 -27514 2964
rect -27480 2930 -27446 2964
rect -27412 2930 -27378 2964
rect -27344 2930 -27310 2964
rect -27276 2930 -27242 2964
rect -27208 2930 -27174 2964
rect -27140 2930 -27106 2964
rect -27072 2930 -27036 2964
rect -29100 2912 -29046 2930
rect -29012 2912 -28958 2930
rect -28924 2912 -28870 2930
rect -28836 2925 -27036 2930
rect -28836 2912 -28189 2925
rect -29114 2895 -28189 2912
rect -28155 2895 -28115 2925
rect -28081 2895 -28041 2925
rect -28007 2895 -27967 2925
rect -27933 2895 -27893 2925
rect -27859 2895 -27819 2925
rect -27785 2895 -27745 2925
rect -27711 2895 -27671 2925
rect -27637 2895 -27597 2925
rect -27563 2895 -27523 2925
rect -27489 2895 -27449 2925
rect -27415 2895 -27375 2925
rect -27341 2895 -27301 2925
rect -27267 2895 -27227 2925
rect -27193 2895 -27153 2925
rect -27119 2895 -27036 2925
rect -29114 2892 -29078 2895
rect -29148 2873 -29078 2892
rect -29044 2873 -29010 2895
rect -29148 2858 -29134 2873
rect -29100 2861 -29078 2873
rect -29012 2861 -29010 2873
rect -28976 2873 -28942 2895
rect -28976 2861 -28958 2873
rect -28908 2861 -28874 2895
rect -28840 2873 -28806 2895
rect -28836 2861 -28806 2873
rect -28772 2861 -28738 2895
rect -28704 2861 -28670 2895
rect -28636 2861 -28602 2895
rect -28568 2861 -28534 2895
rect -28500 2861 -28466 2895
rect -28432 2861 -28398 2895
rect -28364 2861 -28330 2895
rect -28296 2861 -28262 2895
rect -28228 2861 -28194 2895
rect -28155 2891 -28126 2895
rect -28081 2891 -28058 2895
rect -28007 2891 -27990 2895
rect -27933 2891 -27922 2895
rect -27859 2891 -27854 2895
rect -28160 2861 -28126 2891
rect -28092 2861 -28058 2891
rect -28024 2861 -27990 2891
rect -27956 2861 -27922 2891
rect -27888 2861 -27854 2891
rect -27820 2891 -27819 2895
rect -27752 2891 -27745 2895
rect -27684 2891 -27671 2895
rect -27616 2891 -27597 2895
rect -27548 2891 -27523 2895
rect -27480 2891 -27449 2895
rect -27820 2861 -27786 2891
rect -27752 2861 -27718 2891
rect -27684 2861 -27650 2891
rect -27616 2861 -27582 2891
rect -27548 2861 -27514 2891
rect -27480 2861 -27446 2891
rect -27412 2861 -27378 2895
rect -27341 2891 -27310 2895
rect -27267 2891 -27242 2895
rect -27193 2891 -27174 2895
rect -27119 2891 -27106 2895
rect -27344 2861 -27310 2891
rect -27276 2861 -27242 2891
rect -27208 2861 -27174 2891
rect -27140 2861 -27106 2891
rect -27072 2861 -27036 2895
rect -29100 2839 -29046 2861
rect -29012 2839 -28958 2861
rect -28924 2839 -28870 2861
rect -28836 2852 -27036 2861
rect -28836 2839 -28189 2852
rect -29114 2826 -28189 2839
rect -28155 2826 -28115 2852
rect -28081 2826 -28041 2852
rect -28007 2826 -27967 2852
rect -27933 2826 -27893 2852
rect -27859 2826 -27819 2852
rect -27785 2826 -27745 2852
rect -27711 2826 -27671 2852
rect -27637 2826 -27597 2852
rect -27563 2826 -27523 2852
rect -27489 2826 -27449 2852
rect -27415 2826 -27375 2852
rect -27341 2826 -27301 2852
rect -27267 2826 -27227 2852
rect -27193 2826 -27153 2852
rect -27119 2826 -27036 2852
rect -29114 2824 -29078 2826
rect -29148 2800 -29078 2824
rect -29044 2800 -29010 2826
rect -29148 2790 -29134 2800
rect -29100 2792 -29078 2800
rect -29012 2792 -29010 2800
rect -28976 2800 -28942 2826
rect -28976 2792 -28958 2800
rect -28908 2792 -28874 2826
rect -28840 2800 -28806 2826
rect -28836 2792 -28806 2800
rect -28772 2792 -28738 2826
rect -28704 2792 -28670 2826
rect -28636 2792 -28602 2826
rect -28568 2792 -28534 2826
rect -28500 2792 -28466 2826
rect -28432 2792 -28398 2826
rect -28364 2792 -28330 2826
rect -28296 2792 -28262 2826
rect -28228 2792 -28194 2826
rect -28155 2818 -28126 2826
rect -28081 2818 -28058 2826
rect -28007 2818 -27990 2826
rect -27933 2818 -27922 2826
rect -27859 2818 -27854 2826
rect -28160 2792 -28126 2818
rect -28092 2792 -28058 2818
rect -28024 2792 -27990 2818
rect -27956 2792 -27922 2818
rect -27888 2792 -27854 2818
rect -27820 2818 -27819 2826
rect -27752 2818 -27745 2826
rect -27684 2818 -27671 2826
rect -27616 2818 -27597 2826
rect -27548 2818 -27523 2826
rect -27480 2818 -27449 2826
rect -27820 2792 -27786 2818
rect -27752 2792 -27718 2818
rect -27684 2792 -27650 2818
rect -27616 2792 -27582 2818
rect -27548 2792 -27514 2818
rect -27480 2792 -27446 2818
rect -27412 2792 -27378 2826
rect -27341 2818 -27310 2826
rect -27267 2818 -27242 2826
rect -27193 2818 -27174 2826
rect -27119 2818 -27106 2826
rect -27344 2792 -27310 2818
rect -27276 2792 -27242 2818
rect -27208 2792 -27174 2818
rect -27140 2792 -27106 2818
rect -27072 2792 -27036 2826
rect -29100 2766 -29046 2792
rect -29012 2766 -28958 2792
rect -28924 2766 -28870 2792
rect -28836 2779 -27036 2792
rect -28836 2766 -28189 2779
rect -29114 2757 -28189 2766
rect -28155 2757 -28115 2779
rect -28081 2757 -28041 2779
rect -28007 2757 -27967 2779
rect -27933 2757 -27893 2779
rect -27859 2757 -27819 2779
rect -27785 2757 -27745 2779
rect -27711 2757 -27671 2779
rect -27637 2757 -27597 2779
rect -27563 2757 -27523 2779
rect -27489 2757 -27449 2779
rect -27415 2757 -27375 2779
rect -27341 2757 -27301 2779
rect -27267 2757 -27227 2779
rect -27193 2757 -27153 2779
rect -27119 2757 -27036 2779
rect -29114 2756 -29078 2757
rect -29148 2727 -29078 2756
rect -29044 2727 -29010 2757
rect -29148 2722 -29134 2727
rect -29100 2723 -29078 2727
rect -29012 2723 -29010 2727
rect -28976 2727 -28942 2757
rect -28976 2723 -28958 2727
rect -28908 2723 -28874 2757
rect -28840 2727 -28806 2757
rect -28836 2723 -28806 2727
rect -28772 2723 -28738 2757
rect -28704 2723 -28670 2757
rect -28636 2723 -28602 2757
rect -28568 2723 -28534 2757
rect -28500 2723 -28466 2757
rect -28432 2723 -28398 2757
rect -28364 2723 -28330 2757
rect -28296 2723 -28262 2757
rect -28228 2723 -28194 2757
rect -28155 2745 -28126 2757
rect -28081 2745 -28058 2757
rect -28007 2745 -27990 2757
rect -27933 2745 -27922 2757
rect -27859 2745 -27854 2757
rect -28160 2723 -28126 2745
rect -28092 2723 -28058 2745
rect -28024 2723 -27990 2745
rect -27956 2723 -27922 2745
rect -27888 2723 -27854 2745
rect -27820 2745 -27819 2757
rect -27752 2745 -27745 2757
rect -27684 2745 -27671 2757
rect -27616 2745 -27597 2757
rect -27548 2745 -27523 2757
rect -27480 2745 -27449 2757
rect -27820 2723 -27786 2745
rect -27752 2723 -27718 2745
rect -27684 2723 -27650 2745
rect -27616 2723 -27582 2745
rect -27548 2723 -27514 2745
rect -27480 2723 -27446 2745
rect -27412 2723 -27378 2757
rect -27341 2745 -27310 2757
rect -27267 2745 -27242 2757
rect -27193 2745 -27174 2757
rect -27119 2745 -27106 2757
rect -27344 2723 -27310 2745
rect -27276 2723 -27242 2745
rect -27208 2723 -27174 2745
rect -27140 2723 -27106 2745
rect -27072 2723 -27036 2757
rect -29100 2693 -29046 2723
rect -29012 2693 -28958 2723
rect -28924 2693 -28870 2723
rect -28836 2706 -27036 2723
rect -28836 2693 -28189 2706
rect -29114 2688 -28189 2693
rect -28155 2688 -28115 2706
rect -28081 2688 -28041 2706
rect -28007 2688 -27967 2706
rect -27933 2688 -27893 2706
rect -27859 2688 -27819 2706
rect -27785 2688 -27745 2706
rect -27711 2688 -27671 2706
rect -27637 2688 -27597 2706
rect -27563 2688 -27523 2706
rect -27489 2688 -27449 2706
rect -27415 2688 -27375 2706
rect -27341 2688 -27301 2706
rect -27267 2688 -27227 2706
rect -27193 2688 -27153 2706
rect -27119 2688 -27036 2706
rect -29148 2654 -29078 2688
rect -29044 2654 -29010 2688
rect -28976 2654 -28942 2688
rect -28908 2654 -28874 2688
rect -28840 2654 -28806 2688
rect -28772 2654 -28738 2688
rect -28704 2654 -28670 2688
rect -28636 2654 -28602 2688
rect -28568 2654 -28534 2688
rect -28500 2654 -28466 2688
rect -28432 2654 -28398 2688
rect -28364 2654 -28330 2688
rect -28296 2654 -28262 2688
rect -28228 2654 -28194 2688
rect -28155 2672 -28126 2688
rect -28081 2672 -28058 2688
rect -28007 2672 -27990 2688
rect -27933 2672 -27922 2688
rect -27859 2672 -27854 2688
rect -28160 2654 -28126 2672
rect -28092 2654 -28058 2672
rect -28024 2654 -27990 2672
rect -27956 2654 -27922 2672
rect -27888 2654 -27854 2672
rect -27820 2672 -27819 2688
rect -27752 2672 -27745 2688
rect -27684 2672 -27671 2688
rect -27616 2672 -27597 2688
rect -27548 2672 -27523 2688
rect -27480 2672 -27449 2688
rect -27820 2654 -27786 2672
rect -27752 2654 -27718 2672
rect -27684 2654 -27650 2672
rect -27616 2654 -27582 2672
rect -27548 2654 -27514 2672
rect -27480 2654 -27446 2672
rect -27412 2654 -27378 2688
rect -27341 2672 -27310 2688
rect -27267 2672 -27242 2688
rect -27193 2672 -27174 2688
rect -27119 2672 -27106 2688
rect -27344 2654 -27310 2672
rect -27276 2654 -27242 2672
rect -27208 2654 -27174 2672
rect -27140 2654 -27106 2672
rect -27072 2654 -27036 2688
rect -29100 2620 -29046 2654
rect -29012 2620 -28958 2654
rect -28924 2620 -28870 2654
rect -28836 2633 -27036 2654
rect -28836 2620 -28189 2633
rect -29148 2619 -28189 2620
rect -28155 2619 -28115 2633
rect -28081 2619 -28041 2633
rect -28007 2619 -27967 2633
rect -27933 2619 -27893 2633
rect -27859 2619 -27819 2633
rect -27785 2619 -27745 2633
rect -27711 2619 -27671 2633
rect -27637 2619 -27597 2633
rect -27563 2619 -27523 2633
rect -27489 2619 -27449 2633
rect -27415 2619 -27375 2633
rect -27341 2619 -27301 2633
rect -27267 2619 -27227 2633
rect -27193 2619 -27153 2633
rect -27119 2619 -27036 2633
rect -29148 2586 -29078 2619
rect -29114 2585 -29078 2586
rect -29044 2585 -29010 2619
rect -28976 2585 -28942 2619
rect -28908 2585 -28874 2619
rect -28840 2585 -28806 2619
rect -28772 2585 -28738 2619
rect -28704 2585 -28670 2619
rect -28636 2585 -28602 2619
rect -28568 2585 -28534 2619
rect -28500 2585 -28466 2619
rect -28432 2585 -28398 2619
rect -28364 2585 -28330 2619
rect -28296 2585 -28262 2619
rect -28228 2585 -28194 2619
rect -28155 2599 -28126 2619
rect -28081 2599 -28058 2619
rect -28007 2599 -27990 2619
rect -27933 2599 -27922 2619
rect -27859 2599 -27854 2619
rect -28160 2585 -28126 2599
rect -28092 2585 -28058 2599
rect -28024 2585 -27990 2599
rect -27956 2585 -27922 2599
rect -27888 2585 -27854 2599
rect -27820 2599 -27819 2619
rect -27752 2599 -27745 2619
rect -27684 2599 -27671 2619
rect -27616 2599 -27597 2619
rect -27548 2599 -27523 2619
rect -27480 2599 -27449 2619
rect -27820 2585 -27786 2599
rect -27752 2585 -27718 2599
rect -27684 2585 -27650 2599
rect -27616 2585 -27582 2599
rect -27548 2585 -27514 2599
rect -27480 2585 -27446 2599
rect -27412 2585 -27378 2619
rect -27341 2599 -27310 2619
rect -27267 2599 -27242 2619
rect -27193 2599 -27174 2619
rect -27119 2599 -27106 2619
rect -27344 2585 -27310 2599
rect -27276 2585 -27242 2599
rect -27208 2585 -27174 2599
rect -27140 2585 -27106 2599
rect -27072 2585 -27036 2619
rect -29114 2581 -27036 2585
rect -29148 2547 -29134 2552
rect -29100 2550 -29046 2581
rect -29012 2550 -28958 2581
rect -28924 2550 -28870 2581
rect -28836 2560 -27036 2581
rect -746 3510 -712 3512
rect -746 3474 -712 3476
rect -746 3402 -712 3408
rect -746 3330 -712 3340
rect -746 3258 -712 3272
rect -746 3186 -712 3204
rect -746 3114 -712 3136
rect -746 3042 -712 3068
rect -746 2970 -712 3000
rect -746 2898 -712 2932
rect -746 2830 -712 2864
rect -746 2762 -712 2792
rect -746 2694 -712 2720
rect -746 2626 -712 2648
rect -590 3510 -556 3512
rect -590 3474 -556 3476
rect -590 3402 -556 3408
rect -590 3330 -556 3340
rect -590 3258 -556 3272
rect -590 3186 -556 3204
rect -590 3114 -556 3136
rect -590 3042 -556 3068
rect -590 2970 -556 3000
rect -590 2898 -556 2932
rect -590 2830 -556 2864
rect -590 2762 -556 2792
rect -590 2694 -556 2720
rect -590 2626 -556 2648
rect -434 3510 -400 3512
rect -434 3474 -400 3476
rect -434 3402 -400 3408
rect -434 3330 -400 3340
rect -434 3258 -400 3272
rect -434 3186 -400 3204
rect -434 3114 -400 3136
rect -434 3042 -400 3068
rect -434 2970 -400 3000
rect -434 2898 -400 2932
rect -434 2830 -400 2864
rect -434 2762 -400 2792
rect -434 2694 -400 2720
rect -434 2626 -400 2648
rect 168 3510 202 3512
rect 168 3474 202 3476
rect 168 3402 202 3408
rect 168 3330 202 3340
rect 168 3258 202 3272
rect 168 3186 202 3204
rect 168 3114 202 3136
rect 168 3042 202 3068
rect 168 2970 202 3000
rect 168 2898 202 2932
rect 168 2830 202 2864
rect 168 2762 202 2792
rect 168 2694 202 2720
rect 168 2626 202 2648
rect 324 3510 358 3512
rect 324 3474 358 3476
rect 324 3402 358 3408
rect 324 3330 358 3340
rect 324 3258 358 3272
rect 324 3186 358 3204
rect 324 3114 358 3136
rect 324 3042 358 3068
rect 324 2970 358 3000
rect 324 2898 358 2932
rect 324 2830 358 2864
rect 324 2762 358 2792
rect 324 2694 358 2720
rect 324 2626 358 2648
rect 480 3510 514 3512
rect 480 3474 514 3476
rect 480 3402 514 3408
rect 480 3330 514 3340
rect 480 3258 514 3272
rect 480 3186 514 3204
rect 480 3114 514 3136
rect 480 3042 514 3068
rect 480 2970 514 3000
rect 480 2898 514 2932
rect 480 2830 514 2864
rect 480 2762 514 2792
rect 480 2694 514 2720
rect 480 2626 514 2648
rect 616 3510 650 3512
rect 616 3474 650 3476
rect 616 3402 650 3408
rect 616 3330 650 3340
rect 616 3258 650 3272
rect 616 3186 650 3204
rect 616 3114 650 3136
rect 616 3042 650 3068
rect 616 2970 650 3000
rect 616 2898 650 2932
rect 616 2830 650 2864
rect 616 2762 650 2792
rect 616 2694 650 2720
rect 616 2626 650 2648
rect 772 3510 806 3512
rect 772 3474 806 3476
rect 772 3402 806 3408
rect 772 3330 806 3340
rect 772 3258 806 3272
rect 772 3186 806 3204
rect 772 3114 806 3136
rect 772 3042 806 3068
rect 772 2970 806 3000
rect 772 2898 806 2932
rect 772 2830 806 2864
rect 772 2762 806 2792
rect 772 2694 806 2720
rect 772 2626 806 2648
rect 928 3510 962 3512
rect 928 3474 962 3476
rect 928 3402 962 3408
rect 928 3330 962 3340
rect 928 3258 962 3272
rect 928 3186 962 3204
rect 928 3114 962 3136
rect 928 3042 962 3068
rect 928 2970 962 3000
rect 928 2898 962 2932
rect 928 2830 962 2864
rect 928 2762 962 2792
rect 928 2694 962 2720
rect 928 2626 962 2648
rect 1055 3510 1089 3512
rect 1055 3474 1089 3476
rect 1055 3402 1089 3408
rect 1055 3330 1089 3340
rect 1055 3258 1089 3272
rect 1055 3186 1089 3204
rect 1055 3114 1089 3136
rect 1055 3042 1089 3068
rect 1055 2970 1089 3000
rect 1055 2898 1089 2932
rect 1055 2830 1089 2864
rect 1055 2762 1089 2792
rect 1055 2694 1089 2720
rect 1055 2626 1089 2648
rect 1211 3510 1245 3512
rect 1211 3474 1245 3476
rect 1211 3402 1245 3408
rect 1211 3330 1245 3340
rect 1211 3258 1245 3272
rect 1211 3186 1245 3204
rect 1211 3114 1245 3136
rect 1211 3042 1245 3068
rect 1211 2970 1245 3000
rect 1211 2898 1245 2932
rect 1211 2830 1245 2864
rect 1211 2762 1245 2792
rect 1211 2694 1245 2720
rect 1211 2626 1245 2648
rect 1415 3510 1449 3512
rect 1415 3474 1449 3476
rect 1415 3402 1449 3408
rect 1415 3330 1449 3340
rect 1415 3258 1449 3272
rect 1415 3186 1449 3204
rect 1415 3114 1449 3136
rect 1415 3042 1449 3068
rect 1415 2970 1449 3000
rect 1415 2898 1449 2932
rect 1415 2830 1449 2864
rect 1415 2762 1449 2792
rect 1415 2694 1449 2720
rect 1415 2626 1449 2648
rect 1571 3510 1605 3512
rect 1571 3474 1605 3476
rect 1571 3402 1605 3408
rect 1571 3330 1605 3340
rect 1571 3258 1605 3272
rect 1571 3186 1605 3204
rect 1571 3114 1605 3136
rect 1571 3042 1605 3068
rect 1571 2970 1605 3000
rect 1571 2898 1605 2932
rect 1571 2830 1605 2864
rect 1571 2762 1605 2792
rect 1571 2694 1605 2720
rect 1571 2626 1605 2648
rect 1708 3475 1742 3477
rect 1708 3439 1742 3441
rect 1708 3367 1742 3373
rect 1708 3295 1742 3305
rect 1708 3223 1742 3237
rect 1708 3151 1742 3169
rect 1708 3079 1742 3101
rect 1708 3007 1742 3033
rect 1708 2935 1742 2965
rect 1708 2863 1742 2897
rect 1708 2795 1742 2829
rect 1708 2727 1742 2757
rect 1708 2659 1742 2685
rect 1708 2591 1742 2613
rect -28836 2550 -28189 2560
rect -28155 2550 -28115 2560
rect -28081 2550 -28041 2560
rect -28007 2550 -27967 2560
rect -27933 2550 -27893 2560
rect -27859 2550 -27819 2560
rect -27785 2550 -27745 2560
rect -27711 2550 -27671 2560
rect -27637 2550 -27597 2560
rect -27563 2550 -27523 2560
rect -27489 2550 -27449 2560
rect -27415 2550 -27375 2560
rect -27341 2550 -27301 2560
rect -27267 2550 -27227 2560
rect -27193 2550 -27153 2560
rect -27119 2550 -27036 2560
rect -29100 2547 -29078 2550
rect -29012 2547 -29010 2550
rect -29148 2518 -29078 2547
rect -29114 2516 -29078 2518
rect -29044 2516 -29010 2547
rect -28976 2547 -28958 2550
rect -28976 2516 -28942 2547
rect -28908 2516 -28874 2550
rect -28836 2547 -28806 2550
rect -28840 2516 -28806 2547
rect -28772 2516 -28738 2550
rect -28704 2516 -28670 2550
rect -28636 2516 -28602 2550
rect -28568 2516 -28534 2550
rect -28500 2516 -28466 2550
rect -28432 2516 -28398 2550
rect -28364 2516 -28330 2550
rect -28296 2516 -28262 2550
rect -28228 2516 -28194 2550
rect -28155 2526 -28126 2550
rect -28081 2526 -28058 2550
rect -28007 2526 -27990 2550
rect -27933 2526 -27922 2550
rect -27859 2526 -27854 2550
rect -28160 2516 -28126 2526
rect -28092 2516 -28058 2526
rect -28024 2516 -27990 2526
rect -27956 2516 -27922 2526
rect -27888 2516 -27854 2526
rect -27820 2526 -27819 2550
rect -27752 2526 -27745 2550
rect -27684 2526 -27671 2550
rect -27616 2526 -27597 2550
rect -27548 2526 -27523 2550
rect -27480 2526 -27449 2550
rect -27820 2516 -27786 2526
rect -27752 2516 -27718 2526
rect -27684 2516 -27650 2526
rect -27616 2516 -27582 2526
rect -27548 2516 -27514 2526
rect -27480 2516 -27446 2526
rect -27412 2516 -27378 2550
rect -27341 2526 -27310 2550
rect -27267 2526 -27242 2550
rect -27193 2526 -27174 2550
rect -27119 2526 -27106 2550
rect -27344 2516 -27310 2526
rect -27276 2516 -27242 2526
rect -27208 2516 -27174 2526
rect -27140 2516 -27106 2526
rect -27072 2516 -27036 2550
rect 1864 3475 1898 3477
rect 1864 3439 1898 3441
rect 1864 3367 1898 3373
rect 1864 3295 1898 3305
rect 1864 3223 1898 3237
rect 1864 3151 1898 3169
rect 1864 3079 1898 3101
rect 1864 3007 1898 3033
rect 1864 2935 1898 2965
rect 1864 2863 1898 2897
rect 1864 2795 1898 2829
rect 1864 2727 1898 2757
rect 1864 2659 1898 2685
rect 1864 2591 1898 2613
rect 2020 3475 2054 3477
rect 2020 3439 2054 3441
rect 2020 3367 2054 3373
rect 2020 3295 2054 3305
rect 2020 3223 2054 3237
rect 2020 3151 2054 3169
rect 2020 3079 2054 3101
rect 2020 3007 2054 3033
rect 2020 2935 2054 2965
rect 2020 2863 2054 2897
rect 2020 2795 2054 2829
rect 2020 2727 2054 2757
rect 2020 2659 2054 2685
rect 2020 2591 2054 2613
rect 2176 3475 2210 3477
rect 2176 3439 2210 3441
rect 2311 3486 2345 3524
rect 2311 3420 2345 3436
rect 2467 3486 2501 3524
rect 2467 3420 2501 3436
rect 2623 3486 2657 3524
rect 2623 3420 2657 3436
rect 2757 3477 2791 3499
rect 2176 3367 2210 3373
rect 2176 3295 2210 3305
rect 2757 3405 2791 3431
rect 2757 3333 2791 3363
rect 2757 3261 2791 3295
rect 2176 3223 2210 3237
rect 2176 3151 2210 3169
rect 2176 3079 2210 3101
rect 2176 3007 2210 3033
rect 2392 3233 2468 3250
rect 2550 3238 2584 3249
rect 2392 3199 2394 3233
rect 2428 3199 2468 3233
rect 2392 3165 2468 3199
rect 2392 3131 2394 3165
rect 2428 3131 2468 3165
rect 2580 3233 2584 3238
rect 2546 3199 2550 3204
rect 2546 3166 2584 3199
rect 2580 3165 2584 3166
rect 2392 3104 2468 3131
rect 2550 3115 2584 3131
rect 2757 3193 2791 3227
rect 2757 3125 2791 3155
rect 2392 3070 2394 3104
rect 2428 3070 2468 3104
rect 2392 3032 2468 3070
rect 2392 2998 2394 3032
rect 2428 2998 2468 3032
rect 2757 3057 2791 3083
rect 2757 3007 2791 3011
rect 2913 3477 2947 3499
rect 2913 3405 2947 3431
rect 2913 3333 2947 3363
rect 2913 3261 2947 3295
rect 2913 3193 2947 3227
rect 2913 3125 2947 3155
rect 2913 3057 2947 3083
rect 2913 3007 2947 3011
rect 3040 3477 3074 3499
rect 3040 3405 3074 3431
rect 3040 3333 3074 3363
rect 3040 3261 3074 3295
rect 3040 3193 3074 3227
rect 3040 3125 3074 3155
rect 3040 3057 3074 3083
rect 3040 3007 3074 3011
rect 3196 3477 3230 3499
rect 3196 3405 3230 3431
rect 3196 3333 3230 3363
rect 3196 3261 3230 3295
rect 3196 3193 3230 3227
rect 3196 3125 3230 3155
rect 3196 3057 3230 3083
rect 3196 3007 3230 3011
rect 3352 3477 3386 3499
rect 3352 3405 3386 3431
rect 3352 3333 3386 3363
rect 3352 3261 3386 3295
rect 3352 3193 3386 3227
rect 3352 3125 3386 3155
rect 3352 3057 3386 3083
rect 3352 3007 3386 3011
rect 3508 3477 3542 3499
rect 3508 3405 3542 3431
rect 3508 3333 3542 3363
rect 3508 3261 3542 3295
rect 3508 3193 3542 3227
rect 3508 3125 3542 3155
rect 3508 3057 3542 3083
rect 3508 3007 3542 3011
rect 3938 3540 3972 3564
rect 3938 3464 3972 3496
rect 3938 3394 3972 3428
rect 3938 3326 3972 3354
rect 3938 3258 3972 3278
rect 3938 3190 3972 3202
rect 3938 3122 3972 3126
rect 3938 3084 3972 3088
rect 3938 3008 3972 3020
rect 2392 2995 2468 2998
rect 2176 2935 2210 2965
rect 3938 2932 3972 2952
rect 2176 2863 2210 2897
rect 2176 2795 2210 2829
rect 2822 2884 2856 2900
rect 3085 2863 3101 2897
rect 3135 2894 3171 2897
rect 3205 2894 3240 2897
rect 3274 2894 3309 2897
rect 3153 2863 3171 2894
rect 3229 2863 3240 2894
rect 3305 2863 3309 2894
rect 3343 2894 3378 2897
rect 3412 2894 3447 2897
rect 3343 2863 3346 2894
rect 3412 2863 3421 2894
rect 3481 2863 3497 2897
rect 3153 2860 3195 2863
rect 3229 2860 3271 2863
rect 3305 2860 3346 2863
rect 3380 2860 3421 2863
rect 2822 2816 2856 2839
rect 2822 2766 2856 2767
rect 3938 2856 3972 2884
rect 3938 2782 3972 2816
rect 2176 2727 2210 2757
rect 3938 2714 3972 2746
rect 2176 2659 2210 2685
rect 2176 2591 2210 2613
rect 3065 2676 3110 2710
rect 3144 2676 3190 2710
rect 3224 2676 3270 2710
rect 3304 2676 3350 2710
rect 3384 2676 3430 2710
rect 3464 2676 3510 2710
rect 3544 2676 3590 2710
rect 3031 2614 3624 2676
rect 3065 2580 3110 2614
rect 3144 2580 3190 2614
rect 3224 2580 3270 2614
rect 3304 2580 3350 2614
rect 3384 2580 3430 2614
rect 3464 2580 3510 2614
rect 3544 2580 3590 2614
rect 3938 2646 3972 2671
rect 3938 2578 3972 2596
rect -29114 2508 -27036 2516
rect -29148 2474 -29134 2484
rect -29100 2481 -29046 2508
rect -29012 2481 -28958 2508
rect -28924 2481 -28870 2508
rect -28836 2487 -27036 2508
rect -701 2523 -685 2532
rect -651 2523 -590 2532
rect -556 2523 -495 2532
rect -701 2498 -690 2523
rect -651 2498 -617 2523
rect -556 2498 -543 2523
rect -656 2489 -617 2498
rect -583 2489 -543 2498
rect -509 2498 -495 2523
rect -461 2498 -445 2532
rect 248 2524 282 2540
rect 404 2524 438 2540
rect 696 2524 730 2540
rect 852 2524 886 2540
rect 1135 2524 1169 2540
rect 1495 2524 1529 2540
rect -28836 2481 -28189 2487
rect -28155 2481 -28115 2487
rect -28081 2481 -28041 2487
rect -28007 2481 -27967 2487
rect -27933 2481 -27893 2487
rect -27859 2481 -27819 2487
rect -27785 2481 -27745 2487
rect -27711 2481 -27671 2487
rect -27637 2481 -27597 2487
rect -27563 2481 -27523 2487
rect -27489 2481 -27449 2487
rect -27415 2481 -27375 2487
rect -27341 2481 -27301 2487
rect -27267 2481 -27227 2487
rect -27193 2481 -27153 2487
rect -27119 2481 -27036 2487
rect -29100 2474 -29078 2481
rect -29012 2474 -29010 2481
rect -29148 2450 -29078 2474
rect -29114 2447 -29078 2450
rect -29044 2447 -29010 2474
rect -28976 2474 -28958 2481
rect -28976 2447 -28942 2474
rect -28908 2447 -28874 2481
rect -28836 2474 -28806 2481
rect -28840 2447 -28806 2474
rect -28772 2447 -28738 2481
rect -28704 2447 -28670 2481
rect -28636 2447 -28602 2481
rect -28568 2447 -28534 2481
rect -28500 2447 -28466 2481
rect -28432 2447 -28398 2481
rect -28364 2447 -28330 2481
rect -28296 2447 -28262 2481
rect -28228 2447 -28194 2481
rect -28155 2453 -28126 2481
rect -28081 2453 -28058 2481
rect -28007 2453 -27990 2481
rect -27933 2453 -27922 2481
rect -27859 2453 -27854 2481
rect -28160 2447 -28126 2453
rect -28092 2447 -28058 2453
rect -28024 2447 -27990 2453
rect -27956 2447 -27922 2453
rect -27888 2447 -27854 2453
rect -27820 2453 -27819 2481
rect -27752 2453 -27745 2481
rect -27684 2453 -27671 2481
rect -27616 2453 -27597 2481
rect -27548 2453 -27523 2481
rect -27480 2453 -27449 2481
rect -27820 2447 -27786 2453
rect -27752 2447 -27718 2453
rect -27684 2447 -27650 2453
rect -27616 2447 -27582 2453
rect -27548 2447 -27514 2453
rect -27480 2447 -27446 2453
rect -27412 2447 -27378 2481
rect -27341 2453 -27310 2481
rect -27267 2453 -27242 2481
rect -27193 2453 -27174 2481
rect -27119 2453 -27106 2481
rect -27344 2447 -27310 2453
rect -27276 2447 -27242 2453
rect -27208 2447 -27174 2453
rect -27140 2447 -27106 2453
rect -27072 2447 -27036 2481
rect -29114 2435 -27036 2447
rect -29148 2401 -29134 2416
rect -29100 2412 -29046 2435
rect -29012 2412 -28958 2435
rect -28924 2412 -28870 2435
rect -28836 2414 -27036 2435
rect -28836 2412 -28189 2414
rect -28155 2412 -28115 2414
rect -28081 2412 -28041 2414
rect -28007 2412 -27967 2414
rect -27933 2412 -27893 2414
rect -27859 2412 -27819 2414
rect -27785 2412 -27745 2414
rect -27711 2412 -27671 2414
rect -27637 2412 -27597 2414
rect -27563 2412 -27523 2414
rect -27489 2412 -27449 2414
rect -27415 2412 -27375 2414
rect -27341 2412 -27301 2414
rect -27267 2412 -27227 2414
rect -27193 2412 -27153 2414
rect -27119 2412 -27036 2414
rect -29100 2401 -29078 2412
rect -29012 2401 -29010 2412
rect -29148 2382 -29078 2401
rect -29114 2378 -29078 2382
rect -29044 2378 -29010 2401
rect -28976 2401 -28958 2412
rect -28976 2378 -28942 2401
rect -28908 2378 -28874 2412
rect -28836 2401 -28806 2412
rect -28840 2378 -28806 2401
rect -28772 2378 -28738 2412
rect -28704 2378 -28670 2412
rect -28636 2378 -28602 2412
rect -28568 2378 -28534 2412
rect -28500 2378 -28466 2412
rect -28432 2378 -28398 2412
rect -28364 2378 -28330 2412
rect -28296 2378 -28262 2412
rect -28228 2378 -28194 2412
rect -28155 2380 -28126 2412
rect -28081 2380 -28058 2412
rect -28007 2380 -27990 2412
rect -27933 2380 -27922 2412
rect -27859 2380 -27854 2412
rect -28160 2378 -28126 2380
rect -28092 2378 -28058 2380
rect -28024 2378 -27990 2380
rect -27956 2378 -27922 2380
rect -27888 2378 -27854 2380
rect -27820 2380 -27819 2412
rect -27752 2380 -27745 2412
rect -27684 2380 -27671 2412
rect -27616 2380 -27597 2412
rect -27548 2380 -27523 2412
rect -27480 2380 -27449 2412
rect -27820 2378 -27786 2380
rect -27752 2378 -27718 2380
rect -27684 2378 -27650 2380
rect -27616 2378 -27582 2380
rect -27548 2378 -27514 2380
rect -27480 2378 -27446 2380
rect -27412 2378 -27378 2412
rect -27341 2380 -27310 2412
rect -27267 2380 -27242 2412
rect -27193 2380 -27174 2412
rect -27119 2380 -27106 2412
rect -27344 2378 -27310 2380
rect -27276 2378 -27242 2380
rect -27208 2378 -27174 2380
rect -27140 2378 -27106 2380
rect -27072 2378 -27036 2412
rect 281 2469 282 2490
rect 247 2456 282 2469
rect 247 2431 248 2456
rect 281 2406 282 2422
rect 437 2482 438 2490
rect 403 2456 438 2482
rect 403 2444 404 2456
rect 437 2410 438 2422
rect 729 2482 730 2490
rect 695 2456 730 2482
rect 695 2444 696 2456
rect 729 2410 730 2422
rect 885 2482 886 2490
rect 851 2456 886 2482
rect 851 2444 852 2456
rect 885 2410 886 2422
rect 1168 2482 1169 2490
rect 1134 2456 1169 2482
rect 1134 2444 1135 2456
rect 1168 2410 1169 2422
rect 3938 2510 3972 2521
rect 1528 2482 1529 2490
rect 1494 2456 1529 2482
rect 1788 2489 1822 2505
rect 1944 2489 1978 2505
rect 2100 2489 2134 2505
rect 1494 2444 1495 2456
rect 1528 2410 1529 2422
rect 404 2406 438 2410
rect 696 2406 730 2410
rect 852 2406 886 2410
rect 1135 2406 1169 2410
rect 1495 2406 1529 2410
rect 1804 2447 1822 2455
rect 1770 2421 1822 2447
rect 1770 2409 1788 2421
rect -29114 2362 -27036 2378
rect 1804 2375 1822 2387
rect 1977 2447 1978 2455
rect 1943 2421 1978 2447
rect 1943 2409 1944 2421
rect 1977 2375 1978 2387
rect 2133 2447 2134 2455
rect 2099 2421 2134 2447
rect 2099 2409 2100 2421
rect 2133 2375 2134 2387
rect 1788 2371 1822 2375
rect 1944 2371 1978 2375
rect 2100 2371 2134 2375
rect 3938 2442 3972 2446
rect 3938 2374 3972 2408
rect -29148 2328 -29134 2348
rect -29100 2343 -29046 2362
rect -29012 2343 -28958 2362
rect -28924 2343 -28870 2362
rect -28836 2343 -27036 2362
rect -29100 2328 -29078 2343
rect -29012 2328 -29010 2343
rect -29148 2314 -29078 2328
rect -29114 2309 -29078 2314
rect -29044 2309 -29010 2328
rect -28976 2328 -28958 2343
rect -28976 2309 -28942 2328
rect -28908 2309 -28874 2343
rect -28836 2328 -28806 2343
rect -28840 2309 -28806 2328
rect -28772 2309 -28738 2343
rect -28704 2309 -28670 2343
rect -28636 2309 -28602 2343
rect -28568 2309 -28534 2343
rect -28500 2309 -28466 2343
rect -28432 2309 -28398 2343
rect -28364 2309 -28330 2343
rect -28296 2309 -28262 2343
rect -28228 2309 -28194 2343
rect -28160 2341 -28126 2343
rect -28092 2341 -28058 2343
rect -28024 2341 -27990 2343
rect -27956 2341 -27922 2343
rect -27888 2341 -27854 2343
rect -28155 2309 -28126 2341
rect -28081 2309 -28058 2341
rect -28007 2309 -27990 2341
rect -27933 2309 -27922 2341
rect -27859 2309 -27854 2341
rect -27820 2341 -27786 2343
rect -27752 2341 -27718 2343
rect -27684 2341 -27650 2343
rect -27616 2341 -27582 2343
rect -27548 2341 -27514 2343
rect -27480 2341 -27446 2343
rect -27820 2309 -27819 2341
rect -27752 2309 -27745 2341
rect -27684 2309 -27671 2341
rect -27616 2309 -27597 2341
rect -27548 2309 -27523 2341
rect -27480 2309 -27449 2341
rect -27412 2309 -27378 2343
rect -27344 2341 -27310 2343
rect -27276 2341 -27242 2343
rect -27208 2341 -27174 2343
rect -27140 2341 -27106 2343
rect -27341 2309 -27310 2341
rect -27267 2309 -27242 2341
rect -27193 2309 -27174 2341
rect -27119 2309 -27106 2341
rect -27072 2309 -27036 2343
rect -29114 2307 -28189 2309
rect -28155 2307 -28115 2309
rect -28081 2307 -28041 2309
rect -28007 2307 -27967 2309
rect -27933 2307 -27893 2309
rect -27859 2307 -27819 2309
rect -27785 2307 -27745 2309
rect -27711 2307 -27671 2309
rect -27637 2307 -27597 2309
rect -27563 2307 -27523 2309
rect -27489 2307 -27449 2309
rect -27415 2307 -27375 2309
rect -27341 2307 -27301 2309
rect -27267 2307 -27227 2309
rect -27193 2307 -27153 2309
rect -27119 2307 -27036 2309
rect -29114 2289 -27036 2307
rect -29148 2255 -29134 2280
rect -29100 2274 -29046 2289
rect -29012 2274 -28958 2289
rect -28924 2274 -28870 2289
rect -28836 2274 -27036 2289
rect -29100 2255 -29078 2274
rect -29012 2255 -29010 2274
rect -29148 2246 -29078 2255
rect -29114 2240 -29078 2246
rect -29044 2240 -29010 2255
rect -28976 2255 -28958 2274
rect -28976 2240 -28942 2255
rect -28908 2240 -28874 2274
rect -28836 2255 -28806 2274
rect -28840 2240 -28806 2255
rect -28772 2240 -28738 2274
rect -28704 2240 -28670 2274
rect -28636 2240 -28602 2274
rect -28568 2240 -28534 2274
rect -28500 2240 -28466 2274
rect -28432 2240 -28398 2274
rect -28364 2240 -28330 2274
rect -28296 2240 -28262 2274
rect -28228 2240 -28194 2274
rect -28160 2268 -28126 2274
rect -28092 2268 -28058 2274
rect -28024 2268 -27990 2274
rect -27956 2268 -27922 2274
rect -27888 2268 -27854 2274
rect -28155 2240 -28126 2268
rect -28081 2240 -28058 2268
rect -28007 2240 -27990 2268
rect -27933 2240 -27922 2268
rect -27859 2240 -27854 2268
rect -27820 2268 -27786 2274
rect -27752 2268 -27718 2274
rect -27684 2268 -27650 2274
rect -27616 2268 -27582 2274
rect -27548 2268 -27514 2274
rect -27480 2268 -27446 2274
rect -27820 2240 -27819 2268
rect -27752 2240 -27745 2268
rect -27684 2240 -27671 2268
rect -27616 2240 -27597 2268
rect -27548 2240 -27523 2268
rect -27480 2240 -27449 2268
rect -27412 2240 -27378 2274
rect -27344 2268 -27310 2274
rect -27276 2268 -27242 2274
rect -27208 2268 -27174 2274
rect -27140 2268 -27106 2274
rect -27341 2240 -27310 2268
rect -27267 2240 -27242 2268
rect -27193 2240 -27174 2268
rect -27119 2240 -27106 2268
rect -27072 2240 -27036 2274
rect 3938 2306 3972 2340
rect -29114 2234 -28189 2240
rect -28155 2234 -28115 2240
rect -28081 2234 -28041 2240
rect -28007 2234 -27967 2240
rect -27933 2234 -27893 2240
rect -27859 2234 -27819 2240
rect -27785 2234 -27745 2240
rect -27711 2234 -27671 2240
rect -27637 2234 -27597 2240
rect -27563 2234 -27523 2240
rect -27489 2234 -27449 2240
rect -27415 2234 -27375 2240
rect -27341 2234 -27301 2240
rect -27267 2234 -27227 2240
rect -27193 2234 -27153 2240
rect -27119 2234 -27036 2240
rect -29114 2216 -27036 2234
rect -29148 2182 -29134 2212
rect -29100 2205 -29046 2216
rect -29012 2205 -28958 2216
rect -28924 2205 -28870 2216
rect -28836 2205 -27036 2216
rect -29100 2182 -29078 2205
rect -29012 2182 -29010 2205
rect -29148 2178 -29078 2182
rect -29114 2171 -29078 2178
rect -29044 2171 -29010 2182
rect -28976 2182 -28958 2205
rect -28976 2171 -28942 2182
rect -28908 2171 -28874 2205
rect -28836 2182 -28806 2205
rect -28840 2171 -28806 2182
rect -28772 2171 -28738 2205
rect -28704 2171 -28670 2205
rect -28636 2171 -28602 2205
rect -28568 2171 -28534 2205
rect -28500 2171 -28466 2205
rect -28432 2171 -28398 2205
rect -28364 2171 -28330 2205
rect -28296 2171 -28262 2205
rect -28228 2171 -28194 2205
rect -28160 2195 -28126 2205
rect -28092 2195 -28058 2205
rect -28024 2195 -27990 2205
rect -27956 2195 -27922 2205
rect -27888 2195 -27854 2205
rect -28155 2171 -28126 2195
rect -28081 2171 -28058 2195
rect -28007 2171 -27990 2195
rect -27933 2171 -27922 2195
rect -27859 2171 -27854 2195
rect -27820 2195 -27786 2205
rect -27752 2195 -27718 2205
rect -27684 2195 -27650 2205
rect -27616 2195 -27582 2205
rect -27548 2195 -27514 2205
rect -27480 2195 -27446 2205
rect -27820 2171 -27819 2195
rect -27752 2171 -27745 2195
rect -27684 2171 -27671 2195
rect -27616 2171 -27597 2195
rect -27548 2171 -27523 2195
rect -27480 2171 -27449 2195
rect -27412 2171 -27378 2205
rect -27344 2195 -27310 2205
rect -27276 2195 -27242 2205
rect -27208 2195 -27174 2205
rect -27140 2195 -27106 2205
rect -27341 2171 -27310 2195
rect -27267 2171 -27242 2195
rect -27193 2171 -27174 2195
rect -27119 2171 -27106 2195
rect -27072 2171 -27036 2205
rect -29114 2161 -28189 2171
rect -28155 2161 -28115 2171
rect -28081 2161 -28041 2171
rect -28007 2161 -27967 2171
rect -27933 2161 -27893 2171
rect -27859 2161 -27819 2171
rect -27785 2161 -27745 2171
rect -27711 2161 -27671 2171
rect -27637 2161 -27597 2171
rect -27563 2161 -27523 2171
rect -27489 2161 -27449 2171
rect -27415 2161 -27375 2171
rect -27341 2161 -27301 2171
rect -27267 2161 -27227 2171
rect -27193 2161 -27153 2171
rect -27119 2161 -27036 2171
rect -29114 2144 -27036 2161
rect -29148 2143 -27036 2144
rect -29148 2110 -29134 2143
rect -29100 2136 -29046 2143
rect -29012 2136 -28958 2143
rect -28924 2136 -28870 2143
rect -28836 2136 -27036 2143
rect -29100 2109 -29078 2136
rect -29012 2109 -29010 2136
rect -29114 2102 -29078 2109
rect -29044 2102 -29010 2109
rect -28976 2109 -28958 2136
rect -28976 2102 -28942 2109
rect -28908 2102 -28874 2136
rect -28836 2109 -28806 2136
rect -28840 2102 -28806 2109
rect -28772 2102 -28738 2136
rect -28704 2102 -28670 2136
rect -28636 2102 -28602 2136
rect -28568 2102 -28534 2136
rect -28500 2102 -28466 2136
rect -28432 2102 -28398 2136
rect -28364 2102 -28330 2136
rect -28296 2102 -28262 2136
rect -28228 2102 -28194 2136
rect -28160 2122 -28126 2136
rect -28092 2122 -28058 2136
rect -28024 2122 -27990 2136
rect -27956 2122 -27922 2136
rect -27888 2122 -27854 2136
rect -28155 2102 -28126 2122
rect -28081 2102 -28058 2122
rect -28007 2102 -27990 2122
rect -27933 2102 -27922 2122
rect -27859 2102 -27854 2122
rect -27820 2122 -27786 2136
rect -27752 2122 -27718 2136
rect -27684 2122 -27650 2136
rect -27616 2122 -27582 2136
rect -27548 2122 -27514 2136
rect -27480 2122 -27446 2136
rect -27820 2102 -27819 2122
rect -27752 2102 -27745 2122
rect -27684 2102 -27671 2122
rect -27616 2102 -27597 2122
rect -27548 2102 -27523 2122
rect -27480 2102 -27449 2122
rect -27412 2102 -27378 2136
rect -27344 2122 -27310 2136
rect -27276 2122 -27242 2136
rect -27208 2122 -27174 2136
rect -27140 2122 -27106 2136
rect -27341 2102 -27310 2122
rect -27267 2102 -27242 2122
rect -27193 2102 -27174 2122
rect -27119 2102 -27106 2122
rect -27072 2102 -27036 2136
rect -29114 2088 -28189 2102
rect -28155 2088 -28115 2102
rect -28081 2088 -28041 2102
rect -28007 2088 -27967 2102
rect -27933 2088 -27893 2102
rect -27859 2088 -27819 2102
rect -27785 2088 -27745 2102
rect -27711 2088 -27671 2102
rect -27637 2088 -27597 2102
rect -27563 2088 -27523 2102
rect -27489 2088 -27449 2102
rect -27415 2088 -27375 2102
rect -27341 2088 -27301 2102
rect -27267 2088 -27227 2102
rect -27193 2088 -27153 2102
rect -27119 2088 -27036 2102
rect -29114 2076 -27036 2088
rect -29148 2070 -27036 2076
rect -29148 2042 -29134 2070
rect -29100 2067 -29046 2070
rect -29012 2067 -28958 2070
rect -28924 2067 -28870 2070
rect -28836 2067 -27036 2070
rect -29100 2036 -29078 2067
rect -29114 2008 -29078 2036
rect -29148 1997 -29078 2008
rect -29148 1974 -29134 1997
rect -29100 1963 -29078 1997
rect -29114 1940 -29078 1963
rect -29148 1924 -29078 1940
rect -29148 1906 -29134 1924
rect -29100 1890 -29078 1924
rect -29114 1872 -29078 1890
rect -29148 1851 -29078 1872
rect -29148 1838 -29134 1851
rect -29100 1817 -29078 1851
rect -29114 1804 -29078 1817
rect -29148 1778 -29078 1804
rect -29148 1770 -29134 1778
rect -29100 1744 -29078 1778
rect -29114 1736 -29078 1744
rect -29148 1705 -29078 1736
rect -29148 1702 -29134 1705
rect -29100 1671 -29078 1705
rect -29114 1668 -29078 1671
rect -29148 1634 -29078 1668
rect -29114 1632 -29078 1634
rect -29148 1598 -29134 1600
rect -29100 1598 -29078 1632
rect -29148 1566 -29078 1598
rect -29114 1559 -29078 1566
rect -29148 1525 -29134 1532
rect -29100 1525 -29078 1559
rect -29148 1498 -29078 1525
rect -29114 1486 -29078 1498
rect -29148 1452 -29134 1464
rect -29100 1452 -29078 1486
rect -29148 1430 -29078 1452
rect -29114 1413 -29078 1430
rect -29148 1379 -29134 1396
rect -29100 1379 -29078 1413
rect -29148 1362 -29078 1379
rect -29114 1340 -29078 1362
rect -29148 1306 -29134 1328
rect -29100 1306 -29078 1340
rect -29148 1294 -29078 1306
rect -29114 1267 -29078 1294
rect -29148 1233 -29134 1260
rect -29100 1233 -29078 1267
rect -29148 1226 -29078 1233
rect -29114 1194 -29078 1226
rect -29148 1160 -29134 1192
rect -29100 1160 -29078 1194
rect -29148 1158 -29078 1160
rect -29114 1124 -29078 1158
rect -29148 1121 -29078 1124
rect -29148 1090 -29134 1121
rect -29100 1087 -29078 1121
rect -29114 1056 -29078 1087
rect -29148 1048 -29078 1056
rect -29148 1022 -29134 1048
rect -29100 1014 -29078 1048
rect -29114 988 -29078 1014
rect -29148 975 -29078 988
rect -29148 954 -29134 975
rect -29100 941 -29078 975
rect -29114 920 -29078 941
rect -29148 902 -29078 920
rect -29148 886 -29134 902
rect -29100 868 -29078 902
rect -29114 852 -29078 868
rect -29148 829 -29078 852
rect -29148 818 -29134 829
rect -29100 795 -29078 829
rect -29114 784 -29078 795
rect -29148 756 -29078 784
rect -29148 750 -29134 756
rect -29100 722 -29078 756
rect -29114 716 -29078 722
rect -29148 683 -29078 716
rect -29148 682 -29134 683
rect -29100 649 -29078 683
rect -29114 648 -29078 649
rect -29148 614 -29078 648
rect -29114 610 -29078 614
rect -29148 576 -29134 580
rect -29100 576 -29078 610
rect -29148 546 -29078 576
rect -29114 537 -29078 546
rect -29148 503 -29134 512
rect -29100 503 -29078 537
rect -29148 478 -29078 503
rect -29114 464 -29078 478
rect -29148 430 -29134 444
rect -29100 430 -29078 464
rect -29148 410 -29078 430
rect -29114 391 -29078 410
rect -29148 357 -29134 376
rect -29100 357 -29078 391
rect -29148 342 -29078 357
rect -29114 318 -29078 342
rect -29148 284 -29134 308
rect -29100 284 -29078 318
rect -29148 274 -29078 284
rect -29114 245 -29078 274
rect -29148 211 -29134 240
rect -29100 211 -29078 245
rect -29148 206 -29078 211
rect -29114 172 -29078 206
rect -29148 138 -29134 172
rect -29100 138 -29078 172
rect -29114 104 -29078 138
rect -29148 99 -29078 104
rect -29148 70 -29134 99
rect -29100 65 -29078 99
rect -29114 36 -29078 65
rect -29148 26 -29078 36
rect -29148 2 -29134 26
rect -29100 -8 -29078 26
rect -29114 -32 -29078 -8
rect -29148 -47 -29078 -32
rect -29148 -66 -29134 -47
rect -29100 -81 -29078 -47
rect -29114 -100 -29078 -81
rect -29148 -120 -29078 -100
rect -29148 -134 -29134 -120
rect -29100 -154 -29078 -120
rect -29114 -168 -29078 -154
rect -29148 -193 -29078 -168
rect -29148 -202 -29134 -193
rect -29100 -227 -29078 -193
rect -29114 -236 -29078 -227
rect -29148 -266 -29078 -236
rect -29148 -270 -29134 -266
rect -29100 -300 -29078 -266
rect -29114 -304 -29078 -300
rect -29148 -338 -29078 -304
rect -29114 -339 -29078 -338
rect -29148 -373 -29134 -372
rect -29100 -373 -29078 -339
rect -29148 -406 -29078 -373
rect -29114 -412 -29078 -406
rect -29148 -446 -29134 -440
rect -29100 -446 -29078 -412
rect -29148 -474 -29078 -446
rect -29114 -485 -29078 -474
rect -29148 -519 -29134 -508
rect -29100 -519 -29078 -485
rect -29148 -542 -29078 -519
rect -29114 -558 -29078 -542
rect -29148 -592 -29134 -576
rect -29100 -592 -29078 -558
rect -29148 -610 -29078 -592
rect -29114 -631 -29078 -610
rect -29148 -665 -29134 -644
rect -29100 -665 -29078 -631
rect -29148 -678 -29078 -665
rect -29114 -704 -29078 -678
rect -29148 -738 -29134 -712
rect -29100 -738 -29078 -704
rect -29148 -746 -29078 -738
rect -29114 -777 -29078 -746
rect -29148 -811 -29134 -780
rect -29100 -811 -29078 -777
rect -29148 -814 -29078 -811
rect -29114 -848 -29078 -814
rect -29148 -849 -29078 -848
rect -29148 -882 -29134 -849
rect -29100 -883 -29078 -849
rect -29114 -916 -29078 -883
rect -29148 -921 -29078 -916
rect -29148 -950 -29134 -921
rect -29100 -955 -29078 -921
rect -29114 -984 -29078 -955
rect -29148 -993 -29078 -984
rect -29148 -1018 -29134 -993
rect -29100 -1027 -29078 -993
rect -29114 -1052 -29078 -1027
rect -29148 -1065 -29078 -1052
rect -29148 -1086 -29134 -1065
rect -29100 -1099 -29078 -1065
rect -29114 -1120 -29078 -1099
rect -29148 -1137 -29078 -1120
rect -29148 -1154 -29134 -1137
rect -29100 -1171 -29078 -1137
rect -29114 -1188 -29078 -1171
rect -29148 -1209 -29078 -1188
rect -29148 -1222 -29134 -1209
rect -29100 -1243 -29078 -1209
rect -29114 -1256 -29078 -1243
rect -29148 -1281 -29078 -1256
rect -29148 -1290 -29134 -1281
rect -29100 -1315 -29078 -1281
rect -29114 -1324 -29078 -1315
rect -29148 -1353 -29078 -1324
rect -29148 -1358 -29134 -1353
rect -29100 -1387 -29078 -1353
rect -29114 -1392 -29078 -1387
rect -29148 -1425 -29078 -1392
rect -29148 -1426 -29134 -1425
rect -29100 -1459 -29078 -1425
rect -29114 -1460 -29078 -1459
rect -29148 -1494 -29078 -1460
rect -29114 -1497 -29078 -1494
rect -29148 -1531 -29134 -1528
rect -29100 -1531 -29078 -1497
rect -29148 -1562 -29078 -1531
rect -29114 -1569 -29078 -1562
rect -29148 -1603 -29134 -1596
rect -29100 -1603 -29078 -1569
rect -29148 -1630 -29078 -1603
rect -29114 -1641 -29078 -1630
rect -29148 -1675 -29134 -1664
rect -29100 -1675 -29078 -1641
rect -29148 -1698 -29078 -1675
rect -29114 -1713 -29078 -1698
rect -29148 -1747 -29134 -1732
rect -29100 -1747 -29078 -1713
rect -29148 -1766 -29078 -1747
rect -29114 -1785 -29078 -1766
rect -29148 -1819 -29134 -1800
rect -29100 -1819 -29078 -1785
rect -29148 -1834 -29078 -1819
rect -29114 -1857 -29078 -1834
rect -29148 -1891 -29134 -1868
rect -29100 -1891 -29078 -1857
rect -29148 -1902 -29078 -1891
rect -29114 -1929 -29078 -1902
rect -29148 -1963 -29134 -1936
rect -29100 -1963 -29078 -1929
rect -29148 -1970 -29078 -1963
rect -29114 -2001 -29078 -1970
rect -29148 -2035 -29134 -2004
rect -29100 -2035 -29078 -2001
rect -29148 -2038 -29078 -2035
rect -29114 -2072 -29078 -2038
rect -29148 -2073 -29078 -2072
rect -29148 -2106 -29134 -2073
rect -29100 -2107 -29078 -2073
rect -29114 -2140 -29078 -2107
rect -29148 -2145 -29078 -2140
rect -29148 -2174 -29134 -2145
rect -29100 -2179 -29078 -2145
rect -29114 -2208 -29078 -2179
rect -29148 -2217 -29078 -2208
rect -29148 -2242 -29134 -2217
rect -29100 -2251 -29078 -2217
rect -29114 -2276 -29078 -2251
rect -29148 -2289 -29078 -2276
rect -29148 -2310 -29134 -2289
rect -29100 -2323 -29078 -2289
rect -29114 -2344 -29078 -2323
rect -29148 -2361 -29078 -2344
rect -29148 -2378 -29134 -2361
rect -29100 -2395 -29078 -2361
rect -29114 -2412 -29078 -2395
rect -29148 -2433 -29078 -2412
rect -29148 -2446 -29134 -2433
rect -29100 -2467 -29078 -2433
rect -29114 -2480 -29078 -2467
rect -29148 -2505 -29078 -2480
rect -29148 -2514 -29134 -2505
rect -29100 -2539 -29078 -2505
rect -29114 -2548 -29078 -2539
rect -29148 -2577 -29078 -2548
rect -29148 -2582 -29134 -2577
rect -29100 -2611 -29078 -2577
rect -29114 -2616 -29078 -2611
rect -29148 -2649 -29078 -2616
rect -29148 -2650 -29134 -2649
rect -29100 -2683 -29078 -2649
rect -29114 -2684 -29078 -2683
rect -29148 -2718 -29078 -2684
rect -29114 -2721 -29078 -2718
rect -29148 -2755 -29134 -2752
rect -29100 -2755 -29078 -2721
rect -29148 -2786 -29078 -2755
rect -29114 -2793 -29078 -2786
rect -29148 -2827 -29134 -2820
rect -29100 -2827 -29078 -2793
rect -29148 -2854 -29078 -2827
rect -29114 -2865 -29078 -2854
rect -29148 -2899 -29134 -2888
rect -29100 -2899 -29078 -2865
rect -29148 -2922 -29078 -2899
rect -29114 -2937 -29078 -2922
rect -29148 -2971 -29134 -2956
rect -29100 -2971 -29078 -2937
rect -29148 -2990 -29078 -2971
rect -29114 -3009 -29078 -2990
rect -29148 -3043 -29134 -3024
rect -29100 -3043 -29078 -3009
rect -29148 -3058 -29078 -3043
rect -29114 -3081 -29078 -3058
rect -29148 -3115 -29134 -3092
rect -29100 -3115 -29078 -3081
rect -29148 -3126 -29078 -3115
rect -29114 -3153 -29078 -3126
rect -29148 -3187 -29134 -3160
rect -29100 -3187 -29078 -3153
rect -29148 -3194 -29078 -3187
rect -29114 -3225 -29078 -3194
rect -29148 -3259 -29134 -3228
rect -29100 -3259 -29078 -3225
rect -29148 -3262 -29078 -3259
rect -29114 -3296 -29078 -3262
rect -29148 -3297 -29078 -3296
rect -29148 -3330 -29134 -3297
rect -29100 -3331 -29078 -3297
rect -29114 -3364 -29078 -3331
rect -29148 -3369 -29078 -3364
rect -29148 -3398 -29134 -3369
rect -29100 -3403 -29078 -3369
rect -29114 -3432 -29078 -3403
rect -29148 -3441 -29078 -3432
rect -29148 -3466 -29134 -3441
rect -29100 -3475 -29078 -3441
rect -29114 -3500 -29078 -3475
rect -29148 -3513 -29078 -3500
rect -29148 -3534 -29134 -3513
rect -29100 -3547 -29078 -3513
rect -29114 -3568 -29078 -3547
rect -29148 -3585 -29078 -3568
rect -29148 -3602 -29134 -3585
rect -29100 -3619 -29078 -3585
rect -29114 -3636 -29078 -3619
rect -29148 -3657 -29078 -3636
rect -29148 -3670 -29134 -3657
rect -29100 -3691 -29078 -3657
rect -29114 -3704 -29078 -3691
rect -29148 -3729 -29078 -3704
rect -29148 -3738 -29134 -3729
rect -29100 -3763 -29078 -3729
rect -29114 -3772 -29078 -3763
rect -29148 -3801 -29078 -3772
rect -29148 -3806 -29134 -3801
rect -29100 -3835 -29078 -3801
rect -29114 -3840 -29078 -3835
rect -29148 -3873 -29078 -3840
rect -29148 -3874 -29134 -3873
rect -29100 -3907 -29078 -3873
rect -29114 -3908 -29078 -3907
rect -29148 -3942 -29078 -3908
rect -29114 -3945 -29078 -3942
rect -29148 -3979 -29134 -3976
rect -29100 -3979 -29078 -3945
rect -29148 -4010 -29078 -3979
rect -29114 -4017 -29078 -4010
rect -29148 -4051 -29134 -4044
rect -29100 -4051 -29078 -4017
rect -29148 -4078 -29078 -4051
rect -29114 -4089 -29078 -4078
rect -29148 -4123 -29134 -4112
rect -29100 -4123 -29078 -4089
rect -29148 -4146 -29078 -4123
rect -29114 -4161 -29078 -4146
rect -29148 -4195 -29134 -4180
rect -29100 -4195 -29078 -4161
rect -29148 -4214 -29078 -4195
rect -29114 -4233 -29078 -4214
rect -29148 -4267 -29134 -4248
rect -29100 -4267 -29078 -4233
rect -29148 -4282 -29078 -4267
rect -29114 -4305 -29078 -4282
rect -29148 -4339 -29134 -4316
rect -29100 -4339 -29078 -4305
rect -29148 -4350 -29078 -4339
rect -29114 -4377 -29078 -4350
rect -29148 -4411 -29134 -4384
rect -29100 -4411 -29078 -4377
rect -29148 -4418 -29078 -4411
rect -29114 -4449 -29078 -4418
rect -29148 -4483 -29134 -4452
rect -29100 -4483 -29078 -4449
rect -29148 -4486 -29078 -4483
rect -29114 -4520 -29078 -4486
rect -29148 -4521 -29078 -4520
rect -29148 -4554 -29134 -4521
rect -29100 -4555 -29078 -4521
rect -29114 -4588 -29078 -4555
rect -29148 -4593 -29078 -4588
rect -29148 -4622 -29134 -4593
rect -29100 -4627 -29078 -4593
rect -29114 -4656 -29078 -4627
rect -29148 -4665 -29078 -4656
rect -29148 -4690 -29134 -4665
rect -29100 -4699 -29078 -4665
rect -29114 -4724 -29078 -4699
rect -29148 -4737 -29078 -4724
rect -29148 -4758 -29134 -4737
rect -29100 -4771 -29078 -4737
rect -29114 -4792 -29078 -4771
rect -29148 -4809 -29078 -4792
rect -29148 -4826 -29134 -4809
rect -29100 -4843 -29078 -4809
rect -29114 -4860 -29078 -4843
rect -29148 -4881 -29078 -4860
rect -29148 -4894 -29134 -4881
rect -29100 -4915 -29078 -4881
rect -29114 -4928 -29078 -4915
rect -29148 -4953 -29078 -4928
rect -29148 -4962 -29134 -4953
rect -29100 -4987 -29078 -4953
rect -29114 -4996 -29078 -4987
rect -29148 -5025 -29078 -4996
rect -29148 -5030 -29134 -5025
rect -29100 -5059 -29078 -5025
rect -29114 -5064 -29078 -5059
rect -29148 -5097 -29078 -5064
rect -29148 -5098 -29134 -5097
rect -29100 -5131 -29078 -5097
rect -29114 -5132 -29078 -5131
rect -29148 -5166 -29078 -5132
rect -29114 -5169 -29078 -5166
rect -29148 -5203 -29134 -5200
rect -29100 -5203 -29078 -5169
rect -29148 -5234 -29078 -5203
rect -29114 -5241 -29078 -5234
rect -29148 -5275 -29134 -5268
rect -29100 -5275 -29078 -5241
rect -29148 -5302 -29078 -5275
rect -29114 -5313 -29078 -5302
rect -29148 -5347 -29134 -5336
rect -29100 -5347 -29078 -5313
rect -29148 -5370 -29078 -5347
rect -29114 -5385 -29078 -5370
rect -29148 -5419 -29134 -5404
rect -29100 -5419 -29078 -5385
rect -29148 -5438 -29078 -5419
rect -29114 -5457 -29078 -5438
rect -29148 -5491 -29134 -5472
rect -29100 -5491 -29078 -5457
rect -29148 -5506 -29078 -5491
rect -29114 -5529 -29078 -5506
rect -29148 -5563 -29134 -5540
rect -29100 -5563 -29078 -5529
rect -29148 -5574 -29078 -5563
rect -29114 -5601 -29078 -5574
rect -29148 -5635 -29134 -5608
rect -29100 -5635 -29078 -5601
rect -29148 -5642 -29078 -5635
rect -29114 -5673 -29078 -5642
rect -29148 -5707 -29134 -5676
rect -29100 -5707 -29078 -5673
rect -29148 -5710 -29078 -5707
rect -29114 -5744 -29078 -5710
rect -29148 -5745 -29078 -5744
rect -29148 -5778 -29134 -5745
rect -29100 -5779 -29078 -5745
rect -29114 -5812 -29078 -5779
rect -29148 -5817 -29078 -5812
rect -29148 -5846 -29134 -5817
rect -29100 -5851 -29078 -5817
rect -29114 -5880 -29078 -5851
rect -29148 -5889 -29078 -5880
rect -29148 -5914 -29134 -5889
rect -29100 -5923 -29078 -5889
rect -29114 -5948 -29078 -5923
rect -29148 -5961 -29078 -5948
rect -29148 -5982 -29134 -5961
rect -29100 -5995 -29078 -5961
rect -29114 -6016 -29078 -5995
rect -29148 -6033 -29078 -6016
rect -29148 -6050 -29134 -6033
rect -29100 -6067 -29078 -6033
rect -29114 -6084 -29078 -6067
rect -29148 -6105 -29078 -6084
rect -29148 -6118 -29134 -6105
rect -29100 -6139 -29078 -6105
rect -29114 -6152 -29078 -6139
rect -29148 -6177 -29078 -6152
rect -29148 -6186 -29134 -6177
rect -29100 -6211 -29078 -6177
rect -29114 -6220 -29078 -6211
rect -29148 -6249 -29078 -6220
rect -29148 -6254 -29134 -6249
rect -29100 -6283 -29078 -6249
rect -29114 -6288 -29078 -6283
rect -29148 -6321 -29078 -6288
rect -29148 -6322 -29134 -6321
rect -29100 -6355 -29078 -6321
rect -29114 -6356 -29078 -6355
rect -29148 -6390 -29078 -6356
rect -29114 -6393 -29078 -6390
rect -29148 -6427 -29134 -6424
rect -29100 -6427 -29078 -6393
rect -29148 -6458 -29078 -6427
rect -29114 -6465 -29078 -6458
rect -29148 -6499 -29134 -6492
rect -29100 -6499 -29078 -6465
rect -29148 -6526 -29078 -6499
rect -29114 -6537 -29078 -6526
rect -29148 -6571 -29134 -6560
rect -29100 -6571 -29078 -6537
rect -29148 -6594 -29078 -6571
rect -29114 -6609 -29078 -6594
rect -29148 -6643 -29134 -6628
rect -29100 -6643 -29078 -6609
rect -29148 -6662 -29078 -6643
rect -29114 -6681 -29078 -6662
rect -29148 -6715 -29134 -6696
rect -29100 -6715 -29078 -6681
rect -29148 -6730 -29078 -6715
rect -29114 -6753 -29078 -6730
rect -29148 -6787 -29134 -6764
rect -29100 -6787 -29078 -6753
rect -29148 -6798 -29078 -6787
rect -29114 -6825 -29078 -6798
rect -29148 -6859 -29134 -6832
rect -29100 -6859 -29078 -6825
rect -29148 -6866 -29078 -6859
rect -29114 -6897 -29078 -6866
rect -29148 -6931 -29134 -6900
rect -29100 -6931 -29078 -6897
rect -29148 -6934 -29078 -6931
rect -29114 -6968 -29078 -6934
rect -29148 -6969 -29078 -6968
rect -29148 -7002 -29134 -6969
rect -29100 -7003 -29078 -6969
rect -29114 -7036 -29078 -7003
rect -29148 -7041 -29078 -7036
rect -29148 -7070 -29134 -7041
rect -29100 -7075 -29078 -7041
rect -29114 -7104 -29078 -7075
rect -29148 -7113 -29078 -7104
rect -29148 -7138 -29134 -7113
rect -29100 -7147 -29078 -7113
rect -29114 -7172 -29078 -7147
rect -29148 -7185 -29078 -7172
rect -29148 -7206 -29134 -7185
rect -29100 -7219 -29078 -7185
rect -29114 -7240 -29078 -7219
rect -29148 -7257 -29078 -7240
rect -29148 -7274 -29134 -7257
rect -29100 -7291 -29078 -7257
rect -29114 -7308 -29078 -7291
rect -29148 -7329 -29078 -7308
rect -29148 -7342 -29134 -7329
rect -29100 -7363 -29078 -7329
rect -29114 -7376 -29078 -7363
rect -29148 -7401 -29078 -7376
rect -29148 -7410 -29134 -7401
rect -29100 -7435 -29078 -7401
rect -29114 -7444 -29078 -7435
rect -29148 -7473 -29078 -7444
rect -29148 -7478 -29134 -7473
rect -29100 -7507 -29078 -7473
rect -29114 -7512 -29078 -7507
rect -29148 -7545 -29078 -7512
rect -29148 -7546 -29134 -7545
rect -29100 -7579 -29078 -7545
rect -29114 -7580 -29078 -7579
rect -29148 -7614 -29078 -7580
rect -29114 -7617 -29078 -7614
rect -29148 -7651 -29134 -7648
rect -29100 -7651 -29078 -7617
rect -29148 -7682 -29078 -7651
rect -29114 -7689 -29078 -7682
rect -29148 -7723 -29134 -7716
rect -29100 -7723 -29078 -7689
rect -29148 -7750 -29078 -7723
rect -29114 -7761 -29078 -7750
rect -29148 -7795 -29134 -7784
rect -29100 -7795 -29078 -7761
rect -29148 -7818 -29078 -7795
rect -29114 -7833 -29078 -7818
rect -29148 -7867 -29134 -7852
rect -29100 -7867 -29078 -7833
rect -29148 -7886 -29078 -7867
rect -29114 -7905 -29078 -7886
rect -29148 -7939 -29134 -7920
rect -29100 -7939 -29078 -7905
rect -29148 -7954 -29078 -7939
rect -29114 -7977 -29078 -7954
rect -29148 -8011 -29134 -7988
rect -29100 -8011 -29078 -7977
rect -29148 -8022 -29078 -8011
rect -29114 -8049 -29078 -8022
rect -29148 -8083 -29134 -8056
rect -29100 -8083 -29078 -8049
rect -29148 -8090 -29078 -8083
rect -29114 -8121 -29078 -8090
rect -29148 -8155 -29134 -8124
rect -29100 -8155 -29078 -8121
rect -29148 -8158 -29078 -8155
rect -29114 -8192 -29078 -8158
rect -29148 -8193 -29078 -8192
rect -29148 -8226 -29134 -8193
rect -29100 -8227 -29078 -8193
rect -29114 -8260 -29078 -8227
rect -29148 -8265 -29078 -8260
rect -29148 -8294 -29134 -8265
rect -29100 -8299 -29078 -8265
rect -29114 -8328 -29078 -8299
rect -29148 -8337 -29078 -8328
rect -29148 -8362 -29134 -8337
rect -29100 -8371 -29078 -8337
rect -29114 -8396 -29078 -8371
rect -29148 -8409 -29078 -8396
rect -29148 -8430 -29134 -8409
rect -29100 -8443 -29078 -8409
rect -29114 -8464 -29078 -8443
rect -29148 -8481 -29078 -8464
rect -29148 -8498 -29134 -8481
rect -29100 -8515 -29078 -8481
rect -29114 -8532 -29078 -8515
rect -29148 -8553 -29078 -8532
rect -29148 -8566 -29134 -8553
rect -29100 -8587 -29078 -8553
rect -32352 -8678 -32315 -8640
rect -31669 -8643 -31632 -8609
rect -31669 -8677 -31598 -8643
rect -32352 -8712 -32344 -8678
rect -31669 -8711 -31632 -8677
rect -32352 -8750 -32315 -8712
rect -31669 -8745 -31598 -8711
rect -31528 -8659 -31512 -8625
rect -31478 -8659 -31462 -8625
rect -31528 -8685 -31462 -8659
rect -31528 -8731 -31512 -8685
rect -31478 -8731 -31462 -8685
rect -29284 -8627 -29268 -8593
rect -29234 -8627 -29218 -8593
rect -29284 -8665 -29218 -8627
rect -29284 -8731 -29268 -8665
rect -29234 -8731 -29218 -8665
rect -29114 -8600 -29078 -8587
rect -29148 -8625 -29078 -8600
rect -29148 -8634 -29134 -8625
rect -29100 -8659 -29078 -8625
rect -29114 -8668 -29078 -8659
rect -29148 -8697 -29078 -8668
rect -29148 -8702 -29134 -8697
rect -29100 -8731 -29078 -8697
rect -32352 -8784 -32344 -8750
rect -31669 -8779 -31632 -8745
rect -32352 -8822 -32315 -8784
rect -31669 -8813 -31598 -8779
rect -29114 -8736 -29078 -8731
rect -29148 -8769 -29078 -8736
rect -29148 -8803 -29134 -8769
rect -29100 -8803 -29078 -8769
rect -29148 -8813 -29078 -8803
rect -32352 -8856 -32344 -8822
rect -31669 -8847 -31528 -8813
rect -31494 -8847 -31460 -8813
rect -31426 -8847 -31392 -8813
rect -31358 -8847 -31324 -8813
rect -31290 -8847 -31256 -8813
rect -31222 -8847 -31188 -8813
rect -31154 -8847 -31120 -8813
rect -31086 -8847 -31052 -8813
rect -31018 -8847 -30984 -8813
rect -30950 -8847 -30916 -8813
rect -30882 -8847 -30848 -8813
rect -30814 -8847 -30780 -8813
rect -30746 -8847 -30712 -8813
rect -30678 -8847 -30644 -8813
rect -30610 -8847 -30576 -8813
rect -30542 -8847 -30508 -8813
rect -30474 -8847 -30440 -8813
rect -30406 -8847 -30372 -8813
rect -30338 -8847 -30304 -8813
rect -30270 -8847 -30236 -8813
rect -30202 -8847 -30168 -8813
rect -30134 -8847 -30100 -8813
rect -30066 -8847 -30032 -8813
rect -29998 -8847 -29964 -8813
rect -29930 -8847 -29896 -8813
rect -29862 -8847 -29828 -8813
rect -29794 -8847 -29760 -8813
rect -29726 -8847 -29692 -8813
rect -29658 -8847 -29624 -8813
rect -29590 -8847 -29556 -8813
rect -29522 -8847 -29488 -8813
rect -29454 -8847 -29420 -8813
rect -29386 -8847 -29352 -8813
rect -29318 -8847 -29284 -8813
rect -29250 -8847 -29216 -8813
rect -29182 -8841 -29078 -8813
rect -29182 -8847 -29134 -8841
rect -32352 -8918 -32315 -8856
rect -31669 -8875 -29134 -8847
rect -29100 -8847 -29078 -8841
rect -27072 -8847 -27036 2067
rect 244 2169 278 2191
rect 244 2097 278 2123
rect 244 2039 278 2055
rect 1333 2235 1413 2269
rect 1299 2197 1447 2235
rect 2186 2205 2224 2239
rect 3938 2238 3972 2272
rect 4125 3619 4207 3653
rect 4241 3619 4290 3653
rect 4327 3619 4361 3653
rect 4407 3619 4429 3653
rect 4490 3619 4563 3653
rect 4125 3581 4159 3619
rect 4528 3585 4563 3619
rect 4528 3579 4529 3585
rect 4125 3513 4159 3547
rect 4125 3445 4159 3471
rect 4125 3377 4159 3395
rect 4125 3309 4159 3319
rect 4125 3241 4159 3243
rect 4125 3201 4159 3207
rect 4125 3125 4159 3139
rect 4125 3049 4159 3071
rect 4125 2973 4159 3003
rect 4125 2901 4159 2935
rect 4125 2833 4159 2863
rect 4125 2765 4159 2787
rect 4125 2697 4159 2711
rect 4125 2629 4159 2635
rect 4125 2593 4159 2595
rect 4244 3477 4278 3499
rect 4244 3405 4278 3431
rect 4244 3333 4278 3363
rect 4244 3261 4278 3295
rect 4244 3193 4278 3227
rect 4244 3125 4278 3155
rect 4244 3057 4278 3083
rect 4244 2989 4278 3011
rect 4244 2921 4278 2939
rect 4244 2853 4278 2867
rect 4244 2785 4278 2795
rect 4244 2717 4278 2723
rect 4244 2649 4278 2651
rect 4244 2613 4278 2615
rect 4400 3477 4434 3499
rect 4400 3405 4434 3431
rect 4400 3333 4434 3363
rect 4400 3261 4434 3295
rect 4400 3193 4434 3227
rect 4400 3125 4434 3155
rect 4400 3057 4434 3083
rect 4400 2989 4434 3011
rect 4400 2921 4434 2939
rect 4400 2853 4434 2867
rect 4400 2785 4434 2795
rect 4400 2717 4434 2723
rect 4400 2649 4434 2651
rect 4400 2613 4434 2615
rect 4562 3545 4563 3551
rect 4528 3517 4563 3545
rect 4528 3505 4529 3517
rect 4562 3471 4563 3483
rect 4528 3449 4563 3471
rect 4528 3431 4529 3449
rect 4562 3397 4563 3415
rect 4528 3381 4563 3397
rect 4528 3357 4529 3381
rect 4562 3323 4563 3347
rect 4528 3313 4563 3323
rect 4528 3283 4529 3313
rect 4562 3249 4563 3279
rect 4528 3245 4563 3249
rect 4528 3211 4529 3245
rect 4528 3209 4563 3211
rect 4562 3177 4563 3209
rect 4528 3143 4529 3175
rect 4528 3135 4563 3143
rect 4562 3109 4563 3135
rect 4528 3075 4529 3101
rect 4528 3061 4563 3075
rect 4562 3041 4563 3061
rect 4528 3007 4529 3027
rect 4528 2987 4563 3007
rect 4562 2973 4563 2987
rect 4528 2939 4529 2953
rect 4528 2912 4563 2939
rect 4562 2905 4563 2912
rect 4528 2871 4529 2878
rect 4528 2837 4563 2871
rect 4528 2769 4563 2803
rect 4528 2762 4529 2769
rect 4562 2728 4563 2735
rect 4528 2701 4563 2728
rect 4528 2687 4529 2701
rect 4562 2653 4563 2667
rect 4528 2633 4563 2653
rect 4528 2612 4529 2633
rect 4125 2517 4159 2527
rect 4562 2578 4563 2599
rect 4528 2565 4563 2578
rect 4528 2537 4529 2565
rect 4324 2489 4358 2505
rect 4125 2441 4159 2459
rect 4125 2365 4159 2391
rect 4357 2447 4358 2455
rect 4323 2421 4358 2447
rect 4323 2409 4324 2421
rect 4357 2375 4358 2387
rect 4324 2371 4358 2375
rect 4562 2503 4563 2531
rect 4528 2497 4563 2503
rect 4528 2463 4529 2497
rect 4528 2462 4563 2463
rect 4562 2429 4563 2462
rect 4528 2395 4529 2428
rect 4528 2387 4563 2395
rect 4562 2361 4563 2387
rect 4125 2289 4159 2323
rect 4529 2289 4563 2327
rect 4125 2255 4197 2289
rect 4231 2255 4257 2289
rect 4320 2255 4325 2289
rect 4359 2255 4393 2289
rect 4427 2255 4461 2289
rect 4495 2255 4563 2289
rect 4752 3644 4802 3669
rect 4836 3644 4886 3669
rect 4920 3644 4942 3669
rect 5738 3772 5772 3806
rect 5738 3704 5772 3724
rect 4718 3634 4942 3644
rect 4718 3603 4723 3634
rect 4757 3603 4815 3634
rect 4849 3603 4907 3634
rect 4757 3600 4802 3603
rect 4849 3600 4886 3603
rect 4941 3600 4942 3634
rect 4752 3569 4802 3600
rect 4836 3569 4886 3600
rect 4920 3569 4942 3600
rect 4718 3565 4942 3569
rect 4718 3531 4723 3565
rect 4757 3531 4815 3565
rect 4849 3531 4907 3565
rect 4941 3531 4942 3565
rect 4718 3528 4942 3531
rect 4752 3496 4802 3528
rect 4836 3496 4886 3528
rect 4920 3496 4942 3528
rect 4757 3494 4802 3496
rect 4849 3494 4886 3496
rect 4718 3462 4723 3494
rect 4757 3462 4815 3494
rect 4849 3462 4907 3494
rect 4941 3462 4942 3496
rect 4718 3453 4942 3462
rect 4752 3427 4802 3453
rect 4836 3427 4886 3453
rect 4920 3427 4942 3453
rect 4757 3419 4802 3427
rect 4849 3419 4886 3427
rect 4718 3393 4723 3419
rect 4757 3393 4815 3419
rect 4849 3393 4907 3419
rect 4941 3393 4942 3427
rect 4718 3378 4942 3393
rect 4752 3358 4802 3378
rect 4836 3358 4886 3378
rect 4920 3358 4942 3378
rect 4757 3344 4802 3358
rect 4849 3344 4886 3358
rect 4718 3324 4723 3344
rect 4757 3324 4815 3344
rect 4849 3324 4907 3344
rect 4941 3324 4942 3358
rect 4718 3303 4942 3324
rect 4752 3289 4802 3303
rect 4836 3289 4886 3303
rect 4920 3289 4942 3303
rect 4757 3269 4802 3289
rect 4849 3269 4886 3289
rect 4718 3255 4723 3269
rect 4757 3255 4815 3269
rect 4849 3255 4907 3269
rect 4941 3255 4942 3289
rect 4718 3228 4942 3255
rect 4752 3220 4802 3228
rect 4836 3220 4886 3228
rect 4920 3220 4942 3228
rect 4757 3194 4802 3220
rect 4849 3194 4886 3220
rect 4718 3186 4723 3194
rect 4757 3186 4815 3194
rect 4849 3186 4907 3194
rect 4941 3186 4942 3220
rect 4718 3153 4942 3186
rect 4752 3150 4802 3153
rect 4836 3150 4886 3153
rect 4920 3150 4942 3153
rect 4757 3119 4802 3150
rect 4849 3119 4886 3150
rect 4718 3116 4723 3119
rect 4757 3116 4815 3119
rect 4849 3116 4907 3119
rect 4941 3116 4942 3150
rect 4718 3080 4942 3116
rect 4718 3078 4723 3080
rect 4757 3078 4815 3080
rect 4849 3078 4907 3080
rect 4757 3046 4802 3078
rect 4849 3046 4886 3078
rect 4941 3046 4942 3080
rect 4752 3044 4802 3046
rect 4836 3044 4886 3046
rect 4920 3044 4942 3046
rect 4718 3010 4942 3044
rect 4718 3003 4723 3010
rect 4757 3003 4815 3010
rect 4849 3003 4907 3010
rect 4757 2976 4802 3003
rect 4849 2976 4886 3003
rect 4941 2976 4942 3010
rect 4752 2969 4802 2976
rect 4836 2969 4886 2976
rect 4920 2969 4942 2976
rect 4718 2940 4942 2969
rect 4718 2928 4723 2940
rect 4757 2928 4815 2940
rect 4849 2928 4907 2940
rect 4757 2906 4802 2928
rect 4849 2906 4886 2928
rect 4941 2906 4942 2940
rect 4752 2894 4802 2906
rect 4836 2894 4886 2906
rect 4920 2894 4942 2906
rect 4718 2870 4942 2894
rect 4718 2853 4723 2870
rect 4757 2853 4815 2870
rect 4849 2853 4907 2870
rect 4757 2836 4802 2853
rect 4849 2836 4886 2853
rect 4941 2836 4942 2870
rect 4752 2819 4802 2836
rect 4836 2819 4886 2836
rect 4920 2819 4942 2836
rect 4718 2800 4942 2819
rect 4718 2778 4723 2800
rect 4757 2778 4815 2800
rect 4849 2778 4907 2800
rect 4757 2766 4802 2778
rect 4849 2766 4886 2778
rect 4941 2766 4942 2800
rect 4752 2744 4802 2766
rect 4836 2744 4886 2766
rect 4920 2744 4942 2766
rect 4718 2730 4942 2744
rect 4718 2703 4723 2730
rect 4757 2703 4815 2730
rect 4849 2703 4907 2730
rect 4757 2696 4802 2703
rect 4849 2696 4886 2703
rect 4941 2696 4942 2730
rect 4752 2669 4802 2696
rect 4836 2669 4886 2696
rect 4920 2669 4942 2696
rect 4718 2660 4942 2669
rect 4718 2628 4723 2660
rect 4757 2628 4815 2660
rect 4849 2628 4907 2660
rect 4757 2626 4802 2628
rect 4849 2626 4886 2628
rect 4941 2626 4942 2660
rect 4752 2594 4802 2626
rect 4836 2594 4886 2626
rect 4920 2594 4942 2626
rect 4718 2590 4942 2594
rect 4718 2556 4723 2590
rect 4757 2556 4815 2590
rect 4849 2556 4907 2590
rect 4941 2556 4942 2590
rect 4718 2553 4942 2556
rect 4752 2520 4802 2553
rect 4836 2520 4886 2553
rect 4920 2520 4942 2553
rect 4757 2519 4802 2520
rect 4849 2519 4886 2520
rect 4718 2486 4723 2519
rect 4757 2486 4815 2519
rect 4849 2486 4907 2519
rect 4941 2486 4942 2520
rect 4718 2478 4942 2486
rect 4752 2450 4802 2478
rect 4836 2450 4886 2478
rect 4920 2450 4942 2478
rect 4757 2444 4802 2450
rect 4849 2444 4886 2450
rect 4718 2416 4723 2444
rect 4757 2416 4815 2444
rect 4849 2416 4907 2444
rect 4941 2416 4942 2450
rect 4718 2403 4942 2416
rect 4752 2380 4802 2403
rect 4836 2380 4886 2403
rect 4920 2380 4942 2403
rect 4757 2369 4802 2380
rect 4849 2369 4886 2380
rect 4718 2346 4723 2369
rect 4757 2346 4815 2369
rect 4849 2346 4907 2369
rect 4941 2346 4942 2380
rect 4718 2328 4942 2346
rect 4752 2310 4802 2328
rect 4836 2310 4886 2328
rect 4920 2310 4942 2328
rect 4757 2294 4802 2310
rect 4849 2294 4886 2310
rect 4718 2276 4723 2294
rect 4757 2276 4815 2294
rect 4849 2276 4907 2294
rect 4941 2276 4942 2310
rect 4718 2254 4942 2276
rect 5097 3619 5173 3653
rect 5231 3619 5249 3653
rect 5299 3619 5325 3653
rect 5367 3619 5402 3653
rect 5436 3619 5479 3653
rect 5517 3619 5585 3653
rect 5097 3585 5131 3619
rect 5097 3517 5131 3547
rect 5551 3581 5585 3619
rect 5551 3513 5585 3547
rect 5097 3449 5131 3471
rect 5097 3381 5131 3395
rect 5097 3313 5131 3319
rect 5216 3470 5250 3486
rect 5216 3402 5250 3428
rect 5216 3334 5250 3356
rect 5432 3470 5466 3486
rect 5432 3402 5466 3428
rect 5432 3334 5466 3356
rect 5551 3445 5585 3475
rect 5551 3377 5585 3403
rect 5551 3309 5585 3331
rect 5097 3277 5131 3279
rect 5551 3241 5585 3259
rect 5097 3201 5131 3211
rect 5097 3125 5131 3143
rect 5326 3217 5360 3232
rect 5326 3216 5327 3217
rect 5360 3182 5361 3183
rect 5326 3148 5361 3182
rect 5360 3145 5361 3148
rect 5326 3111 5327 3114
rect 5551 3173 5585 3186
rect 5326 3098 5360 3111
rect 5551 3105 5585 3113
rect 5097 3049 5131 3075
rect 5097 2973 5131 3007
rect 5551 3037 5585 3040
rect 5551 3001 5585 3003
rect 5097 2905 5131 2939
rect 5097 2837 5131 2863
rect 5097 2769 5131 2787
rect 5216 2964 5250 2980
rect 5432 2964 5466 2980
rect 5216 2896 5250 2922
rect 5216 2828 5250 2850
rect 5291 2902 5329 2936
rect 5363 2902 5397 2936
rect 5291 2864 5397 2902
rect 5291 2830 5329 2864
rect 5363 2830 5397 2864
rect 5097 2701 5131 2711
rect 5097 2633 5131 2635
rect 5097 2593 5131 2599
rect 5291 2710 5397 2830
rect 5432 2896 5466 2922
rect 5432 2828 5466 2850
rect 5551 2928 5585 2935
rect 5551 2855 5585 2867
rect 5551 2782 5585 2799
rect 5291 2676 5326 2710
rect 5360 2676 5397 2710
rect 5291 2642 5397 2676
rect 5291 2608 5326 2642
rect 5360 2608 5397 2642
rect 5291 2574 5397 2608
rect 5551 2709 5585 2731
rect 5551 2629 5585 2663
rect 5097 2517 5131 2531
rect 5097 2441 5131 2463
rect 5097 2365 5131 2395
rect 5097 2289 5131 2327
rect 5551 2561 5585 2595
rect 5551 2493 5585 2527
rect 5551 2425 5585 2459
rect 5551 2357 5585 2391
rect 5551 2289 5585 2323
rect 5097 2255 5165 2289
rect 5203 2255 5233 2289
rect 5279 2255 5301 2289
rect 5354 2255 5369 2289
rect 5429 2255 5437 2289
rect 5504 2255 5545 2289
rect 5579 2255 5585 2289
rect 5738 3636 5772 3642
rect 5738 3594 5772 3602
rect 5738 3512 5772 3534
rect 5738 3432 5772 3466
rect 5738 3364 5772 3395
rect 5738 3296 5772 3308
rect 5863 3283 5878 3317
rect 5935 3283 5946 3317
rect 5980 3283 5996 3317
rect 6192 3283 6208 3317
rect 6242 3283 6276 3317
rect 6310 3283 6344 3317
rect 6378 3283 6470 3317
rect 6504 3283 6538 3317
rect 6572 3283 6580 3317
rect 6640 3283 6652 3317
rect 6764 3301 6766 3325
rect 5738 3228 5772 3231
rect 5738 3187 5772 3194
rect 6032 3242 6066 3248
rect 6730 3267 6732 3299
rect 6730 3253 6766 3267
rect 6032 3226 6142 3242
rect 6032 3210 6040 3226
rect 6074 3192 6108 3226
rect 6066 3176 6142 3192
rect 6764 3227 6766 3253
rect 6730 3193 6732 3219
rect 6730 3174 6766 3193
rect 6764 3153 6766 3174
rect 5738 3109 5772 3126
rect 5738 3031 5772 3058
rect 5738 2956 5772 2990
rect 5935 3107 6208 3141
rect 6242 3107 6260 3141
rect 6310 3107 6332 3141
rect 6378 3107 6470 3141
rect 6504 3107 6538 3141
rect 6572 3107 6606 3141
rect 6640 3107 6658 3141
rect 6730 3119 6732 3140
rect 5935 2970 5969 3107
rect 6730 3095 6766 3119
rect 6764 3079 6766 3095
rect 6040 3069 6142 3071
rect 6040 3055 6119 3069
rect 6074 3021 6108 3055
rect 6142 3021 6153 3035
rect 6040 3005 6153 3021
rect 5862 2965 5969 2970
rect 6119 2997 6153 3005
rect 5862 2931 5878 2965
rect 5912 2931 5946 2965
rect 5980 2931 5996 2965
rect 6730 3045 6732 3061
rect 6730 3016 6766 3045
rect 6764 3005 6766 3016
rect 6730 2971 6732 2982
rect 6192 2931 6208 2965
rect 6242 2931 6276 2965
rect 6310 2931 6344 2965
rect 6378 2931 6470 2965
rect 6504 2931 6538 2965
rect 6572 2931 6580 2965
rect 6640 2931 6652 2965
rect 6730 2937 6766 2971
rect 6764 2931 6766 2937
rect 5738 2888 5772 2919
rect 5738 2820 5772 2841
rect 6730 2897 6732 2903
rect 6730 2858 6766 2897
rect 5863 2806 5878 2840
rect 5935 2806 5946 2840
rect 5980 2806 5996 2840
rect 6192 2806 6208 2840
rect 6242 2806 6276 2840
rect 6310 2806 6344 2840
rect 6378 2806 6470 2840
rect 6504 2806 6538 2840
rect 6572 2806 6580 2840
rect 6640 2806 6652 2840
rect 6730 2785 6766 2824
rect 6730 2779 6732 2785
rect 5738 2752 5772 2763
rect 6040 2751 6316 2767
rect 6074 2717 6108 2751
rect 6142 2750 6316 2751
rect 6142 2717 6210 2750
rect 6040 2716 6210 2717
rect 6244 2716 6282 2750
rect 6040 2701 6316 2716
rect 6764 2745 6766 2751
rect 6730 2712 6766 2745
rect 5738 2684 5772 2685
rect 6730 2700 6732 2712
rect 6764 2666 6766 2678
rect 5738 2641 5772 2650
rect 5862 2630 5878 2664
rect 5912 2630 5946 2664
rect 5980 2630 6208 2664
rect 6242 2630 6259 2664
rect 6310 2630 6331 2664
rect 6378 2630 6470 2664
rect 6504 2630 6538 2664
rect 6572 2630 6606 2664
rect 6640 2630 6658 2664
rect 6730 2639 6766 2666
rect 6730 2621 6732 2639
rect 6764 2587 6766 2605
rect 5738 2548 5772 2582
rect 6732 2581 6766 2587
rect 4752 2240 4802 2254
rect 4836 2240 4886 2254
rect 4920 2240 4942 2254
rect 4757 2220 4802 2240
rect 4849 2220 4886 2240
rect 480 2169 514 2191
rect 480 2097 514 2123
rect 683 2181 1989 2197
rect 683 2147 1299 2181
rect 1333 2147 1413 2181
rect 1447 2155 1989 2181
rect 3938 2170 3972 2204
rect 1447 2147 2088 2155
rect 683 2120 2088 2147
rect 683 2086 778 2120
rect 812 2086 862 2120
rect 896 2086 946 2120
rect 980 2086 1030 2120
rect 1064 2086 1114 2120
rect 1148 2094 2088 2120
rect 1148 2086 1299 2094
rect 683 2060 1299 2086
rect 1333 2060 1413 2094
rect 1447 2060 2088 2094
rect 3938 2102 3972 2136
rect 4722 2206 4723 2220
rect 4757 2206 4815 2220
rect 4849 2206 4907 2220
rect 4941 2206 4942 2240
rect 4722 2170 4942 2206
rect 4722 2136 4723 2170
rect 4757 2136 4815 2170
rect 4849 2136 4907 2170
rect 4941 2136 4942 2170
rect 4722 2102 4942 2136
rect 5738 2102 5772 2514
rect 3530 2071 3564 2081
rect 3554 2065 3564 2071
rect 3938 2068 4038 2102
rect 4072 2068 4106 2102
rect 4140 2068 4174 2102
rect 4208 2068 4242 2102
rect 4276 2068 4310 2102
rect 4344 2068 4378 2102
rect 4412 2068 4446 2102
rect 4480 2068 4514 2102
rect 4548 2068 4582 2102
rect 4616 2068 4650 2102
rect 4684 2068 4718 2102
rect 4752 2068 4786 2102
rect 4820 2068 4854 2102
rect 4888 2068 4922 2102
rect 4956 2068 4990 2102
rect 5024 2068 5058 2102
rect 5092 2068 5126 2102
rect 5160 2068 5194 2102
rect 5228 2068 5262 2102
rect 5296 2068 5330 2102
rect 5364 2068 5398 2102
rect 5432 2068 5466 2102
rect 5500 2068 5534 2102
rect 5568 2068 5602 2102
rect 5636 2068 5670 2102
rect 5704 2068 5772 2102
rect 683 2059 2088 2060
rect 480 2039 514 2055
rect -823 1987 -763 2023
rect 171 1986 979 1989
rect -176 1982 -160 1983
rect -126 1982 -66 1983
rect -176 1949 -164 1982
rect -126 1949 -90 1982
rect -32 1949 -16 1983
rect 171 1952 184 1986
rect 221 1952 261 1986
rect 296 1952 337 1986
rect 372 1952 411 1986
rect 449 1952 485 1986
rect 526 1952 559 1986
rect 603 1952 633 1986
rect 679 1952 707 1986
rect 755 1952 781 1986
rect 831 1952 855 1986
rect 907 1952 929 1986
rect 963 1952 979 1986
rect 171 1949 979 1952
rect 1035 1949 1051 1983
rect 1104 1949 1125 1983
rect 1179 1949 1199 1983
rect 1254 1949 1273 1983
rect 1328 1949 1347 1983
rect 1402 1949 1421 1983
rect 1476 1949 1495 1983
rect 1550 1949 1569 1983
rect 1624 1949 1643 1983
rect 1698 1949 1718 1983
rect 1772 1949 1793 1983
rect 1827 1949 1843 1983
rect -130 1948 -90 1949
rect -221 1831 -187 1833
rect -221 1795 -187 1797
rect -221 1723 -187 1729
rect -676 1656 -638 1690
rect -530 1631 -496 1669
rect -221 1651 -187 1661
rect -221 1579 -187 1593
rect -221 1507 -187 1525
rect -221 1435 -187 1457
rect -823 1357 -763 1427
rect -221 1363 -187 1389
rect -221 1291 -187 1321
rect -221 1219 -187 1253
rect -221 1151 -187 1185
rect -221 1083 -187 1113
rect -221 1015 -187 1041
rect -221 947 -187 969
rect -5 1831 29 1833
rect -5 1795 29 1797
rect -5 1723 29 1729
rect -5 1651 29 1661
rect -5 1579 29 1593
rect -5 1507 29 1525
rect -5 1435 29 1457
rect -5 1363 29 1389
rect -5 1291 29 1321
rect -5 1219 29 1253
rect -5 1151 29 1185
rect -5 1083 29 1113
rect -5 1015 29 1041
rect -5 947 29 969
rect 126 1831 160 1833
rect 126 1795 160 1797
rect 126 1723 160 1729
rect 126 1651 160 1661
rect 126 1579 160 1593
rect 126 1507 160 1525
rect 126 1435 160 1457
rect 126 1363 160 1389
rect 126 1291 160 1321
rect 126 1219 160 1253
rect 126 1151 160 1185
rect 126 1083 160 1113
rect 126 1015 160 1041
rect 126 947 160 969
rect 342 1831 376 1833
rect 342 1795 376 1797
rect 342 1723 376 1729
rect 342 1651 376 1661
rect 342 1579 376 1593
rect 342 1507 376 1525
rect 342 1435 376 1457
rect 342 1363 376 1389
rect 342 1291 376 1321
rect 342 1219 376 1253
rect 342 1151 376 1185
rect 342 1083 376 1113
rect 342 1015 376 1041
rect 342 947 376 969
rect 558 1831 592 1833
rect 558 1795 592 1797
rect 558 1723 592 1729
rect 558 1651 592 1661
rect 558 1579 592 1593
rect 558 1507 592 1525
rect 558 1435 592 1457
rect 558 1363 592 1389
rect 558 1291 592 1321
rect 558 1219 592 1253
rect 558 1151 592 1185
rect 558 1083 592 1113
rect 558 1015 592 1041
rect 558 947 592 969
rect 774 1831 808 1833
rect 774 1795 808 1797
rect 774 1723 808 1729
rect 774 1651 808 1661
rect 774 1579 808 1593
rect 774 1507 808 1525
rect 774 1435 808 1457
rect 774 1363 808 1389
rect 774 1291 808 1321
rect 774 1219 808 1253
rect 774 1151 808 1185
rect 774 1083 808 1113
rect 774 1015 808 1041
rect 774 947 808 969
rect 990 1831 1024 1833
rect 990 1795 1024 1797
rect 990 1723 1024 1729
rect 990 1651 1024 1661
rect 990 1579 1024 1593
rect 990 1507 1024 1525
rect 990 1435 1024 1457
rect 990 1363 1024 1389
rect 990 1291 1024 1321
rect 990 1219 1024 1253
rect 990 1151 1024 1185
rect 990 1083 1024 1113
rect 990 1015 1024 1041
rect 990 947 1024 969
rect 1206 1831 1240 1833
rect 1206 1795 1240 1797
rect 1206 1723 1240 1729
rect 1206 1651 1240 1661
rect 1206 1579 1240 1593
rect 1206 1507 1240 1525
rect 1206 1435 1240 1457
rect 1206 1363 1240 1389
rect 1206 1291 1240 1321
rect 1206 1219 1240 1253
rect 1206 1151 1240 1185
rect 1206 1083 1240 1113
rect 1206 1015 1240 1041
rect 1206 947 1240 969
rect 1422 1831 1456 1833
rect 1422 1795 1456 1797
rect 1422 1723 1456 1729
rect 1422 1651 1456 1661
rect 1422 1579 1456 1593
rect 1422 1507 1456 1525
rect 1422 1435 1456 1457
rect 1422 1363 1456 1389
rect 1422 1291 1456 1321
rect 1422 1219 1456 1253
rect 1422 1151 1456 1185
rect 1422 1083 1456 1113
rect 1422 1015 1456 1041
rect 1422 947 1456 969
rect 1638 1831 1672 1833
rect 1638 1795 1672 1797
rect 1638 1723 1672 1729
rect 1638 1651 1672 1661
rect 1638 1579 1672 1593
rect 1638 1507 1672 1525
rect 1638 1435 1672 1457
rect 1638 1363 1672 1389
rect 1638 1291 1672 1321
rect 1638 1219 1672 1253
rect 1638 1151 1672 1185
rect 1638 1083 1672 1113
rect 1638 1015 1672 1041
rect 1638 947 1672 969
rect 1854 1831 1888 1833
rect 1854 1795 1888 1797
rect 1854 1723 1888 1729
rect 1854 1651 1888 1661
rect 1854 1579 1888 1593
rect 1854 1507 1888 1525
rect 1854 1435 1888 1457
rect 1854 1363 1888 1389
rect 1854 1291 1888 1321
rect 1854 1219 1888 1253
rect 1854 1151 1888 1185
rect 1854 1083 1888 1113
rect 1854 1015 1888 1041
rect 1854 947 1888 969
rect 1928 832 2088 2059
rect 2127 2053 2240 2065
rect 2161 2049 2240 2053
rect 2161 2019 2206 2049
rect 2127 2015 2206 2019
rect 2489 2049 2523 2065
rect 2127 1981 2240 2015
rect 2161 1947 2206 1981
rect 2127 1931 2240 1947
rect 2522 2007 2523 2015
rect 2488 1981 2523 2007
rect 3520 2031 3530 2037
rect 3520 1999 3564 2031
rect 3554 1997 3564 1999
rect 2488 1969 2489 1981
rect 2742 1983 2758 1989
rect 2792 1983 2853 1989
rect 2742 1955 2751 1983
rect 2792 1955 2850 1983
rect 2887 1955 2948 1989
rect 2982 1955 2998 1989
rect 3054 1955 3070 1989
rect 3104 1955 3165 1989
rect 3199 1983 3260 1989
rect 3294 1983 3310 1989
rect 3202 1955 3260 1983
rect 3301 1955 3310 1983
rect 2785 1949 2850 1955
rect 2884 1949 2948 1955
rect 3104 1949 3168 1955
rect 3202 1949 3267 1955
rect 3530 1947 3564 1963
rect 2522 1935 2523 1947
rect 2489 1931 2523 1935
rect 3934 1922 3950 1956
rect 3991 1933 4029 1967
rect 4063 1933 4064 1956
rect 3984 1922 4064 1933
rect 4098 1922 4114 1956
rect 2697 1837 2731 1839
rect 2131 1820 2165 1824
rect 2131 1748 2165 1774
rect 2131 1676 2165 1706
rect 2131 1604 2165 1638
rect 2131 1536 2165 1570
rect 2131 1468 2165 1498
rect 2131 1400 2165 1426
rect 2131 1332 2165 1354
rect 2287 1820 2321 1824
rect 2287 1748 2321 1774
rect 2287 1676 2321 1706
rect 2287 1604 2321 1638
rect 2287 1536 2321 1570
rect 2287 1468 2321 1498
rect 2287 1400 2321 1426
rect 2287 1332 2321 1354
rect 2414 1820 2448 1824
rect 2414 1748 2448 1774
rect 2414 1676 2448 1706
rect 2414 1604 2448 1638
rect 2414 1536 2448 1570
rect 2414 1468 2448 1498
rect 2414 1400 2448 1426
rect 2414 1332 2448 1354
rect 2570 1820 2604 1824
rect 2570 1748 2604 1774
rect 2570 1676 2604 1706
rect 2570 1604 2604 1638
rect 2570 1536 2604 1570
rect 2570 1468 2604 1498
rect 2570 1400 2604 1426
rect 2570 1332 2604 1354
rect 2697 1801 2731 1803
rect 2697 1729 2731 1735
rect 2697 1657 2731 1667
rect 2697 1585 2731 1599
rect 2697 1513 2731 1531
rect 2697 1441 2731 1463
rect 2697 1369 2731 1395
rect 2697 1297 2731 1327
rect 2697 1225 2731 1259
rect 2697 1157 2731 1191
rect 2697 1089 2731 1119
rect 2697 1021 2731 1047
rect 2697 953 2731 975
rect 2853 1837 2887 1839
rect 2853 1801 2887 1803
rect 2853 1729 2887 1735
rect 2853 1657 2887 1667
rect 2853 1585 2887 1599
rect 2853 1513 2887 1531
rect 2853 1441 2887 1463
rect 2853 1369 2887 1395
rect 2853 1297 2887 1327
rect 2853 1225 2887 1259
rect 2853 1157 2887 1191
rect 2853 1089 2887 1119
rect 2853 1021 2887 1047
rect 2853 953 2887 975
rect 3009 1837 3043 1839
rect 3009 1801 3043 1803
rect 3009 1729 3043 1735
rect 3009 1657 3043 1667
rect 3009 1585 3043 1599
rect 3009 1513 3043 1531
rect 3009 1441 3043 1463
rect 3009 1369 3043 1395
rect 3009 1297 3043 1327
rect 3009 1225 3043 1259
rect 3009 1157 3043 1191
rect 3009 1089 3043 1119
rect 3009 1021 3043 1047
rect 3009 953 3043 975
rect 3165 1837 3199 1839
rect 3165 1801 3199 1803
rect 3165 1729 3199 1735
rect 3165 1657 3199 1667
rect 3165 1585 3199 1599
rect 3165 1513 3199 1531
rect 3165 1441 3199 1463
rect 3165 1369 3199 1395
rect 3165 1297 3199 1327
rect 3165 1225 3199 1259
rect 3165 1157 3199 1191
rect 3165 1089 3199 1119
rect 3165 1021 3199 1047
rect 3165 953 3199 975
rect 3889 1841 3923 1857
rect 3321 1837 3355 1839
rect 3321 1801 3355 1803
rect 3321 1729 3355 1735
rect 3321 1657 3355 1667
rect 3321 1585 3355 1599
rect 3321 1513 3355 1531
rect 3321 1441 3355 1463
rect 3321 1369 3355 1395
rect 3321 1297 3355 1327
rect 3446 1835 3480 1839
rect 3446 1763 3480 1789
rect 3446 1691 3480 1721
rect 3446 1619 3480 1653
rect 3446 1551 3480 1585
rect 3446 1483 3480 1513
rect 3446 1415 3480 1441
rect 3446 1347 3480 1369
rect 3602 1835 3636 1839
rect 3602 1763 3636 1789
rect 3602 1691 3636 1721
rect 3889 1773 3923 1799
rect 3889 1705 3923 1727
rect 4125 1841 4159 1857
rect 4125 1773 4159 1799
rect 4125 1705 4159 1727
rect 3602 1619 3636 1653
rect 3602 1551 3636 1585
rect 3602 1483 3636 1513
rect 3602 1415 3636 1441
rect 3602 1347 3636 1369
rect 3321 1225 3355 1259
rect 3321 1157 3355 1191
rect 3321 1089 3355 1119
rect 3321 1021 3355 1047
rect 3321 953 3355 975
rect 3740 1048 3802 1082
rect 3836 1048 3898 1082
rect 3706 1006 3932 1048
rect 3740 972 3802 1006
rect 3836 972 3898 1006
rect 3706 930 3932 972
rect 3740 896 3802 930
rect 3836 896 3898 930
rect 3706 854 3932 896
rect 184 827 223 832
rect 257 827 296 832
rect 330 827 369 832
rect 403 827 441 832
rect 475 827 513 832
rect 547 827 585 832
rect 619 827 657 832
rect 691 827 729 832
rect 763 827 801 832
rect 835 827 873 832
rect 907 827 945 832
rect 979 827 1017 832
rect 1051 827 1089 832
rect 1123 827 1161 832
rect 1195 827 1233 832
rect 1267 827 1305 832
rect 1339 827 1377 832
rect 1411 827 1449 832
rect 1483 827 1521 832
rect 1555 827 1593 832
rect 1627 827 1665 832
rect 1699 827 1737 832
rect 1771 827 1809 832
rect 1843 827 1881 832
rect 1915 827 1953 832
rect 1987 827 2025 832
rect 2059 827 2097 832
rect 2131 827 2169 832
rect 2203 827 2241 832
rect 2275 827 2313 832
rect 2347 827 2385 832
rect 2419 827 2457 832
rect 2491 827 2529 832
rect 2563 827 2601 832
rect 2635 827 2673 832
rect 2707 827 2745 832
rect 2779 827 2817 832
rect 2851 827 2889 832
rect 2923 827 2961 832
rect 2995 827 3033 832
rect 3067 827 3105 832
rect 3139 827 3177 832
rect 3211 827 3249 832
rect 3283 827 3321 832
rect 144 798 150 827
rect 202 798 223 827
rect 271 798 296 827
rect 340 798 369 827
rect 409 798 441 827
rect 144 793 168 798
rect 202 793 237 798
rect 271 793 306 798
rect 340 793 375 798
rect 409 793 444 798
rect 478 793 513 827
rect 547 793 582 827
rect 619 798 651 827
rect 691 798 720 827
rect 763 798 789 827
rect 835 798 858 827
rect 907 798 927 827
rect 979 798 996 827
rect 1051 798 1065 827
rect 1123 798 1134 827
rect 1195 798 1203 827
rect 1267 798 1272 827
rect 1339 798 1341 827
rect 616 793 651 798
rect 685 793 720 798
rect 754 793 789 798
rect 823 793 858 798
rect 892 793 927 798
rect 961 793 996 798
rect 1030 793 1065 798
rect 1099 793 1134 798
rect 1168 793 1203 798
rect 1237 793 1272 798
rect 1306 793 1341 798
rect 1375 798 1377 827
rect 1444 798 1449 827
rect 1513 798 1521 827
rect 1582 798 1593 827
rect 1651 798 1665 827
rect 1720 798 1737 827
rect 1789 798 1809 827
rect 1858 798 1881 827
rect 1927 798 1953 827
rect 1996 798 2025 827
rect 2065 798 2097 827
rect 1375 793 1410 798
rect 1444 793 1479 798
rect 1513 793 1548 798
rect 1582 793 1617 798
rect 1651 793 1686 798
rect 1720 793 1755 798
rect 1789 793 1824 798
rect 1858 793 1893 798
rect 1927 793 1962 798
rect 1996 793 2031 798
rect 2065 793 2100 798
rect 2134 793 2169 827
rect 2203 793 2238 827
rect 2275 798 2307 827
rect 2347 798 2376 827
rect 2419 798 2445 827
rect 2491 798 2514 827
rect 2563 798 2583 827
rect 2635 798 2652 827
rect 2707 798 2721 827
rect 2779 798 2790 827
rect 2851 798 2859 827
rect 2923 798 2928 827
rect 2995 798 2996 827
rect 2272 793 2307 798
rect 2341 793 2376 798
rect 2410 793 2445 798
rect 2479 793 2514 798
rect 2548 793 2583 798
rect 2617 793 2652 798
rect 2686 793 2721 798
rect 2755 793 2790 798
rect 2824 793 2859 798
rect 2893 793 2928 798
rect 2962 793 2996 798
rect 3030 798 3033 827
rect 3098 798 3105 827
rect 3166 798 3177 827
rect 3234 798 3249 827
rect 3302 798 3321 827
rect 3030 793 3064 798
rect 3098 793 3132 798
rect 3166 793 3200 798
rect 3234 793 3268 798
rect 3302 793 3336 798
rect 3370 793 3394 827
rect 3740 820 3802 854
rect 3836 820 3898 854
rect 3706 778 3932 820
rect 3740 744 3802 778
rect 3836 744 3898 778
rect 3317 704 3318 738
rect 3352 704 3400 738
rect 3434 704 3482 738
rect 3516 704 3517 738
rect 227 640 241 674
rect 295 640 313 674
rect 363 640 385 674
rect 431 640 457 674
rect 499 640 529 674
rect 567 640 601 674
rect 635 640 669 674
rect 707 640 737 674
rect 779 640 805 674
rect 851 640 873 674
rect 923 640 941 674
rect 995 640 1009 674
rect 1067 640 1077 674
rect 1139 640 1145 674
rect 1211 640 1213 674
rect 1247 640 1249 674
rect 1315 640 1321 674
rect 1383 640 1393 674
rect 1451 640 1465 674
rect 1519 640 1537 674
rect 1587 640 1609 674
rect 1655 640 1681 674
rect 1723 640 1753 674
rect 1791 640 1825 674
rect 1859 640 1893 674
rect 1931 640 1961 674
rect 2003 640 2029 674
rect 2075 640 2097 674
rect 2191 612 2225 628
rect 2191 540 2226 578
rect 2191 506 2192 540
rect 2697 611 2731 633
rect 2697 539 2731 565
rect 2191 498 2225 506
rect 2697 481 2731 497
rect 2853 611 2887 633
rect 2853 539 2887 565
rect 2853 481 2887 497
rect 3009 611 3043 633
rect 3009 539 3043 565
rect 3009 481 3043 497
rect 3165 611 3199 633
rect 3165 539 3199 565
rect 3317 635 3517 704
rect 3317 601 3318 635
rect 3352 601 3400 635
rect 3434 601 3482 635
rect 3516 601 3517 635
rect 3317 533 3517 601
rect 3317 499 3318 533
rect 3352 499 3400 533
rect 3434 499 3482 533
rect 3516 499 3517 533
rect 3165 481 3199 497
rect 2191 448 2225 464
rect 227 404 241 438
rect 295 404 313 438
rect 363 404 385 438
rect 431 404 457 438
rect 499 404 529 438
rect 567 404 601 438
rect 635 404 669 438
rect 707 404 737 438
rect 779 404 805 438
rect 851 404 873 438
rect 923 404 941 438
rect 995 404 1009 438
rect 1067 404 1077 438
rect 1139 404 1145 438
rect 1211 404 1213 438
rect 1247 404 1249 438
rect 1315 404 1321 438
rect 1383 404 1393 438
rect 1451 404 1465 438
rect 1519 404 1537 438
rect 1587 404 1609 438
rect 1655 404 1681 438
rect 1723 404 1753 438
rect 1791 404 1825 438
rect 1859 404 1893 438
rect 1931 404 1961 438
rect 2003 404 2029 438
rect 2075 404 2097 438
rect 2742 397 2758 431
rect 2799 397 2828 431
rect 2881 397 2897 431
rect 2963 397 2966 431
rect 3000 397 3010 431
rect 3069 397 3091 431
rect 3138 397 3154 431
rect 227 277 241 311
rect 295 277 313 311
rect 363 277 385 311
rect 431 277 457 311
rect 499 277 529 311
rect 567 277 601 311
rect 635 277 669 311
rect 707 277 737 311
rect 779 277 805 311
rect 851 277 873 311
rect 923 277 941 311
rect 995 277 1009 311
rect 1067 277 1077 311
rect 1139 277 1145 311
rect 1211 277 1213 311
rect 1247 277 1249 311
rect 1315 277 1321 311
rect 1383 277 1393 311
rect 1451 277 1465 311
rect 1519 277 1537 311
rect 1587 277 1609 311
rect 1655 277 1681 311
rect 1723 277 1753 311
rect 1791 277 1825 311
rect 1859 277 1893 311
rect 1931 277 1961 311
rect 2003 277 2029 311
rect 2075 277 2097 311
rect 2191 250 2225 266
rect 2191 208 2225 216
rect 2191 174 2192 208
rect 2191 136 2226 174
rect 2191 86 2225 102
rect 227 41 241 75
rect 295 41 313 75
rect 363 41 385 75
rect 431 41 457 75
rect 499 41 529 75
rect 567 41 601 75
rect 635 41 669 75
rect 707 41 737 75
rect 779 41 805 75
rect 851 41 873 75
rect 923 41 941 75
rect 995 41 1009 75
rect 1067 41 1077 75
rect 1139 41 1145 75
rect 1211 41 1213 75
rect 1247 41 1249 75
rect 1315 41 1321 75
rect 1383 41 1393 75
rect 1451 41 1465 75
rect 1519 41 1537 75
rect 1587 41 1609 75
rect 1655 41 1681 75
rect 1723 41 1753 75
rect 1791 41 1825 75
rect 1859 41 1893 75
rect 1931 41 1961 75
rect 2003 41 2029 75
rect 2075 41 2097 75
rect -11566 -8658 -11500 -8643
rect -11566 -8659 -11540 -8658
rect -11566 -8693 -11550 -8659
rect -11506 -8692 -11500 -8658
rect -11516 -8693 -11500 -8692
rect -11566 -8727 -11500 -8693
rect -11566 -8761 -11550 -8727
rect -11516 -8730 -11500 -8727
rect -11566 -8764 -11540 -8761
rect -11506 -8764 -11500 -8730
rect -11566 -8777 -11500 -8764
rect -29100 -8875 -29046 -8847
rect -29012 -8875 -28958 -8847
rect -28924 -8875 -28870 -8847
rect -28836 -8870 -28189 -8847
rect -28155 -8870 -28115 -8847
rect -28081 -8870 -28041 -8847
rect -28007 -8870 -27967 -8847
rect -27933 -8870 -27893 -8847
rect -27859 -8870 -27819 -8847
rect -27785 -8870 -27745 -8847
rect -27711 -8870 -27671 -8847
rect -27637 -8870 -27597 -8847
rect -27563 -8870 -27523 -8847
rect -27489 -8870 -27449 -8847
rect -27415 -8870 -27375 -8847
rect -27341 -8870 -27301 -8847
rect -27267 -8870 -27227 -8847
rect -27193 -8870 -27153 -8847
rect -27119 -8870 -27036 -8847
rect -28836 -8875 -27036 -8870
rect -31669 -8884 -27036 -8875
rect -31669 -8918 -31632 -8884
rect -27450 -8908 -27415 -8884
rect -32352 -9600 -32338 -8918
rect -27450 -8942 -27449 -8908
rect -27381 -8908 -27346 -8884
rect -27312 -8908 -27277 -8884
rect -27243 -8908 -27208 -8884
rect -27174 -8908 -27139 -8884
rect -27381 -8918 -27375 -8908
rect -27312 -8918 -27301 -8908
rect -27243 -8918 -27227 -8908
rect -27174 -8918 -27153 -8908
rect -27105 -8918 -27070 -8884
rect -27415 -8942 -27375 -8918
rect -27341 -8942 -27301 -8918
rect -27267 -8942 -27227 -8918
rect -27193 -8942 -27153 -8918
rect -27119 -8942 -27036 -8918
rect -27450 -8952 -27036 -8942
rect -27450 -8980 -27415 -8952
rect -27450 -9014 -27449 -8980
rect -27381 -8980 -27346 -8952
rect -27312 -8980 -27277 -8952
rect -27243 -8980 -27208 -8952
rect -27174 -8980 -27139 -8952
rect -27381 -8986 -27375 -8980
rect -27312 -8986 -27301 -8980
rect -27243 -8986 -27227 -8980
rect -27174 -8986 -27153 -8980
rect -27105 -8986 -27070 -8952
rect -27415 -9014 -27375 -8986
rect -27341 -9014 -27301 -8986
rect -27267 -9014 -27227 -8986
rect -27193 -9014 -27153 -8986
rect -27119 -9014 -27036 -8986
rect -27450 -9020 -27036 -9014
rect -27450 -9052 -27415 -9020
rect -27450 -9086 -27449 -9052
rect -27381 -9052 -27346 -9020
rect -27312 -9052 -27277 -9020
rect -27243 -9052 -27208 -9020
rect -27174 -9052 -27139 -9020
rect -27381 -9054 -27375 -9052
rect -27312 -9054 -27301 -9052
rect -27243 -9054 -27227 -9052
rect -27174 -9054 -27153 -9052
rect -27105 -9054 -27070 -9020
rect -27415 -9086 -27375 -9054
rect -27341 -9086 -27301 -9054
rect -27267 -9086 -27227 -9054
rect -27193 -9086 -27153 -9054
rect -27119 -9086 -27036 -9054
rect -27450 -9088 -27036 -9086
rect -27450 -9122 -27415 -9088
rect -27381 -9122 -27346 -9088
rect -27312 -9122 -27277 -9088
rect -27243 -9122 -27208 -9088
rect -27174 -9122 -27139 -9088
rect -27105 -9122 -27070 -9088
rect -27450 -9124 -27036 -9122
rect -27450 -9158 -27449 -9124
rect -27415 -9156 -27375 -9124
rect -27341 -9156 -27301 -9124
rect -27267 -9156 -27227 -9124
rect -27193 -9156 -27153 -9124
rect -27119 -9156 -27036 -9124
rect -27450 -9190 -27415 -9158
rect -27381 -9158 -27375 -9156
rect -27312 -9158 -27301 -9156
rect -27243 -9158 -27227 -9156
rect -27174 -9158 -27153 -9156
rect -27381 -9190 -27346 -9158
rect -27312 -9190 -27277 -9158
rect -27243 -9190 -27208 -9158
rect -27174 -9190 -27139 -9158
rect -27105 -9190 -27070 -9156
rect -27450 -9196 -27036 -9190
rect -27450 -9230 -27449 -9196
rect -27415 -9224 -27375 -9196
rect -27341 -9224 -27301 -9196
rect -27267 -9224 -27227 -9196
rect -27193 -9224 -27153 -9196
rect -27119 -9224 -27036 -9196
rect -27450 -9258 -27415 -9230
rect -27381 -9230 -27375 -9224
rect -27312 -9230 -27301 -9224
rect -27243 -9230 -27227 -9224
rect -27174 -9230 -27153 -9224
rect -27381 -9258 -27346 -9230
rect -27312 -9258 -27277 -9230
rect -27243 -9258 -27208 -9230
rect -27174 -9258 -27139 -9230
rect -27105 -9258 -27070 -9224
rect -27450 -9268 -27036 -9258
rect -27450 -9302 -27449 -9268
rect -27415 -9292 -27375 -9268
rect -27341 -9292 -27301 -9268
rect -27267 -9292 -27227 -9268
rect -27193 -9292 -27153 -9268
rect -27119 -9292 -27036 -9268
rect -27450 -9326 -27415 -9302
rect -27381 -9302 -27375 -9292
rect -27312 -9302 -27301 -9292
rect -27243 -9302 -27227 -9292
rect -27174 -9302 -27153 -9292
rect -27381 -9326 -27346 -9302
rect -27312 -9326 -27277 -9302
rect -27243 -9326 -27208 -9302
rect -27174 -9326 -27139 -9302
rect -27105 -9326 -27070 -9292
rect -27450 -9340 -27036 -9326
rect -27450 -9374 -27449 -9340
rect -27415 -9360 -27375 -9340
rect -27341 -9360 -27301 -9340
rect -27267 -9360 -27227 -9340
rect -27193 -9360 -27153 -9340
rect -27119 -9360 -27036 -9340
rect -27450 -9394 -27415 -9374
rect -27381 -9374 -27375 -9360
rect -27312 -9374 -27301 -9360
rect -27243 -9374 -27227 -9360
rect -27174 -9374 -27153 -9360
rect -27381 -9394 -27346 -9374
rect -27312 -9394 -27277 -9374
rect -27243 -9394 -27208 -9374
rect -27174 -9394 -27139 -9374
rect -27105 -9394 -27070 -9360
rect -27450 -9428 -27036 -9394
rect -27450 -9462 -27415 -9428
rect -27381 -9462 -27346 -9428
rect -27312 -9462 -27277 -9428
rect -27243 -9462 -27208 -9428
rect -27174 -9462 -27139 -9428
rect -27105 -9462 -27070 -9428
rect -27450 -9496 -27036 -9462
rect -27450 -9530 -27415 -9496
rect -27381 -9530 -27346 -9496
rect -27312 -9530 -27277 -9496
rect -27243 -9530 -27208 -9496
rect -27174 -9530 -27139 -9496
rect -27105 -9530 -27070 -9496
rect -27450 -9564 -27036 -9530
rect -27450 -9598 -27415 -9564
rect -27381 -9598 -27346 -9564
rect -27312 -9598 -27277 -9564
rect -27243 -9598 -27208 -9564
rect -27174 -9598 -27139 -9564
rect -27105 -9598 -27070 -9564
rect -30792 -9600 -30753 -9598
rect -30719 -9600 -30680 -9598
rect -30646 -9600 -30607 -9598
rect -30573 -9600 -30534 -9598
rect -30500 -9600 -30461 -9598
rect -30427 -9600 -30388 -9598
rect -30354 -9600 -30315 -9598
rect -30281 -9600 -30242 -9598
rect -30208 -9600 -30169 -9598
rect -30135 -9600 -30096 -9598
rect -30062 -9600 -30023 -9598
rect -29989 -9600 -29950 -9598
rect -29916 -9600 -29877 -9598
rect -29843 -9600 -29804 -9598
rect -29770 -9600 -29731 -9598
rect -29697 -9600 -29658 -9598
rect -29624 -9600 -29585 -9598
rect -29551 -9600 -29512 -9598
rect -29478 -9600 -29439 -9598
rect -29405 -9600 -29366 -9598
rect -29332 -9600 -29293 -9598
rect -29259 -9600 -29220 -9598
rect -29186 -9600 -27036 -9598
rect -32352 -9635 -32315 -9600
rect -31669 -9635 -27036 -9600
<< viali >>
rect -32344 4310 -32315 4332
rect -32315 4310 -32310 4332
rect -32266 4310 -32247 4332
rect -32247 4310 -32232 4332
rect -32188 4310 -32179 4332
rect -32179 4310 -32154 4332
rect -32110 4310 -32077 4332
rect -32077 4310 -32076 4332
rect -32032 4310 -32009 4332
rect -32009 4310 -31998 4332
rect -31954 4310 -31941 4332
rect -31941 4310 -31920 4332
rect -31876 4310 -31873 4332
rect -31873 4310 -31842 4332
rect -31798 4310 -31771 4332
rect -31771 4310 -31764 4332
rect -31718 4310 -31703 4333
rect -31703 4310 -31684 4333
rect -32344 4298 -32310 4310
rect -32266 4298 -32232 4310
rect -32188 4298 -32154 4310
rect -32110 4298 -32076 4310
rect -32032 4298 -31998 4310
rect -31954 4298 -31920 4310
rect -31876 4298 -31842 4310
rect -31798 4298 -31764 4310
rect -31718 4299 -31684 4310
rect -31645 4299 -31611 4333
rect -31572 4299 -31538 4333
rect -31499 4299 -31465 4333
rect -31426 4299 -31392 4333
rect -31353 4299 -31319 4333
rect -31280 4299 -31246 4333
rect -31207 4299 -31173 4333
rect -31134 4299 -31100 4333
rect -31061 4299 -31027 4333
rect -30988 4299 -30954 4333
rect -30915 4299 -30881 4333
rect -30842 4299 -30808 4333
rect -30768 4299 -30734 4333
rect -30694 4299 -30660 4333
rect -30620 4299 -30586 4333
rect -30546 4299 -30512 4333
rect -30472 4299 -30438 4333
rect -30398 4299 -30364 4333
rect -30324 4299 -30290 4333
rect -30250 4299 -30216 4333
rect -30176 4299 -30142 4333
rect -30102 4299 -30068 4333
rect -30028 4299 -29994 4333
rect -29954 4299 -29920 4333
rect -29880 4299 -29846 4333
rect -29806 4299 -29772 4333
rect -29732 4299 -29698 4333
rect -29658 4299 -29624 4333
rect -29584 4299 -29550 4333
rect -29510 4299 -29476 4333
rect -29436 4299 -29402 4333
rect -29362 4299 -29328 4333
rect -29288 4299 -29254 4333
rect -29214 4299 -29180 4333
rect -29134 4299 -29100 4333
rect -29046 4310 -29044 4333
rect -29044 4310 -29012 4333
rect -28958 4310 -28942 4333
rect -28942 4310 -28924 4333
rect -28870 4310 -28840 4333
rect -28840 4310 -28836 4333
rect -29046 4299 -29012 4310
rect -28958 4299 -28924 4310
rect -28870 4299 -28836 4310
rect -32344 4241 -32315 4259
rect -32315 4241 -32310 4259
rect -32266 4241 -32247 4259
rect -32247 4241 -32232 4259
rect -32188 4241 -32179 4259
rect -32179 4241 -32154 4259
rect -32110 4241 -32077 4259
rect -32077 4241 -32076 4259
rect -32032 4241 -32009 4259
rect -32009 4241 -31998 4259
rect -31954 4241 -31941 4259
rect -31941 4241 -31920 4259
rect -31876 4241 -31873 4259
rect -31873 4241 -31842 4259
rect -31798 4241 -31771 4259
rect -31771 4241 -31764 4259
rect -31718 4241 -31703 4261
rect -31703 4241 -31684 4261
rect -31645 4242 -31632 4261
rect -31632 4242 -31611 4261
rect -31572 4242 -31563 4261
rect -31563 4242 -31538 4261
rect -31499 4242 -31494 4261
rect -31494 4242 -31465 4261
rect -31426 4242 -31425 4261
rect -31425 4242 -31392 4261
rect -31353 4242 -31322 4261
rect -31322 4242 -31319 4261
rect -31280 4242 -31253 4261
rect -31253 4242 -31246 4261
rect -31207 4242 -31184 4261
rect -31184 4242 -31173 4261
rect -31134 4242 -31115 4261
rect -31115 4242 -31100 4261
rect -31061 4242 -31046 4261
rect -31046 4242 -31027 4261
rect -30988 4242 -30977 4261
rect -30977 4242 -30954 4261
rect -30915 4242 -30908 4261
rect -30908 4242 -30881 4261
rect -30842 4242 -30839 4261
rect -30839 4242 -30808 4261
rect -30768 4242 -30735 4261
rect -30735 4242 -30734 4261
rect -30694 4242 -30666 4261
rect -30666 4242 -30660 4261
rect -30620 4242 -30597 4261
rect -30597 4242 -30586 4261
rect -30546 4242 -30528 4261
rect -30528 4242 -30512 4261
rect -30472 4242 -30459 4261
rect -30459 4242 -30438 4261
rect -30398 4242 -30390 4261
rect -30390 4242 -30364 4261
rect -30324 4242 -30321 4261
rect -30321 4242 -30290 4261
rect -30250 4242 -30218 4261
rect -30218 4242 -30216 4261
rect -30176 4242 -30149 4261
rect -30149 4242 -30142 4261
rect -30102 4242 -30080 4261
rect -30080 4242 -30068 4261
rect -30028 4242 -30011 4261
rect -30011 4242 -29994 4261
rect -29954 4242 -29942 4261
rect -29942 4242 -29920 4261
rect -29880 4242 -29873 4261
rect -29873 4242 -29846 4261
rect -29806 4242 -29804 4261
rect -29804 4242 -29772 4261
rect -29732 4242 -29700 4261
rect -29700 4242 -29698 4261
rect -29658 4242 -29631 4261
rect -29631 4242 -29624 4261
rect -29584 4242 -29562 4261
rect -29562 4242 -29550 4261
rect -29510 4242 -29493 4261
rect -29493 4242 -29476 4261
rect -29436 4242 -29424 4261
rect -29424 4242 -29402 4261
rect -29362 4242 -29355 4261
rect -29355 4242 -29328 4261
rect -29288 4242 -29286 4261
rect -29286 4242 -29254 4261
rect -29214 4242 -29183 4261
rect -29183 4242 -29180 4261
rect -29134 4242 -29114 4260
rect -29114 4242 -29100 4260
rect -32344 4225 -32310 4241
rect -32266 4225 -32232 4241
rect -32188 4225 -32154 4241
rect -32110 4225 -32076 4241
rect -32032 4225 -31998 4241
rect -31954 4225 -31920 4241
rect -31876 4225 -31842 4241
rect -31798 4225 -31764 4241
rect -31718 4227 -31684 4241
rect -31645 4227 -31611 4242
rect -31572 4227 -31538 4242
rect -31499 4227 -31465 4242
rect -31426 4227 -31392 4242
rect -31353 4227 -31319 4242
rect -31280 4227 -31246 4242
rect -31207 4227 -31173 4242
rect -31134 4227 -31100 4242
rect -31061 4227 -31027 4242
rect -30988 4227 -30954 4242
rect -30915 4227 -30881 4242
rect -30842 4227 -30808 4242
rect -30768 4227 -30734 4242
rect -30694 4227 -30660 4242
rect -30620 4227 -30586 4242
rect -30546 4227 -30512 4242
rect -30472 4227 -30438 4242
rect -30398 4227 -30364 4242
rect -30324 4227 -30290 4242
rect -30250 4227 -30216 4242
rect -30176 4227 -30142 4242
rect -30102 4227 -30068 4242
rect -30028 4227 -29994 4242
rect -29954 4227 -29920 4242
rect -29880 4227 -29846 4242
rect -29806 4227 -29772 4242
rect -29732 4227 -29698 4242
rect -29658 4227 -29624 4242
rect -29584 4227 -29550 4242
rect -29510 4227 -29476 4242
rect -29436 4227 -29402 4242
rect -29362 4227 -29328 4242
rect -29288 4227 -29254 4242
rect -29214 4227 -29180 4242
rect -29134 4226 -29100 4242
rect -29046 4241 -29044 4260
rect -29044 4241 -29012 4260
rect -28958 4241 -28942 4260
rect -28942 4241 -28924 4260
rect -28870 4241 -28840 4260
rect -28840 4241 -28836 4260
rect -29046 4226 -29012 4241
rect -28958 4226 -28924 4241
rect -28870 4226 -28836 4241
rect -28189 4206 -28155 4239
rect -28115 4206 -28081 4239
rect -28041 4206 -28007 4239
rect -27967 4206 -27933 4239
rect -27893 4206 -27859 4239
rect -27819 4206 -27785 4239
rect -27745 4206 -27711 4239
rect -27671 4206 -27637 4239
rect -27597 4206 -27563 4239
rect -27523 4206 -27489 4239
rect -27449 4206 -27415 4239
rect -27375 4206 -27341 4239
rect -27301 4206 -27267 4239
rect -27227 4206 -27193 4239
rect -27153 4206 -27119 4239
rect -32344 4172 -32315 4186
rect -32315 4172 -32310 4186
rect -32266 4172 -32247 4186
rect -32247 4172 -32232 4186
rect -32188 4172 -32179 4186
rect -32179 4172 -32154 4186
rect -32110 4172 -32077 4186
rect -32077 4172 -32076 4186
rect -32032 4172 -32009 4186
rect -32009 4172 -31998 4186
rect -31954 4172 -31941 4186
rect -31941 4172 -31920 4186
rect -31876 4172 -31873 4186
rect -31873 4172 -31842 4186
rect -31798 4172 -31771 4186
rect -31771 4172 -31764 4186
rect -31718 4172 -31703 4189
rect -31703 4172 -31684 4189
rect -31645 4172 -31632 4189
rect -31632 4172 -31611 4189
rect -31572 4172 -31563 4189
rect -31563 4172 -31538 4189
rect -31499 4172 -31494 4189
rect -31494 4172 -31465 4189
rect -31426 4172 -31425 4189
rect -31425 4172 -31392 4189
rect -31353 4172 -31322 4189
rect -31322 4172 -31319 4189
rect -31280 4172 -31253 4189
rect -31253 4172 -31246 4189
rect -31207 4172 -31184 4189
rect -31184 4172 -31173 4189
rect -31134 4172 -31115 4189
rect -31115 4172 -31100 4189
rect -31061 4172 -31046 4189
rect -31046 4172 -31027 4189
rect -30988 4172 -30977 4189
rect -30977 4172 -30954 4189
rect -30915 4172 -30908 4189
rect -30908 4172 -30881 4189
rect -30842 4172 -30839 4189
rect -30839 4172 -30808 4189
rect -30768 4172 -30735 4189
rect -30735 4172 -30734 4189
rect -30694 4172 -30666 4189
rect -30666 4172 -30660 4189
rect -30620 4172 -30597 4189
rect -30597 4172 -30586 4189
rect -30546 4172 -30528 4189
rect -30528 4172 -30512 4189
rect -30472 4172 -30459 4189
rect -30459 4172 -30438 4189
rect -30398 4172 -30390 4189
rect -30390 4172 -30364 4189
rect -30324 4172 -30321 4189
rect -30321 4172 -30290 4189
rect -30250 4172 -30218 4189
rect -30218 4172 -30216 4189
rect -30176 4172 -30149 4189
rect -30149 4172 -30142 4189
rect -30102 4172 -30080 4189
rect -30080 4172 -30068 4189
rect -30028 4172 -30011 4189
rect -30011 4172 -29994 4189
rect -29954 4172 -29942 4189
rect -29942 4172 -29920 4189
rect -29880 4172 -29873 4189
rect -29873 4172 -29846 4189
rect -29806 4172 -29804 4189
rect -29804 4172 -29772 4189
rect -29732 4172 -29700 4189
rect -29700 4172 -29698 4189
rect -29658 4172 -29631 4189
rect -29631 4172 -29624 4189
rect -29584 4172 -29562 4189
rect -29562 4172 -29550 4189
rect -29510 4172 -29493 4189
rect -29493 4172 -29476 4189
rect -29436 4172 -29424 4189
rect -29424 4172 -29402 4189
rect -29362 4172 -29355 4189
rect -29355 4172 -29328 4189
rect -29288 4172 -29286 4189
rect -29286 4172 -29254 4189
rect -29214 4172 -29183 4189
rect -29183 4172 -29180 4189
rect -29134 4172 -29114 4187
rect -29114 4172 -29100 4187
rect -29046 4172 -29044 4187
rect -29044 4172 -29012 4187
rect -28958 4172 -28942 4187
rect -28942 4172 -28924 4187
rect -28870 4172 -28840 4187
rect -28840 4172 -28836 4187
rect -28189 4205 -28160 4206
rect -28160 4205 -28155 4206
rect -28115 4205 -28092 4206
rect -28092 4205 -28081 4206
rect -28041 4205 -28024 4206
rect -28024 4205 -28007 4206
rect -27967 4205 -27956 4206
rect -27956 4205 -27933 4206
rect -27893 4205 -27888 4206
rect -27888 4205 -27859 4206
rect -27819 4205 -27786 4206
rect -27786 4205 -27785 4206
rect -27745 4205 -27718 4206
rect -27718 4205 -27711 4206
rect -27671 4205 -27650 4206
rect -27650 4205 -27637 4206
rect -27597 4205 -27582 4206
rect -27582 4205 -27563 4206
rect -27523 4205 -27514 4206
rect -27514 4205 -27489 4206
rect -27449 4205 -27446 4206
rect -27446 4205 -27415 4206
rect -27375 4205 -27344 4206
rect -27344 4205 -27341 4206
rect -27301 4205 -27276 4206
rect -27276 4205 -27267 4206
rect -27227 4205 -27208 4206
rect -27208 4205 -27193 4206
rect -27153 4205 -27140 4206
rect -27140 4205 -27119 4206
rect -9790 4278 -9756 4312
rect -9790 4210 -9756 4240
rect -9790 4206 -9756 4210
rect -32344 4152 -32310 4172
rect -32266 4152 -32232 4172
rect -32188 4152 -32154 4172
rect -32110 4152 -32076 4172
rect -32032 4152 -31998 4172
rect -31954 4152 -31920 4172
rect -31876 4152 -31842 4172
rect -31798 4152 -31764 4172
rect -31718 4155 -31684 4172
rect -31645 4155 -31611 4172
rect -31572 4155 -31538 4172
rect -31499 4155 -31465 4172
rect -31426 4155 -31392 4172
rect -31353 4155 -31319 4172
rect -31280 4155 -31246 4172
rect -31207 4155 -31173 4172
rect -31134 4155 -31100 4172
rect -31061 4155 -31027 4172
rect -30988 4155 -30954 4172
rect -30915 4155 -30881 4172
rect -30842 4155 -30808 4172
rect -30768 4155 -30734 4172
rect -30694 4155 -30660 4172
rect -30620 4155 -30586 4172
rect -30546 4155 -30512 4172
rect -30472 4155 -30438 4172
rect -30398 4155 -30364 4172
rect -30324 4155 -30290 4172
rect -30250 4155 -30216 4172
rect -30176 4155 -30142 4172
rect -30102 4155 -30068 4172
rect -30028 4155 -29994 4172
rect -29954 4155 -29920 4172
rect -29880 4155 -29846 4172
rect -29806 4155 -29772 4172
rect -29732 4155 -29698 4172
rect -29658 4155 -29624 4172
rect -29584 4155 -29550 4172
rect -29510 4155 -29476 4172
rect -29436 4155 -29402 4172
rect -29362 4155 -29328 4172
rect -29288 4155 -29254 4172
rect -29214 4155 -29180 4172
rect -29134 4153 -29100 4172
rect -29046 4153 -29012 4172
rect -28958 4153 -28924 4172
rect -28870 4153 -28836 4172
rect -28189 4137 -28155 4166
rect -28115 4137 -28081 4166
rect -28041 4137 -28007 4166
rect -27967 4137 -27933 4166
rect -27893 4137 -27859 4166
rect -27819 4137 -27785 4166
rect -27745 4137 -27711 4166
rect -27671 4137 -27637 4166
rect -27597 4137 -27563 4166
rect -27523 4137 -27489 4166
rect -27449 4137 -27415 4166
rect -27375 4137 -27341 4166
rect -27301 4137 -27267 4166
rect -27227 4137 -27193 4166
rect -27153 4137 -27119 4166
rect -32344 4103 -32315 4113
rect -32315 4103 -32310 4113
rect -32266 4103 -32247 4113
rect -32247 4103 -32232 4113
rect -32188 4103 -32179 4113
rect -32179 4103 -32154 4113
rect -32110 4103 -32077 4113
rect -32077 4103 -32076 4113
rect -32032 4103 -32009 4113
rect -32009 4103 -31998 4113
rect -31954 4103 -31941 4113
rect -31941 4103 -31920 4113
rect -31876 4103 -31873 4113
rect -31873 4103 -31842 4113
rect -31798 4103 -31771 4113
rect -31771 4103 -31764 4113
rect -31718 4103 -31703 4117
rect -31703 4103 -31684 4117
rect -32344 4079 -32310 4103
rect -32266 4079 -32232 4103
rect -32188 4079 -32154 4103
rect -32110 4079 -32076 4103
rect -32032 4079 -31998 4103
rect -31954 4079 -31920 4103
rect -31876 4079 -31842 4103
rect -31798 4079 -31764 4103
rect -31718 4083 -31684 4103
rect -31645 4102 -31632 4117
rect -31632 4102 -31611 4117
rect -31572 4102 -31563 4117
rect -31563 4102 -31538 4117
rect -31499 4102 -31494 4117
rect -31494 4102 -31465 4117
rect -31426 4102 -31425 4117
rect -31425 4102 -31392 4117
rect -31353 4102 -31322 4117
rect -31322 4102 -31319 4117
rect -31280 4102 -31253 4117
rect -31253 4102 -31246 4117
rect -31207 4102 -31184 4117
rect -31184 4102 -31173 4117
rect -31134 4102 -31115 4117
rect -31115 4102 -31100 4117
rect -31061 4102 -31046 4117
rect -31046 4102 -31027 4117
rect -30988 4102 -30977 4117
rect -30977 4102 -30954 4117
rect -30915 4102 -30908 4117
rect -30908 4102 -30881 4117
rect -30842 4102 -30839 4117
rect -30839 4102 -30808 4117
rect -30768 4102 -30735 4117
rect -30735 4102 -30734 4117
rect -30694 4102 -30666 4117
rect -30666 4102 -30660 4117
rect -30620 4102 -30597 4117
rect -30597 4102 -30586 4117
rect -30546 4102 -30528 4117
rect -30528 4102 -30512 4117
rect -30472 4102 -30459 4117
rect -30459 4102 -30438 4117
rect -30398 4102 -30390 4117
rect -30390 4102 -30364 4117
rect -30324 4102 -30321 4117
rect -30321 4102 -30290 4117
rect -30250 4102 -30218 4117
rect -30218 4102 -30216 4117
rect -30176 4102 -30149 4117
rect -30149 4102 -30142 4117
rect -30102 4102 -30080 4117
rect -30080 4102 -30068 4117
rect -30028 4102 -30011 4117
rect -30011 4102 -29994 4117
rect -29954 4102 -29942 4117
rect -29942 4102 -29920 4117
rect -29880 4102 -29873 4117
rect -29873 4102 -29846 4117
rect -29806 4102 -29804 4117
rect -29804 4102 -29772 4117
rect -29732 4102 -29700 4117
rect -29700 4102 -29698 4117
rect -29658 4102 -29631 4117
rect -29631 4102 -29624 4117
rect -29584 4102 -29562 4117
rect -29562 4102 -29550 4117
rect -29510 4102 -29493 4117
rect -29493 4102 -29476 4117
rect -29436 4102 -29424 4117
rect -29424 4102 -29402 4117
rect -29362 4102 -29355 4117
rect -29355 4102 -29328 4117
rect -29288 4102 -29286 4117
rect -29286 4102 -29254 4117
rect -29214 4102 -29183 4117
rect -29183 4102 -29180 4117
rect -29134 4102 -29114 4114
rect -29114 4102 -29100 4114
rect -29046 4103 -29044 4114
rect -29044 4103 -29012 4114
rect -28958 4103 -28942 4114
rect -28942 4103 -28924 4114
rect -28870 4103 -28840 4114
rect -28840 4103 -28836 4114
rect -28189 4132 -28160 4137
rect -28160 4132 -28155 4137
rect -28115 4132 -28092 4137
rect -28092 4132 -28081 4137
rect -28041 4132 -28024 4137
rect -28024 4132 -28007 4137
rect -27967 4132 -27956 4137
rect -27956 4132 -27933 4137
rect -27893 4132 -27888 4137
rect -27888 4132 -27859 4137
rect -27819 4132 -27786 4137
rect -27786 4132 -27785 4137
rect -27745 4132 -27718 4137
rect -27718 4132 -27711 4137
rect -27671 4132 -27650 4137
rect -27650 4132 -27637 4137
rect -27597 4132 -27582 4137
rect -27582 4132 -27563 4137
rect -27523 4132 -27514 4137
rect -27514 4132 -27489 4137
rect -27449 4132 -27446 4137
rect -27446 4132 -27415 4137
rect -27375 4132 -27344 4137
rect -27344 4132 -27341 4137
rect -27301 4132 -27276 4137
rect -27276 4132 -27267 4137
rect -27227 4132 -27208 4137
rect -27208 4132 -27193 4137
rect -27153 4132 -27140 4137
rect -27140 4132 -27119 4137
rect -31645 4083 -31611 4102
rect -31572 4083 -31538 4102
rect -31499 4083 -31465 4102
rect -31426 4083 -31392 4102
rect -31353 4083 -31319 4102
rect -31280 4083 -31246 4102
rect -31207 4083 -31173 4102
rect -31134 4083 -31100 4102
rect -31061 4083 -31027 4102
rect -30988 4083 -30954 4102
rect -30915 4083 -30881 4102
rect -30842 4083 -30808 4102
rect -30768 4083 -30734 4102
rect -30694 4083 -30660 4102
rect -30620 4083 -30586 4102
rect -30546 4083 -30512 4102
rect -30472 4083 -30438 4102
rect -30398 4083 -30364 4102
rect -30324 4083 -30290 4102
rect -30250 4083 -30216 4102
rect -30176 4083 -30142 4102
rect -30102 4083 -30068 4102
rect -30028 4083 -29994 4102
rect -29954 4083 -29920 4102
rect -29880 4083 -29846 4102
rect -29806 4083 -29772 4102
rect -29732 4083 -29698 4102
rect -29658 4083 -29624 4102
rect -29584 4083 -29550 4102
rect -29510 4083 -29476 4102
rect -29436 4083 -29402 4102
rect -29362 4083 -29328 4102
rect -29288 4083 -29254 4102
rect -29214 4083 -29180 4102
rect -29134 4080 -29100 4102
rect -29046 4080 -29012 4103
rect -28958 4080 -28924 4103
rect -28870 4080 -28836 4103
rect -28189 4068 -28155 4093
rect -28115 4068 -28081 4093
rect -28041 4068 -28007 4093
rect -27967 4068 -27933 4093
rect -27893 4068 -27859 4093
rect -27819 4068 -27785 4093
rect -27745 4068 -27711 4093
rect -27671 4068 -27637 4093
rect -27597 4068 -27563 4093
rect -27523 4068 -27489 4093
rect -27449 4068 -27415 4093
rect -27375 4068 -27341 4093
rect -27301 4068 -27267 4093
rect -27227 4068 -27193 4093
rect -27153 4068 -27119 4093
rect -32344 4034 -32315 4040
rect -32315 4034 -32310 4040
rect -32266 4034 -32247 4040
rect -32247 4034 -32232 4040
rect -32188 4034 -32179 4040
rect -32179 4034 -32154 4040
rect -32110 4034 -32077 4040
rect -32077 4034 -32076 4040
rect -32032 4034 -32009 4040
rect -32009 4034 -31998 4040
rect -31954 4034 -31941 4040
rect -31941 4034 -31920 4040
rect -31876 4034 -31873 4040
rect -31873 4034 -31842 4040
rect -31798 4034 -31771 4040
rect -31771 4034 -31764 4040
rect -31718 4034 -31703 4045
rect -31703 4034 -31684 4045
rect -32344 4006 -32310 4034
rect -32266 4006 -32232 4034
rect -32188 4006 -32154 4034
rect -32110 4006 -32076 4034
rect -32032 4006 -31998 4034
rect -31954 4006 -31920 4034
rect -31876 4006 -31842 4034
rect -31798 4006 -31764 4034
rect -31718 4011 -31684 4034
rect -31645 4032 -31632 4045
rect -31632 4032 -31611 4045
rect -31572 4032 -31563 4045
rect -31563 4032 -31538 4045
rect -31499 4032 -31494 4045
rect -31494 4032 -31465 4045
rect -31426 4032 -31425 4045
rect -31425 4032 -31392 4045
rect -31353 4032 -31322 4045
rect -31322 4032 -31319 4045
rect -31280 4032 -31253 4045
rect -31253 4032 -31246 4045
rect -31207 4032 -31184 4045
rect -31184 4032 -31173 4045
rect -31134 4032 -31115 4045
rect -31115 4032 -31100 4045
rect -31061 4032 -31046 4045
rect -31046 4032 -31027 4045
rect -30988 4032 -30977 4045
rect -30977 4032 -30954 4045
rect -30915 4032 -30908 4045
rect -30908 4032 -30881 4045
rect -30842 4032 -30839 4045
rect -30839 4032 -30808 4045
rect -30768 4032 -30735 4045
rect -30735 4032 -30734 4045
rect -30694 4032 -30666 4045
rect -30666 4032 -30660 4045
rect -30620 4032 -30597 4045
rect -30597 4032 -30586 4045
rect -30546 4032 -30528 4045
rect -30528 4032 -30512 4045
rect -30472 4032 -30459 4045
rect -30459 4032 -30438 4045
rect -30398 4032 -30390 4045
rect -30390 4032 -30364 4045
rect -30324 4032 -30321 4045
rect -30321 4032 -30290 4045
rect -30250 4032 -30218 4045
rect -30218 4032 -30216 4045
rect -30176 4032 -30149 4045
rect -30149 4032 -30142 4045
rect -30102 4032 -30080 4045
rect -30080 4032 -30068 4045
rect -30028 4032 -30011 4045
rect -30011 4032 -29994 4045
rect -29954 4032 -29942 4045
rect -29942 4032 -29920 4045
rect -29880 4032 -29873 4045
rect -29873 4032 -29846 4045
rect -29806 4032 -29804 4045
rect -29804 4032 -29772 4045
rect -29732 4032 -29700 4045
rect -29700 4032 -29698 4045
rect -29658 4032 -29631 4045
rect -29631 4032 -29624 4045
rect -29584 4032 -29562 4045
rect -29562 4032 -29550 4045
rect -29510 4032 -29493 4045
rect -29493 4032 -29476 4045
rect -29436 4032 -29424 4045
rect -29424 4032 -29402 4045
rect -29362 4032 -29355 4045
rect -29355 4032 -29328 4045
rect -29288 4032 -29286 4045
rect -29286 4032 -29254 4045
rect -29214 4032 -29183 4045
rect -29183 4032 -29180 4045
rect -29134 4032 -29114 4041
rect -29114 4032 -29100 4041
rect -29046 4034 -29044 4041
rect -29044 4034 -29012 4041
rect -28958 4034 -28942 4041
rect -28942 4034 -28924 4041
rect -28870 4034 -28840 4041
rect -28840 4034 -28836 4041
rect -28189 4059 -28160 4068
rect -28160 4059 -28155 4068
rect -28115 4059 -28092 4068
rect -28092 4059 -28081 4068
rect -28041 4059 -28024 4068
rect -28024 4059 -28007 4068
rect -27967 4059 -27956 4068
rect -27956 4059 -27933 4068
rect -27893 4059 -27888 4068
rect -27888 4059 -27859 4068
rect -27819 4059 -27786 4068
rect -27786 4059 -27785 4068
rect -27745 4059 -27718 4068
rect -27718 4059 -27711 4068
rect -27671 4059 -27650 4068
rect -27650 4059 -27637 4068
rect -27597 4059 -27582 4068
rect -27582 4059 -27563 4068
rect -27523 4059 -27514 4068
rect -27514 4059 -27489 4068
rect -27449 4059 -27446 4068
rect -27446 4059 -27415 4068
rect -27375 4059 -27344 4068
rect -27344 4059 -27341 4068
rect -27301 4059 -27276 4068
rect -27276 4059 -27267 4068
rect -27227 4059 -27208 4068
rect -27208 4059 -27193 4068
rect -27153 4059 -27140 4068
rect -27140 4059 -27119 4068
rect -31645 4011 -31611 4032
rect -31572 4011 -31538 4032
rect -31499 4011 -31465 4032
rect -31426 4011 -31392 4032
rect -31353 4011 -31319 4032
rect -31280 4011 -31246 4032
rect -31207 4011 -31173 4032
rect -31134 4011 -31100 4032
rect -31061 4011 -31027 4032
rect -30988 4011 -30954 4032
rect -30915 4011 -30881 4032
rect -30842 4011 -30808 4032
rect -30768 4011 -30734 4032
rect -30694 4011 -30660 4032
rect -30620 4011 -30586 4032
rect -30546 4011 -30512 4032
rect -30472 4011 -30438 4032
rect -30398 4011 -30364 4032
rect -30324 4011 -30290 4032
rect -30250 4011 -30216 4032
rect -30176 4011 -30142 4032
rect -30102 4011 -30068 4032
rect -30028 4011 -29994 4032
rect -29954 4011 -29920 4032
rect -29880 4011 -29846 4032
rect -29806 4011 -29772 4032
rect -29732 4011 -29698 4032
rect -29658 4011 -29624 4032
rect -29584 4011 -29550 4032
rect -29510 4011 -29476 4032
rect -29436 4011 -29402 4032
rect -29362 4011 -29328 4032
rect -29288 4011 -29254 4032
rect -29214 4011 -29180 4032
rect -29134 4007 -29100 4032
rect -29046 4007 -29012 4034
rect -28958 4007 -28924 4034
rect -28870 4007 -28836 4034
rect -28189 3999 -28155 4020
rect -28115 3999 -28081 4020
rect -28041 3999 -28007 4020
rect -27967 3999 -27933 4020
rect -27893 3999 -27859 4020
rect -27819 3999 -27785 4020
rect -27745 3999 -27711 4020
rect -27671 3999 -27637 4020
rect -27597 3999 -27563 4020
rect -27523 3999 -27489 4020
rect -27449 3999 -27415 4020
rect -27375 3999 -27341 4020
rect -27301 3999 -27267 4020
rect -27227 3999 -27193 4020
rect -27153 3999 -27119 4020
rect -32344 3933 -32315 3967
rect -32315 3933 -32310 3967
rect -32266 3933 -32232 3967
rect -32188 3933 -32154 3967
rect -32110 3933 -32076 3967
rect -32032 3933 -31998 3967
rect -31954 3933 -31920 3967
rect -31876 3933 -31842 3967
rect -31798 3933 -31764 3967
rect -31718 3939 -31684 3973
rect -31645 3962 -31632 3973
rect -31632 3962 -31611 3973
rect -31572 3962 -31563 3973
rect -31563 3962 -31538 3973
rect -31499 3962 -31494 3973
rect -31494 3962 -31465 3973
rect -31426 3962 -31425 3973
rect -31425 3962 -31392 3973
rect -31353 3962 -31322 3973
rect -31322 3962 -31319 3973
rect -31280 3962 -31253 3973
rect -31253 3962 -31246 3973
rect -31207 3962 -31184 3973
rect -31184 3962 -31173 3973
rect -31134 3962 -31115 3973
rect -31115 3962 -31100 3973
rect -31061 3962 -31046 3973
rect -31046 3962 -31027 3973
rect -30988 3962 -30977 3973
rect -30977 3962 -30954 3973
rect -30915 3962 -30908 3973
rect -30908 3962 -30881 3973
rect -30842 3962 -30839 3973
rect -30839 3962 -30808 3973
rect -30768 3962 -30735 3973
rect -30735 3962 -30734 3973
rect -30694 3962 -30666 3973
rect -30666 3962 -30660 3973
rect -30620 3962 -30597 3973
rect -30597 3962 -30586 3973
rect -30546 3962 -30528 3973
rect -30528 3962 -30512 3973
rect -30472 3962 -30459 3973
rect -30459 3962 -30438 3973
rect -30398 3962 -30390 3973
rect -30390 3962 -30364 3973
rect -30324 3962 -30321 3973
rect -30321 3962 -30290 3973
rect -30250 3962 -30218 3973
rect -30218 3962 -30216 3973
rect -30176 3962 -30149 3973
rect -30149 3962 -30142 3973
rect -30102 3962 -30080 3973
rect -30080 3962 -30068 3973
rect -30028 3962 -30011 3973
rect -30011 3962 -29994 3973
rect -29954 3962 -29942 3973
rect -29942 3962 -29920 3973
rect -29880 3962 -29873 3973
rect -29873 3962 -29846 3973
rect -29806 3962 -29804 3973
rect -29804 3962 -29772 3973
rect -29732 3962 -29700 3973
rect -29700 3962 -29698 3973
rect -29658 3962 -29631 3973
rect -29631 3962 -29624 3973
rect -29584 3962 -29562 3973
rect -29562 3962 -29550 3973
rect -29510 3962 -29493 3973
rect -29493 3962 -29476 3973
rect -29436 3962 -29424 3973
rect -29424 3962 -29402 3973
rect -29362 3962 -29355 3973
rect -29355 3962 -29328 3973
rect -29288 3962 -29286 3973
rect -29286 3962 -29254 3973
rect -29214 3962 -29183 3973
rect -29183 3962 -29180 3973
rect -29134 3962 -29114 3968
rect -29114 3962 -29100 3968
rect -29046 3965 -29044 3968
rect -29044 3965 -29012 3968
rect -28958 3965 -28942 3968
rect -28942 3965 -28924 3968
rect -28870 3965 -28840 3968
rect -28840 3965 -28836 3968
rect -28189 3986 -28160 3999
rect -28160 3986 -28155 3999
rect -28115 3986 -28092 3999
rect -28092 3986 -28081 3999
rect -28041 3986 -28024 3999
rect -28024 3986 -28007 3999
rect -27967 3986 -27956 3999
rect -27956 3986 -27933 3999
rect -27893 3986 -27888 3999
rect -27888 3986 -27859 3999
rect -27819 3986 -27786 3999
rect -27786 3986 -27785 3999
rect -27745 3986 -27718 3999
rect -27718 3986 -27711 3999
rect -27671 3986 -27650 3999
rect -27650 3986 -27637 3999
rect -27597 3986 -27582 3999
rect -27582 3986 -27563 3999
rect -27523 3986 -27514 3999
rect -27514 3986 -27489 3999
rect -27449 3986 -27446 3999
rect -27446 3986 -27415 3999
rect -27375 3986 -27344 3999
rect -27344 3986 -27341 3999
rect -27301 3986 -27276 3999
rect -27276 3986 -27267 3999
rect -27227 3986 -27208 3999
rect -27208 3986 -27193 3999
rect -27153 3986 -27140 3999
rect -27140 3986 -27119 3999
rect -31645 3939 -31611 3962
rect -31572 3939 -31538 3962
rect -31499 3939 -31465 3962
rect -31426 3939 -31392 3962
rect -31353 3939 -31319 3962
rect -31280 3939 -31246 3962
rect -31207 3939 -31173 3962
rect -31134 3939 -31100 3962
rect -31061 3939 -31027 3962
rect -30988 3939 -30954 3962
rect -30915 3939 -30881 3962
rect -30842 3939 -30808 3962
rect -30768 3939 -30734 3962
rect -30694 3939 -30660 3962
rect -30620 3939 -30586 3962
rect -30546 3939 -30512 3962
rect -30472 3939 -30438 3962
rect -30398 3939 -30364 3962
rect -30324 3939 -30290 3962
rect -30250 3939 -30216 3962
rect -30176 3939 -30142 3962
rect -30102 3939 -30068 3962
rect -30028 3939 -29994 3962
rect -29954 3939 -29920 3962
rect -29880 3939 -29846 3962
rect -29806 3939 -29772 3962
rect -29732 3939 -29698 3962
rect -29658 3939 -29624 3962
rect -29584 3939 -29550 3962
rect -29510 3939 -29476 3962
rect -29436 3939 -29402 3962
rect -29362 3939 -29328 3962
rect -29288 3939 -29254 3962
rect -29214 3939 -29180 3962
rect -29134 3934 -29100 3962
rect -29046 3934 -29012 3965
rect -28958 3934 -28924 3965
rect -28870 3934 -28836 3965
rect -28189 3930 -28155 3947
rect -28115 3930 -28081 3947
rect -28041 3930 -28007 3947
rect -27967 3930 -27933 3947
rect -27893 3930 -27859 3947
rect -27819 3930 -27785 3947
rect -27745 3930 -27711 3947
rect -27671 3930 -27637 3947
rect -27597 3930 -27563 3947
rect -27523 3930 -27489 3947
rect -27449 3930 -27415 3947
rect -27375 3930 -27341 3947
rect -27301 3930 -27267 3947
rect -27227 3930 -27193 3947
rect -27153 3930 -27119 3947
rect -32344 3860 -32315 3894
rect -32315 3860 -32310 3894
rect -32266 3860 -32232 3894
rect -32188 3860 -32154 3894
rect -32110 3860 -32076 3894
rect -32032 3860 -31998 3894
rect -31954 3860 -31920 3894
rect -31876 3860 -31842 3894
rect -31798 3860 -31764 3894
rect -31718 3867 -31684 3901
rect -31645 3892 -31632 3901
rect -31632 3892 -31611 3901
rect -31572 3892 -31563 3901
rect -31563 3892 -31538 3901
rect -31499 3892 -31494 3901
rect -31494 3892 -31465 3901
rect -31426 3892 -31425 3901
rect -31425 3892 -31392 3901
rect -31353 3892 -31322 3901
rect -31322 3892 -31319 3901
rect -31280 3892 -31253 3901
rect -31253 3892 -31246 3901
rect -31207 3892 -31184 3901
rect -31184 3892 -31173 3901
rect -31134 3892 -31115 3901
rect -31115 3892 -31100 3901
rect -31061 3892 -31046 3901
rect -31046 3892 -31027 3901
rect -30988 3892 -30977 3901
rect -30977 3892 -30954 3901
rect -30915 3892 -30908 3901
rect -30908 3892 -30881 3901
rect -30842 3892 -30839 3901
rect -30839 3892 -30808 3901
rect -30768 3892 -30735 3901
rect -30735 3892 -30734 3901
rect -30694 3892 -30666 3901
rect -30666 3892 -30660 3901
rect -30620 3892 -30597 3901
rect -30597 3892 -30586 3901
rect -30546 3892 -30528 3901
rect -30528 3892 -30512 3901
rect -30472 3892 -30459 3901
rect -30459 3892 -30438 3901
rect -30398 3892 -30390 3901
rect -30390 3892 -30364 3901
rect -30324 3892 -30321 3901
rect -30321 3892 -30290 3901
rect -30250 3892 -30218 3901
rect -30218 3892 -30216 3901
rect -30176 3892 -30149 3901
rect -30149 3892 -30142 3901
rect -30102 3892 -30080 3901
rect -30080 3892 -30068 3901
rect -30028 3892 -30011 3901
rect -30011 3892 -29994 3901
rect -29954 3892 -29942 3901
rect -29942 3892 -29920 3901
rect -29880 3892 -29873 3901
rect -29873 3892 -29846 3901
rect -29806 3892 -29804 3901
rect -29804 3892 -29772 3901
rect -29732 3892 -29700 3901
rect -29700 3892 -29698 3901
rect -29658 3892 -29631 3901
rect -29631 3892 -29624 3901
rect -29584 3892 -29562 3901
rect -29562 3892 -29550 3901
rect -29510 3892 -29493 3901
rect -29493 3892 -29476 3901
rect -29436 3892 -29424 3901
rect -29424 3892 -29402 3901
rect -29362 3892 -29355 3901
rect -29355 3892 -29328 3901
rect -29288 3892 -29286 3901
rect -29286 3892 -29254 3901
rect -29214 3892 -29183 3901
rect -29183 3892 -29180 3901
rect -28189 3913 -28160 3930
rect -28160 3913 -28155 3930
rect -28115 3913 -28092 3930
rect -28092 3913 -28081 3930
rect -28041 3913 -28024 3930
rect -28024 3913 -28007 3930
rect -27967 3913 -27956 3930
rect -27956 3913 -27933 3930
rect -27893 3913 -27888 3930
rect -27888 3913 -27859 3930
rect -27819 3913 -27786 3930
rect -27786 3913 -27785 3930
rect -27745 3913 -27718 3930
rect -27718 3913 -27711 3930
rect -27671 3913 -27650 3930
rect -27650 3913 -27637 3930
rect -27597 3913 -27582 3930
rect -27582 3913 -27563 3930
rect -27523 3913 -27514 3930
rect -27514 3913 -27489 3930
rect -27449 3913 -27446 3930
rect -27446 3913 -27415 3930
rect -27375 3913 -27344 3930
rect -27344 3913 -27341 3930
rect -27301 3913 -27276 3930
rect -27276 3913 -27267 3930
rect -27227 3913 -27208 3930
rect -27208 3913 -27193 3930
rect -27153 3913 -27140 3930
rect -27140 3913 -27119 3930
rect -29134 3892 -29114 3895
rect -29114 3892 -29100 3895
rect -31645 3867 -31611 3892
rect -31572 3867 -31538 3892
rect -31499 3867 -31465 3892
rect -31426 3867 -31392 3892
rect -31353 3867 -31319 3892
rect -31280 3867 -31246 3892
rect -31207 3867 -31173 3892
rect -31134 3867 -31100 3892
rect -31061 3867 -31027 3892
rect -30988 3867 -30954 3892
rect -30915 3867 -30881 3892
rect -30842 3867 -30808 3892
rect -30768 3867 -30734 3892
rect -30694 3867 -30660 3892
rect -30620 3867 -30586 3892
rect -30546 3867 -30512 3892
rect -30472 3867 -30438 3892
rect -30398 3867 -30364 3892
rect -30324 3867 -30290 3892
rect -30250 3867 -30216 3892
rect -30176 3867 -30142 3892
rect -30102 3867 -30068 3892
rect -30028 3867 -29994 3892
rect -29954 3867 -29920 3892
rect -29880 3867 -29846 3892
rect -29806 3867 -29772 3892
rect -29732 3867 -29698 3892
rect -29658 3867 -29624 3892
rect -29584 3867 -29550 3892
rect -29510 3867 -29476 3892
rect -29436 3867 -29402 3892
rect -29362 3867 -29328 3892
rect -29288 3867 -29254 3892
rect -29214 3867 -29180 3892
rect -29134 3861 -29100 3892
rect -29046 3861 -29012 3895
rect -28958 3861 -28924 3895
rect -28870 3861 -28836 3895
rect -28189 3861 -28155 3874
rect -28115 3861 -28081 3874
rect -28041 3861 -28007 3874
rect -27967 3861 -27933 3874
rect -27893 3861 -27859 3874
rect -27819 3861 -27785 3874
rect -27745 3861 -27711 3874
rect -27671 3861 -27637 3874
rect -27597 3861 -27563 3874
rect -27523 3861 -27489 3874
rect -27449 3861 -27415 3874
rect -27375 3861 -27341 3874
rect -27301 3861 -27267 3874
rect -27227 3861 -27193 3874
rect -27153 3861 -27119 3874
rect -32344 3787 -32315 3821
rect -32315 3787 -32310 3821
rect -32266 3787 -32232 3821
rect -32188 3787 -32154 3821
rect -32110 3787 -32076 3821
rect -32032 3787 -31998 3821
rect -31954 3787 -31920 3821
rect -31876 3787 -31842 3821
rect -31798 3787 -31764 3821
rect -31718 3795 -31684 3829
rect -31645 3822 -31632 3829
rect -31632 3822 -31611 3829
rect -31572 3822 -31563 3829
rect -31563 3822 -31538 3829
rect -31499 3822 -31494 3829
rect -31494 3822 -31465 3829
rect -31426 3822 -31425 3829
rect -31425 3822 -31392 3829
rect -31353 3822 -31322 3829
rect -31322 3822 -31319 3829
rect -31280 3822 -31253 3829
rect -31253 3822 -31246 3829
rect -31207 3822 -31184 3829
rect -31184 3822 -31173 3829
rect -31134 3822 -31115 3829
rect -31115 3822 -31100 3829
rect -31061 3822 -31046 3829
rect -31046 3822 -31027 3829
rect -30988 3822 -30977 3829
rect -30977 3822 -30954 3829
rect -30915 3822 -30908 3829
rect -30908 3822 -30881 3829
rect -30842 3822 -30839 3829
rect -30839 3822 -30808 3829
rect -30768 3822 -30735 3829
rect -30735 3822 -30734 3829
rect -30694 3822 -30666 3829
rect -30666 3822 -30660 3829
rect -30620 3822 -30597 3829
rect -30597 3822 -30586 3829
rect -30546 3822 -30528 3829
rect -30528 3822 -30512 3829
rect -30472 3822 -30459 3829
rect -30459 3822 -30438 3829
rect -30398 3822 -30390 3829
rect -30390 3822 -30364 3829
rect -30324 3822 -30321 3829
rect -30321 3822 -30290 3829
rect -30250 3822 -30218 3829
rect -30218 3822 -30216 3829
rect -30176 3822 -30149 3829
rect -30149 3822 -30142 3829
rect -30102 3822 -30080 3829
rect -30080 3822 -30068 3829
rect -30028 3822 -30011 3829
rect -30011 3822 -29994 3829
rect -29954 3822 -29942 3829
rect -29942 3822 -29920 3829
rect -29880 3822 -29873 3829
rect -29873 3822 -29846 3829
rect -29806 3822 -29804 3829
rect -29804 3822 -29772 3829
rect -29732 3822 -29700 3829
rect -29700 3822 -29698 3829
rect -29658 3822 -29631 3829
rect -29631 3822 -29624 3829
rect -29584 3822 -29562 3829
rect -29562 3822 -29550 3829
rect -29510 3822 -29493 3829
rect -29493 3822 -29476 3829
rect -29436 3822 -29424 3829
rect -29424 3822 -29402 3829
rect -29362 3822 -29355 3829
rect -29355 3822 -29328 3829
rect -29288 3822 -29286 3829
rect -29286 3822 -29254 3829
rect -29214 3822 -29183 3829
rect -29183 3822 -29180 3829
rect -28189 3840 -28160 3861
rect -28160 3840 -28155 3861
rect -28115 3840 -28092 3861
rect -28092 3840 -28081 3861
rect -28041 3840 -28024 3861
rect -28024 3840 -28007 3861
rect -27967 3840 -27956 3861
rect -27956 3840 -27933 3861
rect -27893 3840 -27888 3861
rect -27888 3840 -27859 3861
rect -27819 3840 -27786 3861
rect -27786 3840 -27785 3861
rect -27745 3840 -27718 3861
rect -27718 3840 -27711 3861
rect -27671 3840 -27650 3861
rect -27650 3840 -27637 3861
rect -27597 3840 -27582 3861
rect -27582 3840 -27563 3861
rect -27523 3840 -27514 3861
rect -27514 3840 -27489 3861
rect -27449 3840 -27446 3861
rect -27446 3840 -27415 3861
rect -27375 3840 -27344 3861
rect -27344 3840 -27341 3861
rect -27301 3840 -27276 3861
rect -27276 3840 -27267 3861
rect -27227 3840 -27208 3861
rect -27208 3840 -27193 3861
rect -27153 3840 -27140 3861
rect -27140 3840 -27119 3861
rect -31645 3795 -31611 3822
rect -31572 3795 -31538 3822
rect -31499 3795 -31465 3822
rect -31426 3795 -31392 3822
rect -31353 3795 -31319 3822
rect -31280 3795 -31246 3822
rect -31207 3795 -31173 3822
rect -31134 3795 -31100 3822
rect -31061 3795 -31027 3822
rect -30988 3795 -30954 3822
rect -30915 3795 -30881 3822
rect -30842 3795 -30808 3822
rect -30768 3795 -30734 3822
rect -30694 3795 -30660 3822
rect -30620 3795 -30586 3822
rect -30546 3795 -30512 3822
rect -30472 3795 -30438 3822
rect -30398 3795 -30364 3822
rect -30324 3795 -30290 3822
rect -30250 3795 -30216 3822
rect -30176 3795 -30142 3822
rect -30102 3795 -30068 3822
rect -30028 3795 -29994 3822
rect -29954 3795 -29920 3822
rect -29880 3795 -29846 3822
rect -29806 3795 -29772 3822
rect -29732 3795 -29698 3822
rect -29658 3795 -29624 3822
rect -29584 3795 -29550 3822
rect -29510 3795 -29476 3822
rect -29436 3795 -29402 3822
rect -29362 3795 -29328 3822
rect -29288 3795 -29254 3822
rect -29214 3795 -29180 3822
rect -29134 3788 -29100 3822
rect -29046 3792 -29012 3822
rect -28958 3792 -28924 3822
rect -28870 3792 -28836 3822
rect -28189 3792 -28155 3801
rect -28115 3792 -28081 3801
rect -28041 3792 -28007 3801
rect -27967 3792 -27933 3801
rect -27893 3792 -27859 3801
rect -27819 3792 -27785 3801
rect -27745 3792 -27711 3801
rect -27671 3792 -27637 3801
rect -27597 3792 -27563 3801
rect -27523 3792 -27489 3801
rect -27449 3792 -27415 3801
rect -27375 3792 -27341 3801
rect -27301 3792 -27267 3801
rect -27227 3792 -27193 3801
rect -27153 3792 -27119 3801
rect -29046 3788 -29044 3792
rect -29044 3788 -29012 3792
rect -32344 3714 -32315 3748
rect -32315 3714 -32310 3748
rect -32266 3714 -32232 3748
rect -32188 3714 -32154 3748
rect -32110 3714 -32076 3748
rect -32032 3714 -31998 3748
rect -31954 3714 -31920 3748
rect -31876 3714 -31842 3748
rect -31798 3714 -31764 3748
rect -31718 3723 -31684 3757
rect -31645 3752 -31632 3757
rect -31632 3752 -31611 3757
rect -31572 3752 -31563 3757
rect -31563 3752 -31538 3757
rect -31499 3752 -31494 3757
rect -31494 3752 -31465 3757
rect -31426 3752 -31425 3757
rect -31425 3752 -31392 3757
rect -31353 3752 -31322 3757
rect -31322 3752 -31319 3757
rect -31280 3752 -31253 3757
rect -31253 3752 -31246 3757
rect -31207 3752 -31184 3757
rect -31184 3752 -31173 3757
rect -31134 3752 -31115 3757
rect -31115 3752 -31100 3757
rect -31061 3752 -31046 3757
rect -31046 3752 -31027 3757
rect -30988 3752 -30977 3757
rect -30977 3752 -30954 3757
rect -30915 3752 -30908 3757
rect -30908 3752 -30881 3757
rect -30842 3752 -30839 3757
rect -30839 3752 -30808 3757
rect -30768 3752 -30735 3757
rect -30735 3752 -30734 3757
rect -30694 3752 -30666 3757
rect -30666 3752 -30660 3757
rect -30620 3752 -30597 3757
rect -30597 3752 -30586 3757
rect -30546 3752 -30528 3757
rect -30528 3752 -30512 3757
rect -30472 3752 -30459 3757
rect -30459 3752 -30438 3757
rect -30398 3752 -30390 3757
rect -30390 3752 -30364 3757
rect -30324 3752 -30321 3757
rect -30321 3752 -30290 3757
rect -30250 3752 -30218 3757
rect -30218 3752 -30216 3757
rect -30176 3752 -30149 3757
rect -30149 3752 -30142 3757
rect -30102 3752 -30080 3757
rect -30080 3752 -30068 3757
rect -30028 3752 -30011 3757
rect -30011 3752 -29994 3757
rect -29954 3752 -29942 3757
rect -29942 3752 -29920 3757
rect -29880 3752 -29873 3757
rect -29873 3752 -29846 3757
rect -29806 3752 -29804 3757
rect -29804 3752 -29772 3757
rect -29732 3752 -29700 3757
rect -29700 3752 -29698 3757
rect -29658 3752 -29631 3757
rect -29631 3752 -29624 3757
rect -29584 3752 -29562 3757
rect -29562 3752 -29550 3757
rect -29510 3752 -29493 3757
rect -29493 3752 -29476 3757
rect -29436 3752 -29424 3757
rect -29424 3752 -29402 3757
rect -29362 3752 -29355 3757
rect -29355 3752 -29328 3757
rect -29288 3752 -29286 3757
rect -29286 3752 -29254 3757
rect -29214 3752 -29183 3757
rect -29183 3752 -29180 3757
rect -28958 3788 -28942 3792
rect -28942 3788 -28924 3792
rect -28870 3788 -28840 3792
rect -28840 3788 -28836 3792
rect -28189 3767 -28160 3792
rect -28160 3767 -28155 3792
rect -28115 3767 -28092 3792
rect -28092 3767 -28081 3792
rect -28041 3767 -28024 3792
rect -28024 3767 -28007 3792
rect -27967 3767 -27956 3792
rect -27956 3767 -27933 3792
rect -27893 3767 -27888 3792
rect -27888 3767 -27859 3792
rect -27819 3767 -27786 3792
rect -27786 3767 -27785 3792
rect -27745 3767 -27718 3792
rect -27718 3767 -27711 3792
rect -27671 3767 -27650 3792
rect -27650 3767 -27637 3792
rect -27597 3767 -27582 3792
rect -27582 3767 -27563 3792
rect -27523 3767 -27514 3792
rect -27514 3767 -27489 3792
rect -27449 3767 -27446 3792
rect -27446 3767 -27415 3792
rect -27375 3767 -27344 3792
rect -27344 3767 -27341 3792
rect -27301 3767 -27276 3792
rect -27276 3767 -27267 3792
rect -27227 3767 -27208 3792
rect -27208 3767 -27193 3792
rect -27153 3767 -27140 3792
rect -27140 3767 -27119 3792
rect -31645 3723 -31611 3752
rect -31572 3723 -31538 3752
rect -31499 3723 -31465 3752
rect -31426 3723 -31392 3752
rect -31353 3723 -31319 3752
rect -31280 3723 -31246 3752
rect -31207 3723 -31173 3752
rect -31134 3723 -31100 3752
rect -31061 3723 -31027 3752
rect -30988 3723 -30954 3752
rect -30915 3723 -30881 3752
rect -30842 3723 -30808 3752
rect -30768 3723 -30734 3752
rect -30694 3723 -30660 3752
rect -30620 3723 -30586 3752
rect -30546 3723 -30512 3752
rect -30472 3723 -30438 3752
rect -30398 3723 -30364 3752
rect -30324 3723 -30290 3752
rect -30250 3723 -30216 3752
rect -30176 3723 -30142 3752
rect -30102 3723 -30068 3752
rect -30028 3723 -29994 3752
rect -29954 3723 -29920 3752
rect -29880 3723 -29846 3752
rect -29806 3723 -29772 3752
rect -29732 3723 -29698 3752
rect -29658 3723 -29624 3752
rect -29584 3723 -29550 3752
rect -29510 3723 -29476 3752
rect -29436 3723 -29402 3752
rect -29362 3723 -29328 3752
rect -29288 3723 -29254 3752
rect -29214 3723 -29180 3752
rect -29134 3716 -29100 3749
rect -29046 3723 -29012 3749
rect -28958 3723 -28924 3749
rect -28870 3723 -28836 3749
rect -28189 3723 -28155 3728
rect -28115 3723 -28081 3728
rect -28041 3723 -28007 3728
rect -27967 3723 -27933 3728
rect -27893 3723 -27859 3728
rect -27819 3723 -27785 3728
rect -27745 3723 -27711 3728
rect -27671 3723 -27637 3728
rect -27597 3723 -27563 3728
rect -27523 3723 -27489 3728
rect -27449 3723 -27415 3728
rect -27375 3723 -27341 3728
rect -27301 3723 -27267 3728
rect -27227 3723 -27193 3728
rect -27153 3723 -27119 3728
rect -32344 3641 -32315 3675
rect -32315 3641 -32310 3675
rect -32266 3641 -32232 3675
rect -32188 3641 -32154 3675
rect -32110 3641 -32076 3675
rect -32032 3641 -31998 3675
rect -31954 3641 -31920 3675
rect -31876 3641 -31842 3675
rect -31798 3641 -31764 3675
rect -31718 3651 -31684 3685
rect -31645 3682 -31632 3685
rect -31632 3682 -31611 3685
rect -31572 3682 -31563 3685
rect -31563 3682 -31538 3685
rect -31499 3682 -31494 3685
rect -31494 3682 -31465 3685
rect -31426 3682 -31425 3685
rect -31425 3682 -31392 3685
rect -31353 3682 -31322 3685
rect -31322 3682 -31319 3685
rect -31280 3682 -31253 3685
rect -31253 3682 -31246 3685
rect -31207 3682 -31184 3685
rect -31184 3682 -31173 3685
rect -31134 3682 -31115 3685
rect -31115 3682 -31100 3685
rect -31061 3682 -31046 3685
rect -31046 3682 -31027 3685
rect -30988 3682 -30977 3685
rect -30977 3682 -30954 3685
rect -30915 3682 -30908 3685
rect -30908 3682 -30881 3685
rect -30842 3682 -30839 3685
rect -30839 3682 -30808 3685
rect -30768 3682 -30735 3685
rect -30735 3682 -30734 3685
rect -30694 3682 -30666 3685
rect -30666 3682 -30660 3685
rect -30620 3682 -30597 3685
rect -30597 3682 -30586 3685
rect -30546 3682 -30528 3685
rect -30528 3682 -30512 3685
rect -30472 3682 -30459 3685
rect -30459 3682 -30438 3685
rect -30398 3682 -30390 3685
rect -30390 3682 -30364 3685
rect -30324 3682 -30321 3685
rect -30321 3682 -30290 3685
rect -30250 3682 -30218 3685
rect -30218 3682 -30216 3685
rect -30176 3682 -30149 3685
rect -30149 3682 -30142 3685
rect -30102 3682 -30080 3685
rect -30080 3682 -30068 3685
rect -30028 3682 -30011 3685
rect -30011 3682 -29994 3685
rect -29954 3682 -29942 3685
rect -29942 3682 -29920 3685
rect -29880 3682 -29873 3685
rect -29873 3682 -29846 3685
rect -29806 3682 -29804 3685
rect -29804 3682 -29772 3685
rect -29732 3682 -29700 3685
rect -29700 3682 -29698 3685
rect -29658 3682 -29631 3685
rect -29631 3682 -29624 3685
rect -29584 3682 -29562 3685
rect -29562 3682 -29550 3685
rect -29510 3682 -29493 3685
rect -29493 3682 -29476 3685
rect -29436 3682 -29424 3685
rect -29424 3682 -29402 3685
rect -29362 3682 -29355 3685
rect -29355 3682 -29328 3685
rect -29288 3682 -29286 3685
rect -29286 3682 -29254 3685
rect -29134 3715 -29114 3716
rect -29114 3715 -29100 3716
rect -29046 3715 -29044 3723
rect -29044 3715 -29012 3723
rect -29214 3682 -29183 3685
rect -29183 3682 -29180 3685
rect -28958 3715 -28942 3723
rect -28942 3715 -28924 3723
rect -28870 3715 -28840 3723
rect -28840 3715 -28836 3723
rect -28189 3694 -28160 3723
rect -28160 3694 -28155 3723
rect -28115 3694 -28092 3723
rect -28092 3694 -28081 3723
rect -28041 3694 -28024 3723
rect -28024 3694 -28007 3723
rect -27967 3694 -27956 3723
rect -27956 3694 -27933 3723
rect -27893 3694 -27888 3723
rect -27888 3694 -27859 3723
rect -27819 3694 -27786 3723
rect -27786 3694 -27785 3723
rect -27745 3694 -27718 3723
rect -27718 3694 -27711 3723
rect -27671 3694 -27650 3723
rect -27650 3694 -27637 3723
rect -27597 3694 -27582 3723
rect -27582 3694 -27563 3723
rect -27523 3694 -27514 3723
rect -27514 3694 -27489 3723
rect -27449 3694 -27446 3723
rect -27446 3694 -27415 3723
rect -27375 3694 -27344 3723
rect -27344 3694 -27341 3723
rect -27301 3694 -27276 3723
rect -27276 3694 -27267 3723
rect -27227 3694 -27208 3723
rect -27208 3694 -27193 3723
rect -27153 3694 -27140 3723
rect -27140 3694 -27119 3723
rect 4010 3806 4044 3840
rect 4082 3806 4106 3840
rect 4106 3806 4116 3840
rect 4154 3806 4174 3840
rect 4174 3806 4188 3840
rect 4226 3806 4242 3840
rect 4242 3806 4260 3840
rect 4298 3806 4310 3840
rect 4310 3806 4332 3840
rect 4370 3806 4378 3840
rect 4378 3806 4404 3840
rect 4442 3806 4446 3840
rect 4446 3806 4476 3840
rect 4514 3806 4548 3840
rect 4586 3806 4616 3840
rect 4616 3806 4620 3840
rect 4658 3806 4684 3840
rect 4684 3806 4692 3840
rect 4730 3806 4752 3840
rect 4752 3806 4764 3840
rect 4802 3806 4820 3840
rect 4820 3806 4836 3840
rect 4874 3806 4888 3840
rect 4888 3806 4908 3840
rect 4946 3806 4956 3840
rect 4956 3806 4980 3840
rect 5018 3806 5024 3840
rect 5024 3806 5052 3840
rect 5090 3806 5092 3840
rect 5092 3806 5124 3840
rect 5162 3806 5194 3840
rect 5194 3806 5196 3840
rect 5234 3806 5262 3840
rect 5262 3806 5268 3840
rect 5306 3806 5330 3840
rect 5330 3806 5340 3840
rect 5378 3806 5398 3840
rect 5398 3806 5412 3840
rect 5450 3806 5466 3840
rect 5466 3806 5484 3840
rect 5522 3806 5534 3840
rect 5534 3806 5556 3840
rect 5594 3806 5602 3840
rect 5602 3806 5628 3840
rect 5666 3806 5670 3840
rect 5670 3806 5700 3840
rect 3938 3734 3972 3768
rect -31645 3651 -31611 3682
rect -31572 3651 -31538 3682
rect -31499 3651 -31465 3682
rect -31426 3651 -31392 3682
rect -31353 3651 -31319 3682
rect -31280 3651 -31246 3682
rect -31207 3651 -31173 3682
rect -31134 3651 -31100 3682
rect -31061 3651 -31027 3682
rect -30988 3651 -30954 3682
rect -30915 3651 -30881 3682
rect -30842 3651 -30808 3682
rect -30768 3651 -30734 3682
rect -30694 3651 -30660 3682
rect -30620 3651 -30586 3682
rect -30546 3651 -30512 3682
rect -30472 3651 -30438 3682
rect -30398 3651 -30364 3682
rect -30324 3651 -30290 3682
rect -30250 3651 -30216 3682
rect -30176 3651 -30142 3682
rect -30102 3651 -30068 3682
rect -30028 3651 -29994 3682
rect -29954 3651 -29920 3682
rect -29880 3651 -29846 3682
rect -29806 3651 -29772 3682
rect -29732 3651 -29698 3682
rect -29658 3651 -29624 3682
rect -29584 3651 -29550 3682
rect -29510 3651 -29476 3682
rect -29436 3651 -29402 3682
rect -29362 3651 -29328 3682
rect -29288 3651 -29254 3682
rect -29214 3651 -29180 3682
rect -29134 3646 -29100 3676
rect -29046 3654 -29012 3676
rect -28958 3654 -28924 3676
rect -28870 3654 -28836 3676
rect -28189 3654 -28155 3655
rect -28115 3654 -28081 3655
rect -28041 3654 -28007 3655
rect -27967 3654 -27933 3655
rect -27893 3654 -27859 3655
rect -27819 3654 -27785 3655
rect -27745 3654 -27711 3655
rect -27671 3654 -27637 3655
rect -27597 3654 -27563 3655
rect -27523 3654 -27489 3655
rect -27449 3654 -27415 3655
rect -27375 3654 -27341 3655
rect -27301 3654 -27267 3655
rect -27227 3654 -27193 3655
rect -27153 3654 -27119 3655
rect -757 3654 -733 3688
rect -733 3654 -723 3688
rect -677 3654 -662 3688
rect -662 3654 -643 3688
rect -597 3654 -591 3688
rect -591 3654 -563 3688
rect -516 3654 -485 3688
rect -485 3654 -482 3688
rect -435 3654 -413 3688
rect -413 3654 -401 3688
rect 171 3654 181 3688
rect 181 3654 205 3688
rect 244 3654 250 3688
rect 250 3654 278 3688
rect 317 3654 319 3688
rect 319 3654 351 3688
rect 390 3654 422 3688
rect 422 3654 424 3688
rect 463 3654 491 3688
rect 491 3654 497 3688
rect 536 3654 560 3688
rect 560 3654 570 3688
rect 609 3654 629 3688
rect 629 3654 643 3688
rect 682 3654 698 3688
rect 698 3654 716 3688
rect 755 3654 767 3688
rect 767 3654 789 3688
rect 828 3654 836 3688
rect 836 3654 862 3688
rect 901 3654 905 3688
rect 905 3654 935 3688
rect 974 3654 1008 3688
rect 1047 3654 1078 3688
rect 1078 3654 1081 3688
rect 1120 3654 1147 3688
rect 1147 3654 1154 3688
rect 1193 3654 1216 3688
rect 1216 3654 1227 3688
rect 1266 3654 1285 3688
rect 1285 3654 1300 3688
rect 1339 3654 1354 3688
rect 1354 3654 1373 3688
rect 1412 3654 1423 3688
rect 1423 3654 1446 3688
rect 1485 3654 1492 3688
rect 1492 3654 1519 3688
rect 1558 3654 1561 3688
rect 1561 3654 1592 3688
rect 1631 3654 1664 3688
rect 1664 3654 1665 3688
rect 1704 3654 1733 3688
rect 1733 3654 1738 3688
rect 1777 3654 1802 3688
rect 1802 3654 1811 3688
rect 1850 3654 1871 3688
rect 1871 3654 1884 3688
rect 1923 3654 1940 3688
rect 1940 3654 1957 3688
rect 1995 3654 2009 3688
rect 2009 3654 2029 3688
rect 2067 3654 2078 3688
rect 2078 3654 2101 3688
rect 2139 3654 2147 3688
rect 2147 3654 2173 3688
rect 2211 3654 2216 3688
rect 2216 3654 2245 3688
rect 2283 3654 2285 3688
rect 2285 3654 2317 3688
rect 2355 3654 2389 3688
rect 2427 3654 2458 3688
rect 2458 3654 2461 3688
rect 2499 3654 2527 3688
rect 2527 3654 2533 3688
rect 2571 3654 2596 3688
rect 2596 3654 2605 3688
rect 2643 3654 2665 3688
rect 2665 3654 2677 3688
rect 2715 3654 2734 3688
rect 2734 3654 2749 3688
rect 2787 3654 2803 3688
rect 2803 3654 2821 3688
rect 2859 3654 2872 3688
rect 2872 3654 2893 3688
rect 2931 3654 2941 3688
rect 2941 3654 2965 3688
rect 3003 3654 3010 3688
rect 3010 3654 3037 3688
rect 3075 3654 3078 3688
rect 3078 3654 3109 3688
rect 3147 3654 3180 3688
rect 3180 3654 3181 3688
rect 3219 3654 3248 3688
rect 3248 3654 3253 3688
rect 3291 3654 3316 3688
rect 3316 3654 3325 3688
rect 3363 3654 3384 3688
rect 3384 3654 3397 3688
rect 3435 3654 3452 3688
rect 3452 3654 3469 3688
rect 3507 3654 3520 3688
rect 3520 3654 3541 3688
rect 3938 3666 3972 3692
rect 3938 3658 3972 3666
rect -32344 3568 -32315 3602
rect -32315 3568 -32310 3602
rect -32266 3568 -32232 3602
rect -32188 3568 -32154 3602
rect -32110 3568 -32076 3602
rect -32032 3568 -31998 3602
rect -31954 3568 -31920 3602
rect -31876 3568 -31842 3602
rect -31798 3568 -31764 3602
rect -31718 3579 -31684 3613
rect -31645 3612 -31632 3613
rect -31632 3612 -31611 3613
rect -31572 3612 -31563 3613
rect -31563 3612 -31538 3613
rect -31499 3612 -31494 3613
rect -31494 3612 -31465 3613
rect -31426 3612 -31425 3613
rect -31425 3612 -31392 3613
rect -31353 3612 -31322 3613
rect -31322 3612 -31319 3613
rect -31280 3612 -31253 3613
rect -31253 3612 -31246 3613
rect -31207 3612 -31184 3613
rect -31184 3612 -31173 3613
rect -31134 3612 -31115 3613
rect -31115 3612 -31100 3613
rect -31061 3612 -31046 3613
rect -31046 3612 -31027 3613
rect -30988 3612 -30977 3613
rect -30977 3612 -30954 3613
rect -30915 3612 -30908 3613
rect -30908 3612 -30881 3613
rect -30842 3612 -30839 3613
rect -30839 3612 -30808 3613
rect -30768 3612 -30735 3613
rect -30735 3612 -30734 3613
rect -30694 3612 -30666 3613
rect -30666 3612 -30660 3613
rect -30620 3612 -30597 3613
rect -30597 3612 -30586 3613
rect -30546 3612 -30528 3613
rect -30528 3612 -30512 3613
rect -30472 3612 -30459 3613
rect -30459 3612 -30438 3613
rect -30398 3612 -30390 3613
rect -30390 3612 -30364 3613
rect -30324 3612 -30321 3613
rect -30321 3612 -30290 3613
rect -30250 3612 -30218 3613
rect -30218 3612 -30216 3613
rect -30176 3612 -30149 3613
rect -30149 3612 -30142 3613
rect -30102 3612 -30080 3613
rect -30080 3612 -30068 3613
rect -30028 3612 -30011 3613
rect -30011 3612 -29994 3613
rect -29954 3612 -29942 3613
rect -29942 3612 -29920 3613
rect -29880 3612 -29873 3613
rect -29873 3612 -29846 3613
rect -29806 3612 -29804 3613
rect -29804 3612 -29772 3613
rect -29732 3612 -29700 3613
rect -29700 3612 -29698 3613
rect -29658 3612 -29631 3613
rect -29631 3612 -29624 3613
rect -29584 3612 -29562 3613
rect -29562 3612 -29550 3613
rect -29510 3612 -29493 3613
rect -29493 3612 -29476 3613
rect -29436 3612 -29424 3613
rect -29424 3612 -29402 3613
rect -29362 3612 -29355 3613
rect -29355 3612 -29328 3613
rect -29288 3612 -29286 3613
rect -29286 3612 -29254 3613
rect -29134 3642 -29114 3646
rect -29114 3642 -29100 3646
rect -29046 3642 -29044 3654
rect -29044 3642 -29012 3654
rect -29214 3612 -29183 3613
rect -29183 3612 -29180 3613
rect -28958 3642 -28942 3654
rect -28942 3642 -28924 3654
rect -28870 3642 -28840 3654
rect -28840 3642 -28836 3654
rect -28189 3621 -28160 3654
rect -28160 3621 -28155 3654
rect -28115 3621 -28092 3654
rect -28092 3621 -28081 3654
rect -28041 3621 -28024 3654
rect -28024 3621 -28007 3654
rect -27967 3621 -27956 3654
rect -27956 3621 -27933 3654
rect -27893 3621 -27888 3654
rect -27888 3621 -27859 3654
rect -27819 3621 -27786 3654
rect -27786 3621 -27785 3654
rect -27745 3621 -27718 3654
rect -27718 3621 -27711 3654
rect -27671 3621 -27650 3654
rect -27650 3621 -27637 3654
rect -27597 3621 -27582 3654
rect -27582 3621 -27563 3654
rect -27523 3621 -27514 3654
rect -27514 3621 -27489 3654
rect -27449 3621 -27446 3654
rect -27446 3621 -27415 3654
rect -27375 3621 -27344 3654
rect -27344 3621 -27341 3654
rect -27301 3621 -27276 3654
rect -27276 3621 -27267 3654
rect -27227 3621 -27208 3654
rect -27208 3621 -27193 3654
rect -27153 3621 -27140 3654
rect -27140 3621 -27119 3654
rect -31645 3579 -31611 3612
rect -31572 3579 -31538 3612
rect -31499 3579 -31465 3612
rect -31426 3579 -31392 3612
rect -31353 3579 -31319 3612
rect -31280 3579 -31246 3612
rect -31207 3579 -31173 3612
rect -31134 3579 -31100 3612
rect -31061 3579 -31027 3612
rect -30988 3579 -30954 3612
rect -30915 3579 -30881 3612
rect -30842 3579 -30808 3612
rect -30768 3579 -30734 3612
rect -30694 3579 -30660 3612
rect -30620 3579 -30586 3612
rect -30546 3579 -30512 3612
rect -30472 3579 -30438 3612
rect -30398 3579 -30364 3612
rect -30324 3579 -30290 3612
rect -30250 3579 -30216 3612
rect -30176 3579 -30142 3612
rect -30102 3579 -30068 3612
rect -30028 3579 -29994 3612
rect -29954 3579 -29920 3612
rect -29880 3579 -29846 3612
rect -29806 3579 -29772 3612
rect -29732 3579 -29698 3612
rect -29658 3579 -29624 3612
rect -29584 3579 -29550 3612
rect -29510 3579 -29476 3612
rect -29436 3579 -29402 3612
rect -29362 3579 -29328 3612
rect -29288 3579 -29254 3612
rect -29214 3579 -29180 3612
rect -29134 3576 -29100 3603
rect -29046 3585 -29012 3603
rect -28958 3585 -28924 3603
rect -28870 3585 -28836 3603
rect -29134 3569 -29114 3576
rect -29114 3569 -29100 3576
rect -29046 3569 -29044 3585
rect -29044 3569 -29012 3585
rect -28958 3569 -28942 3585
rect -28942 3569 -28924 3585
rect -28870 3569 -28840 3585
rect -28840 3569 -28836 3585
rect -28189 3551 -28160 3582
rect -28160 3551 -28155 3582
rect -28115 3551 -28092 3582
rect -28092 3551 -28081 3582
rect -28041 3551 -28024 3582
rect -28024 3551 -28007 3582
rect -27967 3551 -27956 3582
rect -27956 3551 -27933 3582
rect -27893 3551 -27888 3582
rect -27888 3551 -27859 3582
rect -27819 3551 -27786 3582
rect -27786 3551 -27785 3582
rect -27745 3551 -27718 3582
rect -27718 3551 -27711 3582
rect -27671 3551 -27650 3582
rect -27650 3551 -27637 3582
rect -27597 3551 -27582 3582
rect -27582 3551 -27563 3582
rect -27523 3551 -27514 3582
rect -27514 3551 -27489 3582
rect -27449 3551 -27446 3582
rect -27446 3551 -27415 3582
rect -27375 3551 -27344 3582
rect -27344 3551 -27341 3582
rect -27301 3551 -27276 3582
rect -27276 3551 -27267 3582
rect -27227 3551 -27208 3582
rect -27208 3551 -27193 3582
rect -27153 3551 -27140 3582
rect -27140 3551 -27119 3582
rect 4718 3738 4723 3753
rect 4723 3738 4752 3753
rect 4802 3738 4815 3753
rect 4815 3738 4836 3753
rect 4886 3738 4907 3753
rect 4907 3738 4920 3753
rect 4718 3719 4752 3738
rect 4802 3719 4836 3738
rect 4886 3719 4920 3738
rect 4718 3669 4723 3678
rect 4723 3669 4752 3678
rect 4802 3669 4815 3678
rect 4815 3669 4836 3678
rect 4886 3669 4907 3678
rect 4907 3669 4920 3678
rect 3938 3598 3972 3616
rect 3938 3582 3972 3598
rect -28189 3548 -28155 3551
rect -28115 3548 -28081 3551
rect -28041 3548 -28007 3551
rect -27967 3548 -27933 3551
rect -27893 3548 -27859 3551
rect -27819 3548 -27785 3551
rect -27745 3548 -27711 3551
rect -27671 3548 -27637 3551
rect -27597 3548 -27563 3551
rect -27523 3548 -27489 3551
rect -27449 3548 -27415 3551
rect -27375 3548 -27341 3551
rect -27301 3548 -27267 3551
rect -27227 3548 -27193 3551
rect -27153 3548 -27119 3551
rect -32344 3495 -32315 3529
rect -32315 3495 -32310 3529
rect -32266 3495 -32232 3529
rect -32188 3495 -32154 3529
rect -32110 3495 -32076 3529
rect -32032 3495 -31998 3529
rect -31954 3495 -31920 3529
rect -31876 3495 -31842 3529
rect -31798 3495 -31764 3529
rect -31718 3507 -31684 3541
rect -31645 3507 -31611 3541
rect -31572 3507 -31538 3541
rect -31499 3507 -31465 3541
rect -31426 3507 -31392 3541
rect -31353 3507 -31319 3541
rect -31280 3507 -31246 3541
rect -31207 3507 -31173 3541
rect -31134 3507 -31100 3541
rect -31061 3507 -31027 3541
rect -30988 3507 -30954 3541
rect -30915 3507 -30881 3541
rect -30842 3507 -30808 3541
rect -30768 3507 -30734 3541
rect -30694 3507 -30660 3541
rect -30620 3507 -30586 3541
rect -30546 3507 -30512 3541
rect -30472 3507 -30438 3541
rect -30398 3507 -30364 3541
rect -30324 3507 -30290 3541
rect -30250 3507 -30216 3541
rect -30176 3507 -30142 3541
rect -30102 3507 -30068 3541
rect -30028 3507 -29994 3541
rect -29954 3507 -29920 3541
rect -29880 3507 -29846 3541
rect -29806 3507 -29772 3541
rect -29732 3507 -29698 3541
rect -29658 3507 -29624 3541
rect -29584 3507 -29550 3541
rect -29510 3507 -29476 3541
rect -29436 3507 -29402 3541
rect -29362 3507 -29328 3541
rect -29288 3507 -29254 3541
rect -29214 3507 -29180 3541
rect -29134 3506 -29100 3530
rect -29046 3516 -29012 3530
rect -28958 3516 -28924 3530
rect -28870 3516 -28836 3530
rect -29134 3496 -29114 3506
rect -29114 3496 -29100 3506
rect -29046 3496 -29044 3516
rect -29044 3496 -29012 3516
rect -28958 3496 -28942 3516
rect -28942 3496 -28924 3516
rect -28870 3496 -28840 3516
rect -28840 3496 -28836 3516
rect -28189 3482 -28160 3509
rect -28160 3482 -28155 3509
rect -28115 3482 -28092 3509
rect -28092 3482 -28081 3509
rect -28041 3482 -28024 3509
rect -28024 3482 -28007 3509
rect -27967 3482 -27956 3509
rect -27956 3482 -27933 3509
rect -27893 3482 -27888 3509
rect -27888 3482 -27859 3509
rect -27819 3482 -27786 3509
rect -27786 3482 -27785 3509
rect -27745 3482 -27718 3509
rect -27718 3482 -27711 3509
rect -27671 3482 -27650 3509
rect -27650 3482 -27637 3509
rect -27597 3482 -27582 3509
rect -27582 3482 -27563 3509
rect -27523 3482 -27514 3509
rect -27514 3482 -27489 3509
rect -27449 3482 -27446 3509
rect -27446 3482 -27415 3509
rect -27375 3482 -27344 3509
rect -27344 3482 -27341 3509
rect -27301 3482 -27276 3509
rect -27276 3482 -27267 3509
rect -27227 3482 -27208 3509
rect -27208 3482 -27193 3509
rect -27153 3482 -27140 3509
rect -27140 3482 -27119 3509
rect -28189 3475 -28155 3482
rect -28115 3475 -28081 3482
rect -28041 3475 -28007 3482
rect -27967 3475 -27933 3482
rect -27893 3475 -27859 3482
rect -27819 3475 -27785 3482
rect -27745 3475 -27711 3482
rect -27671 3475 -27637 3482
rect -27597 3475 -27563 3482
rect -27523 3475 -27489 3482
rect -27449 3475 -27415 3482
rect -27375 3475 -27341 3482
rect -27301 3475 -27267 3482
rect -27227 3475 -27193 3482
rect -27153 3475 -27119 3482
rect -32344 3422 -32315 3456
rect -32315 3422 -32310 3456
rect -32266 3422 -32232 3456
rect -32188 3422 -32154 3456
rect -32110 3422 -32076 3456
rect -32032 3422 -31998 3456
rect -31954 3422 -31920 3456
rect -31876 3422 -31842 3456
rect -31798 3422 -31764 3456
rect -31718 3435 -31684 3469
rect -31645 3436 -31611 3469
rect -31572 3436 -31538 3469
rect -31499 3436 -31465 3469
rect -31426 3436 -31392 3469
rect -31353 3436 -31319 3469
rect -31280 3436 -31246 3469
rect -31207 3436 -31173 3469
rect -31134 3436 -31100 3469
rect -31061 3436 -31027 3469
rect -30988 3436 -30954 3469
rect -30915 3436 -30881 3469
rect -30842 3436 -30808 3469
rect -30768 3436 -30734 3469
rect -30694 3436 -30660 3469
rect -30620 3436 -30586 3469
rect -30546 3436 -30512 3469
rect -30472 3436 -30438 3469
rect -30398 3436 -30364 3469
rect -30324 3436 -30290 3469
rect -30250 3436 -30216 3469
rect -30176 3436 -30142 3469
rect -30102 3436 -30068 3469
rect -30028 3436 -29994 3469
rect -29954 3436 -29920 3469
rect -29880 3436 -29846 3469
rect -29806 3436 -29772 3469
rect -29732 3436 -29698 3469
rect -29658 3436 -29624 3469
rect -29584 3436 -29550 3469
rect -29510 3436 -29476 3469
rect -29436 3436 -29402 3469
rect -29362 3436 -29328 3469
rect -29288 3436 -29254 3469
rect -29214 3436 -29180 3469
rect -29134 3436 -29100 3457
rect -29046 3447 -29012 3457
rect -28958 3447 -28924 3457
rect -28870 3447 -28836 3457
rect -31645 3435 -31632 3436
rect -31632 3435 -31611 3436
rect -31572 3435 -31563 3436
rect -31563 3435 -31538 3436
rect -31499 3435 -31494 3436
rect -31494 3435 -31465 3436
rect -31426 3435 -31425 3436
rect -31425 3435 -31392 3436
rect -31353 3435 -31322 3436
rect -31322 3435 -31319 3436
rect -31280 3435 -31253 3436
rect -31253 3435 -31246 3436
rect -31207 3435 -31184 3436
rect -31184 3435 -31173 3436
rect -31134 3435 -31115 3436
rect -31115 3435 -31100 3436
rect -31061 3435 -31046 3436
rect -31046 3435 -31027 3436
rect -30988 3435 -30977 3436
rect -30977 3435 -30954 3436
rect -30915 3435 -30908 3436
rect -30908 3435 -30881 3436
rect -30842 3435 -30839 3436
rect -30839 3435 -30808 3436
rect -30768 3435 -30735 3436
rect -30735 3435 -30734 3436
rect -30694 3435 -30666 3436
rect -30666 3435 -30660 3436
rect -30620 3435 -30597 3436
rect -30597 3435 -30586 3436
rect -30546 3435 -30528 3436
rect -30528 3435 -30512 3436
rect -30472 3435 -30459 3436
rect -30459 3435 -30438 3436
rect -30398 3435 -30390 3436
rect -30390 3435 -30364 3436
rect -30324 3435 -30321 3436
rect -30321 3435 -30290 3436
rect -30250 3435 -30218 3436
rect -30218 3435 -30216 3436
rect -30176 3435 -30149 3436
rect -30149 3435 -30142 3436
rect -30102 3435 -30080 3436
rect -30080 3435 -30068 3436
rect -30028 3435 -30011 3436
rect -30011 3435 -29994 3436
rect -29954 3435 -29942 3436
rect -29942 3435 -29920 3436
rect -29880 3435 -29873 3436
rect -29873 3435 -29846 3436
rect -29806 3435 -29804 3436
rect -29804 3435 -29772 3436
rect -29732 3435 -29700 3436
rect -29700 3435 -29698 3436
rect -29658 3435 -29631 3436
rect -29631 3435 -29624 3436
rect -29584 3435 -29562 3436
rect -29562 3435 -29550 3436
rect -29510 3435 -29493 3436
rect -29493 3435 -29476 3436
rect -29436 3435 -29424 3436
rect -29424 3435 -29402 3436
rect -29362 3435 -29355 3436
rect -29355 3435 -29328 3436
rect -29288 3435 -29286 3436
rect -29286 3435 -29254 3436
rect -29214 3435 -29183 3436
rect -29183 3435 -29180 3436
rect -29134 3423 -29114 3436
rect -29114 3423 -29100 3436
rect -29046 3423 -29044 3447
rect -29044 3423 -29012 3447
rect -28958 3423 -28942 3447
rect -28942 3423 -28924 3447
rect -28870 3423 -28840 3447
rect -28840 3423 -28836 3447
rect -28189 3413 -28160 3436
rect -28160 3413 -28155 3436
rect -28115 3413 -28092 3436
rect -28092 3413 -28081 3436
rect -28041 3413 -28024 3436
rect -28024 3413 -28007 3436
rect -27967 3413 -27956 3436
rect -27956 3413 -27933 3436
rect -27893 3413 -27888 3436
rect -27888 3413 -27859 3436
rect -27819 3413 -27786 3436
rect -27786 3413 -27785 3436
rect -27745 3413 -27718 3436
rect -27718 3413 -27711 3436
rect -27671 3413 -27650 3436
rect -27650 3413 -27637 3436
rect -27597 3413 -27582 3436
rect -27582 3413 -27563 3436
rect -27523 3413 -27514 3436
rect -27514 3413 -27489 3436
rect -27449 3413 -27446 3436
rect -27446 3413 -27415 3436
rect -27375 3413 -27344 3436
rect -27344 3413 -27341 3436
rect -27301 3413 -27276 3436
rect -27276 3413 -27267 3436
rect -27227 3413 -27208 3436
rect -27208 3413 -27193 3436
rect -27153 3413 -27140 3436
rect -27140 3413 -27119 3436
rect -28189 3402 -28155 3413
rect -28115 3402 -28081 3413
rect -28041 3402 -28007 3413
rect -27967 3402 -27933 3413
rect -27893 3402 -27859 3413
rect -27819 3402 -27785 3413
rect -27745 3402 -27711 3413
rect -27671 3402 -27637 3413
rect -27597 3402 -27563 3413
rect -27523 3402 -27489 3413
rect -27449 3402 -27415 3413
rect -27375 3402 -27341 3413
rect -27301 3402 -27267 3413
rect -27227 3402 -27193 3413
rect -27153 3402 -27119 3413
rect -32344 3349 -32315 3383
rect -32315 3349 -32310 3383
rect -32266 3349 -32232 3383
rect -32188 3349 -32154 3383
rect -32110 3349 -32076 3383
rect -32032 3349 -31998 3383
rect -31954 3349 -31920 3383
rect -31876 3349 -31842 3383
rect -31798 3349 -31764 3383
rect -31718 3363 -31684 3397
rect -31645 3363 -31611 3397
rect -31572 3363 -31538 3397
rect -31499 3363 -31465 3397
rect -31426 3363 -31392 3397
rect -31353 3363 -31319 3397
rect -31280 3363 -31246 3397
rect -31207 3363 -31173 3397
rect -31134 3363 -31100 3397
rect -31061 3363 -31027 3397
rect -30988 3363 -30954 3397
rect -30915 3363 -30881 3397
rect -30842 3363 -30808 3397
rect -30768 3363 -30734 3397
rect -30694 3363 -30660 3397
rect -30620 3363 -30586 3397
rect -30546 3363 -30512 3397
rect -30472 3363 -30438 3397
rect -30398 3363 -30364 3397
rect -30324 3363 -30290 3397
rect -30250 3363 -30216 3397
rect -30176 3363 -30142 3397
rect -30102 3363 -30068 3397
rect -30028 3363 -29994 3397
rect -29954 3363 -29920 3397
rect -29880 3363 -29846 3397
rect -29806 3363 -29772 3397
rect -29732 3363 -29698 3397
rect -29658 3363 -29624 3397
rect -29584 3363 -29550 3397
rect -29510 3363 -29476 3397
rect -29436 3363 -29402 3397
rect -29362 3363 -29328 3397
rect -29288 3363 -29254 3397
rect -29214 3363 -29180 3397
rect -29134 3350 -29100 3384
rect -29046 3378 -29012 3384
rect -28958 3378 -28924 3384
rect -28870 3378 -28836 3384
rect -29046 3350 -29044 3378
rect -29044 3350 -29012 3378
rect -28958 3350 -28942 3378
rect -28942 3350 -28924 3378
rect -28870 3350 -28840 3378
rect -28840 3350 -28836 3378
rect -28189 3344 -28160 3363
rect -28160 3344 -28155 3363
rect -28115 3344 -28092 3363
rect -28092 3344 -28081 3363
rect -28041 3344 -28024 3363
rect -28024 3344 -28007 3363
rect -27967 3344 -27956 3363
rect -27956 3344 -27933 3363
rect -27893 3344 -27888 3363
rect -27888 3344 -27859 3363
rect -27819 3344 -27786 3363
rect -27786 3344 -27785 3363
rect -27745 3344 -27718 3363
rect -27718 3344 -27711 3363
rect -27671 3344 -27650 3363
rect -27650 3344 -27637 3363
rect -27597 3344 -27582 3363
rect -27582 3344 -27563 3363
rect -27523 3344 -27514 3363
rect -27514 3344 -27489 3363
rect -27449 3344 -27446 3363
rect -27446 3344 -27415 3363
rect -27375 3344 -27344 3363
rect -27344 3344 -27341 3363
rect -27301 3344 -27276 3363
rect -27276 3344 -27267 3363
rect -27227 3344 -27208 3363
rect -27208 3344 -27193 3363
rect -27153 3344 -27140 3363
rect -27140 3344 -27119 3363
rect -32344 3276 -32315 3310
rect -32315 3276 -32310 3310
rect -32266 3276 -32232 3310
rect -32188 3276 -32154 3310
rect -32110 3276 -32076 3310
rect -32032 3276 -31998 3310
rect -31954 3276 -31920 3310
rect -31876 3276 -31842 3310
rect -31798 3276 -31764 3310
rect -28189 3329 -28155 3344
rect -28115 3329 -28081 3344
rect -28041 3329 -28007 3344
rect -27967 3329 -27933 3344
rect -27893 3329 -27859 3344
rect -27819 3329 -27785 3344
rect -27745 3329 -27711 3344
rect -27671 3329 -27637 3344
rect -27597 3329 -27563 3344
rect -27523 3329 -27489 3344
rect -27449 3329 -27415 3344
rect -27375 3329 -27341 3344
rect -27301 3329 -27267 3344
rect -27227 3329 -27193 3344
rect -27153 3329 -27119 3344
rect -32344 3203 -32315 3237
rect -32315 3203 -32310 3237
rect -32266 3203 -32232 3237
rect -32188 3203 -32154 3237
rect -32110 3203 -32076 3237
rect -32032 3203 -31998 3237
rect -31954 3203 -31920 3237
rect -31876 3203 -31842 3237
rect -31798 3203 -31764 3237
rect -32344 3130 -32315 3164
rect -32315 3130 -32310 3164
rect -32266 3130 -32232 3164
rect -32188 3130 -32154 3164
rect -32110 3130 -32076 3164
rect -32032 3130 -31998 3164
rect -31954 3130 -31920 3164
rect -31876 3130 -31842 3164
rect -31798 3130 -31764 3164
rect -32344 3057 -32315 3091
rect -32315 3057 -32310 3091
rect -32266 3057 -32232 3091
rect -32188 3057 -32154 3091
rect -32110 3057 -32076 3091
rect -32032 3057 -31998 3091
rect -31954 3057 -31920 3091
rect -31876 3057 -31842 3091
rect -31798 3057 -31764 3091
rect -32344 2984 -32315 3018
rect -32315 2984 -32310 3018
rect -32266 2984 -32232 3018
rect -32188 2984 -32154 3018
rect -32110 2984 -32076 3018
rect -32032 2984 -31998 3018
rect -31954 2984 -31920 3018
rect -31876 2984 -31842 3018
rect -31798 2984 -31764 3018
rect -32344 2911 -32315 2945
rect -32315 2911 -32310 2945
rect -32266 2911 -32232 2945
rect -32188 2911 -32154 2945
rect -32110 2911 -32076 2945
rect -32032 2911 -31998 2945
rect -31954 2911 -31920 2945
rect -31876 2911 -31842 2945
rect -31798 2911 -31764 2945
rect -32344 2838 -32315 2872
rect -32315 2838 -32310 2872
rect -32266 2838 -32232 2872
rect -32188 2838 -32154 2872
rect -32110 2838 -32076 2872
rect -32032 2838 -31998 2872
rect -31954 2838 -31920 2872
rect -31876 2838 -31842 2872
rect -31798 2838 -31764 2872
rect -32344 2765 -32315 2799
rect -32315 2765 -32310 2799
rect -32266 2765 -32232 2799
rect -32188 2765 -32154 2799
rect -32110 2765 -32076 2799
rect -32032 2765 -31998 2799
rect -31954 2765 -31920 2799
rect -31876 2765 -31842 2799
rect -31798 2765 -31764 2799
rect -32344 2692 -32315 2726
rect -32315 2692 -32310 2726
rect -32266 2692 -32232 2726
rect -32188 2692 -32154 2726
rect -32110 2692 -32076 2726
rect -32032 2692 -31998 2726
rect -31954 2692 -31920 2726
rect -31876 2692 -31842 2726
rect -31798 2692 -31764 2726
rect -32344 2619 -32315 2653
rect -32315 2619 -32310 2653
rect -32266 2619 -32232 2653
rect -32188 2619 -32154 2653
rect -32110 2619 -32076 2653
rect -32032 2619 -31998 2653
rect -31954 2619 -31920 2653
rect -31876 2619 -31842 2653
rect -31798 2619 -31764 2653
rect -32344 2546 -32315 2580
rect -32315 2546 -32310 2580
rect -32266 2546 -32232 2580
rect -32188 2546 -32154 2580
rect -32110 2546 -32076 2580
rect -32032 2546 -31998 2580
rect -31954 2546 -31920 2580
rect -31876 2546 -31842 2580
rect -31798 2546 -31764 2580
rect -32344 2473 -32315 2507
rect -32315 2473 -32310 2507
rect -32266 2473 -32232 2507
rect -32188 2473 -32154 2507
rect -32110 2473 -32076 2507
rect -32032 2473 -31998 2507
rect -31954 2473 -31920 2507
rect -31876 2473 -31842 2507
rect -31798 2473 -31764 2507
rect -32344 2400 -32315 2434
rect -32315 2400 -32310 2434
rect -32266 2400 -32232 2434
rect -32188 2400 -32154 2434
rect -32110 2400 -32076 2434
rect -32032 2400 -31998 2434
rect -31954 2400 -31920 2434
rect -31876 2400 -31842 2434
rect -31798 2400 -31764 2434
rect -32344 2327 -32315 2361
rect -32315 2327 -32310 2361
rect -32266 2327 -32232 2361
rect -32188 2327 -32154 2361
rect -32110 2327 -32076 2361
rect -32032 2327 -31998 2361
rect -31954 2327 -31920 2361
rect -31876 2327 -31842 2361
rect -31798 2327 -31764 2361
rect -32344 2254 -32315 2288
rect -32315 2254 -32310 2288
rect -32266 2254 -32232 2288
rect -32188 2254 -32154 2288
rect -32110 2254 -32076 2288
rect -32032 2254 -31998 2288
rect -31954 2254 -31920 2288
rect -31876 2254 -31842 2288
rect -31798 2254 -31764 2288
rect -32344 2181 -32315 2215
rect -32315 2181 -32310 2215
rect -32266 2181 -32232 2215
rect -32188 2181 -32154 2215
rect -32110 2181 -32076 2215
rect -32032 2181 -31998 2215
rect -31954 2181 -31920 2215
rect -31876 2181 -31842 2215
rect -31798 2181 -31764 2215
rect -32344 2108 -32315 2142
rect -32315 2108 -32310 2142
rect -32266 2108 -32232 2142
rect -32188 2108 -32154 2142
rect -32110 2108 -32076 2142
rect -32032 2108 -31998 2142
rect -31954 2108 -31920 2142
rect -31876 2108 -31842 2142
rect -31798 2108 -31764 2142
rect -32344 2035 -32315 2069
rect -32315 2035 -32310 2069
rect -32266 2035 -32232 2069
rect -32188 2035 -32154 2069
rect -32110 2035 -32076 2069
rect -32032 2035 -31998 2069
rect -31954 2035 -31920 2069
rect -31876 2035 -31842 2069
rect -31798 2035 -31764 2069
rect -32344 1962 -32315 1996
rect -32315 1962 -32310 1996
rect -32266 1962 -32232 1996
rect -32188 1962 -32154 1996
rect -32110 1962 -32076 1996
rect -32032 1962 -31998 1996
rect -31954 1962 -31920 1996
rect -31876 1962 -31842 1996
rect -31798 1962 -31764 1996
rect -32344 1889 -32315 1923
rect -32315 1889 -32310 1923
rect -32266 1889 -32232 1923
rect -32188 1889 -32154 1923
rect -32110 1889 -32076 1923
rect -32032 1889 -31998 1923
rect -31954 1889 -31920 1923
rect -31876 1889 -31842 1923
rect -31798 1889 -31764 1923
rect -32344 1816 -32315 1850
rect -32315 1816 -32310 1850
rect -32266 1816 -32232 1850
rect -32188 1816 -32154 1850
rect -32110 1816 -32076 1850
rect -32032 1816 -31998 1850
rect -31954 1816 -31920 1850
rect -31876 1816 -31842 1850
rect -31798 1816 -31764 1850
rect -32344 1743 -32315 1777
rect -32315 1743 -32310 1777
rect -32266 1743 -32232 1777
rect -32188 1743 -32154 1777
rect -32110 1743 -32076 1777
rect -32032 1743 -31998 1777
rect -31954 1743 -31920 1777
rect -31876 1743 -31842 1777
rect -31798 1743 -31764 1777
rect -32344 1670 -32315 1704
rect -32315 1670 -32310 1704
rect -32266 1670 -32232 1704
rect -32188 1670 -32154 1704
rect -32110 1670 -32076 1704
rect -32032 1670 -31998 1704
rect -31954 1670 -31920 1704
rect -31876 1670 -31842 1704
rect -31798 1670 -31764 1704
rect -32344 1597 -32315 1631
rect -32315 1597 -32310 1631
rect -32266 1597 -32232 1631
rect -32188 1597 -32154 1631
rect -32110 1597 -32076 1631
rect -32032 1597 -31998 1631
rect -31954 1597 -31920 1631
rect -31876 1597 -31842 1631
rect -31798 1597 -31764 1631
rect -32344 1524 -32315 1558
rect -32315 1524 -32310 1558
rect -32266 1524 -32232 1558
rect -32188 1524 -32154 1558
rect -32110 1524 -32076 1558
rect -32032 1524 -31998 1558
rect -31954 1524 -31920 1558
rect -31876 1524 -31842 1558
rect -31798 1524 -31764 1558
rect -32344 1451 -32315 1485
rect -32315 1451 -32310 1485
rect -32266 1451 -32232 1485
rect -32188 1451 -32154 1485
rect -32110 1451 -32076 1485
rect -32032 1451 -31998 1485
rect -31954 1451 -31920 1485
rect -31876 1451 -31842 1485
rect -31798 1451 -31764 1485
rect -32344 1378 -32315 1412
rect -32315 1378 -32310 1412
rect -32266 1378 -32232 1412
rect -32188 1378 -32154 1412
rect -32110 1378 -32076 1412
rect -32032 1378 -31998 1412
rect -31954 1378 -31920 1412
rect -31876 1378 -31842 1412
rect -31798 1378 -31764 1412
rect -32344 1305 -32315 1339
rect -32315 1305 -32310 1339
rect -32266 1305 -32232 1339
rect -32188 1305 -32154 1339
rect -32110 1305 -32076 1339
rect -32032 1305 -31998 1339
rect -31954 1305 -31920 1339
rect -31876 1305 -31842 1339
rect -31798 1305 -31764 1339
rect -32344 1232 -32315 1266
rect -32315 1232 -32310 1266
rect -32266 1232 -32232 1266
rect -32188 1232 -32154 1266
rect -32110 1232 -32076 1266
rect -32032 1232 -31998 1266
rect -31954 1232 -31920 1266
rect -31876 1232 -31842 1266
rect -31798 1232 -31764 1266
rect -32344 1159 -32315 1193
rect -32315 1159 -32310 1193
rect -32266 1159 -32232 1193
rect -32188 1159 -32154 1193
rect -32110 1159 -32076 1193
rect -32032 1159 -31998 1193
rect -31954 1159 -31920 1193
rect -31876 1159 -31842 1193
rect -31798 1159 -31764 1193
rect -32344 1086 -32315 1120
rect -32315 1086 -32310 1120
rect -32266 1086 -32232 1120
rect -32188 1086 -32154 1120
rect -32110 1086 -32076 1120
rect -32032 1086 -31998 1120
rect -31954 1086 -31920 1120
rect -31876 1086 -31842 1120
rect -31798 1086 -31764 1120
rect -32344 1013 -32315 1047
rect -32315 1013 -32310 1047
rect -32266 1013 -32232 1047
rect -32188 1013 -32154 1047
rect -32110 1013 -32076 1047
rect -32032 1013 -31998 1047
rect -31954 1013 -31920 1047
rect -31876 1013 -31842 1047
rect -31798 1013 -31764 1047
rect -32344 940 -32315 974
rect -32315 940 -32310 974
rect -32266 940 -32232 974
rect -32188 940 -32154 974
rect -32110 940 -32076 974
rect -32032 940 -31998 974
rect -31954 940 -31920 974
rect -31876 940 -31842 974
rect -31798 940 -31764 974
rect -32344 867 -32315 901
rect -32315 867 -32310 901
rect -32266 867 -32232 901
rect -32188 867 -32154 901
rect -32110 867 -32076 901
rect -32032 867 -31998 901
rect -31954 867 -31920 901
rect -31876 867 -31842 901
rect -31798 867 -31764 901
rect -32344 794 -32315 828
rect -32315 794 -32310 828
rect -32266 794 -32232 828
rect -32188 794 -32154 828
rect -32110 794 -32076 828
rect -32032 794 -31998 828
rect -31954 794 -31920 828
rect -31876 794 -31842 828
rect -31798 794 -31764 828
rect -32344 721 -32315 755
rect -32315 721 -32310 755
rect -32266 721 -32232 755
rect -32188 721 -32154 755
rect -32110 721 -32076 755
rect -32032 721 -31998 755
rect -31954 721 -31920 755
rect -31876 721 -31842 755
rect -31798 721 -31764 755
rect -32344 648 -32315 682
rect -32315 648 -32310 682
rect -32266 648 -32232 682
rect -32188 648 -32154 682
rect -32110 648 -32076 682
rect -32032 648 -31998 682
rect -31954 648 -31920 682
rect -31876 648 -31842 682
rect -31798 648 -31764 682
rect -32344 576 -32315 610
rect -32315 576 -32310 610
rect -32266 576 -32232 610
rect -32188 576 -32154 610
rect -32110 576 -32076 610
rect -32032 576 -31998 610
rect -31954 576 -31920 610
rect -31876 576 -31842 610
rect -31798 576 -31764 610
rect -32344 504 -32315 538
rect -32315 504 -32310 538
rect -32266 504 -32232 538
rect -32188 504 -32154 538
rect -32110 504 -32076 538
rect -32032 504 -31998 538
rect -31954 504 -31920 538
rect -31876 504 -31842 538
rect -31798 504 -31764 538
rect -32344 432 -32315 466
rect -32315 432 -32310 466
rect -32266 432 -32232 466
rect -32188 432 -32154 466
rect -32110 432 -32076 466
rect -32032 432 -31998 466
rect -31954 432 -31920 466
rect -31876 432 -31842 466
rect -31798 432 -31764 466
rect -32344 360 -32315 394
rect -32315 360 -32310 394
rect -32266 360 -32232 394
rect -32188 360 -32154 394
rect -32110 360 -32076 394
rect -32032 360 -31998 394
rect -31954 360 -31920 394
rect -31876 360 -31842 394
rect -31798 360 -31764 394
rect -32344 288 -32315 322
rect -32315 288 -32310 322
rect -32266 288 -32232 322
rect -32188 288 -32154 322
rect -32110 288 -32076 322
rect -32032 288 -31998 322
rect -31954 288 -31920 322
rect -31876 288 -31842 322
rect -31798 288 -31764 322
rect -32344 216 -32315 250
rect -32315 216 -32310 250
rect -32266 216 -32232 250
rect -32188 216 -32154 250
rect -32110 216 -32076 250
rect -32032 216 -31998 250
rect -31954 216 -31920 250
rect -31876 216 -31842 250
rect -31798 216 -31764 250
rect -32344 144 -32315 178
rect -32315 144 -32310 178
rect -32266 144 -32232 178
rect -32188 144 -32154 178
rect -32110 144 -32076 178
rect -32032 144 -31998 178
rect -31954 144 -31920 178
rect -31876 144 -31842 178
rect -31798 144 -31764 178
rect -32344 72 -32315 106
rect -32315 72 -32310 106
rect -32266 72 -32232 106
rect -32188 72 -32154 106
rect -32110 72 -32076 106
rect -32032 72 -31998 106
rect -31954 72 -31920 106
rect -31876 72 -31842 106
rect -31798 72 -31764 106
rect -32344 0 -32315 34
rect -32315 0 -32310 34
rect -32266 0 -32232 34
rect -32188 0 -32154 34
rect -32110 0 -32076 34
rect -32032 0 -31998 34
rect -31954 0 -31920 34
rect -31876 0 -31842 34
rect -31798 0 -31764 34
rect -32344 -72 -32315 -38
rect -32315 -72 -32310 -38
rect -32266 -72 -32232 -38
rect -32188 -72 -32154 -38
rect -32110 -72 -32076 -38
rect -32032 -72 -31998 -38
rect -31954 -72 -31920 -38
rect -31876 -72 -31842 -38
rect -31798 -72 -31764 -38
rect -32344 -144 -32315 -110
rect -32315 -144 -32310 -110
rect -32266 -144 -32232 -110
rect -32188 -144 -32154 -110
rect -32110 -144 -32076 -110
rect -32032 -144 -31998 -110
rect -31954 -144 -31920 -110
rect -31876 -144 -31842 -110
rect -31798 -144 -31764 -110
rect -32344 -216 -32315 -182
rect -32315 -216 -32310 -182
rect -32266 -216 -32232 -182
rect -32188 -216 -32154 -182
rect -32110 -216 -32076 -182
rect -32032 -216 -31998 -182
rect -31954 -216 -31920 -182
rect -31876 -216 -31842 -182
rect -31798 -216 -31764 -182
rect -32344 -288 -32315 -254
rect -32315 -288 -32310 -254
rect -32266 -288 -32232 -254
rect -32188 -288 -32154 -254
rect -32110 -288 -32076 -254
rect -32032 -288 -31998 -254
rect -31954 -288 -31920 -254
rect -31876 -288 -31842 -254
rect -31798 -288 -31764 -254
rect -32344 -360 -32315 -326
rect -32315 -360 -32310 -326
rect -32266 -360 -32232 -326
rect -32188 -360 -32154 -326
rect -32110 -360 -32076 -326
rect -32032 -360 -31998 -326
rect -31954 -360 -31920 -326
rect -31876 -360 -31842 -326
rect -31798 -360 -31764 -326
rect -32344 -432 -32315 -398
rect -32315 -432 -32310 -398
rect -32266 -432 -32232 -398
rect -32188 -432 -32154 -398
rect -32110 -432 -32076 -398
rect -32032 -432 -31998 -398
rect -31954 -432 -31920 -398
rect -31876 -432 -31842 -398
rect -31798 -432 -31764 -398
rect -32344 -504 -32315 -470
rect -32315 -504 -32310 -470
rect -32266 -504 -32232 -470
rect -32188 -504 -32154 -470
rect -32110 -504 -32076 -470
rect -32032 -504 -31998 -470
rect -31954 -504 -31920 -470
rect -31876 -504 -31842 -470
rect -31798 -504 -31764 -470
rect -32344 -576 -32315 -542
rect -32315 -576 -32310 -542
rect -32266 -576 -32232 -542
rect -32188 -576 -32154 -542
rect -32110 -576 -32076 -542
rect -32032 -576 -31998 -542
rect -31954 -576 -31920 -542
rect -31876 -576 -31842 -542
rect -31798 -576 -31764 -542
rect -32344 -648 -32315 -614
rect -32315 -648 -32310 -614
rect -32266 -648 -32232 -614
rect -32188 -648 -32154 -614
rect -32110 -648 -32076 -614
rect -32032 -648 -31998 -614
rect -31954 -648 -31920 -614
rect -31876 -648 -31842 -614
rect -31798 -648 -31764 -614
rect -32344 -720 -32315 -686
rect -32315 -720 -32310 -686
rect -32266 -720 -32232 -686
rect -32188 -720 -32154 -686
rect -32110 -720 -32076 -686
rect -32032 -720 -31998 -686
rect -31954 -720 -31920 -686
rect -31876 -720 -31842 -686
rect -31798 -720 -31764 -686
rect -32344 -792 -32315 -758
rect -32315 -792 -32310 -758
rect -32266 -792 -32232 -758
rect -32188 -792 -32154 -758
rect -32110 -792 -32076 -758
rect -32032 -792 -31998 -758
rect -31954 -792 -31920 -758
rect -31876 -792 -31842 -758
rect -31798 -792 -31764 -758
rect -32344 -864 -32315 -830
rect -32315 -864 -32310 -830
rect -32266 -864 -32232 -830
rect -32188 -864 -32154 -830
rect -32110 -864 -32076 -830
rect -32032 -864 -31998 -830
rect -31954 -864 -31920 -830
rect -31876 -864 -31842 -830
rect -31798 -864 -31764 -830
rect -32344 -936 -32315 -902
rect -32315 -936 -32310 -902
rect -32266 -936 -32232 -902
rect -32188 -936 -32154 -902
rect -32110 -936 -32076 -902
rect -32032 -936 -31998 -902
rect -31954 -936 -31920 -902
rect -31876 -936 -31842 -902
rect -31798 -936 -31764 -902
rect -32344 -1008 -32315 -974
rect -32315 -1008 -32310 -974
rect -32266 -1008 -32232 -974
rect -32188 -1008 -32154 -974
rect -32110 -1008 -32076 -974
rect -32032 -1008 -31998 -974
rect -31954 -1008 -31920 -974
rect -31876 -1008 -31842 -974
rect -31798 -1008 -31764 -974
rect -32344 -1080 -32315 -1046
rect -32315 -1080 -32310 -1046
rect -32266 -1080 -32232 -1046
rect -32188 -1080 -32154 -1046
rect -32110 -1080 -32076 -1046
rect -32032 -1080 -31998 -1046
rect -31954 -1080 -31920 -1046
rect -31876 -1080 -31842 -1046
rect -31798 -1080 -31764 -1046
rect -32344 -1152 -32315 -1118
rect -32315 -1152 -32310 -1118
rect -32266 -1152 -32232 -1118
rect -32188 -1152 -32154 -1118
rect -32110 -1152 -32076 -1118
rect -32032 -1152 -31998 -1118
rect -31954 -1152 -31920 -1118
rect -31876 -1152 -31842 -1118
rect -31798 -1152 -31764 -1118
rect -32344 -1224 -32315 -1190
rect -32315 -1224 -32310 -1190
rect -32266 -1224 -32232 -1190
rect -32188 -1224 -32154 -1190
rect -32110 -1224 -32076 -1190
rect -32032 -1224 -31998 -1190
rect -31954 -1224 -31920 -1190
rect -31876 -1224 -31842 -1190
rect -31798 -1224 -31764 -1190
rect -32344 -1296 -32315 -1262
rect -32315 -1296 -32310 -1262
rect -32266 -1296 -32232 -1262
rect -32188 -1296 -32154 -1262
rect -32110 -1296 -32076 -1262
rect -32032 -1296 -31998 -1262
rect -31954 -1296 -31920 -1262
rect -31876 -1296 -31842 -1262
rect -31798 -1296 -31764 -1262
rect -32344 -1368 -32315 -1334
rect -32315 -1368 -32310 -1334
rect -32266 -1368 -32232 -1334
rect -32188 -1368 -32154 -1334
rect -32110 -1368 -32076 -1334
rect -32032 -1368 -31998 -1334
rect -31954 -1368 -31920 -1334
rect -31876 -1368 -31842 -1334
rect -31798 -1368 -31764 -1334
rect -32344 -1440 -32315 -1406
rect -32315 -1440 -32310 -1406
rect -32266 -1440 -32232 -1406
rect -32188 -1440 -32154 -1406
rect -32110 -1440 -32076 -1406
rect -32032 -1440 -31998 -1406
rect -31954 -1440 -31920 -1406
rect -31876 -1440 -31842 -1406
rect -31798 -1440 -31764 -1406
rect -32344 -1512 -32315 -1478
rect -32315 -1512 -32310 -1478
rect -32266 -1512 -32232 -1478
rect -32188 -1512 -32154 -1478
rect -32110 -1512 -32076 -1478
rect -32032 -1512 -31998 -1478
rect -31954 -1512 -31920 -1478
rect -31876 -1512 -31842 -1478
rect -31798 -1512 -31764 -1478
rect -32344 -1584 -32315 -1550
rect -32315 -1584 -32310 -1550
rect -32266 -1584 -32232 -1550
rect -32188 -1584 -32154 -1550
rect -32110 -1584 -32076 -1550
rect -32032 -1584 -31998 -1550
rect -31954 -1584 -31920 -1550
rect -31876 -1584 -31842 -1550
rect -31798 -1584 -31764 -1550
rect -32344 -1656 -32315 -1622
rect -32315 -1656 -32310 -1622
rect -32266 -1656 -32232 -1622
rect -32188 -1656 -32154 -1622
rect -32110 -1656 -32076 -1622
rect -32032 -1656 -31998 -1622
rect -31954 -1656 -31920 -1622
rect -31876 -1656 -31842 -1622
rect -31798 -1656 -31764 -1622
rect -32344 -1728 -32315 -1694
rect -32315 -1728 -32310 -1694
rect -32266 -1728 -32232 -1694
rect -32188 -1728 -32154 -1694
rect -32110 -1728 -32076 -1694
rect -32032 -1728 -31998 -1694
rect -31954 -1728 -31920 -1694
rect -31876 -1728 -31842 -1694
rect -31798 -1728 -31764 -1694
rect -32344 -1800 -32315 -1766
rect -32315 -1800 -32310 -1766
rect -32266 -1800 -32232 -1766
rect -32188 -1800 -32154 -1766
rect -32110 -1800 -32076 -1766
rect -32032 -1800 -31998 -1766
rect -31954 -1800 -31920 -1766
rect -31876 -1800 -31842 -1766
rect -31798 -1800 -31764 -1766
rect -32344 -1872 -32315 -1838
rect -32315 -1872 -32310 -1838
rect -32266 -1872 -32232 -1838
rect -32188 -1872 -32154 -1838
rect -32110 -1872 -32076 -1838
rect -32032 -1872 -31998 -1838
rect -31954 -1872 -31920 -1838
rect -31876 -1872 -31842 -1838
rect -31798 -1872 -31764 -1838
rect -32344 -1944 -32315 -1910
rect -32315 -1944 -32310 -1910
rect -32266 -1944 -32232 -1910
rect -32188 -1944 -32154 -1910
rect -32110 -1944 -32076 -1910
rect -32032 -1944 -31998 -1910
rect -31954 -1944 -31920 -1910
rect -31876 -1944 -31842 -1910
rect -31798 -1944 -31764 -1910
rect -32344 -2016 -32315 -1982
rect -32315 -2016 -32310 -1982
rect -32266 -2016 -32232 -1982
rect -32188 -2016 -32154 -1982
rect -32110 -2016 -32076 -1982
rect -32032 -2016 -31998 -1982
rect -31954 -2016 -31920 -1982
rect -31876 -2016 -31842 -1982
rect -31798 -2016 -31764 -1982
rect -32344 -2088 -32315 -2054
rect -32315 -2088 -32310 -2054
rect -32266 -2088 -32232 -2054
rect -32188 -2088 -32154 -2054
rect -32110 -2088 -32076 -2054
rect -32032 -2088 -31998 -2054
rect -31954 -2088 -31920 -2054
rect -31876 -2088 -31842 -2054
rect -31798 -2088 -31764 -2054
rect -32344 -2160 -32315 -2126
rect -32315 -2160 -32310 -2126
rect -32266 -2160 -32232 -2126
rect -32188 -2160 -32154 -2126
rect -32110 -2160 -32076 -2126
rect -32032 -2160 -31998 -2126
rect -31954 -2160 -31920 -2126
rect -31876 -2160 -31842 -2126
rect -31798 -2160 -31764 -2126
rect -32344 -2232 -32315 -2198
rect -32315 -2232 -32310 -2198
rect -32266 -2232 -32232 -2198
rect -32188 -2232 -32154 -2198
rect -32110 -2232 -32076 -2198
rect -32032 -2232 -31998 -2198
rect -31954 -2232 -31920 -2198
rect -31876 -2232 -31842 -2198
rect -31798 -2232 -31764 -2198
rect -32344 -2304 -32315 -2270
rect -32315 -2304 -32310 -2270
rect -32266 -2304 -32232 -2270
rect -32188 -2304 -32154 -2270
rect -32110 -2304 -32076 -2270
rect -32032 -2304 -31998 -2270
rect -31954 -2304 -31920 -2270
rect -31876 -2304 -31842 -2270
rect -31798 -2304 -31764 -2270
rect -32344 -2376 -32315 -2342
rect -32315 -2376 -32310 -2342
rect -32266 -2376 -32232 -2342
rect -32188 -2376 -32154 -2342
rect -32110 -2376 -32076 -2342
rect -32032 -2376 -31998 -2342
rect -31954 -2376 -31920 -2342
rect -31876 -2376 -31842 -2342
rect -31798 -2376 -31764 -2342
rect -32344 -2448 -32315 -2414
rect -32315 -2448 -32310 -2414
rect -32266 -2448 -32232 -2414
rect -32188 -2448 -32154 -2414
rect -32110 -2448 -32076 -2414
rect -32032 -2448 -31998 -2414
rect -31954 -2448 -31920 -2414
rect -31876 -2448 -31842 -2414
rect -31798 -2448 -31764 -2414
rect -32344 -2520 -32315 -2486
rect -32315 -2520 -32310 -2486
rect -32266 -2520 -32232 -2486
rect -32188 -2520 -32154 -2486
rect -32110 -2520 -32076 -2486
rect -32032 -2520 -31998 -2486
rect -31954 -2520 -31920 -2486
rect -31876 -2520 -31842 -2486
rect -31798 -2520 -31764 -2486
rect -32344 -2592 -32315 -2558
rect -32315 -2592 -32310 -2558
rect -32266 -2592 -32232 -2558
rect -32188 -2592 -32154 -2558
rect -32110 -2592 -32076 -2558
rect -32032 -2592 -31998 -2558
rect -31954 -2592 -31920 -2558
rect -31876 -2592 -31842 -2558
rect -31798 -2592 -31764 -2558
rect -32344 -2664 -32315 -2630
rect -32315 -2664 -32310 -2630
rect -32266 -2664 -32232 -2630
rect -32188 -2664 -32154 -2630
rect -32110 -2664 -32076 -2630
rect -32032 -2664 -31998 -2630
rect -31954 -2664 -31920 -2630
rect -31876 -2664 -31842 -2630
rect -31798 -2664 -31764 -2630
rect -32344 -2736 -32315 -2702
rect -32315 -2736 -32310 -2702
rect -32266 -2736 -32232 -2702
rect -32188 -2736 -32154 -2702
rect -32110 -2736 -32076 -2702
rect -32032 -2736 -31998 -2702
rect -31954 -2736 -31920 -2702
rect -31876 -2736 -31842 -2702
rect -31798 -2736 -31764 -2702
rect -32344 -2808 -32315 -2774
rect -32315 -2808 -32310 -2774
rect -32266 -2808 -32232 -2774
rect -32188 -2808 -32154 -2774
rect -32110 -2808 -32076 -2774
rect -32032 -2808 -31998 -2774
rect -31954 -2808 -31920 -2774
rect -31876 -2808 -31842 -2774
rect -31798 -2808 -31764 -2774
rect -32344 -2880 -32315 -2846
rect -32315 -2880 -32310 -2846
rect -32266 -2880 -32232 -2846
rect -32188 -2880 -32154 -2846
rect -32110 -2880 -32076 -2846
rect -32032 -2880 -31998 -2846
rect -31954 -2880 -31920 -2846
rect -31876 -2880 -31842 -2846
rect -31798 -2880 -31764 -2846
rect -32344 -2952 -32315 -2918
rect -32315 -2952 -32310 -2918
rect -32266 -2952 -32232 -2918
rect -32188 -2952 -32154 -2918
rect -32110 -2952 -32076 -2918
rect -32032 -2952 -31998 -2918
rect -31954 -2952 -31920 -2918
rect -31876 -2952 -31842 -2918
rect -31798 -2952 -31764 -2918
rect -32344 -3024 -32315 -2990
rect -32315 -3024 -32310 -2990
rect -32266 -3024 -32232 -2990
rect -32188 -3024 -32154 -2990
rect -32110 -3024 -32076 -2990
rect -32032 -3024 -31998 -2990
rect -31954 -3024 -31920 -2990
rect -31876 -3024 -31842 -2990
rect -31798 -3024 -31764 -2990
rect -32344 -3096 -32315 -3062
rect -32315 -3096 -32310 -3062
rect -32266 -3096 -32232 -3062
rect -32188 -3096 -32154 -3062
rect -32110 -3096 -32076 -3062
rect -32032 -3096 -31998 -3062
rect -31954 -3096 -31920 -3062
rect -31876 -3096 -31842 -3062
rect -31798 -3096 -31764 -3062
rect -32344 -3168 -32315 -3134
rect -32315 -3168 -32310 -3134
rect -32266 -3168 -32232 -3134
rect -32188 -3168 -32154 -3134
rect -32110 -3168 -32076 -3134
rect -32032 -3168 -31998 -3134
rect -31954 -3168 -31920 -3134
rect -31876 -3168 -31842 -3134
rect -31798 -3168 -31764 -3134
rect -32344 -3240 -32315 -3206
rect -32315 -3240 -32310 -3206
rect -32266 -3240 -32232 -3206
rect -32188 -3240 -32154 -3206
rect -32110 -3240 -32076 -3206
rect -32032 -3240 -31998 -3206
rect -31954 -3240 -31920 -3206
rect -31876 -3240 -31842 -3206
rect -31798 -3240 -31764 -3206
rect -32344 -3312 -32315 -3278
rect -32315 -3312 -32310 -3278
rect -32266 -3312 -32232 -3278
rect -32188 -3312 -32154 -3278
rect -32110 -3312 -32076 -3278
rect -32032 -3312 -31998 -3278
rect -31954 -3312 -31920 -3278
rect -31876 -3312 -31842 -3278
rect -31798 -3312 -31764 -3278
rect -32344 -3384 -32315 -3350
rect -32315 -3384 -32310 -3350
rect -32266 -3384 -32232 -3350
rect -32188 -3384 -32154 -3350
rect -32110 -3384 -32076 -3350
rect -32032 -3384 -31998 -3350
rect -31954 -3384 -31920 -3350
rect -31876 -3384 -31842 -3350
rect -31798 -3384 -31764 -3350
rect -32344 -3456 -32315 -3422
rect -32315 -3456 -32310 -3422
rect -32266 -3456 -32232 -3422
rect -32188 -3456 -32154 -3422
rect -32110 -3456 -32076 -3422
rect -32032 -3456 -31998 -3422
rect -31954 -3456 -31920 -3422
rect -31876 -3456 -31842 -3422
rect -31798 -3456 -31764 -3422
rect -32344 -3528 -32315 -3494
rect -32315 -3528 -32310 -3494
rect -32266 -3528 -32232 -3494
rect -32188 -3528 -32154 -3494
rect -32110 -3528 -32076 -3494
rect -32032 -3528 -31998 -3494
rect -31954 -3528 -31920 -3494
rect -31876 -3528 -31842 -3494
rect -31798 -3528 -31764 -3494
rect -32344 -3600 -32315 -3566
rect -32315 -3600 -32310 -3566
rect -32266 -3600 -32232 -3566
rect -32188 -3600 -32154 -3566
rect -32110 -3600 -32076 -3566
rect -32032 -3600 -31998 -3566
rect -31954 -3600 -31920 -3566
rect -31876 -3600 -31842 -3566
rect -31798 -3600 -31764 -3566
rect -32344 -3672 -32315 -3638
rect -32315 -3672 -32310 -3638
rect -32266 -3672 -32232 -3638
rect -32188 -3672 -32154 -3638
rect -32110 -3672 -32076 -3638
rect -32032 -3672 -31998 -3638
rect -31954 -3672 -31920 -3638
rect -31876 -3672 -31842 -3638
rect -31798 -3672 -31764 -3638
rect -32344 -3744 -32315 -3710
rect -32315 -3744 -32310 -3710
rect -32266 -3744 -32232 -3710
rect -32188 -3744 -32154 -3710
rect -32110 -3744 -32076 -3710
rect -32032 -3744 -31998 -3710
rect -31954 -3744 -31920 -3710
rect -31876 -3744 -31842 -3710
rect -31798 -3744 -31764 -3710
rect -32344 -3816 -32315 -3782
rect -32315 -3816 -32310 -3782
rect -32266 -3816 -32232 -3782
rect -32188 -3816 -32154 -3782
rect -32110 -3816 -32076 -3782
rect -32032 -3816 -31998 -3782
rect -31954 -3816 -31920 -3782
rect -31876 -3816 -31842 -3782
rect -31798 -3816 -31764 -3782
rect -32344 -3888 -32315 -3854
rect -32315 -3888 -32310 -3854
rect -32266 -3888 -32232 -3854
rect -32188 -3888 -32154 -3854
rect -32110 -3888 -32076 -3854
rect -32032 -3888 -31998 -3854
rect -31954 -3888 -31920 -3854
rect -31876 -3888 -31842 -3854
rect -31798 -3888 -31764 -3854
rect -32344 -3960 -32315 -3926
rect -32315 -3960 -32310 -3926
rect -32266 -3960 -32232 -3926
rect -32188 -3960 -32154 -3926
rect -32110 -3960 -32076 -3926
rect -32032 -3960 -31998 -3926
rect -31954 -3960 -31920 -3926
rect -31876 -3960 -31842 -3926
rect -31798 -3960 -31764 -3926
rect -32344 -4032 -32315 -3998
rect -32315 -4032 -32310 -3998
rect -32266 -4032 -32232 -3998
rect -32188 -4032 -32154 -3998
rect -32110 -4032 -32076 -3998
rect -32032 -4032 -31998 -3998
rect -31954 -4032 -31920 -3998
rect -31876 -4032 -31842 -3998
rect -31798 -4032 -31764 -3998
rect -32344 -4104 -32315 -4070
rect -32315 -4104 -32310 -4070
rect -32266 -4104 -32232 -4070
rect -32188 -4104 -32154 -4070
rect -32110 -4104 -32076 -4070
rect -32032 -4104 -31998 -4070
rect -31954 -4104 -31920 -4070
rect -31876 -4104 -31842 -4070
rect -31798 -4104 -31764 -4070
rect -32344 -4176 -32315 -4142
rect -32315 -4176 -32310 -4142
rect -32266 -4176 -32232 -4142
rect -32188 -4176 -32154 -4142
rect -32110 -4176 -32076 -4142
rect -32032 -4176 -31998 -4142
rect -31954 -4176 -31920 -4142
rect -31876 -4176 -31842 -4142
rect -31798 -4176 -31764 -4142
rect -32344 -4248 -32315 -4214
rect -32315 -4248 -32310 -4214
rect -32266 -4248 -32232 -4214
rect -32188 -4248 -32154 -4214
rect -32110 -4248 -32076 -4214
rect -32032 -4248 -31998 -4214
rect -31954 -4248 -31920 -4214
rect -31876 -4248 -31842 -4214
rect -31798 -4248 -31764 -4214
rect -32344 -4320 -32315 -4286
rect -32315 -4320 -32310 -4286
rect -32266 -4320 -32232 -4286
rect -32188 -4320 -32154 -4286
rect -32110 -4320 -32076 -4286
rect -32032 -4320 -31998 -4286
rect -31954 -4320 -31920 -4286
rect -31876 -4320 -31842 -4286
rect -31798 -4320 -31764 -4286
rect -32344 -4392 -32315 -4358
rect -32315 -4392 -32310 -4358
rect -32266 -4392 -32232 -4358
rect -32188 -4392 -32154 -4358
rect -32110 -4392 -32076 -4358
rect -32032 -4392 -31998 -4358
rect -31954 -4392 -31920 -4358
rect -31876 -4392 -31842 -4358
rect -31798 -4392 -31764 -4358
rect -32344 -4464 -32315 -4430
rect -32315 -4464 -32310 -4430
rect -32266 -4464 -32232 -4430
rect -32188 -4464 -32154 -4430
rect -32110 -4464 -32076 -4430
rect -32032 -4464 -31998 -4430
rect -31954 -4464 -31920 -4430
rect -31876 -4464 -31842 -4430
rect -31798 -4464 -31764 -4430
rect -32344 -4536 -32315 -4502
rect -32315 -4536 -32310 -4502
rect -32266 -4536 -32232 -4502
rect -32188 -4536 -32154 -4502
rect -32110 -4536 -32076 -4502
rect -32032 -4536 -31998 -4502
rect -31954 -4536 -31920 -4502
rect -31876 -4536 -31842 -4502
rect -31798 -4536 -31764 -4502
rect -32344 -4608 -32315 -4574
rect -32315 -4608 -32310 -4574
rect -32266 -4608 -32232 -4574
rect -32188 -4608 -32154 -4574
rect -32110 -4608 -32076 -4574
rect -32032 -4608 -31998 -4574
rect -31954 -4608 -31920 -4574
rect -31876 -4608 -31842 -4574
rect -31798 -4608 -31764 -4574
rect -32344 -4680 -32315 -4646
rect -32315 -4680 -32310 -4646
rect -32266 -4680 -32232 -4646
rect -32188 -4680 -32154 -4646
rect -32110 -4680 -32076 -4646
rect -32032 -4680 -31998 -4646
rect -31954 -4680 -31920 -4646
rect -31876 -4680 -31842 -4646
rect -31798 -4680 -31764 -4646
rect -32344 -4752 -32315 -4718
rect -32315 -4752 -32310 -4718
rect -32266 -4752 -32232 -4718
rect -32188 -4752 -32154 -4718
rect -32110 -4752 -32076 -4718
rect -32032 -4752 -31998 -4718
rect -31954 -4752 -31920 -4718
rect -31876 -4752 -31842 -4718
rect -31798 -4752 -31764 -4718
rect -32344 -4824 -32315 -4790
rect -32315 -4824 -32310 -4790
rect -32266 -4824 -32232 -4790
rect -32188 -4824 -32154 -4790
rect -32110 -4824 -32076 -4790
rect -32032 -4824 -31998 -4790
rect -31954 -4824 -31920 -4790
rect -31876 -4824 -31842 -4790
rect -31798 -4824 -31764 -4790
rect -32344 -4896 -32315 -4862
rect -32315 -4896 -32310 -4862
rect -32266 -4896 -32232 -4862
rect -32188 -4896 -32154 -4862
rect -32110 -4896 -32076 -4862
rect -32032 -4896 -31998 -4862
rect -31954 -4896 -31920 -4862
rect -31876 -4896 -31842 -4862
rect -31798 -4896 -31764 -4862
rect -32344 -4968 -32315 -4934
rect -32315 -4968 -32310 -4934
rect -32266 -4968 -32232 -4934
rect -32188 -4968 -32154 -4934
rect -32110 -4968 -32076 -4934
rect -32032 -4968 -31998 -4934
rect -31954 -4968 -31920 -4934
rect -31876 -4968 -31842 -4934
rect -31798 -4968 -31764 -4934
rect -32344 -5040 -32315 -5006
rect -32315 -5040 -32310 -5006
rect -32266 -5040 -32232 -5006
rect -32188 -5040 -32154 -5006
rect -32110 -5040 -32076 -5006
rect -32032 -5040 -31998 -5006
rect -31954 -5040 -31920 -5006
rect -31876 -5040 -31842 -5006
rect -31798 -5040 -31764 -5006
rect -32344 -5112 -32315 -5078
rect -32315 -5112 -32310 -5078
rect -32266 -5112 -32232 -5078
rect -32188 -5112 -32154 -5078
rect -32110 -5112 -32076 -5078
rect -32032 -5112 -31998 -5078
rect -31954 -5112 -31920 -5078
rect -31876 -5112 -31842 -5078
rect -31798 -5112 -31764 -5078
rect -32344 -5184 -32315 -5150
rect -32315 -5184 -32310 -5150
rect -32266 -5184 -32232 -5150
rect -32188 -5184 -32154 -5150
rect -32110 -5184 -32076 -5150
rect -32032 -5184 -31998 -5150
rect -31954 -5184 -31920 -5150
rect -31876 -5184 -31842 -5150
rect -31798 -5184 -31764 -5150
rect -32344 -5256 -32315 -5222
rect -32315 -5256 -32310 -5222
rect -32266 -5256 -32232 -5222
rect -32188 -5256 -32154 -5222
rect -32110 -5256 -32076 -5222
rect -32032 -5256 -31998 -5222
rect -31954 -5256 -31920 -5222
rect -31876 -5256 -31842 -5222
rect -31798 -5256 -31764 -5222
rect -32344 -5328 -32315 -5294
rect -32315 -5328 -32310 -5294
rect -32266 -5328 -32232 -5294
rect -32188 -5328 -32154 -5294
rect -32110 -5328 -32076 -5294
rect -32032 -5328 -31998 -5294
rect -31954 -5328 -31920 -5294
rect -31876 -5328 -31842 -5294
rect -31798 -5328 -31764 -5294
rect -32344 -5400 -32315 -5366
rect -32315 -5400 -32310 -5366
rect -32266 -5400 -32232 -5366
rect -32188 -5400 -32154 -5366
rect -32110 -5400 -32076 -5366
rect -32032 -5400 -31998 -5366
rect -31954 -5400 -31920 -5366
rect -31876 -5400 -31842 -5366
rect -31798 -5400 -31764 -5366
rect -32344 -5472 -32315 -5438
rect -32315 -5472 -32310 -5438
rect -32266 -5472 -32232 -5438
rect -32188 -5472 -32154 -5438
rect -32110 -5472 -32076 -5438
rect -32032 -5472 -31998 -5438
rect -31954 -5472 -31920 -5438
rect -31876 -5472 -31842 -5438
rect -31798 -5472 -31764 -5438
rect -32344 -5544 -32315 -5510
rect -32315 -5544 -32310 -5510
rect -32266 -5544 -32232 -5510
rect -32188 -5544 -32154 -5510
rect -32110 -5544 -32076 -5510
rect -32032 -5544 -31998 -5510
rect -31954 -5544 -31920 -5510
rect -31876 -5544 -31842 -5510
rect -31798 -5544 -31764 -5510
rect -32344 -5616 -32315 -5582
rect -32315 -5616 -32310 -5582
rect -32266 -5616 -32232 -5582
rect -32188 -5616 -32154 -5582
rect -32110 -5616 -32076 -5582
rect -32032 -5616 -31998 -5582
rect -31954 -5616 -31920 -5582
rect -31876 -5616 -31842 -5582
rect -31798 -5616 -31764 -5582
rect -32344 -5688 -32315 -5654
rect -32315 -5688 -32310 -5654
rect -32266 -5688 -32232 -5654
rect -32188 -5688 -32154 -5654
rect -32110 -5688 -32076 -5654
rect -32032 -5688 -31998 -5654
rect -31954 -5688 -31920 -5654
rect -31876 -5688 -31842 -5654
rect -31798 -5688 -31764 -5654
rect -32344 -5760 -32315 -5726
rect -32315 -5760 -32310 -5726
rect -32266 -5760 -32232 -5726
rect -32188 -5760 -32154 -5726
rect -32110 -5760 -32076 -5726
rect -32032 -5760 -31998 -5726
rect -31954 -5760 -31920 -5726
rect -31876 -5760 -31842 -5726
rect -31798 -5760 -31764 -5726
rect -32344 -5832 -32315 -5798
rect -32315 -5832 -32310 -5798
rect -32266 -5832 -32232 -5798
rect -32188 -5832 -32154 -5798
rect -32110 -5832 -32076 -5798
rect -32032 -5832 -31998 -5798
rect -31954 -5832 -31920 -5798
rect -31876 -5832 -31842 -5798
rect -31798 -5832 -31764 -5798
rect -32344 -5904 -32315 -5870
rect -32315 -5904 -32310 -5870
rect -32266 -5904 -32232 -5870
rect -32188 -5904 -32154 -5870
rect -32110 -5904 -32076 -5870
rect -32032 -5904 -31998 -5870
rect -31954 -5904 -31920 -5870
rect -31876 -5904 -31842 -5870
rect -31798 -5904 -31764 -5870
rect -32344 -5976 -32315 -5942
rect -32315 -5976 -32310 -5942
rect -32266 -5976 -32232 -5942
rect -32188 -5976 -32154 -5942
rect -32110 -5976 -32076 -5942
rect -32032 -5976 -31998 -5942
rect -31954 -5976 -31920 -5942
rect -31876 -5976 -31842 -5942
rect -31798 -5976 -31764 -5942
rect -32344 -6048 -32315 -6014
rect -32315 -6048 -32310 -6014
rect -32266 -6048 -32232 -6014
rect -32188 -6048 -32154 -6014
rect -32110 -6048 -32076 -6014
rect -32032 -6048 -31998 -6014
rect -31954 -6048 -31920 -6014
rect -31876 -6048 -31842 -6014
rect -31798 -6048 -31764 -6014
rect -32344 -6120 -32315 -6086
rect -32315 -6120 -32310 -6086
rect -32266 -6120 -32232 -6086
rect -32188 -6120 -32154 -6086
rect -32110 -6120 -32076 -6086
rect -32032 -6120 -31998 -6086
rect -31954 -6120 -31920 -6086
rect -31876 -6120 -31842 -6086
rect -31798 -6120 -31764 -6086
rect -32344 -6192 -32315 -6158
rect -32315 -6192 -32310 -6158
rect -32266 -6192 -32232 -6158
rect -32188 -6192 -32154 -6158
rect -32110 -6192 -32076 -6158
rect -32032 -6192 -31998 -6158
rect -31954 -6192 -31920 -6158
rect -31876 -6192 -31842 -6158
rect -31798 -6192 -31764 -6158
rect -32344 -6264 -32315 -6230
rect -32315 -6264 -32310 -6230
rect -32266 -6264 -32232 -6230
rect -32188 -6264 -32154 -6230
rect -32110 -6264 -32076 -6230
rect -32032 -6264 -31998 -6230
rect -31954 -6264 -31920 -6230
rect -31876 -6264 -31842 -6230
rect -31798 -6264 -31764 -6230
rect -32344 -6336 -32315 -6302
rect -32315 -6336 -32310 -6302
rect -32266 -6336 -32232 -6302
rect -32188 -6336 -32154 -6302
rect -32110 -6336 -32076 -6302
rect -32032 -6336 -31998 -6302
rect -31954 -6336 -31920 -6302
rect -31876 -6336 -31842 -6302
rect -31798 -6336 -31764 -6302
rect -32344 -6408 -32315 -6374
rect -32315 -6408 -32310 -6374
rect -32266 -6408 -32232 -6374
rect -32188 -6408 -32154 -6374
rect -32110 -6408 -32076 -6374
rect -32032 -6408 -31998 -6374
rect -31954 -6408 -31920 -6374
rect -31876 -6408 -31842 -6374
rect -31798 -6408 -31764 -6374
rect -32344 -6480 -32315 -6446
rect -32315 -6480 -32310 -6446
rect -32266 -6480 -32232 -6446
rect -32188 -6480 -32154 -6446
rect -32110 -6480 -32076 -6446
rect -32032 -6480 -31998 -6446
rect -31954 -6480 -31920 -6446
rect -31876 -6480 -31842 -6446
rect -31798 -6480 -31764 -6446
rect -32344 -6552 -32315 -6518
rect -32315 -6552 -32310 -6518
rect -32266 -6552 -32232 -6518
rect -32188 -6552 -32154 -6518
rect -32110 -6552 -32076 -6518
rect -32032 -6552 -31998 -6518
rect -31954 -6552 -31920 -6518
rect -31876 -6552 -31842 -6518
rect -31798 -6552 -31764 -6518
rect -32344 -6624 -32315 -6590
rect -32315 -6624 -32310 -6590
rect -32266 -6624 -32232 -6590
rect -32188 -6624 -32154 -6590
rect -32110 -6624 -32076 -6590
rect -32032 -6624 -31998 -6590
rect -31954 -6624 -31920 -6590
rect -31876 -6624 -31842 -6590
rect -31798 -6624 -31764 -6590
rect -32344 -6696 -32315 -6662
rect -32315 -6696 -32310 -6662
rect -32266 -6696 -32232 -6662
rect -32188 -6696 -32154 -6662
rect -32110 -6696 -32076 -6662
rect -32032 -6696 -31998 -6662
rect -31954 -6696 -31920 -6662
rect -31876 -6696 -31842 -6662
rect -31798 -6696 -31764 -6662
rect -32344 -6768 -32315 -6734
rect -32315 -6768 -32310 -6734
rect -32266 -6768 -32232 -6734
rect -32188 -6768 -32154 -6734
rect -32110 -6768 -32076 -6734
rect -32032 -6768 -31998 -6734
rect -31954 -6768 -31920 -6734
rect -31876 -6768 -31842 -6734
rect -31798 -6768 -31764 -6734
rect -32344 -6840 -32315 -6806
rect -32315 -6840 -32310 -6806
rect -32266 -6840 -32232 -6806
rect -32188 -6840 -32154 -6806
rect -32110 -6840 -32076 -6806
rect -32032 -6840 -31998 -6806
rect -31954 -6840 -31920 -6806
rect -31876 -6840 -31842 -6806
rect -31798 -6840 -31764 -6806
rect -32344 -6912 -32315 -6878
rect -32315 -6912 -32310 -6878
rect -32266 -6912 -32232 -6878
rect -32188 -6912 -32154 -6878
rect -32110 -6912 -32076 -6878
rect -32032 -6912 -31998 -6878
rect -31954 -6912 -31920 -6878
rect -31876 -6912 -31842 -6878
rect -31798 -6912 -31764 -6878
rect -32344 -6984 -32315 -6950
rect -32315 -6984 -32310 -6950
rect -32266 -6984 -32232 -6950
rect -32188 -6984 -32154 -6950
rect -32110 -6984 -32076 -6950
rect -32032 -6984 -31998 -6950
rect -31954 -6984 -31920 -6950
rect -31876 -6984 -31842 -6950
rect -31798 -6984 -31764 -6950
rect -32344 -7056 -32315 -7022
rect -32315 -7056 -32310 -7022
rect -32266 -7056 -32232 -7022
rect -32188 -7056 -32154 -7022
rect -32110 -7056 -32076 -7022
rect -32032 -7056 -31998 -7022
rect -31954 -7056 -31920 -7022
rect -31876 -7056 -31842 -7022
rect -31798 -7056 -31764 -7022
rect -32344 -7128 -32315 -7094
rect -32315 -7128 -32310 -7094
rect -32266 -7128 -32232 -7094
rect -32188 -7128 -32154 -7094
rect -32110 -7128 -32076 -7094
rect -32032 -7128 -31998 -7094
rect -31954 -7128 -31920 -7094
rect -31876 -7128 -31842 -7094
rect -31798 -7128 -31764 -7094
rect -32344 -7200 -32315 -7166
rect -32315 -7200 -32310 -7166
rect -32266 -7200 -32232 -7166
rect -32188 -7200 -32154 -7166
rect -32110 -7200 -32076 -7166
rect -32032 -7200 -31998 -7166
rect -31954 -7200 -31920 -7166
rect -31876 -7200 -31842 -7166
rect -31798 -7200 -31764 -7166
rect -32344 -7272 -32315 -7238
rect -32315 -7272 -32310 -7238
rect -32266 -7272 -32232 -7238
rect -32188 -7272 -32154 -7238
rect -32110 -7272 -32076 -7238
rect -32032 -7272 -31998 -7238
rect -31954 -7272 -31920 -7238
rect -31876 -7272 -31842 -7238
rect -31798 -7272 -31764 -7238
rect -32344 -7344 -32315 -7310
rect -32315 -7344 -32310 -7310
rect -32266 -7344 -32232 -7310
rect -32188 -7344 -32154 -7310
rect -32110 -7344 -32076 -7310
rect -32032 -7344 -31998 -7310
rect -31954 -7344 -31920 -7310
rect -31876 -7344 -31842 -7310
rect -31798 -7344 -31764 -7310
rect -32344 -7416 -32315 -7382
rect -32315 -7416 -32310 -7382
rect -32266 -7416 -32232 -7382
rect -32188 -7416 -32154 -7382
rect -32110 -7416 -32076 -7382
rect -32032 -7416 -31998 -7382
rect -31954 -7416 -31920 -7382
rect -31876 -7416 -31842 -7382
rect -31798 -7416 -31764 -7382
rect -32344 -7488 -32315 -7454
rect -32315 -7488 -32310 -7454
rect -32266 -7488 -32232 -7454
rect -32188 -7488 -32154 -7454
rect -32110 -7488 -32076 -7454
rect -32032 -7488 -31998 -7454
rect -31954 -7488 -31920 -7454
rect -31876 -7488 -31842 -7454
rect -31798 -7488 -31764 -7454
rect -32344 -7560 -32315 -7526
rect -32315 -7560 -32310 -7526
rect -32266 -7560 -32232 -7526
rect -32188 -7560 -32154 -7526
rect -32110 -7560 -32076 -7526
rect -32032 -7560 -31998 -7526
rect -31954 -7560 -31920 -7526
rect -31876 -7560 -31842 -7526
rect -31798 -7560 -31764 -7526
rect -32344 -7632 -32315 -7598
rect -32315 -7632 -32310 -7598
rect -32266 -7632 -32232 -7598
rect -32188 -7632 -32154 -7598
rect -32110 -7632 -32076 -7598
rect -32032 -7632 -31998 -7598
rect -31954 -7632 -31920 -7598
rect -31876 -7632 -31842 -7598
rect -31798 -7632 -31764 -7598
rect -32344 -7704 -32315 -7670
rect -32315 -7704 -32310 -7670
rect -32266 -7704 -32232 -7670
rect -32188 -7704 -32154 -7670
rect -32110 -7704 -32076 -7670
rect -32032 -7704 -31998 -7670
rect -31954 -7704 -31920 -7670
rect -31876 -7704 -31842 -7670
rect -31798 -7704 -31764 -7670
rect -32344 -7776 -32315 -7742
rect -32315 -7776 -32310 -7742
rect -32266 -7776 -32232 -7742
rect -32188 -7776 -32154 -7742
rect -32110 -7776 -32076 -7742
rect -32032 -7776 -31998 -7742
rect -31954 -7776 -31920 -7742
rect -31876 -7776 -31842 -7742
rect -31798 -7776 -31764 -7742
rect -32344 -7848 -32315 -7814
rect -32315 -7848 -32310 -7814
rect -32266 -7848 -32232 -7814
rect -32188 -7848 -32154 -7814
rect -32110 -7848 -32076 -7814
rect -32032 -7848 -31998 -7814
rect -31954 -7848 -31920 -7814
rect -31876 -7848 -31842 -7814
rect -31798 -7848 -31764 -7814
rect -32344 -7920 -32315 -7886
rect -32315 -7920 -32310 -7886
rect -32266 -7920 -32232 -7886
rect -32188 -7920 -32154 -7886
rect -32110 -7920 -32076 -7886
rect -32032 -7920 -31998 -7886
rect -31954 -7920 -31920 -7886
rect -31876 -7920 -31842 -7886
rect -31798 -7920 -31764 -7886
rect -32344 -7992 -32315 -7958
rect -32315 -7992 -32310 -7958
rect -32266 -7992 -32232 -7958
rect -32188 -7992 -32154 -7958
rect -32110 -7992 -32076 -7958
rect -32032 -7992 -31998 -7958
rect -31954 -7992 -31920 -7958
rect -31876 -7992 -31842 -7958
rect -31798 -7992 -31764 -7958
rect -32344 -8064 -32315 -8030
rect -32315 -8064 -32310 -8030
rect -32266 -8064 -32232 -8030
rect -32188 -8064 -32154 -8030
rect -32110 -8064 -32076 -8030
rect -32032 -8064 -31998 -8030
rect -31954 -8064 -31920 -8030
rect -31876 -8064 -31842 -8030
rect -31798 -8064 -31764 -8030
rect -32344 -8136 -32315 -8102
rect -32315 -8136 -32310 -8102
rect -32266 -8136 -32232 -8102
rect -32188 -8136 -32154 -8102
rect -32110 -8136 -32076 -8102
rect -32032 -8136 -31998 -8102
rect -31954 -8136 -31920 -8102
rect -31876 -8136 -31842 -8102
rect -31798 -8136 -31764 -8102
rect -32344 -8208 -32315 -8174
rect -32315 -8208 -32310 -8174
rect -32266 -8208 -32232 -8174
rect -32188 -8208 -32154 -8174
rect -32110 -8208 -32076 -8174
rect -32032 -8208 -31998 -8174
rect -31954 -8208 -31920 -8174
rect -31876 -8208 -31842 -8174
rect -31798 -8208 -31764 -8174
rect -32344 -8280 -32315 -8246
rect -32315 -8280 -32310 -8246
rect -32266 -8280 -32232 -8246
rect -32188 -8280 -32154 -8246
rect -32110 -8280 -32076 -8246
rect -32032 -8280 -31998 -8246
rect -31954 -8280 -31920 -8246
rect -31876 -8280 -31842 -8246
rect -31798 -8280 -31764 -8246
rect -32344 -8352 -32315 -8318
rect -32315 -8352 -32310 -8318
rect -32266 -8352 -32232 -8318
rect -32188 -8352 -32154 -8318
rect -32110 -8352 -32076 -8318
rect -32032 -8352 -31998 -8318
rect -31954 -8352 -31920 -8318
rect -31876 -8352 -31842 -8318
rect -31798 -8352 -31764 -8318
rect -32344 -8424 -32315 -8390
rect -32315 -8424 -32310 -8390
rect -32266 -8424 -32232 -8390
rect -32188 -8424 -32154 -8390
rect -32110 -8424 -32076 -8390
rect -32032 -8424 -31998 -8390
rect -31954 -8424 -31920 -8390
rect -31876 -8424 -31842 -8390
rect -31798 -8424 -31764 -8390
rect -32344 -8496 -32315 -8462
rect -32315 -8496 -32310 -8462
rect -32266 -8496 -32232 -8462
rect -32188 -8496 -32154 -8462
rect -32110 -8496 -32076 -8462
rect -32032 -8496 -31998 -8462
rect -31954 -8496 -31920 -8462
rect -31876 -8496 -31842 -8462
rect -31798 -8496 -31764 -8462
rect -32344 -8568 -32315 -8534
rect -32315 -8568 -32310 -8534
rect -32266 -8568 -32232 -8534
rect -32188 -8568 -32154 -8534
rect -32110 -8568 -32076 -8534
rect -32032 -8568 -31998 -8534
rect -31954 -8568 -31920 -8534
rect -31876 -8568 -31842 -8534
rect -31798 -8568 -31764 -8534
rect -32344 -8640 -32315 -8606
rect -32315 -8640 -32310 -8606
rect -32266 -8640 -32232 -8606
rect -32188 -8640 -32154 -8606
rect -32110 -8640 -32076 -8606
rect -32032 -8640 -31998 -8606
rect -31954 -8640 -31920 -8606
rect -31876 -8640 -31842 -8606
rect -31798 -8640 -31764 -8606
rect -29134 3277 -29100 3311
rect -29046 3309 -29012 3311
rect -28958 3309 -28924 3311
rect -28870 3309 -28836 3311
rect -29046 3277 -29044 3309
rect -29044 3277 -29012 3309
rect -28958 3277 -28942 3309
rect -28942 3277 -28924 3309
rect -28870 3277 -28840 3309
rect -28840 3277 -28836 3309
rect -28189 3275 -28160 3290
rect -28160 3275 -28155 3290
rect -28115 3275 -28092 3290
rect -28092 3275 -28081 3290
rect -28041 3275 -28024 3290
rect -28024 3275 -28007 3290
rect -27967 3275 -27956 3290
rect -27956 3275 -27933 3290
rect -27893 3275 -27888 3290
rect -27888 3275 -27859 3290
rect -27819 3275 -27786 3290
rect -27786 3275 -27785 3290
rect -27745 3275 -27718 3290
rect -27718 3275 -27711 3290
rect -27671 3275 -27650 3290
rect -27650 3275 -27637 3290
rect -27597 3275 -27582 3290
rect -27582 3275 -27563 3290
rect -27523 3275 -27514 3290
rect -27514 3275 -27489 3290
rect -27449 3275 -27446 3290
rect -27446 3275 -27415 3290
rect -27375 3275 -27344 3290
rect -27344 3275 -27341 3290
rect -27301 3275 -27276 3290
rect -27276 3275 -27267 3290
rect -27227 3275 -27208 3290
rect -27208 3275 -27193 3290
rect -27153 3275 -27140 3290
rect -27140 3275 -27119 3290
rect -28189 3256 -28155 3275
rect -28115 3256 -28081 3275
rect -28041 3256 -28007 3275
rect -27967 3256 -27933 3275
rect -27893 3256 -27859 3275
rect -27819 3256 -27785 3275
rect -27745 3256 -27711 3275
rect -27671 3256 -27637 3275
rect -27597 3256 -27563 3275
rect -27523 3256 -27489 3275
rect -27449 3256 -27415 3275
rect -27375 3256 -27341 3275
rect -27301 3256 -27267 3275
rect -27227 3256 -27193 3275
rect -27153 3256 -27119 3275
rect -29134 3232 -29114 3238
rect -29114 3232 -29100 3238
rect -29134 3204 -29100 3232
rect -29046 3206 -29044 3238
rect -29044 3206 -29012 3238
rect -28958 3206 -28942 3238
rect -28942 3206 -28924 3238
rect -28870 3206 -28840 3238
rect -28840 3206 -28836 3238
rect -28189 3206 -28160 3217
rect -28160 3206 -28155 3217
rect -28115 3206 -28092 3217
rect -28092 3206 -28081 3217
rect -28041 3206 -28024 3217
rect -28024 3206 -28007 3217
rect -27967 3206 -27956 3217
rect -27956 3206 -27933 3217
rect -27893 3206 -27888 3217
rect -27888 3206 -27859 3217
rect -27819 3206 -27786 3217
rect -27786 3206 -27785 3217
rect -27745 3206 -27718 3217
rect -27718 3206 -27711 3217
rect -27671 3206 -27650 3217
rect -27650 3206 -27637 3217
rect -27597 3206 -27582 3217
rect -27582 3206 -27563 3217
rect -27523 3206 -27514 3217
rect -27514 3206 -27489 3217
rect -27449 3206 -27446 3217
rect -27446 3206 -27415 3217
rect -27375 3206 -27344 3217
rect -27344 3206 -27341 3217
rect -27301 3206 -27276 3217
rect -27276 3206 -27267 3217
rect -27227 3206 -27208 3217
rect -27208 3206 -27193 3217
rect -27153 3206 -27140 3217
rect -27140 3206 -27119 3217
rect -29046 3204 -29012 3206
rect -28958 3204 -28924 3206
rect -28870 3204 -28836 3206
rect -28189 3183 -28155 3206
rect -28115 3183 -28081 3206
rect -28041 3183 -28007 3206
rect -27967 3183 -27933 3206
rect -27893 3183 -27859 3206
rect -27819 3183 -27785 3206
rect -27745 3183 -27711 3206
rect -27671 3183 -27637 3206
rect -27597 3183 -27563 3206
rect -27523 3183 -27489 3206
rect -27449 3183 -27415 3206
rect -27375 3183 -27341 3206
rect -27301 3183 -27267 3206
rect -27227 3183 -27193 3206
rect -27153 3183 -27119 3206
rect -29134 3164 -29114 3165
rect -29114 3164 -29100 3165
rect -29134 3131 -29100 3164
rect -29046 3137 -29044 3165
rect -29044 3137 -29012 3165
rect -28958 3137 -28942 3165
rect -28942 3137 -28924 3165
rect -28870 3137 -28840 3165
rect -28840 3137 -28836 3165
rect -28189 3137 -28160 3144
rect -28160 3137 -28155 3144
rect -28115 3137 -28092 3144
rect -28092 3137 -28081 3144
rect -28041 3137 -28024 3144
rect -28024 3137 -28007 3144
rect -27967 3137 -27956 3144
rect -27956 3137 -27933 3144
rect -27893 3137 -27888 3144
rect -27888 3137 -27859 3144
rect -27819 3137 -27786 3144
rect -27786 3137 -27785 3144
rect -27745 3137 -27718 3144
rect -27718 3137 -27711 3144
rect -27671 3137 -27650 3144
rect -27650 3137 -27637 3144
rect -27597 3137 -27582 3144
rect -27582 3137 -27563 3144
rect -27523 3137 -27514 3144
rect -27514 3137 -27489 3144
rect -27449 3137 -27446 3144
rect -27446 3137 -27415 3144
rect -27375 3137 -27344 3144
rect -27344 3137 -27341 3144
rect -27301 3137 -27276 3144
rect -27276 3137 -27267 3144
rect -27227 3137 -27208 3144
rect -27208 3137 -27193 3144
rect -27153 3137 -27140 3144
rect -27140 3137 -27119 3144
rect -29046 3131 -29012 3137
rect -28958 3131 -28924 3137
rect -28870 3131 -28836 3137
rect -28189 3110 -28155 3137
rect -28115 3110 -28081 3137
rect -28041 3110 -28007 3137
rect -27967 3110 -27933 3137
rect -27893 3110 -27859 3137
rect -27819 3110 -27785 3137
rect -27745 3110 -27711 3137
rect -27671 3110 -27637 3137
rect -27597 3110 -27563 3137
rect -27523 3110 -27489 3137
rect -27449 3110 -27415 3137
rect -27375 3110 -27341 3137
rect -27301 3110 -27267 3137
rect -27227 3110 -27193 3137
rect -27153 3110 -27119 3137
rect -29134 3062 -29100 3092
rect -29046 3068 -29044 3092
rect -29044 3068 -29012 3092
rect -28958 3068 -28942 3092
rect -28942 3068 -28924 3092
rect -28870 3068 -28840 3092
rect -28840 3068 -28836 3092
rect -28189 3068 -28160 3071
rect -28160 3068 -28155 3071
rect -28115 3068 -28092 3071
rect -28092 3068 -28081 3071
rect -28041 3068 -28024 3071
rect -28024 3068 -28007 3071
rect -27967 3068 -27956 3071
rect -27956 3068 -27933 3071
rect -27893 3068 -27888 3071
rect -27888 3068 -27859 3071
rect -27819 3068 -27786 3071
rect -27786 3068 -27785 3071
rect -27745 3068 -27718 3071
rect -27718 3068 -27711 3071
rect -27671 3068 -27650 3071
rect -27650 3068 -27637 3071
rect -27597 3068 -27582 3071
rect -27582 3068 -27563 3071
rect -27523 3068 -27514 3071
rect -27514 3068 -27489 3071
rect -27449 3068 -27446 3071
rect -27446 3068 -27415 3071
rect -27375 3068 -27344 3071
rect -27344 3068 -27341 3071
rect -27301 3068 -27276 3071
rect -27276 3068 -27267 3071
rect -27227 3068 -27208 3071
rect -27208 3068 -27193 3071
rect -27153 3068 -27140 3071
rect -27140 3068 -27119 3071
rect -29134 3058 -29114 3062
rect -29114 3058 -29100 3062
rect -29046 3058 -29012 3068
rect -28958 3058 -28924 3068
rect -28870 3058 -28836 3068
rect -28189 3037 -28155 3068
rect -28115 3037 -28081 3068
rect -28041 3037 -28007 3068
rect -27967 3037 -27933 3068
rect -27893 3037 -27859 3068
rect -27819 3037 -27785 3068
rect -27745 3037 -27711 3068
rect -27671 3037 -27637 3068
rect -27597 3037 -27563 3068
rect -27523 3037 -27489 3068
rect -27449 3037 -27415 3068
rect -27375 3037 -27341 3068
rect -27301 3037 -27267 3068
rect -27227 3037 -27193 3068
rect -27153 3037 -27119 3068
rect -29134 2994 -29100 3019
rect -29046 2999 -29044 3019
rect -29044 2999 -29012 3019
rect -28958 2999 -28942 3019
rect -28942 2999 -28924 3019
rect -28870 2999 -28840 3019
rect -28840 2999 -28836 3019
rect -29134 2985 -29114 2994
rect -29114 2985 -29100 2994
rect -29046 2985 -29012 2999
rect -28958 2985 -28924 2999
rect -28870 2985 -28836 2999
rect -28189 2964 -28155 2998
rect -28115 2964 -28081 2998
rect -28041 2964 -28007 2998
rect -27967 2964 -27933 2998
rect -27893 2964 -27859 2998
rect -27819 2964 -27785 2998
rect -27745 2964 -27711 2998
rect -27671 2964 -27637 2998
rect -27597 2964 -27563 2998
rect -27523 2964 -27489 2998
rect -27449 2964 -27415 2998
rect -27375 2964 -27341 2998
rect -27301 2964 -27267 2998
rect -27227 2964 -27193 2998
rect -27153 2964 -27119 2998
rect -29134 2926 -29100 2946
rect -29046 2930 -29044 2946
rect -29044 2930 -29012 2946
rect -28958 2930 -28942 2946
rect -28942 2930 -28924 2946
rect -28870 2930 -28840 2946
rect -28840 2930 -28836 2946
rect -29134 2912 -29114 2926
rect -29114 2912 -29100 2926
rect -29046 2912 -29012 2930
rect -28958 2912 -28924 2930
rect -28870 2912 -28836 2930
rect -28189 2895 -28155 2925
rect -28115 2895 -28081 2925
rect -28041 2895 -28007 2925
rect -27967 2895 -27933 2925
rect -27893 2895 -27859 2925
rect -27819 2895 -27785 2925
rect -27745 2895 -27711 2925
rect -27671 2895 -27637 2925
rect -27597 2895 -27563 2925
rect -27523 2895 -27489 2925
rect -27449 2895 -27415 2925
rect -27375 2895 -27341 2925
rect -27301 2895 -27267 2925
rect -27227 2895 -27193 2925
rect -27153 2895 -27119 2925
rect -29134 2858 -29100 2873
rect -29046 2861 -29044 2873
rect -29044 2861 -29012 2873
rect -28958 2861 -28942 2873
rect -28942 2861 -28924 2873
rect -28870 2861 -28840 2873
rect -28840 2861 -28836 2873
rect -28189 2891 -28160 2895
rect -28160 2891 -28155 2895
rect -28115 2891 -28092 2895
rect -28092 2891 -28081 2895
rect -28041 2891 -28024 2895
rect -28024 2891 -28007 2895
rect -27967 2891 -27956 2895
rect -27956 2891 -27933 2895
rect -27893 2891 -27888 2895
rect -27888 2891 -27859 2895
rect -27819 2891 -27786 2895
rect -27786 2891 -27785 2895
rect -27745 2891 -27718 2895
rect -27718 2891 -27711 2895
rect -27671 2891 -27650 2895
rect -27650 2891 -27637 2895
rect -27597 2891 -27582 2895
rect -27582 2891 -27563 2895
rect -27523 2891 -27514 2895
rect -27514 2891 -27489 2895
rect -27449 2891 -27446 2895
rect -27446 2891 -27415 2895
rect -27375 2891 -27344 2895
rect -27344 2891 -27341 2895
rect -27301 2891 -27276 2895
rect -27276 2891 -27267 2895
rect -27227 2891 -27208 2895
rect -27208 2891 -27193 2895
rect -27153 2891 -27140 2895
rect -27140 2891 -27119 2895
rect -29134 2839 -29114 2858
rect -29114 2839 -29100 2858
rect -29046 2839 -29012 2861
rect -28958 2839 -28924 2861
rect -28870 2839 -28836 2861
rect -28189 2826 -28155 2852
rect -28115 2826 -28081 2852
rect -28041 2826 -28007 2852
rect -27967 2826 -27933 2852
rect -27893 2826 -27859 2852
rect -27819 2826 -27785 2852
rect -27745 2826 -27711 2852
rect -27671 2826 -27637 2852
rect -27597 2826 -27563 2852
rect -27523 2826 -27489 2852
rect -27449 2826 -27415 2852
rect -27375 2826 -27341 2852
rect -27301 2826 -27267 2852
rect -27227 2826 -27193 2852
rect -27153 2826 -27119 2852
rect -29134 2790 -29100 2800
rect -29046 2792 -29044 2800
rect -29044 2792 -29012 2800
rect -28958 2792 -28942 2800
rect -28942 2792 -28924 2800
rect -28870 2792 -28840 2800
rect -28840 2792 -28836 2800
rect -28189 2818 -28160 2826
rect -28160 2818 -28155 2826
rect -28115 2818 -28092 2826
rect -28092 2818 -28081 2826
rect -28041 2818 -28024 2826
rect -28024 2818 -28007 2826
rect -27967 2818 -27956 2826
rect -27956 2818 -27933 2826
rect -27893 2818 -27888 2826
rect -27888 2818 -27859 2826
rect -27819 2818 -27786 2826
rect -27786 2818 -27785 2826
rect -27745 2818 -27718 2826
rect -27718 2818 -27711 2826
rect -27671 2818 -27650 2826
rect -27650 2818 -27637 2826
rect -27597 2818 -27582 2826
rect -27582 2818 -27563 2826
rect -27523 2818 -27514 2826
rect -27514 2818 -27489 2826
rect -27449 2818 -27446 2826
rect -27446 2818 -27415 2826
rect -27375 2818 -27344 2826
rect -27344 2818 -27341 2826
rect -27301 2818 -27276 2826
rect -27276 2818 -27267 2826
rect -27227 2818 -27208 2826
rect -27208 2818 -27193 2826
rect -27153 2818 -27140 2826
rect -27140 2818 -27119 2826
rect -29134 2766 -29114 2790
rect -29114 2766 -29100 2790
rect -29046 2766 -29012 2792
rect -28958 2766 -28924 2792
rect -28870 2766 -28836 2792
rect -28189 2757 -28155 2779
rect -28115 2757 -28081 2779
rect -28041 2757 -28007 2779
rect -27967 2757 -27933 2779
rect -27893 2757 -27859 2779
rect -27819 2757 -27785 2779
rect -27745 2757 -27711 2779
rect -27671 2757 -27637 2779
rect -27597 2757 -27563 2779
rect -27523 2757 -27489 2779
rect -27449 2757 -27415 2779
rect -27375 2757 -27341 2779
rect -27301 2757 -27267 2779
rect -27227 2757 -27193 2779
rect -27153 2757 -27119 2779
rect -29134 2722 -29100 2727
rect -29046 2723 -29044 2727
rect -29044 2723 -29012 2727
rect -28958 2723 -28942 2727
rect -28942 2723 -28924 2727
rect -28870 2723 -28840 2727
rect -28840 2723 -28836 2727
rect -28189 2745 -28160 2757
rect -28160 2745 -28155 2757
rect -28115 2745 -28092 2757
rect -28092 2745 -28081 2757
rect -28041 2745 -28024 2757
rect -28024 2745 -28007 2757
rect -27967 2745 -27956 2757
rect -27956 2745 -27933 2757
rect -27893 2745 -27888 2757
rect -27888 2745 -27859 2757
rect -27819 2745 -27786 2757
rect -27786 2745 -27785 2757
rect -27745 2745 -27718 2757
rect -27718 2745 -27711 2757
rect -27671 2745 -27650 2757
rect -27650 2745 -27637 2757
rect -27597 2745 -27582 2757
rect -27582 2745 -27563 2757
rect -27523 2745 -27514 2757
rect -27514 2745 -27489 2757
rect -27449 2745 -27446 2757
rect -27446 2745 -27415 2757
rect -27375 2745 -27344 2757
rect -27344 2745 -27341 2757
rect -27301 2745 -27276 2757
rect -27276 2745 -27267 2757
rect -27227 2745 -27208 2757
rect -27208 2745 -27193 2757
rect -27153 2745 -27140 2757
rect -27140 2745 -27119 2757
rect -29134 2693 -29114 2722
rect -29114 2693 -29100 2722
rect -29046 2693 -29012 2723
rect -28958 2693 -28924 2723
rect -28870 2693 -28836 2723
rect -28189 2688 -28155 2706
rect -28115 2688 -28081 2706
rect -28041 2688 -28007 2706
rect -27967 2688 -27933 2706
rect -27893 2688 -27859 2706
rect -27819 2688 -27785 2706
rect -27745 2688 -27711 2706
rect -27671 2688 -27637 2706
rect -27597 2688 -27563 2706
rect -27523 2688 -27489 2706
rect -27449 2688 -27415 2706
rect -27375 2688 -27341 2706
rect -27301 2688 -27267 2706
rect -27227 2688 -27193 2706
rect -27153 2688 -27119 2706
rect -28189 2672 -28160 2688
rect -28160 2672 -28155 2688
rect -28115 2672 -28092 2688
rect -28092 2672 -28081 2688
rect -28041 2672 -28024 2688
rect -28024 2672 -28007 2688
rect -27967 2672 -27956 2688
rect -27956 2672 -27933 2688
rect -27893 2672 -27888 2688
rect -27888 2672 -27859 2688
rect -27819 2672 -27786 2688
rect -27786 2672 -27785 2688
rect -27745 2672 -27718 2688
rect -27718 2672 -27711 2688
rect -27671 2672 -27650 2688
rect -27650 2672 -27637 2688
rect -27597 2672 -27582 2688
rect -27582 2672 -27563 2688
rect -27523 2672 -27514 2688
rect -27514 2672 -27489 2688
rect -27449 2672 -27446 2688
rect -27446 2672 -27415 2688
rect -27375 2672 -27344 2688
rect -27344 2672 -27341 2688
rect -27301 2672 -27276 2688
rect -27276 2672 -27267 2688
rect -27227 2672 -27208 2688
rect -27208 2672 -27193 2688
rect -27153 2672 -27140 2688
rect -27140 2672 -27119 2688
rect -29134 2620 -29114 2654
rect -29114 2620 -29100 2654
rect -29046 2620 -29012 2654
rect -28958 2620 -28924 2654
rect -28870 2620 -28836 2654
rect -28189 2619 -28155 2633
rect -28115 2619 -28081 2633
rect -28041 2619 -28007 2633
rect -27967 2619 -27933 2633
rect -27893 2619 -27859 2633
rect -27819 2619 -27785 2633
rect -27745 2619 -27711 2633
rect -27671 2619 -27637 2633
rect -27597 2619 -27563 2633
rect -27523 2619 -27489 2633
rect -27449 2619 -27415 2633
rect -27375 2619 -27341 2633
rect -27301 2619 -27267 2633
rect -27227 2619 -27193 2633
rect -27153 2619 -27119 2633
rect -28189 2599 -28160 2619
rect -28160 2599 -28155 2619
rect -28115 2599 -28092 2619
rect -28092 2599 -28081 2619
rect -28041 2599 -28024 2619
rect -28024 2599 -28007 2619
rect -27967 2599 -27956 2619
rect -27956 2599 -27933 2619
rect -27893 2599 -27888 2619
rect -27888 2599 -27859 2619
rect -27819 2599 -27786 2619
rect -27786 2599 -27785 2619
rect -27745 2599 -27718 2619
rect -27718 2599 -27711 2619
rect -27671 2599 -27650 2619
rect -27650 2599 -27637 2619
rect -27597 2599 -27582 2619
rect -27582 2599 -27563 2619
rect -27523 2599 -27514 2619
rect -27514 2599 -27489 2619
rect -27449 2599 -27446 2619
rect -27446 2599 -27415 2619
rect -27375 2599 -27344 2619
rect -27344 2599 -27341 2619
rect -27301 2599 -27276 2619
rect -27276 2599 -27267 2619
rect -27227 2599 -27208 2619
rect -27208 2599 -27193 2619
rect -27153 2599 -27140 2619
rect -27140 2599 -27119 2619
rect -29134 2552 -29114 2581
rect -29114 2552 -29100 2581
rect -29134 2547 -29100 2552
rect -29046 2550 -29012 2581
rect -28958 2550 -28924 2581
rect -28870 2550 -28836 2581
rect -746 3512 -712 3546
rect -746 3442 -712 3474
rect -746 3440 -712 3442
rect -746 3374 -712 3402
rect -746 3368 -712 3374
rect -746 3306 -712 3330
rect -746 3296 -712 3306
rect -746 3238 -712 3258
rect -746 3224 -712 3238
rect -746 3170 -712 3186
rect -746 3152 -712 3170
rect -746 3102 -712 3114
rect -746 3080 -712 3102
rect -746 3034 -712 3042
rect -746 3008 -712 3034
rect -746 2966 -712 2970
rect -746 2936 -712 2966
rect -746 2864 -712 2898
rect -746 2796 -712 2826
rect -746 2792 -712 2796
rect -746 2728 -712 2754
rect -746 2720 -712 2728
rect -746 2660 -712 2682
rect -746 2648 -712 2660
rect -746 2592 -712 2610
rect -746 2576 -712 2592
rect -590 3512 -556 3546
rect -590 3442 -556 3474
rect -590 3440 -556 3442
rect -590 3374 -556 3402
rect -590 3368 -556 3374
rect -590 3306 -556 3330
rect -590 3296 -556 3306
rect -590 3238 -556 3258
rect -590 3224 -556 3238
rect -590 3170 -556 3186
rect -590 3152 -556 3170
rect -590 3102 -556 3114
rect -590 3080 -556 3102
rect -590 3034 -556 3042
rect -590 3008 -556 3034
rect -590 2966 -556 2970
rect -590 2936 -556 2966
rect -590 2864 -556 2898
rect -590 2796 -556 2826
rect -590 2792 -556 2796
rect -590 2728 -556 2754
rect -590 2720 -556 2728
rect -590 2660 -556 2682
rect -590 2648 -556 2660
rect -590 2592 -556 2610
rect -590 2576 -556 2592
rect -434 3512 -400 3546
rect -434 3442 -400 3474
rect -434 3440 -400 3442
rect -434 3374 -400 3402
rect -434 3368 -400 3374
rect -434 3306 -400 3330
rect -434 3296 -400 3306
rect -434 3238 -400 3258
rect -434 3224 -400 3238
rect -434 3170 -400 3186
rect -434 3152 -400 3170
rect -434 3102 -400 3114
rect -434 3080 -400 3102
rect -434 3034 -400 3042
rect -434 3008 -400 3034
rect -434 2966 -400 2970
rect -434 2936 -400 2966
rect -434 2864 -400 2898
rect -434 2796 -400 2826
rect -434 2792 -400 2796
rect -434 2728 -400 2754
rect -434 2720 -400 2728
rect -434 2660 -400 2682
rect -434 2648 -400 2660
rect -434 2592 -400 2610
rect -434 2576 -400 2592
rect 168 3512 202 3546
rect 168 3442 202 3474
rect 168 3440 202 3442
rect 168 3374 202 3402
rect 168 3368 202 3374
rect 168 3306 202 3330
rect 168 3296 202 3306
rect 168 3238 202 3258
rect 168 3224 202 3238
rect 168 3170 202 3186
rect 168 3152 202 3170
rect 168 3102 202 3114
rect 168 3080 202 3102
rect 168 3034 202 3042
rect 168 3008 202 3034
rect 168 2966 202 2970
rect 168 2936 202 2966
rect 168 2864 202 2898
rect 168 2796 202 2826
rect 168 2792 202 2796
rect 168 2728 202 2754
rect 168 2720 202 2728
rect 168 2660 202 2682
rect 168 2648 202 2660
rect 168 2592 202 2610
rect 168 2576 202 2592
rect 324 3512 358 3546
rect 324 3442 358 3474
rect 324 3440 358 3442
rect 324 3374 358 3402
rect 324 3368 358 3374
rect 324 3306 358 3330
rect 324 3296 358 3306
rect 324 3238 358 3258
rect 324 3224 358 3238
rect 324 3170 358 3186
rect 324 3152 358 3170
rect 324 3102 358 3114
rect 324 3080 358 3102
rect 324 3034 358 3042
rect 324 3008 358 3034
rect 324 2966 358 2970
rect 324 2936 358 2966
rect 324 2864 358 2898
rect 324 2796 358 2826
rect 324 2792 358 2796
rect 324 2728 358 2754
rect 324 2720 358 2728
rect 324 2660 358 2682
rect 324 2648 358 2660
rect 324 2592 358 2610
rect 324 2576 358 2592
rect 480 3512 514 3546
rect 480 3442 514 3474
rect 480 3440 514 3442
rect 480 3374 514 3402
rect 480 3368 514 3374
rect 480 3306 514 3330
rect 480 3296 514 3306
rect 480 3238 514 3258
rect 480 3224 514 3238
rect 480 3170 514 3186
rect 480 3152 514 3170
rect 480 3102 514 3114
rect 480 3080 514 3102
rect 480 3034 514 3042
rect 480 3008 514 3034
rect 480 2966 514 2970
rect 480 2936 514 2966
rect 480 2864 514 2898
rect 480 2796 514 2826
rect 480 2792 514 2796
rect 480 2728 514 2754
rect 480 2720 514 2728
rect 480 2660 514 2682
rect 480 2648 514 2660
rect 480 2592 514 2610
rect 480 2576 514 2592
rect 616 3512 650 3546
rect 616 3442 650 3474
rect 616 3440 650 3442
rect 616 3374 650 3402
rect 616 3368 650 3374
rect 616 3306 650 3330
rect 616 3296 650 3306
rect 616 3238 650 3258
rect 616 3224 650 3238
rect 616 3170 650 3186
rect 616 3152 650 3170
rect 616 3102 650 3114
rect 616 3080 650 3102
rect 616 3034 650 3042
rect 616 3008 650 3034
rect 616 2966 650 2970
rect 616 2936 650 2966
rect 616 2864 650 2898
rect 616 2796 650 2826
rect 616 2792 650 2796
rect 616 2728 650 2754
rect 616 2720 650 2728
rect 616 2660 650 2682
rect 616 2648 650 2660
rect 616 2592 650 2610
rect 616 2576 650 2592
rect 772 3512 806 3546
rect 772 3442 806 3474
rect 772 3440 806 3442
rect 772 3374 806 3402
rect 772 3368 806 3374
rect 772 3306 806 3330
rect 772 3296 806 3306
rect 772 3238 806 3258
rect 772 3224 806 3238
rect 772 3170 806 3186
rect 772 3152 806 3170
rect 772 3102 806 3114
rect 772 3080 806 3102
rect 772 3034 806 3042
rect 772 3008 806 3034
rect 772 2966 806 2970
rect 772 2936 806 2966
rect 772 2864 806 2898
rect 772 2796 806 2826
rect 772 2792 806 2796
rect 772 2728 806 2754
rect 772 2720 806 2728
rect 772 2660 806 2682
rect 772 2648 806 2660
rect 772 2592 806 2610
rect 772 2576 806 2592
rect 928 3512 962 3546
rect 928 3442 962 3474
rect 928 3440 962 3442
rect 928 3374 962 3402
rect 928 3368 962 3374
rect 928 3306 962 3330
rect 928 3296 962 3306
rect 928 3238 962 3258
rect 928 3224 962 3238
rect 928 3170 962 3186
rect 928 3152 962 3170
rect 928 3102 962 3114
rect 928 3080 962 3102
rect 928 3034 962 3042
rect 928 3008 962 3034
rect 928 2966 962 2970
rect 928 2936 962 2966
rect 928 2864 962 2898
rect 928 2796 962 2826
rect 928 2792 962 2796
rect 928 2728 962 2754
rect 928 2720 962 2728
rect 928 2660 962 2682
rect 928 2648 962 2660
rect 928 2592 962 2610
rect 928 2576 962 2592
rect 1055 3512 1089 3546
rect 1055 3442 1089 3474
rect 1055 3440 1089 3442
rect 1055 3374 1089 3402
rect 1055 3368 1089 3374
rect 1055 3306 1089 3330
rect 1055 3296 1089 3306
rect 1055 3238 1089 3258
rect 1055 3224 1089 3238
rect 1055 3170 1089 3186
rect 1055 3152 1089 3170
rect 1055 3102 1089 3114
rect 1055 3080 1089 3102
rect 1055 3034 1089 3042
rect 1055 3008 1089 3034
rect 1055 2966 1089 2970
rect 1055 2936 1089 2966
rect 1055 2864 1089 2898
rect 1055 2796 1089 2826
rect 1055 2792 1089 2796
rect 1055 2728 1089 2754
rect 1055 2720 1089 2728
rect 1055 2660 1089 2682
rect 1055 2648 1089 2660
rect 1055 2592 1089 2610
rect 1055 2576 1089 2592
rect 1211 3512 1245 3546
rect 1211 3442 1245 3474
rect 1211 3440 1245 3442
rect 1211 3374 1245 3402
rect 1211 3368 1245 3374
rect 1211 3306 1245 3330
rect 1211 3296 1245 3306
rect 1211 3238 1245 3258
rect 1211 3224 1245 3238
rect 1211 3170 1245 3186
rect 1211 3152 1245 3170
rect 1211 3102 1245 3114
rect 1211 3080 1245 3102
rect 1211 3034 1245 3042
rect 1211 3008 1245 3034
rect 1211 2966 1245 2970
rect 1211 2936 1245 2966
rect 1211 2864 1245 2898
rect 1211 2796 1245 2826
rect 1211 2792 1245 2796
rect 1211 2728 1245 2754
rect 1211 2720 1245 2728
rect 1211 2660 1245 2682
rect 1211 2648 1245 2660
rect 1211 2592 1245 2610
rect 1211 2576 1245 2592
rect 1415 3512 1449 3546
rect 1415 3442 1449 3474
rect 1415 3440 1449 3442
rect 1415 3374 1449 3402
rect 1415 3368 1449 3374
rect 1415 3306 1449 3330
rect 1415 3296 1449 3306
rect 1415 3238 1449 3258
rect 1415 3224 1449 3238
rect 1415 3170 1449 3186
rect 1415 3152 1449 3170
rect 1415 3102 1449 3114
rect 1415 3080 1449 3102
rect 1415 3034 1449 3042
rect 1415 3008 1449 3034
rect 1415 2966 1449 2970
rect 1415 2936 1449 2966
rect 1415 2864 1449 2898
rect 1415 2796 1449 2826
rect 1415 2792 1449 2796
rect 1415 2728 1449 2754
rect 1415 2720 1449 2728
rect 1415 2660 1449 2682
rect 1415 2648 1449 2660
rect 1415 2592 1449 2610
rect 1415 2576 1449 2592
rect 1571 3512 1605 3546
rect 2311 3524 2345 3558
rect 1571 3442 1605 3474
rect 1571 3440 1605 3442
rect 1571 3374 1605 3402
rect 1571 3368 1605 3374
rect 1571 3306 1605 3330
rect 1571 3296 1605 3306
rect 1571 3238 1605 3258
rect 1571 3224 1605 3238
rect 1571 3170 1605 3186
rect 1571 3152 1605 3170
rect 1571 3102 1605 3114
rect 1571 3080 1605 3102
rect 1571 3034 1605 3042
rect 1571 3008 1605 3034
rect 1571 2966 1605 2970
rect 1571 2936 1605 2966
rect 1571 2864 1605 2898
rect 1571 2796 1605 2826
rect 1571 2792 1605 2796
rect 1571 2728 1605 2754
rect 1571 2720 1605 2728
rect 1571 2660 1605 2682
rect 1571 2648 1605 2660
rect 1571 2592 1605 2610
rect 1571 2576 1605 2592
rect 1708 3477 1742 3511
rect 1708 3407 1742 3439
rect 1708 3405 1742 3407
rect 1708 3339 1742 3367
rect 1708 3333 1742 3339
rect 1708 3271 1742 3295
rect 1708 3261 1742 3271
rect 1708 3203 1742 3223
rect 1708 3189 1742 3203
rect 1708 3135 1742 3151
rect 1708 3117 1742 3135
rect 1708 3067 1742 3079
rect 1708 3045 1742 3067
rect 1708 2999 1742 3007
rect 1708 2973 1742 2999
rect 1708 2931 1742 2935
rect 1708 2901 1742 2931
rect 1708 2829 1742 2863
rect 1708 2761 1742 2791
rect 1708 2757 1742 2761
rect 1708 2693 1742 2719
rect 1708 2685 1742 2693
rect 1708 2625 1742 2647
rect 1708 2613 1742 2625
rect -28189 2550 -28155 2560
rect -28115 2550 -28081 2560
rect -28041 2550 -28007 2560
rect -27967 2550 -27933 2560
rect -27893 2550 -27859 2560
rect -27819 2550 -27785 2560
rect -27745 2550 -27711 2560
rect -27671 2550 -27637 2560
rect -27597 2550 -27563 2560
rect -27523 2550 -27489 2560
rect -27449 2550 -27415 2560
rect -27375 2550 -27341 2560
rect -27301 2550 -27267 2560
rect -27227 2550 -27193 2560
rect -27153 2550 -27119 2560
rect -29046 2547 -29044 2550
rect -29044 2547 -29012 2550
rect -28958 2547 -28942 2550
rect -28942 2547 -28924 2550
rect -28870 2547 -28840 2550
rect -28840 2547 -28836 2550
rect -28189 2526 -28160 2550
rect -28160 2526 -28155 2550
rect -28115 2526 -28092 2550
rect -28092 2526 -28081 2550
rect -28041 2526 -28024 2550
rect -28024 2526 -28007 2550
rect -27967 2526 -27956 2550
rect -27956 2526 -27933 2550
rect -27893 2526 -27888 2550
rect -27888 2526 -27859 2550
rect -27819 2526 -27786 2550
rect -27786 2526 -27785 2550
rect -27745 2526 -27718 2550
rect -27718 2526 -27711 2550
rect -27671 2526 -27650 2550
rect -27650 2526 -27637 2550
rect -27597 2526 -27582 2550
rect -27582 2526 -27563 2550
rect -27523 2526 -27514 2550
rect -27514 2526 -27489 2550
rect -27449 2526 -27446 2550
rect -27446 2526 -27415 2550
rect -27375 2526 -27344 2550
rect -27344 2526 -27341 2550
rect -27301 2526 -27276 2550
rect -27276 2526 -27267 2550
rect -27227 2526 -27208 2550
rect -27208 2526 -27193 2550
rect -27153 2526 -27140 2550
rect -27140 2526 -27119 2550
rect 1708 2557 1742 2575
rect 1708 2541 1742 2557
rect 1864 3477 1898 3511
rect 1864 3407 1898 3439
rect 1864 3405 1898 3407
rect 1864 3339 1898 3367
rect 1864 3333 1898 3339
rect 1864 3271 1898 3295
rect 1864 3261 1898 3271
rect 1864 3203 1898 3223
rect 1864 3189 1898 3203
rect 1864 3135 1898 3151
rect 1864 3117 1898 3135
rect 1864 3067 1898 3079
rect 1864 3045 1898 3067
rect 1864 2999 1898 3007
rect 1864 2973 1898 2999
rect 1864 2931 1898 2935
rect 1864 2901 1898 2931
rect 1864 2829 1898 2863
rect 1864 2761 1898 2791
rect 1864 2757 1898 2761
rect 1864 2693 1898 2719
rect 1864 2685 1898 2693
rect 1864 2625 1898 2647
rect 1864 2613 1898 2625
rect 1864 2557 1898 2575
rect 1864 2541 1898 2557
rect 2020 3477 2054 3511
rect 2020 3407 2054 3439
rect 2020 3405 2054 3407
rect 2020 3339 2054 3367
rect 2020 3333 2054 3339
rect 2020 3271 2054 3295
rect 2020 3261 2054 3271
rect 2020 3203 2054 3223
rect 2020 3189 2054 3203
rect 2020 3135 2054 3151
rect 2020 3117 2054 3135
rect 2020 3067 2054 3079
rect 2020 3045 2054 3067
rect 2020 2999 2054 3007
rect 2020 2973 2054 2999
rect 2020 2931 2054 2935
rect 2020 2901 2054 2931
rect 2020 2829 2054 2863
rect 2020 2761 2054 2791
rect 2020 2757 2054 2761
rect 2020 2693 2054 2719
rect 2020 2685 2054 2693
rect 2020 2625 2054 2647
rect 2020 2613 2054 2625
rect 2020 2557 2054 2575
rect 2020 2541 2054 2557
rect 2176 3477 2210 3511
rect 2176 3407 2210 3439
rect 2311 3470 2345 3486
rect 2311 3452 2345 3470
rect 2467 3524 2501 3558
rect 2467 3470 2501 3486
rect 2467 3452 2501 3470
rect 2623 3524 2657 3558
rect 2623 3470 2657 3486
rect 2623 3452 2657 3470
rect 2757 3533 2791 3549
rect 2757 3515 2791 3533
rect 2757 3465 2791 3477
rect 2757 3443 2791 3465
rect 2176 3405 2210 3407
rect 2176 3339 2210 3367
rect 2176 3333 2210 3339
rect 2176 3271 2210 3295
rect 2176 3261 2210 3271
rect 2757 3397 2791 3405
rect 2757 3371 2791 3397
rect 2757 3329 2791 3333
rect 2757 3299 2791 3329
rect 2176 3203 2210 3223
rect 2176 3189 2210 3203
rect 2176 3135 2210 3151
rect 2176 3117 2210 3135
rect 2176 3067 2210 3079
rect 2176 3045 2210 3067
rect 2176 2999 2210 3007
rect 2176 2973 2210 2999
rect 2546 3233 2580 3238
rect 2546 3204 2550 3233
rect 2550 3204 2580 3233
rect 2546 3165 2580 3166
rect 2546 3132 2550 3165
rect 2550 3132 2580 3165
rect 2757 3227 2791 3261
rect 2757 3159 2791 3189
rect 2757 3155 2791 3159
rect 2394 3070 2428 3104
rect 2394 2998 2428 3032
rect 2757 3091 2791 3117
rect 2757 3083 2791 3091
rect 2757 3023 2791 3045
rect 2757 3011 2791 3023
rect 2913 3533 2947 3549
rect 2913 3515 2947 3533
rect 2913 3465 2947 3477
rect 2913 3443 2947 3465
rect 2913 3397 2947 3405
rect 2913 3371 2947 3397
rect 2913 3329 2947 3333
rect 2913 3299 2947 3329
rect 2913 3227 2947 3261
rect 2913 3159 2947 3189
rect 2913 3155 2947 3159
rect 2913 3091 2947 3117
rect 2913 3083 2947 3091
rect 2913 3023 2947 3045
rect 2913 3011 2947 3023
rect 3040 3533 3074 3549
rect 3040 3515 3074 3533
rect 3040 3465 3074 3477
rect 3040 3443 3074 3465
rect 3040 3397 3074 3405
rect 3040 3371 3074 3397
rect 3040 3329 3074 3333
rect 3040 3299 3074 3329
rect 3040 3227 3074 3261
rect 3040 3159 3074 3189
rect 3040 3155 3074 3159
rect 3040 3091 3074 3117
rect 3040 3083 3074 3091
rect 3040 3023 3074 3045
rect 3040 3011 3074 3023
rect 3196 3533 3230 3549
rect 3196 3515 3230 3533
rect 3196 3465 3230 3477
rect 3196 3443 3230 3465
rect 3196 3397 3230 3405
rect 3196 3371 3230 3397
rect 3196 3329 3230 3333
rect 3196 3299 3230 3329
rect 3196 3227 3230 3261
rect 3196 3159 3230 3189
rect 3196 3155 3230 3159
rect 3196 3091 3230 3117
rect 3196 3083 3230 3091
rect 3196 3023 3230 3045
rect 3196 3011 3230 3023
rect 3352 3533 3386 3549
rect 3352 3515 3386 3533
rect 3352 3465 3386 3477
rect 3352 3443 3386 3465
rect 3352 3397 3386 3405
rect 3352 3371 3386 3397
rect 3352 3329 3386 3333
rect 3352 3299 3386 3329
rect 3352 3227 3386 3261
rect 3352 3159 3386 3189
rect 3352 3155 3386 3159
rect 3352 3091 3386 3117
rect 3352 3083 3386 3091
rect 3352 3023 3386 3045
rect 3352 3011 3386 3023
rect 3508 3533 3542 3549
rect 3508 3515 3542 3533
rect 3508 3465 3542 3477
rect 3508 3443 3542 3465
rect 3508 3397 3542 3405
rect 3508 3371 3542 3397
rect 3508 3329 3542 3333
rect 3508 3299 3542 3329
rect 3508 3227 3542 3261
rect 3508 3159 3542 3189
rect 3508 3155 3542 3159
rect 3508 3091 3542 3117
rect 3508 3083 3542 3091
rect 3508 3023 3542 3045
rect 3508 3011 3542 3023
rect 3938 3530 3972 3540
rect 3938 3506 3972 3530
rect 3938 3462 3972 3464
rect 3938 3430 3972 3462
rect 3938 3360 3972 3388
rect 3938 3354 3972 3360
rect 3938 3292 3972 3312
rect 3938 3278 3972 3292
rect 3938 3224 3972 3236
rect 3938 3202 3972 3224
rect 3938 3156 3972 3160
rect 3938 3126 3972 3156
rect 3938 3054 3972 3084
rect 3938 3050 3972 3054
rect 2176 2931 2210 2935
rect 2176 2901 2210 2931
rect 3938 2986 3972 3008
rect 3938 2974 3972 2986
rect 3938 2918 3972 2932
rect 2176 2829 2210 2863
rect 2176 2761 2210 2791
rect 3938 2898 3972 2918
rect 2822 2850 2856 2873
rect 3119 2863 3135 2894
rect 3135 2863 3153 2894
rect 3195 2863 3205 2894
rect 3205 2863 3229 2894
rect 3271 2863 3274 2894
rect 3274 2863 3305 2894
rect 3346 2863 3378 2894
rect 3378 2863 3380 2894
rect 3421 2863 3447 2894
rect 3447 2863 3455 2894
rect 3119 2860 3153 2863
rect 3195 2860 3229 2863
rect 3271 2860 3305 2863
rect 3346 2860 3380 2863
rect 3421 2860 3455 2863
rect 2822 2839 2856 2850
rect 2822 2782 2856 2801
rect 2822 2767 2856 2782
rect 3938 2850 3972 2856
rect 3938 2822 3972 2850
rect 2176 2757 2210 2761
rect 2176 2693 2210 2719
rect 3938 2748 3972 2780
rect 3938 2746 3972 2748
rect 2176 2685 2210 2693
rect 2176 2625 2210 2647
rect 2176 2613 2210 2625
rect 3031 2676 3065 2710
rect 3110 2676 3144 2710
rect 3190 2676 3224 2710
rect 3270 2676 3304 2710
rect 3350 2676 3384 2710
rect 3430 2676 3464 2710
rect 3510 2676 3544 2710
rect 3590 2676 3624 2710
rect 3031 2580 3065 2614
rect 3110 2580 3144 2614
rect 3190 2580 3224 2614
rect 3270 2580 3304 2614
rect 3350 2580 3384 2614
rect 3430 2580 3464 2614
rect 3510 2580 3544 2614
rect 3590 2580 3624 2614
rect 3938 2680 3972 2705
rect 3938 2671 3972 2680
rect 3938 2612 3972 2630
rect 3938 2596 3972 2612
rect 2176 2557 2210 2575
rect 2176 2541 2210 2557
rect 3938 2544 3972 2555
rect -29134 2484 -29114 2508
rect -29114 2484 -29100 2508
rect -29134 2474 -29100 2484
rect -29046 2481 -29012 2508
rect -28958 2481 -28924 2508
rect -28870 2481 -28836 2508
rect -690 2498 -685 2523
rect -685 2498 -656 2523
rect -617 2498 -590 2523
rect -590 2498 -583 2523
rect -690 2489 -656 2498
rect -617 2489 -583 2498
rect -543 2489 -509 2523
rect 247 2490 248 2503
rect 248 2490 281 2503
rect -28189 2481 -28155 2487
rect -28115 2481 -28081 2487
rect -28041 2481 -28007 2487
rect -27967 2481 -27933 2487
rect -27893 2481 -27859 2487
rect -27819 2481 -27785 2487
rect -27745 2481 -27711 2487
rect -27671 2481 -27637 2487
rect -27597 2481 -27563 2487
rect -27523 2481 -27489 2487
rect -27449 2481 -27415 2487
rect -27375 2481 -27341 2487
rect -27301 2481 -27267 2487
rect -27227 2481 -27193 2487
rect -27153 2481 -27119 2487
rect -29046 2474 -29044 2481
rect -29044 2474 -29012 2481
rect -28958 2474 -28942 2481
rect -28942 2474 -28924 2481
rect -28870 2474 -28840 2481
rect -28840 2474 -28836 2481
rect -28189 2453 -28160 2481
rect -28160 2453 -28155 2481
rect -28115 2453 -28092 2481
rect -28092 2453 -28081 2481
rect -28041 2453 -28024 2481
rect -28024 2453 -28007 2481
rect -27967 2453 -27956 2481
rect -27956 2453 -27933 2481
rect -27893 2453 -27888 2481
rect -27888 2453 -27859 2481
rect -27819 2453 -27786 2481
rect -27786 2453 -27785 2481
rect -27745 2453 -27718 2481
rect -27718 2453 -27711 2481
rect -27671 2453 -27650 2481
rect -27650 2453 -27637 2481
rect -27597 2453 -27582 2481
rect -27582 2453 -27563 2481
rect -27523 2453 -27514 2481
rect -27514 2453 -27489 2481
rect -27449 2453 -27446 2481
rect -27446 2453 -27415 2481
rect -27375 2453 -27344 2481
rect -27344 2453 -27341 2481
rect -27301 2453 -27276 2481
rect -27276 2453 -27267 2481
rect -27227 2453 -27208 2481
rect -27208 2453 -27193 2481
rect -27153 2453 -27140 2481
rect -27140 2453 -27119 2481
rect -29134 2416 -29114 2435
rect -29114 2416 -29100 2435
rect -29134 2401 -29100 2416
rect -29046 2412 -29012 2435
rect -28958 2412 -28924 2435
rect -28870 2412 -28836 2435
rect -28189 2412 -28155 2414
rect -28115 2412 -28081 2414
rect -28041 2412 -28007 2414
rect -27967 2412 -27933 2414
rect -27893 2412 -27859 2414
rect -27819 2412 -27785 2414
rect -27745 2412 -27711 2414
rect -27671 2412 -27637 2414
rect -27597 2412 -27563 2414
rect -27523 2412 -27489 2414
rect -27449 2412 -27415 2414
rect -27375 2412 -27341 2414
rect -27301 2412 -27267 2414
rect -27227 2412 -27193 2414
rect -27153 2412 -27119 2414
rect -29046 2401 -29044 2412
rect -29044 2401 -29012 2412
rect -28958 2401 -28942 2412
rect -28942 2401 -28924 2412
rect -28870 2401 -28840 2412
rect -28840 2401 -28836 2412
rect -28189 2380 -28160 2412
rect -28160 2380 -28155 2412
rect -28115 2380 -28092 2412
rect -28092 2380 -28081 2412
rect -28041 2380 -28024 2412
rect -28024 2380 -28007 2412
rect -27967 2380 -27956 2412
rect -27956 2380 -27933 2412
rect -27893 2380 -27888 2412
rect -27888 2380 -27859 2412
rect -27819 2380 -27786 2412
rect -27786 2380 -27785 2412
rect -27745 2380 -27718 2412
rect -27718 2380 -27711 2412
rect -27671 2380 -27650 2412
rect -27650 2380 -27637 2412
rect -27597 2380 -27582 2412
rect -27582 2380 -27563 2412
rect -27523 2380 -27514 2412
rect -27514 2380 -27489 2412
rect -27449 2380 -27446 2412
rect -27446 2380 -27415 2412
rect -27375 2380 -27344 2412
rect -27344 2380 -27341 2412
rect -27301 2380 -27276 2412
rect -27276 2380 -27267 2412
rect -27227 2380 -27208 2412
rect -27208 2380 -27193 2412
rect -27153 2380 -27140 2412
rect -27140 2380 -27119 2412
rect 247 2469 281 2490
rect 247 2422 248 2431
rect 248 2422 281 2431
rect 247 2397 281 2422
rect 403 2490 404 2516
rect 404 2490 437 2516
rect 403 2482 437 2490
rect 403 2422 404 2444
rect 404 2422 437 2444
rect 403 2410 437 2422
rect 695 2490 696 2516
rect 696 2490 729 2516
rect 695 2482 729 2490
rect 695 2422 696 2444
rect 696 2422 729 2444
rect 695 2410 729 2422
rect 851 2490 852 2516
rect 852 2490 885 2516
rect 851 2482 885 2490
rect 851 2422 852 2444
rect 852 2422 885 2444
rect 851 2410 885 2422
rect 1134 2490 1135 2516
rect 1135 2490 1168 2516
rect 1134 2482 1168 2490
rect 1134 2422 1135 2444
rect 1135 2422 1168 2444
rect 1134 2410 1168 2422
rect 1494 2490 1495 2516
rect 1495 2490 1528 2516
rect 3938 2521 3972 2544
rect 1494 2482 1528 2490
rect 1494 2422 1495 2444
rect 1495 2422 1528 2444
rect 1494 2410 1528 2422
rect 1770 2455 1788 2481
rect 1788 2455 1804 2481
rect 1770 2447 1804 2455
rect 1770 2387 1788 2409
rect 1788 2387 1804 2409
rect 1770 2375 1804 2387
rect 1943 2455 1944 2481
rect 1944 2455 1977 2481
rect 1943 2447 1977 2455
rect 1943 2387 1944 2409
rect 1944 2387 1977 2409
rect 1943 2375 1977 2387
rect 2099 2455 2100 2481
rect 2100 2455 2133 2481
rect 2099 2447 2133 2455
rect 2099 2387 2100 2409
rect 2100 2387 2133 2409
rect 2099 2375 2133 2387
rect 3938 2476 3972 2480
rect 3938 2446 3972 2476
rect -29134 2348 -29114 2362
rect -29114 2348 -29100 2362
rect -29134 2328 -29100 2348
rect -29046 2343 -29012 2362
rect -28958 2343 -28924 2362
rect -28870 2343 -28836 2362
rect -29046 2328 -29044 2343
rect -29044 2328 -29012 2343
rect -28958 2328 -28942 2343
rect -28942 2328 -28924 2343
rect -28870 2328 -28840 2343
rect -28840 2328 -28836 2343
rect -28189 2309 -28160 2341
rect -28160 2309 -28155 2341
rect -28115 2309 -28092 2341
rect -28092 2309 -28081 2341
rect -28041 2309 -28024 2341
rect -28024 2309 -28007 2341
rect -27967 2309 -27956 2341
rect -27956 2309 -27933 2341
rect -27893 2309 -27888 2341
rect -27888 2309 -27859 2341
rect -27819 2309 -27786 2341
rect -27786 2309 -27785 2341
rect -27745 2309 -27718 2341
rect -27718 2309 -27711 2341
rect -27671 2309 -27650 2341
rect -27650 2309 -27637 2341
rect -27597 2309 -27582 2341
rect -27582 2309 -27563 2341
rect -27523 2309 -27514 2341
rect -27514 2309 -27489 2341
rect -27449 2309 -27446 2341
rect -27446 2309 -27415 2341
rect -27375 2309 -27344 2341
rect -27344 2309 -27341 2341
rect -27301 2309 -27276 2341
rect -27276 2309 -27267 2341
rect -27227 2309 -27208 2341
rect -27208 2309 -27193 2341
rect -27153 2309 -27140 2341
rect -27140 2309 -27119 2341
rect -28189 2307 -28155 2309
rect -28115 2307 -28081 2309
rect -28041 2307 -28007 2309
rect -27967 2307 -27933 2309
rect -27893 2307 -27859 2309
rect -27819 2307 -27785 2309
rect -27745 2307 -27711 2309
rect -27671 2307 -27637 2309
rect -27597 2307 -27563 2309
rect -27523 2307 -27489 2309
rect -27449 2307 -27415 2309
rect -27375 2307 -27341 2309
rect -27301 2307 -27267 2309
rect -27227 2307 -27193 2309
rect -27153 2307 -27119 2309
rect -29134 2280 -29114 2289
rect -29114 2280 -29100 2289
rect -29134 2255 -29100 2280
rect -29046 2274 -29012 2289
rect -28958 2274 -28924 2289
rect -28870 2274 -28836 2289
rect -29046 2255 -29044 2274
rect -29044 2255 -29012 2274
rect -28958 2255 -28942 2274
rect -28942 2255 -28924 2274
rect -28870 2255 -28840 2274
rect -28840 2255 -28836 2274
rect -28189 2240 -28160 2268
rect -28160 2240 -28155 2268
rect -28115 2240 -28092 2268
rect -28092 2240 -28081 2268
rect -28041 2240 -28024 2268
rect -28024 2240 -28007 2268
rect -27967 2240 -27956 2268
rect -27956 2240 -27933 2268
rect -27893 2240 -27888 2268
rect -27888 2240 -27859 2268
rect -27819 2240 -27786 2268
rect -27786 2240 -27785 2268
rect -27745 2240 -27718 2268
rect -27718 2240 -27711 2268
rect -27671 2240 -27650 2268
rect -27650 2240 -27637 2268
rect -27597 2240 -27582 2268
rect -27582 2240 -27563 2268
rect -27523 2240 -27514 2268
rect -27514 2240 -27489 2268
rect -27449 2240 -27446 2268
rect -27446 2240 -27415 2268
rect -27375 2240 -27344 2268
rect -27344 2240 -27341 2268
rect -27301 2240 -27276 2268
rect -27276 2240 -27267 2268
rect -27227 2240 -27208 2268
rect -27208 2240 -27193 2268
rect -27153 2240 -27140 2268
rect -27140 2240 -27119 2268
rect -28189 2234 -28155 2240
rect -28115 2234 -28081 2240
rect -28041 2234 -28007 2240
rect -27967 2234 -27933 2240
rect -27893 2234 -27859 2240
rect -27819 2234 -27785 2240
rect -27745 2234 -27711 2240
rect -27671 2234 -27637 2240
rect -27597 2234 -27563 2240
rect -27523 2234 -27489 2240
rect -27449 2234 -27415 2240
rect -27375 2234 -27341 2240
rect -27301 2234 -27267 2240
rect -27227 2234 -27193 2240
rect -27153 2234 -27119 2240
rect -29134 2212 -29114 2216
rect -29114 2212 -29100 2216
rect -29134 2182 -29100 2212
rect -29046 2205 -29012 2216
rect -28958 2205 -28924 2216
rect -28870 2205 -28836 2216
rect -29046 2182 -29044 2205
rect -29044 2182 -29012 2205
rect -28958 2182 -28942 2205
rect -28942 2182 -28924 2205
rect -28870 2182 -28840 2205
rect -28840 2182 -28836 2205
rect -28189 2171 -28160 2195
rect -28160 2171 -28155 2195
rect -28115 2171 -28092 2195
rect -28092 2171 -28081 2195
rect -28041 2171 -28024 2195
rect -28024 2171 -28007 2195
rect -27967 2171 -27956 2195
rect -27956 2171 -27933 2195
rect -27893 2171 -27888 2195
rect -27888 2171 -27859 2195
rect -27819 2171 -27786 2195
rect -27786 2171 -27785 2195
rect -27745 2171 -27718 2195
rect -27718 2171 -27711 2195
rect -27671 2171 -27650 2195
rect -27650 2171 -27637 2195
rect -27597 2171 -27582 2195
rect -27582 2171 -27563 2195
rect -27523 2171 -27514 2195
rect -27514 2171 -27489 2195
rect -27449 2171 -27446 2195
rect -27446 2171 -27415 2195
rect -27375 2171 -27344 2195
rect -27344 2171 -27341 2195
rect -27301 2171 -27276 2195
rect -27276 2171 -27267 2195
rect -27227 2171 -27208 2195
rect -27208 2171 -27193 2195
rect -27153 2171 -27140 2195
rect -27140 2171 -27119 2195
rect -28189 2161 -28155 2171
rect -28115 2161 -28081 2171
rect -28041 2161 -28007 2171
rect -27967 2161 -27933 2171
rect -27893 2161 -27859 2171
rect -27819 2161 -27785 2171
rect -27745 2161 -27711 2171
rect -27671 2161 -27637 2171
rect -27597 2161 -27563 2171
rect -27523 2161 -27489 2171
rect -27449 2161 -27415 2171
rect -27375 2161 -27341 2171
rect -27301 2161 -27267 2171
rect -27227 2161 -27193 2171
rect -27153 2161 -27119 2171
rect -29134 2110 -29100 2143
rect -29046 2136 -29012 2143
rect -28958 2136 -28924 2143
rect -28870 2136 -28836 2143
rect -29134 2109 -29114 2110
rect -29114 2109 -29100 2110
rect -29046 2109 -29044 2136
rect -29044 2109 -29012 2136
rect -28958 2109 -28942 2136
rect -28942 2109 -28924 2136
rect -28870 2109 -28840 2136
rect -28840 2109 -28836 2136
rect -28189 2102 -28160 2122
rect -28160 2102 -28155 2122
rect -28115 2102 -28092 2122
rect -28092 2102 -28081 2122
rect -28041 2102 -28024 2122
rect -28024 2102 -28007 2122
rect -27967 2102 -27956 2122
rect -27956 2102 -27933 2122
rect -27893 2102 -27888 2122
rect -27888 2102 -27859 2122
rect -27819 2102 -27786 2122
rect -27786 2102 -27785 2122
rect -27745 2102 -27718 2122
rect -27718 2102 -27711 2122
rect -27671 2102 -27650 2122
rect -27650 2102 -27637 2122
rect -27597 2102 -27582 2122
rect -27582 2102 -27563 2122
rect -27523 2102 -27514 2122
rect -27514 2102 -27489 2122
rect -27449 2102 -27446 2122
rect -27446 2102 -27415 2122
rect -27375 2102 -27344 2122
rect -27344 2102 -27341 2122
rect -27301 2102 -27276 2122
rect -27276 2102 -27267 2122
rect -27227 2102 -27208 2122
rect -27208 2102 -27193 2122
rect -27153 2102 -27140 2122
rect -27140 2102 -27119 2122
rect -28189 2088 -28155 2102
rect -28115 2088 -28081 2102
rect -28041 2088 -28007 2102
rect -27967 2088 -27933 2102
rect -27893 2088 -27859 2102
rect -27819 2088 -27785 2102
rect -27745 2088 -27711 2102
rect -27671 2088 -27637 2102
rect -27597 2088 -27563 2102
rect -27523 2088 -27489 2102
rect -27449 2088 -27415 2102
rect -27375 2088 -27341 2102
rect -27301 2088 -27267 2102
rect -27227 2088 -27193 2102
rect -27153 2088 -27119 2102
rect -29134 2042 -29100 2070
rect -29046 2067 -29012 2070
rect -28958 2067 -28924 2070
rect -28870 2067 -28836 2070
rect -29134 2036 -29114 2042
rect -29114 2036 -29100 2042
rect -29046 2036 -29012 2067
rect -28958 2036 -28924 2067
rect -28870 2036 -28836 2067
rect -28189 2015 -28155 2049
rect -28115 2015 -28081 2049
rect -28041 2015 -28007 2049
rect -27967 2015 -27933 2049
rect -27893 2015 -27859 2049
rect -27819 2015 -27785 2049
rect -27745 2015 -27711 2049
rect -27671 2015 -27637 2049
rect -27597 2015 -27563 2049
rect -27523 2015 -27489 2049
rect -27449 2015 -27415 2049
rect -27375 2015 -27341 2049
rect -27301 2015 -27267 2049
rect -27227 2015 -27193 2049
rect -27153 2015 -27119 2049
rect -29134 1974 -29100 1997
rect -29134 1963 -29114 1974
rect -29114 1963 -29100 1974
rect -29046 1963 -29012 1997
rect -28958 1963 -28924 1997
rect -28870 1963 -28836 1997
rect -28189 1942 -28155 1976
rect -28115 1942 -28081 1976
rect -28041 1942 -28007 1976
rect -27967 1942 -27933 1976
rect -27893 1942 -27859 1976
rect -27819 1942 -27785 1976
rect -27745 1942 -27711 1976
rect -27671 1942 -27637 1976
rect -27597 1942 -27563 1976
rect -27523 1942 -27489 1976
rect -27449 1942 -27415 1976
rect -27375 1942 -27341 1976
rect -27301 1942 -27267 1976
rect -27227 1942 -27193 1976
rect -27153 1942 -27119 1976
rect -29134 1906 -29100 1924
rect -29134 1890 -29114 1906
rect -29114 1890 -29100 1906
rect -29046 1890 -29012 1924
rect -28958 1890 -28924 1924
rect -28870 1890 -28836 1924
rect -28189 1869 -28155 1903
rect -28115 1869 -28081 1903
rect -28041 1869 -28007 1903
rect -27967 1869 -27933 1903
rect -27893 1869 -27859 1903
rect -27819 1869 -27785 1903
rect -27745 1869 -27711 1903
rect -27671 1869 -27637 1903
rect -27597 1869 -27563 1903
rect -27523 1869 -27489 1903
rect -27449 1869 -27415 1903
rect -27375 1869 -27341 1903
rect -27301 1869 -27267 1903
rect -27227 1869 -27193 1903
rect -27153 1869 -27119 1903
rect -29134 1838 -29100 1851
rect -29134 1817 -29114 1838
rect -29114 1817 -29100 1838
rect -29046 1817 -29012 1851
rect -28958 1817 -28924 1851
rect -28870 1817 -28836 1851
rect -28189 1796 -28155 1830
rect -28115 1796 -28081 1830
rect -28041 1796 -28007 1830
rect -27967 1796 -27933 1830
rect -27893 1796 -27859 1830
rect -27819 1796 -27785 1830
rect -27745 1796 -27711 1830
rect -27671 1796 -27637 1830
rect -27597 1796 -27563 1830
rect -27523 1796 -27489 1830
rect -27449 1796 -27415 1830
rect -27375 1796 -27341 1830
rect -27301 1796 -27267 1830
rect -27227 1796 -27193 1830
rect -27153 1796 -27119 1830
rect -29134 1770 -29100 1778
rect -29134 1744 -29114 1770
rect -29114 1744 -29100 1770
rect -29046 1744 -29012 1778
rect -28958 1744 -28924 1778
rect -28870 1744 -28836 1778
rect -28189 1723 -28155 1757
rect -28115 1723 -28081 1757
rect -28041 1723 -28007 1757
rect -27967 1723 -27933 1757
rect -27893 1723 -27859 1757
rect -27819 1723 -27785 1757
rect -27745 1723 -27711 1757
rect -27671 1723 -27637 1757
rect -27597 1723 -27563 1757
rect -27523 1723 -27489 1757
rect -27449 1723 -27415 1757
rect -27375 1723 -27341 1757
rect -27301 1723 -27267 1757
rect -27227 1723 -27193 1757
rect -27153 1723 -27119 1757
rect -29134 1702 -29100 1705
rect -29134 1671 -29114 1702
rect -29114 1671 -29100 1702
rect -29046 1671 -29012 1705
rect -28958 1671 -28924 1705
rect -28870 1671 -28836 1705
rect -28189 1650 -28155 1684
rect -28115 1650 -28081 1684
rect -28041 1650 -28007 1684
rect -27967 1650 -27933 1684
rect -27893 1650 -27859 1684
rect -27819 1650 -27785 1684
rect -27745 1650 -27711 1684
rect -27671 1650 -27637 1684
rect -27597 1650 -27563 1684
rect -27523 1650 -27489 1684
rect -27449 1650 -27415 1684
rect -27375 1650 -27341 1684
rect -27301 1650 -27267 1684
rect -27227 1650 -27193 1684
rect -27153 1650 -27119 1684
rect -29134 1600 -29114 1632
rect -29114 1600 -29100 1632
rect -29134 1598 -29100 1600
rect -29046 1598 -29012 1632
rect -28958 1598 -28924 1632
rect -28870 1598 -28836 1632
rect -28189 1577 -28155 1611
rect -28115 1577 -28081 1611
rect -28041 1577 -28007 1611
rect -27967 1577 -27933 1611
rect -27893 1577 -27859 1611
rect -27819 1577 -27785 1611
rect -27745 1577 -27711 1611
rect -27671 1577 -27637 1611
rect -27597 1577 -27563 1611
rect -27523 1577 -27489 1611
rect -27449 1577 -27415 1611
rect -27375 1577 -27341 1611
rect -27301 1577 -27267 1611
rect -27227 1577 -27193 1611
rect -27153 1577 -27119 1611
rect -29134 1532 -29114 1559
rect -29114 1532 -29100 1559
rect -29134 1525 -29100 1532
rect -29046 1525 -29012 1559
rect -28958 1525 -28924 1559
rect -28870 1525 -28836 1559
rect -28189 1504 -28155 1538
rect -28115 1504 -28081 1538
rect -28041 1504 -28007 1538
rect -27967 1504 -27933 1538
rect -27893 1504 -27859 1538
rect -27819 1504 -27785 1538
rect -27745 1504 -27711 1538
rect -27671 1504 -27637 1538
rect -27597 1504 -27563 1538
rect -27523 1504 -27489 1538
rect -27449 1504 -27415 1538
rect -27375 1504 -27341 1538
rect -27301 1504 -27267 1538
rect -27227 1504 -27193 1538
rect -27153 1504 -27119 1538
rect -29134 1464 -29114 1486
rect -29114 1464 -29100 1486
rect -29134 1452 -29100 1464
rect -29046 1452 -29012 1486
rect -28958 1452 -28924 1486
rect -28870 1452 -28836 1486
rect -28189 1431 -28155 1465
rect -28115 1431 -28081 1465
rect -28041 1431 -28007 1465
rect -27967 1431 -27933 1465
rect -27893 1431 -27859 1465
rect -27819 1431 -27785 1465
rect -27745 1431 -27711 1465
rect -27671 1431 -27637 1465
rect -27597 1431 -27563 1465
rect -27523 1431 -27489 1465
rect -27449 1431 -27415 1465
rect -27375 1431 -27341 1465
rect -27301 1431 -27267 1465
rect -27227 1431 -27193 1465
rect -27153 1431 -27119 1465
rect -29134 1396 -29114 1413
rect -29114 1396 -29100 1413
rect -29134 1379 -29100 1396
rect -29046 1379 -29012 1413
rect -28958 1379 -28924 1413
rect -28870 1379 -28836 1413
rect -28189 1358 -28155 1392
rect -28115 1358 -28081 1392
rect -28041 1358 -28007 1392
rect -27967 1358 -27933 1392
rect -27893 1358 -27859 1392
rect -27819 1358 -27785 1392
rect -27745 1358 -27711 1392
rect -27671 1358 -27637 1392
rect -27597 1358 -27563 1392
rect -27523 1358 -27489 1392
rect -27449 1358 -27415 1392
rect -27375 1358 -27341 1392
rect -27301 1358 -27267 1392
rect -27227 1358 -27193 1392
rect -27153 1358 -27119 1392
rect -29134 1328 -29114 1340
rect -29114 1328 -29100 1340
rect -29134 1306 -29100 1328
rect -29046 1306 -29012 1340
rect -28958 1306 -28924 1340
rect -28870 1306 -28836 1340
rect -28189 1285 -28155 1319
rect -28115 1285 -28081 1319
rect -28041 1285 -28007 1319
rect -27967 1285 -27933 1319
rect -27893 1285 -27859 1319
rect -27819 1285 -27785 1319
rect -27745 1285 -27711 1319
rect -27671 1285 -27637 1319
rect -27597 1285 -27563 1319
rect -27523 1285 -27489 1319
rect -27449 1285 -27415 1319
rect -27375 1285 -27341 1319
rect -27301 1285 -27267 1319
rect -27227 1285 -27193 1319
rect -27153 1285 -27119 1319
rect -29134 1260 -29114 1267
rect -29114 1260 -29100 1267
rect -29134 1233 -29100 1260
rect -29046 1233 -29012 1267
rect -28958 1233 -28924 1267
rect -28870 1233 -28836 1267
rect -28189 1212 -28155 1246
rect -28115 1212 -28081 1246
rect -28041 1212 -28007 1246
rect -27967 1212 -27933 1246
rect -27893 1212 -27859 1246
rect -27819 1212 -27785 1246
rect -27745 1212 -27711 1246
rect -27671 1212 -27637 1246
rect -27597 1212 -27563 1246
rect -27523 1212 -27489 1246
rect -27449 1212 -27415 1246
rect -27375 1212 -27341 1246
rect -27301 1212 -27267 1246
rect -27227 1212 -27193 1246
rect -27153 1212 -27119 1246
rect -29134 1192 -29114 1194
rect -29114 1192 -29100 1194
rect -29134 1160 -29100 1192
rect -29046 1160 -29012 1194
rect -28958 1160 -28924 1194
rect -28870 1160 -28836 1194
rect -28189 1139 -28155 1173
rect -28115 1139 -28081 1173
rect -28041 1139 -28007 1173
rect -27967 1139 -27933 1173
rect -27893 1139 -27859 1173
rect -27819 1139 -27785 1173
rect -27745 1139 -27711 1173
rect -27671 1139 -27637 1173
rect -27597 1139 -27563 1173
rect -27523 1139 -27489 1173
rect -27449 1139 -27415 1173
rect -27375 1139 -27341 1173
rect -27301 1139 -27267 1173
rect -27227 1139 -27193 1173
rect -27153 1139 -27119 1173
rect -29134 1090 -29100 1121
rect -29134 1087 -29114 1090
rect -29114 1087 -29100 1090
rect -29046 1087 -29012 1121
rect -28958 1087 -28924 1121
rect -28870 1087 -28836 1121
rect -28189 1066 -28155 1100
rect -28115 1066 -28081 1100
rect -28041 1066 -28007 1100
rect -27967 1066 -27933 1100
rect -27893 1066 -27859 1100
rect -27819 1066 -27785 1100
rect -27745 1066 -27711 1100
rect -27671 1066 -27637 1100
rect -27597 1066 -27563 1100
rect -27523 1066 -27489 1100
rect -27449 1066 -27415 1100
rect -27375 1066 -27341 1100
rect -27301 1066 -27267 1100
rect -27227 1066 -27193 1100
rect -27153 1066 -27119 1100
rect -29134 1022 -29100 1048
rect -29134 1014 -29114 1022
rect -29114 1014 -29100 1022
rect -29046 1014 -29012 1048
rect -28958 1014 -28924 1048
rect -28870 1014 -28836 1048
rect -28189 994 -28155 1028
rect -28115 994 -28081 1028
rect -28041 994 -28007 1028
rect -27967 994 -27933 1028
rect -27893 994 -27859 1028
rect -27819 994 -27785 1028
rect -27745 994 -27711 1028
rect -27671 994 -27637 1028
rect -27597 994 -27563 1028
rect -27523 994 -27489 1028
rect -27449 994 -27415 1028
rect -27375 994 -27341 1028
rect -27301 994 -27267 1028
rect -27227 994 -27193 1028
rect -27153 994 -27119 1028
rect -29134 954 -29100 975
rect -29134 941 -29114 954
rect -29114 941 -29100 954
rect -29046 941 -29012 975
rect -28958 941 -28924 975
rect -28870 941 -28836 975
rect -28189 922 -28155 956
rect -28115 922 -28081 956
rect -28041 922 -28007 956
rect -27967 922 -27933 956
rect -27893 922 -27859 956
rect -27819 922 -27785 956
rect -27745 922 -27711 956
rect -27671 922 -27637 956
rect -27597 922 -27563 956
rect -27523 922 -27489 956
rect -27449 922 -27415 956
rect -27375 922 -27341 956
rect -27301 922 -27267 956
rect -27227 922 -27193 956
rect -27153 922 -27119 956
rect -29134 886 -29100 902
rect -29134 868 -29114 886
rect -29114 868 -29100 886
rect -29046 868 -29012 902
rect -28958 868 -28924 902
rect -28870 868 -28836 902
rect -28189 850 -28155 884
rect -28115 850 -28081 884
rect -28041 850 -28007 884
rect -27967 850 -27933 884
rect -27893 850 -27859 884
rect -27819 850 -27785 884
rect -27745 850 -27711 884
rect -27671 850 -27637 884
rect -27597 850 -27563 884
rect -27523 850 -27489 884
rect -27449 850 -27415 884
rect -27375 850 -27341 884
rect -27301 850 -27267 884
rect -27227 850 -27193 884
rect -27153 850 -27119 884
rect -29134 818 -29100 829
rect -29134 795 -29114 818
rect -29114 795 -29100 818
rect -29046 795 -29012 829
rect -28958 795 -28924 829
rect -28870 795 -28836 829
rect -28189 778 -28155 812
rect -28115 778 -28081 812
rect -28041 778 -28007 812
rect -27967 778 -27933 812
rect -27893 778 -27859 812
rect -27819 778 -27785 812
rect -27745 778 -27711 812
rect -27671 778 -27637 812
rect -27597 778 -27563 812
rect -27523 778 -27489 812
rect -27449 778 -27415 812
rect -27375 778 -27341 812
rect -27301 778 -27267 812
rect -27227 778 -27193 812
rect -27153 778 -27119 812
rect -29134 750 -29100 756
rect -29134 722 -29114 750
rect -29114 722 -29100 750
rect -29046 722 -29012 756
rect -28958 722 -28924 756
rect -28870 722 -28836 756
rect -28189 706 -28155 740
rect -28115 706 -28081 740
rect -28041 706 -28007 740
rect -27967 706 -27933 740
rect -27893 706 -27859 740
rect -27819 706 -27785 740
rect -27745 706 -27711 740
rect -27671 706 -27637 740
rect -27597 706 -27563 740
rect -27523 706 -27489 740
rect -27449 706 -27415 740
rect -27375 706 -27341 740
rect -27301 706 -27267 740
rect -27227 706 -27193 740
rect -27153 706 -27119 740
rect -29134 682 -29100 683
rect -29134 649 -29114 682
rect -29114 649 -29100 682
rect -29046 649 -29012 683
rect -28958 649 -28924 683
rect -28870 649 -28836 683
rect -28189 634 -28155 668
rect -28115 634 -28081 668
rect -28041 634 -28007 668
rect -27967 634 -27933 668
rect -27893 634 -27859 668
rect -27819 634 -27785 668
rect -27745 634 -27711 668
rect -27671 634 -27637 668
rect -27597 634 -27563 668
rect -27523 634 -27489 668
rect -27449 634 -27415 668
rect -27375 634 -27341 668
rect -27301 634 -27267 668
rect -27227 634 -27193 668
rect -27153 634 -27119 668
rect -29134 580 -29114 610
rect -29114 580 -29100 610
rect -29134 576 -29100 580
rect -29046 576 -29012 610
rect -28958 576 -28924 610
rect -28870 576 -28836 610
rect -28189 562 -28155 596
rect -28115 562 -28081 596
rect -28041 562 -28007 596
rect -27967 562 -27933 596
rect -27893 562 -27859 596
rect -27819 562 -27785 596
rect -27745 562 -27711 596
rect -27671 562 -27637 596
rect -27597 562 -27563 596
rect -27523 562 -27489 596
rect -27449 562 -27415 596
rect -27375 562 -27341 596
rect -27301 562 -27267 596
rect -27227 562 -27193 596
rect -27153 562 -27119 596
rect -29134 512 -29114 537
rect -29114 512 -29100 537
rect -29134 503 -29100 512
rect -29046 503 -29012 537
rect -28958 503 -28924 537
rect -28870 503 -28836 537
rect -28189 490 -28155 524
rect -28115 490 -28081 524
rect -28041 490 -28007 524
rect -27967 490 -27933 524
rect -27893 490 -27859 524
rect -27819 490 -27785 524
rect -27745 490 -27711 524
rect -27671 490 -27637 524
rect -27597 490 -27563 524
rect -27523 490 -27489 524
rect -27449 490 -27415 524
rect -27375 490 -27341 524
rect -27301 490 -27267 524
rect -27227 490 -27193 524
rect -27153 490 -27119 524
rect -29134 444 -29114 464
rect -29114 444 -29100 464
rect -29134 430 -29100 444
rect -29046 430 -29012 464
rect -28958 430 -28924 464
rect -28870 430 -28836 464
rect -28189 418 -28155 452
rect -28115 418 -28081 452
rect -28041 418 -28007 452
rect -27967 418 -27933 452
rect -27893 418 -27859 452
rect -27819 418 -27785 452
rect -27745 418 -27711 452
rect -27671 418 -27637 452
rect -27597 418 -27563 452
rect -27523 418 -27489 452
rect -27449 418 -27415 452
rect -27375 418 -27341 452
rect -27301 418 -27267 452
rect -27227 418 -27193 452
rect -27153 418 -27119 452
rect -29134 376 -29114 391
rect -29114 376 -29100 391
rect -29134 357 -29100 376
rect -29046 357 -29012 391
rect -28958 357 -28924 391
rect -28870 357 -28836 391
rect -28189 346 -28155 380
rect -28115 346 -28081 380
rect -28041 346 -28007 380
rect -27967 346 -27933 380
rect -27893 346 -27859 380
rect -27819 346 -27785 380
rect -27745 346 -27711 380
rect -27671 346 -27637 380
rect -27597 346 -27563 380
rect -27523 346 -27489 380
rect -27449 346 -27415 380
rect -27375 346 -27341 380
rect -27301 346 -27267 380
rect -27227 346 -27193 380
rect -27153 346 -27119 380
rect -29134 308 -29114 318
rect -29114 308 -29100 318
rect -29134 284 -29100 308
rect -29046 284 -29012 318
rect -28958 284 -28924 318
rect -28870 284 -28836 318
rect -28189 274 -28155 308
rect -28115 274 -28081 308
rect -28041 274 -28007 308
rect -27967 274 -27933 308
rect -27893 274 -27859 308
rect -27819 274 -27785 308
rect -27745 274 -27711 308
rect -27671 274 -27637 308
rect -27597 274 -27563 308
rect -27523 274 -27489 308
rect -27449 274 -27415 308
rect -27375 274 -27341 308
rect -27301 274 -27267 308
rect -27227 274 -27193 308
rect -27153 274 -27119 308
rect -29134 240 -29114 245
rect -29114 240 -29100 245
rect -29134 211 -29100 240
rect -29046 211 -29012 245
rect -28958 211 -28924 245
rect -28870 211 -28836 245
rect -28189 202 -28155 236
rect -28115 202 -28081 236
rect -28041 202 -28007 236
rect -27967 202 -27933 236
rect -27893 202 -27859 236
rect -27819 202 -27785 236
rect -27745 202 -27711 236
rect -27671 202 -27637 236
rect -27597 202 -27563 236
rect -27523 202 -27489 236
rect -27449 202 -27415 236
rect -27375 202 -27341 236
rect -27301 202 -27267 236
rect -27227 202 -27193 236
rect -27153 202 -27119 236
rect -29134 138 -29100 172
rect -29046 138 -29012 172
rect -28958 138 -28924 172
rect -28870 138 -28836 172
rect -28189 130 -28155 164
rect -28115 130 -28081 164
rect -28041 130 -28007 164
rect -27967 130 -27933 164
rect -27893 130 -27859 164
rect -27819 130 -27785 164
rect -27745 130 -27711 164
rect -27671 130 -27637 164
rect -27597 130 -27563 164
rect -27523 130 -27489 164
rect -27449 130 -27415 164
rect -27375 130 -27341 164
rect -27301 130 -27267 164
rect -27227 130 -27193 164
rect -27153 130 -27119 164
rect -29134 70 -29100 99
rect -29134 65 -29114 70
rect -29114 65 -29100 70
rect -29046 65 -29012 99
rect -28958 65 -28924 99
rect -28870 65 -28836 99
rect -28189 58 -28155 92
rect -28115 58 -28081 92
rect -28041 58 -28007 92
rect -27967 58 -27933 92
rect -27893 58 -27859 92
rect -27819 58 -27785 92
rect -27745 58 -27711 92
rect -27671 58 -27637 92
rect -27597 58 -27563 92
rect -27523 58 -27489 92
rect -27449 58 -27415 92
rect -27375 58 -27341 92
rect -27301 58 -27267 92
rect -27227 58 -27193 92
rect -27153 58 -27119 92
rect -29134 2 -29100 26
rect -29134 -8 -29114 2
rect -29114 -8 -29100 2
rect -29046 -8 -29012 26
rect -28958 -8 -28924 26
rect -28870 -8 -28836 26
rect -28189 -14 -28155 20
rect -28115 -14 -28081 20
rect -28041 -14 -28007 20
rect -27967 -14 -27933 20
rect -27893 -14 -27859 20
rect -27819 -14 -27785 20
rect -27745 -14 -27711 20
rect -27671 -14 -27637 20
rect -27597 -14 -27563 20
rect -27523 -14 -27489 20
rect -27449 -14 -27415 20
rect -27375 -14 -27341 20
rect -27301 -14 -27267 20
rect -27227 -14 -27193 20
rect -27153 -14 -27119 20
rect -29134 -66 -29100 -47
rect -29134 -81 -29114 -66
rect -29114 -81 -29100 -66
rect -29046 -81 -29012 -47
rect -28958 -81 -28924 -47
rect -28870 -81 -28836 -47
rect -28189 -86 -28155 -52
rect -28115 -86 -28081 -52
rect -28041 -86 -28007 -52
rect -27967 -86 -27933 -52
rect -27893 -86 -27859 -52
rect -27819 -86 -27785 -52
rect -27745 -86 -27711 -52
rect -27671 -86 -27637 -52
rect -27597 -86 -27563 -52
rect -27523 -86 -27489 -52
rect -27449 -86 -27415 -52
rect -27375 -86 -27341 -52
rect -27301 -86 -27267 -52
rect -27227 -86 -27193 -52
rect -27153 -86 -27119 -52
rect -29134 -134 -29100 -120
rect -29134 -154 -29114 -134
rect -29114 -154 -29100 -134
rect -29046 -154 -29012 -120
rect -28958 -154 -28924 -120
rect -28870 -154 -28836 -120
rect -28189 -158 -28155 -124
rect -28115 -158 -28081 -124
rect -28041 -158 -28007 -124
rect -27967 -158 -27933 -124
rect -27893 -158 -27859 -124
rect -27819 -158 -27785 -124
rect -27745 -158 -27711 -124
rect -27671 -158 -27637 -124
rect -27597 -158 -27563 -124
rect -27523 -158 -27489 -124
rect -27449 -158 -27415 -124
rect -27375 -158 -27341 -124
rect -27301 -158 -27267 -124
rect -27227 -158 -27193 -124
rect -27153 -158 -27119 -124
rect -29134 -202 -29100 -193
rect -29134 -227 -29114 -202
rect -29114 -227 -29100 -202
rect -29046 -227 -29012 -193
rect -28958 -227 -28924 -193
rect -28870 -227 -28836 -193
rect -28189 -230 -28155 -196
rect -28115 -230 -28081 -196
rect -28041 -230 -28007 -196
rect -27967 -230 -27933 -196
rect -27893 -230 -27859 -196
rect -27819 -230 -27785 -196
rect -27745 -230 -27711 -196
rect -27671 -230 -27637 -196
rect -27597 -230 -27563 -196
rect -27523 -230 -27489 -196
rect -27449 -230 -27415 -196
rect -27375 -230 -27341 -196
rect -27301 -230 -27267 -196
rect -27227 -230 -27193 -196
rect -27153 -230 -27119 -196
rect -29134 -270 -29100 -266
rect -29134 -300 -29114 -270
rect -29114 -300 -29100 -270
rect -29046 -300 -29012 -266
rect -28958 -300 -28924 -266
rect -28870 -300 -28836 -266
rect -28189 -302 -28155 -268
rect -28115 -302 -28081 -268
rect -28041 -302 -28007 -268
rect -27967 -302 -27933 -268
rect -27893 -302 -27859 -268
rect -27819 -302 -27785 -268
rect -27745 -302 -27711 -268
rect -27671 -302 -27637 -268
rect -27597 -302 -27563 -268
rect -27523 -302 -27489 -268
rect -27449 -302 -27415 -268
rect -27375 -302 -27341 -268
rect -27301 -302 -27267 -268
rect -27227 -302 -27193 -268
rect -27153 -302 -27119 -268
rect -29134 -372 -29114 -339
rect -29114 -372 -29100 -339
rect -29134 -373 -29100 -372
rect -29046 -373 -29012 -339
rect -28958 -373 -28924 -339
rect -28870 -373 -28836 -339
rect -28189 -374 -28155 -340
rect -28115 -374 -28081 -340
rect -28041 -374 -28007 -340
rect -27967 -374 -27933 -340
rect -27893 -374 -27859 -340
rect -27819 -374 -27785 -340
rect -27745 -374 -27711 -340
rect -27671 -374 -27637 -340
rect -27597 -374 -27563 -340
rect -27523 -374 -27489 -340
rect -27449 -374 -27415 -340
rect -27375 -374 -27341 -340
rect -27301 -374 -27267 -340
rect -27227 -374 -27193 -340
rect -27153 -374 -27119 -340
rect -29134 -440 -29114 -412
rect -29114 -440 -29100 -412
rect -29134 -446 -29100 -440
rect -29046 -446 -29012 -412
rect -28958 -446 -28924 -412
rect -28870 -446 -28836 -412
rect -28189 -446 -28155 -412
rect -28115 -446 -28081 -412
rect -28041 -446 -28007 -412
rect -27967 -446 -27933 -412
rect -27893 -446 -27859 -412
rect -27819 -446 -27785 -412
rect -27745 -446 -27711 -412
rect -27671 -446 -27637 -412
rect -27597 -446 -27563 -412
rect -27523 -446 -27489 -412
rect -27449 -446 -27415 -412
rect -27375 -446 -27341 -412
rect -27301 -446 -27267 -412
rect -27227 -446 -27193 -412
rect -27153 -446 -27119 -412
rect -29134 -508 -29114 -485
rect -29114 -508 -29100 -485
rect -29134 -519 -29100 -508
rect -29046 -519 -29012 -485
rect -28958 -519 -28924 -485
rect -28870 -519 -28836 -485
rect -28189 -518 -28155 -484
rect -28115 -518 -28081 -484
rect -28041 -518 -28007 -484
rect -27967 -518 -27933 -484
rect -27893 -518 -27859 -484
rect -27819 -518 -27785 -484
rect -27745 -518 -27711 -484
rect -27671 -518 -27637 -484
rect -27597 -518 -27563 -484
rect -27523 -518 -27489 -484
rect -27449 -518 -27415 -484
rect -27375 -518 -27341 -484
rect -27301 -518 -27267 -484
rect -27227 -518 -27193 -484
rect -27153 -518 -27119 -484
rect -29134 -576 -29114 -558
rect -29114 -576 -29100 -558
rect -29134 -592 -29100 -576
rect -29046 -592 -29012 -558
rect -28958 -592 -28924 -558
rect -28870 -592 -28836 -558
rect -28189 -590 -28155 -556
rect -28115 -590 -28081 -556
rect -28041 -590 -28007 -556
rect -27967 -590 -27933 -556
rect -27893 -590 -27859 -556
rect -27819 -590 -27785 -556
rect -27745 -590 -27711 -556
rect -27671 -590 -27637 -556
rect -27597 -590 -27563 -556
rect -27523 -590 -27489 -556
rect -27449 -590 -27415 -556
rect -27375 -590 -27341 -556
rect -27301 -590 -27267 -556
rect -27227 -590 -27193 -556
rect -27153 -590 -27119 -556
rect -29134 -644 -29114 -631
rect -29114 -644 -29100 -631
rect -29134 -665 -29100 -644
rect -29046 -665 -29012 -631
rect -28958 -665 -28924 -631
rect -28870 -665 -28836 -631
rect -28189 -662 -28155 -628
rect -28115 -662 -28081 -628
rect -28041 -662 -28007 -628
rect -27967 -662 -27933 -628
rect -27893 -662 -27859 -628
rect -27819 -662 -27785 -628
rect -27745 -662 -27711 -628
rect -27671 -662 -27637 -628
rect -27597 -662 -27563 -628
rect -27523 -662 -27489 -628
rect -27449 -662 -27415 -628
rect -27375 -662 -27341 -628
rect -27301 -662 -27267 -628
rect -27227 -662 -27193 -628
rect -27153 -662 -27119 -628
rect -29134 -712 -29114 -704
rect -29114 -712 -29100 -704
rect -29134 -738 -29100 -712
rect -29046 -738 -29012 -704
rect -28958 -738 -28924 -704
rect -28870 -738 -28836 -704
rect -28189 -734 -28155 -700
rect -28115 -734 -28081 -700
rect -28041 -734 -28007 -700
rect -27967 -734 -27933 -700
rect -27893 -734 -27859 -700
rect -27819 -734 -27785 -700
rect -27745 -734 -27711 -700
rect -27671 -734 -27637 -700
rect -27597 -734 -27563 -700
rect -27523 -734 -27489 -700
rect -27449 -734 -27415 -700
rect -27375 -734 -27341 -700
rect -27301 -734 -27267 -700
rect -27227 -734 -27193 -700
rect -27153 -734 -27119 -700
rect -29134 -780 -29114 -777
rect -29114 -780 -29100 -777
rect -29134 -811 -29100 -780
rect -29046 -811 -29012 -777
rect -28958 -811 -28924 -777
rect -28870 -811 -28836 -777
rect -28189 -806 -28155 -772
rect -28115 -806 -28081 -772
rect -28041 -806 -28007 -772
rect -27967 -806 -27933 -772
rect -27893 -806 -27859 -772
rect -27819 -806 -27785 -772
rect -27745 -806 -27711 -772
rect -27671 -806 -27637 -772
rect -27597 -806 -27563 -772
rect -27523 -806 -27489 -772
rect -27449 -806 -27415 -772
rect -27375 -806 -27341 -772
rect -27301 -806 -27267 -772
rect -27227 -806 -27193 -772
rect -27153 -806 -27119 -772
rect -29134 -882 -29100 -849
rect -29134 -883 -29114 -882
rect -29114 -883 -29100 -882
rect -29046 -883 -29012 -849
rect -28958 -883 -28924 -849
rect -28870 -883 -28836 -849
rect -28189 -878 -28155 -844
rect -28115 -878 -28081 -844
rect -28041 -878 -28007 -844
rect -27967 -878 -27933 -844
rect -27893 -878 -27859 -844
rect -27819 -878 -27785 -844
rect -27745 -878 -27711 -844
rect -27671 -878 -27637 -844
rect -27597 -878 -27563 -844
rect -27523 -878 -27489 -844
rect -27449 -878 -27415 -844
rect -27375 -878 -27341 -844
rect -27301 -878 -27267 -844
rect -27227 -878 -27193 -844
rect -27153 -878 -27119 -844
rect -29134 -950 -29100 -921
rect -29134 -955 -29114 -950
rect -29114 -955 -29100 -950
rect -29046 -955 -29012 -921
rect -28958 -955 -28924 -921
rect -28870 -955 -28836 -921
rect -28189 -950 -28155 -916
rect -28115 -950 -28081 -916
rect -28041 -950 -28007 -916
rect -27967 -950 -27933 -916
rect -27893 -950 -27859 -916
rect -27819 -950 -27785 -916
rect -27745 -950 -27711 -916
rect -27671 -950 -27637 -916
rect -27597 -950 -27563 -916
rect -27523 -950 -27489 -916
rect -27449 -950 -27415 -916
rect -27375 -950 -27341 -916
rect -27301 -950 -27267 -916
rect -27227 -950 -27193 -916
rect -27153 -950 -27119 -916
rect -29134 -1018 -29100 -993
rect -29134 -1027 -29114 -1018
rect -29114 -1027 -29100 -1018
rect -29046 -1027 -29012 -993
rect -28958 -1027 -28924 -993
rect -28870 -1027 -28836 -993
rect -28189 -1022 -28155 -988
rect -28115 -1022 -28081 -988
rect -28041 -1022 -28007 -988
rect -27967 -1022 -27933 -988
rect -27893 -1022 -27859 -988
rect -27819 -1022 -27785 -988
rect -27745 -1022 -27711 -988
rect -27671 -1022 -27637 -988
rect -27597 -1022 -27563 -988
rect -27523 -1022 -27489 -988
rect -27449 -1022 -27415 -988
rect -27375 -1022 -27341 -988
rect -27301 -1022 -27267 -988
rect -27227 -1022 -27193 -988
rect -27153 -1022 -27119 -988
rect -29134 -1086 -29100 -1065
rect -29134 -1099 -29114 -1086
rect -29114 -1099 -29100 -1086
rect -29046 -1099 -29012 -1065
rect -28958 -1099 -28924 -1065
rect -28870 -1099 -28836 -1065
rect -28189 -1094 -28155 -1060
rect -28115 -1094 -28081 -1060
rect -28041 -1094 -28007 -1060
rect -27967 -1094 -27933 -1060
rect -27893 -1094 -27859 -1060
rect -27819 -1094 -27785 -1060
rect -27745 -1094 -27711 -1060
rect -27671 -1094 -27637 -1060
rect -27597 -1094 -27563 -1060
rect -27523 -1094 -27489 -1060
rect -27449 -1094 -27415 -1060
rect -27375 -1094 -27341 -1060
rect -27301 -1094 -27267 -1060
rect -27227 -1094 -27193 -1060
rect -27153 -1094 -27119 -1060
rect -29134 -1154 -29100 -1137
rect -29134 -1171 -29114 -1154
rect -29114 -1171 -29100 -1154
rect -29046 -1171 -29012 -1137
rect -28958 -1171 -28924 -1137
rect -28870 -1171 -28836 -1137
rect -28189 -1166 -28155 -1132
rect -28115 -1166 -28081 -1132
rect -28041 -1166 -28007 -1132
rect -27967 -1166 -27933 -1132
rect -27893 -1166 -27859 -1132
rect -27819 -1166 -27785 -1132
rect -27745 -1166 -27711 -1132
rect -27671 -1166 -27637 -1132
rect -27597 -1166 -27563 -1132
rect -27523 -1166 -27489 -1132
rect -27449 -1166 -27415 -1132
rect -27375 -1166 -27341 -1132
rect -27301 -1166 -27267 -1132
rect -27227 -1166 -27193 -1132
rect -27153 -1166 -27119 -1132
rect -29134 -1222 -29100 -1209
rect -29134 -1243 -29114 -1222
rect -29114 -1243 -29100 -1222
rect -29046 -1243 -29012 -1209
rect -28958 -1243 -28924 -1209
rect -28870 -1243 -28836 -1209
rect -28189 -1238 -28155 -1204
rect -28115 -1238 -28081 -1204
rect -28041 -1238 -28007 -1204
rect -27967 -1238 -27933 -1204
rect -27893 -1238 -27859 -1204
rect -27819 -1238 -27785 -1204
rect -27745 -1238 -27711 -1204
rect -27671 -1238 -27637 -1204
rect -27597 -1238 -27563 -1204
rect -27523 -1238 -27489 -1204
rect -27449 -1238 -27415 -1204
rect -27375 -1238 -27341 -1204
rect -27301 -1238 -27267 -1204
rect -27227 -1238 -27193 -1204
rect -27153 -1238 -27119 -1204
rect -29134 -1290 -29100 -1281
rect -29134 -1315 -29114 -1290
rect -29114 -1315 -29100 -1290
rect -29046 -1315 -29012 -1281
rect -28958 -1315 -28924 -1281
rect -28870 -1315 -28836 -1281
rect -28189 -1310 -28155 -1276
rect -28115 -1310 -28081 -1276
rect -28041 -1310 -28007 -1276
rect -27967 -1310 -27933 -1276
rect -27893 -1310 -27859 -1276
rect -27819 -1310 -27785 -1276
rect -27745 -1310 -27711 -1276
rect -27671 -1310 -27637 -1276
rect -27597 -1310 -27563 -1276
rect -27523 -1310 -27489 -1276
rect -27449 -1310 -27415 -1276
rect -27375 -1310 -27341 -1276
rect -27301 -1310 -27267 -1276
rect -27227 -1310 -27193 -1276
rect -27153 -1310 -27119 -1276
rect -29134 -1358 -29100 -1353
rect -29134 -1387 -29114 -1358
rect -29114 -1387 -29100 -1358
rect -29046 -1387 -29012 -1353
rect -28958 -1387 -28924 -1353
rect -28870 -1387 -28836 -1353
rect -28189 -1382 -28155 -1348
rect -28115 -1382 -28081 -1348
rect -28041 -1382 -28007 -1348
rect -27967 -1382 -27933 -1348
rect -27893 -1382 -27859 -1348
rect -27819 -1382 -27785 -1348
rect -27745 -1382 -27711 -1348
rect -27671 -1382 -27637 -1348
rect -27597 -1382 -27563 -1348
rect -27523 -1382 -27489 -1348
rect -27449 -1382 -27415 -1348
rect -27375 -1382 -27341 -1348
rect -27301 -1382 -27267 -1348
rect -27227 -1382 -27193 -1348
rect -27153 -1382 -27119 -1348
rect -29134 -1426 -29100 -1425
rect -29134 -1459 -29114 -1426
rect -29114 -1459 -29100 -1426
rect -29046 -1459 -29012 -1425
rect -28958 -1459 -28924 -1425
rect -28870 -1459 -28836 -1425
rect -28189 -1454 -28155 -1420
rect -28115 -1454 -28081 -1420
rect -28041 -1454 -28007 -1420
rect -27967 -1454 -27933 -1420
rect -27893 -1454 -27859 -1420
rect -27819 -1454 -27785 -1420
rect -27745 -1454 -27711 -1420
rect -27671 -1454 -27637 -1420
rect -27597 -1454 -27563 -1420
rect -27523 -1454 -27489 -1420
rect -27449 -1454 -27415 -1420
rect -27375 -1454 -27341 -1420
rect -27301 -1454 -27267 -1420
rect -27227 -1454 -27193 -1420
rect -27153 -1454 -27119 -1420
rect -29134 -1528 -29114 -1497
rect -29114 -1528 -29100 -1497
rect -29134 -1531 -29100 -1528
rect -29046 -1531 -29012 -1497
rect -28958 -1531 -28924 -1497
rect -28870 -1531 -28836 -1497
rect -28189 -1526 -28155 -1492
rect -28115 -1526 -28081 -1492
rect -28041 -1526 -28007 -1492
rect -27967 -1526 -27933 -1492
rect -27893 -1526 -27859 -1492
rect -27819 -1526 -27785 -1492
rect -27745 -1526 -27711 -1492
rect -27671 -1526 -27637 -1492
rect -27597 -1526 -27563 -1492
rect -27523 -1526 -27489 -1492
rect -27449 -1526 -27415 -1492
rect -27375 -1526 -27341 -1492
rect -27301 -1526 -27267 -1492
rect -27227 -1526 -27193 -1492
rect -27153 -1526 -27119 -1492
rect -29134 -1596 -29114 -1569
rect -29114 -1596 -29100 -1569
rect -29134 -1603 -29100 -1596
rect -29046 -1603 -29012 -1569
rect -28958 -1603 -28924 -1569
rect -28870 -1603 -28836 -1569
rect -28189 -1598 -28155 -1564
rect -28115 -1598 -28081 -1564
rect -28041 -1598 -28007 -1564
rect -27967 -1598 -27933 -1564
rect -27893 -1598 -27859 -1564
rect -27819 -1598 -27785 -1564
rect -27745 -1598 -27711 -1564
rect -27671 -1598 -27637 -1564
rect -27597 -1598 -27563 -1564
rect -27523 -1598 -27489 -1564
rect -27449 -1598 -27415 -1564
rect -27375 -1598 -27341 -1564
rect -27301 -1598 -27267 -1564
rect -27227 -1598 -27193 -1564
rect -27153 -1598 -27119 -1564
rect -29134 -1664 -29114 -1641
rect -29114 -1664 -29100 -1641
rect -29134 -1675 -29100 -1664
rect -29046 -1675 -29012 -1641
rect -28958 -1675 -28924 -1641
rect -28870 -1675 -28836 -1641
rect -28189 -1670 -28155 -1636
rect -28115 -1670 -28081 -1636
rect -28041 -1670 -28007 -1636
rect -27967 -1670 -27933 -1636
rect -27893 -1670 -27859 -1636
rect -27819 -1670 -27785 -1636
rect -27745 -1670 -27711 -1636
rect -27671 -1670 -27637 -1636
rect -27597 -1670 -27563 -1636
rect -27523 -1670 -27489 -1636
rect -27449 -1670 -27415 -1636
rect -27375 -1670 -27341 -1636
rect -27301 -1670 -27267 -1636
rect -27227 -1670 -27193 -1636
rect -27153 -1670 -27119 -1636
rect -29134 -1732 -29114 -1713
rect -29114 -1732 -29100 -1713
rect -29134 -1747 -29100 -1732
rect -29046 -1747 -29012 -1713
rect -28958 -1747 -28924 -1713
rect -28870 -1747 -28836 -1713
rect -28189 -1742 -28155 -1708
rect -28115 -1742 -28081 -1708
rect -28041 -1742 -28007 -1708
rect -27967 -1742 -27933 -1708
rect -27893 -1742 -27859 -1708
rect -27819 -1742 -27785 -1708
rect -27745 -1742 -27711 -1708
rect -27671 -1742 -27637 -1708
rect -27597 -1742 -27563 -1708
rect -27523 -1742 -27489 -1708
rect -27449 -1742 -27415 -1708
rect -27375 -1742 -27341 -1708
rect -27301 -1742 -27267 -1708
rect -27227 -1742 -27193 -1708
rect -27153 -1742 -27119 -1708
rect -29134 -1800 -29114 -1785
rect -29114 -1800 -29100 -1785
rect -29134 -1819 -29100 -1800
rect -29046 -1819 -29012 -1785
rect -28958 -1819 -28924 -1785
rect -28870 -1819 -28836 -1785
rect -28189 -1814 -28155 -1780
rect -28115 -1814 -28081 -1780
rect -28041 -1814 -28007 -1780
rect -27967 -1814 -27933 -1780
rect -27893 -1814 -27859 -1780
rect -27819 -1814 -27785 -1780
rect -27745 -1814 -27711 -1780
rect -27671 -1814 -27637 -1780
rect -27597 -1814 -27563 -1780
rect -27523 -1814 -27489 -1780
rect -27449 -1814 -27415 -1780
rect -27375 -1814 -27341 -1780
rect -27301 -1814 -27267 -1780
rect -27227 -1814 -27193 -1780
rect -27153 -1814 -27119 -1780
rect -29134 -1868 -29114 -1857
rect -29114 -1868 -29100 -1857
rect -29134 -1891 -29100 -1868
rect -29046 -1891 -29012 -1857
rect -28958 -1891 -28924 -1857
rect -28870 -1891 -28836 -1857
rect -28189 -1886 -28155 -1852
rect -28115 -1886 -28081 -1852
rect -28041 -1886 -28007 -1852
rect -27967 -1886 -27933 -1852
rect -27893 -1886 -27859 -1852
rect -27819 -1886 -27785 -1852
rect -27745 -1886 -27711 -1852
rect -27671 -1886 -27637 -1852
rect -27597 -1886 -27563 -1852
rect -27523 -1886 -27489 -1852
rect -27449 -1886 -27415 -1852
rect -27375 -1886 -27341 -1852
rect -27301 -1886 -27267 -1852
rect -27227 -1886 -27193 -1852
rect -27153 -1886 -27119 -1852
rect -29134 -1936 -29114 -1929
rect -29114 -1936 -29100 -1929
rect -29134 -1963 -29100 -1936
rect -29046 -1963 -29012 -1929
rect -28958 -1963 -28924 -1929
rect -28870 -1963 -28836 -1929
rect -28189 -1958 -28155 -1924
rect -28115 -1958 -28081 -1924
rect -28041 -1958 -28007 -1924
rect -27967 -1958 -27933 -1924
rect -27893 -1958 -27859 -1924
rect -27819 -1958 -27785 -1924
rect -27745 -1958 -27711 -1924
rect -27671 -1958 -27637 -1924
rect -27597 -1958 -27563 -1924
rect -27523 -1958 -27489 -1924
rect -27449 -1958 -27415 -1924
rect -27375 -1958 -27341 -1924
rect -27301 -1958 -27267 -1924
rect -27227 -1958 -27193 -1924
rect -27153 -1958 -27119 -1924
rect -29134 -2004 -29114 -2001
rect -29114 -2004 -29100 -2001
rect -29134 -2035 -29100 -2004
rect -29046 -2035 -29012 -2001
rect -28958 -2035 -28924 -2001
rect -28870 -2035 -28836 -2001
rect -28189 -2030 -28155 -1996
rect -28115 -2030 -28081 -1996
rect -28041 -2030 -28007 -1996
rect -27967 -2030 -27933 -1996
rect -27893 -2030 -27859 -1996
rect -27819 -2030 -27785 -1996
rect -27745 -2030 -27711 -1996
rect -27671 -2030 -27637 -1996
rect -27597 -2030 -27563 -1996
rect -27523 -2030 -27489 -1996
rect -27449 -2030 -27415 -1996
rect -27375 -2030 -27341 -1996
rect -27301 -2030 -27267 -1996
rect -27227 -2030 -27193 -1996
rect -27153 -2030 -27119 -1996
rect -29134 -2106 -29100 -2073
rect -29134 -2107 -29114 -2106
rect -29114 -2107 -29100 -2106
rect -29046 -2107 -29012 -2073
rect -28958 -2107 -28924 -2073
rect -28870 -2107 -28836 -2073
rect -28189 -2102 -28155 -2068
rect -28115 -2102 -28081 -2068
rect -28041 -2102 -28007 -2068
rect -27967 -2102 -27933 -2068
rect -27893 -2102 -27859 -2068
rect -27819 -2102 -27785 -2068
rect -27745 -2102 -27711 -2068
rect -27671 -2102 -27637 -2068
rect -27597 -2102 -27563 -2068
rect -27523 -2102 -27489 -2068
rect -27449 -2102 -27415 -2068
rect -27375 -2102 -27341 -2068
rect -27301 -2102 -27267 -2068
rect -27227 -2102 -27193 -2068
rect -27153 -2102 -27119 -2068
rect -29134 -2174 -29100 -2145
rect -29134 -2179 -29114 -2174
rect -29114 -2179 -29100 -2174
rect -29046 -2179 -29012 -2145
rect -28958 -2179 -28924 -2145
rect -28870 -2179 -28836 -2145
rect -28189 -2174 -28155 -2140
rect -28115 -2174 -28081 -2140
rect -28041 -2174 -28007 -2140
rect -27967 -2174 -27933 -2140
rect -27893 -2174 -27859 -2140
rect -27819 -2174 -27785 -2140
rect -27745 -2174 -27711 -2140
rect -27671 -2174 -27637 -2140
rect -27597 -2174 -27563 -2140
rect -27523 -2174 -27489 -2140
rect -27449 -2174 -27415 -2140
rect -27375 -2174 -27341 -2140
rect -27301 -2174 -27267 -2140
rect -27227 -2174 -27193 -2140
rect -27153 -2174 -27119 -2140
rect -29134 -2242 -29100 -2217
rect -29134 -2251 -29114 -2242
rect -29114 -2251 -29100 -2242
rect -29046 -2251 -29012 -2217
rect -28958 -2251 -28924 -2217
rect -28870 -2251 -28836 -2217
rect -28189 -2246 -28155 -2212
rect -28115 -2246 -28081 -2212
rect -28041 -2246 -28007 -2212
rect -27967 -2246 -27933 -2212
rect -27893 -2246 -27859 -2212
rect -27819 -2246 -27785 -2212
rect -27745 -2246 -27711 -2212
rect -27671 -2246 -27637 -2212
rect -27597 -2246 -27563 -2212
rect -27523 -2246 -27489 -2212
rect -27449 -2246 -27415 -2212
rect -27375 -2246 -27341 -2212
rect -27301 -2246 -27267 -2212
rect -27227 -2246 -27193 -2212
rect -27153 -2246 -27119 -2212
rect -29134 -2310 -29100 -2289
rect -29134 -2323 -29114 -2310
rect -29114 -2323 -29100 -2310
rect -29046 -2323 -29012 -2289
rect -28958 -2323 -28924 -2289
rect -28870 -2323 -28836 -2289
rect -28189 -2318 -28155 -2284
rect -28115 -2318 -28081 -2284
rect -28041 -2318 -28007 -2284
rect -27967 -2318 -27933 -2284
rect -27893 -2318 -27859 -2284
rect -27819 -2318 -27785 -2284
rect -27745 -2318 -27711 -2284
rect -27671 -2318 -27637 -2284
rect -27597 -2318 -27563 -2284
rect -27523 -2318 -27489 -2284
rect -27449 -2318 -27415 -2284
rect -27375 -2318 -27341 -2284
rect -27301 -2318 -27267 -2284
rect -27227 -2318 -27193 -2284
rect -27153 -2318 -27119 -2284
rect -29134 -2378 -29100 -2361
rect -29134 -2395 -29114 -2378
rect -29114 -2395 -29100 -2378
rect -29046 -2395 -29012 -2361
rect -28958 -2395 -28924 -2361
rect -28870 -2395 -28836 -2361
rect -28189 -2390 -28155 -2356
rect -28115 -2390 -28081 -2356
rect -28041 -2390 -28007 -2356
rect -27967 -2390 -27933 -2356
rect -27893 -2390 -27859 -2356
rect -27819 -2390 -27785 -2356
rect -27745 -2390 -27711 -2356
rect -27671 -2390 -27637 -2356
rect -27597 -2390 -27563 -2356
rect -27523 -2390 -27489 -2356
rect -27449 -2390 -27415 -2356
rect -27375 -2390 -27341 -2356
rect -27301 -2390 -27267 -2356
rect -27227 -2390 -27193 -2356
rect -27153 -2390 -27119 -2356
rect -29134 -2446 -29100 -2433
rect -29134 -2467 -29114 -2446
rect -29114 -2467 -29100 -2446
rect -29046 -2467 -29012 -2433
rect -28958 -2467 -28924 -2433
rect -28870 -2467 -28836 -2433
rect -28189 -2462 -28155 -2428
rect -28115 -2462 -28081 -2428
rect -28041 -2462 -28007 -2428
rect -27967 -2462 -27933 -2428
rect -27893 -2462 -27859 -2428
rect -27819 -2462 -27785 -2428
rect -27745 -2462 -27711 -2428
rect -27671 -2462 -27637 -2428
rect -27597 -2462 -27563 -2428
rect -27523 -2462 -27489 -2428
rect -27449 -2462 -27415 -2428
rect -27375 -2462 -27341 -2428
rect -27301 -2462 -27267 -2428
rect -27227 -2462 -27193 -2428
rect -27153 -2462 -27119 -2428
rect -29134 -2514 -29100 -2505
rect -29134 -2539 -29114 -2514
rect -29114 -2539 -29100 -2514
rect -29046 -2539 -29012 -2505
rect -28958 -2539 -28924 -2505
rect -28870 -2539 -28836 -2505
rect -28189 -2534 -28155 -2500
rect -28115 -2534 -28081 -2500
rect -28041 -2534 -28007 -2500
rect -27967 -2534 -27933 -2500
rect -27893 -2534 -27859 -2500
rect -27819 -2534 -27785 -2500
rect -27745 -2534 -27711 -2500
rect -27671 -2534 -27637 -2500
rect -27597 -2534 -27563 -2500
rect -27523 -2534 -27489 -2500
rect -27449 -2534 -27415 -2500
rect -27375 -2534 -27341 -2500
rect -27301 -2534 -27267 -2500
rect -27227 -2534 -27193 -2500
rect -27153 -2534 -27119 -2500
rect -29134 -2582 -29100 -2577
rect -29134 -2611 -29114 -2582
rect -29114 -2611 -29100 -2582
rect -29046 -2611 -29012 -2577
rect -28958 -2611 -28924 -2577
rect -28870 -2611 -28836 -2577
rect -28189 -2606 -28155 -2572
rect -28115 -2606 -28081 -2572
rect -28041 -2606 -28007 -2572
rect -27967 -2606 -27933 -2572
rect -27893 -2606 -27859 -2572
rect -27819 -2606 -27785 -2572
rect -27745 -2606 -27711 -2572
rect -27671 -2606 -27637 -2572
rect -27597 -2606 -27563 -2572
rect -27523 -2606 -27489 -2572
rect -27449 -2606 -27415 -2572
rect -27375 -2606 -27341 -2572
rect -27301 -2606 -27267 -2572
rect -27227 -2606 -27193 -2572
rect -27153 -2606 -27119 -2572
rect -29134 -2650 -29100 -2649
rect -29134 -2683 -29114 -2650
rect -29114 -2683 -29100 -2650
rect -29046 -2683 -29012 -2649
rect -28958 -2683 -28924 -2649
rect -28870 -2683 -28836 -2649
rect -28189 -2678 -28155 -2644
rect -28115 -2678 -28081 -2644
rect -28041 -2678 -28007 -2644
rect -27967 -2678 -27933 -2644
rect -27893 -2678 -27859 -2644
rect -27819 -2678 -27785 -2644
rect -27745 -2678 -27711 -2644
rect -27671 -2678 -27637 -2644
rect -27597 -2678 -27563 -2644
rect -27523 -2678 -27489 -2644
rect -27449 -2678 -27415 -2644
rect -27375 -2678 -27341 -2644
rect -27301 -2678 -27267 -2644
rect -27227 -2678 -27193 -2644
rect -27153 -2678 -27119 -2644
rect -29134 -2752 -29114 -2721
rect -29114 -2752 -29100 -2721
rect -29134 -2755 -29100 -2752
rect -29046 -2755 -29012 -2721
rect -28958 -2755 -28924 -2721
rect -28870 -2755 -28836 -2721
rect -28189 -2750 -28155 -2716
rect -28115 -2750 -28081 -2716
rect -28041 -2750 -28007 -2716
rect -27967 -2750 -27933 -2716
rect -27893 -2750 -27859 -2716
rect -27819 -2750 -27785 -2716
rect -27745 -2750 -27711 -2716
rect -27671 -2750 -27637 -2716
rect -27597 -2750 -27563 -2716
rect -27523 -2750 -27489 -2716
rect -27449 -2750 -27415 -2716
rect -27375 -2750 -27341 -2716
rect -27301 -2750 -27267 -2716
rect -27227 -2750 -27193 -2716
rect -27153 -2750 -27119 -2716
rect -29134 -2820 -29114 -2793
rect -29114 -2820 -29100 -2793
rect -29134 -2827 -29100 -2820
rect -29046 -2827 -29012 -2793
rect -28958 -2827 -28924 -2793
rect -28870 -2827 -28836 -2793
rect -28189 -2822 -28155 -2788
rect -28115 -2822 -28081 -2788
rect -28041 -2822 -28007 -2788
rect -27967 -2822 -27933 -2788
rect -27893 -2822 -27859 -2788
rect -27819 -2822 -27785 -2788
rect -27745 -2822 -27711 -2788
rect -27671 -2822 -27637 -2788
rect -27597 -2822 -27563 -2788
rect -27523 -2822 -27489 -2788
rect -27449 -2822 -27415 -2788
rect -27375 -2822 -27341 -2788
rect -27301 -2822 -27267 -2788
rect -27227 -2822 -27193 -2788
rect -27153 -2822 -27119 -2788
rect -29134 -2888 -29114 -2865
rect -29114 -2888 -29100 -2865
rect -29134 -2899 -29100 -2888
rect -29046 -2899 -29012 -2865
rect -28958 -2899 -28924 -2865
rect -28870 -2899 -28836 -2865
rect -28189 -2894 -28155 -2860
rect -28115 -2894 -28081 -2860
rect -28041 -2894 -28007 -2860
rect -27967 -2894 -27933 -2860
rect -27893 -2894 -27859 -2860
rect -27819 -2894 -27785 -2860
rect -27745 -2894 -27711 -2860
rect -27671 -2894 -27637 -2860
rect -27597 -2894 -27563 -2860
rect -27523 -2894 -27489 -2860
rect -27449 -2894 -27415 -2860
rect -27375 -2894 -27341 -2860
rect -27301 -2894 -27267 -2860
rect -27227 -2894 -27193 -2860
rect -27153 -2894 -27119 -2860
rect -29134 -2956 -29114 -2937
rect -29114 -2956 -29100 -2937
rect -29134 -2971 -29100 -2956
rect -29046 -2971 -29012 -2937
rect -28958 -2971 -28924 -2937
rect -28870 -2971 -28836 -2937
rect -28189 -2966 -28155 -2932
rect -28115 -2966 -28081 -2932
rect -28041 -2966 -28007 -2932
rect -27967 -2966 -27933 -2932
rect -27893 -2966 -27859 -2932
rect -27819 -2966 -27785 -2932
rect -27745 -2966 -27711 -2932
rect -27671 -2966 -27637 -2932
rect -27597 -2966 -27563 -2932
rect -27523 -2966 -27489 -2932
rect -27449 -2966 -27415 -2932
rect -27375 -2966 -27341 -2932
rect -27301 -2966 -27267 -2932
rect -27227 -2966 -27193 -2932
rect -27153 -2966 -27119 -2932
rect -29134 -3024 -29114 -3009
rect -29114 -3024 -29100 -3009
rect -29134 -3043 -29100 -3024
rect -29046 -3043 -29012 -3009
rect -28958 -3043 -28924 -3009
rect -28870 -3043 -28836 -3009
rect -28189 -3038 -28155 -3004
rect -28115 -3038 -28081 -3004
rect -28041 -3038 -28007 -3004
rect -27967 -3038 -27933 -3004
rect -27893 -3038 -27859 -3004
rect -27819 -3038 -27785 -3004
rect -27745 -3038 -27711 -3004
rect -27671 -3038 -27637 -3004
rect -27597 -3038 -27563 -3004
rect -27523 -3038 -27489 -3004
rect -27449 -3038 -27415 -3004
rect -27375 -3038 -27341 -3004
rect -27301 -3038 -27267 -3004
rect -27227 -3038 -27193 -3004
rect -27153 -3038 -27119 -3004
rect -29134 -3092 -29114 -3081
rect -29114 -3092 -29100 -3081
rect -29134 -3115 -29100 -3092
rect -29046 -3115 -29012 -3081
rect -28958 -3115 -28924 -3081
rect -28870 -3115 -28836 -3081
rect -28189 -3110 -28155 -3076
rect -28115 -3110 -28081 -3076
rect -28041 -3110 -28007 -3076
rect -27967 -3110 -27933 -3076
rect -27893 -3110 -27859 -3076
rect -27819 -3110 -27785 -3076
rect -27745 -3110 -27711 -3076
rect -27671 -3110 -27637 -3076
rect -27597 -3110 -27563 -3076
rect -27523 -3110 -27489 -3076
rect -27449 -3110 -27415 -3076
rect -27375 -3110 -27341 -3076
rect -27301 -3110 -27267 -3076
rect -27227 -3110 -27193 -3076
rect -27153 -3110 -27119 -3076
rect -29134 -3160 -29114 -3153
rect -29114 -3160 -29100 -3153
rect -29134 -3187 -29100 -3160
rect -29046 -3187 -29012 -3153
rect -28958 -3187 -28924 -3153
rect -28870 -3187 -28836 -3153
rect -28189 -3182 -28155 -3148
rect -28115 -3182 -28081 -3148
rect -28041 -3182 -28007 -3148
rect -27967 -3182 -27933 -3148
rect -27893 -3182 -27859 -3148
rect -27819 -3182 -27785 -3148
rect -27745 -3182 -27711 -3148
rect -27671 -3182 -27637 -3148
rect -27597 -3182 -27563 -3148
rect -27523 -3182 -27489 -3148
rect -27449 -3182 -27415 -3148
rect -27375 -3182 -27341 -3148
rect -27301 -3182 -27267 -3148
rect -27227 -3182 -27193 -3148
rect -27153 -3182 -27119 -3148
rect -29134 -3228 -29114 -3225
rect -29114 -3228 -29100 -3225
rect -29134 -3259 -29100 -3228
rect -29046 -3259 -29012 -3225
rect -28958 -3259 -28924 -3225
rect -28870 -3259 -28836 -3225
rect -28189 -3254 -28155 -3220
rect -28115 -3254 -28081 -3220
rect -28041 -3254 -28007 -3220
rect -27967 -3254 -27933 -3220
rect -27893 -3254 -27859 -3220
rect -27819 -3254 -27785 -3220
rect -27745 -3254 -27711 -3220
rect -27671 -3254 -27637 -3220
rect -27597 -3254 -27563 -3220
rect -27523 -3254 -27489 -3220
rect -27449 -3254 -27415 -3220
rect -27375 -3254 -27341 -3220
rect -27301 -3254 -27267 -3220
rect -27227 -3254 -27193 -3220
rect -27153 -3254 -27119 -3220
rect -29134 -3330 -29100 -3297
rect -29134 -3331 -29114 -3330
rect -29114 -3331 -29100 -3330
rect -29046 -3331 -29012 -3297
rect -28958 -3331 -28924 -3297
rect -28870 -3331 -28836 -3297
rect -28189 -3326 -28155 -3292
rect -28115 -3326 -28081 -3292
rect -28041 -3326 -28007 -3292
rect -27967 -3326 -27933 -3292
rect -27893 -3326 -27859 -3292
rect -27819 -3326 -27785 -3292
rect -27745 -3326 -27711 -3292
rect -27671 -3326 -27637 -3292
rect -27597 -3326 -27563 -3292
rect -27523 -3326 -27489 -3292
rect -27449 -3326 -27415 -3292
rect -27375 -3326 -27341 -3292
rect -27301 -3326 -27267 -3292
rect -27227 -3326 -27193 -3292
rect -27153 -3326 -27119 -3292
rect -29134 -3398 -29100 -3369
rect -29134 -3403 -29114 -3398
rect -29114 -3403 -29100 -3398
rect -29046 -3403 -29012 -3369
rect -28958 -3403 -28924 -3369
rect -28870 -3403 -28836 -3369
rect -28189 -3398 -28155 -3364
rect -28115 -3398 -28081 -3364
rect -28041 -3398 -28007 -3364
rect -27967 -3398 -27933 -3364
rect -27893 -3398 -27859 -3364
rect -27819 -3398 -27785 -3364
rect -27745 -3398 -27711 -3364
rect -27671 -3398 -27637 -3364
rect -27597 -3398 -27563 -3364
rect -27523 -3398 -27489 -3364
rect -27449 -3398 -27415 -3364
rect -27375 -3398 -27341 -3364
rect -27301 -3398 -27267 -3364
rect -27227 -3398 -27193 -3364
rect -27153 -3398 -27119 -3364
rect -29134 -3466 -29100 -3441
rect -29134 -3475 -29114 -3466
rect -29114 -3475 -29100 -3466
rect -29046 -3475 -29012 -3441
rect -28958 -3475 -28924 -3441
rect -28870 -3475 -28836 -3441
rect -28189 -3470 -28155 -3436
rect -28115 -3470 -28081 -3436
rect -28041 -3470 -28007 -3436
rect -27967 -3470 -27933 -3436
rect -27893 -3470 -27859 -3436
rect -27819 -3470 -27785 -3436
rect -27745 -3470 -27711 -3436
rect -27671 -3470 -27637 -3436
rect -27597 -3470 -27563 -3436
rect -27523 -3470 -27489 -3436
rect -27449 -3470 -27415 -3436
rect -27375 -3470 -27341 -3436
rect -27301 -3470 -27267 -3436
rect -27227 -3470 -27193 -3436
rect -27153 -3470 -27119 -3436
rect -29134 -3534 -29100 -3513
rect -29134 -3547 -29114 -3534
rect -29114 -3547 -29100 -3534
rect -29046 -3547 -29012 -3513
rect -28958 -3547 -28924 -3513
rect -28870 -3547 -28836 -3513
rect -28189 -3542 -28155 -3508
rect -28115 -3542 -28081 -3508
rect -28041 -3542 -28007 -3508
rect -27967 -3542 -27933 -3508
rect -27893 -3542 -27859 -3508
rect -27819 -3542 -27785 -3508
rect -27745 -3542 -27711 -3508
rect -27671 -3542 -27637 -3508
rect -27597 -3542 -27563 -3508
rect -27523 -3542 -27489 -3508
rect -27449 -3542 -27415 -3508
rect -27375 -3542 -27341 -3508
rect -27301 -3542 -27267 -3508
rect -27227 -3542 -27193 -3508
rect -27153 -3542 -27119 -3508
rect -29134 -3602 -29100 -3585
rect -29134 -3619 -29114 -3602
rect -29114 -3619 -29100 -3602
rect -29046 -3619 -29012 -3585
rect -28958 -3619 -28924 -3585
rect -28870 -3619 -28836 -3585
rect -28189 -3614 -28155 -3580
rect -28115 -3614 -28081 -3580
rect -28041 -3614 -28007 -3580
rect -27967 -3614 -27933 -3580
rect -27893 -3614 -27859 -3580
rect -27819 -3614 -27785 -3580
rect -27745 -3614 -27711 -3580
rect -27671 -3614 -27637 -3580
rect -27597 -3614 -27563 -3580
rect -27523 -3614 -27489 -3580
rect -27449 -3614 -27415 -3580
rect -27375 -3614 -27341 -3580
rect -27301 -3614 -27267 -3580
rect -27227 -3614 -27193 -3580
rect -27153 -3614 -27119 -3580
rect -29134 -3670 -29100 -3657
rect -29134 -3691 -29114 -3670
rect -29114 -3691 -29100 -3670
rect -29046 -3691 -29012 -3657
rect -28958 -3691 -28924 -3657
rect -28870 -3691 -28836 -3657
rect -28189 -3686 -28155 -3652
rect -28115 -3686 -28081 -3652
rect -28041 -3686 -28007 -3652
rect -27967 -3686 -27933 -3652
rect -27893 -3686 -27859 -3652
rect -27819 -3686 -27785 -3652
rect -27745 -3686 -27711 -3652
rect -27671 -3686 -27637 -3652
rect -27597 -3686 -27563 -3652
rect -27523 -3686 -27489 -3652
rect -27449 -3686 -27415 -3652
rect -27375 -3686 -27341 -3652
rect -27301 -3686 -27267 -3652
rect -27227 -3686 -27193 -3652
rect -27153 -3686 -27119 -3652
rect -29134 -3738 -29100 -3729
rect -29134 -3763 -29114 -3738
rect -29114 -3763 -29100 -3738
rect -29046 -3763 -29012 -3729
rect -28958 -3763 -28924 -3729
rect -28870 -3763 -28836 -3729
rect -28189 -3758 -28155 -3724
rect -28115 -3758 -28081 -3724
rect -28041 -3758 -28007 -3724
rect -27967 -3758 -27933 -3724
rect -27893 -3758 -27859 -3724
rect -27819 -3758 -27785 -3724
rect -27745 -3758 -27711 -3724
rect -27671 -3758 -27637 -3724
rect -27597 -3758 -27563 -3724
rect -27523 -3758 -27489 -3724
rect -27449 -3758 -27415 -3724
rect -27375 -3758 -27341 -3724
rect -27301 -3758 -27267 -3724
rect -27227 -3758 -27193 -3724
rect -27153 -3758 -27119 -3724
rect -29134 -3806 -29100 -3801
rect -29134 -3835 -29114 -3806
rect -29114 -3835 -29100 -3806
rect -29046 -3835 -29012 -3801
rect -28958 -3835 -28924 -3801
rect -28870 -3835 -28836 -3801
rect -28189 -3830 -28155 -3796
rect -28115 -3830 -28081 -3796
rect -28041 -3830 -28007 -3796
rect -27967 -3830 -27933 -3796
rect -27893 -3830 -27859 -3796
rect -27819 -3830 -27785 -3796
rect -27745 -3830 -27711 -3796
rect -27671 -3830 -27637 -3796
rect -27597 -3830 -27563 -3796
rect -27523 -3830 -27489 -3796
rect -27449 -3830 -27415 -3796
rect -27375 -3830 -27341 -3796
rect -27301 -3830 -27267 -3796
rect -27227 -3830 -27193 -3796
rect -27153 -3830 -27119 -3796
rect -29134 -3874 -29100 -3873
rect -29134 -3907 -29114 -3874
rect -29114 -3907 -29100 -3874
rect -29046 -3907 -29012 -3873
rect -28958 -3907 -28924 -3873
rect -28870 -3907 -28836 -3873
rect -28189 -3902 -28155 -3868
rect -28115 -3902 -28081 -3868
rect -28041 -3902 -28007 -3868
rect -27967 -3902 -27933 -3868
rect -27893 -3902 -27859 -3868
rect -27819 -3902 -27785 -3868
rect -27745 -3902 -27711 -3868
rect -27671 -3902 -27637 -3868
rect -27597 -3902 -27563 -3868
rect -27523 -3902 -27489 -3868
rect -27449 -3902 -27415 -3868
rect -27375 -3902 -27341 -3868
rect -27301 -3902 -27267 -3868
rect -27227 -3902 -27193 -3868
rect -27153 -3902 -27119 -3868
rect -29134 -3976 -29114 -3945
rect -29114 -3976 -29100 -3945
rect -29134 -3979 -29100 -3976
rect -29046 -3979 -29012 -3945
rect -28958 -3979 -28924 -3945
rect -28870 -3979 -28836 -3945
rect -28189 -3974 -28155 -3940
rect -28115 -3974 -28081 -3940
rect -28041 -3974 -28007 -3940
rect -27967 -3974 -27933 -3940
rect -27893 -3974 -27859 -3940
rect -27819 -3974 -27785 -3940
rect -27745 -3974 -27711 -3940
rect -27671 -3974 -27637 -3940
rect -27597 -3974 -27563 -3940
rect -27523 -3974 -27489 -3940
rect -27449 -3974 -27415 -3940
rect -27375 -3974 -27341 -3940
rect -27301 -3974 -27267 -3940
rect -27227 -3974 -27193 -3940
rect -27153 -3974 -27119 -3940
rect -29134 -4044 -29114 -4017
rect -29114 -4044 -29100 -4017
rect -29134 -4051 -29100 -4044
rect -29046 -4051 -29012 -4017
rect -28958 -4051 -28924 -4017
rect -28870 -4051 -28836 -4017
rect -28189 -4046 -28155 -4012
rect -28115 -4046 -28081 -4012
rect -28041 -4046 -28007 -4012
rect -27967 -4046 -27933 -4012
rect -27893 -4046 -27859 -4012
rect -27819 -4046 -27785 -4012
rect -27745 -4046 -27711 -4012
rect -27671 -4046 -27637 -4012
rect -27597 -4046 -27563 -4012
rect -27523 -4046 -27489 -4012
rect -27449 -4046 -27415 -4012
rect -27375 -4046 -27341 -4012
rect -27301 -4046 -27267 -4012
rect -27227 -4046 -27193 -4012
rect -27153 -4046 -27119 -4012
rect -29134 -4112 -29114 -4089
rect -29114 -4112 -29100 -4089
rect -29134 -4123 -29100 -4112
rect -29046 -4123 -29012 -4089
rect -28958 -4123 -28924 -4089
rect -28870 -4123 -28836 -4089
rect -28189 -4118 -28155 -4084
rect -28115 -4118 -28081 -4084
rect -28041 -4118 -28007 -4084
rect -27967 -4118 -27933 -4084
rect -27893 -4118 -27859 -4084
rect -27819 -4118 -27785 -4084
rect -27745 -4118 -27711 -4084
rect -27671 -4118 -27637 -4084
rect -27597 -4118 -27563 -4084
rect -27523 -4118 -27489 -4084
rect -27449 -4118 -27415 -4084
rect -27375 -4118 -27341 -4084
rect -27301 -4118 -27267 -4084
rect -27227 -4118 -27193 -4084
rect -27153 -4118 -27119 -4084
rect -29134 -4180 -29114 -4161
rect -29114 -4180 -29100 -4161
rect -29134 -4195 -29100 -4180
rect -29046 -4195 -29012 -4161
rect -28958 -4195 -28924 -4161
rect -28870 -4195 -28836 -4161
rect -28189 -4190 -28155 -4156
rect -28115 -4190 -28081 -4156
rect -28041 -4190 -28007 -4156
rect -27967 -4190 -27933 -4156
rect -27893 -4190 -27859 -4156
rect -27819 -4190 -27785 -4156
rect -27745 -4190 -27711 -4156
rect -27671 -4190 -27637 -4156
rect -27597 -4190 -27563 -4156
rect -27523 -4190 -27489 -4156
rect -27449 -4190 -27415 -4156
rect -27375 -4190 -27341 -4156
rect -27301 -4190 -27267 -4156
rect -27227 -4190 -27193 -4156
rect -27153 -4190 -27119 -4156
rect -29134 -4248 -29114 -4233
rect -29114 -4248 -29100 -4233
rect -29134 -4267 -29100 -4248
rect -29046 -4267 -29012 -4233
rect -28958 -4267 -28924 -4233
rect -28870 -4267 -28836 -4233
rect -28189 -4262 -28155 -4228
rect -28115 -4262 -28081 -4228
rect -28041 -4262 -28007 -4228
rect -27967 -4262 -27933 -4228
rect -27893 -4262 -27859 -4228
rect -27819 -4262 -27785 -4228
rect -27745 -4262 -27711 -4228
rect -27671 -4262 -27637 -4228
rect -27597 -4262 -27563 -4228
rect -27523 -4262 -27489 -4228
rect -27449 -4262 -27415 -4228
rect -27375 -4262 -27341 -4228
rect -27301 -4262 -27267 -4228
rect -27227 -4262 -27193 -4228
rect -27153 -4262 -27119 -4228
rect -29134 -4316 -29114 -4305
rect -29114 -4316 -29100 -4305
rect -29134 -4339 -29100 -4316
rect -29046 -4339 -29012 -4305
rect -28958 -4339 -28924 -4305
rect -28870 -4339 -28836 -4305
rect -28189 -4334 -28155 -4300
rect -28115 -4334 -28081 -4300
rect -28041 -4334 -28007 -4300
rect -27967 -4334 -27933 -4300
rect -27893 -4334 -27859 -4300
rect -27819 -4334 -27785 -4300
rect -27745 -4334 -27711 -4300
rect -27671 -4334 -27637 -4300
rect -27597 -4334 -27563 -4300
rect -27523 -4334 -27489 -4300
rect -27449 -4334 -27415 -4300
rect -27375 -4334 -27341 -4300
rect -27301 -4334 -27267 -4300
rect -27227 -4334 -27193 -4300
rect -27153 -4334 -27119 -4300
rect -29134 -4384 -29114 -4377
rect -29114 -4384 -29100 -4377
rect -29134 -4411 -29100 -4384
rect -29046 -4411 -29012 -4377
rect -28958 -4411 -28924 -4377
rect -28870 -4411 -28836 -4377
rect -28189 -4406 -28155 -4372
rect -28115 -4406 -28081 -4372
rect -28041 -4406 -28007 -4372
rect -27967 -4406 -27933 -4372
rect -27893 -4406 -27859 -4372
rect -27819 -4406 -27785 -4372
rect -27745 -4406 -27711 -4372
rect -27671 -4406 -27637 -4372
rect -27597 -4406 -27563 -4372
rect -27523 -4406 -27489 -4372
rect -27449 -4406 -27415 -4372
rect -27375 -4406 -27341 -4372
rect -27301 -4406 -27267 -4372
rect -27227 -4406 -27193 -4372
rect -27153 -4406 -27119 -4372
rect -29134 -4452 -29114 -4449
rect -29114 -4452 -29100 -4449
rect -29134 -4483 -29100 -4452
rect -29046 -4483 -29012 -4449
rect -28958 -4483 -28924 -4449
rect -28870 -4483 -28836 -4449
rect -28189 -4478 -28155 -4444
rect -28115 -4478 -28081 -4444
rect -28041 -4478 -28007 -4444
rect -27967 -4478 -27933 -4444
rect -27893 -4478 -27859 -4444
rect -27819 -4478 -27785 -4444
rect -27745 -4478 -27711 -4444
rect -27671 -4478 -27637 -4444
rect -27597 -4478 -27563 -4444
rect -27523 -4478 -27489 -4444
rect -27449 -4478 -27415 -4444
rect -27375 -4478 -27341 -4444
rect -27301 -4478 -27267 -4444
rect -27227 -4478 -27193 -4444
rect -27153 -4478 -27119 -4444
rect -29134 -4554 -29100 -4521
rect -29134 -4555 -29114 -4554
rect -29114 -4555 -29100 -4554
rect -29046 -4555 -29012 -4521
rect -28958 -4555 -28924 -4521
rect -28870 -4555 -28836 -4521
rect -28189 -4550 -28155 -4516
rect -28115 -4550 -28081 -4516
rect -28041 -4550 -28007 -4516
rect -27967 -4550 -27933 -4516
rect -27893 -4550 -27859 -4516
rect -27819 -4550 -27785 -4516
rect -27745 -4550 -27711 -4516
rect -27671 -4550 -27637 -4516
rect -27597 -4550 -27563 -4516
rect -27523 -4550 -27489 -4516
rect -27449 -4550 -27415 -4516
rect -27375 -4550 -27341 -4516
rect -27301 -4550 -27267 -4516
rect -27227 -4550 -27193 -4516
rect -27153 -4550 -27119 -4516
rect -29134 -4622 -29100 -4593
rect -29134 -4627 -29114 -4622
rect -29114 -4627 -29100 -4622
rect -29046 -4627 -29012 -4593
rect -28958 -4627 -28924 -4593
rect -28870 -4627 -28836 -4593
rect -28189 -4622 -28155 -4588
rect -28115 -4622 -28081 -4588
rect -28041 -4622 -28007 -4588
rect -27967 -4622 -27933 -4588
rect -27893 -4622 -27859 -4588
rect -27819 -4622 -27785 -4588
rect -27745 -4622 -27711 -4588
rect -27671 -4622 -27637 -4588
rect -27597 -4622 -27563 -4588
rect -27523 -4622 -27489 -4588
rect -27449 -4622 -27415 -4588
rect -27375 -4622 -27341 -4588
rect -27301 -4622 -27267 -4588
rect -27227 -4622 -27193 -4588
rect -27153 -4622 -27119 -4588
rect -29134 -4690 -29100 -4665
rect -29134 -4699 -29114 -4690
rect -29114 -4699 -29100 -4690
rect -29046 -4699 -29012 -4665
rect -28958 -4699 -28924 -4665
rect -28870 -4699 -28836 -4665
rect -28189 -4694 -28155 -4660
rect -28115 -4694 -28081 -4660
rect -28041 -4694 -28007 -4660
rect -27967 -4694 -27933 -4660
rect -27893 -4694 -27859 -4660
rect -27819 -4694 -27785 -4660
rect -27745 -4694 -27711 -4660
rect -27671 -4694 -27637 -4660
rect -27597 -4694 -27563 -4660
rect -27523 -4694 -27489 -4660
rect -27449 -4694 -27415 -4660
rect -27375 -4694 -27341 -4660
rect -27301 -4694 -27267 -4660
rect -27227 -4694 -27193 -4660
rect -27153 -4694 -27119 -4660
rect -29134 -4758 -29100 -4737
rect -29134 -4771 -29114 -4758
rect -29114 -4771 -29100 -4758
rect -29046 -4771 -29012 -4737
rect -28958 -4771 -28924 -4737
rect -28870 -4771 -28836 -4737
rect -28189 -4766 -28155 -4732
rect -28115 -4766 -28081 -4732
rect -28041 -4766 -28007 -4732
rect -27967 -4766 -27933 -4732
rect -27893 -4766 -27859 -4732
rect -27819 -4766 -27785 -4732
rect -27745 -4766 -27711 -4732
rect -27671 -4766 -27637 -4732
rect -27597 -4766 -27563 -4732
rect -27523 -4766 -27489 -4732
rect -27449 -4766 -27415 -4732
rect -27375 -4766 -27341 -4732
rect -27301 -4766 -27267 -4732
rect -27227 -4766 -27193 -4732
rect -27153 -4766 -27119 -4732
rect -29134 -4826 -29100 -4809
rect -29134 -4843 -29114 -4826
rect -29114 -4843 -29100 -4826
rect -29046 -4843 -29012 -4809
rect -28958 -4843 -28924 -4809
rect -28870 -4843 -28836 -4809
rect -28189 -4838 -28155 -4804
rect -28115 -4838 -28081 -4804
rect -28041 -4838 -28007 -4804
rect -27967 -4838 -27933 -4804
rect -27893 -4838 -27859 -4804
rect -27819 -4838 -27785 -4804
rect -27745 -4838 -27711 -4804
rect -27671 -4838 -27637 -4804
rect -27597 -4838 -27563 -4804
rect -27523 -4838 -27489 -4804
rect -27449 -4838 -27415 -4804
rect -27375 -4838 -27341 -4804
rect -27301 -4838 -27267 -4804
rect -27227 -4838 -27193 -4804
rect -27153 -4838 -27119 -4804
rect -29134 -4894 -29100 -4881
rect -29134 -4915 -29114 -4894
rect -29114 -4915 -29100 -4894
rect -29046 -4915 -29012 -4881
rect -28958 -4915 -28924 -4881
rect -28870 -4915 -28836 -4881
rect -28189 -4910 -28155 -4876
rect -28115 -4910 -28081 -4876
rect -28041 -4910 -28007 -4876
rect -27967 -4910 -27933 -4876
rect -27893 -4910 -27859 -4876
rect -27819 -4910 -27785 -4876
rect -27745 -4910 -27711 -4876
rect -27671 -4910 -27637 -4876
rect -27597 -4910 -27563 -4876
rect -27523 -4910 -27489 -4876
rect -27449 -4910 -27415 -4876
rect -27375 -4910 -27341 -4876
rect -27301 -4910 -27267 -4876
rect -27227 -4910 -27193 -4876
rect -27153 -4910 -27119 -4876
rect -29134 -4962 -29100 -4953
rect -29134 -4987 -29114 -4962
rect -29114 -4987 -29100 -4962
rect -29046 -4987 -29012 -4953
rect -28958 -4987 -28924 -4953
rect -28870 -4987 -28836 -4953
rect -28189 -4982 -28155 -4948
rect -28115 -4982 -28081 -4948
rect -28041 -4982 -28007 -4948
rect -27967 -4982 -27933 -4948
rect -27893 -4982 -27859 -4948
rect -27819 -4982 -27785 -4948
rect -27745 -4982 -27711 -4948
rect -27671 -4982 -27637 -4948
rect -27597 -4982 -27563 -4948
rect -27523 -4982 -27489 -4948
rect -27449 -4982 -27415 -4948
rect -27375 -4982 -27341 -4948
rect -27301 -4982 -27267 -4948
rect -27227 -4982 -27193 -4948
rect -27153 -4982 -27119 -4948
rect -29134 -5030 -29100 -5025
rect -29134 -5059 -29114 -5030
rect -29114 -5059 -29100 -5030
rect -29046 -5059 -29012 -5025
rect -28958 -5059 -28924 -5025
rect -28870 -5059 -28836 -5025
rect -28189 -5054 -28155 -5020
rect -28115 -5054 -28081 -5020
rect -28041 -5054 -28007 -5020
rect -27967 -5054 -27933 -5020
rect -27893 -5054 -27859 -5020
rect -27819 -5054 -27785 -5020
rect -27745 -5054 -27711 -5020
rect -27671 -5054 -27637 -5020
rect -27597 -5054 -27563 -5020
rect -27523 -5054 -27489 -5020
rect -27449 -5054 -27415 -5020
rect -27375 -5054 -27341 -5020
rect -27301 -5054 -27267 -5020
rect -27227 -5054 -27193 -5020
rect -27153 -5054 -27119 -5020
rect -29134 -5098 -29100 -5097
rect -29134 -5131 -29114 -5098
rect -29114 -5131 -29100 -5098
rect -29046 -5131 -29012 -5097
rect -28958 -5131 -28924 -5097
rect -28870 -5131 -28836 -5097
rect -28189 -5126 -28155 -5092
rect -28115 -5126 -28081 -5092
rect -28041 -5126 -28007 -5092
rect -27967 -5126 -27933 -5092
rect -27893 -5126 -27859 -5092
rect -27819 -5126 -27785 -5092
rect -27745 -5126 -27711 -5092
rect -27671 -5126 -27637 -5092
rect -27597 -5126 -27563 -5092
rect -27523 -5126 -27489 -5092
rect -27449 -5126 -27415 -5092
rect -27375 -5126 -27341 -5092
rect -27301 -5126 -27267 -5092
rect -27227 -5126 -27193 -5092
rect -27153 -5126 -27119 -5092
rect -29134 -5200 -29114 -5169
rect -29114 -5200 -29100 -5169
rect -29134 -5203 -29100 -5200
rect -29046 -5203 -29012 -5169
rect -28958 -5203 -28924 -5169
rect -28870 -5203 -28836 -5169
rect -28189 -5198 -28155 -5164
rect -28115 -5198 -28081 -5164
rect -28041 -5198 -28007 -5164
rect -27967 -5198 -27933 -5164
rect -27893 -5198 -27859 -5164
rect -27819 -5198 -27785 -5164
rect -27745 -5198 -27711 -5164
rect -27671 -5198 -27637 -5164
rect -27597 -5198 -27563 -5164
rect -27523 -5198 -27489 -5164
rect -27449 -5198 -27415 -5164
rect -27375 -5198 -27341 -5164
rect -27301 -5198 -27267 -5164
rect -27227 -5198 -27193 -5164
rect -27153 -5198 -27119 -5164
rect -29134 -5268 -29114 -5241
rect -29114 -5268 -29100 -5241
rect -29134 -5275 -29100 -5268
rect -29046 -5275 -29012 -5241
rect -28958 -5275 -28924 -5241
rect -28870 -5275 -28836 -5241
rect -28189 -5270 -28155 -5236
rect -28115 -5270 -28081 -5236
rect -28041 -5270 -28007 -5236
rect -27967 -5270 -27933 -5236
rect -27893 -5270 -27859 -5236
rect -27819 -5270 -27785 -5236
rect -27745 -5270 -27711 -5236
rect -27671 -5270 -27637 -5236
rect -27597 -5270 -27563 -5236
rect -27523 -5270 -27489 -5236
rect -27449 -5270 -27415 -5236
rect -27375 -5270 -27341 -5236
rect -27301 -5270 -27267 -5236
rect -27227 -5270 -27193 -5236
rect -27153 -5270 -27119 -5236
rect -29134 -5336 -29114 -5313
rect -29114 -5336 -29100 -5313
rect -29134 -5347 -29100 -5336
rect -29046 -5347 -29012 -5313
rect -28958 -5347 -28924 -5313
rect -28870 -5347 -28836 -5313
rect -28189 -5342 -28155 -5308
rect -28115 -5342 -28081 -5308
rect -28041 -5342 -28007 -5308
rect -27967 -5342 -27933 -5308
rect -27893 -5342 -27859 -5308
rect -27819 -5342 -27785 -5308
rect -27745 -5342 -27711 -5308
rect -27671 -5342 -27637 -5308
rect -27597 -5342 -27563 -5308
rect -27523 -5342 -27489 -5308
rect -27449 -5342 -27415 -5308
rect -27375 -5342 -27341 -5308
rect -27301 -5342 -27267 -5308
rect -27227 -5342 -27193 -5308
rect -27153 -5342 -27119 -5308
rect -29134 -5404 -29114 -5385
rect -29114 -5404 -29100 -5385
rect -29134 -5419 -29100 -5404
rect -29046 -5419 -29012 -5385
rect -28958 -5419 -28924 -5385
rect -28870 -5419 -28836 -5385
rect -28189 -5414 -28155 -5380
rect -28115 -5414 -28081 -5380
rect -28041 -5414 -28007 -5380
rect -27967 -5414 -27933 -5380
rect -27893 -5414 -27859 -5380
rect -27819 -5414 -27785 -5380
rect -27745 -5414 -27711 -5380
rect -27671 -5414 -27637 -5380
rect -27597 -5414 -27563 -5380
rect -27523 -5414 -27489 -5380
rect -27449 -5414 -27415 -5380
rect -27375 -5414 -27341 -5380
rect -27301 -5414 -27267 -5380
rect -27227 -5414 -27193 -5380
rect -27153 -5414 -27119 -5380
rect -29134 -5472 -29114 -5457
rect -29114 -5472 -29100 -5457
rect -29134 -5491 -29100 -5472
rect -29046 -5491 -29012 -5457
rect -28958 -5491 -28924 -5457
rect -28870 -5491 -28836 -5457
rect -28189 -5486 -28155 -5452
rect -28115 -5486 -28081 -5452
rect -28041 -5486 -28007 -5452
rect -27967 -5486 -27933 -5452
rect -27893 -5486 -27859 -5452
rect -27819 -5486 -27785 -5452
rect -27745 -5486 -27711 -5452
rect -27671 -5486 -27637 -5452
rect -27597 -5486 -27563 -5452
rect -27523 -5486 -27489 -5452
rect -27449 -5486 -27415 -5452
rect -27375 -5486 -27341 -5452
rect -27301 -5486 -27267 -5452
rect -27227 -5486 -27193 -5452
rect -27153 -5486 -27119 -5452
rect -29134 -5540 -29114 -5529
rect -29114 -5540 -29100 -5529
rect -29134 -5563 -29100 -5540
rect -29046 -5563 -29012 -5529
rect -28958 -5563 -28924 -5529
rect -28870 -5563 -28836 -5529
rect -28189 -5558 -28155 -5524
rect -28115 -5558 -28081 -5524
rect -28041 -5558 -28007 -5524
rect -27967 -5558 -27933 -5524
rect -27893 -5558 -27859 -5524
rect -27819 -5558 -27785 -5524
rect -27745 -5558 -27711 -5524
rect -27671 -5558 -27637 -5524
rect -27597 -5558 -27563 -5524
rect -27523 -5558 -27489 -5524
rect -27449 -5558 -27415 -5524
rect -27375 -5558 -27341 -5524
rect -27301 -5558 -27267 -5524
rect -27227 -5558 -27193 -5524
rect -27153 -5558 -27119 -5524
rect -29134 -5608 -29114 -5601
rect -29114 -5608 -29100 -5601
rect -29134 -5635 -29100 -5608
rect -29046 -5635 -29012 -5601
rect -28958 -5635 -28924 -5601
rect -28870 -5635 -28836 -5601
rect -28189 -5630 -28155 -5596
rect -28115 -5630 -28081 -5596
rect -28041 -5630 -28007 -5596
rect -27967 -5630 -27933 -5596
rect -27893 -5630 -27859 -5596
rect -27819 -5630 -27785 -5596
rect -27745 -5630 -27711 -5596
rect -27671 -5630 -27637 -5596
rect -27597 -5630 -27563 -5596
rect -27523 -5630 -27489 -5596
rect -27449 -5630 -27415 -5596
rect -27375 -5630 -27341 -5596
rect -27301 -5630 -27267 -5596
rect -27227 -5630 -27193 -5596
rect -27153 -5630 -27119 -5596
rect -29134 -5676 -29114 -5673
rect -29114 -5676 -29100 -5673
rect -29134 -5707 -29100 -5676
rect -29046 -5707 -29012 -5673
rect -28958 -5707 -28924 -5673
rect -28870 -5707 -28836 -5673
rect -28189 -5702 -28155 -5668
rect -28115 -5702 -28081 -5668
rect -28041 -5702 -28007 -5668
rect -27967 -5702 -27933 -5668
rect -27893 -5702 -27859 -5668
rect -27819 -5702 -27785 -5668
rect -27745 -5702 -27711 -5668
rect -27671 -5702 -27637 -5668
rect -27597 -5702 -27563 -5668
rect -27523 -5702 -27489 -5668
rect -27449 -5702 -27415 -5668
rect -27375 -5702 -27341 -5668
rect -27301 -5702 -27267 -5668
rect -27227 -5702 -27193 -5668
rect -27153 -5702 -27119 -5668
rect -29134 -5778 -29100 -5745
rect -29134 -5779 -29114 -5778
rect -29114 -5779 -29100 -5778
rect -29046 -5779 -29012 -5745
rect -28958 -5779 -28924 -5745
rect -28870 -5779 -28836 -5745
rect -28189 -5774 -28155 -5740
rect -28115 -5774 -28081 -5740
rect -28041 -5774 -28007 -5740
rect -27967 -5774 -27933 -5740
rect -27893 -5774 -27859 -5740
rect -27819 -5774 -27785 -5740
rect -27745 -5774 -27711 -5740
rect -27671 -5774 -27637 -5740
rect -27597 -5774 -27563 -5740
rect -27523 -5774 -27489 -5740
rect -27449 -5774 -27415 -5740
rect -27375 -5774 -27341 -5740
rect -27301 -5774 -27267 -5740
rect -27227 -5774 -27193 -5740
rect -27153 -5774 -27119 -5740
rect -29134 -5846 -29100 -5817
rect -29134 -5851 -29114 -5846
rect -29114 -5851 -29100 -5846
rect -29046 -5851 -29012 -5817
rect -28958 -5851 -28924 -5817
rect -28870 -5851 -28836 -5817
rect -28189 -5846 -28155 -5812
rect -28115 -5846 -28081 -5812
rect -28041 -5846 -28007 -5812
rect -27967 -5846 -27933 -5812
rect -27893 -5846 -27859 -5812
rect -27819 -5846 -27785 -5812
rect -27745 -5846 -27711 -5812
rect -27671 -5846 -27637 -5812
rect -27597 -5846 -27563 -5812
rect -27523 -5846 -27489 -5812
rect -27449 -5846 -27415 -5812
rect -27375 -5846 -27341 -5812
rect -27301 -5846 -27267 -5812
rect -27227 -5846 -27193 -5812
rect -27153 -5846 -27119 -5812
rect -29134 -5914 -29100 -5889
rect -29134 -5923 -29114 -5914
rect -29114 -5923 -29100 -5914
rect -29046 -5923 -29012 -5889
rect -28958 -5923 -28924 -5889
rect -28870 -5923 -28836 -5889
rect -28189 -5918 -28155 -5884
rect -28115 -5918 -28081 -5884
rect -28041 -5918 -28007 -5884
rect -27967 -5918 -27933 -5884
rect -27893 -5918 -27859 -5884
rect -27819 -5918 -27785 -5884
rect -27745 -5918 -27711 -5884
rect -27671 -5918 -27637 -5884
rect -27597 -5918 -27563 -5884
rect -27523 -5918 -27489 -5884
rect -27449 -5918 -27415 -5884
rect -27375 -5918 -27341 -5884
rect -27301 -5918 -27267 -5884
rect -27227 -5918 -27193 -5884
rect -27153 -5918 -27119 -5884
rect -29134 -5982 -29100 -5961
rect -29134 -5995 -29114 -5982
rect -29114 -5995 -29100 -5982
rect -29046 -5995 -29012 -5961
rect -28958 -5995 -28924 -5961
rect -28870 -5995 -28836 -5961
rect -28189 -5990 -28155 -5956
rect -28115 -5990 -28081 -5956
rect -28041 -5990 -28007 -5956
rect -27967 -5990 -27933 -5956
rect -27893 -5990 -27859 -5956
rect -27819 -5990 -27785 -5956
rect -27745 -5990 -27711 -5956
rect -27671 -5990 -27637 -5956
rect -27597 -5990 -27563 -5956
rect -27523 -5990 -27489 -5956
rect -27449 -5990 -27415 -5956
rect -27375 -5990 -27341 -5956
rect -27301 -5990 -27267 -5956
rect -27227 -5990 -27193 -5956
rect -27153 -5990 -27119 -5956
rect -29134 -6050 -29100 -6033
rect -29134 -6067 -29114 -6050
rect -29114 -6067 -29100 -6050
rect -29046 -6067 -29012 -6033
rect -28958 -6067 -28924 -6033
rect -28870 -6067 -28836 -6033
rect -28189 -6062 -28155 -6028
rect -28115 -6062 -28081 -6028
rect -28041 -6062 -28007 -6028
rect -27967 -6062 -27933 -6028
rect -27893 -6062 -27859 -6028
rect -27819 -6062 -27785 -6028
rect -27745 -6062 -27711 -6028
rect -27671 -6062 -27637 -6028
rect -27597 -6062 -27563 -6028
rect -27523 -6062 -27489 -6028
rect -27449 -6062 -27415 -6028
rect -27375 -6062 -27341 -6028
rect -27301 -6062 -27267 -6028
rect -27227 -6062 -27193 -6028
rect -27153 -6062 -27119 -6028
rect -29134 -6118 -29100 -6105
rect -29134 -6139 -29114 -6118
rect -29114 -6139 -29100 -6118
rect -29046 -6139 -29012 -6105
rect -28958 -6139 -28924 -6105
rect -28870 -6139 -28836 -6105
rect -28189 -6134 -28155 -6100
rect -28115 -6134 -28081 -6100
rect -28041 -6134 -28007 -6100
rect -27967 -6134 -27933 -6100
rect -27893 -6134 -27859 -6100
rect -27819 -6134 -27785 -6100
rect -27745 -6134 -27711 -6100
rect -27671 -6134 -27637 -6100
rect -27597 -6134 -27563 -6100
rect -27523 -6134 -27489 -6100
rect -27449 -6134 -27415 -6100
rect -27375 -6134 -27341 -6100
rect -27301 -6134 -27267 -6100
rect -27227 -6134 -27193 -6100
rect -27153 -6134 -27119 -6100
rect -29134 -6186 -29100 -6177
rect -29134 -6211 -29114 -6186
rect -29114 -6211 -29100 -6186
rect -29046 -6211 -29012 -6177
rect -28958 -6211 -28924 -6177
rect -28870 -6211 -28836 -6177
rect -28189 -6206 -28155 -6172
rect -28115 -6206 -28081 -6172
rect -28041 -6206 -28007 -6172
rect -27967 -6206 -27933 -6172
rect -27893 -6206 -27859 -6172
rect -27819 -6206 -27785 -6172
rect -27745 -6206 -27711 -6172
rect -27671 -6206 -27637 -6172
rect -27597 -6206 -27563 -6172
rect -27523 -6206 -27489 -6172
rect -27449 -6206 -27415 -6172
rect -27375 -6206 -27341 -6172
rect -27301 -6206 -27267 -6172
rect -27227 -6206 -27193 -6172
rect -27153 -6206 -27119 -6172
rect -29134 -6254 -29100 -6249
rect -29134 -6283 -29114 -6254
rect -29114 -6283 -29100 -6254
rect -29046 -6283 -29012 -6249
rect -28958 -6283 -28924 -6249
rect -28870 -6283 -28836 -6249
rect -28189 -6278 -28155 -6244
rect -28115 -6278 -28081 -6244
rect -28041 -6278 -28007 -6244
rect -27967 -6278 -27933 -6244
rect -27893 -6278 -27859 -6244
rect -27819 -6278 -27785 -6244
rect -27745 -6278 -27711 -6244
rect -27671 -6278 -27637 -6244
rect -27597 -6278 -27563 -6244
rect -27523 -6278 -27489 -6244
rect -27449 -6278 -27415 -6244
rect -27375 -6278 -27341 -6244
rect -27301 -6278 -27267 -6244
rect -27227 -6278 -27193 -6244
rect -27153 -6278 -27119 -6244
rect -29134 -6322 -29100 -6321
rect -29134 -6355 -29114 -6322
rect -29114 -6355 -29100 -6322
rect -29046 -6355 -29012 -6321
rect -28958 -6355 -28924 -6321
rect -28870 -6355 -28836 -6321
rect -28189 -6350 -28155 -6316
rect -28115 -6350 -28081 -6316
rect -28041 -6350 -28007 -6316
rect -27967 -6350 -27933 -6316
rect -27893 -6350 -27859 -6316
rect -27819 -6350 -27785 -6316
rect -27745 -6350 -27711 -6316
rect -27671 -6350 -27637 -6316
rect -27597 -6350 -27563 -6316
rect -27523 -6350 -27489 -6316
rect -27449 -6350 -27415 -6316
rect -27375 -6350 -27341 -6316
rect -27301 -6350 -27267 -6316
rect -27227 -6350 -27193 -6316
rect -27153 -6350 -27119 -6316
rect -29134 -6424 -29114 -6393
rect -29114 -6424 -29100 -6393
rect -29134 -6427 -29100 -6424
rect -29046 -6427 -29012 -6393
rect -28958 -6427 -28924 -6393
rect -28870 -6427 -28836 -6393
rect -28189 -6422 -28155 -6388
rect -28115 -6422 -28081 -6388
rect -28041 -6422 -28007 -6388
rect -27967 -6422 -27933 -6388
rect -27893 -6422 -27859 -6388
rect -27819 -6422 -27785 -6388
rect -27745 -6422 -27711 -6388
rect -27671 -6422 -27637 -6388
rect -27597 -6422 -27563 -6388
rect -27523 -6422 -27489 -6388
rect -27449 -6422 -27415 -6388
rect -27375 -6422 -27341 -6388
rect -27301 -6422 -27267 -6388
rect -27227 -6422 -27193 -6388
rect -27153 -6422 -27119 -6388
rect -29134 -6492 -29114 -6465
rect -29114 -6492 -29100 -6465
rect -29134 -6499 -29100 -6492
rect -29046 -6499 -29012 -6465
rect -28958 -6499 -28924 -6465
rect -28870 -6499 -28836 -6465
rect -28189 -6494 -28155 -6460
rect -28115 -6494 -28081 -6460
rect -28041 -6494 -28007 -6460
rect -27967 -6494 -27933 -6460
rect -27893 -6494 -27859 -6460
rect -27819 -6494 -27785 -6460
rect -27745 -6494 -27711 -6460
rect -27671 -6494 -27637 -6460
rect -27597 -6494 -27563 -6460
rect -27523 -6494 -27489 -6460
rect -27449 -6494 -27415 -6460
rect -27375 -6494 -27341 -6460
rect -27301 -6494 -27267 -6460
rect -27227 -6494 -27193 -6460
rect -27153 -6494 -27119 -6460
rect -29134 -6560 -29114 -6537
rect -29114 -6560 -29100 -6537
rect -29134 -6571 -29100 -6560
rect -29046 -6571 -29012 -6537
rect -28958 -6571 -28924 -6537
rect -28870 -6571 -28836 -6537
rect -28189 -6566 -28155 -6532
rect -28115 -6566 -28081 -6532
rect -28041 -6566 -28007 -6532
rect -27967 -6566 -27933 -6532
rect -27893 -6566 -27859 -6532
rect -27819 -6566 -27785 -6532
rect -27745 -6566 -27711 -6532
rect -27671 -6566 -27637 -6532
rect -27597 -6566 -27563 -6532
rect -27523 -6566 -27489 -6532
rect -27449 -6566 -27415 -6532
rect -27375 -6566 -27341 -6532
rect -27301 -6566 -27267 -6532
rect -27227 -6566 -27193 -6532
rect -27153 -6566 -27119 -6532
rect -29134 -6628 -29114 -6609
rect -29114 -6628 -29100 -6609
rect -29134 -6643 -29100 -6628
rect -29046 -6643 -29012 -6609
rect -28958 -6643 -28924 -6609
rect -28870 -6643 -28836 -6609
rect -28189 -6638 -28155 -6604
rect -28115 -6638 -28081 -6604
rect -28041 -6638 -28007 -6604
rect -27967 -6638 -27933 -6604
rect -27893 -6638 -27859 -6604
rect -27819 -6638 -27785 -6604
rect -27745 -6638 -27711 -6604
rect -27671 -6638 -27637 -6604
rect -27597 -6638 -27563 -6604
rect -27523 -6638 -27489 -6604
rect -27449 -6638 -27415 -6604
rect -27375 -6638 -27341 -6604
rect -27301 -6638 -27267 -6604
rect -27227 -6638 -27193 -6604
rect -27153 -6638 -27119 -6604
rect -29134 -6696 -29114 -6681
rect -29114 -6696 -29100 -6681
rect -29134 -6715 -29100 -6696
rect -29046 -6715 -29012 -6681
rect -28958 -6715 -28924 -6681
rect -28870 -6715 -28836 -6681
rect -28189 -6710 -28155 -6676
rect -28115 -6710 -28081 -6676
rect -28041 -6710 -28007 -6676
rect -27967 -6710 -27933 -6676
rect -27893 -6710 -27859 -6676
rect -27819 -6710 -27785 -6676
rect -27745 -6710 -27711 -6676
rect -27671 -6710 -27637 -6676
rect -27597 -6710 -27563 -6676
rect -27523 -6710 -27489 -6676
rect -27449 -6710 -27415 -6676
rect -27375 -6710 -27341 -6676
rect -27301 -6710 -27267 -6676
rect -27227 -6710 -27193 -6676
rect -27153 -6710 -27119 -6676
rect -29134 -6764 -29114 -6753
rect -29114 -6764 -29100 -6753
rect -29134 -6787 -29100 -6764
rect -29046 -6787 -29012 -6753
rect -28958 -6787 -28924 -6753
rect -28870 -6787 -28836 -6753
rect -28189 -6782 -28155 -6748
rect -28115 -6782 -28081 -6748
rect -28041 -6782 -28007 -6748
rect -27967 -6782 -27933 -6748
rect -27893 -6782 -27859 -6748
rect -27819 -6782 -27785 -6748
rect -27745 -6782 -27711 -6748
rect -27671 -6782 -27637 -6748
rect -27597 -6782 -27563 -6748
rect -27523 -6782 -27489 -6748
rect -27449 -6782 -27415 -6748
rect -27375 -6782 -27341 -6748
rect -27301 -6782 -27267 -6748
rect -27227 -6782 -27193 -6748
rect -27153 -6782 -27119 -6748
rect -29134 -6832 -29114 -6825
rect -29114 -6832 -29100 -6825
rect -29134 -6859 -29100 -6832
rect -29046 -6859 -29012 -6825
rect -28958 -6859 -28924 -6825
rect -28870 -6859 -28836 -6825
rect -28189 -6854 -28155 -6820
rect -28115 -6854 -28081 -6820
rect -28041 -6854 -28007 -6820
rect -27967 -6854 -27933 -6820
rect -27893 -6854 -27859 -6820
rect -27819 -6854 -27785 -6820
rect -27745 -6854 -27711 -6820
rect -27671 -6854 -27637 -6820
rect -27597 -6854 -27563 -6820
rect -27523 -6854 -27489 -6820
rect -27449 -6854 -27415 -6820
rect -27375 -6854 -27341 -6820
rect -27301 -6854 -27267 -6820
rect -27227 -6854 -27193 -6820
rect -27153 -6854 -27119 -6820
rect -29134 -6900 -29114 -6897
rect -29114 -6900 -29100 -6897
rect -29134 -6931 -29100 -6900
rect -29046 -6931 -29012 -6897
rect -28958 -6931 -28924 -6897
rect -28870 -6931 -28836 -6897
rect -28189 -6926 -28155 -6892
rect -28115 -6926 -28081 -6892
rect -28041 -6926 -28007 -6892
rect -27967 -6926 -27933 -6892
rect -27893 -6926 -27859 -6892
rect -27819 -6926 -27785 -6892
rect -27745 -6926 -27711 -6892
rect -27671 -6926 -27637 -6892
rect -27597 -6926 -27563 -6892
rect -27523 -6926 -27489 -6892
rect -27449 -6926 -27415 -6892
rect -27375 -6926 -27341 -6892
rect -27301 -6926 -27267 -6892
rect -27227 -6926 -27193 -6892
rect -27153 -6926 -27119 -6892
rect -29134 -7002 -29100 -6969
rect -29134 -7003 -29114 -7002
rect -29114 -7003 -29100 -7002
rect -29046 -7003 -29012 -6969
rect -28958 -7003 -28924 -6969
rect -28870 -7003 -28836 -6969
rect -28189 -6998 -28155 -6964
rect -28115 -6998 -28081 -6964
rect -28041 -6998 -28007 -6964
rect -27967 -6998 -27933 -6964
rect -27893 -6998 -27859 -6964
rect -27819 -6998 -27785 -6964
rect -27745 -6998 -27711 -6964
rect -27671 -6998 -27637 -6964
rect -27597 -6998 -27563 -6964
rect -27523 -6998 -27489 -6964
rect -27449 -6998 -27415 -6964
rect -27375 -6998 -27341 -6964
rect -27301 -6998 -27267 -6964
rect -27227 -6998 -27193 -6964
rect -27153 -6998 -27119 -6964
rect -29134 -7070 -29100 -7041
rect -29134 -7075 -29114 -7070
rect -29114 -7075 -29100 -7070
rect -29046 -7075 -29012 -7041
rect -28958 -7075 -28924 -7041
rect -28870 -7075 -28836 -7041
rect -28189 -7070 -28155 -7036
rect -28115 -7070 -28081 -7036
rect -28041 -7070 -28007 -7036
rect -27967 -7070 -27933 -7036
rect -27893 -7070 -27859 -7036
rect -27819 -7070 -27785 -7036
rect -27745 -7070 -27711 -7036
rect -27671 -7070 -27637 -7036
rect -27597 -7070 -27563 -7036
rect -27523 -7070 -27489 -7036
rect -27449 -7070 -27415 -7036
rect -27375 -7070 -27341 -7036
rect -27301 -7070 -27267 -7036
rect -27227 -7070 -27193 -7036
rect -27153 -7070 -27119 -7036
rect -29134 -7138 -29100 -7113
rect -29134 -7147 -29114 -7138
rect -29114 -7147 -29100 -7138
rect -29046 -7147 -29012 -7113
rect -28958 -7147 -28924 -7113
rect -28870 -7147 -28836 -7113
rect -28189 -7142 -28155 -7108
rect -28115 -7142 -28081 -7108
rect -28041 -7142 -28007 -7108
rect -27967 -7142 -27933 -7108
rect -27893 -7142 -27859 -7108
rect -27819 -7142 -27785 -7108
rect -27745 -7142 -27711 -7108
rect -27671 -7142 -27637 -7108
rect -27597 -7142 -27563 -7108
rect -27523 -7142 -27489 -7108
rect -27449 -7142 -27415 -7108
rect -27375 -7142 -27341 -7108
rect -27301 -7142 -27267 -7108
rect -27227 -7142 -27193 -7108
rect -27153 -7142 -27119 -7108
rect -29134 -7206 -29100 -7185
rect -29134 -7219 -29114 -7206
rect -29114 -7219 -29100 -7206
rect -29046 -7219 -29012 -7185
rect -28958 -7219 -28924 -7185
rect -28870 -7219 -28836 -7185
rect -28189 -7214 -28155 -7180
rect -28115 -7214 -28081 -7180
rect -28041 -7214 -28007 -7180
rect -27967 -7214 -27933 -7180
rect -27893 -7214 -27859 -7180
rect -27819 -7214 -27785 -7180
rect -27745 -7214 -27711 -7180
rect -27671 -7214 -27637 -7180
rect -27597 -7214 -27563 -7180
rect -27523 -7214 -27489 -7180
rect -27449 -7214 -27415 -7180
rect -27375 -7214 -27341 -7180
rect -27301 -7214 -27267 -7180
rect -27227 -7214 -27193 -7180
rect -27153 -7214 -27119 -7180
rect -29134 -7274 -29100 -7257
rect -29134 -7291 -29114 -7274
rect -29114 -7291 -29100 -7274
rect -29046 -7291 -29012 -7257
rect -28958 -7291 -28924 -7257
rect -28870 -7291 -28836 -7257
rect -28189 -7286 -28155 -7252
rect -28115 -7286 -28081 -7252
rect -28041 -7286 -28007 -7252
rect -27967 -7286 -27933 -7252
rect -27893 -7286 -27859 -7252
rect -27819 -7286 -27785 -7252
rect -27745 -7286 -27711 -7252
rect -27671 -7286 -27637 -7252
rect -27597 -7286 -27563 -7252
rect -27523 -7286 -27489 -7252
rect -27449 -7286 -27415 -7252
rect -27375 -7286 -27341 -7252
rect -27301 -7286 -27267 -7252
rect -27227 -7286 -27193 -7252
rect -27153 -7286 -27119 -7252
rect -29134 -7342 -29100 -7329
rect -29134 -7363 -29114 -7342
rect -29114 -7363 -29100 -7342
rect -29046 -7363 -29012 -7329
rect -28958 -7363 -28924 -7329
rect -28870 -7363 -28836 -7329
rect -28189 -7358 -28155 -7324
rect -28115 -7358 -28081 -7324
rect -28041 -7358 -28007 -7324
rect -27967 -7358 -27933 -7324
rect -27893 -7358 -27859 -7324
rect -27819 -7358 -27785 -7324
rect -27745 -7358 -27711 -7324
rect -27671 -7358 -27637 -7324
rect -27597 -7358 -27563 -7324
rect -27523 -7358 -27489 -7324
rect -27449 -7358 -27415 -7324
rect -27375 -7358 -27341 -7324
rect -27301 -7358 -27267 -7324
rect -27227 -7358 -27193 -7324
rect -27153 -7358 -27119 -7324
rect -29134 -7410 -29100 -7401
rect -29134 -7435 -29114 -7410
rect -29114 -7435 -29100 -7410
rect -29046 -7435 -29012 -7401
rect -28958 -7435 -28924 -7401
rect -28870 -7435 -28836 -7401
rect -28189 -7430 -28155 -7396
rect -28115 -7430 -28081 -7396
rect -28041 -7430 -28007 -7396
rect -27967 -7430 -27933 -7396
rect -27893 -7430 -27859 -7396
rect -27819 -7430 -27785 -7396
rect -27745 -7430 -27711 -7396
rect -27671 -7430 -27637 -7396
rect -27597 -7430 -27563 -7396
rect -27523 -7430 -27489 -7396
rect -27449 -7430 -27415 -7396
rect -27375 -7430 -27341 -7396
rect -27301 -7430 -27267 -7396
rect -27227 -7430 -27193 -7396
rect -27153 -7430 -27119 -7396
rect -29134 -7478 -29100 -7473
rect -29134 -7507 -29114 -7478
rect -29114 -7507 -29100 -7478
rect -29046 -7507 -29012 -7473
rect -28958 -7507 -28924 -7473
rect -28870 -7507 -28836 -7473
rect -28189 -7502 -28155 -7468
rect -28115 -7502 -28081 -7468
rect -28041 -7502 -28007 -7468
rect -27967 -7502 -27933 -7468
rect -27893 -7502 -27859 -7468
rect -27819 -7502 -27785 -7468
rect -27745 -7502 -27711 -7468
rect -27671 -7502 -27637 -7468
rect -27597 -7502 -27563 -7468
rect -27523 -7502 -27489 -7468
rect -27449 -7502 -27415 -7468
rect -27375 -7502 -27341 -7468
rect -27301 -7502 -27267 -7468
rect -27227 -7502 -27193 -7468
rect -27153 -7502 -27119 -7468
rect -29134 -7546 -29100 -7545
rect -29134 -7579 -29114 -7546
rect -29114 -7579 -29100 -7546
rect -29046 -7579 -29012 -7545
rect -28958 -7579 -28924 -7545
rect -28870 -7579 -28836 -7545
rect -28189 -7574 -28155 -7540
rect -28115 -7574 -28081 -7540
rect -28041 -7574 -28007 -7540
rect -27967 -7574 -27933 -7540
rect -27893 -7574 -27859 -7540
rect -27819 -7574 -27785 -7540
rect -27745 -7574 -27711 -7540
rect -27671 -7574 -27637 -7540
rect -27597 -7574 -27563 -7540
rect -27523 -7574 -27489 -7540
rect -27449 -7574 -27415 -7540
rect -27375 -7574 -27341 -7540
rect -27301 -7574 -27267 -7540
rect -27227 -7574 -27193 -7540
rect -27153 -7574 -27119 -7540
rect -29134 -7648 -29114 -7617
rect -29114 -7648 -29100 -7617
rect -29134 -7651 -29100 -7648
rect -29046 -7651 -29012 -7617
rect -28958 -7651 -28924 -7617
rect -28870 -7651 -28836 -7617
rect -28189 -7646 -28155 -7612
rect -28115 -7646 -28081 -7612
rect -28041 -7646 -28007 -7612
rect -27967 -7646 -27933 -7612
rect -27893 -7646 -27859 -7612
rect -27819 -7646 -27785 -7612
rect -27745 -7646 -27711 -7612
rect -27671 -7646 -27637 -7612
rect -27597 -7646 -27563 -7612
rect -27523 -7646 -27489 -7612
rect -27449 -7646 -27415 -7612
rect -27375 -7646 -27341 -7612
rect -27301 -7646 -27267 -7612
rect -27227 -7646 -27193 -7612
rect -27153 -7646 -27119 -7612
rect -29134 -7716 -29114 -7689
rect -29114 -7716 -29100 -7689
rect -29134 -7723 -29100 -7716
rect -29046 -7723 -29012 -7689
rect -28958 -7723 -28924 -7689
rect -28870 -7723 -28836 -7689
rect -28189 -7718 -28155 -7684
rect -28115 -7718 -28081 -7684
rect -28041 -7718 -28007 -7684
rect -27967 -7718 -27933 -7684
rect -27893 -7718 -27859 -7684
rect -27819 -7718 -27785 -7684
rect -27745 -7718 -27711 -7684
rect -27671 -7718 -27637 -7684
rect -27597 -7718 -27563 -7684
rect -27523 -7718 -27489 -7684
rect -27449 -7718 -27415 -7684
rect -27375 -7718 -27341 -7684
rect -27301 -7718 -27267 -7684
rect -27227 -7718 -27193 -7684
rect -27153 -7718 -27119 -7684
rect -29134 -7784 -29114 -7761
rect -29114 -7784 -29100 -7761
rect -29134 -7795 -29100 -7784
rect -29046 -7795 -29012 -7761
rect -28958 -7795 -28924 -7761
rect -28870 -7795 -28836 -7761
rect -28189 -7790 -28155 -7756
rect -28115 -7790 -28081 -7756
rect -28041 -7790 -28007 -7756
rect -27967 -7790 -27933 -7756
rect -27893 -7790 -27859 -7756
rect -27819 -7790 -27785 -7756
rect -27745 -7790 -27711 -7756
rect -27671 -7790 -27637 -7756
rect -27597 -7790 -27563 -7756
rect -27523 -7790 -27489 -7756
rect -27449 -7790 -27415 -7756
rect -27375 -7790 -27341 -7756
rect -27301 -7790 -27267 -7756
rect -27227 -7790 -27193 -7756
rect -27153 -7790 -27119 -7756
rect -29134 -7852 -29114 -7833
rect -29114 -7852 -29100 -7833
rect -29134 -7867 -29100 -7852
rect -29046 -7867 -29012 -7833
rect -28958 -7867 -28924 -7833
rect -28870 -7867 -28836 -7833
rect -28189 -7862 -28155 -7828
rect -28115 -7862 -28081 -7828
rect -28041 -7862 -28007 -7828
rect -27967 -7862 -27933 -7828
rect -27893 -7862 -27859 -7828
rect -27819 -7862 -27785 -7828
rect -27745 -7862 -27711 -7828
rect -27671 -7862 -27637 -7828
rect -27597 -7862 -27563 -7828
rect -27523 -7862 -27489 -7828
rect -27449 -7862 -27415 -7828
rect -27375 -7862 -27341 -7828
rect -27301 -7862 -27267 -7828
rect -27227 -7862 -27193 -7828
rect -27153 -7862 -27119 -7828
rect -29134 -7920 -29114 -7905
rect -29114 -7920 -29100 -7905
rect -29134 -7939 -29100 -7920
rect -29046 -7939 -29012 -7905
rect -28958 -7939 -28924 -7905
rect -28870 -7939 -28836 -7905
rect -28189 -7934 -28155 -7900
rect -28115 -7934 -28081 -7900
rect -28041 -7934 -28007 -7900
rect -27967 -7934 -27933 -7900
rect -27893 -7934 -27859 -7900
rect -27819 -7934 -27785 -7900
rect -27745 -7934 -27711 -7900
rect -27671 -7934 -27637 -7900
rect -27597 -7934 -27563 -7900
rect -27523 -7934 -27489 -7900
rect -27449 -7934 -27415 -7900
rect -27375 -7934 -27341 -7900
rect -27301 -7934 -27267 -7900
rect -27227 -7934 -27193 -7900
rect -27153 -7934 -27119 -7900
rect -29134 -7988 -29114 -7977
rect -29114 -7988 -29100 -7977
rect -29134 -8011 -29100 -7988
rect -29046 -8011 -29012 -7977
rect -28958 -8011 -28924 -7977
rect -28870 -8011 -28836 -7977
rect -28189 -8006 -28155 -7972
rect -28115 -8006 -28081 -7972
rect -28041 -8006 -28007 -7972
rect -27967 -8006 -27933 -7972
rect -27893 -8006 -27859 -7972
rect -27819 -8006 -27785 -7972
rect -27745 -8006 -27711 -7972
rect -27671 -8006 -27637 -7972
rect -27597 -8006 -27563 -7972
rect -27523 -8006 -27489 -7972
rect -27449 -8006 -27415 -7972
rect -27375 -8006 -27341 -7972
rect -27301 -8006 -27267 -7972
rect -27227 -8006 -27193 -7972
rect -27153 -8006 -27119 -7972
rect -29134 -8056 -29114 -8049
rect -29114 -8056 -29100 -8049
rect -29134 -8083 -29100 -8056
rect -29046 -8083 -29012 -8049
rect -28958 -8083 -28924 -8049
rect -28870 -8083 -28836 -8049
rect -28189 -8078 -28155 -8044
rect -28115 -8078 -28081 -8044
rect -28041 -8078 -28007 -8044
rect -27967 -8078 -27933 -8044
rect -27893 -8078 -27859 -8044
rect -27819 -8078 -27785 -8044
rect -27745 -8078 -27711 -8044
rect -27671 -8078 -27637 -8044
rect -27597 -8078 -27563 -8044
rect -27523 -8078 -27489 -8044
rect -27449 -8078 -27415 -8044
rect -27375 -8078 -27341 -8044
rect -27301 -8078 -27267 -8044
rect -27227 -8078 -27193 -8044
rect -27153 -8078 -27119 -8044
rect -29134 -8124 -29114 -8121
rect -29114 -8124 -29100 -8121
rect -29134 -8155 -29100 -8124
rect -29046 -8155 -29012 -8121
rect -28958 -8155 -28924 -8121
rect -28870 -8155 -28836 -8121
rect -28189 -8150 -28155 -8116
rect -28115 -8150 -28081 -8116
rect -28041 -8150 -28007 -8116
rect -27967 -8150 -27933 -8116
rect -27893 -8150 -27859 -8116
rect -27819 -8150 -27785 -8116
rect -27745 -8150 -27711 -8116
rect -27671 -8150 -27637 -8116
rect -27597 -8150 -27563 -8116
rect -27523 -8150 -27489 -8116
rect -27449 -8150 -27415 -8116
rect -27375 -8150 -27341 -8116
rect -27301 -8150 -27267 -8116
rect -27227 -8150 -27193 -8116
rect -27153 -8150 -27119 -8116
rect -29134 -8226 -29100 -8193
rect -29134 -8227 -29114 -8226
rect -29114 -8227 -29100 -8226
rect -29046 -8227 -29012 -8193
rect -28958 -8227 -28924 -8193
rect -28870 -8227 -28836 -8193
rect -28189 -8222 -28155 -8188
rect -28115 -8222 -28081 -8188
rect -28041 -8222 -28007 -8188
rect -27967 -8222 -27933 -8188
rect -27893 -8222 -27859 -8188
rect -27819 -8222 -27785 -8188
rect -27745 -8222 -27711 -8188
rect -27671 -8222 -27637 -8188
rect -27597 -8222 -27563 -8188
rect -27523 -8222 -27489 -8188
rect -27449 -8222 -27415 -8188
rect -27375 -8222 -27341 -8188
rect -27301 -8222 -27267 -8188
rect -27227 -8222 -27193 -8188
rect -27153 -8222 -27119 -8188
rect -29134 -8294 -29100 -8265
rect -29134 -8299 -29114 -8294
rect -29114 -8299 -29100 -8294
rect -29046 -8299 -29012 -8265
rect -28958 -8299 -28924 -8265
rect -28870 -8299 -28836 -8265
rect -28189 -8294 -28155 -8260
rect -28115 -8294 -28081 -8260
rect -28041 -8294 -28007 -8260
rect -27967 -8294 -27933 -8260
rect -27893 -8294 -27859 -8260
rect -27819 -8294 -27785 -8260
rect -27745 -8294 -27711 -8260
rect -27671 -8294 -27637 -8260
rect -27597 -8294 -27563 -8260
rect -27523 -8294 -27489 -8260
rect -27449 -8294 -27415 -8260
rect -27375 -8294 -27341 -8260
rect -27301 -8294 -27267 -8260
rect -27227 -8294 -27193 -8260
rect -27153 -8294 -27119 -8260
rect -29134 -8362 -29100 -8337
rect -29134 -8371 -29114 -8362
rect -29114 -8371 -29100 -8362
rect -29046 -8371 -29012 -8337
rect -28958 -8371 -28924 -8337
rect -28870 -8371 -28836 -8337
rect -28189 -8366 -28155 -8332
rect -28115 -8366 -28081 -8332
rect -28041 -8366 -28007 -8332
rect -27967 -8366 -27933 -8332
rect -27893 -8366 -27859 -8332
rect -27819 -8366 -27785 -8332
rect -27745 -8366 -27711 -8332
rect -27671 -8366 -27637 -8332
rect -27597 -8366 -27563 -8332
rect -27523 -8366 -27489 -8332
rect -27449 -8366 -27415 -8332
rect -27375 -8366 -27341 -8332
rect -27301 -8366 -27267 -8332
rect -27227 -8366 -27193 -8332
rect -27153 -8366 -27119 -8332
rect -29134 -8430 -29100 -8409
rect -29134 -8443 -29114 -8430
rect -29114 -8443 -29100 -8430
rect -29046 -8443 -29012 -8409
rect -28958 -8443 -28924 -8409
rect -28870 -8443 -28836 -8409
rect -28189 -8438 -28155 -8404
rect -28115 -8438 -28081 -8404
rect -28041 -8438 -28007 -8404
rect -27967 -8438 -27933 -8404
rect -27893 -8438 -27859 -8404
rect -27819 -8438 -27785 -8404
rect -27745 -8438 -27711 -8404
rect -27671 -8438 -27637 -8404
rect -27597 -8438 -27563 -8404
rect -27523 -8438 -27489 -8404
rect -27449 -8438 -27415 -8404
rect -27375 -8438 -27341 -8404
rect -27301 -8438 -27267 -8404
rect -27227 -8438 -27193 -8404
rect -27153 -8438 -27119 -8404
rect -29134 -8498 -29100 -8481
rect -29134 -8515 -29114 -8498
rect -29114 -8515 -29100 -8498
rect -29046 -8515 -29012 -8481
rect -28958 -8515 -28924 -8481
rect -28870 -8515 -28836 -8481
rect -28189 -8510 -28155 -8476
rect -28115 -8510 -28081 -8476
rect -28041 -8510 -28007 -8476
rect -27967 -8510 -27933 -8476
rect -27893 -8510 -27859 -8476
rect -27819 -8510 -27785 -8476
rect -27745 -8510 -27711 -8476
rect -27671 -8510 -27637 -8476
rect -27597 -8510 -27563 -8476
rect -27523 -8510 -27489 -8476
rect -27449 -8510 -27415 -8476
rect -27375 -8510 -27341 -8476
rect -27301 -8510 -27267 -8476
rect -27227 -8510 -27193 -8476
rect -27153 -8510 -27119 -8476
rect -29134 -8566 -29100 -8553
rect -29134 -8587 -29114 -8566
rect -29114 -8587 -29100 -8566
rect -29046 -8587 -29012 -8553
rect -28958 -8587 -28924 -8553
rect -28870 -8587 -28836 -8553
rect -28189 -8582 -28155 -8548
rect -28115 -8582 -28081 -8548
rect -28041 -8582 -28007 -8548
rect -27967 -8582 -27933 -8548
rect -27893 -8582 -27859 -8548
rect -27819 -8582 -27785 -8548
rect -27745 -8582 -27711 -8548
rect -27671 -8582 -27637 -8548
rect -27597 -8582 -27563 -8548
rect -27523 -8582 -27489 -8548
rect -27449 -8582 -27415 -8548
rect -27375 -8582 -27341 -8548
rect -27301 -8582 -27267 -8548
rect -27227 -8582 -27193 -8548
rect -27153 -8582 -27119 -8548
rect -32344 -8712 -32315 -8678
rect -32315 -8712 -32310 -8678
rect -32266 -8712 -32232 -8678
rect -32188 -8712 -32154 -8678
rect -32110 -8712 -32076 -8678
rect -32032 -8712 -31998 -8678
rect -31954 -8712 -31920 -8678
rect -31876 -8712 -31842 -8678
rect -31798 -8712 -31764 -8678
rect -31512 -8659 -31478 -8625
rect -31512 -8719 -31478 -8697
rect -31512 -8731 -31478 -8719
rect -29268 -8627 -29234 -8593
rect -29268 -8697 -29234 -8665
rect -29268 -8699 -29234 -8697
rect -29134 -8634 -29100 -8625
rect -29134 -8659 -29114 -8634
rect -29114 -8659 -29100 -8634
rect -29046 -8659 -29012 -8625
rect -28958 -8659 -28924 -8625
rect -28870 -8659 -28836 -8625
rect -28189 -8654 -28155 -8620
rect -28115 -8654 -28081 -8620
rect -28041 -8654 -28007 -8620
rect -27967 -8654 -27933 -8620
rect -27893 -8654 -27859 -8620
rect -27819 -8654 -27785 -8620
rect -27745 -8654 -27711 -8620
rect -27671 -8654 -27637 -8620
rect -27597 -8654 -27563 -8620
rect -27523 -8654 -27489 -8620
rect -27449 -8654 -27415 -8620
rect -27375 -8654 -27341 -8620
rect -27301 -8654 -27267 -8620
rect -27227 -8654 -27193 -8620
rect -27153 -8654 -27119 -8620
rect -29134 -8702 -29100 -8697
rect -29134 -8731 -29114 -8702
rect -29114 -8731 -29100 -8702
rect -29046 -8731 -29012 -8697
rect -28958 -8731 -28924 -8697
rect -28870 -8731 -28836 -8697
rect -28189 -8726 -28155 -8692
rect -28115 -8726 -28081 -8692
rect -28041 -8726 -28007 -8692
rect -27967 -8726 -27933 -8692
rect -27893 -8726 -27859 -8692
rect -27819 -8726 -27785 -8692
rect -27745 -8726 -27711 -8692
rect -27671 -8726 -27637 -8692
rect -27597 -8726 -27563 -8692
rect -27523 -8726 -27489 -8692
rect -27449 -8726 -27415 -8692
rect -27375 -8726 -27341 -8692
rect -27301 -8726 -27267 -8692
rect -27227 -8726 -27193 -8692
rect -27153 -8726 -27119 -8692
rect -32344 -8784 -32315 -8750
rect -32315 -8784 -32310 -8750
rect -32266 -8784 -32232 -8750
rect -32188 -8784 -32154 -8750
rect -32110 -8784 -32076 -8750
rect -32032 -8784 -31998 -8750
rect -31954 -8784 -31920 -8750
rect -31876 -8784 -31842 -8750
rect -31798 -8784 -31764 -8750
rect -29134 -8803 -29100 -8769
rect -29046 -8803 -29012 -8769
rect -28958 -8803 -28924 -8769
rect -28870 -8803 -28836 -8769
rect -28189 -8798 -28155 -8764
rect -28115 -8798 -28081 -8764
rect -28041 -8798 -28007 -8764
rect -27967 -8798 -27933 -8764
rect -27893 -8798 -27859 -8764
rect -27819 -8798 -27785 -8764
rect -27745 -8798 -27711 -8764
rect -27671 -8798 -27637 -8764
rect -27597 -8798 -27563 -8764
rect -27523 -8798 -27489 -8764
rect -27449 -8798 -27415 -8764
rect -27375 -8798 -27341 -8764
rect -27301 -8798 -27267 -8764
rect -27227 -8798 -27193 -8764
rect -27153 -8798 -27119 -8764
rect -32344 -8856 -32315 -8822
rect -32315 -8856 -32310 -8822
rect -32266 -8856 -32232 -8822
rect -32188 -8856 -32154 -8822
rect -32110 -8856 -32076 -8822
rect -32032 -8856 -31998 -8822
rect -31954 -8856 -31920 -8822
rect -31876 -8856 -31842 -8822
rect -31798 -8856 -31764 -8822
rect -29134 -8875 -29100 -8841
rect -29046 -8847 -29012 -8841
rect -28958 -8847 -28924 -8841
rect -28870 -8847 -28836 -8841
rect -28189 -8847 -28155 -8836
rect -28115 -8847 -28081 -8836
rect -28041 -8847 -28007 -8836
rect -27967 -8847 -27933 -8836
rect -27893 -8847 -27859 -8836
rect -27819 -8847 -27785 -8836
rect -27745 -8847 -27711 -8836
rect -27671 -8847 -27637 -8836
rect -27597 -8847 -27563 -8836
rect -27523 -8847 -27489 -8836
rect -27449 -8847 -27415 -8836
rect -27375 -8847 -27341 -8836
rect -27301 -8847 -27267 -8836
rect -27227 -8847 -27193 -8836
rect -27153 -8847 -27119 -8836
rect 244 2225 278 2241
rect 244 2207 278 2225
rect 244 2157 278 2169
rect 244 2135 278 2157
rect 244 2089 278 2097
rect 244 2063 278 2089
rect 480 2225 514 2241
rect 480 2207 514 2225
rect 1299 2235 1333 2269
rect 1413 2235 1447 2269
rect 2152 2205 2186 2239
rect 2224 2205 2258 2239
rect 4207 3619 4241 3653
rect 4290 3619 4293 3653
rect 4293 3619 4324 3653
rect 4373 3619 4395 3653
rect 4395 3619 4407 3653
rect 4456 3619 4463 3653
rect 4463 3619 4490 3653
rect 4125 3547 4159 3581
rect 4528 3551 4529 3579
rect 4529 3551 4562 3579
rect 4125 3479 4159 3505
rect 4125 3471 4159 3479
rect 4125 3411 4159 3429
rect 4125 3395 4159 3411
rect 4125 3343 4159 3353
rect 4125 3319 4159 3343
rect 4125 3275 4159 3277
rect 4125 3243 4159 3275
rect 4125 3173 4159 3201
rect 4125 3167 4159 3173
rect 4125 3105 4159 3125
rect 4125 3091 4159 3105
rect 4125 3037 4159 3049
rect 4125 3015 4159 3037
rect 4125 2969 4159 2973
rect 4125 2939 4159 2969
rect 4125 2867 4159 2897
rect 4125 2863 4159 2867
rect 4125 2799 4159 2821
rect 4125 2787 4159 2799
rect 4125 2731 4159 2745
rect 4125 2711 4159 2731
rect 4125 2663 4159 2669
rect 4125 2635 4159 2663
rect 4125 2561 4159 2593
rect 4244 3533 4278 3549
rect 4244 3515 4278 3533
rect 4244 3465 4278 3477
rect 4244 3443 4278 3465
rect 4244 3397 4278 3405
rect 4244 3371 4278 3397
rect 4244 3329 4278 3333
rect 4244 3299 4278 3329
rect 4244 3227 4278 3261
rect 4244 3159 4278 3189
rect 4244 3155 4278 3159
rect 4244 3091 4278 3117
rect 4244 3083 4278 3091
rect 4244 3023 4278 3045
rect 4244 3011 4278 3023
rect 4244 2955 4278 2973
rect 4244 2939 4278 2955
rect 4244 2887 4278 2901
rect 4244 2867 4278 2887
rect 4244 2819 4278 2829
rect 4244 2795 4278 2819
rect 4244 2751 4278 2757
rect 4244 2723 4278 2751
rect 4244 2683 4278 2685
rect 4244 2651 4278 2683
rect 4244 2579 4278 2613
rect 4400 3533 4434 3549
rect 4400 3515 4434 3533
rect 4400 3465 4434 3477
rect 4400 3443 4434 3465
rect 4400 3397 4434 3405
rect 4400 3371 4434 3397
rect 4400 3329 4434 3333
rect 4400 3299 4434 3329
rect 4400 3227 4434 3261
rect 4400 3159 4434 3189
rect 4400 3155 4434 3159
rect 4400 3091 4434 3117
rect 4400 3083 4434 3091
rect 4400 3023 4434 3045
rect 4400 3011 4434 3023
rect 4400 2955 4434 2973
rect 4400 2939 4434 2955
rect 4400 2887 4434 2901
rect 4400 2867 4434 2887
rect 4400 2819 4434 2829
rect 4400 2795 4434 2819
rect 4400 2751 4434 2757
rect 4400 2723 4434 2751
rect 4400 2683 4434 2685
rect 4400 2651 4434 2683
rect 4400 2579 4434 2613
rect 4528 3545 4562 3551
rect 4528 3483 4529 3505
rect 4529 3483 4562 3505
rect 4528 3471 4562 3483
rect 4528 3415 4529 3431
rect 4529 3415 4562 3431
rect 4528 3397 4562 3415
rect 4528 3347 4529 3357
rect 4529 3347 4562 3357
rect 4528 3323 4562 3347
rect 4528 3279 4529 3283
rect 4529 3279 4562 3283
rect 4528 3249 4562 3279
rect 4528 3177 4562 3209
rect 4528 3175 4529 3177
rect 4529 3175 4562 3177
rect 4528 3109 4562 3135
rect 4528 3101 4529 3109
rect 4529 3101 4562 3109
rect 4528 3041 4562 3061
rect 4528 3027 4529 3041
rect 4529 3027 4562 3041
rect 4528 2973 4562 2987
rect 4528 2953 4529 2973
rect 4529 2953 4562 2973
rect 4528 2905 4562 2912
rect 4528 2878 4529 2905
rect 4529 2878 4562 2905
rect 4528 2803 4529 2837
rect 4529 2803 4562 2837
rect 4528 2735 4529 2762
rect 4529 2735 4562 2762
rect 4528 2728 4562 2735
rect 4528 2667 4529 2687
rect 4529 2667 4562 2687
rect 4528 2653 4562 2667
rect 4528 2599 4529 2612
rect 4529 2599 4562 2612
rect 4125 2559 4159 2561
rect 4125 2493 4159 2517
rect 4528 2578 4562 2599
rect 4528 2531 4529 2537
rect 4529 2531 4562 2537
rect 4125 2483 4159 2493
rect 4125 2425 4159 2441
rect 4125 2407 4159 2425
rect 4323 2455 4324 2481
rect 4324 2455 4357 2481
rect 4323 2447 4357 2455
rect 4323 2387 4324 2409
rect 4324 2387 4357 2409
rect 4323 2375 4357 2387
rect 4528 2503 4562 2531
rect 4528 2429 4562 2462
rect 4528 2428 4529 2429
rect 4529 2428 4562 2429
rect 4125 2357 4159 2365
rect 4125 2331 4159 2357
rect 4528 2361 4562 2387
rect 4528 2353 4529 2361
rect 4529 2353 4562 2361
rect 4197 2255 4231 2289
rect 4286 2255 4291 2289
rect 4291 2255 4320 2289
rect 4718 3644 4752 3669
rect 4802 3644 4836 3669
rect 4886 3644 4920 3669
rect 5738 3738 5772 3758
rect 5738 3724 5772 3738
rect 5738 3670 5772 3676
rect 4718 3600 4723 3603
rect 4723 3600 4752 3603
rect 4802 3600 4815 3603
rect 4815 3600 4836 3603
rect 4886 3600 4907 3603
rect 4907 3600 4920 3603
rect 4718 3569 4752 3600
rect 4802 3569 4836 3600
rect 4886 3569 4920 3600
rect 4718 3496 4752 3528
rect 4802 3496 4836 3528
rect 4886 3496 4920 3528
rect 4718 3494 4723 3496
rect 4723 3494 4752 3496
rect 4802 3494 4815 3496
rect 4815 3494 4836 3496
rect 4886 3494 4907 3496
rect 4907 3494 4920 3496
rect 4718 3427 4752 3453
rect 4802 3427 4836 3453
rect 4886 3427 4920 3453
rect 4718 3419 4723 3427
rect 4723 3419 4752 3427
rect 4802 3419 4815 3427
rect 4815 3419 4836 3427
rect 4886 3419 4907 3427
rect 4907 3419 4920 3427
rect 4718 3358 4752 3378
rect 4802 3358 4836 3378
rect 4886 3358 4920 3378
rect 4718 3344 4723 3358
rect 4723 3344 4752 3358
rect 4802 3344 4815 3358
rect 4815 3344 4836 3358
rect 4886 3344 4907 3358
rect 4907 3344 4920 3358
rect 4718 3289 4752 3303
rect 4802 3289 4836 3303
rect 4886 3289 4920 3303
rect 4718 3269 4723 3289
rect 4723 3269 4752 3289
rect 4802 3269 4815 3289
rect 4815 3269 4836 3289
rect 4886 3269 4907 3289
rect 4907 3269 4920 3289
rect 4718 3220 4752 3228
rect 4802 3220 4836 3228
rect 4886 3220 4920 3228
rect 4718 3194 4723 3220
rect 4723 3194 4752 3220
rect 4802 3194 4815 3220
rect 4815 3194 4836 3220
rect 4886 3194 4907 3220
rect 4907 3194 4920 3220
rect 4718 3150 4752 3153
rect 4802 3150 4836 3153
rect 4886 3150 4920 3153
rect 4718 3119 4723 3150
rect 4723 3119 4752 3150
rect 4802 3119 4815 3150
rect 4815 3119 4836 3150
rect 4886 3119 4907 3150
rect 4907 3119 4920 3150
rect 4718 3046 4723 3078
rect 4723 3046 4752 3078
rect 4802 3046 4815 3078
rect 4815 3046 4836 3078
rect 4886 3046 4907 3078
rect 4907 3046 4920 3078
rect 4718 3044 4752 3046
rect 4802 3044 4836 3046
rect 4886 3044 4920 3046
rect 4718 2976 4723 3003
rect 4723 2976 4752 3003
rect 4802 2976 4815 3003
rect 4815 2976 4836 3003
rect 4886 2976 4907 3003
rect 4907 2976 4920 3003
rect 4718 2969 4752 2976
rect 4802 2969 4836 2976
rect 4886 2969 4920 2976
rect 4718 2906 4723 2928
rect 4723 2906 4752 2928
rect 4802 2906 4815 2928
rect 4815 2906 4836 2928
rect 4886 2906 4907 2928
rect 4907 2906 4920 2928
rect 4718 2894 4752 2906
rect 4802 2894 4836 2906
rect 4886 2894 4920 2906
rect 4718 2836 4723 2853
rect 4723 2836 4752 2853
rect 4802 2836 4815 2853
rect 4815 2836 4836 2853
rect 4886 2836 4907 2853
rect 4907 2836 4920 2853
rect 4718 2819 4752 2836
rect 4802 2819 4836 2836
rect 4886 2819 4920 2836
rect 4718 2766 4723 2778
rect 4723 2766 4752 2778
rect 4802 2766 4815 2778
rect 4815 2766 4836 2778
rect 4886 2766 4907 2778
rect 4907 2766 4920 2778
rect 4718 2744 4752 2766
rect 4802 2744 4836 2766
rect 4886 2744 4920 2766
rect 4718 2696 4723 2703
rect 4723 2696 4752 2703
rect 4802 2696 4815 2703
rect 4815 2696 4836 2703
rect 4886 2696 4907 2703
rect 4907 2696 4920 2703
rect 4718 2669 4752 2696
rect 4802 2669 4836 2696
rect 4886 2669 4920 2696
rect 4718 2626 4723 2628
rect 4723 2626 4752 2628
rect 4802 2626 4815 2628
rect 4815 2626 4836 2628
rect 4886 2626 4907 2628
rect 4907 2626 4920 2628
rect 4718 2594 4752 2626
rect 4802 2594 4836 2626
rect 4886 2594 4920 2626
rect 4718 2520 4752 2553
rect 4802 2520 4836 2553
rect 4886 2520 4920 2553
rect 4718 2519 4723 2520
rect 4723 2519 4752 2520
rect 4802 2519 4815 2520
rect 4815 2519 4836 2520
rect 4886 2519 4907 2520
rect 4907 2519 4920 2520
rect 4718 2450 4752 2478
rect 4802 2450 4836 2478
rect 4886 2450 4920 2478
rect 4718 2444 4723 2450
rect 4723 2444 4752 2450
rect 4802 2444 4815 2450
rect 4815 2444 4836 2450
rect 4886 2444 4907 2450
rect 4907 2444 4920 2450
rect 4718 2380 4752 2403
rect 4802 2380 4836 2403
rect 4886 2380 4920 2403
rect 4718 2369 4723 2380
rect 4723 2369 4752 2380
rect 4802 2369 4815 2380
rect 4815 2369 4836 2380
rect 4886 2369 4907 2380
rect 4907 2369 4920 2380
rect 4718 2310 4752 2328
rect 4802 2310 4836 2328
rect 4886 2310 4920 2328
rect 4718 2294 4723 2310
rect 4723 2294 4752 2310
rect 4802 2294 4815 2310
rect 4815 2294 4836 2310
rect 4886 2294 4907 2310
rect 4907 2294 4920 2310
rect 5173 3619 5197 3653
rect 5197 3619 5207 3653
rect 5249 3619 5265 3653
rect 5265 3619 5283 3653
rect 5325 3619 5333 3653
rect 5333 3619 5359 3653
rect 5402 3619 5436 3653
rect 5479 3619 5483 3653
rect 5483 3619 5513 3653
rect 5097 3551 5131 3581
rect 5097 3547 5131 3551
rect 5097 3483 5131 3505
rect 5551 3547 5585 3581
rect 5097 3471 5131 3483
rect 5097 3415 5131 3429
rect 5097 3395 5131 3415
rect 5097 3347 5131 3353
rect 5097 3319 5131 3347
rect 5216 3436 5250 3462
rect 5216 3428 5250 3436
rect 5216 3368 5250 3390
rect 5216 3356 5250 3368
rect 5216 3300 5250 3318
rect 5216 3284 5250 3300
rect 5432 3436 5466 3462
rect 5432 3428 5466 3436
rect 5432 3368 5466 3390
rect 5432 3356 5466 3368
rect 5432 3300 5466 3318
rect 5432 3284 5466 3300
rect 5551 3479 5585 3509
rect 5551 3475 5585 3479
rect 5551 3411 5585 3437
rect 5551 3403 5585 3411
rect 5551 3343 5585 3365
rect 5551 3331 5585 3343
rect 5097 3245 5131 3277
rect 5097 3243 5131 3245
rect 5551 3275 5585 3293
rect 5551 3259 5585 3275
rect 5097 3177 5131 3201
rect 5097 3167 5131 3177
rect 5097 3109 5131 3125
rect 5097 3091 5131 3109
rect 5327 3216 5361 3217
rect 5327 3183 5360 3216
rect 5360 3183 5361 3216
rect 5327 3114 5360 3145
rect 5360 3114 5361 3145
rect 5327 3111 5361 3114
rect 5551 3207 5585 3220
rect 5551 3186 5585 3207
rect 5551 3139 5585 3147
rect 5551 3113 5585 3139
rect 5097 3041 5131 3049
rect 5097 3015 5131 3041
rect 5551 3071 5585 3074
rect 5551 3040 5585 3071
rect 5097 2939 5131 2973
rect 5097 2871 5131 2897
rect 5097 2863 5131 2871
rect 5097 2803 5131 2821
rect 5097 2787 5131 2803
rect 5216 2930 5250 2956
rect 5216 2922 5250 2930
rect 5216 2862 5250 2884
rect 5216 2850 5250 2862
rect 5216 2794 5250 2812
rect 5216 2778 5250 2794
rect 5329 2902 5363 2936
rect 5329 2830 5363 2864
rect 5097 2735 5131 2745
rect 5097 2711 5131 2735
rect 5097 2667 5131 2669
rect 5097 2635 5131 2667
rect 5097 2565 5131 2593
rect 5432 2930 5466 2956
rect 5432 2922 5466 2930
rect 5432 2862 5466 2884
rect 5432 2850 5466 2862
rect 5432 2794 5466 2812
rect 5432 2778 5466 2794
rect 5551 2969 5585 3001
rect 5551 2967 5585 2969
rect 5551 2901 5585 2928
rect 5551 2894 5585 2901
rect 5551 2833 5585 2855
rect 5551 2821 5585 2833
rect 5551 2765 5585 2782
rect 5551 2748 5585 2765
rect 5551 2697 5585 2709
rect 5551 2675 5585 2697
rect 5097 2559 5131 2565
rect 5097 2497 5131 2517
rect 5097 2483 5131 2497
rect 5097 2429 5131 2441
rect 5097 2407 5131 2429
rect 5097 2361 5131 2365
rect 5097 2331 5131 2361
rect 5169 2255 5199 2289
rect 5199 2255 5203 2289
rect 5245 2255 5267 2289
rect 5267 2255 5279 2289
rect 5320 2255 5335 2289
rect 5335 2255 5354 2289
rect 5395 2255 5403 2289
rect 5403 2255 5429 2289
rect 5470 2255 5471 2289
rect 5471 2255 5504 2289
rect 5545 2255 5579 2289
rect 5738 3642 5772 3670
rect 5738 3568 5772 3594
rect 5738 3560 5772 3568
rect 5738 3500 5772 3512
rect 5738 3478 5772 3500
rect 5738 3398 5772 3429
rect 5738 3395 5772 3398
rect 5738 3330 5772 3342
rect 5738 3308 5772 3330
rect 5829 3283 5863 3317
rect 5901 3283 5912 3317
rect 5912 3283 5935 3317
rect 6580 3283 6606 3317
rect 6606 3283 6614 3317
rect 6652 3283 6686 3317
rect 6730 3301 6764 3333
rect 6730 3299 6732 3301
rect 6732 3299 6764 3301
rect 5738 3262 5772 3265
rect 5738 3231 5772 3262
rect 5738 3160 5772 3187
rect 6032 3248 6066 3282
rect 6032 3192 6040 3210
rect 6040 3192 6066 3210
rect 6032 3176 6066 3192
rect 6730 3227 6764 3253
rect 6730 3219 6732 3227
rect 6732 3219 6764 3227
rect 5738 3153 5772 3160
rect 6730 3153 6764 3174
rect 5738 3092 5772 3109
rect 5738 3075 5772 3092
rect 5738 3024 5772 3031
rect 5738 2997 5772 3024
rect 6260 3107 6276 3141
rect 6276 3107 6294 3141
rect 6332 3107 6344 3141
rect 6344 3107 6366 3141
rect 6730 3140 6732 3153
rect 6732 3140 6764 3153
rect 6730 3079 6764 3095
rect 6119 3055 6153 3069
rect 6119 3035 6142 3055
rect 6142 3035 6153 3055
rect 5738 2922 5772 2953
rect 6119 2963 6153 2997
rect 6730 3061 6732 3079
rect 6732 3061 6764 3079
rect 6730 3005 6764 3016
rect 6730 2982 6732 3005
rect 6732 2982 6764 3005
rect 6580 2931 6606 2965
rect 6606 2931 6614 2965
rect 6652 2931 6686 2965
rect 6730 2931 6764 2937
rect 5738 2919 5772 2922
rect 5738 2854 5772 2875
rect 5738 2841 5772 2854
rect 6730 2903 6732 2931
rect 6732 2903 6764 2931
rect 5829 2806 5863 2840
rect 5901 2806 5912 2840
rect 5912 2806 5935 2840
rect 6580 2806 6606 2840
rect 6606 2806 6614 2840
rect 6652 2806 6686 2840
rect 6730 2824 6732 2858
rect 6732 2824 6764 2858
rect 5738 2786 5772 2797
rect 5738 2763 5772 2786
rect 5738 2718 5772 2719
rect 5738 2685 5772 2718
rect 6210 2716 6244 2750
rect 6282 2716 6316 2750
rect 6730 2751 6732 2779
rect 6732 2751 6764 2779
rect 6730 2745 6764 2751
rect 6730 2678 6732 2700
rect 6732 2678 6764 2700
rect 6730 2666 6764 2678
rect 5738 2616 5772 2641
rect 6259 2630 6276 2664
rect 6276 2630 6293 2664
rect 6331 2630 6344 2664
rect 6344 2630 6365 2664
rect 5738 2607 5772 2616
rect 6730 2605 6732 2621
rect 6732 2605 6764 2621
rect 6730 2587 6764 2605
rect 4718 2240 4752 2254
rect 4802 2240 4836 2254
rect 4886 2240 4920 2254
rect 4718 2220 4723 2240
rect 4723 2220 4752 2240
rect 4802 2220 4815 2240
rect 4815 2220 4836 2240
rect 4886 2220 4907 2240
rect 4907 2220 4920 2240
rect 480 2157 514 2169
rect 480 2135 514 2157
rect 480 2089 514 2097
rect 480 2063 514 2089
rect 1299 2147 1333 2181
rect 1413 2147 1447 2181
rect 778 2086 812 2120
rect 862 2086 896 2120
rect 946 2086 980 2120
rect 1030 2086 1064 2120
rect 1114 2086 1148 2120
rect 1299 2060 1333 2094
rect 1413 2060 1447 2094
rect 3520 2065 3554 2071
rect -164 1949 -160 1982
rect -160 1949 -130 1982
rect -90 1949 -66 1982
rect -66 1949 -56 1982
rect 184 1952 187 1986
rect 187 1952 218 1986
rect 261 1952 262 1986
rect 262 1952 295 1986
rect 338 1952 371 1986
rect 371 1952 372 1986
rect 415 1952 445 1986
rect 445 1952 449 1986
rect 492 1952 519 1986
rect 519 1952 526 1986
rect 569 1952 593 1986
rect 593 1952 603 1986
rect 645 1952 667 1986
rect 667 1952 679 1986
rect 721 1952 741 1986
rect 741 1952 755 1986
rect 797 1952 815 1986
rect 815 1952 831 1986
rect 873 1952 889 1986
rect 889 1952 907 1986
rect 1070 1949 1085 1983
rect 1085 1949 1104 1983
rect 1145 1949 1159 1983
rect 1159 1949 1179 1983
rect 1220 1949 1233 1983
rect 1233 1949 1254 1983
rect 1294 1949 1307 1983
rect 1307 1949 1328 1983
rect 1368 1949 1381 1983
rect 1381 1949 1402 1983
rect 1442 1949 1455 1983
rect 1455 1949 1476 1983
rect 1516 1949 1529 1983
rect 1529 1949 1550 1983
rect 1590 1949 1603 1983
rect 1603 1949 1624 1983
rect 1664 1949 1677 1983
rect 1677 1949 1698 1983
rect 1738 1949 1752 1983
rect 1752 1949 1772 1983
rect -164 1948 -130 1949
rect -90 1948 -56 1949
rect -221 1833 -187 1867
rect -221 1763 -187 1795
rect -221 1761 -187 1763
rect -710 1656 -676 1690
rect -638 1656 -604 1690
rect -530 1669 -496 1703
rect -530 1597 -496 1631
rect -221 1695 -187 1723
rect -221 1689 -187 1695
rect -221 1627 -187 1651
rect -221 1617 -187 1627
rect -221 1559 -187 1579
rect -221 1545 -187 1559
rect -221 1491 -187 1507
rect -221 1473 -187 1491
rect -221 1423 -187 1435
rect -221 1401 -187 1423
rect -221 1355 -187 1363
rect -221 1329 -187 1355
rect -221 1287 -187 1291
rect -221 1257 -187 1287
rect -221 1185 -187 1219
rect -221 1117 -187 1147
rect -221 1113 -187 1117
rect -221 1049 -187 1075
rect -221 1041 -187 1049
rect -221 981 -187 1003
rect -221 969 -187 981
rect -221 913 -187 931
rect -221 897 -187 913
rect -5 1833 29 1867
rect -5 1763 29 1795
rect -5 1761 29 1763
rect -5 1695 29 1723
rect -5 1689 29 1695
rect -5 1627 29 1651
rect -5 1617 29 1627
rect -5 1559 29 1579
rect -5 1545 29 1559
rect -5 1491 29 1507
rect -5 1473 29 1491
rect -5 1423 29 1435
rect -5 1401 29 1423
rect -5 1355 29 1363
rect -5 1329 29 1355
rect -5 1287 29 1291
rect -5 1257 29 1287
rect -5 1185 29 1219
rect -5 1117 29 1147
rect -5 1113 29 1117
rect -5 1049 29 1075
rect -5 1041 29 1049
rect -5 981 29 1003
rect -5 969 29 981
rect -5 913 29 931
rect -5 897 29 913
rect 126 1833 160 1867
rect 126 1763 160 1795
rect 126 1761 160 1763
rect 126 1695 160 1723
rect 126 1689 160 1695
rect 126 1627 160 1651
rect 126 1617 160 1627
rect 126 1559 160 1579
rect 126 1545 160 1559
rect 126 1491 160 1507
rect 126 1473 160 1491
rect 126 1423 160 1435
rect 126 1401 160 1423
rect 126 1355 160 1363
rect 126 1329 160 1355
rect 126 1287 160 1291
rect 126 1257 160 1287
rect 126 1185 160 1219
rect 126 1117 160 1147
rect 126 1113 160 1117
rect 126 1049 160 1075
rect 126 1041 160 1049
rect 126 981 160 1003
rect 126 969 160 981
rect 126 913 160 931
rect 126 897 160 913
rect 342 1833 376 1867
rect 342 1763 376 1795
rect 342 1761 376 1763
rect 342 1695 376 1723
rect 342 1689 376 1695
rect 342 1627 376 1651
rect 342 1617 376 1627
rect 342 1559 376 1579
rect 342 1545 376 1559
rect 342 1491 376 1507
rect 342 1473 376 1491
rect 342 1423 376 1435
rect 342 1401 376 1423
rect 342 1355 376 1363
rect 342 1329 376 1355
rect 342 1287 376 1291
rect 342 1257 376 1287
rect 342 1185 376 1219
rect 342 1117 376 1147
rect 342 1113 376 1117
rect 342 1049 376 1075
rect 342 1041 376 1049
rect 342 981 376 1003
rect 342 969 376 981
rect 342 913 376 931
rect 342 897 376 913
rect 558 1833 592 1867
rect 558 1763 592 1795
rect 558 1761 592 1763
rect 558 1695 592 1723
rect 558 1689 592 1695
rect 558 1627 592 1651
rect 558 1617 592 1627
rect 558 1559 592 1579
rect 558 1545 592 1559
rect 558 1491 592 1507
rect 558 1473 592 1491
rect 558 1423 592 1435
rect 558 1401 592 1423
rect 558 1355 592 1363
rect 558 1329 592 1355
rect 558 1287 592 1291
rect 558 1257 592 1287
rect 558 1185 592 1219
rect 558 1117 592 1147
rect 558 1113 592 1117
rect 558 1049 592 1075
rect 558 1041 592 1049
rect 558 981 592 1003
rect 558 969 592 981
rect 558 913 592 931
rect 558 897 592 913
rect 774 1833 808 1867
rect 774 1763 808 1795
rect 774 1761 808 1763
rect 774 1695 808 1723
rect 774 1689 808 1695
rect 774 1627 808 1651
rect 774 1617 808 1627
rect 774 1559 808 1579
rect 774 1545 808 1559
rect 774 1491 808 1507
rect 774 1473 808 1491
rect 774 1423 808 1435
rect 774 1401 808 1423
rect 774 1355 808 1363
rect 774 1329 808 1355
rect 774 1287 808 1291
rect 774 1257 808 1287
rect 774 1185 808 1219
rect 774 1117 808 1147
rect 774 1113 808 1117
rect 774 1049 808 1075
rect 774 1041 808 1049
rect 774 981 808 1003
rect 774 969 808 981
rect 774 913 808 931
rect 774 897 808 913
rect 990 1833 1024 1867
rect 990 1763 1024 1795
rect 990 1761 1024 1763
rect 990 1695 1024 1723
rect 990 1689 1024 1695
rect 990 1627 1024 1651
rect 990 1617 1024 1627
rect 990 1559 1024 1579
rect 990 1545 1024 1559
rect 990 1491 1024 1507
rect 990 1473 1024 1491
rect 990 1423 1024 1435
rect 990 1401 1024 1423
rect 990 1355 1024 1363
rect 990 1329 1024 1355
rect 990 1287 1024 1291
rect 990 1257 1024 1287
rect 990 1185 1024 1219
rect 990 1117 1024 1147
rect 990 1113 1024 1117
rect 990 1049 1024 1075
rect 990 1041 1024 1049
rect 990 981 1024 1003
rect 990 969 1024 981
rect 990 913 1024 931
rect 990 897 1024 913
rect 1206 1833 1240 1867
rect 1206 1763 1240 1795
rect 1206 1761 1240 1763
rect 1206 1695 1240 1723
rect 1206 1689 1240 1695
rect 1206 1627 1240 1651
rect 1206 1617 1240 1627
rect 1206 1559 1240 1579
rect 1206 1545 1240 1559
rect 1206 1491 1240 1507
rect 1206 1473 1240 1491
rect 1206 1423 1240 1435
rect 1206 1401 1240 1423
rect 1206 1355 1240 1363
rect 1206 1329 1240 1355
rect 1206 1287 1240 1291
rect 1206 1257 1240 1287
rect 1206 1185 1240 1219
rect 1206 1117 1240 1147
rect 1206 1113 1240 1117
rect 1206 1049 1240 1075
rect 1206 1041 1240 1049
rect 1206 981 1240 1003
rect 1206 969 1240 981
rect 1206 913 1240 931
rect 1206 897 1240 913
rect 1422 1833 1456 1867
rect 1422 1763 1456 1795
rect 1422 1761 1456 1763
rect 1422 1695 1456 1723
rect 1422 1689 1456 1695
rect 1422 1627 1456 1651
rect 1422 1617 1456 1627
rect 1422 1559 1456 1579
rect 1422 1545 1456 1559
rect 1422 1491 1456 1507
rect 1422 1473 1456 1491
rect 1422 1423 1456 1435
rect 1422 1401 1456 1423
rect 1422 1355 1456 1363
rect 1422 1329 1456 1355
rect 1422 1287 1456 1291
rect 1422 1257 1456 1287
rect 1422 1185 1456 1219
rect 1422 1117 1456 1147
rect 1422 1113 1456 1117
rect 1422 1049 1456 1075
rect 1422 1041 1456 1049
rect 1422 981 1456 1003
rect 1422 969 1456 981
rect 1422 913 1456 931
rect 1422 897 1456 913
rect 1638 1833 1672 1867
rect 1638 1763 1672 1795
rect 1638 1761 1672 1763
rect 1638 1695 1672 1723
rect 1638 1689 1672 1695
rect 1638 1627 1672 1651
rect 1638 1617 1672 1627
rect 1638 1559 1672 1579
rect 1638 1545 1672 1559
rect 1638 1491 1672 1507
rect 1638 1473 1672 1491
rect 1638 1423 1672 1435
rect 1638 1401 1672 1423
rect 1638 1355 1672 1363
rect 1638 1329 1672 1355
rect 1638 1287 1672 1291
rect 1638 1257 1672 1287
rect 1638 1185 1672 1219
rect 1638 1117 1672 1147
rect 1638 1113 1672 1117
rect 1638 1049 1672 1075
rect 1638 1041 1672 1049
rect 1638 981 1672 1003
rect 1638 969 1672 981
rect 1638 913 1672 931
rect 1638 897 1672 913
rect 1854 1833 1888 1867
rect 1854 1763 1888 1795
rect 1854 1761 1888 1763
rect 1854 1695 1888 1723
rect 1854 1689 1888 1695
rect 1854 1627 1888 1651
rect 1854 1617 1888 1627
rect 1854 1559 1888 1579
rect 1854 1545 1888 1559
rect 1854 1491 1888 1507
rect 1854 1473 1888 1491
rect 1854 1423 1888 1435
rect 1854 1401 1888 1423
rect 1854 1355 1888 1363
rect 1854 1329 1888 1355
rect 1854 1287 1888 1291
rect 1854 1257 1888 1287
rect 1854 1185 1888 1219
rect 1854 1117 1888 1147
rect 1854 1113 1888 1117
rect 1854 1049 1888 1075
rect 1854 1041 1888 1049
rect 1854 981 1888 1003
rect 1854 969 1888 981
rect 1854 913 1888 931
rect 1854 897 1888 913
rect 2127 2019 2161 2053
rect 2127 1947 2161 1981
rect 2488 2015 2489 2041
rect 2489 2015 2522 2041
rect 2488 2007 2522 2015
rect 3520 2037 3530 2065
rect 3530 2037 3554 2065
rect 3520 1997 3554 1999
rect 2488 1947 2489 1969
rect 2489 1947 2522 1969
rect 2751 1955 2758 1983
rect 2758 1955 2785 1983
rect 2850 1955 2853 1983
rect 2853 1955 2884 1983
rect 2948 1955 2982 1983
rect 3070 1955 3104 1983
rect 3168 1955 3199 1983
rect 3199 1955 3202 1983
rect 3267 1955 3294 1983
rect 3294 1955 3301 1983
rect 3520 1965 3530 1997
rect 3530 1965 3554 1997
rect 2751 1949 2785 1955
rect 2850 1949 2884 1955
rect 2948 1949 2982 1955
rect 3070 1949 3104 1955
rect 3168 1949 3202 1955
rect 3267 1949 3301 1955
rect 3957 1956 3991 1967
rect 2488 1935 2522 1947
rect 3957 1933 3984 1956
rect 3984 1933 3991 1956
rect 4029 1933 4063 1967
rect 2697 1839 2731 1873
rect 2131 1808 2165 1820
rect 2131 1786 2165 1808
rect 2131 1740 2165 1748
rect 2131 1714 2165 1740
rect 2131 1672 2165 1676
rect 2131 1642 2165 1672
rect 2131 1570 2165 1604
rect 2131 1502 2165 1532
rect 2131 1498 2165 1502
rect 2131 1434 2165 1460
rect 2131 1426 2165 1434
rect 2131 1366 2165 1388
rect 2131 1354 2165 1366
rect 2131 1298 2165 1316
rect 2131 1282 2165 1298
rect 2287 1808 2321 1820
rect 2287 1786 2321 1808
rect 2287 1740 2321 1748
rect 2287 1714 2321 1740
rect 2287 1672 2321 1676
rect 2287 1642 2321 1672
rect 2287 1570 2321 1604
rect 2287 1502 2321 1532
rect 2287 1498 2321 1502
rect 2287 1434 2321 1460
rect 2287 1426 2321 1434
rect 2287 1366 2321 1388
rect 2287 1354 2321 1366
rect 2287 1298 2321 1316
rect 2287 1282 2321 1298
rect 2414 1808 2448 1820
rect 2414 1786 2448 1808
rect 2414 1740 2448 1748
rect 2414 1714 2448 1740
rect 2414 1672 2448 1676
rect 2414 1642 2448 1672
rect 2414 1570 2448 1604
rect 2414 1502 2448 1532
rect 2414 1498 2448 1502
rect 2414 1434 2448 1460
rect 2414 1426 2448 1434
rect 2414 1366 2448 1388
rect 2414 1354 2448 1366
rect 2414 1298 2448 1316
rect 2414 1282 2448 1298
rect 2570 1808 2604 1820
rect 2570 1786 2604 1808
rect 2570 1740 2604 1748
rect 2570 1714 2604 1740
rect 2570 1672 2604 1676
rect 2570 1642 2604 1672
rect 2570 1570 2604 1604
rect 2570 1502 2604 1532
rect 2570 1498 2604 1502
rect 2570 1434 2604 1460
rect 2570 1426 2604 1434
rect 2570 1366 2604 1388
rect 2570 1354 2604 1366
rect 2570 1298 2604 1316
rect 2570 1282 2604 1298
rect 2697 1769 2731 1801
rect 2697 1767 2731 1769
rect 2697 1701 2731 1729
rect 2697 1695 2731 1701
rect 2697 1633 2731 1657
rect 2697 1623 2731 1633
rect 2697 1565 2731 1585
rect 2697 1551 2731 1565
rect 2697 1497 2731 1513
rect 2697 1479 2731 1497
rect 2697 1429 2731 1441
rect 2697 1407 2731 1429
rect 2697 1361 2731 1369
rect 2697 1335 2731 1361
rect 2697 1293 2731 1297
rect 2697 1263 2731 1293
rect 2697 1191 2731 1225
rect 2697 1123 2731 1153
rect 2697 1119 2731 1123
rect 2697 1055 2731 1081
rect 2697 1047 2731 1055
rect 2697 987 2731 1009
rect 2697 975 2731 987
rect 2697 919 2731 937
rect 2697 903 2731 919
rect 2853 1839 2887 1873
rect 2853 1769 2887 1801
rect 2853 1767 2887 1769
rect 2853 1701 2887 1729
rect 2853 1695 2887 1701
rect 2853 1633 2887 1657
rect 2853 1623 2887 1633
rect 2853 1565 2887 1585
rect 2853 1551 2887 1565
rect 2853 1497 2887 1513
rect 2853 1479 2887 1497
rect 2853 1429 2887 1441
rect 2853 1407 2887 1429
rect 2853 1361 2887 1369
rect 2853 1335 2887 1361
rect 2853 1293 2887 1297
rect 2853 1263 2887 1293
rect 2853 1191 2887 1225
rect 2853 1123 2887 1153
rect 2853 1119 2887 1123
rect 2853 1055 2887 1081
rect 2853 1047 2887 1055
rect 2853 987 2887 1009
rect 2853 975 2887 987
rect 2853 919 2887 937
rect 2853 903 2887 919
rect 3009 1839 3043 1873
rect 3009 1769 3043 1801
rect 3009 1767 3043 1769
rect 3009 1701 3043 1729
rect 3009 1695 3043 1701
rect 3009 1633 3043 1657
rect 3009 1623 3043 1633
rect 3009 1565 3043 1585
rect 3009 1551 3043 1565
rect 3009 1497 3043 1513
rect 3009 1479 3043 1497
rect 3009 1429 3043 1441
rect 3009 1407 3043 1429
rect 3009 1361 3043 1369
rect 3009 1335 3043 1361
rect 3009 1293 3043 1297
rect 3009 1263 3043 1293
rect 3009 1191 3043 1225
rect 3009 1123 3043 1153
rect 3009 1119 3043 1123
rect 3009 1055 3043 1081
rect 3009 1047 3043 1055
rect 3009 987 3043 1009
rect 3009 975 3043 987
rect 3009 919 3043 937
rect 3009 903 3043 919
rect 3165 1839 3199 1873
rect 3165 1769 3199 1801
rect 3165 1767 3199 1769
rect 3165 1701 3199 1729
rect 3165 1695 3199 1701
rect 3165 1633 3199 1657
rect 3165 1623 3199 1633
rect 3165 1565 3199 1585
rect 3165 1551 3199 1565
rect 3165 1497 3199 1513
rect 3165 1479 3199 1497
rect 3165 1429 3199 1441
rect 3165 1407 3199 1429
rect 3165 1361 3199 1369
rect 3165 1335 3199 1361
rect 3165 1293 3199 1297
rect 3165 1263 3199 1293
rect 3165 1191 3199 1225
rect 3165 1123 3199 1153
rect 3165 1119 3199 1123
rect 3165 1055 3199 1081
rect 3165 1047 3199 1055
rect 3165 987 3199 1009
rect 3165 975 3199 987
rect 3165 919 3199 937
rect 3165 903 3199 919
rect 3321 1839 3355 1873
rect 3321 1769 3355 1801
rect 3321 1767 3355 1769
rect 3321 1701 3355 1729
rect 3321 1695 3355 1701
rect 3321 1633 3355 1657
rect 3321 1623 3355 1633
rect 3321 1565 3355 1585
rect 3321 1551 3355 1565
rect 3321 1497 3355 1513
rect 3321 1479 3355 1497
rect 3321 1429 3355 1441
rect 3321 1407 3355 1429
rect 3321 1361 3355 1369
rect 3321 1335 3355 1361
rect 3446 1823 3480 1835
rect 3446 1801 3480 1823
rect 3446 1755 3480 1763
rect 3446 1729 3480 1755
rect 3446 1687 3480 1691
rect 3446 1657 3480 1687
rect 3446 1585 3480 1619
rect 3446 1517 3480 1547
rect 3446 1513 3480 1517
rect 3446 1449 3480 1475
rect 3446 1441 3480 1449
rect 3446 1381 3480 1403
rect 3446 1369 3480 1381
rect 3446 1313 3480 1331
rect 3446 1297 3480 1313
rect 3602 1823 3636 1835
rect 3602 1801 3636 1823
rect 3602 1755 3636 1763
rect 3602 1729 3636 1755
rect 3602 1687 3636 1691
rect 3602 1657 3636 1687
rect 3889 1807 3923 1833
rect 3889 1799 3923 1807
rect 3889 1739 3923 1761
rect 3889 1727 3923 1739
rect 3889 1671 3923 1689
rect 3889 1655 3923 1671
rect 4125 1807 4159 1833
rect 4125 1799 4159 1807
rect 4125 1739 4159 1761
rect 4125 1727 4159 1739
rect 4125 1671 4159 1689
rect 4125 1655 4159 1671
rect 3602 1585 3636 1619
rect 3602 1517 3636 1547
rect 3602 1513 3636 1517
rect 3602 1449 3636 1475
rect 3602 1441 3636 1449
rect 3602 1381 3636 1403
rect 3602 1369 3636 1381
rect 3602 1313 3636 1331
rect 3602 1297 3636 1313
rect 3321 1293 3355 1297
rect 3321 1263 3355 1293
rect 3321 1191 3355 1225
rect 3321 1123 3355 1153
rect 3321 1119 3355 1123
rect 3321 1055 3355 1081
rect 3321 1047 3355 1055
rect 3321 987 3355 1009
rect 3321 975 3355 987
rect 3321 919 3355 937
rect 3321 903 3355 919
rect 3706 1048 3740 1082
rect 3802 1048 3836 1082
rect 3898 1048 3932 1082
rect 3706 972 3740 1006
rect 3802 972 3836 1006
rect 3898 972 3932 1006
rect 3706 896 3740 930
rect 3802 896 3836 930
rect 3898 896 3932 930
rect 150 827 184 832
rect 223 827 257 832
rect 296 827 330 832
rect 369 827 403 832
rect 441 827 475 832
rect 513 827 547 832
rect 585 827 619 832
rect 657 827 691 832
rect 729 827 763 832
rect 801 827 835 832
rect 873 827 907 832
rect 945 827 979 832
rect 1017 827 1051 832
rect 1089 827 1123 832
rect 1161 827 1195 832
rect 1233 827 1267 832
rect 1305 827 1339 832
rect 1377 827 1411 832
rect 1449 827 1483 832
rect 1521 827 1555 832
rect 1593 827 1627 832
rect 1665 827 1699 832
rect 1737 827 1771 832
rect 1809 827 1843 832
rect 1881 827 1915 832
rect 1953 827 1987 832
rect 2025 827 2059 832
rect 2097 827 2131 832
rect 2169 827 2203 832
rect 2241 827 2275 832
rect 2313 827 2347 832
rect 2385 827 2419 832
rect 2457 827 2491 832
rect 2529 827 2563 832
rect 2601 827 2635 832
rect 2673 827 2707 832
rect 2745 827 2779 832
rect 2817 827 2851 832
rect 2889 827 2923 832
rect 2961 827 2995 832
rect 3033 827 3067 832
rect 3105 827 3139 832
rect 3177 827 3211 832
rect 3249 827 3283 832
rect 3321 827 3355 832
rect 150 798 168 827
rect 168 798 184 827
rect 223 798 237 827
rect 237 798 257 827
rect 296 798 306 827
rect 306 798 330 827
rect 369 798 375 827
rect 375 798 403 827
rect 441 798 444 827
rect 444 798 475 827
rect 513 798 547 827
rect 585 798 616 827
rect 616 798 619 827
rect 657 798 685 827
rect 685 798 691 827
rect 729 798 754 827
rect 754 798 763 827
rect 801 798 823 827
rect 823 798 835 827
rect 873 798 892 827
rect 892 798 907 827
rect 945 798 961 827
rect 961 798 979 827
rect 1017 798 1030 827
rect 1030 798 1051 827
rect 1089 798 1099 827
rect 1099 798 1123 827
rect 1161 798 1168 827
rect 1168 798 1195 827
rect 1233 798 1237 827
rect 1237 798 1267 827
rect 1305 798 1306 827
rect 1306 798 1339 827
rect 1377 798 1410 827
rect 1410 798 1411 827
rect 1449 798 1479 827
rect 1479 798 1483 827
rect 1521 798 1548 827
rect 1548 798 1555 827
rect 1593 798 1617 827
rect 1617 798 1627 827
rect 1665 798 1686 827
rect 1686 798 1699 827
rect 1737 798 1755 827
rect 1755 798 1771 827
rect 1809 798 1824 827
rect 1824 798 1843 827
rect 1881 798 1893 827
rect 1893 798 1915 827
rect 1953 798 1962 827
rect 1962 798 1987 827
rect 2025 798 2031 827
rect 2031 798 2059 827
rect 2097 798 2100 827
rect 2100 798 2131 827
rect 2169 798 2203 827
rect 2241 798 2272 827
rect 2272 798 2275 827
rect 2313 798 2341 827
rect 2341 798 2347 827
rect 2385 798 2410 827
rect 2410 798 2419 827
rect 2457 798 2479 827
rect 2479 798 2491 827
rect 2529 798 2548 827
rect 2548 798 2563 827
rect 2601 798 2617 827
rect 2617 798 2635 827
rect 2673 798 2686 827
rect 2686 798 2707 827
rect 2745 798 2755 827
rect 2755 798 2779 827
rect 2817 798 2824 827
rect 2824 798 2851 827
rect 2889 798 2893 827
rect 2893 798 2923 827
rect 2961 798 2962 827
rect 2962 798 2995 827
rect 3033 798 3064 827
rect 3064 798 3067 827
rect 3105 798 3132 827
rect 3132 798 3139 827
rect 3177 798 3200 827
rect 3200 798 3211 827
rect 3249 798 3268 827
rect 3268 798 3283 827
rect 3321 798 3336 827
rect 3336 798 3355 827
rect 3706 820 3740 854
rect 3802 820 3836 854
rect 3898 820 3932 854
rect 3706 744 3740 778
rect 3802 744 3836 778
rect 3898 744 3932 778
rect 3318 704 3352 738
rect 3400 704 3434 738
rect 3482 704 3516 738
rect 169 640 193 674
rect 193 640 203 674
rect 241 640 261 674
rect 261 640 275 674
rect 313 640 329 674
rect 329 640 347 674
rect 385 640 397 674
rect 397 640 419 674
rect 457 640 465 674
rect 465 640 491 674
rect 529 640 533 674
rect 533 640 563 674
rect 601 640 635 674
rect 673 640 703 674
rect 703 640 707 674
rect 745 640 771 674
rect 771 640 779 674
rect 817 640 839 674
rect 839 640 851 674
rect 889 640 907 674
rect 907 640 923 674
rect 961 640 975 674
rect 975 640 995 674
rect 1033 640 1043 674
rect 1043 640 1067 674
rect 1105 640 1111 674
rect 1111 640 1139 674
rect 1177 640 1179 674
rect 1179 640 1211 674
rect 1249 640 1281 674
rect 1281 640 1283 674
rect 1321 640 1349 674
rect 1349 640 1355 674
rect 1393 640 1417 674
rect 1417 640 1427 674
rect 1465 640 1485 674
rect 1485 640 1499 674
rect 1537 640 1553 674
rect 1553 640 1571 674
rect 1609 640 1621 674
rect 1621 640 1643 674
rect 1681 640 1689 674
rect 1689 640 1715 674
rect 1753 640 1757 674
rect 1757 640 1787 674
rect 1825 640 1859 674
rect 1897 640 1927 674
rect 1927 640 1931 674
rect 1969 640 1995 674
rect 1995 640 2003 674
rect 2041 640 2063 674
rect 2063 640 2075 674
rect 2113 640 2131 674
rect 2131 640 2147 674
rect 2697 667 2731 683
rect 2697 649 2731 667
rect 2192 578 2225 612
rect 2225 578 2226 612
rect 2192 506 2226 540
rect 2697 599 2731 611
rect 2697 577 2731 599
rect 2697 531 2731 539
rect 2697 505 2731 531
rect 2853 667 2887 683
rect 2853 649 2887 667
rect 2853 599 2887 611
rect 2853 577 2887 599
rect 2853 531 2887 539
rect 2853 505 2887 531
rect 3009 667 3043 683
rect 3009 649 3043 667
rect 3009 599 3043 611
rect 3009 577 3043 599
rect 3009 531 3043 539
rect 3009 505 3043 531
rect 3165 667 3199 683
rect 3165 649 3199 667
rect 3165 599 3199 611
rect 3165 577 3199 599
rect 3165 531 3199 539
rect 3165 505 3199 531
rect 3318 601 3352 635
rect 3400 601 3434 635
rect 3482 601 3516 635
rect 3318 499 3352 533
rect 3400 499 3434 533
rect 3482 499 3516 533
rect 169 404 193 438
rect 193 404 203 438
rect 241 404 261 438
rect 261 404 275 438
rect 313 404 329 438
rect 329 404 347 438
rect 385 404 397 438
rect 397 404 419 438
rect 457 404 465 438
rect 465 404 491 438
rect 529 404 533 438
rect 533 404 563 438
rect 601 404 635 438
rect 673 404 703 438
rect 703 404 707 438
rect 745 404 771 438
rect 771 404 779 438
rect 817 404 839 438
rect 839 404 851 438
rect 889 404 907 438
rect 907 404 923 438
rect 961 404 975 438
rect 975 404 995 438
rect 1033 404 1043 438
rect 1043 404 1067 438
rect 1105 404 1111 438
rect 1111 404 1139 438
rect 1177 404 1179 438
rect 1179 404 1211 438
rect 1249 404 1281 438
rect 1281 404 1283 438
rect 1321 404 1349 438
rect 1349 404 1355 438
rect 1393 404 1417 438
rect 1417 404 1427 438
rect 1465 404 1485 438
rect 1485 404 1499 438
rect 1537 404 1553 438
rect 1553 404 1571 438
rect 1609 404 1621 438
rect 1621 404 1643 438
rect 1681 404 1689 438
rect 1689 404 1715 438
rect 1753 404 1757 438
rect 1757 404 1787 438
rect 1825 404 1859 438
rect 1897 404 1927 438
rect 1927 404 1931 438
rect 1969 404 1995 438
rect 1995 404 2003 438
rect 2041 404 2063 438
rect 2063 404 2075 438
rect 2113 404 2131 438
rect 2131 404 2147 438
rect 2765 397 2792 431
rect 2792 397 2799 431
rect 2847 397 2862 431
rect 2862 397 2881 431
rect 2929 397 2931 431
rect 2931 397 2963 431
rect 3010 397 3035 431
rect 3035 397 3044 431
rect 3091 397 3104 431
rect 3104 397 3125 431
rect 169 277 193 311
rect 193 277 203 311
rect 241 277 261 311
rect 261 277 275 311
rect 313 277 329 311
rect 329 277 347 311
rect 385 277 397 311
rect 397 277 419 311
rect 457 277 465 311
rect 465 277 491 311
rect 529 277 533 311
rect 533 277 563 311
rect 601 277 635 311
rect 673 277 703 311
rect 703 277 707 311
rect 745 277 771 311
rect 771 277 779 311
rect 817 277 839 311
rect 839 277 851 311
rect 889 277 907 311
rect 907 277 923 311
rect 961 277 975 311
rect 975 277 995 311
rect 1033 277 1043 311
rect 1043 277 1067 311
rect 1105 277 1111 311
rect 1111 277 1139 311
rect 1177 277 1179 311
rect 1179 277 1211 311
rect 1249 277 1281 311
rect 1281 277 1283 311
rect 1321 277 1349 311
rect 1349 277 1355 311
rect 1393 277 1417 311
rect 1417 277 1427 311
rect 1465 277 1485 311
rect 1485 277 1499 311
rect 1537 277 1553 311
rect 1553 277 1571 311
rect 1609 277 1621 311
rect 1621 277 1643 311
rect 1681 277 1689 311
rect 1689 277 1715 311
rect 1753 277 1757 311
rect 1757 277 1787 311
rect 1825 277 1859 311
rect 1897 277 1927 311
rect 1927 277 1931 311
rect 1969 277 1995 311
rect 1995 277 2003 311
rect 2041 277 2063 311
rect 2063 277 2075 311
rect 2113 277 2131 311
rect 2131 277 2147 311
rect 2192 174 2226 208
rect 2192 102 2225 136
rect 2225 102 2226 136
rect 169 41 193 75
rect 193 41 203 75
rect 241 41 261 75
rect 261 41 275 75
rect 313 41 329 75
rect 329 41 347 75
rect 385 41 397 75
rect 397 41 419 75
rect 457 41 465 75
rect 465 41 491 75
rect 529 41 533 75
rect 533 41 563 75
rect 601 41 635 75
rect 673 41 703 75
rect 703 41 707 75
rect 745 41 771 75
rect 771 41 779 75
rect 817 41 839 75
rect 839 41 851 75
rect 889 41 907 75
rect 907 41 923 75
rect 961 41 975 75
rect 975 41 995 75
rect 1033 41 1043 75
rect 1043 41 1067 75
rect 1105 41 1111 75
rect 1111 41 1139 75
rect 1177 41 1179 75
rect 1179 41 1211 75
rect 1249 41 1281 75
rect 1281 41 1283 75
rect 1321 41 1349 75
rect 1349 41 1355 75
rect 1393 41 1417 75
rect 1417 41 1427 75
rect 1465 41 1485 75
rect 1485 41 1499 75
rect 1537 41 1553 75
rect 1553 41 1571 75
rect 1609 41 1621 75
rect 1621 41 1643 75
rect 1681 41 1689 75
rect 1689 41 1715 75
rect 1753 41 1757 75
rect 1757 41 1787 75
rect 1825 41 1859 75
rect 1897 41 1927 75
rect 1927 41 1931 75
rect 1969 41 1995 75
rect 1995 41 2003 75
rect 2041 41 2063 75
rect 2063 41 2075 75
rect 2113 41 2131 75
rect 2131 41 2147 75
rect -11540 -8659 -11506 -8658
rect -11540 -8692 -11516 -8659
rect -11516 -8692 -11506 -8659
rect -11540 -8761 -11516 -8730
rect -11516 -8761 -11506 -8730
rect -11540 -8764 -11506 -8761
rect -29046 -8875 -29012 -8847
rect -28958 -8875 -28924 -8847
rect -28870 -8875 -28836 -8847
rect -28189 -8870 -28155 -8847
rect -28115 -8870 -28081 -8847
rect -28041 -8870 -28007 -8847
rect -27967 -8870 -27933 -8847
rect -27893 -8870 -27859 -8847
rect -27819 -8870 -27785 -8847
rect -27745 -8870 -27711 -8847
rect -27671 -8870 -27637 -8847
rect -27597 -8870 -27563 -8847
rect -27523 -8870 -27489 -8847
rect -27449 -8870 -27415 -8847
rect -27375 -8870 -27341 -8847
rect -27301 -8870 -27267 -8847
rect -27227 -8870 -27193 -8847
rect -27153 -8870 -27119 -8847
rect -32338 -9600 -32315 -8918
rect -32315 -9600 -31669 -8918
rect -31669 -9598 -31632 -8918
rect -31632 -9598 -30792 -8918
rect -30753 -8952 -30719 -8918
rect -30680 -8952 -30646 -8918
rect -30607 -8952 -30573 -8918
rect -30534 -8952 -30500 -8918
rect -30461 -8952 -30427 -8918
rect -30388 -8952 -30354 -8918
rect -30315 -8952 -30281 -8918
rect -30242 -8952 -30208 -8918
rect -30169 -8952 -30135 -8918
rect -30096 -8952 -30062 -8918
rect -30023 -8952 -29989 -8918
rect -29950 -8952 -29916 -8918
rect -29877 -8952 -29843 -8918
rect -29804 -8952 -29770 -8918
rect -29731 -8952 -29697 -8918
rect -29658 -8952 -29624 -8918
rect -29585 -8952 -29551 -8918
rect -29512 -8952 -29478 -8918
rect -29439 -8952 -29405 -8918
rect -29366 -8952 -29332 -8918
rect -29293 -8952 -29259 -8918
rect -29220 -8952 -29186 -8918
rect -29134 -8947 -29100 -8913
rect -29046 -8947 -29012 -8913
rect -28958 -8947 -28924 -8913
rect -28870 -8947 -28836 -8913
rect -28189 -8942 -28155 -8908
rect -28115 -8942 -28081 -8908
rect -28041 -8942 -28007 -8908
rect -27967 -8942 -27933 -8908
rect -27893 -8942 -27859 -8908
rect -27819 -8942 -27785 -8908
rect -27745 -8942 -27711 -8908
rect -27671 -8942 -27637 -8908
rect -27597 -8942 -27563 -8908
rect -27523 -8942 -27489 -8908
rect -27449 -8942 -27415 -8908
rect -27375 -8918 -27346 -8908
rect -27346 -8918 -27341 -8908
rect -27301 -8918 -27277 -8908
rect -27277 -8918 -27267 -8908
rect -27227 -8918 -27208 -8908
rect -27208 -8918 -27193 -8908
rect -27153 -8918 -27139 -8908
rect -27139 -8918 -27119 -8908
rect -27375 -8942 -27341 -8918
rect -27301 -8942 -27267 -8918
rect -27227 -8942 -27193 -8918
rect -27153 -8942 -27119 -8918
rect -30753 -9024 -30719 -8990
rect -30680 -9024 -30646 -8990
rect -30607 -9024 -30573 -8990
rect -30534 -9024 -30500 -8990
rect -30461 -9024 -30427 -8990
rect -30388 -9024 -30354 -8990
rect -30315 -9024 -30281 -8990
rect -30242 -9024 -30208 -8990
rect -30169 -9024 -30135 -8990
rect -30096 -9024 -30062 -8990
rect -30023 -9024 -29989 -8990
rect -29950 -9024 -29916 -8990
rect -29877 -9024 -29843 -8990
rect -29804 -9024 -29770 -8990
rect -29731 -9024 -29697 -8990
rect -29658 -9024 -29624 -8990
rect -29585 -9024 -29551 -8990
rect -29512 -9024 -29478 -8990
rect -29439 -9024 -29405 -8990
rect -29366 -9024 -29332 -8990
rect -29293 -9024 -29259 -8990
rect -29220 -9024 -29186 -8990
rect -29134 -9019 -29100 -8985
rect -29046 -9019 -29012 -8985
rect -28958 -9019 -28924 -8985
rect -28870 -9019 -28836 -8985
rect -28189 -9014 -28155 -8980
rect -28115 -9014 -28081 -8980
rect -28041 -9014 -28007 -8980
rect -27967 -9014 -27933 -8980
rect -27893 -9014 -27859 -8980
rect -27819 -9014 -27785 -8980
rect -27745 -9014 -27711 -8980
rect -27671 -9014 -27637 -8980
rect -27597 -9014 -27563 -8980
rect -27523 -9014 -27489 -8980
rect -27449 -9014 -27415 -8980
rect -27375 -8986 -27346 -8980
rect -27346 -8986 -27341 -8980
rect -27301 -8986 -27277 -8980
rect -27277 -8986 -27267 -8980
rect -27227 -8986 -27208 -8980
rect -27208 -8986 -27193 -8980
rect -27153 -8986 -27139 -8980
rect -27139 -8986 -27119 -8980
rect -27375 -9014 -27341 -8986
rect -27301 -9014 -27267 -8986
rect -27227 -9014 -27193 -8986
rect -27153 -9014 -27119 -8986
rect -30753 -9096 -30719 -9062
rect -30680 -9096 -30646 -9062
rect -30607 -9096 -30573 -9062
rect -30534 -9096 -30500 -9062
rect -30461 -9096 -30427 -9062
rect -30388 -9096 -30354 -9062
rect -30315 -9096 -30281 -9062
rect -30242 -9096 -30208 -9062
rect -30169 -9096 -30135 -9062
rect -30096 -9096 -30062 -9062
rect -30023 -9096 -29989 -9062
rect -29950 -9096 -29916 -9062
rect -29877 -9096 -29843 -9062
rect -29804 -9096 -29770 -9062
rect -29731 -9096 -29697 -9062
rect -29658 -9096 -29624 -9062
rect -29585 -9096 -29551 -9062
rect -29512 -9096 -29478 -9062
rect -29439 -9096 -29405 -9062
rect -29366 -9096 -29332 -9062
rect -29293 -9096 -29259 -9062
rect -29220 -9096 -29186 -9062
rect -29134 -9091 -29100 -9057
rect -29046 -9091 -29012 -9057
rect -28958 -9091 -28924 -9057
rect -28870 -9091 -28836 -9057
rect -28189 -9086 -28155 -9052
rect -28115 -9086 -28081 -9052
rect -28041 -9086 -28007 -9052
rect -27967 -9086 -27933 -9052
rect -27893 -9086 -27859 -9052
rect -27819 -9086 -27785 -9052
rect -27745 -9086 -27711 -9052
rect -27671 -9086 -27637 -9052
rect -27597 -9086 -27563 -9052
rect -27523 -9086 -27489 -9052
rect -27449 -9086 -27415 -9052
rect -27375 -9054 -27346 -9052
rect -27346 -9054 -27341 -9052
rect -27301 -9054 -27277 -9052
rect -27277 -9054 -27267 -9052
rect -27227 -9054 -27208 -9052
rect -27208 -9054 -27193 -9052
rect -27153 -9054 -27139 -9052
rect -27139 -9054 -27119 -9052
rect -27375 -9086 -27341 -9054
rect -27301 -9086 -27267 -9054
rect -27227 -9086 -27193 -9054
rect -27153 -9086 -27119 -9054
rect -30753 -9168 -30719 -9134
rect -30680 -9168 -30646 -9134
rect -30607 -9168 -30573 -9134
rect -30534 -9168 -30500 -9134
rect -30461 -9168 -30427 -9134
rect -30388 -9168 -30354 -9134
rect -30315 -9168 -30281 -9134
rect -30242 -9168 -30208 -9134
rect -30169 -9168 -30135 -9134
rect -30096 -9168 -30062 -9134
rect -30023 -9168 -29989 -9134
rect -29950 -9168 -29916 -9134
rect -29877 -9168 -29843 -9134
rect -29804 -9168 -29770 -9134
rect -29731 -9168 -29697 -9134
rect -29658 -9168 -29624 -9134
rect -29585 -9168 -29551 -9134
rect -29512 -9168 -29478 -9134
rect -29439 -9168 -29405 -9134
rect -29366 -9168 -29332 -9134
rect -29293 -9168 -29259 -9134
rect -29220 -9168 -29186 -9134
rect -29134 -9163 -29100 -9129
rect -29046 -9163 -29012 -9129
rect -28958 -9163 -28924 -9129
rect -28870 -9163 -28836 -9129
rect -28189 -9158 -28155 -9124
rect -28115 -9158 -28081 -9124
rect -28041 -9158 -28007 -9124
rect -27967 -9158 -27933 -9124
rect -27893 -9158 -27859 -9124
rect -27819 -9158 -27785 -9124
rect -27745 -9158 -27711 -9124
rect -27671 -9158 -27637 -9124
rect -27597 -9158 -27563 -9124
rect -27523 -9158 -27489 -9124
rect -27449 -9158 -27415 -9124
rect -27375 -9156 -27341 -9124
rect -27301 -9156 -27267 -9124
rect -27227 -9156 -27193 -9124
rect -27153 -9156 -27119 -9124
rect -27375 -9158 -27346 -9156
rect -27346 -9158 -27341 -9156
rect -27301 -9158 -27277 -9156
rect -27277 -9158 -27267 -9156
rect -27227 -9158 -27208 -9156
rect -27208 -9158 -27193 -9156
rect -27153 -9158 -27139 -9156
rect -27139 -9158 -27119 -9156
rect -30753 -9240 -30719 -9206
rect -30680 -9240 -30646 -9206
rect -30607 -9240 -30573 -9206
rect -30534 -9240 -30500 -9206
rect -30461 -9240 -30427 -9206
rect -30388 -9240 -30354 -9206
rect -30315 -9240 -30281 -9206
rect -30242 -9240 -30208 -9206
rect -30169 -9240 -30135 -9206
rect -30096 -9240 -30062 -9206
rect -30023 -9240 -29989 -9206
rect -29950 -9240 -29916 -9206
rect -29877 -9240 -29843 -9206
rect -29804 -9240 -29770 -9206
rect -29731 -9240 -29697 -9206
rect -29658 -9240 -29624 -9206
rect -29585 -9240 -29551 -9206
rect -29512 -9240 -29478 -9206
rect -29439 -9240 -29405 -9206
rect -29366 -9240 -29332 -9206
rect -29293 -9240 -29259 -9206
rect -29220 -9240 -29186 -9206
rect -29134 -9235 -29100 -9201
rect -29046 -9235 -29012 -9201
rect -28958 -9235 -28924 -9201
rect -28870 -9235 -28836 -9201
rect -28189 -9230 -28155 -9196
rect -28115 -9230 -28081 -9196
rect -28041 -9230 -28007 -9196
rect -27967 -9230 -27933 -9196
rect -27893 -9230 -27859 -9196
rect -27819 -9230 -27785 -9196
rect -27745 -9230 -27711 -9196
rect -27671 -9230 -27637 -9196
rect -27597 -9230 -27563 -9196
rect -27523 -9230 -27489 -9196
rect -27449 -9230 -27415 -9196
rect -27375 -9224 -27341 -9196
rect -27301 -9224 -27267 -9196
rect -27227 -9224 -27193 -9196
rect -27153 -9224 -27119 -9196
rect -27375 -9230 -27346 -9224
rect -27346 -9230 -27341 -9224
rect -27301 -9230 -27277 -9224
rect -27277 -9230 -27267 -9224
rect -27227 -9230 -27208 -9224
rect -27208 -9230 -27193 -9224
rect -27153 -9230 -27139 -9224
rect -27139 -9230 -27119 -9224
rect -30753 -9312 -30719 -9278
rect -30680 -9312 -30646 -9278
rect -30607 -9312 -30573 -9278
rect -30534 -9312 -30500 -9278
rect -30461 -9312 -30427 -9278
rect -30388 -9312 -30354 -9278
rect -30315 -9312 -30281 -9278
rect -30242 -9312 -30208 -9278
rect -30169 -9312 -30135 -9278
rect -30096 -9312 -30062 -9278
rect -30023 -9312 -29989 -9278
rect -29950 -9312 -29916 -9278
rect -29877 -9312 -29843 -9278
rect -29804 -9312 -29770 -9278
rect -29731 -9312 -29697 -9278
rect -29658 -9312 -29624 -9278
rect -29585 -9312 -29551 -9278
rect -29512 -9312 -29478 -9278
rect -29439 -9312 -29405 -9278
rect -29366 -9312 -29332 -9278
rect -29293 -9312 -29259 -9278
rect -29220 -9312 -29186 -9278
rect -29134 -9307 -29100 -9273
rect -29046 -9307 -29012 -9273
rect -28958 -9307 -28924 -9273
rect -28870 -9307 -28836 -9273
rect -28189 -9302 -28155 -9268
rect -28115 -9302 -28081 -9268
rect -28041 -9302 -28007 -9268
rect -27967 -9302 -27933 -9268
rect -27893 -9302 -27859 -9268
rect -27819 -9302 -27785 -9268
rect -27745 -9302 -27711 -9268
rect -27671 -9302 -27637 -9268
rect -27597 -9302 -27563 -9268
rect -27523 -9302 -27489 -9268
rect -27449 -9302 -27415 -9268
rect -27375 -9292 -27341 -9268
rect -27301 -9292 -27267 -9268
rect -27227 -9292 -27193 -9268
rect -27153 -9292 -27119 -9268
rect -27375 -9302 -27346 -9292
rect -27346 -9302 -27341 -9292
rect -27301 -9302 -27277 -9292
rect -27277 -9302 -27267 -9292
rect -27227 -9302 -27208 -9292
rect -27208 -9302 -27193 -9292
rect -27153 -9302 -27139 -9292
rect -27139 -9302 -27119 -9292
rect -30753 -9384 -30719 -9350
rect -30680 -9384 -30646 -9350
rect -30607 -9384 -30573 -9350
rect -30534 -9384 -30500 -9350
rect -30461 -9384 -30427 -9350
rect -30388 -9384 -30354 -9350
rect -30315 -9384 -30281 -9350
rect -30242 -9384 -30208 -9350
rect -30169 -9384 -30135 -9350
rect -30096 -9384 -30062 -9350
rect -30023 -9384 -29989 -9350
rect -29950 -9384 -29916 -9350
rect -29877 -9384 -29843 -9350
rect -29804 -9384 -29770 -9350
rect -29731 -9384 -29697 -9350
rect -29658 -9384 -29624 -9350
rect -29585 -9384 -29551 -9350
rect -29512 -9384 -29478 -9350
rect -29439 -9384 -29405 -9350
rect -29366 -9384 -29332 -9350
rect -29293 -9384 -29259 -9350
rect -29220 -9384 -29186 -9350
rect -29134 -9379 -29100 -9345
rect -29046 -9379 -29012 -9345
rect -28958 -9379 -28924 -9345
rect -28870 -9379 -28836 -9345
rect -28189 -9374 -28155 -9340
rect -28115 -9374 -28081 -9340
rect -28041 -9374 -28007 -9340
rect -27967 -9374 -27933 -9340
rect -27893 -9374 -27859 -9340
rect -27819 -9374 -27785 -9340
rect -27745 -9374 -27711 -9340
rect -27671 -9374 -27637 -9340
rect -27597 -9374 -27563 -9340
rect -27523 -9374 -27489 -9340
rect -27449 -9374 -27415 -9340
rect -27375 -9360 -27341 -9340
rect -27301 -9360 -27267 -9340
rect -27227 -9360 -27193 -9340
rect -27153 -9360 -27119 -9340
rect -27375 -9374 -27346 -9360
rect -27346 -9374 -27341 -9360
rect -27301 -9374 -27277 -9360
rect -27277 -9374 -27267 -9360
rect -27227 -9374 -27208 -9360
rect -27208 -9374 -27193 -9360
rect -27153 -9374 -27139 -9360
rect -27139 -9374 -27119 -9360
rect -30753 -9456 -30719 -9422
rect -30680 -9456 -30646 -9422
rect -30607 -9456 -30573 -9422
rect -30534 -9456 -30500 -9422
rect -30461 -9456 -30427 -9422
rect -30388 -9456 -30354 -9422
rect -30315 -9456 -30281 -9422
rect -30242 -9456 -30208 -9422
rect -30169 -9456 -30135 -9422
rect -30096 -9456 -30062 -9422
rect -30023 -9456 -29989 -9422
rect -29950 -9456 -29916 -9422
rect -29877 -9456 -29843 -9422
rect -29804 -9456 -29770 -9422
rect -29731 -9456 -29697 -9422
rect -29658 -9456 -29624 -9422
rect -29585 -9456 -29551 -9422
rect -29512 -9456 -29478 -9422
rect -29439 -9456 -29405 -9422
rect -29366 -9456 -29332 -9422
rect -29293 -9456 -29259 -9422
rect -29220 -9456 -29186 -9422
rect -29134 -9451 -29100 -9417
rect -29046 -9451 -29012 -9417
rect -28958 -9451 -28924 -9417
rect -28870 -9451 -28836 -9417
rect -30753 -9528 -30719 -9494
rect -30680 -9528 -30646 -9494
rect -30607 -9528 -30573 -9494
rect -30534 -9528 -30500 -9494
rect -30461 -9528 -30427 -9494
rect -30388 -9528 -30354 -9494
rect -30315 -9528 -30281 -9494
rect -30242 -9528 -30208 -9494
rect -30169 -9528 -30135 -9494
rect -30096 -9528 -30062 -9494
rect -30023 -9528 -29989 -9494
rect -29950 -9528 -29916 -9494
rect -29877 -9528 -29843 -9494
rect -29804 -9528 -29770 -9494
rect -29731 -9528 -29697 -9494
rect -29658 -9528 -29624 -9494
rect -29585 -9528 -29551 -9494
rect -29512 -9528 -29478 -9494
rect -29439 -9528 -29405 -9494
rect -29366 -9528 -29332 -9494
rect -29293 -9528 -29259 -9494
rect -29220 -9528 -29186 -9494
rect -29134 -9523 -29100 -9489
rect -29046 -9523 -29012 -9489
rect -28958 -9523 -28924 -9489
rect -28870 -9523 -28836 -9489
rect -30753 -9598 -30719 -9566
rect -30680 -9598 -30646 -9566
rect -30607 -9598 -30573 -9566
rect -30534 -9598 -30500 -9566
rect -30461 -9598 -30427 -9566
rect -30388 -9598 -30354 -9566
rect -30315 -9598 -30281 -9566
rect -30242 -9598 -30208 -9566
rect -30169 -9598 -30135 -9566
rect -30096 -9598 -30062 -9566
rect -30023 -9598 -29989 -9566
rect -29950 -9598 -29916 -9566
rect -29877 -9598 -29843 -9566
rect -29804 -9598 -29770 -9566
rect -29731 -9598 -29697 -9566
rect -29658 -9598 -29624 -9566
rect -29585 -9598 -29551 -9566
rect -29512 -9598 -29478 -9566
rect -29439 -9598 -29405 -9566
rect -29366 -9598 -29332 -9566
rect -29293 -9598 -29259 -9566
rect -29220 -9598 -29186 -9566
rect -29134 -9595 -29100 -9561
rect -29046 -9595 -29012 -9561
rect -28958 -9595 -28924 -9561
rect -28870 -9595 -28836 -9561
rect -31669 -9600 -30792 -9598
rect -30753 -9600 -30719 -9598
rect -30680 -9600 -30646 -9598
rect -30607 -9600 -30573 -9598
rect -30534 -9600 -30500 -9598
rect -30461 -9600 -30427 -9598
rect -30388 -9600 -30354 -9598
rect -30315 -9600 -30281 -9598
rect -30242 -9600 -30208 -9598
rect -30169 -9600 -30135 -9598
rect -30096 -9600 -30062 -9598
rect -30023 -9600 -29989 -9598
rect -29950 -9600 -29916 -9598
rect -29877 -9600 -29843 -9598
rect -29804 -9600 -29770 -9598
rect -29731 -9600 -29697 -9598
rect -29658 -9600 -29624 -9598
rect -29585 -9600 -29551 -9598
rect -29512 -9600 -29478 -9598
rect -29439 -9600 -29405 -9598
rect -29366 -9600 -29332 -9598
rect -29293 -9600 -29259 -9598
rect -29220 -9600 -29186 -9598
<< metal1 >>
rect -28202 4843 -28196 4895
rect -28144 4843 -28132 4895
rect -28080 4843 -28068 4895
rect -28016 4843 -28004 4895
rect -27952 4843 -27940 4895
rect -27888 4843 -27876 4895
rect -27824 4843 -27812 4895
rect -27760 4843 -27748 4895
rect -27696 4843 -27684 4895
rect -27632 4843 -27620 4895
rect -27568 4843 -27555 4895
rect -27503 4843 -27490 4895
rect -27438 4843 -27425 4895
rect -27373 4843 -27360 4895
rect -27308 4843 -27295 4895
rect -27243 4843 -27230 4895
rect -27178 4843 -27165 4895
rect -27113 4843 -27106 4895
rect -28202 4773 -27106 4843
rect -28202 4721 -28196 4773
rect -28144 4721 -28132 4773
rect -28080 4721 -28068 4773
rect -28016 4721 -28004 4773
rect -27952 4721 -27940 4773
rect -27888 4721 -27876 4773
rect -27824 4721 -27812 4773
rect -27760 4721 -27748 4773
rect -27696 4721 -27684 4773
rect -27632 4721 -27620 4773
rect -27568 4721 -27555 4773
rect -27503 4721 -27490 4773
rect -27438 4721 -27425 4773
rect -27373 4721 -27360 4773
rect -27308 4721 -27295 4773
rect -27243 4721 -27230 4773
rect -27178 4721 -27165 4773
rect -27113 4721 -27106 4773
rect -32350 4333 -28830 4345
rect -32350 4332 -31718 4333
rect -32350 4298 -32344 4332
rect -32310 4298 -32266 4332
rect -32232 4298 -32188 4332
rect -32154 4298 -32110 4332
rect -32076 4298 -32032 4332
rect -31998 4298 -31954 4332
rect -31920 4298 -31876 4332
rect -31842 4298 -31798 4332
rect -31764 4299 -31718 4332
rect -31684 4299 -31645 4333
rect -31611 4299 -31572 4333
rect -31538 4299 -31499 4333
rect -31465 4299 -31426 4333
rect -31392 4299 -31353 4333
rect -31319 4299 -31280 4333
rect -31246 4299 -31207 4333
rect -31173 4299 -31134 4333
rect -31100 4299 -31061 4333
rect -31027 4299 -30988 4333
rect -30954 4299 -30915 4333
rect -30881 4299 -30842 4333
rect -30808 4299 -30768 4333
rect -30734 4299 -30694 4333
rect -30660 4299 -30620 4333
rect -30586 4299 -30546 4333
rect -30512 4299 -30472 4333
rect -30438 4299 -30398 4333
rect -30364 4299 -30324 4333
rect -30290 4299 -30250 4333
rect -30216 4299 -30176 4333
rect -30142 4299 -30102 4333
rect -30068 4299 -30028 4333
rect -29994 4299 -29954 4333
rect -29920 4299 -29880 4333
rect -29846 4299 -29806 4333
rect -29772 4299 -29732 4333
rect -29698 4299 -29658 4333
rect -29624 4299 -29584 4333
rect -29550 4299 -29510 4333
rect -29476 4299 -29436 4333
rect -29402 4299 -29362 4333
rect -29328 4299 -29288 4333
rect -29254 4299 -29214 4333
rect -29180 4299 -29134 4333
rect -29100 4299 -29046 4333
rect -29012 4299 -28958 4333
rect -28924 4299 -28870 4333
rect -28836 4299 -28830 4333
rect -31764 4298 -28830 4299
rect -32350 4261 -28830 4298
rect -32350 4259 -31718 4261
rect -32350 4225 -32344 4259
rect -32310 4225 -32266 4259
rect -32232 4225 -32188 4259
rect -32154 4225 -32110 4259
rect -32076 4225 -32032 4259
rect -31998 4225 -31954 4259
rect -31920 4225 -31876 4259
rect -31842 4225 -31798 4259
rect -31764 4227 -31718 4259
rect -31684 4227 -31645 4261
rect -31611 4227 -31572 4261
rect -31538 4227 -31499 4261
rect -31465 4227 -31426 4261
rect -31392 4227 -31353 4261
rect -31319 4227 -31280 4261
rect -31246 4227 -31207 4261
rect -31173 4227 -31134 4261
rect -31100 4227 -31061 4261
rect -31027 4227 -30988 4261
rect -30954 4227 -30915 4261
rect -30881 4227 -30842 4261
rect -30808 4227 -30768 4261
rect -30734 4227 -30694 4261
rect -30660 4227 -30620 4261
rect -30586 4227 -30546 4261
rect -30512 4227 -30472 4261
rect -30438 4227 -30398 4261
rect -30364 4227 -30324 4261
rect -30290 4227 -30250 4261
rect -30216 4227 -30176 4261
rect -30142 4227 -30102 4261
rect -30068 4227 -30028 4261
rect -29994 4227 -29954 4261
rect -29920 4227 -29880 4261
rect -29846 4227 -29806 4261
rect -29772 4227 -29732 4261
rect -29698 4227 -29658 4261
rect -29624 4227 -29584 4261
rect -29550 4227 -29510 4261
rect -29476 4227 -29436 4261
rect -29402 4227 -29362 4261
rect -29328 4227 -29288 4261
rect -29254 4227 -29214 4261
rect -29180 4260 -28830 4261
rect -29180 4227 -29134 4260
rect -31764 4226 -29134 4227
rect -29100 4226 -29046 4260
rect -29012 4226 -28958 4260
rect -28924 4226 -28870 4260
rect -28836 4226 -28830 4260
rect -31764 4225 -28830 4226
rect -32350 4189 -28830 4225
rect -32350 4186 -31718 4189
rect -32350 4152 -32344 4186
rect -32310 4152 -32266 4186
rect -32232 4152 -32188 4186
rect -32154 4152 -32110 4186
rect -32076 4152 -32032 4186
rect -31998 4152 -31954 4186
rect -31920 4152 -31876 4186
rect -31842 4152 -31798 4186
rect -31764 4155 -31718 4186
rect -31684 4155 -31645 4189
rect -31611 4155 -31572 4189
rect -31538 4155 -31499 4189
rect -31465 4155 -31426 4189
rect -31392 4155 -31353 4189
rect -31319 4155 -31280 4189
rect -31246 4155 -31207 4189
rect -31173 4155 -31134 4189
rect -31100 4155 -31061 4189
rect -31027 4155 -30988 4189
rect -30954 4155 -30915 4189
rect -30881 4155 -30842 4189
rect -30808 4155 -30768 4189
rect -30734 4155 -30694 4189
rect -30660 4155 -30620 4189
rect -30586 4155 -30546 4189
rect -30512 4155 -30472 4189
rect -30438 4155 -30398 4189
rect -30364 4155 -30324 4189
rect -30290 4155 -30250 4189
rect -30216 4155 -30176 4189
rect -30142 4155 -30102 4189
rect -30068 4155 -30028 4189
rect -29994 4155 -29954 4189
rect -29920 4155 -29880 4189
rect -29846 4155 -29806 4189
rect -29772 4155 -29732 4189
rect -29698 4155 -29658 4189
rect -29624 4155 -29584 4189
rect -29550 4155 -29510 4189
rect -29476 4155 -29436 4189
rect -29402 4155 -29362 4189
rect -29328 4155 -29288 4189
rect -29254 4155 -29214 4189
rect -29180 4187 -28830 4189
rect -29180 4155 -29134 4187
rect -31764 4153 -29134 4155
rect -29100 4153 -29046 4187
rect -29012 4153 -28958 4187
rect -28924 4153 -28870 4187
rect -28836 4153 -28830 4187
rect -31764 4152 -28830 4153
rect -32350 4117 -28830 4152
rect -32350 4113 -31718 4117
rect -32350 4079 -32344 4113
rect -32310 4079 -32266 4113
rect -32232 4079 -32188 4113
rect -32154 4079 -32110 4113
rect -32076 4079 -32032 4113
rect -31998 4079 -31954 4113
rect -31920 4079 -31876 4113
rect -31842 4079 -31798 4113
rect -31764 4083 -31718 4113
rect -31684 4083 -31645 4117
rect -31611 4083 -31572 4117
rect -31538 4083 -31499 4117
rect -31465 4083 -31426 4117
rect -31392 4083 -31353 4117
rect -31319 4083 -31280 4117
rect -31246 4083 -31207 4117
rect -31173 4083 -31134 4117
rect -31100 4083 -31061 4117
rect -31027 4083 -30988 4117
rect -30954 4083 -30915 4117
rect -30881 4083 -30842 4117
rect -30808 4083 -30768 4117
rect -30734 4083 -30694 4117
rect -30660 4083 -30620 4117
rect -30586 4083 -30546 4117
rect -30512 4083 -30472 4117
rect -30438 4083 -30398 4117
rect -30364 4083 -30324 4117
rect -30290 4083 -30250 4117
rect -30216 4083 -30176 4117
rect -30142 4083 -30102 4117
rect -30068 4083 -30028 4117
rect -29994 4083 -29954 4117
rect -29920 4083 -29880 4117
rect -29846 4083 -29806 4117
rect -29772 4083 -29732 4117
rect -29698 4083 -29658 4117
rect -29624 4083 -29584 4117
rect -29550 4083 -29510 4117
rect -29476 4083 -29436 4117
rect -29402 4083 -29362 4117
rect -29328 4083 -29288 4117
rect -29254 4083 -29214 4117
rect -29180 4114 -28830 4117
rect -29180 4083 -29134 4114
rect -31764 4080 -29134 4083
rect -29100 4080 -29046 4114
rect -29012 4080 -28958 4114
rect -28924 4080 -28870 4114
rect -28836 4080 -28830 4114
rect -31764 4079 -28830 4080
rect -32350 4045 -28830 4079
rect -32350 4040 -31718 4045
rect -32350 4006 -32344 4040
rect -32310 4006 -32266 4040
rect -32232 4006 -32188 4040
rect -32154 4006 -32110 4040
rect -32076 4006 -32032 4040
rect -31998 4006 -31954 4040
rect -31920 4006 -31876 4040
rect -31842 4006 -31798 4040
rect -31764 4011 -31718 4040
rect -31684 4011 -31645 4045
rect -31611 4011 -31572 4045
rect -31538 4011 -31499 4045
rect -31465 4011 -31426 4045
rect -31392 4011 -31353 4045
rect -31319 4011 -31280 4045
rect -31246 4011 -31207 4045
rect -31173 4011 -31134 4045
rect -31100 4011 -31061 4045
rect -31027 4011 -30988 4045
rect -30954 4011 -30915 4045
rect -30881 4011 -30842 4045
rect -30808 4011 -30768 4045
rect -30734 4011 -30694 4045
rect -30660 4011 -30620 4045
rect -30586 4011 -30546 4045
rect -30512 4011 -30472 4045
rect -30438 4011 -30398 4045
rect -30364 4011 -30324 4045
rect -30290 4011 -30250 4045
rect -30216 4011 -30176 4045
rect -30142 4011 -30102 4045
rect -30068 4011 -30028 4045
rect -29994 4011 -29954 4045
rect -29920 4011 -29880 4045
rect -29846 4011 -29806 4045
rect -29772 4011 -29732 4045
rect -29698 4011 -29658 4045
rect -29624 4011 -29584 4045
rect -29550 4011 -29510 4045
rect -29476 4011 -29436 4045
rect -29402 4011 -29362 4045
rect -29328 4011 -29288 4045
rect -29254 4011 -29214 4045
rect -29180 4041 -28830 4045
rect -29180 4011 -29134 4041
rect -31764 4007 -29134 4011
rect -29100 4007 -29046 4041
rect -29012 4007 -28958 4041
rect -28924 4007 -28870 4041
rect -28836 4007 -28830 4041
rect -31764 4006 -28830 4007
rect -32350 3973 -28830 4006
rect -32350 3967 -31718 3973
rect -32350 3933 -32344 3967
rect -32310 3933 -32266 3967
rect -32232 3933 -32188 3967
rect -32154 3933 -32110 3967
rect -32076 3933 -32032 3967
rect -31998 3933 -31954 3967
rect -31920 3933 -31876 3967
rect -31842 3933 -31798 3967
rect -31764 3939 -31718 3967
rect -31684 3939 -31645 3973
rect -31611 3939 -31572 3973
rect -31538 3939 -31499 3973
rect -31465 3939 -31426 3973
rect -31392 3939 -31353 3973
rect -31319 3939 -31280 3973
rect -31246 3939 -31207 3973
rect -31173 3939 -31134 3973
rect -31100 3939 -31061 3973
rect -31027 3939 -30988 3973
rect -30954 3939 -30915 3973
rect -30881 3939 -30842 3973
rect -30808 3939 -30768 3973
rect -30734 3939 -30694 3973
rect -30660 3939 -30620 3973
rect -30586 3939 -30546 3973
rect -30512 3939 -30472 3973
rect -30438 3939 -30398 3973
rect -30364 3939 -30324 3973
rect -30290 3939 -30250 3973
rect -30216 3939 -30176 3973
rect -30142 3939 -30102 3973
rect -30068 3939 -30028 3973
rect -29994 3939 -29954 3973
rect -29920 3939 -29880 3973
rect -29846 3939 -29806 3973
rect -29772 3939 -29732 3973
rect -29698 3939 -29658 3973
rect -29624 3939 -29584 3973
rect -29550 3939 -29510 3973
rect -29476 3939 -29436 3973
rect -29402 3939 -29362 3973
rect -29328 3939 -29288 3973
rect -29254 3939 -29214 3973
rect -29180 3968 -28830 3973
rect -29180 3939 -29134 3968
rect -31764 3934 -29134 3939
rect -29100 3934 -29046 3968
rect -29012 3934 -28958 3968
rect -28924 3934 -28870 3968
rect -28836 3934 -28830 3968
rect -31764 3933 -28830 3934
rect -32350 3901 -28830 3933
rect -32350 3894 -31718 3901
rect -32350 3860 -32344 3894
rect -32310 3860 -32266 3894
rect -32232 3860 -32188 3894
rect -32154 3860 -32110 3894
rect -32076 3860 -32032 3894
rect -31998 3860 -31954 3894
rect -31920 3860 -31876 3894
rect -31842 3860 -31798 3894
rect -31764 3867 -31718 3894
rect -31684 3867 -31645 3901
rect -31611 3867 -31572 3901
rect -31538 3867 -31499 3901
rect -31465 3867 -31426 3901
rect -31392 3867 -31353 3901
rect -31319 3867 -31280 3901
rect -31246 3867 -31207 3901
rect -31173 3867 -31134 3901
rect -31100 3867 -31061 3901
rect -31027 3867 -30988 3901
rect -30954 3867 -30915 3901
rect -30881 3867 -30842 3901
rect -30808 3867 -30768 3901
rect -30734 3867 -30694 3901
rect -30660 3867 -30620 3901
rect -30586 3867 -30546 3901
rect -30512 3867 -30472 3901
rect -30438 3867 -30398 3901
rect -30364 3867 -30324 3901
rect -30290 3867 -30250 3901
rect -30216 3867 -30176 3901
rect -30142 3867 -30102 3901
rect -30068 3867 -30028 3901
rect -29994 3867 -29954 3901
rect -29920 3867 -29880 3901
rect -29846 3867 -29806 3901
rect -29772 3867 -29732 3901
rect -29698 3867 -29658 3901
rect -29624 3867 -29584 3901
rect -29550 3867 -29510 3901
rect -29476 3867 -29436 3901
rect -29402 3867 -29362 3901
rect -29328 3867 -29288 3901
rect -29254 3867 -29214 3901
rect -29180 3895 -28830 3901
rect -29180 3867 -29134 3895
rect -31764 3861 -29134 3867
rect -29100 3861 -29046 3895
rect -29012 3861 -28958 3895
rect -28924 3861 -28870 3895
rect -28836 3861 -28830 3895
rect -31764 3860 -28830 3861
rect -32350 3829 -28830 3860
rect -32350 3821 -31718 3829
rect -32350 3787 -32344 3821
rect -32310 3787 -32266 3821
rect -32232 3787 -32188 3821
rect -32154 3787 -32110 3821
rect -32076 3787 -32032 3821
rect -31998 3787 -31954 3821
rect -31920 3787 -31876 3821
rect -31842 3787 -31798 3821
rect -31764 3795 -31718 3821
rect -31684 3795 -31645 3829
rect -31611 3795 -31572 3829
rect -31538 3795 -31499 3829
rect -31465 3795 -31426 3829
rect -31392 3795 -31353 3829
rect -31319 3795 -31280 3829
rect -31246 3795 -31207 3829
rect -31173 3795 -31134 3829
rect -31100 3795 -31061 3829
rect -31027 3795 -30988 3829
rect -30954 3795 -30915 3829
rect -30881 3795 -30842 3829
rect -30808 3795 -30768 3829
rect -30734 3795 -30694 3829
rect -30660 3795 -30620 3829
rect -30586 3795 -30546 3829
rect -30512 3795 -30472 3829
rect -30438 3795 -30398 3829
rect -30364 3795 -30324 3829
rect -30290 3795 -30250 3829
rect -30216 3795 -30176 3829
rect -30142 3795 -30102 3829
rect -30068 3795 -30028 3829
rect -29994 3795 -29954 3829
rect -29920 3795 -29880 3829
rect -29846 3795 -29806 3829
rect -29772 3795 -29732 3829
rect -29698 3795 -29658 3829
rect -29624 3795 -29584 3829
rect -29550 3795 -29510 3829
rect -29476 3795 -29436 3829
rect -29402 3795 -29362 3829
rect -29328 3795 -29288 3829
rect -29254 3795 -29214 3829
rect -29180 3822 -28830 3829
rect -29180 3795 -29134 3822
rect -31764 3788 -29134 3795
rect -29100 3788 -29046 3822
rect -29012 3788 -28958 3822
rect -28924 3788 -28870 3822
rect -28836 3788 -28830 3822
rect -31764 3787 -28830 3788
rect -32350 3757 -28830 3787
rect -32350 3748 -31718 3757
rect -32350 3714 -32344 3748
rect -32310 3714 -32266 3748
rect -32232 3714 -32188 3748
rect -32154 3714 -32110 3748
rect -32076 3714 -32032 3748
rect -31998 3714 -31954 3748
rect -31920 3714 -31876 3748
rect -31842 3714 -31798 3748
rect -31764 3723 -31718 3748
rect -31684 3723 -31645 3757
rect -31611 3723 -31572 3757
rect -31538 3723 -31499 3757
rect -31465 3723 -31426 3757
rect -31392 3723 -31353 3757
rect -31319 3723 -31280 3757
rect -31246 3723 -31207 3757
rect -31173 3723 -31134 3757
rect -31100 3723 -31061 3757
rect -31027 3723 -30988 3757
rect -30954 3723 -30915 3757
rect -30881 3723 -30842 3757
rect -30808 3723 -30768 3757
rect -30734 3723 -30694 3757
rect -30660 3723 -30620 3757
rect -30586 3723 -30546 3757
rect -30512 3723 -30472 3757
rect -30438 3723 -30398 3757
rect -30364 3723 -30324 3757
rect -30290 3723 -30250 3757
rect -30216 3723 -30176 3757
rect -30142 3723 -30102 3757
rect -30068 3723 -30028 3757
rect -29994 3723 -29954 3757
rect -29920 3723 -29880 3757
rect -29846 3723 -29806 3757
rect -29772 3723 -29732 3757
rect -29698 3723 -29658 3757
rect -29624 3723 -29584 3757
rect -29550 3723 -29510 3757
rect -29476 3723 -29436 3757
rect -29402 3723 -29362 3757
rect -29328 3723 -29288 3757
rect -29254 3723 -29214 3757
rect -29180 3749 -28830 3757
rect -29180 3723 -29134 3749
rect -31764 3715 -29134 3723
rect -29100 3715 -29046 3749
rect -29012 3715 -28958 3749
rect -28924 3715 -28870 3749
rect -28836 3715 -28830 3749
rect -31764 3714 -28830 3715
rect -32350 3685 -28830 3714
rect -32350 3675 -31718 3685
rect -32350 3641 -32344 3675
rect -32310 3641 -32266 3675
rect -32232 3641 -32188 3675
rect -32154 3641 -32110 3675
rect -32076 3641 -32032 3675
rect -31998 3641 -31954 3675
rect -31920 3641 -31876 3675
rect -31842 3641 -31798 3675
rect -31764 3651 -31718 3675
rect -31684 3651 -31645 3685
rect -31611 3651 -31572 3685
rect -31538 3651 -31499 3685
rect -31465 3651 -31426 3685
rect -31392 3651 -31353 3685
rect -31319 3651 -31280 3685
rect -31246 3651 -31207 3685
rect -31173 3651 -31134 3685
rect -31100 3651 -31061 3685
rect -31027 3651 -30988 3685
rect -30954 3651 -30915 3685
rect -30881 3651 -30842 3685
rect -30808 3651 -30768 3685
rect -30734 3651 -30694 3685
rect -30660 3651 -30620 3685
rect -30586 3651 -30546 3685
rect -30512 3651 -30472 3685
rect -30438 3651 -30398 3685
rect -30364 3651 -30324 3685
rect -30290 3651 -30250 3685
rect -30216 3651 -30176 3685
rect -30142 3651 -30102 3685
rect -30068 3651 -30028 3685
rect -29994 3651 -29954 3685
rect -29920 3651 -29880 3685
rect -29846 3651 -29806 3685
rect -29772 3651 -29732 3685
rect -29698 3651 -29658 3685
rect -29624 3651 -29584 3685
rect -29550 3651 -29510 3685
rect -29476 3651 -29436 3685
rect -29402 3651 -29362 3685
rect -29328 3651 -29288 3685
rect -29254 3651 -29214 3685
rect -29180 3676 -28830 3685
rect -29180 3651 -29134 3676
rect -31764 3642 -29134 3651
rect -29100 3642 -29046 3676
rect -29012 3642 -28958 3676
rect -28924 3642 -28870 3676
rect -28836 3642 -28830 3676
rect -31764 3641 -28830 3642
rect -32350 3613 -28830 3641
rect -32350 3602 -31718 3613
rect -32350 3568 -32344 3602
rect -32310 3568 -32266 3602
rect -32232 3568 -32188 3602
rect -32154 3568 -32110 3602
rect -32076 3568 -32032 3602
rect -31998 3568 -31954 3602
rect -31920 3568 -31876 3602
rect -31842 3568 -31798 3602
rect -31764 3579 -31718 3602
rect -31684 3579 -31645 3613
rect -31611 3579 -31572 3613
rect -31538 3579 -31499 3613
rect -31465 3579 -31426 3613
rect -31392 3579 -31353 3613
rect -31319 3579 -31280 3613
rect -31246 3579 -31207 3613
rect -31173 3579 -31134 3613
rect -31100 3579 -31061 3613
rect -31027 3579 -30988 3613
rect -30954 3579 -30915 3613
rect -30881 3579 -30842 3613
rect -30808 3579 -30768 3613
rect -30734 3579 -30694 3613
rect -30660 3579 -30620 3613
rect -30586 3579 -30546 3613
rect -30512 3579 -30472 3613
rect -30438 3579 -30398 3613
rect -30364 3579 -30324 3613
rect -30290 3579 -30250 3613
rect -30216 3579 -30176 3613
rect -30142 3579 -30102 3613
rect -30068 3579 -30028 3613
rect -29994 3579 -29954 3613
rect -29920 3579 -29880 3613
rect -29846 3579 -29806 3613
rect -29772 3579 -29732 3613
rect -29698 3579 -29658 3613
rect -29624 3579 -29584 3613
rect -29550 3579 -29510 3613
rect -29476 3579 -29436 3613
rect -29402 3579 -29362 3613
rect -29328 3579 -29288 3613
rect -29254 3579 -29214 3613
rect -29180 3603 -28830 3613
rect -29180 3579 -29134 3603
rect -31764 3569 -29134 3579
rect -29100 3569 -29046 3603
rect -29012 3569 -28958 3603
rect -28924 3569 -28870 3603
rect -28836 3569 -28830 3603
rect -31764 3568 -28830 3569
rect -32350 3541 -28830 3568
rect -32350 3529 -31718 3541
rect -32350 3495 -32344 3529
rect -32310 3495 -32266 3529
rect -32232 3495 -32188 3529
rect -32154 3495 -32110 3529
rect -32076 3495 -32032 3529
rect -31998 3495 -31954 3529
rect -31920 3495 -31876 3529
rect -31842 3495 -31798 3529
rect -31764 3507 -31718 3529
rect -31684 3507 -31645 3541
rect -31611 3507 -31572 3541
rect -31538 3507 -31499 3541
rect -31465 3507 -31426 3541
rect -31392 3507 -31353 3541
rect -31319 3507 -31280 3541
rect -31246 3507 -31207 3541
rect -31173 3507 -31134 3541
rect -31100 3507 -31061 3541
rect -31027 3507 -30988 3541
rect -30954 3507 -30915 3541
rect -30881 3507 -30842 3541
rect -30808 3507 -30768 3541
rect -30734 3507 -30694 3541
rect -30660 3507 -30620 3541
rect -30586 3507 -30546 3541
rect -30512 3507 -30472 3541
rect -30438 3507 -30398 3541
rect -30364 3507 -30324 3541
rect -30290 3507 -30250 3541
rect -30216 3507 -30176 3541
rect -30142 3507 -30102 3541
rect -30068 3507 -30028 3541
rect -29994 3507 -29954 3541
rect -29920 3507 -29880 3541
rect -29846 3507 -29806 3541
rect -29772 3507 -29732 3541
rect -29698 3507 -29658 3541
rect -29624 3507 -29584 3541
rect -29550 3507 -29510 3541
rect -29476 3507 -29436 3541
rect -29402 3507 -29362 3541
rect -29328 3507 -29288 3541
rect -29254 3507 -29214 3541
rect -29180 3530 -28830 3541
rect -29180 3507 -29134 3530
rect -31764 3496 -29134 3507
rect -29100 3496 -29046 3530
rect -29012 3496 -28958 3530
rect -28924 3496 -28870 3530
rect -28836 3496 -28830 3530
rect -31764 3495 -28830 3496
rect -32350 3469 -28830 3495
rect -32350 3456 -31718 3469
rect -32350 3422 -32344 3456
rect -32310 3422 -32266 3456
rect -32232 3422 -32188 3456
rect -32154 3422 -32110 3456
rect -32076 3422 -32032 3456
rect -31998 3422 -31954 3456
rect -31920 3422 -31876 3456
rect -31842 3422 -31798 3456
rect -31764 3435 -31718 3456
rect -31684 3435 -31645 3469
rect -31611 3435 -31572 3469
rect -31538 3435 -31499 3469
rect -31465 3435 -31426 3469
rect -31392 3435 -31353 3469
rect -31319 3435 -31280 3469
rect -31246 3435 -31207 3469
rect -31173 3435 -31134 3469
rect -31100 3435 -31061 3469
rect -31027 3435 -30988 3469
rect -30954 3435 -30915 3469
rect -30881 3435 -30842 3469
rect -30808 3435 -30768 3469
rect -30734 3435 -30694 3469
rect -30660 3435 -30620 3469
rect -30586 3435 -30546 3469
rect -30512 3435 -30472 3469
rect -30438 3435 -30398 3469
rect -30364 3435 -30324 3469
rect -30290 3435 -30250 3469
rect -30216 3435 -30176 3469
rect -30142 3435 -30102 3469
rect -30068 3435 -30028 3469
rect -29994 3435 -29954 3469
rect -29920 3435 -29880 3469
rect -29846 3435 -29806 3469
rect -29772 3435 -29732 3469
rect -29698 3435 -29658 3469
rect -29624 3435 -29584 3469
rect -29550 3435 -29510 3469
rect -29476 3435 -29436 3469
rect -29402 3435 -29362 3469
rect -29328 3435 -29288 3469
rect -29254 3435 -29214 3469
rect -29180 3457 -28830 3469
rect -29180 3435 -29134 3457
rect -31764 3423 -29134 3435
rect -29100 3423 -29046 3457
rect -29012 3423 -28958 3457
rect -28924 3423 -28870 3457
rect -28836 3423 -28830 3457
rect -31764 3422 -28830 3423
rect -32350 3397 -28830 3422
rect -32350 3383 -31718 3397
rect -32350 3349 -32344 3383
rect -32310 3349 -32266 3383
rect -32232 3349 -32188 3383
rect -32154 3349 -32110 3383
rect -32076 3349 -32032 3383
rect -31998 3349 -31954 3383
rect -31920 3349 -31876 3383
rect -31842 3349 -31798 3383
rect -31764 3363 -31718 3383
rect -31684 3363 -31645 3397
rect -31611 3363 -31572 3397
rect -31538 3363 -31499 3397
rect -31465 3363 -31426 3397
rect -31392 3363 -31353 3397
rect -31319 3363 -31280 3397
rect -31246 3363 -31207 3397
rect -31173 3363 -31134 3397
rect -31100 3363 -31061 3397
rect -31027 3363 -30988 3397
rect -30954 3363 -30915 3397
rect -30881 3363 -30842 3397
rect -30808 3363 -30768 3397
rect -30734 3363 -30694 3397
rect -30660 3363 -30620 3397
rect -30586 3363 -30546 3397
rect -30512 3363 -30472 3397
rect -30438 3363 -30398 3397
rect -30364 3363 -30324 3397
rect -30290 3363 -30250 3397
rect -30216 3363 -30176 3397
rect -30142 3363 -30102 3397
rect -30068 3363 -30028 3397
rect -29994 3363 -29954 3397
rect -29920 3363 -29880 3397
rect -29846 3363 -29806 3397
rect -29772 3363 -29732 3397
rect -29698 3363 -29658 3397
rect -29624 3363 -29584 3397
rect -29550 3363 -29510 3397
rect -29476 3363 -29436 3397
rect -29402 3363 -29362 3397
rect -29328 3363 -29288 3397
rect -29254 3363 -29214 3397
rect -29180 3384 -28830 3397
rect -29180 3363 -29134 3384
rect -31764 3352 -29134 3363
rect -31764 3350 -31544 3352
tri -31544 3350 -31542 3352 nw
tri -29656 3350 -29654 3352 ne
rect -29654 3350 -29134 3352
rect -29100 3350 -29046 3384
rect -29012 3350 -28958 3384
rect -28924 3350 -28870 3384
rect -28836 3350 -28830 3384
rect -31764 3349 -31565 3350
rect -32350 3329 -31565 3349
tri -31565 3329 -31544 3350 nw
tri -29654 3329 -29633 3350 ne
rect -29633 3329 -28830 3350
rect -32350 3311 -31583 3329
tri -31583 3311 -31565 3329 nw
tri -29633 3311 -29615 3329 ne
rect -29615 3311 -28830 3329
rect -32350 3310 -31617 3311
rect -32350 3276 -32344 3310
rect -32310 3276 -32266 3310
rect -32232 3276 -32188 3310
rect -32154 3276 -32110 3310
rect -32076 3276 -32032 3310
rect -31998 3276 -31954 3310
rect -31920 3276 -31876 3310
rect -31842 3276 -31798 3310
rect -31764 3277 -31617 3310
tri -31617 3277 -31583 3311 nw
tri -29615 3277 -29581 3311 ne
rect -29581 3277 -29134 3311
rect -29100 3277 -29046 3311
rect -29012 3277 -28958 3311
rect -28924 3277 -28870 3311
rect -28836 3277 -28830 3311
rect -31764 3276 -31638 3277
rect -32350 3256 -31638 3276
tri -31638 3256 -31617 3277 nw
tri -29581 3256 -29560 3277 ne
rect -29560 3256 -28830 3277
rect -32350 3238 -31656 3256
tri -31656 3238 -31638 3256 nw
tri -29560 3238 -29542 3256 ne
rect -29542 3238 -28830 3256
rect -32350 3237 -31690 3238
rect -32350 3203 -32344 3237
rect -32310 3203 -32266 3237
rect -32232 3203 -32188 3237
rect -32154 3203 -32110 3237
rect -32076 3203 -32032 3237
rect -31998 3203 -31954 3237
rect -31920 3203 -31876 3237
rect -31842 3203 -31798 3237
rect -31764 3204 -31690 3237
tri -31690 3204 -31656 3238 nw
tri -29542 3204 -29508 3238 ne
rect -29508 3204 -29134 3238
rect -29100 3204 -29046 3238
rect -29012 3204 -28958 3238
rect -28924 3204 -28870 3238
rect -28836 3204 -28830 3238
rect -31764 3203 -31711 3204
rect -32350 3183 -31711 3203
tri -31711 3183 -31690 3204 nw
tri -29508 3183 -29487 3204 ne
rect -29487 3183 -28830 3204
rect -32350 3165 -31729 3183
tri -31729 3165 -31711 3183 nw
tri -29487 3165 -29469 3183 ne
rect -29469 3165 -28830 3183
rect -32350 3164 -31758 3165
rect -32350 3130 -32344 3164
rect -32310 3130 -32266 3164
rect -32232 3130 -32188 3164
rect -32154 3130 -32110 3164
rect -32076 3130 -32032 3164
rect -31998 3130 -31954 3164
rect -31920 3130 -31876 3164
rect -31842 3130 -31798 3164
rect -31764 3130 -31758 3164
tri -31758 3136 -31729 3165 nw
tri -29469 3136 -29440 3165 ne
rect -29440 3136 -29134 3165
tri -29440 3131 -29435 3136 ne
rect -29435 3131 -29134 3136
rect -29100 3131 -29046 3165
rect -29012 3131 -28958 3165
rect -28924 3131 -28870 3165
rect -28836 3131 -28830 3165
rect -32350 3091 -31758 3130
tri -29435 3110 -29414 3131 ne
rect -29414 3110 -28830 3131
tri -29414 3092 -29396 3110 ne
rect -29396 3092 -28830 3110
rect -32350 3057 -32344 3091
rect -32310 3057 -32266 3091
rect -32232 3057 -32188 3091
rect -32154 3057 -32110 3091
rect -32076 3057 -32032 3091
rect -31998 3057 -31954 3091
rect -31920 3057 -31876 3091
rect -31842 3057 -31798 3091
rect -31764 3057 -31758 3091
tri -29396 3058 -29362 3092 ne
rect -29362 3058 -29134 3092
rect -29100 3058 -29046 3092
rect -29012 3058 -28958 3092
rect -28924 3058 -28870 3092
rect -28836 3058 -28830 3092
rect -32350 3018 -31758 3057
tri -29362 3037 -29341 3058 ne
rect -29341 3037 -28830 3058
tri -29341 3019 -29323 3037 ne
rect -29323 3019 -28830 3037
rect -32350 2984 -32344 3018
rect -32310 2984 -32266 3018
rect -32232 2984 -32188 3018
rect -32154 2984 -32110 3018
rect -32076 2984 -32032 3018
rect -31998 2984 -31954 3018
rect -31920 2984 -31876 3018
rect -31842 2984 -31798 3018
rect -31764 2984 -31758 3018
tri -29323 2985 -29289 3019 ne
rect -29289 2985 -29134 3019
rect -29100 2985 -29046 3019
rect -29012 2985 -28958 3019
rect -28924 2985 -28870 3019
rect -28836 2985 -28830 3019
rect -32350 2945 -31758 2984
tri -29289 2964 -29268 2985 ne
rect -29268 2964 -28830 2985
tri -29268 2946 -29250 2964 ne
rect -29250 2946 -28830 2964
rect -32350 2911 -32344 2945
rect -32310 2911 -32266 2945
rect -32232 2911 -32188 2945
rect -32154 2911 -32110 2945
rect -32076 2911 -32032 2945
rect -31998 2911 -31954 2945
rect -31920 2911 -31876 2945
rect -31842 2911 -31798 2945
rect -31764 2911 -31758 2945
tri -29250 2912 -29216 2946 ne
rect -29216 2912 -29134 2946
rect -29100 2912 -29046 2946
rect -29012 2912 -28958 2946
rect -28924 2912 -28870 2946
rect -28836 2912 -28830 2946
rect -32350 2872 -31758 2911
tri -29216 2891 -29195 2912 ne
rect -29195 2891 -28830 2912
tri -29195 2873 -29177 2891 ne
rect -29177 2873 -28830 2891
rect -32350 2838 -32344 2872
rect -32310 2838 -32266 2872
rect -32232 2838 -32188 2872
rect -32154 2838 -32110 2872
rect -32076 2838 -32032 2872
rect -31998 2838 -31954 2872
rect -31920 2838 -31876 2872
rect -31842 2838 -31798 2872
rect -31764 2838 -31758 2872
tri -29177 2839 -29143 2873 ne
rect -29143 2839 -29134 2873
rect -29100 2839 -29046 2873
rect -29012 2839 -28958 2873
rect -28924 2839 -28870 2873
rect -28836 2839 -28830 2873
rect -32350 2799 -31758 2838
tri -29143 2836 -29140 2839 ne
rect -32350 2765 -32344 2799
rect -32310 2765 -32266 2799
rect -32232 2765 -32188 2799
rect -32154 2765 -32110 2799
rect -32076 2765 -32032 2799
rect -31998 2765 -31954 2799
rect -31920 2765 -31876 2799
rect -31842 2765 -31798 2799
rect -31764 2765 -31758 2799
rect -32350 2726 -31758 2765
rect -32350 2692 -32344 2726
rect -32310 2692 -32266 2726
rect -32232 2692 -32188 2726
rect -32154 2692 -32110 2726
rect -32076 2692 -32032 2726
rect -31998 2692 -31954 2726
rect -31920 2692 -31876 2726
rect -31842 2692 -31798 2726
rect -31764 2692 -31758 2726
rect -32350 2653 -31758 2692
rect -32350 2619 -32344 2653
rect -32310 2619 -32266 2653
rect -32232 2619 -32188 2653
rect -32154 2619 -32110 2653
rect -32076 2619 -32032 2653
rect -31998 2619 -31954 2653
rect -31920 2619 -31876 2653
rect -31842 2619 -31798 2653
rect -31764 2619 -31758 2653
rect -32350 2580 -31758 2619
rect -32350 2546 -32344 2580
rect -32310 2546 -32266 2580
rect -32232 2546 -32188 2580
rect -32154 2546 -32110 2580
rect -32076 2546 -32032 2580
rect -31998 2546 -31954 2580
rect -31920 2546 -31876 2580
rect -31842 2546 -31798 2580
rect -31764 2546 -31758 2580
rect -32350 2507 -31758 2546
rect -32350 2473 -32344 2507
rect -32310 2473 -32266 2507
rect -32232 2473 -32188 2507
rect -32154 2473 -32110 2507
rect -32076 2473 -32032 2507
rect -31998 2473 -31954 2507
rect -31920 2473 -31876 2507
rect -31842 2473 -31798 2507
rect -31764 2473 -31758 2507
rect -32350 2434 -31758 2473
rect -32350 2400 -32344 2434
rect -32310 2400 -32266 2434
rect -32232 2400 -32188 2434
rect -32154 2400 -32110 2434
rect -32076 2400 -32032 2434
rect -31998 2400 -31954 2434
rect -31920 2400 -31876 2434
rect -31842 2400 -31798 2434
rect -31764 2400 -31758 2434
rect -32350 2361 -31758 2400
rect -32350 2327 -32344 2361
rect -32310 2327 -32266 2361
rect -32232 2327 -32188 2361
rect -32154 2327 -32110 2361
rect -32076 2327 -32032 2361
rect -31998 2327 -31954 2361
rect -31920 2327 -31876 2361
rect -31842 2327 -31798 2361
rect -31764 2327 -31758 2361
rect -32350 2288 -31758 2327
rect -32350 2254 -32344 2288
rect -32310 2254 -32266 2288
rect -32232 2254 -32188 2288
rect -32154 2254 -32110 2288
rect -32076 2254 -32032 2288
rect -31998 2254 -31954 2288
rect -31920 2254 -31876 2288
rect -31842 2254 -31798 2288
rect -31764 2254 -31758 2288
rect -32350 2215 -31758 2254
rect -32350 2181 -32344 2215
rect -32310 2181 -32266 2215
rect -32232 2181 -32188 2215
rect -32154 2181 -32110 2215
rect -32076 2181 -32032 2215
rect -31998 2181 -31954 2215
rect -31920 2181 -31876 2215
rect -31842 2181 -31798 2215
rect -31764 2181 -31758 2215
rect -32350 2142 -31758 2181
rect -32350 2108 -32344 2142
rect -32310 2108 -32266 2142
rect -32232 2108 -32188 2142
rect -32154 2108 -32110 2142
rect -32076 2108 -32032 2142
rect -31998 2108 -31954 2142
rect -31920 2108 -31876 2142
rect -31842 2108 -31798 2142
rect -31764 2108 -31758 2142
rect -32350 2069 -31758 2108
rect -32350 2035 -32344 2069
rect -32310 2035 -32266 2069
rect -32232 2035 -32188 2069
rect -32154 2035 -32110 2069
rect -32076 2035 -32032 2069
rect -31998 2035 -31954 2069
rect -31920 2035 -31876 2069
rect -31842 2035 -31798 2069
rect -31764 2035 -31758 2069
rect -32350 1996 -31758 2035
rect -32350 1962 -32344 1996
rect -32310 1962 -32266 1996
rect -32232 1962 -32188 1996
rect -32154 1962 -32110 1996
rect -32076 1962 -32032 1996
rect -31998 1962 -31954 1996
rect -31920 1962 -31876 1996
rect -31842 1962 -31798 1996
rect -31764 1962 -31758 1996
rect -32350 1923 -31758 1962
rect -32350 1889 -32344 1923
rect -32310 1889 -32266 1923
rect -32232 1889 -32188 1923
rect -32154 1889 -32110 1923
rect -32076 1889 -32032 1923
rect -31998 1889 -31954 1923
rect -31920 1889 -31876 1923
rect -31842 1889 -31798 1923
rect -31764 1889 -31758 1923
rect -32350 1850 -31758 1889
rect -32350 1816 -32344 1850
rect -32310 1816 -32266 1850
rect -32232 1816 -32188 1850
rect -32154 1816 -32110 1850
rect -32076 1816 -32032 1850
rect -31998 1816 -31954 1850
rect -31920 1816 -31876 1850
rect -31842 1816 -31798 1850
rect -31764 1816 -31758 1850
rect -32350 1777 -31758 1816
rect -32350 1743 -32344 1777
rect -32310 1743 -32266 1777
rect -32232 1743 -32188 1777
rect -32154 1743 -32110 1777
rect -32076 1743 -32032 1777
rect -31998 1743 -31954 1777
rect -31920 1743 -31876 1777
rect -31842 1743 -31798 1777
rect -31764 1743 -31758 1777
rect -32350 1704 -31758 1743
rect -32350 1670 -32344 1704
rect -32310 1670 -32266 1704
rect -32232 1670 -32188 1704
rect -32154 1670 -32110 1704
rect -32076 1670 -32032 1704
rect -31998 1670 -31954 1704
rect -31920 1670 -31876 1704
rect -31842 1670 -31798 1704
rect -31764 1670 -31758 1704
rect -32350 1631 -31758 1670
rect -32350 1597 -32344 1631
rect -32310 1597 -32266 1631
rect -32232 1597 -32188 1631
rect -32154 1597 -32110 1631
rect -32076 1597 -32032 1631
rect -31998 1597 -31954 1631
rect -31920 1597 -31876 1631
rect -31842 1597 -31798 1631
rect -31764 1597 -31758 1631
rect -32350 1558 -31758 1597
rect -32350 1524 -32344 1558
rect -32310 1524 -32266 1558
rect -32232 1524 -32188 1558
rect -32154 1524 -32110 1558
rect -32076 1524 -32032 1558
rect -31998 1524 -31954 1558
rect -31920 1524 -31876 1558
rect -31842 1524 -31798 1558
rect -31764 1524 -31758 1558
rect -32350 1485 -31758 1524
rect -32350 1451 -32344 1485
rect -32310 1451 -32266 1485
rect -32232 1451 -32188 1485
rect -32154 1451 -32110 1485
rect -32076 1451 -32032 1485
rect -31998 1451 -31954 1485
rect -31920 1451 -31876 1485
rect -31842 1451 -31798 1485
rect -31764 1451 -31758 1485
rect -32350 1412 -31758 1451
rect -32350 1378 -32344 1412
rect -32310 1378 -32266 1412
rect -32232 1378 -32188 1412
rect -32154 1378 -32110 1412
rect -32076 1378 -32032 1412
rect -31998 1378 -31954 1412
rect -31920 1378 -31876 1412
rect -31842 1378 -31798 1412
rect -31764 1378 -31758 1412
rect -32350 1339 -31758 1378
rect -32350 1305 -32344 1339
rect -32310 1305 -32266 1339
rect -32232 1305 -32188 1339
rect -32154 1305 -32110 1339
rect -32076 1305 -32032 1339
rect -31998 1305 -31954 1339
rect -31920 1305 -31876 1339
rect -31842 1305 -31798 1339
rect -31764 1305 -31758 1339
rect -32350 1266 -31758 1305
rect -32350 1232 -32344 1266
rect -32310 1232 -32266 1266
rect -32232 1232 -32188 1266
rect -32154 1232 -32110 1266
rect -32076 1232 -32032 1266
rect -31998 1232 -31954 1266
rect -31920 1232 -31876 1266
rect -31842 1232 -31798 1266
rect -31764 1232 -31758 1266
rect -32350 1193 -31758 1232
rect -32350 1159 -32344 1193
rect -32310 1159 -32266 1193
rect -32232 1159 -32188 1193
rect -32154 1159 -32110 1193
rect -32076 1159 -32032 1193
rect -31998 1159 -31954 1193
rect -31920 1159 -31876 1193
rect -31842 1159 -31798 1193
rect -31764 1159 -31758 1193
rect -32350 1120 -31758 1159
rect -32350 1086 -32344 1120
rect -32310 1086 -32266 1120
rect -32232 1086 -32188 1120
rect -32154 1086 -32110 1120
rect -32076 1086 -32032 1120
rect -31998 1086 -31954 1120
rect -31920 1086 -31876 1120
rect -31842 1086 -31798 1120
rect -31764 1086 -31758 1120
rect -32350 1047 -31758 1086
rect -32350 1013 -32344 1047
rect -32310 1013 -32266 1047
rect -32232 1013 -32188 1047
rect -32154 1013 -32110 1047
rect -32076 1013 -32032 1047
rect -31998 1013 -31954 1047
rect -31920 1013 -31876 1047
rect -31842 1013 -31798 1047
rect -31764 1013 -31758 1047
rect -32350 974 -31758 1013
rect -32350 940 -32344 974
rect -32310 940 -32266 974
rect -32232 940 -32188 974
rect -32154 940 -32110 974
rect -32076 940 -32032 974
rect -31998 940 -31954 974
rect -31920 940 -31876 974
rect -31842 940 -31798 974
rect -31764 940 -31758 974
rect -32350 901 -31758 940
rect -32350 867 -32344 901
rect -32310 867 -32266 901
rect -32232 867 -32188 901
rect -32154 867 -32110 901
rect -32076 867 -32032 901
rect -31998 867 -31954 901
rect -31920 867 -31876 901
rect -31842 867 -31798 901
rect -31764 867 -31758 901
rect -32350 828 -31758 867
rect -32350 794 -32344 828
rect -32310 794 -32266 828
rect -32232 794 -32188 828
rect -32154 794 -32110 828
rect -32076 794 -32032 828
rect -31998 794 -31954 828
rect -31920 794 -31876 828
rect -31842 794 -31798 828
rect -31764 794 -31758 828
rect -32350 755 -31758 794
rect -32350 721 -32344 755
rect -32310 721 -32266 755
rect -32232 721 -32188 755
rect -32154 721 -32110 755
rect -32076 721 -32032 755
rect -31998 721 -31954 755
rect -31920 721 -31876 755
rect -31842 721 -31798 755
rect -31764 721 -31758 755
rect -32350 682 -31758 721
rect -32350 648 -32344 682
rect -32310 648 -32266 682
rect -32232 648 -32188 682
rect -32154 648 -32110 682
rect -32076 648 -32032 682
rect -31998 648 -31954 682
rect -31920 648 -31876 682
rect -31842 648 -31798 682
rect -31764 648 -31758 682
rect -32350 610 -31758 648
rect -32350 576 -32344 610
rect -32310 576 -32266 610
rect -32232 576 -32188 610
rect -32154 576 -32110 610
rect -32076 576 -32032 610
rect -31998 576 -31954 610
rect -31920 576 -31876 610
rect -31842 576 -31798 610
rect -31764 576 -31758 610
rect -32350 538 -31758 576
rect -32350 504 -32344 538
rect -32310 504 -32266 538
rect -32232 504 -32188 538
rect -32154 504 -32110 538
rect -32076 504 -32032 538
rect -31998 504 -31954 538
rect -31920 504 -31876 538
rect -31842 504 -31798 538
rect -31764 504 -31758 538
rect -32350 501 -31758 504
rect -32350 466 -32338 501
rect -32350 432 -32344 466
rect -32286 449 -32273 501
rect -32221 449 -32208 501
rect -32156 466 -32143 501
rect -32091 466 -32078 501
rect -32026 466 -32013 501
rect -31961 466 -31948 501
rect -32154 449 -32143 466
rect -31961 449 -31954 466
rect -31896 449 -31882 501
rect -31830 449 -31816 501
rect -32310 437 -32266 449
rect -32232 437 -32188 449
rect -32154 437 -32110 449
rect -32076 437 -32032 449
rect -31998 437 -31954 449
rect -31920 437 -31876 449
rect -31842 437 -31798 449
rect -32350 394 -32338 432
rect -32350 360 -32344 394
rect -32286 385 -32273 437
rect -32221 385 -32208 437
rect -32154 432 -32143 437
rect -31961 432 -31954 437
rect -32156 394 -32143 432
rect -32091 394 -32078 432
rect -32026 394 -32013 432
rect -31961 394 -31948 432
rect -32154 385 -32143 394
rect -31961 385 -31954 394
rect -31896 385 -31882 437
rect -31830 385 -31816 437
rect -32310 373 -32266 385
rect -32232 373 -32188 385
rect -32154 373 -32110 385
rect -32076 373 -32032 385
rect -31998 373 -31954 385
rect -31920 373 -31876 385
rect -31842 373 -31798 385
rect -32350 322 -32338 360
rect -32350 288 -32344 322
rect -32286 321 -32273 373
rect -32221 321 -32208 373
rect -32154 360 -32143 373
rect -31961 360 -31954 373
rect -32156 322 -32143 360
rect -32091 322 -32078 360
rect -32026 322 -32013 360
rect -31961 322 -31948 360
rect -32154 321 -32143 322
rect -31961 321 -31954 322
rect -31896 321 -31882 373
rect -31830 321 -31816 373
rect -32310 309 -32266 321
rect -32232 309 -32188 321
rect -32154 309 -32110 321
rect -32076 309 -32032 321
rect -31998 309 -31954 321
rect -31920 309 -31876 321
rect -31842 309 -31798 321
rect -32350 257 -32338 288
rect -32286 257 -32273 309
rect -32221 257 -32208 309
rect -32154 288 -32143 309
rect -31961 288 -31954 309
rect -32156 257 -32143 288
rect -32091 257 -32078 288
rect -32026 257 -32013 288
rect -31961 257 -31948 288
rect -31896 257 -31882 309
rect -31830 257 -31816 309
rect -31764 257 -31758 501
rect -32350 250 -31758 257
rect -32350 216 -32344 250
rect -32310 245 -32266 250
rect -32232 245 -32188 250
rect -32154 245 -32110 250
rect -32076 245 -32032 250
rect -31998 245 -31954 250
rect -31920 245 -31876 250
rect -31842 245 -31798 250
rect -32350 193 -32338 216
rect -32286 193 -32273 245
rect -32221 193 -32208 245
rect -32154 216 -32143 245
rect -31961 216 -31954 245
rect -32156 193 -32143 216
rect -32091 193 -32078 216
rect -32026 193 -32013 216
rect -31961 193 -31948 216
rect -31896 193 -31882 245
rect -31830 193 -31816 245
rect -31764 193 -31758 250
rect -32350 181 -31758 193
rect -32350 178 -32338 181
rect -32350 144 -32344 178
rect -32350 129 -32338 144
rect -32286 129 -32273 181
rect -32221 129 -32208 181
rect -32156 178 -32143 181
rect -32091 178 -32078 181
rect -32026 178 -32013 181
rect -31961 178 -31948 181
rect -32154 144 -32143 178
rect -31961 144 -31954 178
rect -32156 129 -32143 144
rect -32091 129 -32078 144
rect -32026 129 -32013 144
rect -31961 129 -31948 144
rect -31896 129 -31882 181
rect -31830 129 -31816 181
rect -31764 129 -31758 181
rect -32350 117 -31758 129
rect -32350 106 -32338 117
rect -32350 72 -32344 106
rect -32350 65 -32338 72
rect -32286 65 -32273 117
rect -32221 65 -32208 117
rect -32156 106 -32143 117
rect -32091 106 -32078 117
rect -32026 106 -32013 117
rect -31961 106 -31948 117
rect -32154 72 -32143 106
rect -31961 72 -31954 106
rect -32156 65 -32143 72
rect -32091 65 -32078 72
rect -32026 65 -32013 72
rect -31961 65 -31948 72
rect -31896 65 -31882 117
rect -31830 65 -31816 117
rect -31764 65 -31758 117
rect -32350 53 -31758 65
rect -32350 34 -32338 53
rect -32350 0 -32344 34
rect -32286 1 -32273 53
rect -32221 1 -32208 53
rect -32156 34 -32143 53
rect -32091 34 -32078 53
rect -32026 34 -32013 53
rect -31961 34 -31948 53
rect -32154 1 -32143 34
rect -31961 1 -31954 34
rect -31896 1 -31882 53
rect -31830 1 -31816 53
rect -32310 0 -32266 1
rect -32232 0 -32188 1
rect -32154 0 -32110 1
rect -32076 0 -32032 1
rect -31998 0 -31954 1
rect -31920 0 -31876 1
rect -31842 0 -31798 1
rect -31764 0 -31758 53
rect -32350 -11 -31758 0
rect -32350 -38 -32338 -11
rect -32350 -72 -32344 -38
rect -32286 -63 -32273 -11
rect -32221 -63 -32208 -11
rect -32156 -38 -32143 -11
rect -32091 -38 -32078 -11
rect -32026 -38 -32013 -11
rect -31961 -38 -31948 -11
rect -32154 -63 -32143 -38
rect -31961 -63 -31954 -38
rect -31896 -63 -31882 -11
rect -31830 -63 -31816 -11
rect -32310 -72 -32266 -63
rect -32232 -72 -32188 -63
rect -32154 -72 -32110 -63
rect -32076 -72 -32032 -63
rect -31998 -72 -31954 -63
rect -31920 -72 -31876 -63
rect -31842 -72 -31798 -63
rect -31764 -72 -31758 -11
rect -32350 -75 -31758 -72
rect -32350 -110 -32338 -75
rect -32350 -144 -32344 -110
rect -32286 -127 -32273 -75
rect -32221 -127 -32208 -75
rect -32156 -110 -32143 -75
rect -32091 -110 -32078 -75
rect -32026 -110 -32013 -75
rect -31961 -110 -31948 -75
rect -32154 -127 -32143 -110
rect -31961 -127 -31954 -110
rect -31896 -127 -31882 -75
rect -31830 -127 -31816 -75
rect -32310 -139 -32266 -127
rect -32232 -139 -32188 -127
rect -32154 -139 -32110 -127
rect -32076 -139 -32032 -127
rect -31998 -139 -31954 -127
rect -31920 -139 -31876 -127
rect -31842 -139 -31798 -127
rect -32350 -182 -32338 -144
rect -32350 -216 -32344 -182
rect -32286 -191 -32273 -139
rect -32221 -191 -32208 -139
rect -32154 -144 -32143 -139
rect -31961 -144 -31954 -139
rect -32156 -182 -32143 -144
rect -32091 -182 -32078 -144
rect -32026 -182 -32013 -144
rect -31961 -182 -31948 -144
rect -32154 -191 -32143 -182
rect -31961 -191 -31954 -182
rect -31896 -191 -31882 -139
rect -31830 -191 -31816 -139
rect -32310 -203 -32266 -191
rect -32232 -203 -32188 -191
rect -32154 -203 -32110 -191
rect -32076 -203 -32032 -191
rect -31998 -203 -31954 -191
rect -31920 -203 -31876 -191
rect -31842 -203 -31798 -191
rect -32350 -254 -32338 -216
rect -32350 -288 -32344 -254
rect -32286 -255 -32273 -203
rect -32221 -255 -32208 -203
rect -32154 -216 -32143 -203
rect -31961 -216 -31954 -203
rect -32156 -254 -32143 -216
rect -32091 -254 -32078 -216
rect -32026 -254 -32013 -216
rect -31961 -254 -31948 -216
rect -32154 -255 -32143 -254
rect -31961 -255 -31954 -254
rect -31896 -255 -31882 -203
rect -31830 -255 -31816 -203
rect -32310 -267 -32266 -255
rect -32232 -267 -32188 -255
rect -32154 -267 -32110 -255
rect -32076 -267 -32032 -255
rect -31998 -267 -31954 -255
rect -31920 -267 -31876 -255
rect -31842 -267 -31798 -255
rect -32350 -319 -32338 -288
rect -32286 -319 -32273 -267
rect -32221 -319 -32208 -267
rect -32154 -288 -32143 -267
rect -31961 -288 -31954 -267
rect -32156 -319 -32143 -288
rect -32091 -319 -32078 -288
rect -32026 -319 -32013 -288
rect -31961 -319 -31948 -288
rect -31896 -319 -31882 -267
rect -31830 -319 -31816 -267
rect -31764 -319 -31758 -75
rect -32350 -326 -31758 -319
rect -32350 -360 -32344 -326
rect -32310 -331 -32266 -326
rect -32232 -331 -32188 -326
rect -32154 -331 -32110 -326
rect -32076 -331 -32032 -326
rect -31998 -331 -31954 -326
rect -31920 -331 -31876 -326
rect -31842 -331 -31798 -326
rect -32350 -383 -32338 -360
rect -32286 -383 -32273 -331
rect -32221 -383 -32208 -331
rect -32154 -360 -32143 -331
rect -31961 -360 -31954 -331
rect -32156 -383 -32143 -360
rect -32091 -383 -32078 -360
rect -32026 -383 -32013 -360
rect -31961 -383 -31948 -360
rect -31896 -383 -31882 -331
rect -31830 -383 -31816 -331
rect -31764 -383 -31758 -326
rect -32350 -398 -31758 -383
rect -32350 -432 -32344 -398
rect -32310 -432 -32266 -398
rect -32232 -432 -32188 -398
rect -32154 -432 -32110 -398
rect -32076 -432 -32032 -398
rect -31998 -432 -31954 -398
rect -31920 -432 -31876 -398
rect -31842 -432 -31798 -398
rect -31764 -432 -31758 -398
rect -32350 -470 -31758 -432
rect -32350 -504 -32344 -470
rect -32310 -504 -32266 -470
rect -32232 -504 -32188 -470
rect -32154 -504 -32110 -470
rect -32076 -504 -32032 -470
rect -31998 -504 -31954 -470
rect -31920 -504 -31876 -470
rect -31842 -504 -31798 -470
rect -31764 -504 -31758 -470
rect -32350 -542 -31758 -504
rect -32350 -576 -32344 -542
rect -32310 -576 -32266 -542
rect -32232 -576 -32188 -542
rect -32154 -576 -32110 -542
rect -32076 -576 -32032 -542
rect -31998 -576 -31954 -542
rect -31920 -576 -31876 -542
rect -31842 -576 -31798 -542
rect -31764 -576 -31758 -542
rect -32350 -614 -31758 -576
rect -32350 -648 -32344 -614
rect -32310 -648 -32266 -614
rect -32232 -648 -32188 -614
rect -32154 -648 -32110 -614
rect -32076 -648 -32032 -614
rect -31998 -648 -31954 -614
rect -31920 -648 -31876 -614
rect -31842 -648 -31798 -614
rect -31764 -648 -31758 -614
rect -32350 -686 -31758 -648
rect -32350 -720 -32344 -686
rect -32310 -720 -32266 -686
rect -32232 -720 -32188 -686
rect -32154 -720 -32110 -686
rect -32076 -720 -32032 -686
rect -31998 -720 -31954 -686
rect -31920 -720 -31876 -686
rect -31842 -720 -31798 -686
rect -31764 -720 -31758 -686
rect -32350 -758 -31758 -720
rect -32350 -792 -32344 -758
rect -32310 -792 -32266 -758
rect -32232 -792 -32188 -758
rect -32154 -792 -32110 -758
rect -32076 -792 -32032 -758
rect -31998 -792 -31954 -758
rect -31920 -792 -31876 -758
rect -31842 -792 -31798 -758
rect -31764 -792 -31758 -758
rect -32350 -830 -31758 -792
rect -32350 -864 -32344 -830
rect -32310 -864 -32266 -830
rect -32232 -864 -32188 -830
rect -32154 -864 -32110 -830
rect -32076 -864 -32032 -830
rect -31998 -864 -31954 -830
rect -31920 -864 -31876 -830
rect -31842 -864 -31798 -830
rect -31764 -864 -31758 -830
rect -32350 -902 -31758 -864
rect -32350 -936 -32344 -902
rect -32310 -936 -32266 -902
rect -32232 -936 -32188 -902
rect -32154 -936 -32110 -902
rect -32076 -936 -32032 -902
rect -31998 -936 -31954 -902
rect -31920 -936 -31876 -902
rect -31842 -936 -31798 -902
rect -31764 -936 -31758 -902
rect -32350 -974 -31758 -936
rect -32350 -1008 -32344 -974
rect -32310 -1008 -32266 -974
rect -32232 -1008 -32188 -974
rect -32154 -1008 -32110 -974
rect -32076 -1008 -32032 -974
rect -31998 -1008 -31954 -974
rect -31920 -1008 -31876 -974
rect -31842 -1008 -31798 -974
rect -31764 -1008 -31758 -974
rect -32350 -1046 -31758 -1008
rect -32350 -1080 -32344 -1046
rect -32310 -1080 -32266 -1046
rect -32232 -1080 -32188 -1046
rect -32154 -1080 -32110 -1046
rect -32076 -1080 -32032 -1046
rect -31998 -1080 -31954 -1046
rect -31920 -1080 -31876 -1046
rect -31842 -1080 -31798 -1046
rect -31764 -1080 -31758 -1046
rect -32350 -1118 -31758 -1080
rect -32350 -1152 -32344 -1118
rect -32310 -1152 -32266 -1118
rect -32232 -1152 -32188 -1118
rect -32154 -1152 -32110 -1118
rect -32076 -1152 -32032 -1118
rect -31998 -1152 -31954 -1118
rect -31920 -1152 -31876 -1118
rect -31842 -1152 -31798 -1118
rect -31764 -1152 -31758 -1118
rect -32350 -1190 -31758 -1152
rect -32350 -1224 -32344 -1190
rect -32310 -1224 -32266 -1190
rect -32232 -1224 -32188 -1190
rect -32154 -1224 -32110 -1190
rect -32076 -1224 -32032 -1190
rect -31998 -1224 -31954 -1190
rect -31920 -1224 -31876 -1190
rect -31842 -1224 -31798 -1190
rect -31764 -1224 -31758 -1190
rect -32350 -1262 -31758 -1224
rect -32350 -1296 -32344 -1262
rect -32310 -1296 -32266 -1262
rect -32232 -1296 -32188 -1262
rect -32154 -1296 -32110 -1262
rect -32076 -1296 -32032 -1262
rect -31998 -1296 -31954 -1262
rect -31920 -1296 -31876 -1262
rect -31842 -1296 -31798 -1262
rect -31764 -1296 -31758 -1262
rect -32350 -1334 -31758 -1296
rect -32350 -1368 -32344 -1334
rect -32310 -1368 -32266 -1334
rect -32232 -1368 -32188 -1334
rect -32154 -1368 -32110 -1334
rect -32076 -1368 -32032 -1334
rect -31998 -1368 -31954 -1334
rect -31920 -1368 -31876 -1334
rect -31842 -1368 -31798 -1334
rect -31764 -1368 -31758 -1334
rect -32350 -1406 -31758 -1368
rect -32350 -1440 -32344 -1406
rect -32310 -1440 -32266 -1406
rect -32232 -1440 -32188 -1406
rect -32154 -1440 -32110 -1406
rect -32076 -1440 -32032 -1406
rect -31998 -1440 -31954 -1406
rect -31920 -1440 -31876 -1406
rect -31842 -1440 -31798 -1406
rect -31764 -1440 -31758 -1406
rect -32350 -1478 -31758 -1440
rect -32350 -1512 -32344 -1478
rect -32310 -1512 -32266 -1478
rect -32232 -1512 -32188 -1478
rect -32154 -1512 -32110 -1478
rect -32076 -1512 -32032 -1478
rect -31998 -1512 -31954 -1478
rect -31920 -1512 -31876 -1478
rect -31842 -1512 -31798 -1478
rect -31764 -1512 -31758 -1478
rect -32350 -1550 -31758 -1512
rect -32350 -1584 -32344 -1550
rect -32310 -1584 -32266 -1550
rect -32232 -1584 -32188 -1550
rect -32154 -1584 -32110 -1550
rect -32076 -1584 -32032 -1550
rect -31998 -1584 -31954 -1550
rect -31920 -1584 -31876 -1550
rect -31842 -1584 -31798 -1550
rect -31764 -1584 -31758 -1550
rect -32350 -1622 -31758 -1584
rect -32350 -1656 -32344 -1622
rect -32310 -1656 -32266 -1622
rect -32232 -1656 -32188 -1622
rect -32154 -1656 -32110 -1622
rect -32076 -1656 -32032 -1622
rect -31998 -1656 -31954 -1622
rect -31920 -1656 -31876 -1622
rect -31842 -1656 -31798 -1622
rect -31764 -1656 -31758 -1622
rect -32350 -1694 -31758 -1656
rect -32350 -1728 -32344 -1694
rect -32310 -1728 -32266 -1694
rect -32232 -1728 -32188 -1694
rect -32154 -1728 -32110 -1694
rect -32076 -1728 -32032 -1694
rect -31998 -1728 -31954 -1694
rect -31920 -1728 -31876 -1694
rect -31842 -1728 -31798 -1694
rect -31764 -1728 -31758 -1694
rect -32350 -1766 -31758 -1728
rect -32350 -1800 -32344 -1766
rect -32310 -1800 -32266 -1766
rect -32232 -1800 -32188 -1766
rect -32154 -1800 -32110 -1766
rect -32076 -1800 -32032 -1766
rect -31998 -1800 -31954 -1766
rect -31920 -1800 -31876 -1766
rect -31842 -1800 -31798 -1766
rect -31764 -1800 -31758 -1766
rect -32350 -1838 -31758 -1800
rect -32350 -1872 -32344 -1838
rect -32310 -1872 -32266 -1838
rect -32232 -1872 -32188 -1838
rect -32154 -1872 -32110 -1838
rect -32076 -1872 -32032 -1838
rect -31998 -1872 -31954 -1838
rect -31920 -1872 -31876 -1838
rect -31842 -1872 -31798 -1838
rect -31764 -1872 -31758 -1838
rect -32350 -1910 -31758 -1872
rect -32350 -1944 -32344 -1910
rect -32310 -1944 -32266 -1910
rect -32232 -1944 -32188 -1910
rect -32154 -1944 -32110 -1910
rect -32076 -1944 -32032 -1910
rect -31998 -1944 -31954 -1910
rect -31920 -1944 -31876 -1910
rect -31842 -1944 -31798 -1910
rect -31764 -1944 -31758 -1910
rect -32350 -1982 -31758 -1944
rect -32350 -2016 -32344 -1982
rect -32310 -2016 -32266 -1982
rect -32232 -2016 -32188 -1982
rect -32154 -2016 -32110 -1982
rect -32076 -2016 -32032 -1982
rect -31998 -2016 -31954 -1982
rect -31920 -2016 -31876 -1982
rect -31842 -2016 -31798 -1982
rect -31764 -2016 -31758 -1982
rect -32350 -2054 -31758 -2016
rect -32350 -2088 -32344 -2054
rect -32310 -2088 -32266 -2054
rect -32232 -2088 -32188 -2054
rect -32154 -2088 -32110 -2054
rect -32076 -2088 -32032 -2054
rect -31998 -2088 -31954 -2054
rect -31920 -2088 -31876 -2054
rect -31842 -2088 -31798 -2054
rect -31764 -2088 -31758 -2054
rect -32350 -2126 -31758 -2088
rect -32350 -2160 -32344 -2126
rect -32310 -2160 -32266 -2126
rect -32232 -2160 -32188 -2126
rect -32154 -2160 -32110 -2126
rect -32076 -2160 -32032 -2126
rect -31998 -2160 -31954 -2126
rect -31920 -2160 -31876 -2126
rect -31842 -2160 -31798 -2126
rect -31764 -2160 -31758 -2126
rect -32350 -2198 -31758 -2160
rect -32350 -2232 -32344 -2198
rect -32310 -2232 -32266 -2198
rect -32232 -2232 -32188 -2198
rect -32154 -2232 -32110 -2198
rect -32076 -2232 -32032 -2198
rect -31998 -2232 -31954 -2198
rect -31920 -2232 -31876 -2198
rect -31842 -2232 -31798 -2198
rect -31764 -2232 -31758 -2198
rect -32350 -2270 -31758 -2232
rect -32350 -2304 -32344 -2270
rect -32310 -2304 -32266 -2270
rect -32232 -2304 -32188 -2270
rect -32154 -2304 -32110 -2270
rect -32076 -2304 -32032 -2270
rect -31998 -2304 -31954 -2270
rect -31920 -2304 -31876 -2270
rect -31842 -2304 -31798 -2270
rect -31764 -2304 -31758 -2270
rect -32350 -2342 -31758 -2304
rect -32350 -2376 -32344 -2342
rect -32310 -2376 -32266 -2342
rect -32232 -2376 -32188 -2342
rect -32154 -2376 -32110 -2342
rect -32076 -2376 -32032 -2342
rect -31998 -2376 -31954 -2342
rect -31920 -2376 -31876 -2342
rect -31842 -2376 -31798 -2342
rect -31764 -2376 -31758 -2342
rect -32350 -2414 -31758 -2376
rect -32350 -2448 -32344 -2414
rect -32310 -2448 -32266 -2414
rect -32232 -2448 -32188 -2414
rect -32154 -2448 -32110 -2414
rect -32076 -2448 -32032 -2414
rect -31998 -2448 -31954 -2414
rect -31920 -2448 -31876 -2414
rect -31842 -2448 -31798 -2414
rect -31764 -2448 -31758 -2414
rect -32350 -2486 -31758 -2448
rect -32350 -2520 -32344 -2486
rect -32310 -2520 -32266 -2486
rect -32232 -2520 -32188 -2486
rect -32154 -2520 -32110 -2486
rect -32076 -2520 -32032 -2486
rect -31998 -2520 -31954 -2486
rect -31920 -2520 -31876 -2486
rect -31842 -2520 -31798 -2486
rect -31764 -2520 -31758 -2486
rect -32350 -2558 -31758 -2520
rect -32350 -2592 -32344 -2558
rect -32310 -2592 -32266 -2558
rect -32232 -2592 -32188 -2558
rect -32154 -2592 -32110 -2558
rect -32076 -2592 -32032 -2558
rect -31998 -2592 -31954 -2558
rect -31920 -2592 -31876 -2558
rect -31842 -2592 -31798 -2558
rect -31764 -2592 -31758 -2558
rect -32350 -2630 -31758 -2592
rect -32350 -2664 -32344 -2630
rect -32310 -2664 -32266 -2630
rect -32232 -2664 -32188 -2630
rect -32154 -2664 -32110 -2630
rect -32076 -2664 -32032 -2630
rect -31998 -2664 -31954 -2630
rect -31920 -2664 -31876 -2630
rect -31842 -2664 -31798 -2630
rect -31764 -2664 -31758 -2630
rect -32350 -2702 -31758 -2664
rect -32350 -2736 -32344 -2702
rect -32310 -2736 -32266 -2702
rect -32232 -2736 -32188 -2702
rect -32154 -2736 -32110 -2702
rect -32076 -2736 -32032 -2702
rect -31998 -2736 -31954 -2702
rect -31920 -2736 -31876 -2702
rect -31842 -2736 -31798 -2702
rect -31764 -2736 -31758 -2702
rect -32350 -2774 -31758 -2736
rect -32350 -2808 -32344 -2774
rect -32310 -2808 -32266 -2774
rect -32232 -2808 -32188 -2774
rect -32154 -2808 -32110 -2774
rect -32076 -2808 -32032 -2774
rect -31998 -2808 -31954 -2774
rect -31920 -2808 -31876 -2774
rect -31842 -2808 -31798 -2774
rect -31764 -2808 -31758 -2774
rect -32350 -2846 -31758 -2808
rect -32350 -2880 -32344 -2846
rect -32310 -2880 -32266 -2846
rect -32232 -2880 -32188 -2846
rect -32154 -2880 -32110 -2846
rect -32076 -2880 -32032 -2846
rect -31998 -2880 -31954 -2846
rect -31920 -2880 -31876 -2846
rect -31842 -2880 -31798 -2846
rect -31764 -2880 -31758 -2846
rect -32350 -2918 -31758 -2880
rect -32350 -2952 -32344 -2918
rect -32310 -2952 -32266 -2918
rect -32232 -2952 -32188 -2918
rect -32154 -2952 -32110 -2918
rect -32076 -2952 -32032 -2918
rect -31998 -2952 -31954 -2918
rect -31920 -2952 -31876 -2918
rect -31842 -2952 -31798 -2918
rect -31764 -2952 -31758 -2918
rect -32350 -2990 -31758 -2952
rect -32350 -3024 -32344 -2990
rect -32310 -3024 -32266 -2990
rect -32232 -3024 -32188 -2990
rect -32154 -3024 -32110 -2990
rect -32076 -3024 -32032 -2990
rect -31998 -3024 -31954 -2990
rect -31920 -3024 -31876 -2990
rect -31842 -3024 -31798 -2990
rect -31764 -3024 -31758 -2990
rect -32350 -3062 -31758 -3024
rect -32350 -3096 -32344 -3062
rect -32310 -3096 -32266 -3062
rect -32232 -3096 -32188 -3062
rect -32154 -3096 -32110 -3062
rect -32076 -3096 -32032 -3062
rect -31998 -3096 -31954 -3062
rect -31920 -3096 -31876 -3062
rect -31842 -3096 -31798 -3062
rect -31764 -3096 -31758 -3062
rect -32350 -3134 -31758 -3096
rect -32350 -3168 -32344 -3134
rect -32310 -3168 -32266 -3134
rect -32232 -3168 -32188 -3134
rect -32154 -3168 -32110 -3134
rect -32076 -3168 -32032 -3134
rect -31998 -3168 -31954 -3134
rect -31920 -3168 -31876 -3134
rect -31842 -3168 -31798 -3134
rect -31764 -3168 -31758 -3134
rect -32350 -3206 -31758 -3168
rect -32350 -3240 -32344 -3206
rect -32310 -3240 -32266 -3206
rect -32232 -3240 -32188 -3206
rect -32154 -3240 -32110 -3206
rect -32076 -3240 -32032 -3206
rect -31998 -3240 -31954 -3206
rect -31920 -3240 -31876 -3206
rect -31842 -3240 -31798 -3206
rect -31764 -3240 -31758 -3206
rect -32350 -3278 -31758 -3240
rect -32350 -3312 -32344 -3278
rect -32310 -3312 -32266 -3278
rect -32232 -3312 -32188 -3278
rect -32154 -3312 -32110 -3278
rect -32076 -3312 -32032 -3278
rect -31998 -3312 -31954 -3278
rect -31920 -3312 -31876 -3278
rect -31842 -3312 -31798 -3278
rect -31764 -3312 -31758 -3278
rect -32350 -3350 -31758 -3312
rect -32350 -3384 -32344 -3350
rect -32310 -3384 -32266 -3350
rect -32232 -3384 -32188 -3350
rect -32154 -3384 -32110 -3350
rect -32076 -3384 -32032 -3350
rect -31998 -3384 -31954 -3350
rect -31920 -3384 -31876 -3350
rect -31842 -3384 -31798 -3350
rect -31764 -3384 -31758 -3350
rect -32350 -3422 -31758 -3384
rect -32350 -3456 -32344 -3422
rect -32310 -3456 -32266 -3422
rect -32232 -3456 -32188 -3422
rect -32154 -3456 -32110 -3422
rect -32076 -3456 -32032 -3422
rect -31998 -3456 -31954 -3422
rect -31920 -3456 -31876 -3422
rect -31842 -3456 -31798 -3422
rect -31764 -3456 -31758 -3422
rect -32350 -3494 -31758 -3456
rect -32350 -3528 -32344 -3494
rect -32310 -3528 -32266 -3494
rect -32232 -3528 -32188 -3494
rect -32154 -3528 -32110 -3494
rect -32076 -3528 -32032 -3494
rect -31998 -3528 -31954 -3494
rect -31920 -3528 -31876 -3494
rect -31842 -3528 -31798 -3494
rect -31764 -3528 -31758 -3494
rect -32350 -3566 -31758 -3528
rect -32350 -3600 -32344 -3566
rect -32310 -3600 -32266 -3566
rect -32232 -3600 -32188 -3566
rect -32154 -3600 -32110 -3566
rect -32076 -3600 -32032 -3566
rect -31998 -3600 -31954 -3566
rect -31920 -3600 -31876 -3566
rect -31842 -3600 -31798 -3566
rect -31764 -3600 -31758 -3566
rect -32350 -3638 -31758 -3600
rect -32350 -3672 -32344 -3638
rect -32310 -3672 -32266 -3638
rect -32232 -3672 -32188 -3638
rect -32154 -3672 -32110 -3638
rect -32076 -3672 -32032 -3638
rect -31998 -3672 -31954 -3638
rect -31920 -3672 -31876 -3638
rect -31842 -3672 -31798 -3638
rect -31764 -3672 -31758 -3638
rect -32350 -3710 -31758 -3672
rect -32350 -3744 -32344 -3710
rect -32310 -3744 -32266 -3710
rect -32232 -3744 -32188 -3710
rect -32154 -3744 -32110 -3710
rect -32076 -3744 -32032 -3710
rect -31998 -3744 -31954 -3710
rect -31920 -3744 -31876 -3710
rect -31842 -3744 -31798 -3710
rect -31764 -3744 -31758 -3710
rect -32350 -3782 -31758 -3744
rect -32350 -3816 -32344 -3782
rect -32310 -3816 -32266 -3782
rect -32232 -3816 -32188 -3782
rect -32154 -3816 -32110 -3782
rect -32076 -3816 -32032 -3782
rect -31998 -3816 -31954 -3782
rect -31920 -3816 -31876 -3782
rect -31842 -3816 -31798 -3782
rect -31764 -3816 -31758 -3782
rect -32350 -3854 -31758 -3816
rect -32350 -3888 -32344 -3854
rect -32310 -3888 -32266 -3854
rect -32232 -3888 -32188 -3854
rect -32154 -3888 -32110 -3854
rect -32076 -3888 -32032 -3854
rect -31998 -3888 -31954 -3854
rect -31920 -3888 -31876 -3854
rect -31842 -3888 -31798 -3854
rect -31764 -3888 -31758 -3854
rect -32350 -3926 -31758 -3888
rect -32350 -3960 -32344 -3926
rect -32310 -3960 -32266 -3926
rect -32232 -3960 -32188 -3926
rect -32154 -3960 -32110 -3926
rect -32076 -3960 -32032 -3926
rect -31998 -3960 -31954 -3926
rect -31920 -3960 -31876 -3926
rect -31842 -3960 -31798 -3926
rect -31764 -3960 -31758 -3926
rect -32350 -3998 -31758 -3960
rect -32350 -4032 -32344 -3998
rect -32310 -4032 -32266 -3998
rect -32232 -4032 -32188 -3998
rect -32154 -4032 -32110 -3998
rect -32076 -4032 -32032 -3998
rect -31998 -4032 -31954 -3998
rect -31920 -4032 -31876 -3998
rect -31842 -4032 -31798 -3998
rect -31764 -4032 -31758 -3998
rect -32350 -4070 -31758 -4032
rect -32350 -4104 -32344 -4070
rect -32310 -4104 -32266 -4070
rect -32232 -4104 -32188 -4070
rect -32154 -4104 -32110 -4070
rect -32076 -4104 -32032 -4070
rect -31998 -4104 -31954 -4070
rect -31920 -4104 -31876 -4070
rect -31842 -4104 -31798 -4070
rect -31764 -4104 -31758 -4070
rect -32350 -4142 -31758 -4104
rect -32350 -4176 -32344 -4142
rect -32310 -4176 -32266 -4142
rect -32232 -4176 -32188 -4142
rect -32154 -4176 -32110 -4142
rect -32076 -4176 -32032 -4142
rect -31998 -4176 -31954 -4142
rect -31920 -4176 -31876 -4142
rect -31842 -4176 -31798 -4142
rect -31764 -4176 -31758 -4142
rect -32350 -4214 -31758 -4176
rect -32350 -4248 -32344 -4214
rect -32310 -4248 -32266 -4214
rect -32232 -4248 -32188 -4214
rect -32154 -4248 -32110 -4214
rect -32076 -4248 -32032 -4214
rect -31998 -4248 -31954 -4214
rect -31920 -4248 -31876 -4214
rect -31842 -4248 -31798 -4214
rect -31764 -4248 -31758 -4214
rect -32350 -4286 -31758 -4248
rect -32350 -4320 -32344 -4286
rect -32310 -4320 -32266 -4286
rect -32232 -4320 -32188 -4286
rect -32154 -4320 -32110 -4286
rect -32076 -4320 -32032 -4286
rect -31998 -4320 -31954 -4286
rect -31920 -4320 -31876 -4286
rect -31842 -4320 -31798 -4286
rect -31764 -4320 -31758 -4286
rect -32350 -4358 -31758 -4320
rect -32350 -4392 -32344 -4358
rect -32310 -4392 -32266 -4358
rect -32232 -4392 -32188 -4358
rect -32154 -4392 -32110 -4358
rect -32076 -4392 -32032 -4358
rect -31998 -4392 -31954 -4358
rect -31920 -4392 -31876 -4358
rect -31842 -4392 -31798 -4358
rect -31764 -4392 -31758 -4358
rect -32350 -4430 -31758 -4392
rect -32350 -4464 -32344 -4430
rect -32310 -4464 -32266 -4430
rect -32232 -4464 -32188 -4430
rect -32154 -4464 -32110 -4430
rect -32076 -4464 -32032 -4430
rect -31998 -4464 -31954 -4430
rect -31920 -4464 -31876 -4430
rect -31842 -4464 -31798 -4430
rect -31764 -4464 -31758 -4430
rect -32350 -4502 -31758 -4464
rect -32350 -4536 -32344 -4502
rect -32310 -4536 -32266 -4502
rect -32232 -4536 -32188 -4502
rect -32154 -4536 -32110 -4502
rect -32076 -4536 -32032 -4502
rect -31998 -4536 -31954 -4502
rect -31920 -4536 -31876 -4502
rect -31842 -4536 -31798 -4502
rect -31764 -4536 -31758 -4502
rect -32350 -4574 -31758 -4536
rect -32350 -4608 -32344 -4574
rect -32310 -4608 -32266 -4574
rect -32232 -4608 -32188 -4574
rect -32154 -4608 -32110 -4574
rect -32076 -4608 -32032 -4574
rect -31998 -4608 -31954 -4574
rect -31920 -4608 -31876 -4574
rect -31842 -4608 -31798 -4574
rect -31764 -4608 -31758 -4574
rect -32350 -4646 -31758 -4608
rect -32350 -4680 -32344 -4646
rect -32310 -4680 -32266 -4646
rect -32232 -4680 -32188 -4646
rect -32154 -4680 -32110 -4646
rect -32076 -4680 -32032 -4646
rect -31998 -4680 -31954 -4646
rect -31920 -4680 -31876 -4646
rect -31842 -4680 -31798 -4646
rect -31764 -4680 -31758 -4646
rect -32350 -4718 -31758 -4680
rect -32350 -4752 -32344 -4718
rect -32310 -4752 -32266 -4718
rect -32232 -4752 -32188 -4718
rect -32154 -4752 -32110 -4718
rect -32076 -4752 -32032 -4718
rect -31998 -4752 -31954 -4718
rect -31920 -4752 -31876 -4718
rect -31842 -4752 -31798 -4718
rect -31764 -4752 -31758 -4718
rect -32350 -4790 -31758 -4752
rect -32350 -4824 -32344 -4790
rect -32310 -4824 -32266 -4790
rect -32232 -4824 -32188 -4790
rect -32154 -4824 -32110 -4790
rect -32076 -4824 -32032 -4790
rect -31998 -4824 -31954 -4790
rect -31920 -4824 -31876 -4790
rect -31842 -4824 -31798 -4790
rect -31764 -4824 -31758 -4790
rect -32350 -4862 -31758 -4824
rect -32350 -4896 -32344 -4862
rect -32310 -4896 -32266 -4862
rect -32232 -4896 -32188 -4862
rect -32154 -4896 -32110 -4862
rect -32076 -4896 -32032 -4862
rect -31998 -4896 -31954 -4862
rect -31920 -4896 -31876 -4862
rect -31842 -4896 -31798 -4862
rect -31764 -4896 -31758 -4862
rect -32350 -4934 -31758 -4896
rect -32350 -4968 -32344 -4934
rect -32310 -4968 -32266 -4934
rect -32232 -4968 -32188 -4934
rect -32154 -4968 -32110 -4934
rect -32076 -4968 -32032 -4934
rect -31998 -4968 -31954 -4934
rect -31920 -4968 -31876 -4934
rect -31842 -4968 -31798 -4934
rect -31764 -4968 -31758 -4934
rect -32350 -5006 -31758 -4968
rect -32350 -5040 -32344 -5006
rect -32310 -5040 -32266 -5006
rect -32232 -5040 -32188 -5006
rect -32154 -5040 -32110 -5006
rect -32076 -5040 -32032 -5006
rect -31998 -5040 -31954 -5006
rect -31920 -5040 -31876 -5006
rect -31842 -5040 -31798 -5006
rect -31764 -5040 -31758 -5006
rect -32350 -5078 -31758 -5040
rect -32350 -5112 -32344 -5078
rect -32310 -5112 -32266 -5078
rect -32232 -5112 -32188 -5078
rect -32154 -5112 -32110 -5078
rect -32076 -5112 -32032 -5078
rect -31998 -5112 -31954 -5078
rect -31920 -5112 -31876 -5078
rect -31842 -5112 -31798 -5078
rect -31764 -5112 -31758 -5078
rect -32350 -5150 -31758 -5112
rect -32350 -5184 -32344 -5150
rect -32310 -5184 -32266 -5150
rect -32232 -5184 -32188 -5150
rect -32154 -5184 -32110 -5150
rect -32076 -5184 -32032 -5150
rect -31998 -5184 -31954 -5150
rect -31920 -5184 -31876 -5150
rect -31842 -5184 -31798 -5150
rect -31764 -5184 -31758 -5150
rect -32350 -5222 -31758 -5184
rect -32350 -5256 -32344 -5222
rect -32310 -5256 -32266 -5222
rect -32232 -5256 -32188 -5222
rect -32154 -5256 -32110 -5222
rect -32076 -5256 -32032 -5222
rect -31998 -5256 -31954 -5222
rect -31920 -5256 -31876 -5222
rect -31842 -5256 -31798 -5222
rect -31764 -5256 -31758 -5222
rect -32350 -5294 -31758 -5256
rect -32350 -5328 -32344 -5294
rect -32310 -5328 -32266 -5294
rect -32232 -5328 -32188 -5294
rect -32154 -5328 -32110 -5294
rect -32076 -5328 -32032 -5294
rect -31998 -5328 -31954 -5294
rect -31920 -5328 -31876 -5294
rect -31842 -5328 -31798 -5294
rect -31764 -5328 -31758 -5294
rect -32350 -5366 -31758 -5328
rect -32350 -5400 -32344 -5366
rect -32310 -5400 -32266 -5366
rect -32232 -5400 -32188 -5366
rect -32154 -5400 -32110 -5366
rect -32076 -5400 -32032 -5366
rect -31998 -5400 -31954 -5366
rect -31920 -5400 -31876 -5366
rect -31842 -5400 -31798 -5366
rect -31764 -5400 -31758 -5366
rect -32350 -5438 -31758 -5400
rect -32350 -5472 -32344 -5438
rect -32310 -5472 -32266 -5438
rect -32232 -5472 -32188 -5438
rect -32154 -5472 -32110 -5438
rect -32076 -5472 -32032 -5438
rect -31998 -5472 -31954 -5438
rect -31920 -5472 -31876 -5438
rect -31842 -5472 -31798 -5438
rect -31764 -5472 -31758 -5438
rect -32350 -5510 -31758 -5472
rect -32350 -5544 -32344 -5510
rect -32310 -5544 -32266 -5510
rect -32232 -5544 -32188 -5510
rect -32154 -5544 -32110 -5510
rect -32076 -5544 -32032 -5510
rect -31998 -5544 -31954 -5510
rect -31920 -5544 -31876 -5510
rect -31842 -5544 -31798 -5510
rect -31764 -5544 -31758 -5510
rect -32350 -5582 -31758 -5544
rect -32350 -5616 -32344 -5582
rect -32310 -5616 -32266 -5582
rect -32232 -5616 -32188 -5582
rect -32154 -5616 -32110 -5582
rect -32076 -5616 -32032 -5582
rect -31998 -5616 -31954 -5582
rect -31920 -5616 -31876 -5582
rect -31842 -5616 -31798 -5582
rect -31764 -5616 -31758 -5582
rect -32350 -5654 -31758 -5616
rect -32350 -5688 -32344 -5654
rect -32310 -5688 -32266 -5654
rect -32232 -5688 -32188 -5654
rect -32154 -5688 -32110 -5654
rect -32076 -5688 -32032 -5654
rect -31998 -5688 -31954 -5654
rect -31920 -5688 -31876 -5654
rect -31842 -5688 -31798 -5654
rect -31764 -5688 -31758 -5654
rect -32350 -5726 -31758 -5688
rect -32350 -5760 -32344 -5726
rect -32310 -5760 -32266 -5726
rect -32232 -5760 -32188 -5726
rect -32154 -5760 -32110 -5726
rect -32076 -5760 -32032 -5726
rect -31998 -5760 -31954 -5726
rect -31920 -5760 -31876 -5726
rect -31842 -5760 -31798 -5726
rect -31764 -5760 -31758 -5726
rect -32350 -5798 -31758 -5760
rect -32350 -5832 -32344 -5798
rect -32310 -5832 -32266 -5798
rect -32232 -5832 -32188 -5798
rect -32154 -5832 -32110 -5798
rect -32076 -5832 -32032 -5798
rect -31998 -5832 -31954 -5798
rect -31920 -5832 -31876 -5798
rect -31842 -5832 -31798 -5798
rect -31764 -5832 -31758 -5798
rect -32350 -5870 -31758 -5832
rect -32350 -5904 -32344 -5870
rect -32310 -5904 -32266 -5870
rect -32232 -5904 -32188 -5870
rect -32154 -5904 -32110 -5870
rect -32076 -5904 -32032 -5870
rect -31998 -5904 -31954 -5870
rect -31920 -5904 -31876 -5870
rect -31842 -5904 -31798 -5870
rect -31764 -5904 -31758 -5870
rect -32350 -5942 -31758 -5904
rect -32350 -5976 -32344 -5942
rect -32310 -5976 -32266 -5942
rect -32232 -5976 -32188 -5942
rect -32154 -5976 -32110 -5942
rect -32076 -5976 -32032 -5942
rect -31998 -5976 -31954 -5942
rect -31920 -5976 -31876 -5942
rect -31842 -5976 -31798 -5942
rect -31764 -5976 -31758 -5942
rect -32350 -6014 -31758 -5976
rect -32350 -6048 -32344 -6014
rect -32310 -6048 -32266 -6014
rect -32232 -6048 -32188 -6014
rect -32154 -6048 -32110 -6014
rect -32076 -6048 -32032 -6014
rect -31998 -6048 -31954 -6014
rect -31920 -6048 -31876 -6014
rect -31842 -6048 -31798 -6014
rect -31764 -6048 -31758 -6014
rect -32350 -6086 -31758 -6048
rect -32350 -6120 -32344 -6086
rect -32310 -6120 -32266 -6086
rect -32232 -6120 -32188 -6086
rect -32154 -6120 -32110 -6086
rect -32076 -6120 -32032 -6086
rect -31998 -6120 -31954 -6086
rect -31920 -6120 -31876 -6086
rect -31842 -6120 -31798 -6086
rect -31764 -6120 -31758 -6086
rect -32350 -6158 -31758 -6120
rect -32350 -6192 -32344 -6158
rect -32310 -6192 -32266 -6158
rect -32232 -6192 -32188 -6158
rect -32154 -6192 -32110 -6158
rect -32076 -6192 -32032 -6158
rect -31998 -6192 -31954 -6158
rect -31920 -6192 -31876 -6158
rect -31842 -6192 -31798 -6158
rect -31764 -6192 -31758 -6158
rect -32350 -6230 -31758 -6192
rect -32350 -6264 -32344 -6230
rect -32310 -6264 -32266 -6230
rect -32232 -6264 -32188 -6230
rect -32154 -6264 -32110 -6230
rect -32076 -6264 -32032 -6230
rect -31998 -6264 -31954 -6230
rect -31920 -6264 -31876 -6230
rect -31842 -6264 -31798 -6230
rect -31764 -6264 -31758 -6230
rect -32350 -6302 -31758 -6264
rect -32350 -6336 -32344 -6302
rect -32310 -6336 -32266 -6302
rect -32232 -6336 -32188 -6302
rect -32154 -6336 -32110 -6302
rect -32076 -6336 -32032 -6302
rect -31998 -6336 -31954 -6302
rect -31920 -6336 -31876 -6302
rect -31842 -6336 -31798 -6302
rect -31764 -6336 -31758 -6302
rect -32350 -6374 -31758 -6336
rect -32350 -6408 -32344 -6374
rect -32310 -6408 -32266 -6374
rect -32232 -6408 -32188 -6374
rect -32154 -6408 -32110 -6374
rect -32076 -6408 -32032 -6374
rect -31998 -6408 -31954 -6374
rect -31920 -6408 -31876 -6374
rect -31842 -6408 -31798 -6374
rect -31764 -6408 -31758 -6374
rect -32350 -6446 -31758 -6408
rect -32350 -6480 -32344 -6446
rect -32310 -6480 -32266 -6446
rect -32232 -6480 -32188 -6446
rect -32154 -6480 -32110 -6446
rect -32076 -6480 -32032 -6446
rect -31998 -6480 -31954 -6446
rect -31920 -6480 -31876 -6446
rect -31842 -6480 -31798 -6446
rect -31764 -6480 -31758 -6446
rect -32350 -6518 -31758 -6480
rect -32350 -6552 -32344 -6518
rect -32310 -6552 -32266 -6518
rect -32232 -6552 -32188 -6518
rect -32154 -6552 -32110 -6518
rect -32076 -6552 -32032 -6518
rect -31998 -6552 -31954 -6518
rect -31920 -6552 -31876 -6518
rect -31842 -6552 -31798 -6518
rect -31764 -6552 -31758 -6518
rect -32350 -6590 -31758 -6552
rect -32350 -6624 -32344 -6590
rect -32310 -6624 -32266 -6590
rect -32232 -6624 -32188 -6590
rect -32154 -6624 -32110 -6590
rect -32076 -6624 -32032 -6590
rect -31998 -6624 -31954 -6590
rect -31920 -6624 -31876 -6590
rect -31842 -6624 -31798 -6590
rect -31764 -6624 -31758 -6590
rect -32350 -6662 -31758 -6624
rect -32350 -6696 -32344 -6662
rect -32310 -6696 -32266 -6662
rect -32232 -6696 -32188 -6662
rect -32154 -6696 -32110 -6662
rect -32076 -6696 -32032 -6662
rect -31998 -6696 -31954 -6662
rect -31920 -6696 -31876 -6662
rect -31842 -6696 -31798 -6662
rect -31764 -6696 -31758 -6662
rect -32350 -6734 -31758 -6696
rect -32350 -6768 -32344 -6734
rect -32310 -6768 -32266 -6734
rect -32232 -6768 -32188 -6734
rect -32154 -6768 -32110 -6734
rect -32076 -6768 -32032 -6734
rect -31998 -6768 -31954 -6734
rect -31920 -6768 -31876 -6734
rect -31842 -6768 -31798 -6734
rect -31764 -6768 -31758 -6734
rect -32350 -6806 -31758 -6768
rect -32350 -6840 -32344 -6806
rect -32310 -6840 -32266 -6806
rect -32232 -6840 -32188 -6806
rect -32154 -6840 -32110 -6806
rect -32076 -6840 -32032 -6806
rect -31998 -6840 -31954 -6806
rect -31920 -6840 -31876 -6806
rect -31842 -6840 -31798 -6806
rect -31764 -6840 -31758 -6806
rect -32350 -6878 -31758 -6840
rect -32350 -6912 -32344 -6878
rect -32310 -6912 -32266 -6878
rect -32232 -6912 -32188 -6878
rect -32154 -6912 -32110 -6878
rect -32076 -6912 -32032 -6878
rect -31998 -6912 -31954 -6878
rect -31920 -6912 -31876 -6878
rect -31842 -6912 -31798 -6878
rect -31764 -6912 -31758 -6878
rect -32350 -6950 -31758 -6912
rect -32350 -6984 -32344 -6950
rect -32310 -6984 -32266 -6950
rect -32232 -6984 -32188 -6950
rect -32154 -6984 -32110 -6950
rect -32076 -6984 -32032 -6950
rect -31998 -6984 -31954 -6950
rect -31920 -6984 -31876 -6950
rect -31842 -6984 -31798 -6950
rect -31764 -6984 -31758 -6950
rect -32350 -7022 -31758 -6984
rect -32350 -7056 -32344 -7022
rect -32310 -7056 -32266 -7022
rect -32232 -7056 -32188 -7022
rect -32154 -7056 -32110 -7022
rect -32076 -7056 -32032 -7022
rect -31998 -7056 -31954 -7022
rect -31920 -7056 -31876 -7022
rect -31842 -7056 -31798 -7022
rect -31764 -7056 -31758 -7022
rect -32350 -7094 -31758 -7056
rect -32350 -7128 -32344 -7094
rect -32310 -7128 -32266 -7094
rect -32232 -7128 -32188 -7094
rect -32154 -7128 -32110 -7094
rect -32076 -7128 -32032 -7094
rect -31998 -7128 -31954 -7094
rect -31920 -7128 -31876 -7094
rect -31842 -7128 -31798 -7094
rect -31764 -7128 -31758 -7094
rect -32350 -7166 -31758 -7128
rect -32350 -7200 -32344 -7166
rect -32310 -7200 -32266 -7166
rect -32232 -7200 -32188 -7166
rect -32154 -7200 -32110 -7166
rect -32076 -7200 -32032 -7166
rect -31998 -7200 -31954 -7166
rect -31920 -7200 -31876 -7166
rect -31842 -7200 -31798 -7166
rect -31764 -7200 -31758 -7166
rect -32350 -7238 -31758 -7200
rect -32350 -7272 -32344 -7238
rect -32310 -7272 -32266 -7238
rect -32232 -7272 -32188 -7238
rect -32154 -7272 -32110 -7238
rect -32076 -7272 -32032 -7238
rect -31998 -7272 -31954 -7238
rect -31920 -7272 -31876 -7238
rect -31842 -7272 -31798 -7238
rect -31764 -7272 -31758 -7238
rect -32350 -7310 -31758 -7272
rect -32350 -7344 -32344 -7310
rect -32310 -7344 -32266 -7310
rect -32232 -7344 -32188 -7310
rect -32154 -7344 -32110 -7310
rect -32076 -7344 -32032 -7310
rect -31998 -7344 -31954 -7310
rect -31920 -7344 -31876 -7310
rect -31842 -7344 -31798 -7310
rect -31764 -7344 -31758 -7310
rect -32350 -7382 -31758 -7344
rect -32350 -7416 -32344 -7382
rect -32310 -7416 -32266 -7382
rect -32232 -7416 -32188 -7382
rect -32154 -7416 -32110 -7382
rect -32076 -7416 -32032 -7382
rect -31998 -7416 -31954 -7382
rect -31920 -7416 -31876 -7382
rect -31842 -7416 -31798 -7382
rect -31764 -7416 -31758 -7382
rect -32350 -7454 -31758 -7416
rect -32350 -7488 -32344 -7454
rect -32310 -7488 -32266 -7454
rect -32232 -7488 -32188 -7454
rect -32154 -7488 -32110 -7454
rect -32076 -7488 -32032 -7454
rect -31998 -7488 -31954 -7454
rect -31920 -7488 -31876 -7454
rect -31842 -7488 -31798 -7454
rect -31764 -7488 -31758 -7454
rect -32350 -7526 -31758 -7488
rect -32350 -7560 -32344 -7526
rect -32310 -7560 -32266 -7526
rect -32232 -7560 -32188 -7526
rect -32154 -7560 -32110 -7526
rect -32076 -7560 -32032 -7526
rect -31998 -7560 -31954 -7526
rect -31920 -7560 -31876 -7526
rect -31842 -7560 -31798 -7526
rect -31764 -7560 -31758 -7526
rect -32350 -7598 -31758 -7560
rect -32350 -7632 -32344 -7598
rect -32310 -7632 -32266 -7598
rect -32232 -7632 -32188 -7598
rect -32154 -7632 -32110 -7598
rect -32076 -7632 -32032 -7598
rect -31998 -7632 -31954 -7598
rect -31920 -7632 -31876 -7598
rect -31842 -7632 -31798 -7598
rect -31764 -7632 -31758 -7598
rect -32350 -7670 -31758 -7632
rect -32350 -7704 -32344 -7670
rect -32310 -7704 -32266 -7670
rect -32232 -7704 -32188 -7670
rect -32154 -7704 -32110 -7670
rect -32076 -7704 -32032 -7670
rect -31998 -7704 -31954 -7670
rect -31920 -7704 -31876 -7670
rect -31842 -7704 -31798 -7670
rect -31764 -7704 -31758 -7670
rect -32350 -7742 -31758 -7704
rect -32350 -7776 -32344 -7742
rect -32310 -7776 -32266 -7742
rect -32232 -7776 -32188 -7742
rect -32154 -7776 -32110 -7742
rect -32076 -7776 -32032 -7742
rect -31998 -7776 -31954 -7742
rect -31920 -7776 -31876 -7742
rect -31842 -7776 -31798 -7742
rect -31764 -7776 -31758 -7742
rect -32350 -7814 -31758 -7776
rect -32350 -7848 -32344 -7814
rect -32310 -7848 -32266 -7814
rect -32232 -7848 -32188 -7814
rect -32154 -7848 -32110 -7814
rect -32076 -7848 -32032 -7814
rect -31998 -7848 -31954 -7814
rect -31920 -7848 -31876 -7814
rect -31842 -7848 -31798 -7814
rect -31764 -7848 -31758 -7814
rect -32350 -7886 -31758 -7848
rect -32350 -7920 -32344 -7886
rect -32310 -7920 -32266 -7886
rect -32232 -7920 -32188 -7886
rect -32154 -7920 -32110 -7886
rect -32076 -7920 -32032 -7886
rect -31998 -7920 -31954 -7886
rect -31920 -7920 -31876 -7886
rect -31842 -7920 -31798 -7886
rect -31764 -7920 -31758 -7886
rect -32350 -7958 -31758 -7920
rect -32350 -7992 -32344 -7958
rect -32310 -7992 -32266 -7958
rect -32232 -7992 -32188 -7958
rect -32154 -7992 -32110 -7958
rect -32076 -7992 -32032 -7958
rect -31998 -7992 -31954 -7958
rect -31920 -7992 -31876 -7958
rect -31842 -7992 -31798 -7958
rect -31764 -7992 -31758 -7958
rect -32350 -8030 -31758 -7992
rect -32350 -8064 -32344 -8030
rect -32310 -8064 -32266 -8030
rect -32232 -8064 -32188 -8030
rect -32154 -8064 -32110 -8030
rect -32076 -8064 -32032 -8030
rect -31998 -8064 -31954 -8030
rect -31920 -8064 -31876 -8030
rect -31842 -8064 -31798 -8030
rect -31764 -8064 -31758 -8030
rect -32350 -8102 -31758 -8064
rect -32350 -8136 -32344 -8102
rect -32310 -8136 -32266 -8102
rect -32232 -8136 -32188 -8102
rect -32154 -8136 -32110 -8102
rect -32076 -8136 -32032 -8102
rect -31998 -8136 -31954 -8102
rect -31920 -8136 -31876 -8102
rect -31842 -8136 -31798 -8102
rect -31764 -8136 -31758 -8102
rect -32350 -8174 -31758 -8136
rect -32350 -8208 -32344 -8174
rect -32310 -8208 -32266 -8174
rect -32232 -8208 -32188 -8174
rect -32154 -8208 -32110 -8174
rect -32076 -8208 -32032 -8174
rect -31998 -8208 -31954 -8174
rect -31920 -8208 -31876 -8174
rect -31842 -8208 -31798 -8174
rect -31764 -8208 -31758 -8174
rect -32350 -8246 -31758 -8208
rect -32350 -8280 -32344 -8246
rect -32310 -8280 -32266 -8246
rect -32232 -8280 -32188 -8246
rect -32154 -8280 -32110 -8246
rect -32076 -8280 -32032 -8246
rect -31998 -8280 -31954 -8246
rect -31920 -8280 -31876 -8246
rect -31842 -8280 -31798 -8246
rect -31764 -8280 -31758 -8246
rect -32350 -8318 -31758 -8280
rect -32350 -8352 -32344 -8318
rect -32310 -8352 -32266 -8318
rect -32232 -8352 -32188 -8318
rect -32154 -8352 -32110 -8318
rect -32076 -8352 -32032 -8318
rect -31998 -8352 -31954 -8318
rect -31920 -8352 -31876 -8318
rect -31842 -8352 -31798 -8318
rect -31764 -8352 -31758 -8318
rect -32350 -8390 -31758 -8352
rect -32350 -8424 -32344 -8390
rect -32310 -8424 -32266 -8390
rect -32232 -8424 -32188 -8390
rect -32154 -8424 -32110 -8390
rect -32076 -8424 -32032 -8390
rect -31998 -8424 -31954 -8390
rect -31920 -8424 -31876 -8390
rect -31842 -8424 -31798 -8390
rect -31764 -8424 -31758 -8390
rect -32350 -8462 -31758 -8424
rect -32350 -8496 -32344 -8462
rect -32310 -8496 -32266 -8462
rect -32232 -8496 -32188 -8462
rect -32154 -8496 -32110 -8462
rect -32076 -8496 -32032 -8462
rect -31998 -8496 -31954 -8462
rect -31920 -8496 -31876 -8462
rect -31842 -8496 -31798 -8462
rect -31764 -8496 -31758 -8462
rect -32350 -8534 -31758 -8496
rect -32350 -8568 -32344 -8534
rect -32310 -8568 -32266 -8534
rect -32232 -8568 -32188 -8534
rect -32154 -8568 -32110 -8534
rect -32076 -8568 -32032 -8534
rect -31998 -8568 -31954 -8534
rect -31920 -8568 -31876 -8534
rect -31842 -8568 -31798 -8534
rect -31764 -8568 -31758 -8534
rect -32350 -8606 -31758 -8568
rect -29140 2800 -28830 2839
rect -29140 2766 -29134 2800
rect -29100 2766 -29046 2800
rect -29012 2766 -28958 2800
rect -28924 2766 -28870 2800
rect -28836 2766 -28830 2800
rect -29140 2727 -28830 2766
rect -29140 2693 -29134 2727
rect -29100 2693 -29046 2727
rect -29012 2693 -28958 2727
rect -28924 2693 -28870 2727
rect -28836 2693 -28830 2727
rect -29140 2654 -28830 2693
rect -29140 2620 -29134 2654
rect -29100 2620 -29046 2654
rect -29012 2620 -28958 2654
rect -28924 2620 -28870 2654
rect -28836 2620 -28830 2654
rect -29140 2581 -28830 2620
rect -29140 2547 -29134 2581
rect -29100 2547 -29046 2581
rect -29012 2547 -28958 2581
rect -28924 2547 -28870 2581
rect -28836 2547 -28830 2581
rect -29140 2508 -28830 2547
rect -29140 2474 -29134 2508
rect -29100 2474 -29046 2508
rect -29012 2474 -28958 2508
rect -28924 2474 -28870 2508
rect -28836 2474 -28830 2508
rect -29140 2435 -28830 2474
rect -29140 2401 -29134 2435
rect -29100 2401 -29046 2435
rect -29012 2401 -28958 2435
rect -28924 2401 -28870 2435
rect -28836 2401 -28830 2435
rect -29140 2362 -28830 2401
rect -29140 2328 -29134 2362
rect -29100 2328 -29046 2362
rect -29012 2328 -28958 2362
rect -28924 2328 -28870 2362
rect -28836 2328 -28830 2362
rect -29140 2289 -28830 2328
rect -29140 2255 -29134 2289
rect -29100 2255 -29046 2289
rect -29012 2255 -28958 2289
rect -28924 2255 -28870 2289
rect -28836 2255 -28830 2289
rect -29140 2216 -28830 2255
rect -29140 2182 -29134 2216
rect -29100 2182 -29046 2216
rect -29012 2182 -28958 2216
rect -28924 2182 -28870 2216
rect -28836 2182 -28830 2216
rect -29140 2143 -28830 2182
rect -29140 2109 -29134 2143
rect -29100 2109 -29046 2143
rect -29012 2109 -28958 2143
rect -28924 2109 -28870 2143
rect -28836 2109 -28830 2143
rect -29140 2070 -28830 2109
rect -29140 2036 -29134 2070
rect -29100 2036 -29046 2070
rect -29012 2036 -28958 2070
rect -28924 2036 -28870 2070
rect -28836 2036 -28830 2070
rect -29140 1997 -28830 2036
rect -29140 1963 -29134 1997
rect -29100 1963 -29046 1997
rect -29012 1963 -28958 1997
rect -28924 1963 -28870 1997
rect -28836 1963 -28830 1997
rect -29140 1924 -28830 1963
rect -29140 1890 -29134 1924
rect -29100 1890 -29046 1924
rect -29012 1890 -28958 1924
rect -28924 1890 -28870 1924
rect -28836 1890 -28830 1924
rect -29140 1851 -28830 1890
rect -29140 1817 -29134 1851
rect -29100 1817 -29046 1851
rect -29012 1817 -28958 1851
rect -28924 1817 -28870 1851
rect -28836 1817 -28830 1851
rect -29140 1778 -28830 1817
rect -29140 1744 -29134 1778
rect -29100 1744 -29046 1778
rect -29012 1744 -28958 1778
rect -28924 1744 -28870 1778
rect -28836 1744 -28830 1778
rect -29140 1705 -28830 1744
rect -29140 1671 -29134 1705
rect -29100 1671 -29046 1705
rect -29012 1671 -28958 1705
rect -28924 1671 -28870 1705
rect -28836 1671 -28830 1705
rect -29140 1632 -28830 1671
rect -29140 1598 -29134 1632
rect -29100 1598 -29046 1632
rect -29012 1598 -28958 1632
rect -28924 1598 -28870 1632
rect -28836 1598 -28830 1632
rect -29140 1559 -28830 1598
rect -29140 1525 -29134 1559
rect -29100 1525 -29046 1559
rect -29012 1525 -28958 1559
rect -28924 1525 -28870 1559
rect -28836 1525 -28830 1559
rect -29140 1486 -28830 1525
rect -29140 1452 -29134 1486
rect -29100 1452 -29046 1486
rect -29012 1452 -28958 1486
rect -28924 1452 -28870 1486
rect -28836 1452 -28830 1486
rect -29140 1413 -28830 1452
rect -29140 1379 -29134 1413
rect -29100 1379 -29046 1413
rect -29012 1379 -28958 1413
rect -28924 1379 -28870 1413
rect -28836 1379 -28830 1413
rect -29140 1340 -28830 1379
rect -29140 1306 -29134 1340
rect -29100 1306 -29046 1340
rect -29012 1306 -28958 1340
rect -28924 1306 -28870 1340
rect -28836 1306 -28830 1340
rect -29140 1267 -28830 1306
rect -29140 1233 -29134 1267
rect -29100 1233 -29046 1267
rect -29012 1233 -28958 1267
rect -28924 1233 -28870 1267
rect -28836 1233 -28830 1267
rect -29140 1194 -28830 1233
rect -29140 1160 -29134 1194
rect -29100 1160 -29046 1194
rect -29012 1160 -28958 1194
rect -28924 1160 -28870 1194
rect -28836 1160 -28830 1194
rect -29140 1121 -28830 1160
rect -29140 1087 -29134 1121
rect -29100 1087 -29046 1121
rect -29012 1087 -28958 1121
rect -28924 1087 -28870 1121
rect -28836 1087 -28830 1121
rect -29140 1048 -28830 1087
rect -29140 1014 -29134 1048
rect -29100 1014 -29046 1048
rect -29012 1014 -28958 1048
rect -28924 1014 -28870 1048
rect -28836 1014 -28830 1048
rect -29140 975 -28830 1014
rect -29140 941 -29134 975
rect -29100 941 -29046 975
rect -29012 941 -28958 975
rect -28924 941 -28870 975
rect -28836 941 -28830 975
rect -29140 902 -28830 941
rect -29140 868 -29134 902
rect -29100 868 -29046 902
rect -29012 868 -28958 902
rect -28924 868 -28870 902
rect -28836 868 -28830 902
rect -29140 829 -28830 868
rect -29140 795 -29134 829
rect -29100 795 -29046 829
rect -29012 795 -28958 829
rect -28924 795 -28870 829
rect -28836 795 -28830 829
rect -29140 756 -28830 795
rect -29140 722 -29134 756
rect -29100 722 -29046 756
rect -29012 722 -28958 756
rect -28924 722 -28870 756
rect -28836 722 -28830 756
rect -29140 683 -28830 722
rect -29140 649 -29134 683
rect -29100 649 -29046 683
rect -29012 649 -28958 683
rect -28924 649 -28870 683
rect -28836 649 -28830 683
rect -29140 610 -28830 649
rect -29140 576 -29134 610
rect -29100 576 -29046 610
rect -29012 576 -28958 610
rect -28924 576 -28870 610
rect -28836 576 -28830 610
rect -29140 537 -28830 576
rect -29140 503 -29134 537
rect -29100 503 -29046 537
rect -29012 503 -28958 537
rect -28924 503 -28870 537
rect -28836 503 -28830 537
rect -29140 495 -28830 503
rect -29140 443 -29135 495
rect -29083 443 -29053 495
rect -29001 443 -28971 495
rect -28919 443 -28889 495
rect -28837 464 -28830 495
rect -29140 430 -29134 443
rect -29100 430 -29046 443
rect -29012 430 -28958 443
rect -28924 430 -28870 443
rect -28836 430 -28830 464
rect -29140 378 -29135 430
rect -29083 378 -29053 430
rect -29001 378 -28971 430
rect -28919 378 -28889 430
rect -28837 391 -28830 430
rect -29140 365 -29134 378
rect -29100 365 -29046 378
rect -29012 365 -28958 378
rect -28924 365 -28870 378
rect -29140 313 -29135 365
rect -29083 313 -29053 365
rect -29001 313 -28971 365
rect -28919 313 -28889 365
rect -28836 357 -28830 391
rect -28837 318 -28830 357
rect -29140 301 -29134 313
rect -29100 301 -29046 313
rect -29012 301 -28958 313
rect -28924 301 -28870 313
rect -29140 249 -29135 301
rect -29083 249 -29053 301
rect -29001 249 -28971 301
rect -28919 249 -28889 301
rect -28836 284 -28830 318
rect -28837 249 -28830 284
rect -29140 245 -28830 249
rect -29140 237 -29134 245
rect -29100 237 -29046 245
rect -29012 237 -28958 245
rect -28924 237 -28870 245
rect -29140 185 -29135 237
rect -29083 185 -29053 237
rect -29001 185 -28971 237
rect -28919 185 -28889 237
rect -28836 211 -28830 245
rect -28837 185 -28830 211
rect -29140 173 -28830 185
rect -29140 121 -29135 173
rect -29083 121 -29053 173
rect -29001 121 -28971 173
rect -28919 121 -28889 173
rect -28837 172 -28830 173
rect -28836 138 -28830 172
rect -28837 121 -28830 138
rect -29140 109 -28830 121
rect -29140 57 -29135 109
rect -29083 57 -29053 109
rect -29001 57 -28971 109
rect -28919 57 -28889 109
rect -28837 99 -28830 109
rect -28836 65 -28830 99
rect -28837 57 -28830 65
rect -29140 45 -28830 57
rect -29140 -7 -29135 45
rect -29083 -7 -29053 45
rect -29001 -7 -28971 45
rect -28919 -7 -28889 45
rect -28837 26 -28830 45
rect -29140 -8 -29134 -7
rect -29100 -8 -29046 -7
rect -29012 -8 -28958 -7
rect -28924 -8 -28870 -7
rect -28836 -8 -28830 26
rect -29140 -19 -28830 -8
rect -29140 -71 -29135 -19
rect -29083 -71 -29053 -19
rect -29001 -71 -28971 -19
rect -28919 -71 -28889 -19
rect -28837 -47 -28830 -19
rect -29140 -81 -29134 -71
rect -29100 -81 -29046 -71
rect -29012 -81 -28958 -71
rect -28924 -81 -28870 -71
rect -28836 -81 -28830 -47
rect -29140 -83 -28830 -81
rect -29140 -135 -29135 -83
rect -29083 -135 -29053 -83
rect -29001 -135 -28971 -83
rect -28919 -135 -28889 -83
rect -28837 -120 -28830 -83
rect -29140 -147 -29134 -135
rect -29100 -147 -29046 -135
rect -29012 -147 -28958 -135
rect -28924 -147 -28870 -135
rect -29140 -199 -29135 -147
rect -29083 -199 -29053 -147
rect -29001 -199 -28971 -147
rect -28919 -199 -28889 -147
rect -28836 -154 -28830 -120
rect -28837 -193 -28830 -154
rect -29140 -211 -29134 -199
rect -29100 -211 -29046 -199
rect -29012 -211 -28958 -199
rect -28924 -211 -28870 -199
rect -29140 -263 -29135 -211
rect -29083 -263 -29053 -211
rect -29001 -263 -28971 -211
rect -28919 -263 -28889 -211
rect -28836 -227 -28830 -193
rect -28837 -263 -28830 -227
rect -29140 -266 -28830 -263
rect -29140 -275 -29134 -266
rect -29100 -275 -29046 -266
rect -29012 -275 -28958 -266
rect -28924 -275 -28870 -266
rect -29140 -327 -29135 -275
rect -29083 -327 -29053 -275
rect -29001 -327 -28971 -275
rect -28919 -327 -28889 -275
rect -28836 -300 -28830 -266
rect -28837 -327 -28830 -300
rect -29140 -339 -28830 -327
rect -29140 -391 -29135 -339
rect -29083 -391 -29053 -339
rect -29001 -391 -28971 -339
rect -28919 -391 -28889 -339
rect -28836 -373 -28830 -339
rect -28837 -391 -28830 -373
rect -29140 -412 -28830 -391
rect -29140 -446 -29134 -412
rect -29100 -446 -29046 -412
rect -29012 -446 -28958 -412
rect -28924 -446 -28870 -412
rect -28836 -446 -28830 -412
rect -29140 -485 -28830 -446
rect -29140 -519 -29134 -485
rect -29100 -519 -29046 -485
rect -29012 -519 -28958 -485
rect -28924 -519 -28870 -485
rect -28836 -519 -28830 -485
rect -29140 -558 -28830 -519
rect -29140 -592 -29134 -558
rect -29100 -592 -29046 -558
rect -29012 -592 -28958 -558
rect -28924 -592 -28870 -558
rect -28836 -592 -28830 -558
rect -29140 -631 -28830 -592
rect -29140 -665 -29134 -631
rect -29100 -665 -29046 -631
rect -29012 -665 -28958 -631
rect -28924 -665 -28870 -631
rect -28836 -665 -28830 -631
rect -29140 -704 -28830 -665
rect -29140 -738 -29134 -704
rect -29100 -738 -29046 -704
rect -29012 -738 -28958 -704
rect -28924 -738 -28870 -704
rect -28836 -738 -28830 -704
rect -29140 -777 -28830 -738
rect -29140 -811 -29134 -777
rect -29100 -811 -29046 -777
rect -29012 -811 -28958 -777
rect -28924 -811 -28870 -777
rect -28836 -811 -28830 -777
rect -29140 -849 -28830 -811
rect -29140 -883 -29134 -849
rect -29100 -883 -29046 -849
rect -29012 -883 -28958 -849
rect -28924 -883 -28870 -849
rect -28836 -883 -28830 -849
rect -29140 -921 -28830 -883
rect -29140 -955 -29134 -921
rect -29100 -955 -29046 -921
rect -29012 -955 -28958 -921
rect -28924 -955 -28870 -921
rect -28836 -955 -28830 -921
rect -29140 -993 -28830 -955
rect -29140 -1027 -29134 -993
rect -29100 -1027 -29046 -993
rect -29012 -1027 -28958 -993
rect -28924 -1027 -28870 -993
rect -28836 -1027 -28830 -993
rect -29140 -1065 -28830 -1027
rect -29140 -1099 -29134 -1065
rect -29100 -1099 -29046 -1065
rect -29012 -1099 -28958 -1065
rect -28924 -1099 -28870 -1065
rect -28836 -1099 -28830 -1065
rect -29140 -1137 -28830 -1099
rect -29140 -1171 -29134 -1137
rect -29100 -1171 -29046 -1137
rect -29012 -1171 -28958 -1137
rect -28924 -1171 -28870 -1137
rect -28836 -1171 -28830 -1137
rect -29140 -1209 -28830 -1171
rect -29140 -1243 -29134 -1209
rect -29100 -1243 -29046 -1209
rect -29012 -1243 -28958 -1209
rect -28924 -1243 -28870 -1209
rect -28836 -1243 -28830 -1209
rect -29140 -1281 -28830 -1243
rect -29140 -1315 -29134 -1281
rect -29100 -1315 -29046 -1281
rect -29012 -1315 -28958 -1281
rect -28924 -1315 -28870 -1281
rect -28836 -1315 -28830 -1281
rect -29140 -1353 -28830 -1315
rect -29140 -1387 -29134 -1353
rect -29100 -1387 -29046 -1353
rect -29012 -1387 -28958 -1353
rect -28924 -1387 -28870 -1353
rect -28836 -1387 -28830 -1353
rect -29140 -1425 -28830 -1387
rect -29140 -1459 -29134 -1425
rect -29100 -1459 -29046 -1425
rect -29012 -1459 -28958 -1425
rect -28924 -1459 -28870 -1425
rect -28836 -1459 -28830 -1425
rect -29140 -1497 -28830 -1459
rect -29140 -1531 -29134 -1497
rect -29100 -1531 -29046 -1497
rect -29012 -1531 -28958 -1497
rect -28924 -1531 -28870 -1497
rect -28836 -1531 -28830 -1497
rect -29140 -1569 -28830 -1531
rect -29140 -1603 -29134 -1569
rect -29100 -1603 -29046 -1569
rect -29012 -1603 -28958 -1569
rect -28924 -1603 -28870 -1569
rect -28836 -1603 -28830 -1569
rect -29140 -1641 -28830 -1603
rect -29140 -1675 -29134 -1641
rect -29100 -1675 -29046 -1641
rect -29012 -1675 -28958 -1641
rect -28924 -1675 -28870 -1641
rect -28836 -1675 -28830 -1641
rect -29140 -1713 -28830 -1675
rect -29140 -1747 -29134 -1713
rect -29100 -1747 -29046 -1713
rect -29012 -1747 -28958 -1713
rect -28924 -1747 -28870 -1713
rect -28836 -1747 -28830 -1713
rect -29140 -1785 -28830 -1747
rect -29140 -1819 -29134 -1785
rect -29100 -1819 -29046 -1785
rect -29012 -1819 -28958 -1785
rect -28924 -1819 -28870 -1785
rect -28836 -1819 -28830 -1785
rect -29140 -1857 -28830 -1819
rect -29140 -1891 -29134 -1857
rect -29100 -1891 -29046 -1857
rect -29012 -1891 -28958 -1857
rect -28924 -1891 -28870 -1857
rect -28836 -1891 -28830 -1857
rect -29140 -1929 -28830 -1891
rect -29140 -1963 -29134 -1929
rect -29100 -1963 -29046 -1929
rect -29012 -1963 -28958 -1929
rect -28924 -1963 -28870 -1929
rect -28836 -1963 -28830 -1929
rect -29140 -2001 -28830 -1963
rect -29140 -2035 -29134 -2001
rect -29100 -2035 -29046 -2001
rect -29012 -2035 -28958 -2001
rect -28924 -2035 -28870 -2001
rect -28836 -2035 -28830 -2001
rect -29140 -2073 -28830 -2035
rect -29140 -2107 -29134 -2073
rect -29100 -2107 -29046 -2073
rect -29012 -2107 -28958 -2073
rect -28924 -2107 -28870 -2073
rect -28836 -2107 -28830 -2073
rect -29140 -2145 -28830 -2107
rect -29140 -2179 -29134 -2145
rect -29100 -2179 -29046 -2145
rect -29012 -2179 -28958 -2145
rect -28924 -2179 -28870 -2145
rect -28836 -2179 -28830 -2145
rect -29140 -2217 -28830 -2179
rect -29140 -2251 -29134 -2217
rect -29100 -2251 -29046 -2217
rect -29012 -2251 -28958 -2217
rect -28924 -2251 -28870 -2217
rect -28836 -2251 -28830 -2217
rect -29140 -2289 -28830 -2251
rect -29140 -2323 -29134 -2289
rect -29100 -2323 -29046 -2289
rect -29012 -2323 -28958 -2289
rect -28924 -2323 -28870 -2289
rect -28836 -2323 -28830 -2289
rect -29140 -2361 -28830 -2323
rect -29140 -2395 -29134 -2361
rect -29100 -2395 -29046 -2361
rect -29012 -2395 -28958 -2361
rect -28924 -2395 -28870 -2361
rect -28836 -2395 -28830 -2361
rect -29140 -2433 -28830 -2395
rect -29140 -2467 -29134 -2433
rect -29100 -2467 -29046 -2433
rect -29012 -2467 -28958 -2433
rect -28924 -2467 -28870 -2433
rect -28836 -2467 -28830 -2433
rect -29140 -2505 -28830 -2467
rect -29140 -2539 -29134 -2505
rect -29100 -2539 -29046 -2505
rect -29012 -2539 -28958 -2505
rect -28924 -2539 -28870 -2505
rect -28836 -2539 -28830 -2505
rect -29140 -2577 -28830 -2539
rect -29140 -2611 -29134 -2577
rect -29100 -2611 -29046 -2577
rect -29012 -2611 -28958 -2577
rect -28924 -2611 -28870 -2577
rect -28836 -2611 -28830 -2577
rect -29140 -2649 -28830 -2611
rect -29140 -2683 -29134 -2649
rect -29100 -2683 -29046 -2649
rect -29012 -2683 -28958 -2649
rect -28924 -2683 -28870 -2649
rect -28836 -2683 -28830 -2649
rect -29140 -2721 -28830 -2683
rect -29140 -2755 -29134 -2721
rect -29100 -2755 -29046 -2721
rect -29012 -2755 -28958 -2721
rect -28924 -2755 -28870 -2721
rect -28836 -2755 -28830 -2721
rect -29140 -2793 -28830 -2755
rect -29140 -2827 -29134 -2793
rect -29100 -2827 -29046 -2793
rect -29012 -2827 -28958 -2793
rect -28924 -2827 -28870 -2793
rect -28836 -2827 -28830 -2793
rect -29140 -2865 -28830 -2827
rect -29140 -2899 -29134 -2865
rect -29100 -2899 -29046 -2865
rect -29012 -2899 -28958 -2865
rect -28924 -2899 -28870 -2865
rect -28836 -2899 -28830 -2865
rect -29140 -2937 -28830 -2899
rect -29140 -2971 -29134 -2937
rect -29100 -2971 -29046 -2937
rect -29012 -2971 -28958 -2937
rect -28924 -2971 -28870 -2937
rect -28836 -2971 -28830 -2937
rect -29140 -3009 -28830 -2971
rect -29140 -3043 -29134 -3009
rect -29100 -3043 -29046 -3009
rect -29012 -3043 -28958 -3009
rect -28924 -3043 -28870 -3009
rect -28836 -3043 -28830 -3009
rect -29140 -3081 -28830 -3043
rect -29140 -3115 -29134 -3081
rect -29100 -3115 -29046 -3081
rect -29012 -3115 -28958 -3081
rect -28924 -3115 -28870 -3081
rect -28836 -3115 -28830 -3081
rect -29140 -3153 -28830 -3115
rect -29140 -3187 -29134 -3153
rect -29100 -3187 -29046 -3153
rect -29012 -3187 -28958 -3153
rect -28924 -3187 -28870 -3153
rect -28836 -3187 -28830 -3153
rect -29140 -3225 -28830 -3187
rect -29140 -3259 -29134 -3225
rect -29100 -3259 -29046 -3225
rect -29012 -3259 -28958 -3225
rect -28924 -3259 -28870 -3225
rect -28836 -3259 -28830 -3225
rect -29140 -3297 -28830 -3259
rect -29140 -3331 -29134 -3297
rect -29100 -3331 -29046 -3297
rect -29012 -3331 -28958 -3297
rect -28924 -3331 -28870 -3297
rect -28836 -3331 -28830 -3297
rect -29140 -3369 -28830 -3331
rect -29140 -3403 -29134 -3369
rect -29100 -3403 -29046 -3369
rect -29012 -3403 -28958 -3369
rect -28924 -3403 -28870 -3369
rect -28836 -3403 -28830 -3369
rect -29140 -3441 -28830 -3403
rect -29140 -3475 -29134 -3441
rect -29100 -3475 -29046 -3441
rect -29012 -3475 -28958 -3441
rect -28924 -3475 -28870 -3441
rect -28836 -3475 -28830 -3441
rect -29140 -3513 -28830 -3475
rect -29140 -3547 -29134 -3513
rect -29100 -3547 -29046 -3513
rect -29012 -3547 -28958 -3513
rect -28924 -3547 -28870 -3513
rect -28836 -3547 -28830 -3513
rect -29140 -3585 -28830 -3547
rect -29140 -3619 -29134 -3585
rect -29100 -3619 -29046 -3585
rect -29012 -3619 -28958 -3585
rect -28924 -3619 -28870 -3585
rect -28836 -3619 -28830 -3585
rect -29140 -3657 -28830 -3619
rect -29140 -3691 -29134 -3657
rect -29100 -3691 -29046 -3657
rect -29012 -3691 -28958 -3657
rect -28924 -3691 -28870 -3657
rect -28836 -3691 -28830 -3657
rect -29140 -3729 -28830 -3691
rect -29140 -3763 -29134 -3729
rect -29100 -3763 -29046 -3729
rect -29012 -3763 -28958 -3729
rect -28924 -3763 -28870 -3729
rect -28836 -3763 -28830 -3729
rect -29140 -3801 -28830 -3763
rect -29140 -3835 -29134 -3801
rect -29100 -3835 -29046 -3801
rect -29012 -3835 -28958 -3801
rect -28924 -3835 -28870 -3801
rect -28836 -3835 -28830 -3801
rect -29140 -3873 -28830 -3835
rect -29140 -3907 -29134 -3873
rect -29100 -3907 -29046 -3873
rect -29012 -3907 -28958 -3873
rect -28924 -3907 -28870 -3873
rect -28836 -3907 -28830 -3873
rect -29140 -3945 -28830 -3907
rect -29140 -3979 -29134 -3945
rect -29100 -3979 -29046 -3945
rect -29012 -3979 -28958 -3945
rect -28924 -3979 -28870 -3945
rect -28836 -3979 -28830 -3945
rect -29140 -4017 -28830 -3979
rect -29140 -4051 -29134 -4017
rect -29100 -4051 -29046 -4017
rect -29012 -4051 -28958 -4017
rect -28924 -4051 -28870 -4017
rect -28836 -4051 -28830 -4017
rect -29140 -4089 -28830 -4051
rect -29140 -4123 -29134 -4089
rect -29100 -4123 -29046 -4089
rect -29012 -4123 -28958 -4089
rect -28924 -4123 -28870 -4089
rect -28836 -4123 -28830 -4089
rect -29140 -4161 -28830 -4123
rect -29140 -4195 -29134 -4161
rect -29100 -4195 -29046 -4161
rect -29012 -4195 -28958 -4161
rect -28924 -4195 -28870 -4161
rect -28836 -4195 -28830 -4161
rect -29140 -4233 -28830 -4195
rect -29140 -4267 -29134 -4233
rect -29100 -4267 -29046 -4233
rect -29012 -4267 -28958 -4233
rect -28924 -4267 -28870 -4233
rect -28836 -4267 -28830 -4233
rect -29140 -4305 -28830 -4267
rect -29140 -4339 -29134 -4305
rect -29100 -4339 -29046 -4305
rect -29012 -4339 -28958 -4305
rect -28924 -4339 -28870 -4305
rect -28836 -4339 -28830 -4305
rect -29140 -4377 -28830 -4339
rect -29140 -4411 -29134 -4377
rect -29100 -4411 -29046 -4377
rect -29012 -4411 -28958 -4377
rect -28924 -4411 -28870 -4377
rect -28836 -4411 -28830 -4377
rect -29140 -4449 -28830 -4411
rect -29140 -4483 -29134 -4449
rect -29100 -4483 -29046 -4449
rect -29012 -4483 -28958 -4449
rect -28924 -4483 -28870 -4449
rect -28836 -4483 -28830 -4449
rect -29140 -4521 -28830 -4483
rect -29140 -4555 -29134 -4521
rect -29100 -4555 -29046 -4521
rect -29012 -4555 -28958 -4521
rect -28924 -4555 -28870 -4521
rect -28836 -4555 -28830 -4521
rect -29140 -4593 -28830 -4555
rect -29140 -4627 -29134 -4593
rect -29100 -4627 -29046 -4593
rect -29012 -4627 -28958 -4593
rect -28924 -4627 -28870 -4593
rect -28836 -4627 -28830 -4593
rect -29140 -4665 -28830 -4627
rect -29140 -4699 -29134 -4665
rect -29100 -4699 -29046 -4665
rect -29012 -4699 -28958 -4665
rect -28924 -4699 -28870 -4665
rect -28836 -4699 -28830 -4665
rect -29140 -4737 -28830 -4699
rect -29140 -4771 -29134 -4737
rect -29100 -4771 -29046 -4737
rect -29012 -4771 -28958 -4737
rect -28924 -4771 -28870 -4737
rect -28836 -4771 -28830 -4737
rect -29140 -4809 -28830 -4771
rect -29140 -4843 -29134 -4809
rect -29100 -4843 -29046 -4809
rect -29012 -4843 -28958 -4809
rect -28924 -4843 -28870 -4809
rect -28836 -4843 -28830 -4809
rect -29140 -4881 -28830 -4843
rect -29140 -4915 -29134 -4881
rect -29100 -4915 -29046 -4881
rect -29012 -4915 -28958 -4881
rect -28924 -4915 -28870 -4881
rect -28836 -4915 -28830 -4881
rect -29140 -4953 -28830 -4915
rect -29140 -4987 -29134 -4953
rect -29100 -4987 -29046 -4953
rect -29012 -4987 -28958 -4953
rect -28924 -4987 -28870 -4953
rect -28836 -4987 -28830 -4953
rect -29140 -5025 -28830 -4987
rect -29140 -5059 -29134 -5025
rect -29100 -5059 -29046 -5025
rect -29012 -5059 -28958 -5025
rect -28924 -5059 -28870 -5025
rect -28836 -5059 -28830 -5025
rect -29140 -5097 -28830 -5059
rect -29140 -5131 -29134 -5097
rect -29100 -5131 -29046 -5097
rect -29012 -5131 -28958 -5097
rect -28924 -5131 -28870 -5097
rect -28836 -5131 -28830 -5097
rect -29140 -5169 -28830 -5131
rect -29140 -5203 -29134 -5169
rect -29100 -5203 -29046 -5169
rect -29012 -5203 -28958 -5169
rect -28924 -5203 -28870 -5169
rect -28836 -5203 -28830 -5169
rect -29140 -5241 -28830 -5203
rect -29140 -5275 -29134 -5241
rect -29100 -5275 -29046 -5241
rect -29012 -5275 -28958 -5241
rect -28924 -5275 -28870 -5241
rect -28836 -5275 -28830 -5241
rect -29140 -5313 -28830 -5275
rect -29140 -5347 -29134 -5313
rect -29100 -5347 -29046 -5313
rect -29012 -5347 -28958 -5313
rect -28924 -5347 -28870 -5313
rect -28836 -5347 -28830 -5313
rect -29140 -5385 -28830 -5347
rect -29140 -5419 -29134 -5385
rect -29100 -5419 -29046 -5385
rect -29012 -5419 -28958 -5385
rect -28924 -5419 -28870 -5385
rect -28836 -5419 -28830 -5385
rect -29140 -5457 -28830 -5419
rect -29140 -5491 -29134 -5457
rect -29100 -5491 -29046 -5457
rect -29012 -5491 -28958 -5457
rect -28924 -5491 -28870 -5457
rect -28836 -5491 -28830 -5457
rect -29140 -5529 -28830 -5491
rect -29140 -5563 -29134 -5529
rect -29100 -5563 -29046 -5529
rect -29012 -5563 -28958 -5529
rect -28924 -5563 -28870 -5529
rect -28836 -5563 -28830 -5529
rect -29140 -5601 -28830 -5563
rect -29140 -5635 -29134 -5601
rect -29100 -5635 -29046 -5601
rect -29012 -5635 -28958 -5601
rect -28924 -5635 -28870 -5601
rect -28836 -5635 -28830 -5601
rect -29140 -5673 -28830 -5635
rect -29140 -5707 -29134 -5673
rect -29100 -5707 -29046 -5673
rect -29012 -5707 -28958 -5673
rect -28924 -5707 -28870 -5673
rect -28836 -5707 -28830 -5673
rect -29140 -5745 -28830 -5707
rect -29140 -5779 -29134 -5745
rect -29100 -5779 -29046 -5745
rect -29012 -5779 -28958 -5745
rect -28924 -5779 -28870 -5745
rect -28836 -5779 -28830 -5745
rect -29140 -5817 -28830 -5779
rect -29140 -5851 -29134 -5817
rect -29100 -5851 -29046 -5817
rect -29012 -5851 -28958 -5817
rect -28924 -5851 -28870 -5817
rect -28836 -5851 -28830 -5817
rect -29140 -5889 -28830 -5851
rect -29140 -5923 -29134 -5889
rect -29100 -5923 -29046 -5889
rect -29012 -5923 -28958 -5889
rect -28924 -5923 -28870 -5889
rect -28836 -5923 -28830 -5889
rect -29140 -5961 -28830 -5923
rect -29140 -5995 -29134 -5961
rect -29100 -5995 -29046 -5961
rect -29012 -5995 -28958 -5961
rect -28924 -5995 -28870 -5961
rect -28836 -5995 -28830 -5961
rect -29140 -6033 -28830 -5995
rect -29140 -6067 -29134 -6033
rect -29100 -6067 -29046 -6033
rect -29012 -6067 -28958 -6033
rect -28924 -6067 -28870 -6033
rect -28836 -6067 -28830 -6033
rect -29140 -6105 -28830 -6067
rect -29140 -6139 -29134 -6105
rect -29100 -6139 -29046 -6105
rect -29012 -6139 -28958 -6105
rect -28924 -6139 -28870 -6105
rect -28836 -6139 -28830 -6105
rect -29140 -6177 -28830 -6139
rect -29140 -6211 -29134 -6177
rect -29100 -6211 -29046 -6177
rect -29012 -6211 -28958 -6177
rect -28924 -6211 -28870 -6177
rect -28836 -6211 -28830 -6177
rect -29140 -6249 -28830 -6211
rect -29140 -6283 -29134 -6249
rect -29100 -6283 -29046 -6249
rect -29012 -6283 -28958 -6249
rect -28924 -6283 -28870 -6249
rect -28836 -6283 -28830 -6249
rect -29140 -6321 -28830 -6283
rect -29140 -6355 -29134 -6321
rect -29100 -6355 -29046 -6321
rect -29012 -6355 -28958 -6321
rect -28924 -6355 -28870 -6321
rect -28836 -6355 -28830 -6321
rect -29140 -6393 -28830 -6355
rect -29140 -6427 -29134 -6393
rect -29100 -6427 -29046 -6393
rect -29012 -6427 -28958 -6393
rect -28924 -6427 -28870 -6393
rect -28836 -6427 -28830 -6393
rect -29140 -6465 -28830 -6427
rect -29140 -6499 -29134 -6465
rect -29100 -6499 -29046 -6465
rect -29012 -6499 -28958 -6465
rect -28924 -6499 -28870 -6465
rect -28836 -6499 -28830 -6465
rect -29140 -6537 -28830 -6499
rect -29140 -6571 -29134 -6537
rect -29100 -6571 -29046 -6537
rect -29012 -6571 -28958 -6537
rect -28924 -6571 -28870 -6537
rect -28836 -6571 -28830 -6537
rect -29140 -6609 -28830 -6571
rect -29140 -6643 -29134 -6609
rect -29100 -6643 -29046 -6609
rect -29012 -6643 -28958 -6609
rect -28924 -6643 -28870 -6609
rect -28836 -6643 -28830 -6609
rect -29140 -6681 -28830 -6643
rect -29140 -6715 -29134 -6681
rect -29100 -6715 -29046 -6681
rect -29012 -6715 -28958 -6681
rect -28924 -6715 -28870 -6681
rect -28836 -6715 -28830 -6681
rect -29140 -6753 -28830 -6715
rect -29140 -6787 -29134 -6753
rect -29100 -6787 -29046 -6753
rect -29012 -6787 -28958 -6753
rect -28924 -6787 -28870 -6753
rect -28836 -6787 -28830 -6753
rect -29140 -6825 -28830 -6787
rect -29140 -6859 -29134 -6825
rect -29100 -6859 -29046 -6825
rect -29012 -6859 -28958 -6825
rect -28924 -6859 -28870 -6825
rect -28836 -6859 -28830 -6825
rect -29140 -6897 -28830 -6859
rect -29140 -6931 -29134 -6897
rect -29100 -6931 -29046 -6897
rect -29012 -6931 -28958 -6897
rect -28924 -6931 -28870 -6897
rect -28836 -6931 -28830 -6897
rect -29140 -6969 -28830 -6931
rect -29140 -7003 -29134 -6969
rect -29100 -7003 -29046 -6969
rect -29012 -7003 -28958 -6969
rect -28924 -7003 -28870 -6969
rect -28836 -7003 -28830 -6969
rect -29140 -7041 -28830 -7003
rect -29140 -7075 -29134 -7041
rect -29100 -7075 -29046 -7041
rect -29012 -7075 -28958 -7041
rect -28924 -7075 -28870 -7041
rect -28836 -7075 -28830 -7041
rect -29140 -7113 -28830 -7075
rect -29140 -7147 -29134 -7113
rect -29100 -7147 -29046 -7113
rect -29012 -7147 -28958 -7113
rect -28924 -7147 -28870 -7113
rect -28836 -7147 -28830 -7113
rect -29140 -7185 -28830 -7147
rect -29140 -7219 -29134 -7185
rect -29100 -7219 -29046 -7185
rect -29012 -7219 -28958 -7185
rect -28924 -7219 -28870 -7185
rect -28836 -7219 -28830 -7185
rect -29140 -7257 -28830 -7219
rect -29140 -7291 -29134 -7257
rect -29100 -7291 -29046 -7257
rect -29012 -7291 -28958 -7257
rect -28924 -7291 -28870 -7257
rect -28836 -7291 -28830 -7257
rect -29140 -7329 -28830 -7291
rect -29140 -7363 -29134 -7329
rect -29100 -7363 -29046 -7329
rect -29012 -7363 -28958 -7329
rect -28924 -7363 -28870 -7329
rect -28836 -7363 -28830 -7329
rect -29140 -7401 -28830 -7363
rect -29140 -7435 -29134 -7401
rect -29100 -7435 -29046 -7401
rect -29012 -7435 -28958 -7401
rect -28924 -7435 -28870 -7401
rect -28836 -7435 -28830 -7401
rect -29140 -7473 -28830 -7435
rect -29140 -7507 -29134 -7473
rect -29100 -7507 -29046 -7473
rect -29012 -7507 -28958 -7473
rect -28924 -7507 -28870 -7473
rect -28836 -7507 -28830 -7473
rect -29140 -7545 -28830 -7507
rect -29140 -7579 -29134 -7545
rect -29100 -7579 -29046 -7545
rect -29012 -7579 -28958 -7545
rect -28924 -7579 -28870 -7545
rect -28836 -7579 -28830 -7545
rect -29140 -7617 -28830 -7579
rect -29140 -7651 -29134 -7617
rect -29100 -7651 -29046 -7617
rect -29012 -7651 -28958 -7617
rect -28924 -7651 -28870 -7617
rect -28836 -7651 -28830 -7617
rect -29140 -7689 -28830 -7651
rect -29140 -7723 -29134 -7689
rect -29100 -7723 -29046 -7689
rect -29012 -7723 -28958 -7689
rect -28924 -7723 -28870 -7689
rect -28836 -7723 -28830 -7689
rect -29140 -7761 -28830 -7723
rect -29140 -7795 -29134 -7761
rect -29100 -7795 -29046 -7761
rect -29012 -7795 -28958 -7761
rect -28924 -7795 -28870 -7761
rect -28836 -7795 -28830 -7761
rect -29140 -7833 -28830 -7795
rect -29140 -7867 -29134 -7833
rect -29100 -7867 -29046 -7833
rect -29012 -7867 -28958 -7833
rect -28924 -7867 -28870 -7833
rect -28836 -7867 -28830 -7833
rect -29140 -7905 -28830 -7867
rect -29140 -7939 -29134 -7905
rect -29100 -7939 -29046 -7905
rect -29012 -7939 -28958 -7905
rect -28924 -7939 -28870 -7905
rect -28836 -7939 -28830 -7905
rect -29140 -7977 -28830 -7939
rect -29140 -8011 -29134 -7977
rect -29100 -8011 -29046 -7977
rect -29012 -8011 -28958 -7977
rect -28924 -8011 -28870 -7977
rect -28836 -8011 -28830 -7977
rect -29140 -8049 -28830 -8011
rect -29140 -8083 -29134 -8049
rect -29100 -8083 -29046 -8049
rect -29012 -8083 -28958 -8049
rect -28924 -8083 -28870 -8049
rect -28836 -8083 -28830 -8049
rect -29140 -8121 -28830 -8083
rect -29140 -8155 -29134 -8121
rect -29100 -8155 -29046 -8121
rect -29012 -8155 -28958 -8121
rect -28924 -8155 -28870 -8121
rect -28836 -8155 -28830 -8121
rect -29140 -8193 -28830 -8155
rect -29140 -8227 -29134 -8193
rect -29100 -8227 -29046 -8193
rect -29012 -8227 -28958 -8193
rect -28924 -8227 -28870 -8193
rect -28836 -8227 -28830 -8193
rect -29140 -8265 -28830 -8227
rect -29140 -8299 -29134 -8265
rect -29100 -8299 -29046 -8265
rect -29012 -8299 -28958 -8265
rect -28924 -8299 -28870 -8265
rect -28836 -8299 -28830 -8265
rect -29140 -8337 -28830 -8299
rect -29140 -8371 -29134 -8337
rect -29100 -8371 -29046 -8337
rect -29012 -8371 -28958 -8337
rect -28924 -8371 -28870 -8337
rect -28836 -8371 -28830 -8337
rect -29140 -8409 -28830 -8371
rect -29140 -8443 -29134 -8409
rect -29100 -8443 -29046 -8409
rect -29012 -8443 -28958 -8409
rect -28924 -8443 -28870 -8409
rect -28836 -8443 -28830 -8409
rect -29140 -8481 -28830 -8443
rect -29140 -8515 -29134 -8481
rect -29100 -8515 -29046 -8481
rect -29012 -8515 -28958 -8481
rect -28924 -8515 -28870 -8481
rect -28836 -8515 -28830 -8481
rect -29140 -8553 -28830 -8515
rect -32350 -8640 -32344 -8606
rect -32310 -8640 -32266 -8606
rect -32232 -8640 -32188 -8606
rect -32154 -8640 -32110 -8606
rect -32076 -8640 -32032 -8606
rect -31998 -8640 -31954 -8606
rect -31920 -8640 -31876 -8606
rect -31842 -8640 -31798 -8606
rect -31764 -8640 -31758 -8606
rect -29280 -8589 -29228 -8579
rect -32350 -8678 -31758 -8640
rect -32350 -8712 -32344 -8678
rect -32310 -8712 -32266 -8678
rect -32232 -8712 -32188 -8678
rect -32154 -8712 -32110 -8678
rect -32076 -8712 -32032 -8678
rect -31998 -8712 -31954 -8678
rect -31920 -8712 -31876 -8678
rect -31842 -8712 -31798 -8678
rect -31764 -8697 -31758 -8678
rect -31521 -8625 -31469 -8611
rect -31521 -8689 -31469 -8677
tri -31758 -8697 -31750 -8689 sw
rect -31764 -8712 -31750 -8697
rect -32350 -8731 -31750 -8712
tri -31750 -8731 -31716 -8697 sw
rect -29280 -8653 -29228 -8641
rect -29280 -8711 -29228 -8705
rect -29140 -8587 -29134 -8553
rect -29100 -8587 -29046 -8553
rect -29012 -8587 -28958 -8553
rect -28924 -8587 -28870 -8553
rect -28836 -8587 -28830 -8553
rect -29140 -8625 -28830 -8587
rect -29140 -8659 -29134 -8625
rect -29100 -8659 -29046 -8625
rect -29012 -8659 -28958 -8625
rect -28924 -8659 -28870 -8625
rect -28836 -8659 -28830 -8625
rect -29140 -8697 -28830 -8659
tri -29153 -8731 -29140 -8718 se
rect -29140 -8731 -29134 -8697
rect -29100 -8731 -29046 -8697
rect -29012 -8731 -28958 -8697
rect -28924 -8731 -28870 -8697
rect -28836 -8731 -28830 -8697
rect -32350 -8750 -31716 -8731
rect -32350 -8784 -32344 -8750
rect -32310 -8784 -32266 -8750
rect -32232 -8784 -32188 -8750
rect -32154 -8784 -32110 -8750
rect -32076 -8784 -32032 -8750
rect -31998 -8784 -31954 -8750
rect -31920 -8784 -31876 -8750
rect -31842 -8784 -31798 -8750
rect -31764 -8764 -31716 -8750
tri -31716 -8764 -31683 -8731 sw
rect -31521 -8747 -31469 -8741
tri -29169 -8747 -29153 -8731 se
rect -29153 -8747 -28830 -8731
tri -29186 -8764 -29169 -8747 se
rect -29169 -8764 -28830 -8747
rect -31764 -8769 -31683 -8764
tri -31683 -8769 -31678 -8764 sw
tri -29191 -8769 -29186 -8764 se
rect -29186 -8769 -28830 -8764
rect -31764 -8784 -31678 -8769
rect -32350 -8803 -31678 -8784
tri -31678 -8803 -31644 -8769 sw
tri -29225 -8803 -29191 -8769 se
rect -29191 -8803 -29134 -8769
rect -29100 -8803 -29046 -8769
rect -29012 -8803 -28958 -8769
rect -28924 -8803 -28870 -8769
rect -28836 -8803 -28830 -8769
rect -32350 -8822 -31644 -8803
rect -32350 -8856 -32344 -8822
rect -32310 -8856 -32266 -8822
rect -32232 -8856 -32188 -8822
rect -32154 -8856 -32110 -8822
rect -32076 -8856 -32032 -8822
rect -31998 -8856 -31954 -8822
rect -31920 -8856 -31876 -8822
rect -31842 -8856 -31798 -8822
rect -31764 -8836 -31644 -8822
tri -31644 -8836 -31611 -8803 sw
tri -29258 -8836 -29225 -8803 se
rect -29225 -8836 -28830 -8803
rect -31764 -8841 -31611 -8836
tri -31611 -8841 -31606 -8836 sw
tri -29263 -8841 -29258 -8836 se
rect -29258 -8841 -28830 -8836
rect -31764 -8856 -31606 -8841
rect -32350 -8875 -31606 -8856
tri -31606 -8875 -31572 -8841 sw
tri -29297 -8875 -29263 -8841 se
rect -29263 -8875 -29134 -8841
rect -29100 -8875 -29046 -8841
rect -29012 -8875 -28958 -8841
rect -28924 -8875 -28870 -8841
rect -28836 -8875 -28830 -8841
rect -32350 -8908 -31572 -8875
tri -31572 -8908 -31539 -8875 sw
tri -29330 -8908 -29297 -8875 se
rect -29297 -8908 -28830 -8875
rect -32350 -8911 -31539 -8908
tri -31539 -8911 -31536 -8908 sw
tri -29333 -8911 -29330 -8908 se
rect -29330 -8911 -28830 -8908
rect -32350 -8913 -28830 -8911
rect -32350 -8918 -29134 -8913
rect -32350 -9600 -32338 -8918
rect -30792 -8952 -30753 -8918
rect -30719 -8952 -30680 -8918
rect -30646 -8952 -30607 -8918
rect -30573 -8952 -30534 -8918
rect -30500 -8952 -30461 -8918
rect -30427 -8952 -30388 -8918
rect -30354 -8952 -30315 -8918
rect -30281 -8952 -30242 -8918
rect -30208 -8952 -30169 -8918
rect -30135 -8952 -30096 -8918
rect -30062 -8952 -30023 -8918
rect -29989 -8952 -29950 -8918
rect -29916 -8952 -29877 -8918
rect -29843 -8952 -29804 -8918
rect -29770 -8952 -29731 -8918
rect -29697 -8952 -29658 -8918
rect -29624 -8952 -29585 -8918
rect -29551 -8952 -29512 -8918
rect -29478 -8952 -29439 -8918
rect -29405 -8952 -29366 -8918
rect -29332 -8952 -29293 -8918
rect -29259 -8952 -29220 -8918
rect -29186 -8947 -29134 -8918
rect -29100 -8947 -29046 -8913
rect -29012 -8947 -28958 -8913
rect -28924 -8947 -28870 -8913
rect -28836 -8947 -28830 -8913
rect -29186 -8952 -28830 -8947
rect -30792 -8985 -28830 -8952
rect -30792 -8990 -29134 -8985
rect -30792 -9024 -30753 -8990
rect -30719 -9024 -30680 -8990
rect -30646 -9024 -30607 -8990
rect -30573 -9024 -30534 -8990
rect -30500 -9024 -30461 -8990
rect -30427 -9024 -30388 -8990
rect -30354 -9024 -30315 -8990
rect -30281 -9024 -30242 -8990
rect -30208 -9024 -30169 -8990
rect -30135 -9024 -30096 -8990
rect -30062 -9024 -30023 -8990
rect -29989 -9024 -29950 -8990
rect -29916 -9024 -29877 -8990
rect -29843 -9024 -29804 -8990
rect -29770 -9024 -29731 -8990
rect -29697 -9024 -29658 -8990
rect -29624 -9024 -29585 -8990
rect -29551 -9024 -29512 -8990
rect -29478 -9024 -29439 -8990
rect -29405 -9024 -29366 -8990
rect -29332 -9024 -29293 -8990
rect -29259 -9024 -29220 -8990
rect -29186 -9019 -29134 -8990
rect -29100 -9019 -29046 -8985
rect -29012 -9019 -28958 -8985
rect -28924 -9019 -28870 -8985
rect -28836 -9019 -28830 -8985
rect -29186 -9024 -28830 -9019
rect -30792 -9057 -28830 -9024
rect -30792 -9062 -29134 -9057
rect -30792 -9096 -30753 -9062
rect -30719 -9096 -30680 -9062
rect -30646 -9096 -30607 -9062
rect -30573 -9096 -30534 -9062
rect -30500 -9096 -30461 -9062
rect -30427 -9096 -30388 -9062
rect -30354 -9096 -30315 -9062
rect -30281 -9096 -30242 -9062
rect -30208 -9096 -30169 -9062
rect -30135 -9096 -30096 -9062
rect -30062 -9096 -30023 -9062
rect -29989 -9096 -29950 -9062
rect -29916 -9096 -29877 -9062
rect -29843 -9096 -29804 -9062
rect -29770 -9096 -29731 -9062
rect -29697 -9096 -29658 -9062
rect -29624 -9096 -29585 -9062
rect -29551 -9096 -29512 -9062
rect -29478 -9096 -29439 -9062
rect -29405 -9096 -29366 -9062
rect -29332 -9096 -29293 -9062
rect -29259 -9096 -29220 -9062
rect -29186 -9091 -29134 -9062
rect -29100 -9091 -29046 -9057
rect -29012 -9091 -28958 -9057
rect -28924 -9091 -28870 -9057
rect -28836 -9091 -28830 -9057
rect -29186 -9096 -28830 -9091
rect -30792 -9129 -28830 -9096
rect -30792 -9134 -29134 -9129
rect -30792 -9168 -30753 -9134
rect -30719 -9168 -30680 -9134
rect -30646 -9168 -30607 -9134
rect -30573 -9168 -30534 -9134
rect -30500 -9168 -30461 -9134
rect -30427 -9168 -30388 -9134
rect -30354 -9168 -30315 -9134
rect -30281 -9168 -30242 -9134
rect -30208 -9168 -30169 -9134
rect -30135 -9168 -30096 -9134
rect -30062 -9168 -30023 -9134
rect -29989 -9168 -29950 -9134
rect -29916 -9168 -29877 -9134
rect -29843 -9168 -29804 -9134
rect -29770 -9168 -29731 -9134
rect -29697 -9168 -29658 -9134
rect -29624 -9168 -29585 -9134
rect -29551 -9168 -29512 -9134
rect -29478 -9168 -29439 -9134
rect -29405 -9168 -29366 -9134
rect -29332 -9168 -29293 -9134
rect -29259 -9168 -29220 -9134
rect -29186 -9163 -29134 -9134
rect -29100 -9163 -29046 -9129
rect -29012 -9163 -28958 -9129
rect -28924 -9163 -28870 -9129
rect -28836 -9163 -28830 -9129
rect -29186 -9168 -28830 -9163
rect -30792 -9201 -28830 -9168
rect -30792 -9206 -29134 -9201
rect -30792 -9240 -30753 -9206
rect -30719 -9240 -30680 -9206
rect -30646 -9240 -30607 -9206
rect -30573 -9240 -30534 -9206
rect -30500 -9240 -30461 -9206
rect -30427 -9240 -30388 -9206
rect -30354 -9240 -30315 -9206
rect -30281 -9240 -30242 -9206
rect -30208 -9240 -30169 -9206
rect -30135 -9240 -30096 -9206
rect -30062 -9240 -30023 -9206
rect -29989 -9240 -29950 -9206
rect -29916 -9240 -29877 -9206
rect -29843 -9240 -29804 -9206
rect -29770 -9240 -29731 -9206
rect -29697 -9240 -29658 -9206
rect -29624 -9240 -29585 -9206
rect -29551 -9240 -29512 -9206
rect -29478 -9240 -29439 -9206
rect -29405 -9240 -29366 -9206
rect -29332 -9240 -29293 -9206
rect -29259 -9240 -29220 -9206
rect -29186 -9235 -29134 -9206
rect -29100 -9235 -29046 -9201
rect -29012 -9235 -28958 -9201
rect -28924 -9235 -28870 -9201
rect -28836 -9235 -28830 -9201
rect -29186 -9240 -28830 -9235
rect -30792 -9273 -28830 -9240
rect -30792 -9278 -29134 -9273
rect -30792 -9312 -30753 -9278
rect -30719 -9312 -30680 -9278
rect -30646 -9312 -30607 -9278
rect -30573 -9312 -30534 -9278
rect -30500 -9312 -30461 -9278
rect -30427 -9312 -30388 -9278
rect -30354 -9312 -30315 -9278
rect -30281 -9312 -30242 -9278
rect -30208 -9312 -30169 -9278
rect -30135 -9312 -30096 -9278
rect -30062 -9312 -30023 -9278
rect -29989 -9312 -29950 -9278
rect -29916 -9312 -29877 -9278
rect -29843 -9312 -29804 -9278
rect -29770 -9312 -29731 -9278
rect -29697 -9312 -29658 -9278
rect -29624 -9312 -29585 -9278
rect -29551 -9312 -29512 -9278
rect -29478 -9312 -29439 -9278
rect -29405 -9312 -29366 -9278
rect -29332 -9312 -29293 -9278
rect -29259 -9312 -29220 -9278
rect -29186 -9307 -29134 -9278
rect -29100 -9307 -29046 -9273
rect -29012 -9307 -28958 -9273
rect -28924 -9307 -28870 -9273
rect -28836 -9307 -28830 -9273
rect -29186 -9312 -28830 -9307
rect -30792 -9345 -28830 -9312
rect -30792 -9350 -29134 -9345
rect -30792 -9384 -30753 -9350
rect -30719 -9384 -30680 -9350
rect -30646 -9384 -30607 -9350
rect -30573 -9384 -30534 -9350
rect -30500 -9384 -30461 -9350
rect -30427 -9384 -30388 -9350
rect -30354 -9384 -30315 -9350
rect -30281 -9384 -30242 -9350
rect -30208 -9384 -30169 -9350
rect -30135 -9384 -30096 -9350
rect -30062 -9384 -30023 -9350
rect -29989 -9384 -29950 -9350
rect -29916 -9384 -29877 -9350
rect -29843 -9384 -29804 -9350
rect -29770 -9384 -29731 -9350
rect -29697 -9384 -29658 -9350
rect -29624 -9384 -29585 -9350
rect -29551 -9384 -29512 -9350
rect -29478 -9384 -29439 -9350
rect -29405 -9384 -29366 -9350
rect -29332 -9384 -29293 -9350
rect -29259 -9384 -29220 -9350
rect -29186 -9379 -29134 -9350
rect -29100 -9379 -29046 -9345
rect -29012 -9379 -28958 -9345
rect -28924 -9379 -28870 -9345
rect -28836 -9379 -28830 -9345
rect -29186 -9384 -28830 -9379
rect -30792 -9417 -28830 -9384
rect -28202 4239 -27106 4721
rect -21227 4644 -21221 4696
rect -21169 4644 -21145 4696
rect -21093 4644 -21069 4696
rect -21017 4644 -20993 4696
rect -20941 4644 -20917 4696
rect -20865 4644 -20841 4696
rect -20789 4644 -20783 4696
rect -21227 4570 -20783 4644
rect -21227 4518 -21221 4570
rect -21169 4518 -21145 4570
rect -21093 4518 -21069 4570
rect -21017 4518 -20993 4570
rect -20941 4518 -20917 4570
rect -20865 4518 -20841 4570
rect -20789 4518 -20783 4570
rect -28202 4205 -28189 4239
rect -28155 4205 -28115 4239
rect -28081 4205 -28041 4239
rect -28007 4205 -27967 4239
rect -27933 4205 -27893 4239
rect -27859 4205 -27819 4239
rect -27785 4205 -27745 4239
rect -27711 4205 -27671 4239
rect -27637 4205 -27597 4239
rect -27563 4205 -27523 4239
rect -27489 4205 -27449 4239
rect -27415 4205 -27375 4239
rect -27341 4205 -27301 4239
rect -27267 4205 -27227 4239
rect -27193 4205 -27153 4239
rect -27119 4205 -27106 4239
rect -28202 4166 -27106 4205
rect -28202 4132 -28189 4166
rect -28155 4132 -28115 4166
rect -28081 4132 -28041 4166
rect -28007 4132 -27967 4166
rect -27933 4132 -27893 4166
rect -27859 4132 -27819 4166
rect -27785 4132 -27745 4166
rect -27711 4132 -27671 4166
rect -27637 4132 -27597 4166
rect -27563 4132 -27523 4166
rect -27489 4132 -27449 4166
rect -27415 4132 -27375 4166
rect -27341 4132 -27301 4166
rect -27267 4132 -27227 4166
rect -27193 4132 -27153 4166
rect -27119 4132 -27106 4166
rect -28202 4093 -27106 4132
rect -28202 4059 -28189 4093
rect -28155 4059 -28115 4093
rect -28081 4059 -28041 4093
rect -28007 4059 -27967 4093
rect -27933 4059 -27893 4093
rect -27859 4059 -27819 4093
rect -27785 4059 -27745 4093
rect -27711 4059 -27671 4093
rect -27637 4059 -27597 4093
rect -27563 4059 -27523 4093
rect -27489 4059 -27449 4093
rect -27415 4059 -27375 4093
rect -27341 4059 -27301 4093
rect -27267 4059 -27227 4093
rect -27193 4059 -27153 4093
rect -27119 4059 -27106 4093
rect -28202 4020 -27106 4059
rect -28202 3986 -28189 4020
rect -28155 3986 -28115 4020
rect -28081 3986 -28041 4020
rect -28007 3986 -27967 4020
rect -27933 3986 -27893 4020
rect -27859 3986 -27819 4020
rect -27785 3986 -27745 4020
rect -27711 3986 -27671 4020
rect -27637 3986 -27597 4020
rect -27563 3986 -27523 4020
rect -27489 3986 -27449 4020
rect -27415 3986 -27375 4020
rect -27341 3986 -27301 4020
rect -27267 3986 -27227 4020
rect -27193 3986 -27153 4020
rect -27119 3986 -27106 4020
rect -28202 3947 -27106 3986
rect -28202 3913 -28189 3947
rect -28155 3913 -28115 3947
rect -28081 3913 -28041 3947
rect -28007 3913 -27967 3947
rect -27933 3913 -27893 3947
rect -27859 3913 -27819 3947
rect -27785 3913 -27745 3947
rect -27711 3913 -27671 3947
rect -27637 3913 -27597 3947
rect -27563 3913 -27523 3947
rect -27489 3913 -27449 3947
rect -27415 3913 -27375 3947
rect -27341 3913 -27301 3947
rect -27267 3913 -27227 3947
rect -27193 3913 -27153 3947
rect -27119 3913 -27106 3947
rect -28202 3874 -27106 3913
rect -28202 3840 -28189 3874
rect -28155 3840 -28115 3874
rect -28081 3840 -28041 3874
rect -28007 3840 -27967 3874
rect -27933 3840 -27893 3874
rect -27859 3840 -27819 3874
rect -27785 3840 -27745 3874
rect -27711 3840 -27671 3874
rect -27637 3840 -27597 3874
rect -27563 3840 -27523 3874
rect -27489 3840 -27449 3874
rect -27415 3840 -27375 3874
rect -27341 3840 -27301 3874
rect -27267 3840 -27227 3874
rect -27193 3840 -27153 3874
rect -27119 3840 -27106 3874
rect -28202 3801 -27106 3840
rect -28202 3767 -28189 3801
rect -28155 3767 -28115 3801
rect -28081 3767 -28041 3801
rect -28007 3767 -27967 3801
rect -27933 3767 -27893 3801
rect -27859 3767 -27819 3801
rect -27785 3767 -27745 3801
rect -27711 3767 -27671 3801
rect -27637 3767 -27597 3801
rect -27563 3767 -27523 3801
rect -27489 3767 -27449 3801
rect -27415 3767 -27375 3801
rect -27341 3767 -27301 3801
rect -27267 3767 -27227 3801
rect -27193 3767 -27153 3801
rect -27119 3767 -27106 3801
rect -28202 3728 -27106 3767
rect -28202 3694 -28189 3728
rect -28155 3694 -28115 3728
rect -28081 3694 -28041 3728
rect -28007 3694 -27967 3728
rect -27933 3694 -27893 3728
rect -27859 3694 -27819 3728
rect -27785 3694 -27745 3728
rect -27711 3694 -27671 3728
rect -27637 3694 -27597 3728
rect -27563 3694 -27523 3728
rect -27489 3694 -27449 3728
rect -27415 3694 -27375 3728
rect -27341 3694 -27301 3728
rect -27267 3694 -27227 3728
rect -27193 3694 -27153 3728
rect -27119 3694 -27106 3728
rect -28202 3655 -27106 3694
rect -28202 3621 -28189 3655
rect -28155 3621 -28115 3655
rect -28081 3621 -28041 3655
rect -28007 3621 -27967 3655
rect -27933 3621 -27893 3655
rect -27859 3621 -27819 3655
rect -27785 3621 -27745 3655
rect -27711 3621 -27671 3655
rect -27637 3621 -27597 3655
rect -27563 3621 -27523 3655
rect -27489 3621 -27449 3655
rect -27415 3621 -27375 3655
rect -27341 3621 -27301 3655
rect -27267 3621 -27227 3655
rect -27193 3621 -27153 3655
rect -27119 3621 -27106 3655
rect -28202 3582 -27106 3621
rect -28202 3548 -28189 3582
rect -28155 3548 -28115 3582
rect -28081 3548 -28041 3582
rect -28007 3548 -27967 3582
rect -27933 3548 -27893 3582
rect -27859 3548 -27819 3582
rect -27785 3548 -27745 3582
rect -27711 3548 -27671 3582
rect -27637 3548 -27597 3582
rect -27563 3548 -27523 3582
rect -27489 3548 -27449 3582
rect -27415 3548 -27375 3582
rect -27341 3548 -27301 3582
rect -27267 3548 -27227 3582
rect -27193 3548 -27153 3582
rect -27119 3548 -27106 3582
rect -28202 3509 -27106 3548
rect -28202 3475 -28189 3509
rect -28155 3475 -28115 3509
rect -28081 3475 -28041 3509
rect -28007 3475 -27967 3509
rect -27933 3475 -27893 3509
rect -27859 3475 -27819 3509
rect -27785 3475 -27745 3509
rect -27711 3475 -27671 3509
rect -27637 3475 -27597 3509
rect -27563 3475 -27523 3509
rect -27489 3475 -27449 3509
rect -27415 3475 -27375 3509
rect -27341 3475 -27301 3509
rect -27267 3475 -27227 3509
rect -27193 3475 -27153 3509
rect -27119 3475 -27106 3509
rect -28202 3436 -27106 3475
rect -28202 3402 -28189 3436
rect -28155 3402 -28115 3436
rect -28081 3402 -28041 3436
rect -28007 3402 -27967 3436
rect -27933 3402 -27893 3436
rect -27859 3402 -27819 3436
rect -27785 3402 -27745 3436
rect -27711 3402 -27671 3436
rect -27637 3402 -27597 3436
rect -27563 3402 -27523 3436
rect -27489 3402 -27449 3436
rect -27415 3402 -27375 3436
rect -27341 3402 -27301 3436
rect -27267 3402 -27227 3436
rect -27193 3402 -27153 3436
rect -27119 3402 -27106 3436
rect -28202 3363 -27106 3402
rect -28202 3329 -28189 3363
rect -28155 3329 -28115 3363
rect -28081 3329 -28041 3363
rect -28007 3329 -27967 3363
rect -27933 3329 -27893 3363
rect -27859 3329 -27819 3363
rect -27785 3329 -27745 3363
rect -27711 3329 -27671 3363
rect -27637 3329 -27597 3363
rect -27563 3329 -27523 3363
rect -27489 3329 -27449 3363
rect -27415 3329 -27375 3363
rect -27341 3329 -27301 3363
rect -27267 3329 -27227 3363
rect -27193 3329 -27153 3363
rect -27119 3329 -27106 3363
rect -28202 3290 -27106 3329
rect -28202 3256 -28189 3290
rect -28155 3256 -28115 3290
rect -28081 3256 -28041 3290
rect -28007 3256 -27967 3290
rect -27933 3256 -27893 3290
rect -27859 3256 -27819 3290
rect -27785 3256 -27745 3290
rect -27711 3256 -27671 3290
rect -27637 3256 -27597 3290
rect -27563 3256 -27523 3290
rect -27489 3256 -27449 3290
rect -27415 3256 -27375 3290
rect -27341 3256 -27301 3290
rect -27267 3256 -27227 3290
rect -27193 3256 -27153 3290
rect -27119 3256 -27106 3290
rect -28202 3217 -27106 3256
rect -28202 3183 -28189 3217
rect -28155 3183 -28115 3217
rect -28081 3183 -28041 3217
rect -28007 3183 -27967 3217
rect -27933 3183 -27893 3217
rect -27859 3183 -27819 3217
rect -27785 3183 -27745 3217
rect -27711 3183 -27671 3217
rect -27637 3183 -27597 3217
rect -27563 3183 -27523 3217
rect -27489 3183 -27449 3217
rect -27415 3183 -27375 3217
rect -27341 3183 -27301 3217
rect -27267 3183 -27227 3217
rect -27193 3183 -27153 3217
rect -27119 3183 -27106 3217
rect -28202 3144 -27106 3183
rect -28202 3110 -28189 3144
rect -28155 3110 -28115 3144
rect -28081 3110 -28041 3144
rect -28007 3110 -27967 3144
rect -27933 3110 -27893 3144
rect -27859 3110 -27819 3144
rect -27785 3110 -27745 3144
rect -27711 3110 -27671 3144
rect -27637 3110 -27597 3144
rect -27563 3110 -27523 3144
rect -27489 3110 -27449 3144
rect -27415 3110 -27375 3144
rect -27341 3110 -27301 3144
rect -27267 3110 -27227 3144
rect -27193 3110 -27153 3144
rect -27119 3110 -27106 3144
rect -28202 3071 -27106 3110
rect -28202 3037 -28189 3071
rect -28155 3037 -28115 3071
rect -28081 3037 -28041 3071
rect -28007 3037 -27967 3071
rect -27933 3037 -27893 3071
rect -27859 3037 -27819 3071
rect -27785 3037 -27745 3071
rect -27711 3037 -27671 3071
rect -27637 3037 -27597 3071
rect -27563 3037 -27523 3071
rect -27489 3037 -27449 3071
rect -27415 3037 -27375 3071
rect -27341 3037 -27301 3071
rect -27267 3037 -27227 3071
rect -27193 3037 -27153 3071
rect -27119 3037 -27106 3071
rect -28202 2998 -27106 3037
rect -28202 2964 -28189 2998
rect -28155 2964 -28115 2998
rect -28081 2964 -28041 2998
rect -28007 2964 -27967 2998
rect -27933 2964 -27893 2998
rect -27859 2964 -27819 2998
rect -27785 2964 -27745 2998
rect -27711 2964 -27671 2998
rect -27637 2964 -27597 2998
rect -27563 2964 -27523 2998
rect -27489 2964 -27449 2998
rect -27415 2964 -27375 2998
rect -27341 2964 -27301 2998
rect -27267 2964 -27227 2998
rect -27193 2964 -27153 2998
rect -27119 2964 -27106 2998
rect -28202 2925 -27106 2964
rect -28202 2891 -28189 2925
rect -28155 2891 -28115 2925
rect -28081 2891 -28041 2925
rect -28007 2891 -27967 2925
rect -27933 2891 -27893 2925
rect -27859 2891 -27819 2925
rect -27785 2891 -27745 2925
rect -27711 2891 -27671 2925
rect -27637 2891 -27597 2925
rect -27563 2891 -27523 2925
rect -27489 2891 -27449 2925
rect -27415 2891 -27375 2925
rect -27341 2891 -27301 2925
rect -27267 2891 -27227 2925
rect -27193 2891 -27153 2925
rect -27119 2891 -27106 2925
rect -28202 2852 -27106 2891
rect -28202 2818 -28189 2852
rect -28155 2818 -28115 2852
rect -28081 2818 -28041 2852
rect -28007 2818 -27967 2852
rect -27933 2818 -27893 2852
rect -27859 2818 -27819 2852
rect -27785 2818 -27745 2852
rect -27711 2818 -27671 2852
rect -27637 2818 -27597 2852
rect -27563 2818 -27523 2852
rect -27489 2818 -27449 2852
rect -27415 2818 -27375 2852
rect -27341 2818 -27301 2852
rect -27267 2818 -27227 2852
rect -27193 2818 -27153 2852
rect -27119 2818 -27106 2852
rect -28202 2779 -27106 2818
rect -28202 2745 -28189 2779
rect -28155 2745 -28115 2779
rect -28081 2745 -28041 2779
rect -28007 2745 -27967 2779
rect -27933 2745 -27893 2779
rect -27859 2745 -27819 2779
rect -27785 2745 -27745 2779
rect -27711 2745 -27671 2779
rect -27637 2745 -27597 2779
rect -27563 2745 -27523 2779
rect -27489 2745 -27449 2779
rect -27415 2745 -27375 2779
rect -27341 2745 -27301 2779
rect -27267 2745 -27227 2779
rect -27193 2745 -27153 2779
rect -27119 2745 -27106 2779
rect -28202 2706 -27106 2745
rect -28202 2672 -28189 2706
rect -28155 2672 -28115 2706
rect -28081 2672 -28041 2706
rect -28007 2672 -27967 2706
rect -27933 2672 -27893 2706
rect -27859 2672 -27819 2706
rect -27785 2672 -27745 2706
rect -27711 2672 -27671 2706
rect -27637 2672 -27597 2706
rect -27563 2672 -27523 2706
rect -27489 2672 -27449 2706
rect -27415 2672 -27375 2706
rect -27341 2672 -27301 2706
rect -27267 2672 -27227 2706
rect -27193 2672 -27153 2706
rect -27119 2672 -27106 2706
rect -28202 2633 -27106 2672
rect -28202 2599 -28189 2633
rect -28155 2599 -28115 2633
rect -28081 2599 -28041 2633
rect -28007 2599 -27967 2633
rect -27933 2599 -27893 2633
rect -27859 2599 -27819 2633
rect -27785 2599 -27745 2633
rect -27711 2599 -27671 2633
rect -27637 2599 -27597 2633
rect -27563 2599 -27523 2633
rect -27489 2599 -27449 2633
rect -27415 2599 -27375 2633
rect -27341 2599 -27301 2633
rect -27267 2599 -27227 2633
rect -27193 2599 -27153 2633
rect -27119 2599 -27106 2633
rect -28202 2560 -27106 2599
rect -28202 2526 -28189 2560
rect -28155 2526 -28115 2560
rect -28081 2526 -28041 2560
rect -28007 2526 -27967 2560
rect -27933 2526 -27893 2560
rect -27859 2526 -27819 2560
rect -27785 2526 -27745 2560
rect -27711 2526 -27671 2560
rect -27637 2526 -27597 2560
rect -27563 2526 -27523 2560
rect -27489 2526 -27449 2560
rect -27415 2526 -27375 2560
rect -27341 2526 -27301 2560
rect -27267 2526 -27227 2560
rect -27193 2526 -27153 2560
rect -27119 2526 -27106 2560
rect -28202 2487 -27106 2526
rect -28202 2453 -28189 2487
rect -28155 2453 -28115 2487
rect -28081 2453 -28041 2487
rect -28007 2453 -27967 2487
rect -27933 2453 -27893 2487
rect -27859 2453 -27819 2487
rect -27785 2453 -27745 2487
rect -27711 2453 -27671 2487
rect -27637 2453 -27597 2487
rect -27563 2453 -27523 2487
rect -27489 2453 -27449 2487
rect -27415 2453 -27375 2487
rect -27341 2453 -27301 2487
rect -27267 2453 -27227 2487
rect -27193 2453 -27153 2487
rect -27119 2453 -27106 2487
rect -28202 2414 -27106 2453
rect -28202 2380 -28189 2414
rect -28155 2380 -28115 2414
rect -28081 2380 -28041 2414
rect -28007 2380 -27967 2414
rect -27933 2380 -27893 2414
rect -27859 2380 -27819 2414
rect -27785 2380 -27745 2414
rect -27711 2380 -27671 2414
rect -27637 2380 -27597 2414
rect -27563 2380 -27523 2414
rect -27489 2380 -27449 2414
rect -27415 2380 -27375 2414
rect -27341 2380 -27301 2414
rect -27267 2380 -27227 2414
rect -27193 2380 -27153 2414
rect -27119 2380 -27106 2414
rect -28202 2341 -27106 2380
rect -28202 2307 -28189 2341
rect -28155 2307 -28115 2341
rect -28081 2307 -28041 2341
rect -28007 2307 -27967 2341
rect -27933 2307 -27893 2341
rect -27859 2307 -27819 2341
rect -27785 2307 -27745 2341
rect -27711 2307 -27671 2341
rect -27637 2307 -27597 2341
rect -27563 2307 -27523 2341
rect -27489 2307 -27449 2341
rect -27415 2307 -27375 2341
rect -27341 2307 -27301 2341
rect -27267 2307 -27227 2341
rect -27193 2307 -27153 2341
rect -27119 2307 -27106 2341
rect -28202 2268 -27106 2307
rect -28202 2234 -28189 2268
rect -28155 2234 -28115 2268
rect -28081 2234 -28041 2268
rect -28007 2234 -27967 2268
rect -27933 2234 -27893 2268
rect -27859 2234 -27819 2268
rect -27785 2234 -27745 2268
rect -27711 2234 -27671 2268
rect -27637 2234 -27597 2268
rect -27563 2234 -27523 2268
rect -27489 2234 -27449 2268
rect -27415 2234 -27375 2268
rect -27341 2234 -27301 2268
rect -27267 2234 -27227 2268
rect -27193 2234 -27153 2268
rect -27119 2234 -27106 2268
rect -28202 2195 -27106 2234
rect -28202 2161 -28189 2195
rect -28155 2161 -28115 2195
rect -28081 2161 -28041 2195
rect -28007 2161 -27967 2195
rect -27933 2161 -27893 2195
rect -27859 2161 -27819 2195
rect -27785 2161 -27745 2195
rect -27711 2161 -27671 2195
rect -27637 2161 -27597 2195
rect -27563 2161 -27523 2195
rect -27489 2161 -27449 2195
rect -27415 2161 -27375 2195
rect -27341 2161 -27301 2195
rect -27267 2161 -27227 2195
rect -27193 2161 -27153 2195
rect -27119 2161 -27106 2195
rect -28202 2122 -27106 2161
rect -28202 2088 -28189 2122
rect -28155 2088 -28115 2122
rect -28081 2088 -28041 2122
rect -28007 2088 -27967 2122
rect -27933 2088 -27893 2122
rect -27859 2088 -27819 2122
rect -27785 2088 -27745 2122
rect -27711 2088 -27671 2122
rect -27637 2088 -27597 2122
rect -27563 2088 -27523 2122
rect -27489 2088 -27449 2122
rect -27415 2088 -27375 2122
rect -27341 2088 -27301 2122
rect -27267 2088 -27227 2122
rect -27193 2088 -27153 2122
rect -27119 2088 -27106 2122
rect -28202 2049 -27106 2088
rect -28202 2015 -28189 2049
rect -28155 2015 -28115 2049
rect -28081 2015 -28041 2049
rect -28007 2015 -27967 2049
rect -27933 2015 -27893 2049
rect -27859 2015 -27819 2049
rect -27785 2015 -27745 2049
rect -27711 2015 -27671 2049
rect -27637 2015 -27597 2049
rect -27563 2015 -27523 2049
rect -27489 2015 -27449 2049
rect -27415 2015 -27375 2049
rect -27341 2015 -27301 2049
rect -27267 2015 -27227 2049
rect -27193 2015 -27153 2049
rect -27119 2015 -27106 2049
rect -28202 1976 -27106 2015
rect -28202 1942 -28189 1976
rect -28155 1942 -28115 1976
rect -28081 1942 -28041 1976
rect -28007 1942 -27967 1976
rect -27933 1942 -27893 1976
rect -27859 1942 -27819 1976
rect -27785 1942 -27745 1976
rect -27711 1942 -27671 1976
rect -27637 1942 -27597 1976
rect -27563 1942 -27523 1976
rect -27489 1942 -27449 1976
rect -27415 1942 -27375 1976
rect -27341 1942 -27301 1976
rect -27267 1942 -27227 1976
rect -27193 1942 -27153 1976
rect -27119 1942 -27106 1976
rect -28202 1903 -27106 1942
rect -28202 1869 -28189 1903
rect -28155 1869 -28115 1903
rect -28081 1869 -28041 1903
rect -28007 1869 -27967 1903
rect -27933 1869 -27893 1903
rect -27859 1869 -27819 1903
rect -27785 1869 -27745 1903
rect -27711 1869 -27671 1903
rect -27637 1869 -27597 1903
rect -27563 1869 -27523 1903
rect -27489 1869 -27449 1903
rect -27415 1869 -27375 1903
rect -27341 1869 -27301 1903
rect -27267 1869 -27227 1903
rect -27193 1869 -27153 1903
rect -27119 1869 -27106 1903
rect -28202 1830 -27106 1869
rect -28202 1796 -28189 1830
rect -28155 1796 -28115 1830
rect -28081 1796 -28041 1830
rect -28007 1796 -27967 1830
rect -27933 1796 -27893 1830
rect -27859 1796 -27819 1830
rect -27785 1796 -27745 1830
rect -27711 1796 -27671 1830
rect -27637 1796 -27597 1830
rect -27563 1796 -27523 1830
rect -27489 1796 -27449 1830
rect -27415 1796 -27375 1830
rect -27341 1796 -27301 1830
rect -27267 1796 -27227 1830
rect -27193 1796 -27153 1830
rect -27119 1796 -27106 1830
rect -28202 1757 -27106 1796
rect -28202 1723 -28189 1757
rect -28155 1723 -28115 1757
rect -28081 1723 -28041 1757
rect -28007 1723 -27967 1757
rect -27933 1723 -27893 1757
rect -27859 1723 -27819 1757
rect -27785 1723 -27745 1757
rect -27711 1723 -27671 1757
rect -27637 1723 -27597 1757
rect -27563 1723 -27523 1757
rect -27489 1723 -27449 1757
rect -27415 1723 -27375 1757
rect -27341 1723 -27301 1757
rect -27267 1723 -27227 1757
rect -27193 1723 -27153 1757
rect -27119 1723 -27106 1757
rect -28202 1684 -27106 1723
rect -28202 1650 -28189 1684
rect -28155 1650 -28115 1684
rect -28081 1650 -28041 1684
rect -28007 1650 -27967 1684
rect -27933 1650 -27893 1684
rect -27859 1650 -27819 1684
rect -27785 1650 -27745 1684
rect -27711 1650 -27671 1684
rect -27637 1650 -27597 1684
rect -27563 1650 -27523 1684
rect -27489 1650 -27449 1684
rect -27415 1650 -27375 1684
rect -27341 1650 -27301 1684
rect -27267 1650 -27227 1684
rect -27193 1650 -27153 1684
rect -27119 1650 -27106 1684
rect -28202 1611 -27106 1650
rect -28202 1577 -28189 1611
rect -28155 1577 -28115 1611
rect -28081 1577 -28041 1611
rect -28007 1577 -27967 1611
rect -27933 1577 -27893 1611
rect -27859 1577 -27819 1611
rect -27785 1577 -27745 1611
rect -27711 1577 -27671 1611
rect -27637 1577 -27597 1611
rect -27563 1577 -27523 1611
rect -27489 1577 -27449 1611
rect -27415 1577 -27375 1611
rect -27341 1577 -27301 1611
rect -27267 1577 -27227 1611
rect -27193 1577 -27153 1611
rect -27119 1577 -27106 1611
rect -28202 1538 -27106 1577
rect -28202 1504 -28189 1538
rect -28155 1504 -28115 1538
rect -28081 1504 -28041 1538
rect -28007 1504 -27967 1538
rect -27933 1504 -27893 1538
rect -27859 1504 -27819 1538
rect -27785 1504 -27745 1538
rect -27711 1504 -27671 1538
rect -27637 1504 -27597 1538
rect -27563 1504 -27523 1538
rect -27489 1504 -27449 1538
rect -27415 1504 -27375 1538
rect -27341 1504 -27301 1538
rect -27267 1504 -27227 1538
rect -27193 1504 -27153 1538
rect -27119 1504 -27106 1538
rect -28202 1465 -27106 1504
rect -28202 1431 -28189 1465
rect -28155 1431 -28115 1465
rect -28081 1431 -28041 1465
rect -28007 1431 -27967 1465
rect -27933 1431 -27893 1465
rect -27859 1431 -27819 1465
rect -27785 1431 -27745 1465
rect -27711 1431 -27671 1465
rect -27637 1431 -27597 1465
rect -27563 1431 -27523 1465
rect -27489 1431 -27449 1465
rect -27415 1431 -27375 1465
rect -27341 1431 -27301 1465
rect -27267 1431 -27227 1465
rect -27193 1431 -27153 1465
rect -27119 1431 -27106 1465
rect -28202 1392 -27106 1431
rect -28202 1358 -28189 1392
rect -28155 1358 -28115 1392
rect -28081 1358 -28041 1392
rect -28007 1358 -27967 1392
rect -27933 1358 -27893 1392
rect -27859 1358 -27819 1392
rect -27785 1358 -27745 1392
rect -27711 1358 -27671 1392
rect -27637 1358 -27597 1392
rect -27563 1358 -27523 1392
rect -27489 1358 -27449 1392
rect -27415 1358 -27375 1392
rect -27341 1358 -27301 1392
rect -27267 1358 -27227 1392
rect -27193 1358 -27153 1392
rect -27119 1358 -27106 1392
rect -28202 1319 -27106 1358
rect -28202 1285 -28189 1319
rect -28155 1285 -28115 1319
rect -28081 1285 -28041 1319
rect -28007 1285 -27967 1319
rect -27933 1285 -27893 1319
rect -27859 1285 -27819 1319
rect -27785 1285 -27745 1319
rect -27711 1285 -27671 1319
rect -27637 1285 -27597 1319
rect -27563 1285 -27523 1319
rect -27489 1285 -27449 1319
rect -27415 1285 -27375 1319
rect -27341 1285 -27301 1319
rect -27267 1285 -27227 1319
rect -27193 1285 -27153 1319
rect -27119 1285 -27106 1319
rect -28202 1246 -27106 1285
rect -28202 1212 -28189 1246
rect -28155 1212 -28115 1246
rect -28081 1212 -28041 1246
rect -28007 1212 -27967 1246
rect -27933 1212 -27893 1246
rect -27859 1212 -27819 1246
rect -27785 1212 -27745 1246
rect -27711 1212 -27671 1246
rect -27637 1212 -27597 1246
rect -27563 1212 -27523 1246
rect -27489 1212 -27449 1246
rect -27415 1212 -27375 1246
rect -27341 1212 -27301 1246
rect -27267 1212 -27227 1246
rect -27193 1212 -27153 1246
rect -27119 1212 -27106 1246
rect -28202 1173 -27106 1212
rect -28202 1139 -28189 1173
rect -28155 1139 -28115 1173
rect -28081 1139 -28041 1173
rect -28007 1139 -27967 1173
rect -27933 1139 -27893 1173
rect -27859 1139 -27819 1173
rect -27785 1139 -27745 1173
rect -27711 1139 -27671 1173
rect -27637 1139 -27597 1173
rect -27563 1139 -27523 1173
rect -27489 1139 -27449 1173
rect -27415 1139 -27375 1173
rect -27341 1139 -27301 1173
rect -27267 1139 -27227 1173
rect -27193 1139 -27153 1173
rect -27119 1139 -27106 1173
rect -28202 1100 -27106 1139
rect -28202 1066 -28189 1100
rect -28155 1066 -28115 1100
rect -28081 1066 -28041 1100
rect -28007 1066 -27967 1100
rect -27933 1066 -27893 1100
rect -27859 1066 -27819 1100
rect -27785 1066 -27745 1100
rect -27711 1066 -27671 1100
rect -27637 1066 -27597 1100
rect -27563 1066 -27523 1100
rect -27489 1066 -27449 1100
rect -27415 1066 -27375 1100
rect -27341 1066 -27301 1100
rect -27267 1066 -27227 1100
rect -27193 1066 -27153 1100
rect -27119 1066 -27106 1100
rect -28202 1028 -27106 1066
rect -28202 994 -28189 1028
rect -28155 994 -28115 1028
rect -28081 994 -28041 1028
rect -28007 994 -27967 1028
rect -27933 994 -27893 1028
rect -27859 994 -27819 1028
rect -27785 994 -27745 1028
rect -27711 994 -27671 1028
rect -27637 994 -27597 1028
rect -27563 994 -27523 1028
rect -27489 994 -27449 1028
rect -27415 994 -27375 1028
rect -27341 994 -27301 1028
rect -27267 994 -27227 1028
rect -27193 994 -27153 1028
rect -27119 994 -27106 1028
rect -28202 956 -27106 994
rect -28202 922 -28189 956
rect -28155 922 -28115 956
rect -28081 922 -28041 956
rect -28007 922 -27967 956
rect -27933 922 -27893 956
rect -27859 922 -27819 956
rect -27785 922 -27745 956
rect -27711 922 -27671 956
rect -27637 922 -27597 956
rect -27563 922 -27523 956
rect -27489 922 -27449 956
rect -27415 922 -27375 956
rect -27341 922 -27301 956
rect -27267 922 -27227 956
rect -27193 922 -27153 956
rect -27119 922 -27106 956
rect -28202 884 -27106 922
rect -28202 850 -28189 884
rect -28155 850 -28115 884
rect -28081 850 -28041 884
rect -28007 850 -27967 884
rect -27933 850 -27893 884
rect -27859 850 -27819 884
rect -27785 850 -27745 884
rect -27711 850 -27671 884
rect -27637 850 -27597 884
rect -27563 850 -27523 884
rect -27489 850 -27449 884
rect -27415 850 -27375 884
rect -27341 850 -27301 884
rect -27267 850 -27227 884
rect -27193 850 -27153 884
rect -27119 850 -27106 884
rect -28202 812 -27106 850
rect -28202 778 -28189 812
rect -28155 778 -28115 812
rect -28081 778 -28041 812
rect -28007 778 -27967 812
rect -27933 778 -27893 812
rect -27859 778 -27819 812
rect -27785 778 -27745 812
rect -27711 778 -27671 812
rect -27637 778 -27597 812
rect -27563 778 -27523 812
rect -27489 778 -27449 812
rect -27415 778 -27375 812
rect -27341 778 -27301 812
rect -27267 778 -27227 812
rect -27193 778 -27153 812
rect -27119 778 -27106 812
rect -28202 740 -27106 778
rect -28202 706 -28189 740
rect -28155 706 -28115 740
rect -28081 706 -28041 740
rect -28007 706 -27967 740
rect -27933 706 -27893 740
rect -27859 706 -27819 740
rect -27785 706 -27745 740
rect -27711 706 -27671 740
rect -27637 706 -27597 740
rect -27563 706 -27523 740
rect -27489 706 -27449 740
rect -27415 706 -27375 740
rect -27341 706 -27301 740
rect -27267 706 -27227 740
rect -27193 706 -27153 740
rect -27119 706 -27106 740
rect -28202 668 -27106 706
rect -28202 634 -28189 668
rect -28155 634 -28115 668
rect -28081 634 -28041 668
rect -28007 634 -27967 668
rect -27933 634 -27893 668
rect -27859 634 -27819 668
rect -27785 634 -27745 668
rect -27711 634 -27671 668
rect -27637 634 -27597 668
rect -27563 634 -27523 668
rect -27489 634 -27449 668
rect -27415 634 -27375 668
rect -27341 634 -27301 668
rect -27267 634 -27227 668
rect -27193 634 -27153 668
rect -27119 634 -27106 668
rect -28202 596 -27106 634
rect -28202 562 -28189 596
rect -28155 562 -28115 596
rect -28081 562 -28041 596
rect -28007 562 -27967 596
rect -27933 562 -27893 596
rect -27859 562 -27819 596
rect -27785 562 -27745 596
rect -27711 562 -27671 596
rect -27637 562 -27597 596
rect -27563 562 -27523 596
rect -27489 562 -27449 596
rect -27415 562 -27375 596
rect -27341 562 -27301 596
rect -27267 562 -27227 596
rect -27193 562 -27153 596
rect -27119 562 -27106 596
rect -28202 524 -27106 562
rect -28202 490 -28189 524
rect -28155 490 -28115 524
rect -28081 490 -28041 524
rect -28007 490 -27967 524
rect -27933 490 -27893 524
rect -27859 490 -27819 524
rect -27785 490 -27745 524
rect -27711 490 -27671 524
rect -27637 490 -27597 524
rect -27563 490 -27523 524
rect -27489 490 -27449 524
rect -27415 490 -27375 524
rect -27341 490 -27301 524
rect -27267 490 -27227 524
rect -27193 490 -27153 524
rect -27119 490 -27106 524
rect -28202 488 -27106 490
rect -28202 452 -28188 488
rect -28202 418 -28189 452
rect -28136 436 -28122 488
rect -28070 436 -28056 488
rect -28004 436 -27990 488
rect -27938 452 -27924 488
rect -27872 452 -27858 488
rect -27806 452 -27792 488
rect -27740 452 -27726 488
rect -27674 452 -27659 488
rect -27607 452 -27592 488
rect -27933 436 -27924 452
rect -27859 436 -27858 452
rect -27674 436 -27671 452
rect -27607 436 -27597 452
rect -27540 436 -27525 488
rect -27473 436 -27458 488
rect -27406 436 -27391 488
rect -27339 436 -27324 488
rect -27272 452 -27257 488
rect -27205 452 -27190 488
rect -27138 452 -27106 488
rect -27267 436 -27257 452
rect -27193 436 -27190 452
rect -28155 420 -28115 436
rect -28081 420 -28041 436
rect -28007 420 -27967 436
rect -27933 420 -27893 436
rect -27859 420 -27819 436
rect -27785 420 -27745 436
rect -27711 420 -27671 436
rect -27637 420 -27597 436
rect -27563 420 -27523 436
rect -27489 420 -27449 436
rect -27415 420 -27375 436
rect -27341 420 -27301 436
rect -27267 420 -27227 436
rect -27193 420 -27153 436
rect -28202 380 -28188 418
rect -28202 346 -28189 380
rect -28136 368 -28122 420
rect -28070 368 -28056 420
rect -28004 368 -27990 420
rect -27933 418 -27924 420
rect -27859 418 -27858 420
rect -27674 418 -27671 420
rect -27607 418 -27597 420
rect -27938 380 -27924 418
rect -27872 380 -27858 418
rect -27806 380 -27792 418
rect -27740 380 -27726 418
rect -27674 380 -27659 418
rect -27607 380 -27592 418
rect -27933 368 -27924 380
rect -27859 368 -27858 380
rect -27674 368 -27671 380
rect -27607 368 -27597 380
rect -27540 368 -27525 420
rect -27473 368 -27458 420
rect -27406 368 -27391 420
rect -27339 368 -27324 420
rect -27267 418 -27257 420
rect -27193 418 -27190 420
rect -27119 418 -27106 452
rect -27272 380 -27257 418
rect -27205 380 -27190 418
rect -27138 380 -27106 418
rect -27267 368 -27257 380
rect -27193 368 -27190 380
rect -28155 352 -28115 368
rect -28081 352 -28041 368
rect -28007 352 -27967 368
rect -27933 352 -27893 368
rect -27859 352 -27819 368
rect -27785 352 -27745 368
rect -27711 352 -27671 368
rect -27637 352 -27597 368
rect -27563 352 -27523 368
rect -27489 352 -27449 368
rect -27415 352 -27375 368
rect -27341 352 -27301 368
rect -27267 352 -27227 368
rect -27193 352 -27153 368
rect -28202 308 -28188 346
rect -28202 274 -28189 308
rect -28136 300 -28122 352
rect -28070 300 -28056 352
rect -28004 300 -27990 352
rect -27933 346 -27924 352
rect -27859 346 -27858 352
rect -27674 346 -27671 352
rect -27607 346 -27597 352
rect -27938 308 -27924 346
rect -27872 308 -27858 346
rect -27806 308 -27792 346
rect -27740 308 -27726 346
rect -27674 308 -27659 346
rect -27607 308 -27592 346
rect -27933 300 -27924 308
rect -27859 300 -27858 308
rect -27674 300 -27671 308
rect -27607 300 -27597 308
rect -27540 300 -27525 352
rect -27473 300 -27458 352
rect -27406 300 -27391 352
rect -27339 300 -27324 352
rect -27267 346 -27257 352
rect -27193 346 -27190 352
rect -27119 346 -27106 380
rect -27272 308 -27257 346
rect -27205 308 -27190 346
rect -27138 308 -27106 346
rect -27267 300 -27257 308
rect -27193 300 -27190 308
rect -28155 284 -28115 300
rect -28081 284 -28041 300
rect -28007 284 -27967 300
rect -27933 284 -27893 300
rect -27859 284 -27819 300
rect -27785 284 -27745 300
rect -27711 284 -27671 300
rect -27637 284 -27597 300
rect -27563 284 -27523 300
rect -27489 284 -27449 300
rect -27415 284 -27375 300
rect -27341 284 -27301 300
rect -27267 284 -27227 300
rect -27193 284 -27153 300
rect -28202 236 -28188 274
rect -28202 202 -28189 236
rect -28136 232 -28122 284
rect -28070 232 -28056 284
rect -28004 232 -27990 284
rect -27933 274 -27924 284
rect -27859 274 -27858 284
rect -27674 274 -27671 284
rect -27607 274 -27597 284
rect -27938 236 -27924 274
rect -27872 236 -27858 274
rect -27806 236 -27792 274
rect -27740 236 -27726 274
rect -27674 236 -27659 274
rect -27607 236 -27592 274
rect -27933 232 -27924 236
rect -27859 232 -27858 236
rect -27674 232 -27671 236
rect -27607 232 -27597 236
rect -27540 232 -27525 284
rect -27473 232 -27458 284
rect -27406 232 -27391 284
rect -27339 232 -27324 284
rect -27267 274 -27257 284
rect -27193 274 -27190 284
rect -27119 274 -27106 308
rect -27272 236 -27257 274
rect -27205 236 -27190 274
rect -27138 236 -27106 274
rect -27267 232 -27257 236
rect -27193 232 -27190 236
rect -28155 216 -28115 232
rect -28081 216 -28041 232
rect -28007 216 -27967 232
rect -27933 216 -27893 232
rect -27859 216 -27819 232
rect -27785 216 -27745 232
rect -27711 216 -27671 232
rect -27637 216 -27597 232
rect -27563 216 -27523 232
rect -27489 216 -27449 232
rect -27415 216 -27375 232
rect -27341 216 -27301 232
rect -27267 216 -27227 232
rect -27193 216 -27153 232
rect -28202 164 -28188 202
rect -28136 164 -28122 216
rect -28070 164 -28056 216
rect -28004 164 -27990 216
rect -27933 202 -27924 216
rect -27859 202 -27858 216
rect -27674 202 -27671 216
rect -27607 202 -27597 216
rect -27938 164 -27924 202
rect -27872 164 -27858 202
rect -27806 164 -27792 202
rect -27740 164 -27726 202
rect -27674 164 -27659 202
rect -27607 164 -27592 202
rect -27540 164 -27525 216
rect -27473 164 -27458 216
rect -27406 164 -27391 216
rect -27339 164 -27324 216
rect -27267 202 -27257 216
rect -27193 202 -27190 216
rect -27119 202 -27106 236
rect -27272 164 -27257 202
rect -27205 164 -27190 202
rect -27138 164 -27106 202
rect -28202 130 -28189 164
rect -28155 148 -28115 164
rect -28081 148 -28041 164
rect -28007 148 -27967 164
rect -27933 148 -27893 164
rect -27859 148 -27819 164
rect -27785 148 -27745 164
rect -27711 148 -27671 164
rect -27637 148 -27597 164
rect -27563 148 -27523 164
rect -27489 148 -27449 164
rect -27415 148 -27375 164
rect -27341 148 -27301 164
rect -27267 148 -27227 164
rect -27193 148 -27153 164
rect -28202 96 -28188 130
rect -28136 96 -28122 148
rect -28070 96 -28056 148
rect -28004 96 -27990 148
rect -27933 130 -27924 148
rect -27859 130 -27858 148
rect -27674 130 -27671 148
rect -27607 130 -27597 148
rect -27938 96 -27924 130
rect -27872 96 -27858 130
rect -27806 96 -27792 130
rect -27740 96 -27726 130
rect -27674 96 -27659 130
rect -27607 96 -27592 130
rect -27540 96 -27525 148
rect -27473 96 -27458 148
rect -27406 96 -27391 148
rect -27339 96 -27324 148
rect -27267 130 -27257 148
rect -27193 130 -27190 148
rect -27119 130 -27106 164
rect -27272 96 -27257 130
rect -27205 96 -27190 130
rect -27138 96 -27106 130
rect -28202 92 -27106 96
rect -28202 58 -28189 92
rect -28155 80 -28115 92
rect -28081 80 -28041 92
rect -28007 80 -27967 92
rect -27933 80 -27893 92
rect -27859 80 -27819 92
rect -27785 80 -27745 92
rect -27711 80 -27671 92
rect -27637 80 -27597 92
rect -27563 80 -27523 92
rect -27489 80 -27449 92
rect -27415 80 -27375 92
rect -27341 80 -27301 92
rect -27267 80 -27227 92
rect -27193 80 -27153 92
rect -28202 28 -28188 58
rect -28136 28 -28122 80
rect -28070 28 -28056 80
rect -28004 28 -27990 80
rect -27933 58 -27924 80
rect -27859 58 -27858 80
rect -27674 58 -27671 80
rect -27607 58 -27597 80
rect -27938 28 -27924 58
rect -27872 28 -27858 58
rect -27806 28 -27792 58
rect -27740 28 -27726 58
rect -27674 28 -27659 58
rect -27607 28 -27592 58
rect -27540 28 -27525 80
rect -27473 28 -27458 80
rect -27406 28 -27391 80
rect -27339 28 -27324 80
rect -27267 58 -27257 80
rect -27193 58 -27190 80
rect -27119 58 -27106 92
rect -27272 28 -27257 58
rect -27205 28 -27190 58
rect -27138 28 -27106 58
rect -28202 20 -27106 28
rect -28202 -14 -28189 20
rect -28155 12 -28115 20
rect -28081 12 -28041 20
rect -28007 12 -27967 20
rect -27933 12 -27893 20
rect -27859 12 -27819 20
rect -27785 12 -27745 20
rect -27711 12 -27671 20
rect -27637 12 -27597 20
rect -27563 12 -27523 20
rect -27489 12 -27449 20
rect -27415 12 -27375 20
rect -27341 12 -27301 20
rect -27267 12 -27227 20
rect -27193 12 -27153 20
rect -28202 -40 -28188 -14
rect -28136 -40 -28122 12
rect -28070 -40 -28056 12
rect -28004 -40 -27990 12
rect -27933 -14 -27924 12
rect -27859 -14 -27858 12
rect -27674 -14 -27671 12
rect -27607 -14 -27597 12
rect -27938 -40 -27924 -14
rect -27872 -40 -27858 -14
rect -27806 -40 -27792 -14
rect -27740 -40 -27726 -14
rect -27674 -40 -27659 -14
rect -27607 -40 -27592 -14
rect -27540 -40 -27525 12
rect -27473 -40 -27458 12
rect -27406 -40 -27391 12
rect -27339 -40 -27324 12
rect -27267 -14 -27257 12
rect -27193 -14 -27190 12
rect -27119 -14 -27106 20
rect -27272 -40 -27257 -14
rect -27205 -40 -27190 -14
rect -27138 -40 -27106 -14
rect -28202 -52 -27106 -40
rect -28202 -86 -28189 -52
rect -28155 -56 -28115 -52
rect -28081 -56 -28041 -52
rect -28007 -56 -27967 -52
rect -27933 -56 -27893 -52
rect -27859 -56 -27819 -52
rect -27785 -56 -27745 -52
rect -27711 -56 -27671 -52
rect -27637 -56 -27597 -52
rect -27563 -56 -27523 -52
rect -27489 -56 -27449 -52
rect -27415 -56 -27375 -52
rect -27341 -56 -27301 -52
rect -27267 -56 -27227 -52
rect -27193 -56 -27153 -52
rect -28202 -108 -28188 -86
rect -28136 -108 -28122 -56
rect -28070 -108 -28056 -56
rect -28004 -108 -27990 -56
rect -27933 -86 -27924 -56
rect -27859 -86 -27858 -56
rect -27674 -86 -27671 -56
rect -27607 -86 -27597 -56
rect -27938 -108 -27924 -86
rect -27872 -108 -27858 -86
rect -27806 -108 -27792 -86
rect -27740 -108 -27726 -86
rect -27674 -108 -27659 -86
rect -27607 -108 -27592 -86
rect -27540 -108 -27525 -56
rect -27473 -108 -27458 -56
rect -27406 -108 -27391 -56
rect -27339 -108 -27324 -56
rect -27267 -86 -27257 -56
rect -27193 -86 -27190 -56
rect -27119 -86 -27106 -52
rect -27272 -108 -27257 -86
rect -27205 -108 -27190 -86
rect -27138 -108 -27106 -86
rect -28202 -124 -27106 -108
rect -28202 -158 -28189 -124
rect -28202 -176 -28188 -158
rect -28136 -176 -28122 -124
rect -28070 -176 -28056 -124
rect -28004 -176 -27990 -124
rect -27933 -158 -27924 -124
rect -27859 -158 -27858 -124
rect -27674 -158 -27671 -124
rect -27607 -158 -27597 -124
rect -27938 -176 -27924 -158
rect -27872 -176 -27858 -158
rect -27806 -176 -27792 -158
rect -27740 -176 -27726 -158
rect -27674 -176 -27659 -158
rect -27607 -176 -27592 -158
rect -27540 -176 -27525 -124
rect -27473 -176 -27458 -124
rect -27406 -176 -27391 -124
rect -27339 -176 -27324 -124
rect -27267 -158 -27257 -124
rect -27193 -158 -27190 -124
rect -27119 -158 -27106 -124
rect -27272 -176 -27257 -158
rect -27205 -176 -27190 -158
rect -27138 -176 -27106 -158
rect -28202 -192 -27106 -176
rect -28202 -196 -28188 -192
rect -28202 -230 -28189 -196
rect -28202 -244 -28188 -230
rect -28136 -244 -28122 -192
rect -28070 -244 -28056 -192
rect -28004 -244 -27990 -192
rect -27938 -196 -27924 -192
rect -27872 -196 -27858 -192
rect -27806 -196 -27792 -192
rect -27740 -196 -27726 -192
rect -27674 -196 -27659 -192
rect -27607 -196 -27592 -192
rect -27933 -230 -27924 -196
rect -27859 -230 -27858 -196
rect -27674 -230 -27671 -196
rect -27607 -230 -27597 -196
rect -27938 -244 -27924 -230
rect -27872 -244 -27858 -230
rect -27806 -244 -27792 -230
rect -27740 -244 -27726 -230
rect -27674 -244 -27659 -230
rect -27607 -244 -27592 -230
rect -27540 -244 -27525 -192
rect -27473 -244 -27458 -192
rect -27406 -244 -27391 -192
rect -27339 -244 -27324 -192
rect -27272 -196 -27257 -192
rect -27205 -196 -27190 -192
rect -27138 -196 -27106 -192
rect -27267 -230 -27257 -196
rect -27193 -230 -27190 -196
rect -27119 -230 -27106 -196
rect -27272 -244 -27257 -230
rect -27205 -244 -27190 -230
rect -27138 -244 -27106 -230
rect -28202 -260 -27106 -244
rect -28202 -268 -28188 -260
rect -28202 -302 -28189 -268
rect -28202 -312 -28188 -302
rect -28136 -312 -28122 -260
rect -28070 -312 -28056 -260
rect -28004 -312 -27990 -260
rect -27938 -268 -27924 -260
rect -27872 -268 -27858 -260
rect -27806 -268 -27792 -260
rect -27740 -268 -27726 -260
rect -27674 -268 -27659 -260
rect -27607 -268 -27592 -260
rect -27933 -302 -27924 -268
rect -27859 -302 -27858 -268
rect -27674 -302 -27671 -268
rect -27607 -302 -27597 -268
rect -27938 -312 -27924 -302
rect -27872 -312 -27858 -302
rect -27806 -312 -27792 -302
rect -27740 -312 -27726 -302
rect -27674 -312 -27659 -302
rect -27607 -312 -27592 -302
rect -27540 -312 -27525 -260
rect -27473 -312 -27458 -260
rect -27406 -312 -27391 -260
rect -27339 -312 -27324 -260
rect -27272 -268 -27257 -260
rect -27205 -268 -27190 -260
rect -27138 -268 -27106 -260
rect -27267 -302 -27257 -268
rect -27193 -302 -27190 -268
rect -27119 -302 -27106 -268
rect -27272 -312 -27257 -302
rect -27205 -312 -27190 -302
rect -27138 -312 -27106 -302
rect -28202 -328 -27106 -312
rect -28202 -340 -28188 -328
rect -28202 -374 -28189 -340
rect -28202 -380 -28188 -374
rect -28136 -380 -28122 -328
rect -28070 -380 -28056 -328
rect -28004 -380 -27990 -328
rect -27938 -340 -27924 -328
rect -27872 -340 -27858 -328
rect -27806 -340 -27792 -328
rect -27740 -340 -27726 -328
rect -27674 -340 -27659 -328
rect -27607 -340 -27592 -328
rect -27933 -374 -27924 -340
rect -27859 -374 -27858 -340
rect -27674 -374 -27671 -340
rect -27607 -374 -27597 -340
rect -27938 -380 -27924 -374
rect -27872 -380 -27858 -374
rect -27806 -380 -27792 -374
rect -27740 -380 -27726 -374
rect -27674 -380 -27659 -374
rect -27607 -380 -27592 -374
rect -27540 -380 -27525 -328
rect -27473 -380 -27458 -328
rect -27406 -380 -27391 -328
rect -27339 -380 -27324 -328
rect -27272 -340 -27257 -328
rect -27205 -340 -27190 -328
rect -27138 -340 -27106 -328
rect -27267 -374 -27257 -340
rect -27193 -374 -27190 -340
rect -27119 -374 -27106 -340
rect -27272 -380 -27257 -374
rect -27205 -380 -27190 -374
rect -27138 -380 -27106 -374
rect -28202 -412 -27106 -380
rect -28202 -446 -28189 -412
rect -28155 -446 -28115 -412
rect -28081 -446 -28041 -412
rect -28007 -446 -27967 -412
rect -27933 -446 -27893 -412
rect -27859 -446 -27819 -412
rect -27785 -446 -27745 -412
rect -27711 -446 -27671 -412
rect -27637 -446 -27597 -412
rect -27563 -446 -27523 -412
rect -27489 -446 -27449 -412
rect -27415 -446 -27375 -412
rect -27341 -446 -27301 -412
rect -27267 -446 -27227 -412
rect -27193 -446 -27153 -412
rect -27119 -446 -27106 -412
rect -28202 -484 -27106 -446
rect -28202 -518 -28189 -484
rect -28155 -518 -28115 -484
rect -28081 -518 -28041 -484
rect -28007 -518 -27967 -484
rect -27933 -518 -27893 -484
rect -27859 -518 -27819 -484
rect -27785 -518 -27745 -484
rect -27711 -518 -27671 -484
rect -27637 -518 -27597 -484
rect -27563 -518 -27523 -484
rect -27489 -518 -27449 -484
rect -27415 -518 -27375 -484
rect -27341 -518 -27301 -484
rect -27267 -518 -27227 -484
rect -27193 -518 -27153 -484
rect -27119 -518 -27106 -484
rect -28202 -556 -27106 -518
rect -28202 -590 -28189 -556
rect -28155 -590 -28115 -556
rect -28081 -590 -28041 -556
rect -28007 -590 -27967 -556
rect -27933 -590 -27893 -556
rect -27859 -590 -27819 -556
rect -27785 -590 -27745 -556
rect -27711 -590 -27671 -556
rect -27637 -590 -27597 -556
rect -27563 -590 -27523 -556
rect -27489 -590 -27449 -556
rect -27415 -590 -27375 -556
rect -27341 -590 -27301 -556
rect -27267 -590 -27227 -556
rect -27193 -590 -27153 -556
rect -27119 -590 -27106 -556
rect -28202 -628 -27106 -590
rect -28202 -662 -28189 -628
rect -28155 -662 -28115 -628
rect -28081 -662 -28041 -628
rect -28007 -662 -27967 -628
rect -27933 -662 -27893 -628
rect -27859 -662 -27819 -628
rect -27785 -662 -27745 -628
rect -27711 -662 -27671 -628
rect -27637 -662 -27597 -628
rect -27563 -662 -27523 -628
rect -27489 -662 -27449 -628
rect -27415 -662 -27375 -628
rect -27341 -662 -27301 -628
rect -27267 -662 -27227 -628
rect -27193 -662 -27153 -628
rect -27119 -662 -27106 -628
rect -28202 -700 -27106 -662
rect -28202 -734 -28189 -700
rect -28155 -734 -28115 -700
rect -28081 -734 -28041 -700
rect -28007 -734 -27967 -700
rect -27933 -734 -27893 -700
rect -27859 -734 -27819 -700
rect -27785 -734 -27745 -700
rect -27711 -734 -27671 -700
rect -27637 -734 -27597 -700
rect -27563 -734 -27523 -700
rect -27489 -734 -27449 -700
rect -27415 -734 -27375 -700
rect -27341 -734 -27301 -700
rect -27267 -734 -27227 -700
rect -27193 -734 -27153 -700
rect -27119 -734 -27106 -700
rect -28202 -772 -27106 -734
rect -28202 -806 -28189 -772
rect -28155 -806 -28115 -772
rect -28081 -806 -28041 -772
rect -28007 -806 -27967 -772
rect -27933 -806 -27893 -772
rect -27859 -806 -27819 -772
rect -27785 -806 -27745 -772
rect -27711 -806 -27671 -772
rect -27637 -806 -27597 -772
rect -27563 -806 -27523 -772
rect -27489 -806 -27449 -772
rect -27415 -806 -27375 -772
rect -27341 -806 -27301 -772
rect -27267 -806 -27227 -772
rect -27193 -806 -27153 -772
rect -27119 -806 -27106 -772
rect -28202 -844 -27106 -806
rect -28202 -878 -28189 -844
rect -28155 -878 -28115 -844
rect -28081 -878 -28041 -844
rect -28007 -878 -27967 -844
rect -27933 -878 -27893 -844
rect -27859 -878 -27819 -844
rect -27785 -878 -27745 -844
rect -27711 -878 -27671 -844
rect -27637 -878 -27597 -844
rect -27563 -878 -27523 -844
rect -27489 -878 -27449 -844
rect -27415 -878 -27375 -844
rect -27341 -878 -27301 -844
rect -27267 -878 -27227 -844
rect -27193 -878 -27153 -844
rect -27119 -878 -27106 -844
rect -28202 -916 -27106 -878
rect -28202 -950 -28189 -916
rect -28155 -950 -28115 -916
rect -28081 -950 -28041 -916
rect -28007 -950 -27967 -916
rect -27933 -950 -27893 -916
rect -27859 -950 -27819 -916
rect -27785 -950 -27745 -916
rect -27711 -950 -27671 -916
rect -27637 -950 -27597 -916
rect -27563 -950 -27523 -916
rect -27489 -950 -27449 -916
rect -27415 -950 -27375 -916
rect -27341 -950 -27301 -916
rect -27267 -950 -27227 -916
rect -27193 -950 -27153 -916
rect -27119 -950 -27106 -916
rect -28202 -988 -27106 -950
rect -28202 -1022 -28189 -988
rect -28155 -1022 -28115 -988
rect -28081 -1022 -28041 -988
rect -28007 -1022 -27967 -988
rect -27933 -1022 -27893 -988
rect -27859 -1022 -27819 -988
rect -27785 -1022 -27745 -988
rect -27711 -1022 -27671 -988
rect -27637 -1022 -27597 -988
rect -27563 -1022 -27523 -988
rect -27489 -1022 -27449 -988
rect -27415 -1022 -27375 -988
rect -27341 -1022 -27301 -988
rect -27267 -1022 -27227 -988
rect -27193 -1022 -27153 -988
rect -27119 -1022 -27106 -988
rect -28202 -1060 -27106 -1022
rect -9796 4312 -9750 4324
rect -9796 4278 -9790 4312
rect -9756 4278 -9750 4312
rect -9796 4240 -9750 4278
rect -9796 4206 -9790 4240
rect -9756 4206 -9750 4240
rect -9796 -1015 -9750 4206
rect 3932 3840 5778 3846
rect 3932 3806 4010 3840
rect 4044 3806 4082 3840
rect 4116 3806 4154 3840
rect 4188 3806 4226 3840
rect 4260 3806 4298 3840
rect 4332 3806 4370 3840
rect 4404 3806 4442 3840
rect 4476 3806 4514 3840
rect 4548 3806 4586 3840
rect 4620 3806 4658 3840
rect 4692 3806 4730 3840
rect 4764 3806 4802 3840
rect 4836 3806 4874 3840
rect 4908 3806 4946 3840
rect 4980 3806 5018 3840
rect 5052 3806 5090 3840
rect 5124 3806 5162 3840
rect 5196 3806 5234 3840
rect 5268 3806 5306 3840
rect 5340 3806 5378 3840
rect 5412 3806 5450 3840
rect 5484 3806 5522 3840
rect 5556 3806 5594 3840
rect 5628 3806 5666 3840
rect 5700 3806 5778 3840
rect 3932 3800 5778 3806
rect 3932 3768 3978 3800
rect 3932 3734 3938 3768
rect 3972 3734 3978 3768
rect -793 3648 -787 3700
rect -735 3688 -717 3700
rect -665 3688 -646 3700
rect -594 3688 -575 3700
rect -523 3688 -504 3700
rect -452 3694 -446 3700
rect -452 3688 -389 3694
rect -723 3654 -717 3688
rect -523 3654 -516 3688
rect -452 3654 -435 3688
rect -401 3654 -389 3688
rect -735 3648 -717 3654
rect -665 3648 -646 3654
rect -594 3648 -575 3654
rect -523 3648 -504 3654
rect -452 3648 -389 3654
rect -597 3617 -545 3648
rect 159 3645 170 3697
rect 222 3645 235 3697
rect 287 3645 300 3697
rect 352 3645 365 3697
rect 417 3688 430 3697
rect 482 3688 495 3697
rect 547 3688 560 3697
rect 612 3688 625 3697
rect 677 3688 690 3697
rect 424 3654 430 3688
rect 677 3654 682 3688
rect 417 3645 430 3654
rect 482 3645 495 3654
rect 547 3645 560 3654
rect 612 3645 625 3654
rect 677 3645 690 3654
rect 742 3645 755 3697
rect 807 3645 820 3697
rect 872 3645 885 3697
rect 937 3645 950 3697
rect 1002 3688 1015 3697
rect 1067 3688 1080 3697
rect 1132 3688 1145 3697
rect 1197 3688 1210 3697
rect 1262 3688 1275 3697
rect 1327 3688 1340 3697
rect 1008 3654 1015 3688
rect 1262 3654 1266 3688
rect 1327 3654 1339 3688
rect 1002 3645 1015 3654
rect 1067 3645 1080 3654
rect 1132 3645 1145 3654
rect 1197 3645 1210 3654
rect 1262 3645 1275 3654
rect 1327 3645 1340 3654
rect 1392 3645 1405 3697
rect 1457 3645 1470 3697
rect 1522 3645 1535 3697
rect 1587 3688 1600 3697
rect 1652 3688 1665 3697
rect 1717 3688 1730 3697
rect 1782 3688 1795 3697
rect 1847 3688 1860 3697
rect 1912 3688 1925 3697
rect 1592 3654 1600 3688
rect 1847 3654 1850 3688
rect 1912 3654 1923 3688
rect 1587 3645 1600 3654
rect 1652 3645 1665 3654
rect 1717 3645 1730 3654
rect 1782 3645 1795 3654
rect 1847 3645 1860 3654
rect 1912 3645 1925 3654
rect 1977 3645 1990 3697
rect 2042 3645 2055 3697
rect 2107 3645 2120 3697
rect 2172 3688 2185 3697
rect 2237 3688 2250 3697
rect 2302 3688 2315 3697
rect 2367 3688 2380 3697
rect 2432 3688 2445 3697
rect 2497 3688 2510 3697
rect 2562 3688 2575 3697
rect 2173 3654 2185 3688
rect 2245 3654 2250 3688
rect 2497 3654 2499 3688
rect 2562 3654 2571 3688
rect 2172 3645 2185 3654
rect 2237 3645 2250 3654
rect 2302 3645 2315 3654
rect 2367 3645 2380 3654
rect 2432 3645 2445 3654
rect 2497 3645 2510 3654
rect 2562 3645 2575 3654
rect 2627 3645 2640 3697
rect 2692 3645 2705 3697
rect 2757 3645 2770 3697
rect 2822 3645 2835 3697
rect 2887 3688 2900 3697
rect 2952 3688 2965 3697
rect 3017 3688 3030 3697
rect 3082 3688 3095 3697
rect 3147 3688 3160 3697
rect 3212 3688 3224 3697
rect 2893 3654 2900 3688
rect 3212 3654 3219 3688
rect 2887 3645 2900 3654
rect 2952 3645 2965 3654
rect 3017 3645 3030 3654
rect 3082 3645 3095 3654
rect 3147 3645 3160 3654
rect 3212 3645 3224 3654
rect 3276 3645 3288 3697
rect 3340 3645 3352 3697
rect 3404 3645 3416 3697
rect 3468 3688 3480 3697
rect 3532 3688 3553 3697
rect 3469 3654 3480 3688
rect 3541 3654 3553 3688
rect 3468 3645 3480 3654
rect 3532 3645 3553 3654
rect 3932 3692 3978 3734
rect 3932 3658 3938 3692
rect 3972 3658 3978 3692
rect 4712 3753 4926 3800
rect 4712 3719 4718 3753
rect 4752 3719 4802 3753
rect 4836 3719 4886 3753
rect 4920 3719 4926 3753
rect 4712 3678 4926 3719
rect 5732 3758 5778 3800
rect 5732 3724 5738 3758
rect 5772 3724 5778 3758
rect 3932 3616 3978 3658
rect 3932 3582 3938 3616
rect 3972 3582 3978 3616
rect -929 3546 -706 3558
rect -929 3512 -746 3546
rect -712 3512 -706 3546
rect -929 3474 -706 3512
rect -929 3440 -746 3474
rect -712 3440 -706 3474
rect -929 3402 -706 3440
rect -929 3368 -746 3402
rect -712 3368 -706 3402
rect -929 3330 -706 3368
rect -929 3296 -746 3330
rect -712 3296 -706 3330
rect -929 3258 -706 3296
rect -929 3224 -746 3258
rect -712 3224 -706 3258
rect -929 3186 -706 3224
rect -929 3152 -746 3186
rect -712 3152 -706 3186
rect -929 3114 -706 3152
rect -929 3080 -746 3114
rect -712 3080 -706 3114
rect -929 3042 -706 3080
rect -929 3008 -746 3042
rect -712 3008 -706 3042
rect -929 2970 -706 3008
rect -929 2936 -746 2970
rect -712 2936 -706 2970
rect -929 2898 -706 2936
rect -929 2864 -746 2898
rect -712 2864 -706 2898
rect -929 2826 -706 2864
rect -929 2792 -746 2826
rect -712 2792 -706 2826
rect -929 2754 -706 2792
rect -929 2720 -746 2754
rect -712 2720 -706 2754
rect -929 2682 -706 2720
rect -929 2648 -746 2682
rect -712 2648 -706 2682
rect -929 2610 -706 2648
rect -929 2576 -746 2610
rect -712 2576 -706 2610
rect -929 2564 -706 2576
rect -597 3550 -545 3565
rect -597 3483 -545 3498
rect -597 3416 -545 3431
rect -597 3349 -545 3364
rect -597 3296 -590 3297
rect -556 3296 -545 3297
rect -597 3283 -545 3296
rect -597 3224 -590 3231
rect -556 3224 -545 3231
rect -597 3217 -545 3224
rect -597 3152 -590 3165
rect -556 3152 -545 3165
rect -597 3151 -545 3152
rect -597 3085 -590 3099
rect -556 3085 -545 3099
rect -597 3019 -590 3033
rect -556 3019 -545 3033
rect -597 2953 -590 2967
rect -556 2953 -545 2967
rect -597 2898 -545 2901
rect -597 2887 -590 2898
rect -556 2887 -545 2898
rect -597 2826 -545 2835
rect -597 2821 -590 2826
rect -556 2821 -545 2826
rect -597 2755 -545 2769
rect -597 2689 -545 2703
rect -597 2623 -545 2637
rect -597 2564 -545 2571
rect -440 3546 -258 3558
rect -440 3512 -434 3546
rect -400 3512 -258 3546
rect -440 3474 -258 3512
rect -440 3440 -434 3474
rect -400 3440 -258 3474
rect -440 3402 -258 3440
rect -440 3368 -434 3402
rect -400 3368 -258 3402
rect -440 3330 -258 3368
rect -440 3296 -434 3330
rect -400 3296 -258 3330
rect -440 3258 -258 3296
rect -440 3224 -434 3258
rect -400 3224 -258 3258
rect -440 3186 -258 3224
rect -440 3152 -434 3186
rect -400 3152 -258 3186
rect -440 3114 -258 3152
rect -440 3080 -434 3114
rect -400 3080 -258 3114
rect -440 3042 -258 3080
rect -440 3008 -434 3042
rect -400 3008 -258 3042
rect -440 2970 -258 3008
rect -440 2936 -434 2970
rect -400 2936 -258 2970
rect -440 2898 -258 2936
rect -440 2864 -434 2898
rect -400 2864 -258 2898
rect -440 2826 -258 2864
rect -440 2792 -434 2826
rect -400 2792 -258 2826
rect -440 2754 -258 2792
rect -440 2720 -434 2754
rect -400 2720 -258 2754
rect -440 2682 -258 2720
rect -440 2648 -434 2682
rect -400 2648 -258 2682
rect -440 2610 -258 2648
rect -440 2576 -434 2610
rect -400 2576 -258 2610
rect -440 2564 -258 2576
rect -929 2541 -775 2564
tri -775 2541 -752 2564 nw
tri -440 2541 -417 2564 ne
rect -417 2541 -258 2564
rect -929 2529 -787 2541
tri -787 2529 -775 2541 nw
tri -417 2529 -405 2541 ne
rect -405 2529 -258 2541
rect -929 2523 -793 2529
tri -793 2523 -787 2529 nw
rect -702 2523 -459 2529
rect -929 2489 -827 2523
tri -827 2489 -793 2523 nw
rect -702 2489 -690 2523
rect -656 2489 -617 2523
rect -583 2489 -543 2523
rect -509 2489 -459 2523
tri -405 2521 -397 2529 ne
rect -397 2521 -258 2529
tri -397 2517 -393 2521 ne
rect -393 2517 -258 2521
tri -393 2516 -392 2517 ne
rect -392 2516 -258 2517
tri -392 2503 -379 2516 ne
rect -379 2503 -258 2516
rect -929 2469 -847 2489
tri -847 2469 -827 2489 nw
rect -702 2483 -459 2489
tri -595 2469 -581 2483 ne
rect -581 2469 -459 2483
tri -379 2469 -345 2503 ne
rect -345 2469 -258 2503
rect -929 2447 -869 2469
tri -869 2447 -847 2469 nw
tri -581 2447 -559 2469 ne
rect -559 2447 -459 2469
tri -345 2447 -323 2469 ne
rect -323 2447 -258 2469
rect -929 2446 -870 2447
tri -870 2446 -869 2447 nw
tri -559 2446 -558 2447 ne
rect -558 2446 -459 2447
tri -323 2446 -322 2447 ne
rect -322 2446 -258 2447
rect -929 2444 -872 2446
tri -872 2444 -870 2446 nw
tri -558 2444 -556 2446 ne
rect -556 2444 -459 2446
tri -322 2444 -320 2446 ne
rect -320 2444 -258 2446
rect -1709 2213 -1703 2265
rect -1651 2213 -1639 2265
rect -1587 2213 -1581 2265
tri -1679 2207 -1673 2213 ne
rect -1673 2207 -1581 2213
tri -1673 2205 -1671 2207 ne
rect -1671 2205 -1581 2207
tri -1671 2181 -1647 2205 ne
rect -1647 2181 -1581 2205
tri -1647 2178 -1644 2181 ne
rect -1644 2178 -1581 2181
rect -1761 2172 -1709 2178
tri -1644 2169 -1635 2178 ne
rect -1635 2169 -1581 2178
tri -1635 2161 -1627 2169 ne
rect -1761 2108 -1709 2120
tri -1827 -493 -1761 -427 se
rect -1761 -441 -1709 2056
tri -1761 -493 -1709 -441 nw
tri -1893 -559 -1827 -493 se
tri -1827 -559 -1761 -493 nw
tri -1630 -559 -1627 -556 se
rect -1627 -559 -1581 2169
rect -929 714 -873 2444
tri -873 2443 -872 2444 nw
tri -556 2443 -555 2444 ne
rect -555 2443 -459 2444
tri -555 2431 -543 2443 ne
rect -543 2431 -459 2443
tri -320 2434 -310 2444 ne
tri -543 2413 -525 2431 ne
rect -525 2413 -459 2431
tri -525 2397 -509 2413 ne
rect -509 2397 -459 2413
tri -459 2397 -443 2413 sw
tri -509 2375 -487 2397 ne
rect -487 2375 -443 2397
tri -443 2375 -421 2397 sw
tri -487 2365 -477 2375 ne
rect -477 2365 -421 2375
tri -421 2365 -411 2375 sw
tri -477 2359 -471 2365 ne
rect -471 2359 -411 2365
tri -411 2359 -405 2365 sw
tri -471 2347 -459 2359 ne
rect -459 2347 -405 2359
tri -459 2331 -443 2347 ne
rect -443 2331 -405 2347
tri -405 2331 -377 2359 sw
tri -443 2328 -440 2331 ne
rect -440 2328 -377 2331
tri -377 2328 -374 2331 sw
tri -440 2294 -406 2328 ne
rect -406 2294 -374 2328
tri -374 2294 -340 2328 sw
tri -406 2293 -405 2294 ne
rect -405 2293 -340 2294
tri -340 2293 -339 2294 sw
tri -405 2289 -401 2293 ne
rect -401 2289 -339 2293
tri -401 2273 -385 2289 ne
rect -841 2271 -457 2272
rect -841 2219 -805 2271
rect -753 2219 -739 2271
rect -687 2219 -673 2271
rect -621 2219 -606 2271
rect -554 2219 -539 2271
rect -487 2219 -457 2271
rect -841 2177 -457 2219
rect -841 2125 -805 2177
rect -753 2125 -739 2177
rect -687 2125 -673 2177
rect -621 2125 -606 2177
rect -554 2125 -539 2177
rect -487 2125 -457 2177
rect -841 2089 -457 2125
tri -407 1873 -385 1895 se
rect -385 1875 -339 2289
rect -385 1873 -341 1875
tri -341 1873 -339 1875 nw
tri -411 1869 -407 1873 se
rect -407 1869 -345 1873
tri -345 1869 -341 1873 nw
tri -413 1867 -411 1869 se
rect -411 1867 -347 1869
tri -347 1867 -345 1869 nw
tri -447 1833 -413 1867 se
rect -413 1833 -381 1867
tri -381 1833 -347 1867 nw
tri -451 1829 -447 1833 se
rect -447 1829 -385 1833
tri -385 1829 -381 1833 nw
tri -460 1820 -451 1829 se
rect -451 1820 -394 1829
tri -394 1820 -385 1829 nw
tri -485 1795 -460 1820 se
rect -460 1795 -419 1820
tri -419 1795 -394 1820 nw
tri -517 1763 -485 1795 se
rect -485 1763 -451 1795
tri -451 1763 -419 1795 nw
tri -519 1761 -517 1763 se
rect -517 1761 -453 1763
tri -453 1761 -451 1763 nw
tri -532 1748 -519 1761 se
rect -519 1748 -466 1761
tri -466 1748 -453 1761 nw
tri -536 1744 -532 1748 se
rect -532 1744 -470 1748
tri -470 1744 -466 1748 nw
rect -536 1741 -473 1744
tri -473 1741 -470 1744 nw
rect -536 1703 -490 1741
tri -490 1724 -473 1741 nw
rect -722 1647 -716 1699
rect -664 1647 -650 1699
rect -598 1647 -592 1699
rect -536 1669 -530 1703
rect -496 1669 -490 1703
rect -536 1631 -490 1669
rect -536 1597 -530 1631
rect -496 1597 -490 1631
rect -536 1585 -490 1597
rect -731 1400 -440 1423
rect -731 1348 -725 1400
rect -673 1348 -650 1400
rect -598 1348 -574 1400
rect -522 1348 -498 1400
rect -446 1348 -440 1400
rect -731 1325 -440 1348
rect -310 1299 -258 2444
rect 162 3546 208 3558
rect 162 3512 168 3546
rect 202 3512 208 3546
rect 162 3474 208 3512
rect 162 3440 168 3474
rect 202 3440 208 3474
rect 162 3402 208 3440
rect 162 3368 168 3402
rect 202 3368 208 3402
rect 315 3557 367 3563
rect 315 3493 367 3505
rect 315 3440 324 3441
rect 358 3440 367 3441
rect 315 3429 367 3440
rect 315 3371 324 3377
tri 315 3368 318 3371 ne
rect 318 3368 324 3371
rect 358 3371 367 3377
rect 358 3368 364 3371
tri 364 3368 367 3371 nw
rect 474 3546 520 3558
rect 474 3512 480 3546
rect 514 3512 520 3546
rect 474 3474 520 3512
rect 474 3440 480 3474
rect 514 3440 520 3474
rect 474 3402 520 3440
rect 474 3368 480 3402
rect 514 3368 520 3402
rect 162 3330 208 3368
rect 162 3296 168 3330
rect 202 3296 208 3330
rect 162 3258 208 3296
rect 162 3224 168 3258
rect 202 3224 208 3258
rect 162 3186 208 3224
rect 162 3152 168 3186
rect 202 3152 208 3186
rect 162 3114 208 3152
rect 162 3080 168 3114
rect 202 3080 208 3114
rect 162 3042 208 3080
rect 162 3008 168 3042
rect 202 3008 208 3042
rect 162 2970 208 3008
rect 162 2936 168 2970
rect 202 2936 208 2970
rect 162 2898 208 2936
rect 162 2864 168 2898
rect 202 2864 208 2898
rect 162 2826 208 2864
rect 162 2792 168 2826
rect 202 2792 208 2826
rect 162 2754 208 2792
rect 162 2720 168 2754
rect 202 2720 208 2754
rect 162 2682 208 2720
rect 162 2648 168 2682
rect 202 2648 208 2682
rect 162 2610 208 2648
rect 162 2576 168 2610
rect 202 2576 208 2610
rect -11 2432 41 2438
rect -11 2368 41 2380
rect -176 1942 -170 1994
rect -118 1942 -102 1994
rect -50 1942 -44 1994
rect -227 1867 -181 1879
rect -227 1833 -221 1867
rect -187 1833 -181 1867
rect -227 1795 -181 1833
rect -227 1761 -221 1795
rect -187 1761 -181 1795
rect -227 1723 -181 1761
rect -227 1689 -221 1723
rect -187 1689 -181 1723
rect -227 1651 -181 1689
rect -227 1617 -221 1651
rect -187 1617 -181 1651
rect -227 1579 -181 1617
rect -227 1545 -221 1579
rect -187 1545 -181 1579
tri -230 1524 -227 1527 se
rect -227 1524 -181 1545
rect -11 1867 41 2316
rect 162 2294 208 2576
rect 318 3330 364 3368
rect 318 3296 324 3330
rect 358 3296 364 3330
rect 318 3258 364 3296
rect 318 3224 324 3258
rect 358 3224 364 3258
rect 318 3186 364 3224
rect 318 3152 324 3186
rect 358 3152 364 3186
rect 318 3114 364 3152
rect 318 3080 324 3114
rect 358 3080 364 3114
rect 318 3042 364 3080
rect 318 3008 324 3042
rect 358 3008 364 3042
rect 318 2970 364 3008
rect 318 2936 324 2970
rect 358 2936 364 2970
rect 318 2898 364 2936
rect 318 2864 324 2898
rect 358 2864 364 2898
rect 318 2826 364 2864
rect 318 2792 324 2826
rect 358 2792 364 2826
rect 318 2754 364 2792
rect 318 2720 324 2754
rect 358 2720 364 2754
rect 318 2682 364 2720
rect 318 2648 324 2682
rect 358 2648 364 2682
rect 318 2610 364 2648
rect 318 2576 324 2610
rect 358 2576 364 2610
rect 318 2564 364 2576
rect 474 3330 520 3368
rect 474 3296 480 3330
rect 514 3296 520 3330
rect 474 3258 520 3296
rect 610 3546 656 3558
rect 610 3512 616 3546
rect 650 3512 656 3546
rect 610 3474 656 3512
rect 610 3440 616 3474
rect 650 3440 656 3474
rect 610 3402 656 3440
rect 610 3368 616 3402
rect 650 3368 656 3402
rect 610 3330 656 3368
rect 610 3296 616 3330
rect 650 3296 656 3330
rect 474 3224 480 3258
rect 514 3224 520 3258
rect 474 3186 520 3224
rect 474 3152 480 3186
rect 514 3152 520 3186
tri 607 3281 610 3284 se
rect 610 3281 656 3296
rect 766 3546 812 3558
rect 766 3512 772 3546
rect 806 3512 812 3546
rect 766 3474 812 3512
rect 766 3440 772 3474
rect 806 3440 812 3474
rect 766 3402 812 3440
rect 766 3368 772 3402
rect 806 3368 812 3402
rect 919 3557 971 3563
rect 919 3493 971 3505
rect 919 3440 928 3441
rect 962 3440 971 3441
rect 919 3429 971 3440
rect 919 3371 928 3377
tri 919 3368 922 3371 ne
rect 922 3368 928 3371
rect 962 3371 971 3377
rect 962 3368 968 3371
tri 968 3368 971 3371 nw
rect 1049 3546 1095 3558
rect 1049 3512 1055 3546
rect 1089 3512 1095 3546
rect 1049 3474 1095 3512
rect 1049 3440 1055 3474
rect 1089 3440 1095 3474
rect 1049 3402 1095 3440
rect 1049 3368 1055 3402
rect 1089 3368 1095 3402
rect 766 3330 812 3368
rect 766 3296 772 3330
rect 806 3296 812 3330
tri 656 3281 659 3284 sw
rect 607 3275 659 3281
rect 607 3211 659 3223
rect 607 3153 616 3159
tri 607 3152 608 3153 ne
rect 608 3152 616 3153
rect 650 3153 659 3159
rect 650 3152 658 3153
tri 658 3152 659 3153 nw
rect 766 3258 812 3296
rect 766 3224 772 3258
rect 806 3224 812 3258
rect 766 3186 812 3224
rect 766 3152 772 3186
rect 806 3152 812 3186
rect 474 3114 520 3152
tri 608 3151 609 3152 ne
rect 609 3151 657 3152
tri 657 3151 658 3152 nw
tri 609 3150 610 3151 ne
rect 474 3080 480 3114
rect 514 3080 520 3114
rect 474 3042 520 3080
rect 474 3008 480 3042
rect 514 3008 520 3042
rect 474 2970 520 3008
rect 474 2936 480 2970
rect 514 2936 520 2970
rect 474 2898 520 2936
rect 474 2864 480 2898
rect 514 2864 520 2898
rect 474 2826 520 2864
rect 474 2792 480 2826
rect 514 2792 520 2826
rect 474 2754 520 2792
rect 474 2720 480 2754
rect 514 2720 520 2754
rect 474 2682 520 2720
rect 474 2648 480 2682
rect 514 2648 520 2682
rect 474 2610 520 2648
rect 474 2576 480 2610
rect 514 2576 520 2610
rect 391 2520 443 2528
rect 241 2503 287 2515
rect 241 2469 247 2503
rect 281 2469 287 2503
rect 241 2431 287 2469
rect 241 2397 247 2431
rect 281 2397 287 2431
rect 391 2456 443 2468
rect 391 2398 443 2404
rect 474 2410 520 2576
rect 610 3114 656 3151
tri 656 3150 657 3151 nw
rect 610 3080 616 3114
rect 650 3080 656 3114
rect 766 3114 812 3152
rect 610 3042 656 3080
rect 610 3008 616 3042
rect 650 3008 656 3042
rect 610 2970 656 3008
rect 610 2936 616 2970
rect 650 2936 656 2970
tri 763 3095 766 3098 se
rect 766 3095 772 3114
rect 763 3089 772 3095
rect 806 3095 812 3114
rect 922 3330 968 3368
rect 922 3296 928 3330
rect 962 3296 968 3330
rect 922 3258 968 3296
rect 1049 3330 1095 3368
rect 1049 3296 1055 3330
rect 1089 3296 1095 3330
rect 922 3224 928 3258
rect 962 3224 968 3258
rect 922 3186 968 3224
rect 922 3152 928 3186
rect 962 3152 968 3186
tri 1046 3281 1049 3284 se
rect 1049 3281 1095 3296
rect 1205 3546 1251 3558
rect 1205 3512 1211 3546
rect 1245 3512 1251 3546
rect 1205 3474 1251 3512
rect 1205 3440 1211 3474
rect 1245 3440 1251 3474
rect 1205 3402 1251 3440
rect 1205 3368 1211 3402
rect 1245 3368 1251 3402
rect 1406 3557 1458 3563
rect 1406 3493 1458 3505
rect 1406 3440 1415 3441
rect 1449 3440 1458 3441
rect 1406 3429 1458 3440
rect 1406 3371 1415 3377
tri 1406 3368 1409 3371 ne
rect 1409 3368 1415 3371
rect 1449 3371 1458 3377
rect 1449 3368 1455 3371
tri 1455 3368 1458 3371 nw
rect 1565 3546 1611 3558
rect 1565 3512 1571 3546
rect 1605 3512 1611 3546
rect 1565 3474 1611 3512
rect 1565 3440 1571 3474
rect 1605 3440 1611 3474
rect 1565 3402 1611 3440
rect 1565 3368 1571 3402
rect 1605 3368 1611 3402
rect 1699 3557 1751 3563
rect 2305 3558 2351 3570
rect 2305 3524 2311 3558
rect 2345 3524 2351 3558
rect 1699 3493 1708 3505
rect 1742 3493 1751 3505
rect 1699 3439 1751 3441
rect 1699 3429 1708 3439
rect 1742 3429 1751 3439
rect 1699 3371 1751 3377
tri 1699 3368 1702 3371 ne
rect 1205 3330 1251 3368
rect 1205 3296 1211 3330
rect 1245 3296 1251 3330
tri 1095 3281 1098 3284 sw
rect 1046 3275 1098 3281
rect 1046 3211 1098 3223
rect 1046 3153 1055 3159
tri 1046 3152 1047 3153 ne
rect 1047 3152 1055 3153
rect 1089 3153 1098 3159
rect 1089 3152 1097 3153
tri 1097 3152 1098 3153 nw
rect 1205 3258 1251 3296
rect 1205 3224 1211 3258
rect 1245 3224 1251 3258
rect 1205 3186 1251 3224
rect 1205 3152 1211 3186
rect 1245 3152 1251 3186
rect 922 3114 968 3152
tri 1047 3151 1048 3152 ne
rect 1048 3151 1096 3152
tri 1096 3151 1097 3152 nw
tri 1048 3150 1049 3151 ne
tri 812 3095 815 3098 sw
rect 806 3089 815 3095
rect 763 3025 772 3037
rect 806 3025 815 3037
rect 763 2970 815 2973
rect 763 2967 772 2970
tri 763 2964 766 2967 ne
rect 610 2898 656 2936
rect 610 2864 616 2898
rect 650 2864 656 2898
rect 610 2826 656 2864
rect 610 2792 616 2826
rect 650 2792 656 2826
rect 610 2754 656 2792
rect 610 2720 616 2754
rect 650 2720 656 2754
rect 610 2682 656 2720
rect 610 2648 616 2682
rect 650 2648 656 2682
rect 610 2610 656 2648
rect 610 2576 616 2610
rect 650 2576 656 2610
rect 610 2564 656 2576
rect 766 2936 772 2967
rect 806 2967 815 2970
rect 806 2936 812 2967
tri 812 2964 815 2967 nw
rect 922 3080 928 3114
rect 962 3080 968 3114
rect 922 3042 968 3080
rect 922 3008 928 3042
rect 962 3008 968 3042
rect 922 2970 968 3008
rect 766 2898 812 2936
rect 766 2864 772 2898
rect 806 2864 812 2898
rect 766 2826 812 2864
rect 766 2792 772 2826
rect 806 2792 812 2826
rect 766 2754 812 2792
rect 766 2720 772 2754
rect 806 2720 812 2754
rect 766 2682 812 2720
rect 766 2648 772 2682
rect 806 2648 812 2682
rect 766 2610 812 2648
rect 766 2576 772 2610
rect 806 2576 812 2610
rect 766 2564 812 2576
rect 922 2936 928 2970
rect 962 2936 968 2970
rect 922 2898 968 2936
rect 922 2864 928 2898
rect 962 2864 968 2898
rect 922 2826 968 2864
rect 922 2792 928 2826
rect 962 2792 968 2826
rect 922 2754 968 2792
rect 922 2720 928 2754
rect 962 2720 968 2754
rect 922 2682 968 2720
rect 922 2648 928 2682
rect 962 2648 968 2682
rect 922 2610 968 2648
rect 922 2576 928 2610
rect 962 2576 968 2610
rect 922 2564 968 2576
rect 1049 3114 1095 3151
tri 1095 3150 1096 3151 nw
rect 1049 3080 1055 3114
rect 1089 3080 1095 3114
rect 1049 3042 1095 3080
rect 1049 3008 1055 3042
rect 1089 3008 1095 3042
rect 1049 2970 1095 3008
rect 1049 2936 1055 2970
rect 1089 2936 1095 2970
rect 1049 2898 1095 2936
rect 1049 2864 1055 2898
rect 1089 2864 1095 2898
rect 1205 3114 1251 3152
rect 1205 3080 1211 3114
rect 1245 3080 1251 3114
rect 1205 3042 1251 3080
rect 1205 3008 1211 3042
rect 1245 3008 1251 3042
rect 1205 2970 1251 3008
rect 1205 2936 1211 2970
rect 1245 2936 1251 2970
rect 1205 2898 1251 2936
rect 1049 2826 1095 2864
rect 1049 2792 1055 2826
rect 1089 2792 1095 2826
rect 1049 2754 1095 2792
rect 1049 2720 1055 2754
rect 1089 2720 1095 2754
rect 1049 2682 1095 2720
rect 1049 2648 1055 2682
rect 1089 2648 1095 2682
rect 1049 2610 1095 2648
rect 1049 2576 1055 2610
rect 1089 2576 1095 2610
rect 1049 2564 1095 2576
rect 1124 2883 1176 2889
rect 1124 2819 1176 2831
tri 682 2521 689 2528 se
rect 689 2521 735 2528
tri 678 2517 682 2521 se
rect 682 2517 735 2521
tri 677 2516 678 2517 se
rect 678 2516 735 2517
tri 648 2487 677 2516 se
rect 677 2487 695 2516
rect 607 2435 613 2487
rect 665 2435 677 2487
tri 652 2419 668 2435 ne
rect 668 2419 695 2435
tri 520 2410 529 2419 sw
tri 668 2410 677 2419 ne
rect 677 2410 695 2419
rect 729 2410 735 2516
rect 474 2409 529 2410
tri 529 2409 530 2410 sw
tri 677 2409 678 2410 ne
rect 678 2409 735 2410
rect 474 2398 530 2409
tri 530 2398 541 2409 sw
tri 678 2398 689 2409 ne
rect 689 2398 735 2409
rect 845 2516 891 2528
rect 845 2482 851 2516
rect 885 2482 891 2516
rect 845 2444 891 2482
rect 845 2410 851 2444
rect 885 2410 891 2444
rect 1124 2516 1176 2767
rect 1124 2482 1134 2516
rect 1168 2482 1176 2516
rect 1124 2444 1176 2482
tri 891 2410 921 2440 sw
rect 1124 2410 1134 2444
rect 1168 2410 1176 2444
rect 845 2409 921 2410
tri 921 2409 922 2410 sw
rect 241 2385 287 2397
rect 474 2385 541 2398
tri 541 2385 554 2398 sw
rect 845 2387 922 2409
tri 922 2387 944 2409 sw
rect 474 2375 554 2385
tri 554 2375 564 2385 sw
rect 474 2365 564 2375
tri 564 2365 574 2375 sw
rect 474 2362 574 2365
tri 574 2362 577 2365 sw
tri 208 2294 239 2325 sw
rect 474 2310 480 2362
rect 532 2310 544 2362
rect 596 2310 602 2362
rect 845 2335 851 2387
rect 903 2335 915 2387
rect 967 2335 973 2387
tri 1095 2335 1124 2364 se
rect 1124 2342 1176 2410
rect 1124 2335 1165 2342
tri 1091 2331 1095 2335 se
rect 1095 2331 1165 2335
tri 1165 2331 1176 2342 nw
rect 1205 2864 1211 2898
rect 1245 2864 1251 2898
rect 1205 2826 1251 2864
rect 1205 2792 1211 2826
rect 1245 2792 1251 2826
rect 1205 2754 1251 2792
rect 1205 2720 1211 2754
rect 1245 2720 1251 2754
rect 1205 2682 1251 2720
rect 1205 2648 1211 2682
rect 1245 2648 1251 2682
rect 1205 2610 1251 2648
rect 1205 2576 1211 2610
rect 1245 2576 1251 2610
tri 1088 2328 1091 2331 se
rect 1091 2328 1162 2331
tri 1162 2328 1165 2331 nw
tri 1070 2310 1088 2328 se
rect 1088 2310 1128 2328
tri 1054 2294 1070 2310 se
rect 1070 2294 1128 2310
tri 1128 2294 1162 2328 nw
rect 162 2289 239 2294
tri 239 2289 244 2294 sw
tri 1051 2291 1054 2294 se
rect 1054 2291 1125 2294
tri 1125 2291 1128 2294 nw
tri 708 2289 710 2291 se
rect 710 2289 1123 2291
tri 1123 2289 1125 2291 nw
rect 162 2269 244 2289
tri 244 2269 264 2289 sw
tri 688 2269 708 2289 se
rect 708 2269 1103 2289
tri 1103 2269 1123 2289 nw
rect 162 2255 264 2269
tri 264 2255 278 2269 sw
tri 674 2255 688 2269 se
rect 688 2255 1073 2269
rect 162 2253 278 2255
tri 278 2253 280 2255 sw
tri 672 2253 674 2255 se
rect 674 2253 1073 2255
rect 162 2241 284 2253
rect 162 2207 244 2241
rect 278 2207 284 2241
rect 162 2169 284 2207
rect 162 2135 244 2169
rect 278 2135 284 2169
rect 162 2097 284 2135
rect 474 2241 520 2253
rect 474 2207 480 2241
rect 514 2207 520 2241
tri 654 2235 672 2253 se
rect 672 2239 1073 2253
tri 1073 2239 1103 2269 nw
rect 672 2235 728 2239
tri 728 2235 732 2239 nw
tri 636 2217 654 2235 se
rect 654 2217 710 2235
tri 710 2217 728 2235 nw
rect 474 2169 520 2207
tri 624 2205 636 2217 se
rect 636 2205 698 2217
tri 698 2205 710 2217 nw
rect 474 2135 480 2169
rect 514 2135 520 2169
tri 617 2198 624 2205 se
rect 624 2198 691 2205
tri 691 2198 698 2205 nw
rect 617 2181 674 2198
tri 674 2181 691 2198 nw
rect 474 2129 520 2135
tri 520 2129 531 2140 sw
tri 468 2120 474 2126 se
rect 474 2120 531 2129
tri 531 2120 540 2129 sw
tri 445 2097 468 2120 se
rect 468 2097 540 2120
rect 162 2063 244 2097
rect 278 2063 284 2097
rect 162 2051 284 2063
tri 440 2092 445 2097 se
rect 445 2092 480 2097
rect 514 2092 540 2097
tri 540 2092 568 2120 sw
rect 440 2040 446 2092
rect 498 2040 510 2063
rect 562 2040 568 2092
rect 617 2026 669 2181
tri 669 2176 674 2181 nw
rect 765 2077 771 2129
rect 823 2077 837 2129
rect 889 2120 904 2129
rect 956 2120 971 2129
rect 1023 2120 1038 2129
rect 896 2086 904 2120
rect 1023 2086 1030 2120
rect 889 2077 904 2086
rect 956 2077 971 2086
rect 1023 2077 1038 2086
rect 1090 2077 1105 2129
rect 1157 2077 1163 2129
tri 1202 2030 1205 2033 se
rect 1205 2030 1251 2576
rect 1409 3330 1455 3368
rect 1409 3296 1415 3330
rect 1449 3296 1455 3330
rect 1409 3258 1455 3296
rect 1409 3224 1415 3258
rect 1449 3224 1455 3258
rect 1409 3186 1455 3224
rect 1409 3152 1415 3186
rect 1449 3152 1455 3186
rect 1409 3114 1455 3152
rect 1409 3080 1415 3114
rect 1449 3080 1455 3114
rect 1409 3042 1455 3080
rect 1409 3008 1415 3042
rect 1449 3008 1455 3042
rect 1409 2970 1455 3008
rect 1409 2936 1415 2970
rect 1449 2936 1455 2970
rect 1409 2898 1455 2936
rect 1409 2864 1415 2898
rect 1449 2864 1455 2898
rect 1409 2826 1455 2864
rect 1409 2792 1415 2826
rect 1449 2792 1455 2826
rect 1409 2754 1455 2792
rect 1409 2720 1415 2754
rect 1449 2720 1455 2754
rect 1409 2682 1455 2720
rect 1409 2648 1415 2682
rect 1449 2648 1455 2682
rect 1409 2610 1455 2648
rect 1409 2576 1415 2610
rect 1449 2576 1455 2610
rect 1409 2564 1455 2576
rect 1565 3330 1611 3368
rect 1565 3296 1571 3330
rect 1605 3296 1611 3330
rect 1565 3258 1611 3296
rect 1565 3224 1571 3258
rect 1605 3224 1611 3258
rect 1565 3186 1611 3224
rect 1565 3152 1571 3186
rect 1605 3152 1611 3186
rect 1565 3114 1611 3152
rect 1565 3080 1571 3114
rect 1605 3080 1611 3114
rect 1565 3042 1611 3080
rect 1565 3008 1571 3042
rect 1605 3008 1611 3042
rect 1565 2970 1611 3008
rect 1565 2936 1571 2970
rect 1605 2936 1611 2970
rect 1565 2898 1611 2936
rect 1565 2864 1571 2898
rect 1605 2864 1611 2898
rect 1565 2826 1611 2864
rect 1565 2792 1571 2826
rect 1605 2792 1611 2826
rect 1565 2754 1611 2792
rect 1565 2720 1571 2754
rect 1605 2720 1611 2754
rect 1565 2682 1611 2720
rect 1565 2648 1571 2682
rect 1605 2648 1611 2682
rect 1565 2610 1611 2648
rect 1565 2576 1571 2610
rect 1605 2576 1611 2610
tri 1481 2521 1488 2528 se
rect 1488 2521 1534 2528
tri 1477 2517 1481 2521 se
rect 1481 2517 1534 2521
tri 1476 2516 1477 2517 se
rect 1477 2516 1534 2517
tri 1473 2513 1476 2516 se
rect 1476 2513 1494 2516
rect 1406 2461 1412 2513
rect 1464 2461 1476 2513
rect 1528 2461 1534 2516
tri 1450 2447 1464 2461 ne
rect 1464 2447 1534 2461
tri 1464 2446 1465 2447 ne
rect 1465 2446 1534 2447
tri 1465 2444 1467 2446 ne
rect 1467 2444 1534 2446
tri 1467 2423 1488 2444 ne
rect 1488 2410 1494 2444
rect 1528 2410 1534 2444
rect 1293 2269 1453 2281
rect 1293 2235 1299 2269
rect 1333 2235 1413 2269
rect 1447 2235 1453 2269
rect 1293 2181 1453 2235
rect 1293 2147 1299 2181
rect 1333 2147 1413 2181
rect 1447 2147 1453 2181
rect 1293 2127 1453 2147
rect 1293 2060 1299 2127
rect 1351 2075 1395 2127
rect 1333 2060 1413 2075
rect 1447 2060 1453 2127
rect 1293 2048 1453 2060
rect 1488 2113 1534 2410
rect 1565 2205 1611 2576
rect 1702 3367 1748 3371
tri 1748 3368 1751 3371 nw
rect 1858 3511 1904 3523
rect 1858 3477 1864 3511
rect 1898 3477 1904 3511
rect 1858 3439 1904 3477
rect 1858 3405 1864 3439
rect 1898 3405 1904 3439
rect 1702 3333 1708 3367
rect 1742 3333 1748 3367
rect 1702 3295 1748 3333
rect 1702 3261 1708 3295
rect 1742 3261 1748 3295
rect 1702 3223 1748 3261
rect 1702 3189 1708 3223
rect 1742 3189 1748 3223
rect 1702 3151 1748 3189
rect 1702 3117 1708 3151
rect 1742 3117 1748 3151
rect 1702 3079 1748 3117
rect 1702 3045 1708 3079
rect 1742 3045 1748 3079
rect 1702 3007 1748 3045
rect 1702 2973 1708 3007
rect 1742 2973 1748 3007
rect 1702 2935 1748 2973
rect 1702 2901 1708 2935
rect 1742 2901 1748 2935
rect 1702 2863 1748 2901
rect 1702 2829 1708 2863
rect 1742 2829 1748 2863
rect 1702 2791 1748 2829
rect 1702 2757 1708 2791
rect 1742 2757 1748 2791
rect 1702 2719 1748 2757
rect 1702 2685 1708 2719
rect 1742 2685 1748 2719
rect 1702 2647 1748 2685
rect 1702 2613 1708 2647
rect 1742 2613 1748 2647
rect 1702 2575 1748 2613
rect 1702 2541 1708 2575
rect 1742 2541 1748 2575
rect 1702 2529 1748 2541
rect 1858 3367 1904 3405
rect 1858 3333 1864 3367
rect 1898 3333 1904 3367
rect 1858 3295 1904 3333
rect 1858 3261 1864 3295
rect 1898 3261 1904 3295
rect 1858 3223 1904 3261
rect 1858 3189 1864 3223
rect 1898 3189 1904 3223
rect 1858 3151 1904 3189
rect 1858 3117 1864 3151
rect 1898 3117 1904 3151
rect 1858 3079 1904 3117
rect 1858 3045 1864 3079
rect 1898 3045 1904 3079
rect 1858 3007 1904 3045
rect 1858 2973 1864 3007
rect 1898 2973 1904 3007
rect 1858 2935 1904 2973
rect 1858 2901 1864 2935
rect 1898 2901 1904 2935
rect 1858 2863 1904 2901
rect 1858 2829 1864 2863
rect 1898 2829 1904 2863
rect 1858 2791 1904 2829
rect 1858 2757 1864 2791
rect 1898 2757 1904 2791
rect 1858 2719 1904 2757
rect 2014 3511 2060 3523
rect 2014 3477 2020 3511
rect 2054 3477 2060 3511
rect 2014 3439 2060 3477
rect 2014 3405 2020 3439
rect 2054 3405 2060 3439
rect 2014 3367 2060 3405
rect 2014 3333 2020 3367
rect 2054 3333 2060 3367
rect 2014 3295 2060 3333
rect 2014 3261 2020 3295
rect 2054 3261 2060 3295
rect 2014 3223 2060 3261
rect 2014 3189 2020 3223
rect 2054 3189 2060 3223
rect 2014 3151 2060 3189
rect 2014 3117 2020 3151
rect 2054 3117 2060 3151
rect 2014 3079 2060 3117
rect 2014 3045 2020 3079
rect 2054 3045 2060 3079
rect 2014 3007 2060 3045
rect 2014 2973 2020 3007
rect 2054 2973 2060 3007
rect 2014 2935 2060 2973
rect 2014 2901 2020 2935
rect 2054 2901 2060 2935
rect 2014 2863 2060 2901
rect 2014 2829 2020 2863
rect 2054 2829 2060 2863
rect 2014 2791 2060 2829
rect 2014 2757 2020 2791
rect 2054 2757 2060 2791
rect 1858 2685 1864 2719
rect 1898 2685 1904 2719
rect 1858 2647 1904 2685
rect 1858 2613 1864 2647
rect 1898 2613 1904 2647
rect 1858 2575 1904 2613
rect 1858 2541 1864 2575
rect 1898 2541 1904 2575
rect 1764 2481 1810 2493
rect 1764 2447 1770 2481
rect 1804 2447 1810 2481
tri 1750 2409 1764 2423 se
rect 1764 2409 1810 2447
tri 1728 2387 1750 2409 se
rect 1750 2387 1770 2409
rect 1682 2335 1688 2387
rect 1740 2335 1752 2387
rect 1804 2335 1810 2409
tri 1855 2331 1858 2334 se
rect 1858 2331 1904 2541
rect 1933 2744 1985 2750
rect 1933 2680 1985 2692
rect 1933 2481 1985 2628
rect 1933 2447 1943 2481
rect 1977 2447 1985 2481
rect 1933 2409 1985 2447
rect 1933 2375 1943 2409
rect 1977 2375 1985 2409
rect 1933 2363 1985 2375
rect 2014 2719 2060 2757
rect 2014 2685 2020 2719
rect 2054 2685 2060 2719
rect 2014 2647 2060 2685
rect 2014 2613 2020 2647
rect 2054 2613 2060 2647
rect 2014 2575 2060 2613
rect 2014 2541 2020 2575
rect 2054 2541 2060 2575
tri 1852 2328 1855 2331 se
rect 1855 2328 1904 2331
tri 1831 2307 1852 2328 se
rect 1852 2307 1904 2328
rect 1776 2255 1782 2307
rect 1834 2255 1846 2307
rect 1898 2255 1904 2307
tri 2003 2255 2014 2266 se
rect 2014 2255 2060 2541
rect 2170 3511 2216 3523
rect 2170 3477 2176 3511
rect 2210 3477 2216 3511
rect 2170 3439 2216 3477
rect 2170 3405 2176 3439
rect 2210 3405 2216 3439
rect 2170 3367 2216 3405
rect 2170 3333 2176 3367
rect 2210 3333 2216 3367
rect 2170 3295 2216 3333
rect 2170 3261 2176 3295
rect 2210 3261 2216 3295
rect 2170 3223 2216 3261
rect 2170 3189 2176 3223
rect 2210 3189 2216 3223
rect 2170 3151 2216 3189
rect 2170 3117 2176 3151
rect 2210 3117 2216 3151
rect 2170 3079 2216 3117
rect 2170 3045 2176 3079
rect 2210 3045 2216 3079
rect 2305 3486 2351 3524
rect 2305 3452 2311 3486
rect 2345 3452 2351 3486
rect 2305 3372 2351 3452
rect 2458 3562 2510 3570
rect 2458 3498 2510 3510
rect 2458 3440 2510 3446
rect 2617 3558 2663 3570
rect 2617 3524 2623 3558
rect 2657 3524 2663 3558
rect 2617 3486 2663 3524
rect 2617 3452 2623 3486
rect 2657 3452 2663 3486
tri 2351 3372 2366 3387 sw
rect 2305 3371 2366 3372
tri 2366 3371 2367 3372 sw
rect 2305 3354 2367 3371
tri 2367 3354 2384 3371 sw
rect 2305 3353 2384 3354
tri 2384 3353 2385 3354 sw
rect 2305 3333 2385 3353
tri 2385 3333 2405 3353 sw
rect 2305 3323 2405 3333
tri 2405 3323 2415 3333 sw
rect 2305 3279 2586 3323
rect 2305 3278 2395 3279
tri 2395 3278 2396 3279 nw
tri 2505 3278 2506 3279 ne
rect 2506 3278 2586 3279
rect 2305 3277 2394 3278
tri 2394 3277 2395 3278 nw
tri 2506 3277 2507 3278 ne
rect 2507 3277 2586 3278
rect 2305 3261 2378 3277
tri 2378 3261 2394 3277 nw
tri 2507 3261 2523 3277 ne
rect 2523 3261 2586 3277
rect 2305 3250 2367 3261
tri 2367 3250 2378 3261 nw
tri 2523 3250 2534 3261 ne
rect 2534 3250 2586 3261
rect 2305 3238 2355 3250
tri 2355 3238 2367 3250 nw
tri 2534 3244 2540 3250 ne
rect 2540 3238 2586 3250
tri 2304 3050 2305 3051 se
rect 2305 3050 2351 3238
tri 2351 3234 2355 3238 nw
rect 2540 3204 2546 3238
rect 2580 3204 2586 3238
rect 2540 3166 2586 3204
rect 2540 3132 2546 3166
rect 2580 3132 2586 3166
tri 2303 3049 2304 3050 se
rect 2304 3049 2351 3050
rect 2170 3007 2216 3045
rect 2170 2973 2176 3007
rect 2210 2973 2216 3007
rect 2170 2935 2216 2973
rect 2170 2901 2176 2935
rect 2210 2901 2216 2935
tri 2299 3045 2303 3049 se
rect 2303 3045 2351 3049
rect 2299 3039 2351 3045
rect 2299 2975 2351 2987
rect 2388 3104 2434 3121
rect 2540 3120 2586 3132
rect 2388 3070 2394 3104
rect 2428 3083 2434 3104
tri 2434 3083 2436 3085 sw
rect 2428 3076 2436 3083
tri 2436 3076 2443 3083 sw
rect 2428 3070 2443 3076
rect 2388 3067 2443 3070
tri 2443 3067 2452 3076 sw
tri 2608 3067 2617 3076 se
rect 2617 3067 2663 3452
rect 2748 3561 2800 3567
rect 3031 3561 3083 3567
rect 3343 3561 3395 3567
rect 2748 3496 2800 3509
rect 2748 3443 2757 3444
rect 2791 3443 2800 3444
rect 2748 3430 2800 3443
rect 2748 3372 2757 3378
tri 2748 3371 2749 3372 ne
rect 2749 3371 2757 3372
rect 2791 3372 2800 3378
rect 2791 3371 2799 3372
tri 2799 3371 2800 3372 nw
rect 2907 3549 2953 3561
rect 2907 3515 2913 3549
rect 2947 3515 2953 3549
rect 2907 3477 2953 3515
rect 2907 3443 2913 3477
rect 2947 3443 2953 3477
rect 2907 3405 2953 3443
rect 2907 3371 2913 3405
rect 2947 3371 2953 3405
rect 3031 3496 3083 3509
rect 3031 3443 3040 3444
rect 3074 3443 3083 3444
rect 3031 3430 3083 3443
rect 3031 3372 3040 3378
tri 3031 3371 3032 3372 ne
rect 3032 3371 3040 3372
rect 3074 3372 3083 3378
rect 3074 3371 3082 3372
tri 3082 3371 3083 3372 nw
rect 3190 3549 3236 3561
rect 3190 3515 3196 3549
rect 3230 3515 3236 3549
rect 3190 3477 3236 3515
rect 3190 3443 3196 3477
rect 3230 3443 3236 3477
rect 3190 3405 3236 3443
rect 3190 3371 3196 3405
rect 3230 3371 3236 3405
rect 3343 3496 3395 3509
rect 3343 3443 3352 3444
rect 3386 3443 3395 3444
rect 3343 3430 3395 3443
rect 3343 3372 3352 3378
tri 3343 3371 3344 3372 ne
rect 3344 3371 3352 3372
rect 3386 3372 3395 3378
rect 3386 3371 3394 3372
tri 3394 3371 3395 3372 nw
rect 3502 3549 3548 3561
rect 3502 3515 3508 3549
rect 3542 3515 3548 3549
rect 3502 3477 3548 3515
rect 3502 3443 3508 3477
rect 3542 3443 3548 3477
rect 3502 3405 3548 3443
rect 3932 3540 3978 3582
rect 3932 3506 3938 3540
rect 3972 3506 3978 3540
rect 3932 3464 3978 3506
rect 3932 3430 3938 3464
rect 3972 3430 3978 3464
rect 3502 3371 3508 3405
rect 3542 3371 3548 3405
tri 3912 3395 3932 3415 se
rect 3932 3395 3978 3430
tri 3905 3388 3912 3395 se
rect 3912 3388 3978 3395
tri 2749 3369 2751 3371 ne
rect 2388 3050 2452 3067
tri 2452 3050 2469 3067 sw
tri 2591 3050 2608 3067 se
rect 2608 3050 2663 3067
rect 2388 3049 2469 3050
tri 2469 3049 2470 3050 sw
tri 2590 3049 2591 3050 se
rect 2591 3049 2663 3050
rect 2388 3045 2470 3049
tri 2470 3045 2474 3049 sw
tri 2586 3045 2590 3049 se
rect 2590 3045 2663 3049
rect 2388 3032 2474 3045
rect 2388 2998 2394 3032
rect 2428 3027 2474 3032
tri 2474 3027 2492 3045 sw
tri 2568 3027 2586 3045 se
rect 2586 3027 2663 3045
rect 2428 2998 2663 3027
rect 2751 3333 2797 3371
tri 2797 3369 2799 3371 nw
rect 2751 3299 2757 3333
rect 2791 3299 2797 3333
rect 2751 3261 2797 3299
rect 2751 3227 2757 3261
rect 2791 3227 2797 3261
rect 2751 3189 2797 3227
rect 2751 3155 2757 3189
rect 2791 3155 2797 3189
rect 2751 3117 2797 3155
rect 2751 3083 2757 3117
rect 2791 3083 2797 3117
rect 2751 3045 2797 3083
rect 2751 3011 2757 3045
rect 2791 3011 2797 3045
rect 2751 2999 2797 3011
rect 2907 3333 2953 3371
tri 3032 3369 3034 3371 ne
rect 2907 3299 2913 3333
rect 2947 3299 2953 3333
rect 2907 3261 2953 3299
rect 2907 3227 2913 3261
rect 2947 3227 2953 3261
rect 2907 3189 2953 3227
rect 2907 3155 2913 3189
rect 2947 3155 2953 3189
rect 2907 3117 2953 3155
rect 2907 3083 2913 3117
rect 2947 3083 2953 3117
rect 2907 3045 2953 3083
rect 2907 3011 2913 3045
rect 2947 3011 2953 3045
rect 2388 2981 2663 2998
tri 2565 2974 2572 2981 ne
rect 2572 2974 2663 2981
tri 2572 2973 2573 2974 ne
rect 2573 2973 2663 2974
tri 2573 2969 2577 2973 ne
rect 2577 2969 2663 2973
tri 2577 2939 2607 2969 ne
rect 2607 2939 2663 2969
tri 2607 2932 2614 2939 ne
rect 2614 2932 2663 2939
tri 2614 2929 2617 2932 ne
rect 2299 2917 2351 2923
tri 2299 2911 2305 2917 ne
rect 2170 2863 2216 2901
rect 2170 2829 2176 2863
rect 2210 2829 2216 2863
rect 2170 2791 2216 2829
rect 2170 2757 2176 2791
rect 2210 2757 2216 2791
rect 2170 2719 2216 2757
rect 2170 2685 2176 2719
rect 2210 2685 2216 2719
rect 2170 2647 2216 2685
rect 2170 2613 2176 2647
rect 2210 2635 2216 2647
tri 2216 2635 2223 2642 sw
rect 2305 2635 2351 2917
tri 2351 2635 2371 2655 sw
rect 2210 2630 2223 2635
tri 2223 2630 2228 2635 sw
tri 2305 2630 2310 2635 ne
rect 2310 2630 2371 2635
tri 2371 2630 2376 2635 sw
rect 2210 2614 2228 2630
tri 2228 2614 2244 2630 sw
tri 2310 2620 2320 2630 ne
rect 2320 2620 2376 2630
tri 2376 2620 2386 2630 sw
tri 2320 2614 2326 2620 ne
rect 2326 2614 2386 2620
tri 2386 2614 2392 2620 sw
rect 2210 2613 2244 2614
rect 2170 2590 2244 2613
tri 2244 2590 2268 2614 sw
tri 2326 2590 2350 2614 ne
rect 2350 2590 2392 2614
tri 2392 2590 2416 2614 sw
rect 2170 2580 2268 2590
tri 2268 2580 2278 2590 sw
tri 2350 2589 2351 2590 ne
rect 2351 2589 2416 2590
tri 2351 2580 2360 2589 ne
rect 2360 2580 2416 2589
tri 2416 2580 2426 2590 sw
rect 2170 2575 2278 2580
rect 2170 2541 2176 2575
rect 2210 2564 2278 2575
tri 2278 2564 2294 2580 sw
tri 2360 2564 2376 2580 ne
rect 2376 2564 2426 2580
tri 2426 2564 2442 2580 sw
rect 2210 2559 2294 2564
tri 2294 2559 2299 2564 sw
tri 2376 2559 2381 2564 ne
rect 2381 2559 2442 2564
tri 2442 2559 2447 2564 sw
rect 2210 2555 2299 2559
tri 2299 2555 2303 2559 sw
tri 2381 2555 2385 2559 ne
rect 2385 2555 2447 2559
tri 2447 2555 2451 2559 sw
rect 2210 2541 2303 2555
rect 2170 2529 2303 2541
tri 2303 2529 2329 2555 sw
tri 2385 2554 2386 2555 ne
rect 2386 2554 2451 2555
tri 2451 2554 2452 2555 sw
tri 2386 2529 2411 2554 ne
rect 2411 2529 2452 2554
tri 2452 2529 2477 2554 sw
tri 2255 2521 2263 2529 ne
rect 2263 2521 2329 2529
tri 2329 2521 2337 2529 sw
tri 2411 2521 2419 2529 ne
rect 2419 2521 2477 2529
tri 2477 2521 2485 2529 sw
tri 2263 2517 2267 2521 ne
rect 2267 2517 2337 2521
tri 2337 2517 2341 2521 sw
tri 2419 2517 2423 2521 ne
rect 2423 2517 2485 2521
tri 2485 2517 2489 2521 sw
tri 2267 2516 2268 2517 ne
rect 2268 2516 2341 2517
tri 2341 2516 2342 2517 sw
tri 2423 2516 2424 2517 ne
rect 2424 2516 2489 2517
tri 2489 2516 2490 2517 sw
tri 2268 2493 2291 2516 ne
rect 2291 2493 2342 2516
tri 2342 2493 2365 2516 sw
tri 2424 2493 2447 2516 ne
rect 2447 2493 2490 2516
tri 2490 2493 2513 2516 sw
rect 2093 2491 2215 2493
tri 2215 2491 2217 2493 sw
tri 2291 2491 2293 2493 ne
rect 2293 2491 2365 2493
tri 2365 2491 2367 2493 sw
tri 2447 2491 2449 2493 ne
rect 2449 2491 2513 2493
tri 2513 2491 2515 2493 sw
rect 2093 2487 2217 2491
tri 2217 2487 2221 2491 sw
tri 2293 2487 2297 2491 ne
rect 2297 2487 2367 2491
tri 2367 2487 2371 2491 sw
tri 2449 2488 2452 2491 ne
rect 2452 2488 2515 2491
tri 2515 2488 2518 2491 sw
tri 2452 2487 2453 2488 ne
rect 2453 2487 2518 2488
tri 2518 2487 2519 2488 sw
rect 2093 2435 2099 2487
rect 2151 2435 2163 2487
rect 2215 2483 2221 2487
tri 2221 2483 2225 2487 sw
tri 2297 2483 2301 2487 ne
rect 2301 2483 2371 2487
tri 2371 2483 2375 2487 sw
tri 2453 2483 2457 2487 ne
rect 2457 2483 2519 2487
tri 2519 2483 2523 2487 sw
rect 2215 2481 2225 2483
tri 2225 2481 2227 2483 sw
tri 2301 2481 2303 2483 ne
rect 2303 2481 2375 2483
tri 2375 2481 2377 2483 sw
tri 2457 2481 2459 2483 ne
rect 2459 2481 2523 2483
tri 2523 2481 2525 2483 sw
rect 2215 2480 2227 2481
tri 2227 2480 2228 2481 sw
tri 2303 2480 2304 2481 ne
rect 2304 2480 2377 2481
tri 2377 2480 2378 2481 sw
tri 2459 2480 2460 2481 ne
rect 2460 2480 2525 2481
tri 2525 2480 2526 2481 sw
rect 2215 2446 2228 2480
tri 2228 2446 2262 2480 sw
tri 2304 2446 2338 2480 ne
rect 2338 2446 2378 2480
tri 2378 2446 2412 2480 sw
tri 2460 2446 2494 2480 ne
rect 2494 2446 2526 2480
tri 2526 2446 2560 2480 sw
rect 2617 2449 2663 2932
rect 2734 2917 2740 2969
rect 2792 2917 2804 2969
rect 2856 2917 2862 2969
tri 2734 2898 2753 2917 ne
rect 2753 2898 2862 2917
tri 2753 2897 2754 2898 ne
rect 2754 2897 2862 2898
tri 2754 2894 2757 2897 ne
rect 2757 2894 2862 2897
tri 2757 2885 2766 2894 ne
rect 2766 2885 2862 2894
tri 2766 2873 2778 2885 ne
rect 2778 2873 2862 2885
tri 2778 2839 2812 2873 ne
rect 2812 2839 2822 2873
rect 2856 2839 2862 2873
tri 2812 2835 2816 2839 ne
rect 2816 2801 2862 2839
rect 2816 2767 2822 2801
rect 2856 2767 2862 2801
tri 2617 2446 2620 2449 ne
rect 2620 2446 2663 2449
tri 2663 2446 2686 2469 sw
rect 2816 2447 2862 2767
rect 2907 2932 2953 3011
rect 3034 3333 3080 3371
tri 3080 3369 3082 3371 nw
rect 3034 3299 3040 3333
rect 3074 3299 3080 3333
rect 3034 3261 3080 3299
rect 3034 3227 3040 3261
rect 3074 3227 3080 3261
rect 3190 3333 3236 3371
tri 3344 3369 3346 3371 ne
rect 3190 3299 3196 3333
rect 3230 3299 3236 3333
rect 3190 3261 3236 3299
rect 3034 3189 3080 3227
rect 3034 3155 3040 3189
rect 3074 3155 3080 3189
rect 3034 3117 3080 3155
rect 3034 3083 3040 3117
rect 3074 3083 3080 3117
tri 3187 3234 3190 3237 se
rect 3190 3234 3196 3261
rect 3187 3228 3196 3234
rect 3230 3236 3236 3261
rect 3346 3333 3392 3371
tri 3392 3369 3394 3371 nw
rect 3346 3299 3352 3333
rect 3386 3299 3392 3333
rect 3346 3261 3392 3299
tri 3236 3236 3237 3237 sw
rect 3230 3234 3237 3236
tri 3237 3234 3239 3236 sw
rect 3230 3228 3239 3234
rect 3187 3164 3196 3176
rect 3230 3164 3239 3176
rect 3187 3106 3196 3112
tri 3187 3103 3190 3106 ne
rect 3034 3045 3080 3083
rect 3034 3011 3040 3045
rect 3074 3011 3080 3045
rect 3034 2999 3080 3011
rect 3190 3083 3196 3106
rect 3230 3106 3239 3112
rect 3230 3104 3237 3106
tri 3237 3104 3239 3106 nw
rect 3346 3227 3352 3261
rect 3386 3227 3392 3261
rect 3502 3333 3548 3371
tri 3886 3369 3905 3388 se
rect 3905 3369 3938 3388
tri 3884 3367 3886 3369 se
rect 3886 3367 3938 3369
tri 3657 3354 3670 3367 se
rect 3670 3354 3938 3367
rect 3972 3354 3978 3388
tri 3656 3353 3657 3354 se
rect 3657 3353 3978 3354
rect 3502 3299 3508 3333
rect 3542 3299 3548 3333
tri 3622 3319 3656 3353 se
rect 3656 3319 3978 3353
tri 3615 3312 3622 3319 se
rect 3622 3312 3978 3319
rect 3502 3261 3548 3299
rect 3346 3189 3392 3227
rect 3346 3155 3352 3189
rect 3386 3155 3392 3189
rect 3346 3117 3392 3155
rect 3230 3083 3236 3104
tri 3236 3103 3237 3104 nw
rect 3190 3045 3236 3083
rect 3190 3011 3196 3045
rect 3230 3011 3236 3045
rect 3190 2999 3236 3011
rect 3346 3083 3352 3117
rect 3386 3083 3392 3117
tri 3500 3234 3502 3236 se
rect 3502 3234 3508 3261
rect 3500 3228 3508 3234
rect 3542 3236 3548 3261
tri 3586 3283 3615 3312 se
rect 3615 3283 3938 3312
rect 3586 3279 3938 3283
rect 3586 3278 3707 3279
tri 3707 3278 3708 3279 nw
tri 3876 3278 3877 3279 ne
rect 3877 3278 3938 3279
rect 3972 3278 3978 3312
rect 3586 3277 3706 3278
tri 3706 3277 3707 3278 nw
tri 3877 3277 3878 3278 ne
rect 3878 3277 3978 3278
tri 3548 3236 3550 3238 sw
rect 3542 3234 3550 3236
tri 3550 3234 3552 3236 sw
rect 3542 3228 3552 3234
rect 3500 3164 3508 3176
rect 3542 3164 3552 3176
rect 3500 3106 3508 3112
tri 3500 3104 3502 3106 ne
rect 3346 3045 3392 3083
rect 3346 3011 3352 3045
rect 3386 3011 3392 3045
rect 3346 2999 3392 3011
rect 3502 3083 3508 3106
rect 3542 3106 3552 3112
rect 3542 3104 3550 3106
tri 3550 3104 3552 3106 nw
rect 3542 3083 3548 3104
tri 3548 3102 3550 3104 nw
rect 3502 3045 3548 3083
rect 3502 3011 3508 3045
rect 3542 3011 3548 3045
rect 3502 2999 3548 3011
tri 2953 2932 2956 2935 sw
rect 2907 2900 2956 2932
tri 2956 2900 2988 2932 sw
rect 2907 2894 3467 2900
rect 2907 2860 3119 2894
rect 3153 2860 3195 2894
rect 3229 2860 3271 2894
rect 3305 2860 3346 2894
rect 3380 2860 3421 2894
rect 3455 2860 3467 2894
rect 2907 2854 3467 2860
rect 2907 2822 2957 2854
tri 2957 2822 2989 2854 nw
tri 3561 2822 3586 2847 se
rect 3586 2822 3675 3277
tri 3675 3246 3706 3277 nw
tri 3878 3246 3909 3277 ne
rect 3909 3246 3978 3277
tri 3909 3243 3912 3246 ne
rect 3912 3243 3978 3246
rect 4119 3653 4568 3659
rect 4119 3619 4207 3653
rect 4241 3619 4290 3653
rect 4324 3619 4373 3653
rect 4407 3619 4456 3653
rect 4490 3619 4568 3653
rect 4119 3613 4568 3619
rect 4119 3603 4301 3613
tri 4301 3603 4311 3613 nw
rect 4119 3581 4284 3603
tri 4284 3586 4301 3603 nw
rect 4119 3547 4125 3581
rect 4159 3549 4284 3581
rect 4522 3579 4568 3613
rect 4159 3547 4244 3549
rect 4119 3515 4244 3547
rect 4278 3515 4284 3549
rect 4119 3505 4284 3515
rect 4119 3471 4125 3505
rect 4159 3477 4284 3505
rect 4159 3471 4244 3477
rect 4119 3443 4244 3471
rect 4278 3443 4284 3477
rect 4119 3429 4284 3443
rect 4119 3395 4125 3429
rect 4159 3405 4284 3429
rect 4159 3395 4244 3405
rect 4119 3371 4244 3395
rect 4278 3371 4284 3405
rect 4119 3353 4284 3371
rect 4119 3319 4125 3353
rect 4159 3333 4284 3353
rect 4159 3319 4244 3333
rect 4119 3299 4244 3319
rect 4278 3299 4284 3333
rect 4119 3277 4284 3299
rect 4119 3243 4125 3277
rect 4159 3261 4284 3277
rect 4159 3243 4244 3261
tri 3912 3238 3917 3243 ne
rect 3917 3238 3981 3243
tri 3917 3236 3919 3238 ne
rect 3919 3237 3981 3238
rect 3919 3236 3929 3237
tri 3919 3226 3929 3236 ne
rect 3929 3160 3981 3185
rect 3929 3126 3938 3160
rect 3972 3126 3981 3160
rect 3929 3125 3981 3126
rect 3929 3067 3938 3073
rect 2907 2821 2956 2822
tri 2956 2821 2957 2822 nw
tri 3560 2821 3561 2822 se
rect 3561 2821 3675 2822
rect 2907 2483 2953 2821
tri 2953 2818 2956 2821 nw
tri 3557 2818 3560 2821 se
rect 3560 2818 3675 2821
tri 3526 2787 3557 2818 se
rect 3557 2787 3675 2818
tri 3519 2780 3526 2787 se
rect 3526 2780 3675 2787
tri 3485 2746 3519 2780 se
rect 3519 2746 3675 2780
tri 3484 2745 3485 2746 se
rect 3485 2745 3675 2746
tri 3455 2716 3484 2745 se
rect 3484 2716 3675 2745
rect 3019 2710 3675 2716
rect 3019 2676 3031 2710
rect 3065 2676 3110 2710
rect 3144 2676 3190 2710
rect 3224 2676 3270 2710
rect 3304 2676 3350 2710
rect 3384 2676 3430 2710
rect 3464 2676 3510 2710
rect 3544 2676 3590 2710
rect 3624 2676 3675 2710
rect 3019 2614 3675 2676
rect 3019 2580 3031 2614
rect 3065 2580 3110 2614
rect 3144 2580 3190 2614
rect 3224 2580 3270 2614
rect 3304 2580 3350 2614
rect 3384 2580 3430 2614
rect 3464 2580 3510 2614
rect 3544 2580 3590 2614
rect 3624 2580 3675 2614
rect 3019 2574 3675 2580
rect 3932 3050 3938 3067
rect 3972 3067 3981 3073
rect 4119 3227 4244 3243
rect 4278 3227 4284 3261
rect 4119 3201 4284 3227
rect 4119 3167 4125 3201
rect 4159 3189 4284 3201
rect 4159 3167 4244 3189
rect 4119 3155 4244 3167
rect 4278 3155 4284 3189
rect 4119 3125 4284 3155
rect 4119 3091 4125 3125
rect 4159 3117 4284 3125
rect 4159 3091 4244 3117
rect 4119 3083 4244 3091
rect 4278 3083 4284 3117
rect 3972 3050 3978 3067
rect 3932 3008 3978 3050
rect 3932 2974 3938 3008
rect 3972 2974 3978 3008
rect 3932 2932 3978 2974
rect 3932 2898 3938 2932
rect 3972 2898 3978 2932
rect 3932 2856 3978 2898
rect 3932 2822 3938 2856
rect 3972 2822 3978 2856
rect 3932 2780 3978 2822
rect 3932 2746 3938 2780
rect 3972 2746 3978 2780
rect 3932 2705 3978 2746
rect 3932 2671 3938 2705
rect 3972 2671 3978 2705
rect 3932 2630 3978 2671
rect 3932 2596 3938 2630
rect 3972 2596 3978 2630
rect 3932 2555 3978 2596
rect 3932 2521 3938 2555
rect 3972 2521 3978 2555
tri 2953 2483 2957 2487 sw
rect 2907 2481 2957 2483
tri 2957 2481 2959 2483 sw
rect 2907 2480 2959 2481
tri 2959 2480 2960 2481 sw
rect 3932 2480 3978 2521
rect 2907 2467 2960 2480
tri 2960 2467 2973 2480 sw
tri 2816 2446 2817 2447 ne
rect 2817 2446 2862 2447
tri 2862 2446 2883 2467 sw
tri 2907 2458 2916 2467 ne
rect 2916 2458 2973 2467
tri 2973 2458 2982 2467 sw
tri 2916 2454 2920 2458 ne
rect 2920 2454 3506 2458
tri 3506 2454 3510 2458 sw
tri 2920 2446 2928 2454 ne
rect 2928 2446 3510 2454
tri 3510 2446 3518 2454 sw
rect 3932 2446 3938 2480
rect 3972 2446 3978 2480
rect 2215 2442 2262 2446
tri 2262 2442 2266 2446 sw
tri 2338 2442 2342 2446 ne
rect 2342 2444 2412 2446
tri 2412 2444 2414 2446 sw
tri 2494 2444 2496 2446 ne
rect 2496 2444 2560 2446
tri 2560 2444 2562 2446 sw
tri 2620 2444 2622 2446 ne
rect 2622 2444 2686 2446
tri 2686 2444 2688 2446 sw
tri 2817 2444 2819 2446 ne
rect 2819 2444 2883 2446
tri 2883 2444 2885 2446 sw
tri 2928 2444 2930 2446 ne
rect 2930 2444 3518 2446
tri 3518 2444 3520 2446 sw
rect 2342 2442 2414 2444
tri 2414 2442 2416 2444 sw
tri 2496 2442 2498 2444 ne
rect 2498 2442 2562 2444
tri 2562 2442 2564 2444 sw
tri 2622 2442 2624 2444 ne
rect 2624 2442 2688 2444
tri 2688 2442 2690 2444 sw
tri 2819 2442 2821 2444 ne
rect 2821 2442 2885 2444
rect 2215 2441 2266 2442
tri 2266 2441 2267 2442 sw
tri 2342 2441 2343 2442 ne
rect 2343 2441 2416 2442
tri 2416 2441 2417 2442 sw
tri 2498 2441 2499 2442 ne
rect 2499 2441 2564 2442
tri 2564 2441 2565 2442 sw
tri 2624 2441 2625 2442 ne
rect 2625 2441 2690 2442
tri 2690 2441 2691 2442 sw
tri 2821 2441 2822 2442 ne
rect 2822 2441 2885 2442
tri 2885 2441 2888 2444 sw
tri 2930 2441 2933 2444 ne
rect 2933 2441 3520 2444
tri 3520 2441 3523 2444 sw
rect 2215 2435 2267 2441
rect 2093 2409 2267 2435
rect 2093 2375 2099 2409
rect 2133 2407 2267 2409
tri 2267 2407 2301 2441 sw
tri 2343 2407 2377 2441 ne
rect 2377 2422 2417 2441
tri 2417 2422 2436 2441 sw
tri 2499 2422 2518 2441 ne
rect 2518 2422 2565 2441
tri 2565 2422 2584 2441 sw
tri 2625 2432 2634 2441 ne
rect 2634 2432 2691 2441
tri 2691 2432 2700 2441 sw
tri 2822 2432 2831 2441 ne
rect 2831 2432 2888 2441
tri 2634 2422 2644 2432 ne
rect 2644 2422 2700 2432
tri 2700 2422 2710 2432 sw
tri 2831 2422 2841 2432 ne
rect 2841 2422 2888 2432
tri 2888 2422 2907 2441 sw
tri 2933 2422 2952 2441 ne
rect 2952 2434 3523 2441
tri 3523 2434 3530 2441 sw
rect 3932 2434 3978 2446
rect 4119 3049 4284 3083
rect 4119 3015 4125 3049
rect 4159 3045 4284 3049
rect 4159 3015 4244 3045
rect 4119 3011 4244 3015
rect 4278 3011 4284 3045
rect 4119 2973 4284 3011
rect 4119 2939 4125 2973
rect 4159 2939 4244 2973
rect 4278 2939 4284 2973
rect 4119 2901 4284 2939
rect 4119 2897 4244 2901
rect 4119 2863 4125 2897
rect 4159 2867 4244 2897
rect 4278 2867 4284 2901
rect 4159 2863 4284 2867
rect 4119 2829 4284 2863
rect 4119 2821 4244 2829
rect 4119 2787 4125 2821
rect 4159 2795 4244 2821
rect 4278 2795 4284 2829
rect 4159 2787 4284 2795
rect 4119 2757 4284 2787
rect 4119 2745 4244 2757
rect 4119 2711 4125 2745
rect 4159 2723 4244 2745
rect 4278 2723 4284 2757
rect 4159 2711 4284 2723
rect 4119 2685 4284 2711
rect 4119 2669 4244 2685
rect 4119 2635 4125 2669
rect 4159 2651 4244 2669
rect 4278 2651 4284 2685
rect 4159 2635 4284 2651
rect 4119 2613 4284 2635
rect 4119 2593 4244 2613
rect 4119 2559 4125 2593
rect 4159 2579 4244 2593
rect 4278 2579 4284 2613
rect 4159 2567 4284 2579
rect 4394 3549 4440 3561
rect 4394 3515 4400 3549
rect 4434 3515 4440 3549
rect 4394 3477 4440 3515
rect 4394 3443 4400 3477
rect 4434 3443 4440 3477
rect 4394 3405 4440 3443
rect 4394 3371 4400 3405
rect 4434 3371 4440 3405
rect 4394 3333 4440 3371
rect 4394 3299 4400 3333
rect 4434 3299 4440 3333
rect 4394 3261 4440 3299
rect 4394 3227 4400 3261
rect 4434 3227 4440 3261
rect 4394 3189 4440 3227
rect 4394 3155 4400 3189
rect 4434 3155 4440 3189
rect 4394 3117 4440 3155
rect 4394 3083 4400 3117
rect 4434 3083 4440 3117
rect 4394 3045 4440 3083
rect 4394 3011 4400 3045
rect 4434 3011 4440 3045
rect 4394 2973 4440 3011
rect 4394 2939 4400 2973
rect 4434 2939 4440 2973
rect 4394 2901 4440 2939
rect 4394 2867 4400 2901
rect 4434 2867 4440 2901
rect 4394 2829 4440 2867
rect 4394 2795 4400 2829
rect 4434 2795 4440 2829
rect 4394 2757 4440 2795
rect 4394 2723 4400 2757
rect 4434 2723 4440 2757
rect 4394 2685 4440 2723
rect 4394 2651 4400 2685
rect 4434 2651 4440 2685
rect 4394 2613 4440 2651
rect 4394 2579 4400 2613
rect 4434 2579 4440 2613
rect 4159 2559 4258 2567
tri 4258 2559 4266 2567 nw
rect 4119 2553 4252 2559
tri 4252 2553 4258 2559 nw
rect 4119 2537 4236 2553
tri 4236 2537 4252 2553 nw
rect 4119 2517 4202 2537
rect 4119 2483 4125 2517
rect 4159 2503 4202 2517
tri 4202 2503 4236 2537 nw
rect 4159 2493 4192 2503
tri 4192 2493 4202 2503 nw
rect 4159 2483 4187 2493
tri 4187 2488 4192 2493 nw
tri 4312 2488 4317 2493 se
rect 4317 2488 4363 2493
tri 4311 2487 4312 2488 se
rect 4312 2487 4363 2488
rect 4119 2441 4187 2483
rect 2952 2422 3530 2434
rect 2377 2407 2436 2422
tri 2436 2407 2451 2422 sw
tri 2518 2407 2533 2422 ne
rect 2533 2407 2584 2422
tri 2584 2407 2599 2422 sw
tri 2644 2407 2659 2422 ne
rect 2659 2407 2710 2422
tri 2710 2407 2725 2422 sw
tri 2841 2407 2856 2422 ne
rect 2856 2421 2907 2422
tri 2907 2421 2908 2422 sw
tri 2952 2421 2953 2422 ne
rect 2953 2421 3530 2422
rect 2856 2407 2908 2421
tri 2908 2407 2922 2421 sw
tri 2953 2412 2962 2421 ne
rect 2962 2412 3530 2421
tri 3486 2407 3491 2412 ne
rect 3491 2407 3530 2412
tri 3530 2407 3557 2434 sw
rect 4119 2407 4125 2441
rect 4159 2407 4187 2441
rect 4235 2435 4241 2487
rect 4293 2435 4305 2487
rect 4357 2435 4363 2487
tri 4257 2428 4264 2435 ne
rect 4264 2428 4363 2435
tri 4264 2409 4283 2428 ne
rect 4283 2409 4363 2428
rect 2133 2402 2301 2407
tri 2301 2402 2306 2407 sw
tri 2377 2402 2382 2407 ne
rect 2382 2402 2451 2407
tri 2451 2402 2456 2407 sw
tri 2533 2402 2538 2407 ne
rect 2538 2402 2599 2407
tri 2599 2402 2604 2407 sw
tri 2659 2403 2663 2407 ne
rect 2663 2403 2725 2407
tri 2663 2402 2664 2403 ne
rect 2664 2402 2725 2403
tri 2725 2402 2730 2407 sw
tri 2856 2402 2861 2407 ne
rect 2861 2402 2922 2407
tri 2922 2402 2927 2407 sw
tri 3491 2402 3496 2407 ne
rect 3496 2402 3557 2407
tri 3557 2402 3562 2407 sw
rect 2133 2375 2306 2402
tri 2306 2375 2333 2402 sw
tri 2382 2375 2409 2402 ne
rect 2409 2401 2456 2402
tri 2456 2401 2457 2402 sw
tri 2538 2401 2539 2402 ne
rect 2539 2401 2604 2402
tri 2604 2401 2605 2402 sw
tri 2664 2401 2665 2402 ne
rect 2665 2401 2730 2402
tri 2730 2401 2731 2402 sw
tri 2861 2401 2862 2402 ne
rect 2862 2401 2927 2402
rect 2409 2378 2457 2401
tri 2457 2378 2480 2401 sw
tri 2539 2378 2562 2401 ne
rect 2562 2378 2605 2401
tri 2605 2378 2628 2401 sw
tri 2665 2378 2688 2401 ne
rect 2688 2378 2731 2401
tri 2731 2378 2754 2401 sw
tri 2862 2378 2885 2401 ne
rect 2885 2387 2927 2401
tri 2927 2387 2942 2402 sw
tri 3496 2388 3510 2402 ne
rect 3510 2388 3562 2402
tri 3562 2388 3576 2402 sw
tri 3510 2387 3511 2388 ne
rect 3511 2387 3576 2388
tri 3576 2387 3577 2388 sw
rect 2885 2378 2942 2387
tri 2942 2378 2951 2387 sw
tri 3511 2378 3520 2387 ne
rect 3520 2378 3577 2387
tri 3577 2378 3586 2387 sw
rect 2409 2375 2480 2378
tri 2480 2375 2483 2378 sw
tri 2562 2375 2565 2378 ne
rect 2565 2375 2628 2378
tri 2628 2375 2631 2378 sw
tri 2688 2375 2691 2378 ne
rect 2691 2375 2754 2378
tri 2754 2375 2757 2378 sw
tri 2885 2375 2888 2378 ne
rect 2888 2375 3470 2378
tri 3470 2375 3473 2378 sw
tri 3520 2375 3523 2378 ne
rect 3523 2375 3586 2378
tri 3586 2375 3589 2378 sw
rect 2093 2368 2333 2375
tri 2333 2368 2340 2375 sw
tri 2409 2368 2416 2375 ne
rect 2416 2368 2483 2375
tri 2483 2368 2490 2375 sw
tri 2565 2368 2572 2375 ne
rect 2572 2368 2631 2375
tri 2631 2368 2638 2375 sw
tri 2691 2368 2698 2375 ne
rect 2698 2368 2757 2375
tri 2757 2368 2764 2375 sw
tri 2888 2368 2895 2375 ne
rect 2895 2368 3473 2375
rect 2093 2365 2340 2368
tri 2340 2365 2343 2368 sw
tri 2416 2365 2419 2368 ne
rect 2419 2365 2490 2368
tri 2490 2365 2493 2368 sw
tri 2572 2365 2575 2368 ne
rect 2575 2365 2638 2368
tri 2638 2365 2641 2368 sw
tri 2698 2366 2700 2368 ne
rect 2700 2366 2764 2368
tri 2764 2366 2766 2368 sw
tri 2895 2366 2897 2368 ne
rect 2897 2366 3473 2368
tri 2700 2365 2701 2366 ne
rect 2701 2365 2766 2366
tri 2766 2365 2767 2366 sw
tri 2897 2365 2898 2366 ne
rect 2898 2365 3473 2366
tri 3473 2365 3483 2375 sw
tri 3523 2365 3533 2375 ne
rect 3533 2365 3589 2375
tri 3589 2365 3599 2375 sw
rect 2093 2363 2343 2365
tri 2343 2363 2345 2365 sw
tri 2419 2363 2421 2365 ne
rect 2421 2363 2493 2365
tri 2493 2363 2495 2365 sw
tri 2575 2363 2577 2365 ne
rect 2577 2363 2641 2365
tri 2641 2363 2643 2365 sw
tri 2701 2363 2703 2365 ne
rect 2703 2363 2767 2365
tri 2767 2363 2769 2365 sw
tri 2898 2363 2900 2365 ne
rect 2900 2363 3483 2365
tri 3483 2363 3485 2365 sw
tri 3533 2363 3535 2365 ne
rect 3535 2363 3599 2365
tri 3599 2363 3601 2365 sw
tri 2271 2331 2303 2363 ne
rect 2303 2331 2345 2363
tri 2345 2331 2377 2363 sw
tri 2421 2331 2453 2363 ne
rect 2453 2354 2495 2363
tri 2495 2354 2504 2363 sw
tri 2577 2356 2584 2363 ne
rect 2584 2356 2643 2363
tri 2643 2356 2650 2363 sw
tri 2703 2356 2710 2363 ne
rect 2710 2356 2769 2363
tri 2769 2356 2776 2363 sw
tri 2900 2356 2907 2363 ne
rect 2907 2356 3485 2363
tri 2584 2354 2586 2356 ne
rect 2586 2354 2650 2356
tri 2650 2354 2652 2356 sw
tri 2710 2354 2712 2356 ne
rect 2712 2354 2776 2356
tri 2776 2354 2778 2356 sw
tri 2907 2354 2909 2356 ne
rect 2909 2354 3485 2356
tri 3485 2354 3494 2363 sw
tri 3535 2354 3544 2363 ne
rect 3544 2354 3601 2363
tri 3601 2354 3610 2363 sw
rect 2453 2332 2504 2354
tri 2504 2332 2526 2354 sw
tri 2586 2332 2608 2354 ne
rect 2608 2332 2652 2354
tri 2652 2332 2674 2354 sw
tri 2712 2332 2734 2354 ne
rect 2734 2332 2778 2354
tri 2778 2332 2800 2354 sw
tri 2909 2332 2931 2354 ne
rect 2931 2338 3494 2354
tri 3494 2338 3510 2354 sw
tri 3544 2338 3560 2354 ne
rect 3560 2338 3610 2354
rect 2931 2332 3510 2338
rect 2453 2331 2526 2332
tri 2526 2331 2527 2332 sw
tri 2608 2331 2609 2332 ne
rect 2609 2331 2674 2332
tri 2674 2331 2675 2332 sw
tri 2734 2331 2735 2332 ne
rect 2735 2331 2800 2332
tri 2800 2331 2801 2332 sw
tri 3450 2331 3451 2332 ne
rect 3451 2331 3510 2332
tri 3510 2331 3517 2338 sw
tri 3560 2331 3567 2338 ne
rect 3567 2331 3610 2338
tri 3610 2331 3633 2354 sw
rect 3945 2335 3953 2387
rect 4005 2335 4017 2387
rect 4069 2335 4075 2387
tri 2303 2328 2306 2331 ne
rect 2306 2328 2377 2331
tri 2377 2328 2380 2331 sw
tri 2453 2328 2456 2331 ne
rect 2456 2328 2527 2331
tri 2527 2328 2530 2331 sw
tri 2609 2328 2612 2331 ne
rect 2612 2328 2675 2331
tri 2675 2328 2678 2331 sw
tri 2735 2328 2738 2331 ne
rect 2738 2328 2801 2331
tri 2801 2328 2804 2331 sw
tri 3451 2328 3454 2331 ne
rect 3454 2328 3517 2331
tri 3517 2328 3520 2331 sw
tri 3567 2328 3570 2331 ne
rect 3570 2328 3633 2331
tri 3633 2328 3636 2331 sw
tri 2306 2294 2340 2328 ne
rect 2340 2294 2380 2328
tri 2380 2294 2414 2328 sw
tri 2456 2294 2490 2328 ne
rect 2490 2294 2530 2328
tri 2530 2294 2564 2328 sw
tri 2612 2294 2646 2328 ne
rect 2646 2306 2678 2328
tri 2678 2306 2700 2328 sw
tri 2738 2306 2760 2328 ne
rect 2760 2306 2804 2328
rect 2646 2300 2700 2306
tri 2700 2300 2706 2306 sw
tri 2760 2300 2766 2306 ne
rect 2766 2300 2804 2306
tri 2804 2300 2832 2328 sw
tri 3454 2300 3482 2328 ne
rect 3482 2322 3520 2328
tri 3520 2322 3526 2328 sw
tri 3570 2322 3576 2328 ne
rect 3576 2322 3636 2328
tri 3636 2322 3642 2328 sw
rect 3482 2300 3526 2322
rect 2646 2294 2706 2300
tri 2706 2294 2712 2300 sw
tri 2766 2294 2772 2300 ne
rect 2772 2294 3137 2300
tri 3137 2294 3143 2300 sw
tri 3482 2294 3488 2300 ne
rect 3488 2294 3526 2300
tri 3526 2294 3554 2322 sw
tri 3576 2302 3596 2322 ne
tri 2340 2289 2345 2294 ne
rect 2345 2289 2414 2294
tri 2414 2289 2419 2294 sw
tri 2490 2289 2495 2294 ne
rect 2495 2289 2564 2294
tri 2564 2289 2569 2294 sw
tri 2646 2290 2650 2294 ne
rect 2650 2290 2712 2294
tri 2712 2290 2716 2294 sw
tri 2772 2290 2776 2294 ne
rect 2776 2290 3143 2294
tri 3143 2290 3147 2294 sw
tri 3488 2290 3492 2294 ne
rect 3492 2290 3554 2294
tri 2650 2289 2651 2290 ne
rect 2651 2289 2716 2290
tri 2716 2289 2717 2290 sw
tri 2776 2289 2777 2290 ne
rect 2777 2289 3147 2290
tri 3147 2289 3148 2290 sw
tri 3492 2289 3493 2290 ne
rect 3493 2289 3554 2290
tri 3554 2289 3559 2294 sw
tri 2345 2255 2379 2289 ne
rect 2379 2255 2419 2289
tri 2419 2255 2453 2289 sw
tri 2495 2255 2529 2289 ne
rect 2529 2288 2569 2289
tri 2569 2288 2570 2289 sw
tri 2651 2288 2652 2289 ne
rect 2652 2288 2717 2289
tri 2717 2288 2718 2289 sw
tri 2777 2288 2778 2289 ne
rect 2778 2288 3148 2289
tri 3148 2288 3149 2289 sw
tri 3493 2288 3494 2289 ne
rect 3494 2288 3559 2289
tri 3559 2288 3560 2289 sw
rect 2529 2268 2570 2288
tri 2570 2268 2590 2288 sw
tri 2652 2268 2672 2288 ne
rect 2672 2268 2718 2288
tri 2718 2268 2738 2288 sw
tri 2778 2268 2798 2288 ne
rect 2798 2268 3149 2288
tri 3149 2268 3169 2288 sw
tri 3494 2268 3514 2288 ne
rect 2529 2255 2590 2268
tri 2590 2255 2603 2268 sw
tri 2672 2255 2685 2268 ne
rect 2685 2255 2738 2268
tri 2738 2255 2751 2268 sw
tri 2798 2255 2811 2268 ne
rect 2811 2255 3169 2268
tri 3169 2255 3182 2268 sw
tri 2002 2254 2003 2255 se
rect 2003 2254 2060 2255
tri 2379 2254 2380 2255 ne
rect 2380 2254 2453 2255
tri 2453 2254 2454 2255 sw
tri 2529 2254 2530 2255 ne
rect 2530 2254 2603 2255
tri 2603 2254 2604 2255 sw
tri 2685 2254 2686 2255 ne
rect 2686 2254 2751 2255
tri 2751 2254 2752 2255 sw
tri 2811 2254 2812 2255 ne
rect 2812 2254 3182 2255
tri 3182 2254 3183 2255 sw
tri 1996 2248 2002 2254 se
rect 2002 2248 2060 2254
tri 2380 2248 2386 2254 ne
rect 2386 2249 2454 2254
tri 2454 2249 2459 2254 sw
tri 2530 2249 2535 2254 ne
rect 2535 2249 2604 2254
tri 2604 2249 2609 2254 sw
tri 2686 2249 2691 2254 ne
rect 2691 2249 2752 2254
tri 2752 2249 2757 2254 sw
tri 3071 2249 3076 2254 ne
rect 3076 2249 3183 2254
tri 3183 2249 3188 2254 sw
rect 2386 2248 2459 2249
tri 2459 2248 2460 2249 sw
tri 2535 2248 2536 2249 ne
rect 2536 2248 2609 2249
tri 2609 2248 2610 2249 sw
tri 2691 2248 2692 2249 ne
rect 2692 2248 2757 2249
tri 2757 2248 2758 2249 sw
tri 3076 2248 3077 2249 ne
rect 3077 2248 3188 2249
tri 3188 2248 3189 2249 sw
tri 1987 2239 1996 2248 se
rect 1996 2239 2060 2248
tri 1975 2227 1987 2239 se
rect 1987 2227 2060 2239
tri 1611 2205 1631 2225 sw
rect 1565 2196 1631 2205
tri 1631 2196 1640 2205 sw
rect 1565 2159 1640 2196
tri 1565 2147 1577 2159 ne
rect 1577 2147 1640 2159
tri 1640 2147 1689 2196 sw
rect 1932 2175 1938 2227
rect 1990 2175 2002 2227
rect 2054 2175 2060 2227
rect 2140 2196 2146 2248
rect 2198 2196 2212 2248
rect 2264 2220 2324 2248
tri 2324 2220 2352 2248 sw
tri 2386 2220 2414 2248 ne
rect 2414 2220 2460 2248
tri 2460 2220 2488 2248 sw
tri 2536 2220 2564 2248 ne
rect 2564 2224 2610 2248
tri 2610 2224 2634 2248 sw
tri 2692 2224 2716 2248 ne
rect 2716 2224 2758 2248
tri 2758 2224 2782 2248 sw
tri 3077 2224 3101 2248 ne
rect 3101 2224 3189 2248
tri 3189 2224 3213 2248 sw
rect 2564 2220 2634 2224
tri 2634 2220 2638 2224 sw
tri 2716 2220 2720 2224 ne
rect 2720 2220 2803 2224
rect 2264 2201 2352 2220
tri 2352 2201 2371 2220 sw
tri 2414 2201 2433 2220 ne
rect 2433 2201 2488 2220
tri 2488 2201 2507 2220 sw
rect 2564 2201 2638 2220
tri 2638 2201 2657 2220 sw
tri 2720 2201 2739 2220 ne
rect 2739 2201 2803 2220
rect 2264 2196 2371 2201
tri 2371 2196 2376 2201 sw
tri 2433 2196 2438 2201 ne
rect 2438 2196 2507 2201
tri 2507 2196 2512 2201 sw
rect 2564 2196 2657 2201
tri 2657 2196 2662 2201 sw
tri 2739 2196 2744 2201 ne
rect 2744 2196 2803 2201
tri 2302 2175 2323 2196 ne
rect 2323 2192 2376 2196
tri 2376 2192 2380 2196 sw
tri 2438 2192 2442 2196 ne
rect 2442 2192 2512 2196
rect 2323 2180 2380 2192
tri 2380 2180 2392 2192 sw
tri 2442 2180 2454 2192 ne
rect 2454 2180 2512 2192
tri 2512 2180 2528 2196 sw
rect 2323 2175 2392 2180
tri 2323 2147 2351 2175 ne
rect 2351 2149 2392 2175
tri 2392 2149 2423 2180 sw
tri 2454 2158 2476 2180 ne
rect 2351 2147 2423 2149
tri 1577 2122 1602 2147 ne
rect 1602 2127 2236 2147
tri 2236 2127 2256 2147 sw
tri 2351 2127 2371 2147 ne
rect 1602 2122 2256 2127
tri 2256 2122 2261 2127 sw
tri 1602 2117 1607 2122 ne
rect 1607 2117 2261 2122
tri 1534 2113 1538 2117 sw
tri 1607 2113 1611 2117 ne
rect 1611 2113 2261 2117
rect 1488 2101 1538 2113
tri 1538 2101 1550 2113 sw
tri 1611 2101 1623 2113 ne
rect 1623 2101 2261 2113
rect 1488 2071 1550 2101
tri 1550 2071 1580 2101 sw
tri 2216 2071 2246 2101 ne
rect 2246 2071 2261 2101
tri 2261 2071 2312 2122 sw
rect 1488 2065 1580 2071
tri 1580 2065 1586 2071 sw
tri 2246 2065 2252 2071 ne
rect 2252 2065 2312 2071
tri 2312 2065 2318 2071 sw
rect 1488 2053 2167 2065
tri 2252 2056 2261 2065 ne
rect 2261 2056 2318 2065
tri 2318 2056 2327 2065 sw
rect 1488 2052 2127 2053
tri 1488 2048 1492 2052 ne
rect 1492 2048 2127 2052
tri 669 2026 673 2030 sw
tri 1198 2026 1202 2030 se
rect 1202 2026 1251 2030
tri 612 2021 617 2026 se
rect 617 2021 673 2026
tri 673 2021 678 2026 sw
tri 1193 2021 1198 2026 se
rect 1198 2021 1251 2026
tri 1492 2021 1519 2048 ne
rect 1519 2021 2127 2048
tri 610 2019 612 2021 se
rect 612 2019 678 2021
tri 678 2019 680 2021 sw
tri 1191 2019 1193 2021 se
rect 1193 2019 1251 2021
tri 1251 2019 1253 2021 sw
tri 1519 2019 1521 2021 ne
rect 1521 2019 2127 2021
rect 2161 2019 2167 2053
tri 2261 2041 2276 2056 ne
rect 2276 2041 2327 2056
tri 2276 2036 2281 2041 ne
tri 598 2007 610 2019 se
rect 610 2007 680 2019
tri 680 2007 692 2019 sw
tri 1179 2007 1191 2019 se
rect 1191 2007 1253 2019
tri 1253 2007 1265 2019 sw
tri 2037 2007 2049 2019 ne
rect 2049 2007 2167 2019
tri 590 1999 598 2007 se
rect 598 1999 692 2007
tri 692 1999 700 2007 sw
tri 1171 1999 1179 2007 se
rect 1179 1999 1265 2007
tri 1265 1999 1273 2007 sw
tri 2049 1999 2057 2007 ne
rect 2057 1999 2167 2007
tri 583 1992 590 1999 se
rect 590 1992 700 1999
tri 700 1992 707 1999 sw
tri 1164 1992 1171 1999 se
rect 1171 1992 1273 1999
tri 1273 1992 1280 1999 sw
tri 2057 1992 2064 1999 ne
rect 2064 1992 2167 1999
rect 172 1986 919 1992
tri 1161 1989 1164 1992 se
rect 1164 1989 1280 1992
tri 1280 1989 1283 1992 sw
tri 2064 1989 2067 1992 ne
rect 2067 1989 2167 1992
rect 172 1952 184 1986
rect 218 1952 261 1986
rect 295 1952 338 1986
rect 372 1952 415 1986
rect 449 1952 492 1986
rect 526 1952 569 1986
rect 603 1952 645 1986
rect 679 1952 721 1986
rect 755 1952 797 1986
rect 831 1952 873 1986
rect 907 1952 919 1986
rect 172 1946 919 1952
rect 1058 1983 1754 1989
rect 1058 1949 1070 1983
rect 1104 1949 1145 1983
rect 1179 1949 1220 1983
rect 1254 1949 1294 1983
rect 1328 1949 1368 1983
rect 1402 1949 1442 1983
rect 1476 1949 1516 1983
rect 1550 1949 1590 1983
rect 1624 1949 1664 1983
rect 1698 1949 1738 1983
rect 1058 1943 1754 1949
tri 1742 1937 1748 1943 ne
rect 1748 1937 1754 1943
rect 1806 1937 1821 1989
rect 1873 1937 1888 1989
rect 1940 1937 1955 1989
rect 2007 1937 2013 1989
tri 2067 1983 2073 1989 ne
rect 2073 1983 2167 1989
tri 2073 1981 2075 1983 ne
rect 2075 1981 2167 1983
tri 2075 1947 2109 1981 ne
rect 2109 1947 2127 1981
rect 2161 1947 2167 1981
tri 1926 1935 1928 1937 ne
rect 1928 1935 2013 1937
tri 2109 1935 2121 1947 ne
rect 2121 1935 2167 1947
tri 1928 1933 1930 1935 ne
rect 1930 1933 2013 1935
tri 1930 1896 1967 1933 ne
rect -11 1833 -5 1867
rect 29 1833 41 1867
rect -11 1795 41 1833
rect -11 1761 -5 1795
rect 29 1761 41 1795
rect -11 1723 41 1761
rect -11 1689 -5 1723
rect 29 1689 41 1723
rect -11 1651 41 1689
rect -11 1617 -5 1651
rect 29 1617 41 1651
rect -11 1579 41 1617
rect -11 1545 -5 1579
rect 29 1545 41 1579
tri -181 1524 -178 1527 sw
rect -230 1518 -178 1524
rect -230 1454 -178 1466
rect -230 1401 -221 1402
rect -187 1401 -178 1402
rect -230 1396 -178 1401
tri -230 1393 -227 1396 ne
rect -310 1235 -258 1247
rect -310 1177 -258 1183
rect -227 1363 -181 1396
tri -181 1393 -178 1396 nw
rect -11 1507 41 1545
rect 120 1867 166 1879
rect 120 1833 126 1867
rect 160 1833 166 1867
rect 120 1795 166 1833
rect 120 1761 126 1795
rect 160 1761 166 1795
rect 120 1723 166 1761
rect 120 1689 126 1723
rect 160 1689 166 1723
rect 336 1867 382 1879
rect 336 1833 342 1867
rect 376 1833 382 1867
rect 336 1795 382 1833
rect 336 1761 342 1795
rect 376 1761 382 1795
rect 336 1723 382 1761
rect 120 1651 166 1689
rect 120 1617 126 1651
rect 160 1617 166 1651
rect 120 1579 166 1617
rect 120 1545 126 1579
rect 160 1545 166 1579
tri 333 1699 336 1702 se
rect 336 1699 342 1723
rect 333 1693 342 1699
rect 376 1699 382 1723
rect 552 1867 598 1879
rect 552 1833 558 1867
rect 592 1833 598 1867
rect 552 1795 598 1833
rect 552 1761 558 1795
rect 592 1761 598 1795
rect 552 1723 598 1761
tri 382 1699 385 1702 sw
rect 376 1693 385 1699
rect 333 1629 342 1641
rect 376 1629 385 1641
rect 333 1571 342 1577
tri 333 1568 336 1571 ne
rect -11 1473 -5 1507
rect 29 1473 41 1507
rect -11 1435 41 1473
rect -11 1401 -5 1435
rect 29 1401 41 1435
rect -227 1329 -221 1363
rect -187 1329 -181 1363
rect -227 1291 -181 1329
rect -227 1257 -221 1291
rect -187 1257 -181 1291
rect -227 1219 -181 1257
rect -227 1185 -221 1219
rect -187 1185 -181 1219
rect -227 1147 -181 1185
rect -227 1113 -221 1147
rect -187 1113 -181 1147
rect -227 1075 -181 1113
rect -227 1041 -221 1075
rect -187 1041 -181 1075
rect -227 1003 -181 1041
rect -227 969 -221 1003
rect -187 969 -181 1003
rect -227 931 -181 969
rect -227 897 -221 931
rect -187 897 -181 931
rect -227 885 -181 897
rect -11 1363 41 1401
tri 117 1524 120 1527 se
rect 120 1524 166 1545
rect 336 1545 342 1571
rect 376 1571 385 1577
rect 376 1545 382 1571
tri 382 1568 385 1571 nw
rect 552 1689 558 1723
rect 592 1689 598 1723
rect 552 1651 598 1689
rect 552 1617 558 1651
rect 592 1617 598 1651
rect 552 1579 598 1617
tri 166 1524 169 1527 sw
rect 117 1518 169 1524
rect 117 1454 169 1466
rect 117 1401 126 1402
rect 160 1401 169 1402
rect 117 1396 169 1401
tri 117 1393 120 1396 ne
rect -11 1329 -5 1363
rect 29 1329 41 1363
rect -11 1291 41 1329
rect -11 1257 -5 1291
rect 29 1257 41 1291
rect -11 1219 41 1257
rect -11 1185 -5 1219
rect 29 1185 41 1219
rect -11 1147 41 1185
rect -11 1113 -5 1147
rect 29 1113 41 1147
rect -11 1075 41 1113
rect -11 1041 -5 1075
rect 29 1041 41 1075
rect -11 1003 41 1041
rect -11 969 -5 1003
rect 29 969 41 1003
rect -11 931 41 969
rect -11 897 -5 931
rect 29 897 41 931
rect -11 885 41 897
rect 120 1363 166 1396
tri 166 1393 169 1396 nw
rect 336 1507 382 1545
rect 552 1545 558 1579
rect 592 1545 598 1579
rect 336 1473 342 1507
rect 376 1473 382 1507
rect 336 1435 382 1473
rect 336 1401 342 1435
rect 376 1401 382 1435
rect 120 1329 126 1363
rect 160 1329 166 1363
rect 120 1291 166 1329
rect 120 1257 126 1291
rect 160 1257 166 1291
rect 120 1219 166 1257
rect 120 1185 126 1219
rect 160 1185 166 1219
rect 120 1147 166 1185
rect 120 1113 126 1147
rect 160 1113 166 1147
rect 120 1075 166 1113
rect 120 1041 126 1075
rect 160 1041 166 1075
rect 120 1003 166 1041
rect 120 969 126 1003
rect 160 969 166 1003
rect 120 931 166 969
rect 120 897 126 931
rect 160 897 166 931
rect 120 885 166 897
rect 336 1363 382 1401
tri 549 1524 552 1527 se
rect 552 1524 598 1545
rect 768 1867 814 1879
rect 768 1833 774 1867
rect 808 1833 814 1867
rect 768 1795 814 1833
rect 768 1761 774 1795
rect 808 1761 814 1795
rect 768 1723 814 1761
rect 768 1689 774 1723
rect 808 1689 814 1723
rect 768 1651 814 1689
rect 768 1617 774 1651
rect 808 1617 814 1651
rect 768 1579 814 1617
rect 768 1545 774 1579
rect 808 1545 814 1579
tri 598 1524 601 1527 sw
rect 549 1518 601 1524
rect 549 1454 601 1466
rect 549 1401 558 1402
rect 592 1401 601 1402
rect 549 1396 601 1401
tri 549 1393 552 1396 ne
rect 336 1329 342 1363
rect 376 1329 382 1363
rect 336 1291 382 1329
rect 336 1257 342 1291
rect 376 1257 382 1291
rect 336 1219 382 1257
rect 336 1185 342 1219
rect 376 1185 382 1219
rect 336 1147 382 1185
rect 336 1113 342 1147
rect 376 1113 382 1147
rect 336 1075 382 1113
rect 336 1041 342 1075
rect 376 1041 382 1075
rect 336 1003 382 1041
rect 336 969 342 1003
rect 376 969 382 1003
rect 336 931 382 969
rect 336 897 342 931
rect 376 897 382 931
rect 336 885 382 897
rect 552 1363 598 1396
tri 598 1393 601 1396 nw
rect 768 1507 814 1545
rect 984 1867 1030 1879
rect 984 1833 990 1867
rect 1024 1833 1030 1867
rect 984 1795 1030 1833
rect 984 1761 990 1795
rect 1024 1761 1030 1795
rect 984 1723 1030 1761
tri 1197 1869 1200 1872 se
rect 1200 1869 1246 1879
tri 1246 1869 1249 1872 sw
rect 1197 1867 1249 1869
rect 1197 1863 1206 1867
rect 1240 1863 1249 1867
rect 1197 1799 1249 1811
rect 1197 1741 1249 1747
tri 1197 1738 1200 1741 ne
rect 984 1689 990 1723
rect 1024 1689 1030 1723
rect 984 1651 1030 1689
rect 984 1617 990 1651
rect 1024 1617 1030 1651
rect 984 1579 1030 1617
rect 984 1545 990 1579
rect 1024 1545 1030 1579
rect 768 1473 774 1507
rect 808 1473 814 1507
rect 768 1435 814 1473
rect 768 1401 774 1435
rect 808 1401 814 1435
rect 552 1329 558 1363
rect 592 1329 598 1363
rect 552 1291 598 1329
rect 552 1257 558 1291
rect 592 1257 598 1291
rect 552 1219 598 1257
rect 552 1185 558 1219
rect 592 1185 598 1219
rect 552 1147 598 1185
rect 552 1113 558 1147
rect 592 1113 598 1147
rect 552 1075 598 1113
rect 768 1363 814 1401
tri 981 1524 984 1527 se
rect 984 1524 1030 1545
rect 1200 1723 1246 1741
tri 1246 1738 1249 1741 nw
rect 1416 1867 1462 1879
rect 1416 1833 1422 1867
rect 1456 1833 1462 1867
rect 1416 1795 1462 1833
rect 1416 1761 1422 1795
rect 1456 1761 1462 1795
rect 1200 1689 1206 1723
rect 1240 1689 1246 1723
rect 1200 1651 1246 1689
rect 1200 1617 1206 1651
rect 1240 1617 1246 1651
rect 1200 1579 1246 1617
rect 1200 1545 1206 1579
rect 1240 1545 1246 1579
tri 1030 1524 1033 1527 sw
rect 981 1518 1033 1524
rect 981 1454 1033 1466
rect 981 1401 990 1402
rect 1024 1401 1033 1402
rect 981 1396 1033 1401
tri 981 1393 984 1396 ne
rect 768 1329 774 1363
rect 808 1329 814 1363
rect 768 1291 814 1329
rect 768 1257 774 1291
rect 808 1257 814 1291
rect 768 1219 814 1257
rect 768 1185 774 1219
rect 808 1185 814 1219
rect 768 1147 814 1185
rect 768 1113 774 1147
rect 808 1113 814 1147
rect 552 1041 558 1075
rect 592 1041 598 1075
rect 552 1003 598 1041
rect 552 969 558 1003
rect 592 969 598 1003
rect 552 931 598 969
rect 552 897 558 931
rect 592 897 598 931
rect 552 885 598 897
tri 765 1083 768 1086 se
rect 768 1083 814 1113
rect 984 1363 1030 1396
tri 1030 1393 1033 1396 nw
rect 1200 1507 1246 1545
rect 1416 1723 1462 1761
tri 1629 1869 1632 1872 se
rect 1632 1869 1678 1879
tri 1678 1869 1681 1872 sw
rect 1629 1867 1681 1869
rect 1629 1863 1638 1867
rect 1672 1863 1681 1867
rect 1629 1799 1681 1811
rect 1629 1741 1681 1747
tri 1629 1738 1632 1741 ne
rect 1416 1689 1422 1723
rect 1456 1689 1462 1723
rect 1416 1651 1462 1689
rect 1416 1617 1422 1651
rect 1456 1617 1462 1651
rect 1416 1579 1462 1617
rect 1416 1545 1422 1579
rect 1456 1545 1462 1579
rect 1200 1473 1206 1507
rect 1240 1473 1246 1507
rect 1200 1435 1246 1473
rect 1200 1401 1206 1435
rect 1240 1401 1246 1435
rect 984 1329 990 1363
rect 1024 1329 1030 1363
rect 984 1291 1030 1329
rect 984 1257 990 1291
rect 1024 1257 1030 1291
rect 984 1219 1030 1257
rect 984 1185 990 1219
rect 1024 1185 1030 1219
rect 984 1147 1030 1185
rect 984 1113 990 1147
rect 1024 1113 1030 1147
tri 814 1083 817 1086 sw
rect 765 1077 817 1083
rect 765 1013 817 1025
rect 765 949 817 961
rect 765 885 817 897
rect 984 1075 1030 1113
rect 984 1041 990 1075
rect 1024 1041 1030 1075
rect 984 1003 1030 1041
rect 984 969 990 1003
rect 1024 969 1030 1003
rect 984 931 1030 969
rect 984 897 990 931
rect 1024 897 1030 931
rect 984 885 1030 897
rect 1200 1363 1246 1401
tri 1413 1524 1416 1527 se
rect 1416 1524 1462 1545
rect 1632 1723 1678 1741
tri 1678 1738 1681 1741 nw
rect 1848 1867 1894 1879
rect 1848 1833 1854 1867
rect 1888 1833 1894 1867
rect 1848 1795 1894 1833
rect 1848 1761 1854 1795
rect 1888 1761 1894 1795
rect 1632 1689 1638 1723
rect 1672 1689 1678 1723
rect 1632 1651 1678 1689
rect 1632 1617 1638 1651
rect 1672 1617 1678 1651
rect 1632 1579 1678 1617
rect 1632 1545 1638 1579
rect 1672 1545 1678 1579
tri 1462 1524 1465 1527 sw
rect 1413 1518 1465 1524
rect 1413 1454 1465 1466
rect 1413 1401 1422 1402
rect 1456 1401 1465 1402
rect 1413 1396 1465 1401
tri 1413 1393 1416 1396 ne
rect 1200 1329 1206 1363
rect 1240 1329 1246 1363
rect 1200 1291 1246 1329
rect 1200 1257 1206 1291
rect 1240 1257 1246 1291
rect 1200 1219 1246 1257
rect 1200 1185 1206 1219
rect 1240 1185 1246 1219
rect 1200 1147 1246 1185
rect 1200 1113 1206 1147
rect 1240 1113 1246 1147
rect 1200 1075 1246 1113
rect 1200 1041 1206 1075
rect 1240 1041 1246 1075
rect 1200 1003 1246 1041
rect 1200 969 1206 1003
rect 1240 969 1246 1003
rect 1200 931 1246 969
rect 1200 897 1206 931
rect 1240 897 1246 931
rect 1200 885 1246 897
rect 1416 1363 1462 1396
tri 1462 1393 1465 1396 nw
rect 1632 1507 1678 1545
rect 1848 1723 1894 1761
rect 1848 1689 1854 1723
rect 1888 1689 1894 1723
rect 1848 1651 1894 1689
rect 1848 1617 1854 1651
rect 1888 1617 1894 1651
rect 1848 1579 1894 1617
rect 1848 1545 1854 1579
rect 1888 1545 1894 1579
tri 1964 1699 1967 1702 se
rect 1967 1699 2013 1933
rect 2125 1820 2171 1832
rect 2125 1786 2131 1820
rect 2165 1786 2171 1820
rect 2125 1748 2171 1786
rect 2125 1714 2131 1748
rect 2165 1714 2171 1748
tri 2013 1699 2016 1702 sw
rect 1964 1693 2016 1699
rect 1964 1629 2016 1641
rect 1964 1571 2016 1577
tri 1964 1570 1965 1571 ne
rect 1965 1570 2015 1571
tri 2015 1570 2016 1571 nw
rect 2125 1676 2171 1714
rect 2125 1642 2131 1676
rect 2165 1642 2171 1676
rect 2125 1604 2171 1642
rect 2125 1570 2131 1604
rect 2165 1570 2171 1604
tri 1965 1568 1967 1570 ne
rect 1632 1473 1638 1507
rect 1672 1473 1678 1507
rect 1632 1435 1678 1473
rect 1632 1401 1638 1435
rect 1672 1401 1678 1435
rect 1416 1329 1422 1363
rect 1456 1329 1462 1363
rect 1416 1291 1462 1329
rect 1416 1257 1422 1291
rect 1456 1257 1462 1291
rect 1416 1219 1462 1257
rect 1416 1185 1422 1219
rect 1456 1185 1462 1219
rect 1416 1147 1462 1185
rect 1416 1113 1422 1147
rect 1456 1113 1462 1147
rect 1416 1075 1462 1113
rect 1416 1041 1422 1075
rect 1456 1041 1462 1075
rect 1416 1003 1462 1041
rect 1416 969 1422 1003
rect 1456 969 1462 1003
rect 1416 931 1462 969
rect 1416 897 1422 931
rect 1456 897 1462 931
rect 1416 885 1462 897
rect 1632 1363 1678 1401
tri 1845 1524 1848 1527 se
rect 1848 1524 1894 1545
tri 1894 1524 1897 1527 sw
rect 1845 1518 1897 1524
rect 1845 1454 1897 1466
rect 1845 1401 1854 1402
rect 1888 1401 1897 1402
rect 1845 1396 1897 1401
tri 1845 1393 1848 1396 ne
rect 1632 1329 1638 1363
rect 1672 1329 1678 1363
rect 1632 1291 1678 1329
rect 1632 1257 1638 1291
rect 1672 1257 1678 1291
rect 1632 1219 1678 1257
rect 1632 1185 1638 1219
rect 1672 1185 1678 1219
rect 1632 1147 1678 1185
rect 1632 1113 1638 1147
rect 1672 1113 1678 1147
rect 1632 1075 1678 1113
rect 1632 1041 1638 1075
rect 1672 1041 1678 1075
rect 1632 1003 1678 1041
rect 1632 969 1638 1003
rect 1672 969 1678 1003
rect 1632 931 1678 969
rect 1632 897 1638 931
rect 1672 897 1678 931
rect 1632 885 1678 897
rect 1848 1363 1894 1396
tri 1894 1393 1897 1396 nw
rect 1848 1329 1854 1363
rect 1888 1329 1894 1363
rect 1848 1291 1894 1329
rect 1848 1257 1854 1291
rect 1888 1257 1894 1291
rect 1967 1267 2013 1570
tri 2013 1568 2015 1570 nw
rect 2125 1532 2171 1570
rect 2125 1498 2131 1532
rect 2165 1498 2171 1532
rect 2125 1460 2171 1498
rect 2125 1426 2131 1460
rect 2165 1426 2171 1460
rect 2125 1388 2171 1426
rect 2125 1354 2131 1388
rect 2165 1354 2171 1388
rect 2125 1316 2171 1354
rect 2125 1282 2131 1316
rect 2165 1282 2171 1316
rect 1848 1219 1894 1257
rect 1848 1185 1854 1219
rect 1888 1185 1894 1219
rect 1848 1147 1894 1185
rect 1848 1113 1854 1147
rect 1888 1113 1894 1147
rect 1848 1075 1894 1113
rect 2125 1083 2171 1282
rect 2281 1820 2327 2041
rect 2371 1894 2423 2147
rect 2476 2059 2528 2180
rect 2476 1995 2528 2007
rect 2476 1935 2488 1943
rect 2522 1935 2528 1943
rect 2476 1923 2528 1935
rect 2564 2172 2662 2196
tri 2662 2172 2686 2196 sw
tri 2744 2172 2768 2196 ne
rect 2768 2172 2803 2196
rect 2855 2172 2867 2224
rect 2919 2172 2925 2224
tri 3101 2220 3105 2224 ne
rect 3105 2220 3213 2224
tri 3213 2220 3217 2224 sw
tri 3105 2215 3110 2220 ne
rect 3110 2210 3217 2220
tri 3217 2210 3227 2220 sw
rect 2564 2158 2686 2172
tri 2686 2158 2700 2172 sw
rect 3110 2158 3116 2210
rect 3168 2158 3180 2210
rect 3232 2158 3238 2210
rect 2564 2079 2700 2158
tri 2700 2079 2779 2158 sw
rect 2564 2071 3123 2079
tri 3123 2071 3131 2079 sw
rect 3514 2071 3560 2288
rect 2564 2037 3131 2071
tri 3131 2037 3165 2071 sw
rect 3514 2037 3520 2071
rect 3554 2037 3560 2071
rect 2564 2033 3165 2037
rect 2564 1999 2617 2033
tri 2617 1999 2651 2033 nw
tri 3014 1999 3048 2033 ne
rect 3048 1999 3165 2033
tri 3165 1999 3203 2037 sw
rect 3514 1999 3560 2037
rect 2564 1995 2613 1999
tri 2613 1995 2617 1999 nw
tri 3048 1995 3052 1999 ne
rect 3052 1995 3203 1999
tri 3203 1995 3207 1999 sw
tri 2423 1894 2445 1916 sw
tri 2371 1885 2380 1894 ne
rect 2380 1885 2445 1894
tri 2445 1885 2454 1894 sw
tri 2380 1873 2392 1885 ne
rect 2392 1873 2454 1885
tri 2392 1857 2408 1873 ne
rect 2281 1786 2287 1820
rect 2321 1786 2327 1820
rect 2281 1748 2327 1786
rect 2281 1714 2287 1748
rect 2321 1714 2327 1748
rect 2281 1676 2327 1714
rect 2281 1642 2287 1676
rect 2321 1642 2327 1676
rect 2281 1604 2327 1642
rect 2281 1570 2287 1604
rect 2321 1570 2327 1604
rect 2281 1532 2327 1570
rect 2281 1498 2287 1532
rect 2321 1498 2327 1532
rect 2281 1460 2327 1498
rect 2281 1426 2287 1460
rect 2321 1426 2327 1460
rect 2281 1388 2327 1426
rect 2281 1354 2287 1388
rect 2321 1354 2327 1388
rect 2281 1316 2327 1354
rect 2281 1282 2287 1316
rect 2321 1282 2327 1316
rect 2281 1270 2327 1282
rect 2408 1820 2454 1873
rect 2408 1786 2414 1820
rect 2448 1786 2454 1820
rect 2408 1748 2454 1786
rect 2408 1714 2414 1748
rect 2448 1714 2454 1748
rect 2408 1676 2454 1714
rect 2408 1642 2414 1676
rect 2448 1642 2454 1676
rect 2408 1604 2454 1642
rect 2408 1570 2414 1604
rect 2448 1570 2454 1604
rect 2408 1532 2454 1570
rect 2408 1498 2414 1532
rect 2448 1498 2454 1532
rect 2408 1460 2454 1498
rect 2408 1426 2414 1460
rect 2448 1426 2454 1460
rect 2408 1388 2454 1426
rect 2408 1354 2414 1388
rect 2448 1354 2454 1388
rect 2408 1316 2454 1354
rect 2408 1282 2414 1316
rect 2448 1282 2454 1316
rect 2408 1083 2454 1282
rect 2564 1820 2610 1995
tri 2610 1992 2613 1995 nw
tri 3052 1992 3055 1995 ne
rect 3055 1992 3249 1995
tri 3055 1989 3058 1992 ne
rect 2685 1937 2691 1989
rect 2743 1983 2755 1989
rect 2807 1983 2994 1989
rect 2743 1949 2751 1983
rect 2807 1949 2850 1983
rect 2884 1949 2948 1983
rect 2982 1949 2994 1983
rect 2743 1937 2755 1949
rect 2807 1943 2994 1949
rect 3058 1983 3249 1992
rect 3058 1949 3070 1983
rect 3104 1949 3168 1983
rect 3202 1949 3249 1983
rect 3058 1943 3249 1949
rect 3301 1943 3313 1995
rect 3365 1943 3371 1995
rect 3514 1965 3520 1999
rect 3554 1965 3560 1999
rect 3514 1953 3560 1965
rect 2807 1937 2813 1943
tri 2813 1937 2819 1943 nw
rect 2564 1786 2570 1820
rect 2604 1786 2610 1820
rect 2564 1748 2610 1786
rect 2564 1714 2570 1748
rect 2604 1714 2610 1748
rect 2564 1676 2610 1714
rect 2564 1642 2570 1676
rect 2604 1642 2610 1676
rect 2564 1604 2610 1642
rect 2564 1570 2570 1604
rect 2604 1570 2610 1604
rect 2564 1532 2610 1570
rect 2564 1498 2570 1532
rect 2604 1498 2610 1532
rect 2564 1460 2610 1498
rect 2564 1426 2570 1460
rect 2604 1426 2610 1460
rect 2564 1388 2610 1426
rect 2564 1354 2570 1388
rect 2604 1354 2610 1388
rect 2564 1316 2610 1354
rect 2564 1282 2570 1316
rect 2604 1282 2610 1316
rect 2564 1270 2610 1282
rect 2691 1873 2737 1885
rect 2691 1839 2697 1873
rect 2731 1839 2737 1873
rect 2691 1801 2737 1839
rect 2691 1767 2697 1801
rect 2731 1767 2737 1801
rect 2691 1729 2737 1767
rect 2691 1695 2697 1729
rect 2731 1695 2737 1729
rect 2844 1873 2896 1885
rect 2844 1839 2853 1873
rect 2887 1839 2896 1873
rect 2844 1836 2896 1839
rect 2844 1772 2853 1784
rect 2887 1772 2896 1784
rect 2844 1714 2853 1720
tri 2844 1711 2847 1714 ne
rect 2691 1657 2737 1695
rect 2691 1623 2697 1657
rect 2731 1623 2737 1657
rect 2691 1585 2737 1623
rect 2691 1551 2697 1585
rect 2731 1551 2737 1585
rect 2691 1513 2737 1551
rect 2691 1479 2697 1513
rect 2731 1479 2737 1513
rect 2691 1441 2737 1479
rect 2691 1407 2697 1441
rect 2731 1407 2737 1441
rect 2691 1369 2737 1407
rect 2691 1335 2697 1369
rect 2731 1335 2737 1369
rect 2691 1297 2737 1335
rect 2691 1263 2697 1297
rect 2731 1263 2737 1297
rect 2691 1225 2737 1263
rect 2691 1191 2697 1225
rect 2731 1191 2737 1225
rect 2691 1153 2737 1191
rect 2691 1119 2697 1153
rect 2731 1119 2737 1153
rect 2691 1083 2737 1119
rect 2847 1695 2853 1714
rect 2887 1714 2896 1720
rect 2887 1695 2893 1714
tri 2893 1711 2896 1714 nw
rect 3003 1873 3049 1885
rect 3003 1839 3009 1873
rect 3043 1839 3049 1873
rect 3003 1801 3049 1839
rect 3003 1767 3009 1801
rect 3043 1767 3049 1801
rect 3003 1729 3049 1767
rect 2847 1657 2893 1695
rect 2847 1623 2853 1657
rect 2887 1623 2893 1657
rect 2847 1585 2893 1623
rect 2847 1551 2853 1585
rect 2887 1551 2893 1585
rect 2847 1513 2893 1551
rect 2847 1479 2853 1513
rect 2887 1479 2893 1513
rect 2847 1441 2893 1479
rect 2847 1407 2853 1441
rect 2887 1407 2893 1441
rect 2847 1369 2893 1407
rect 2847 1335 2853 1369
rect 2887 1335 2893 1369
rect 2847 1297 2893 1335
rect 2847 1263 2853 1297
rect 2887 1263 2893 1297
rect 2847 1225 2893 1263
rect 2847 1191 2853 1225
rect 2887 1191 2893 1225
rect 2847 1153 2893 1191
rect 2847 1119 2853 1153
rect 2887 1119 2893 1153
rect 1848 1041 1854 1075
rect 1888 1041 1894 1075
rect 1848 1003 1894 1041
rect 1848 969 1854 1003
rect 1888 969 1894 1003
rect 1848 931 1894 969
rect 1848 897 1854 931
rect 1888 897 1894 931
rect 1848 885 1894 897
rect 2122 1077 2174 1083
rect 2122 1013 2174 1025
rect 2122 949 2174 961
rect 2122 891 2174 897
rect 2404 1077 2456 1083
rect 2404 1013 2456 1025
rect 2404 949 2456 961
rect 2404 891 2456 897
rect 2688 1081 2740 1083
rect 2688 1077 2697 1081
rect 2731 1077 2740 1081
rect 2688 1013 2740 1025
rect 2688 949 2740 961
rect 2688 891 2740 897
rect 2847 1081 2893 1119
rect 3003 1695 3009 1729
rect 3043 1695 3049 1729
rect 3156 1873 3208 1885
rect 3156 1839 3165 1873
rect 3199 1839 3208 1873
rect 3156 1836 3208 1839
rect 3156 1772 3165 1784
rect 3199 1772 3208 1784
rect 3156 1714 3165 1720
tri 3156 1711 3159 1714 ne
rect 3003 1657 3049 1695
rect 3003 1623 3009 1657
rect 3043 1623 3049 1657
rect 3003 1585 3049 1623
rect 3003 1551 3009 1585
rect 3043 1551 3049 1585
rect 3003 1513 3049 1551
rect 3003 1479 3009 1513
rect 3043 1479 3049 1513
rect 3003 1441 3049 1479
rect 3003 1407 3009 1441
rect 3043 1407 3049 1441
rect 3003 1369 3049 1407
rect 3003 1335 3009 1369
rect 3043 1335 3049 1369
rect 3003 1297 3049 1335
rect 3003 1263 3009 1297
rect 3043 1263 3049 1297
rect 3003 1225 3049 1263
rect 3003 1191 3009 1225
rect 3043 1191 3049 1225
rect 3003 1153 3049 1191
rect 3003 1119 3009 1153
rect 3043 1119 3049 1153
rect 2847 1047 2853 1081
rect 2887 1047 2893 1081
rect 2847 1009 2893 1047
rect 2847 975 2853 1009
rect 2887 975 2893 1009
rect 2847 937 2893 975
rect 2847 903 2853 937
rect 2887 903 2893 937
rect 2847 891 2893 903
tri 3000 1083 3003 1086 se
rect 3003 1083 3049 1119
rect 3159 1695 3165 1714
rect 3199 1714 3208 1720
rect 3199 1695 3205 1714
tri 3205 1711 3208 1714 nw
rect 3315 1873 3512 1885
rect 3315 1839 3321 1873
rect 3355 1839 3512 1873
rect 3315 1835 3512 1839
rect 3315 1801 3446 1835
rect 3480 1801 3512 1835
rect 3315 1767 3321 1801
rect 3355 1767 3512 1801
rect 3315 1763 3512 1767
rect 3315 1729 3446 1763
rect 3480 1729 3512 1763
rect 3159 1657 3205 1695
rect 3159 1623 3165 1657
rect 3199 1623 3205 1657
rect 3159 1585 3205 1623
rect 3159 1551 3165 1585
rect 3199 1551 3205 1585
rect 3159 1513 3205 1551
rect 3159 1479 3165 1513
rect 3199 1479 3205 1513
rect 3159 1441 3205 1479
rect 3159 1407 3165 1441
rect 3199 1407 3205 1441
rect 3159 1369 3205 1407
rect 3159 1335 3165 1369
rect 3199 1335 3205 1369
rect 3159 1297 3205 1335
rect 3159 1263 3165 1297
rect 3199 1263 3205 1297
rect 3159 1225 3205 1263
rect 3159 1191 3165 1225
rect 3199 1191 3205 1225
rect 3159 1153 3205 1191
rect 3159 1119 3165 1153
rect 3199 1119 3205 1153
tri 3049 1083 3052 1086 sw
rect 3000 1081 3052 1083
rect 3000 1077 3009 1081
rect 3043 1077 3052 1081
rect 3000 1013 3052 1025
rect 3000 949 3052 961
rect 3000 891 3052 897
rect 3159 1081 3205 1119
rect 3159 1047 3165 1081
rect 3199 1047 3205 1081
rect 3159 1009 3205 1047
rect 3159 975 3165 1009
rect 3199 975 3205 1009
rect 3159 937 3205 975
rect 3159 903 3165 937
rect 3199 903 3205 937
rect 3315 1695 3321 1729
rect 3355 1695 3512 1729
rect 3315 1691 3512 1695
rect 3315 1657 3446 1691
rect 3480 1657 3512 1691
rect 3315 1623 3321 1657
rect 3355 1623 3512 1657
rect 3315 1619 3512 1623
rect 3315 1585 3446 1619
rect 3480 1585 3512 1619
rect 3315 1551 3321 1585
rect 3355 1551 3512 1585
rect 3315 1547 3512 1551
rect 3315 1513 3446 1547
rect 3480 1513 3512 1547
rect 3315 1479 3321 1513
rect 3355 1479 3512 1513
rect 3315 1475 3512 1479
rect 3315 1441 3446 1475
rect 3480 1441 3512 1475
rect 3315 1407 3321 1441
rect 3355 1407 3512 1441
rect 3315 1403 3512 1407
rect 3315 1369 3446 1403
rect 3480 1369 3512 1403
rect 3315 1335 3321 1369
rect 3355 1335 3512 1369
rect 3315 1331 3512 1335
rect 3315 1297 3446 1331
rect 3480 1297 3512 1331
rect 3315 1263 3321 1297
rect 3355 1263 3512 1297
rect 3315 1225 3512 1263
rect 3315 1191 3321 1225
rect 3355 1191 3512 1225
rect 3315 1153 3512 1191
rect 3315 1119 3321 1153
rect 3355 1119 3512 1153
rect 3315 1081 3512 1119
rect 3315 1077 3321 1081
rect 3355 1077 3512 1081
rect 3367 1025 3436 1077
rect 3488 1025 3512 1077
rect 3315 1013 3512 1025
rect 3367 1001 3512 1013
rect 3367 961 3436 1001
rect 3315 949 3436 961
rect 3488 949 3512 1001
tri 3288 903 3315 930 se
rect 3367 924 3512 949
rect 3159 891 3205 903
tri 3281 896 3288 903 se
rect 3288 897 3315 903
rect 3367 897 3436 924
rect 3288 896 3436 897
tri 3276 891 3281 896 se
rect 3281 891 3436 896
tri 3270 885 3276 891 se
rect 3276 885 3436 891
tri 3239 854 3270 885 se
rect 3270 872 3436 885
rect 3488 872 3512 924
rect 3270 854 3512 872
tri 3226 841 3239 854 se
rect 3239 847 3512 854
rect 3239 841 3436 847
rect 138 832 169 841
rect 221 832 234 841
rect 286 832 299 841
rect 138 798 150 832
rect 221 798 223 832
rect 286 798 296 832
rect 138 789 169 798
rect 221 789 234 798
rect 286 789 299 798
rect 351 789 363 841
rect 415 789 427 841
rect 479 789 491 841
rect 543 832 555 841
rect 607 832 619 841
rect 671 832 683 841
rect 735 832 747 841
rect 799 832 811 841
rect 863 832 875 841
rect 547 798 555 832
rect 799 798 801 832
rect 863 798 873 832
rect 543 789 555 798
rect 607 789 619 798
rect 671 789 683 798
rect 735 789 747 798
rect 799 789 811 798
rect 863 789 875 798
rect 927 789 939 841
rect 991 789 1003 841
rect 1055 789 1067 841
rect 1119 832 1131 841
rect 1183 832 1195 841
rect 1247 832 1259 841
rect 1311 832 1323 841
rect 1375 832 1387 841
rect 1439 832 1451 841
rect 1123 798 1131 832
rect 1375 798 1377 832
rect 1439 798 1449 832
rect 1119 789 1131 798
rect 1183 789 1195 798
rect 1247 789 1259 798
rect 1311 789 1323 798
rect 1375 789 1387 798
rect 1439 789 1451 798
rect 1503 789 1515 841
rect 1567 789 1579 841
rect 1631 789 1643 841
rect 1695 832 1707 841
rect 1759 832 1771 841
rect 1823 832 1835 841
rect 1887 832 1899 841
rect 1951 832 1963 841
rect 2015 832 2027 841
rect 1699 798 1707 832
rect 1951 798 1953 832
rect 2015 798 2025 832
rect 1695 789 1707 798
rect 1759 789 1771 798
rect 1823 789 1835 798
rect 1887 789 1899 798
rect 1951 789 1963 798
rect 2015 789 2027 798
rect 2079 789 2091 841
rect 2143 789 2155 841
rect 2207 789 2219 841
rect 2271 832 2283 841
rect 2335 832 2347 841
rect 2399 832 2411 841
rect 2463 832 2475 841
rect 2527 832 2539 841
rect 2591 832 2603 841
rect 2275 798 2283 832
rect 2527 798 2529 832
rect 2591 798 2601 832
rect 2271 789 2283 798
rect 2335 789 2347 798
rect 2399 789 2411 798
rect 2463 789 2475 798
rect 2527 789 2539 798
rect 2591 789 2603 798
rect 2655 789 2667 841
rect 2719 789 2731 841
rect 2783 789 2795 841
rect 2847 832 2859 841
rect 2911 832 2923 841
rect 2975 832 2987 841
rect 3039 832 3051 841
rect 3103 832 3115 841
rect 3167 832 3179 841
rect 2851 798 2859 832
rect 3103 798 3105 832
rect 3167 798 3177 832
rect 2847 789 2859 798
rect 2911 789 2923 798
rect 2975 789 2987 798
rect 3039 789 3051 798
rect 3103 789 3115 798
rect 3167 789 3179 798
rect 3231 789 3243 841
rect 3295 789 3307 841
rect 3359 795 3436 841
rect 3488 795 3512 847
rect 3359 789 3512 795
tri 3212 778 3223 789 ne
rect 3223 778 3512 789
tri 3223 744 3257 778 ne
rect 3257 750 3512 778
rect 3596 1835 3642 2322
rect 3945 1967 4075 2335
rect 4119 2375 4187 2407
tri 4283 2380 4312 2409 ne
rect 4312 2380 4323 2409
tri 4187 2375 4192 2380 sw
tri 4312 2375 4317 2380 ne
rect 4317 2375 4323 2380
rect 4357 2375 4363 2409
rect 4119 2365 4192 2375
rect 4119 2331 4125 2365
rect 4159 2363 4192 2365
tri 4192 2363 4204 2375 sw
rect 4317 2363 4363 2375
rect 4159 2353 4204 2363
tri 4204 2353 4214 2363 sw
rect 4159 2331 4214 2353
tri 4214 2331 4236 2353 sw
rect 4119 2328 4236 2331
tri 4236 2328 4239 2331 sw
rect 4119 2295 4239 2328
tri 4239 2295 4272 2328 sw
rect 4119 2289 4332 2295
rect 4119 2255 4197 2289
rect 4231 2255 4286 2289
rect 4320 2255 4332 2289
rect 4119 2249 4332 2255
rect 4119 2230 4253 2249
tri 4253 2230 4272 2249 nw
tri 4119 2220 4129 2230 ne
rect 4129 2220 4243 2230
tri 4243 2220 4253 2230 nw
tri 4129 2208 4141 2220 ne
rect 4141 2208 4231 2220
tri 4231 2208 4243 2220 nw
rect 3945 1933 3957 1967
rect 3991 1933 4029 1967
rect 4063 1933 4075 1967
rect 3945 1927 4075 1933
tri 3945 1923 3949 1927 ne
rect 3949 1923 4054 1927
tri 3949 1916 3956 1923 ne
rect 3956 1916 4054 1923
tri 3956 1894 3978 1916 ne
rect 3978 1894 4054 1916
tri 4054 1906 4075 1927 nw
tri 3978 1885 3987 1894 ne
rect 3987 1885 4054 1894
tri 3987 1876 3996 1885 ne
rect 3883 1842 3929 1845
rect 3596 1801 3602 1835
rect 3636 1801 3642 1835
rect 3596 1763 3642 1801
rect 3596 1729 3602 1763
rect 3636 1729 3642 1763
rect 3596 1691 3642 1729
rect 3879 1836 3931 1842
rect 3879 1772 3931 1784
rect 3879 1714 3931 1720
rect 3596 1657 3602 1691
rect 3636 1657 3642 1691
rect 3596 1619 3642 1657
rect 3596 1585 3602 1619
rect 3636 1585 3642 1619
rect 3596 1547 3642 1585
rect 3596 1513 3602 1547
rect 3636 1513 3642 1547
rect 3596 1475 3642 1513
rect 3596 1441 3602 1475
rect 3636 1441 3642 1475
rect 3596 1403 3642 1441
rect 3596 1369 3602 1403
rect 3636 1369 3642 1403
rect 3596 1331 3642 1369
rect 3596 1297 3602 1331
rect 3636 1297 3642 1331
rect 3257 744 3523 750
tri 3257 738 3263 744 ne
rect 3263 738 3523 744
tri 3263 724 3277 738 ne
rect 3277 724 3318 738
tri -929 704 -919 714 ne
rect -919 704 -873 714
tri -873 704 -853 724 sw
tri 3277 722 3279 724 ne
rect 3279 722 3318 724
rect 2687 716 2739 722
tri -919 683 -898 704 ne
rect -898 683 -853 704
tri -853 683 -832 704 sw
rect 3000 716 3052 722
tri -898 680 -895 683 ne
rect -895 680 -832 683
tri -832 680 -829 683 sw
tri -895 674 -889 680 ne
rect -889 674 1291 680
rect 1343 674 1372 680
rect 1424 674 2159 680
tri -889 658 -873 674 ne
rect -873 658 169 674
tri -873 640 -855 658 ne
rect -855 640 169 658
rect 203 640 241 674
rect 275 640 313 674
rect 347 640 385 674
rect 419 640 457 674
rect 491 640 529 674
rect 563 640 601 674
rect 635 640 673 674
rect 707 640 745 674
rect 779 640 817 674
rect 851 640 889 674
rect 923 640 961 674
rect 995 640 1033 674
rect 1067 640 1105 674
rect 1139 640 1177 674
rect 1211 640 1249 674
rect 1283 640 1291 674
rect 1355 640 1372 674
rect 1427 640 1465 674
rect 1499 640 1537 674
rect 1571 640 1609 674
rect 1643 640 1681 674
rect 1715 640 1753 674
rect 1787 640 1825 674
rect 1859 640 1897 674
rect 1931 640 1969 674
rect 2003 640 2041 674
rect 2075 640 2113 674
rect 2147 640 2159 674
tri -855 635 -850 640 ne
rect -850 635 1291 640
tri -850 634 -849 635 ne
rect -849 634 1291 635
tri 1279 628 1285 634 ne
rect 1285 628 1291 634
rect 1343 628 1372 640
rect 1424 634 2159 640
rect 2687 652 2697 664
rect 2731 652 2739 664
rect 1424 628 1430 634
tri 1430 628 1436 634 nw
rect 2186 612 2232 624
rect 2186 578 2192 612
rect 2226 611 2232 612
tri 2232 611 2245 624 sw
rect 2226 594 2245 611
tri 2245 594 2262 611 sw
rect 2687 594 2697 600
rect 2226 578 2262 594
rect 2186 577 2262 578
tri 2262 577 2279 594 sw
tri 2687 590 2691 594 ne
rect 2691 577 2697 594
rect 2731 594 2739 600
rect 2731 577 2737 594
tri 2737 592 2739 594 nw
rect 2847 683 2893 695
rect 2847 649 2853 683
rect 2887 649 2893 683
rect 2847 611 2893 649
rect 60 515 66 567
rect 118 515 130 567
rect 182 515 840 567
rect 2186 555 2279 577
tri 2279 555 2301 577 sw
rect 2186 540 2465 555
rect 2186 506 2192 540
rect 2226 539 2465 540
tri 2465 539 2481 555 sw
rect 2691 539 2737 577
rect 2847 577 2853 611
rect 2887 577 2893 611
tri 3279 704 3297 722 ne
rect 3297 704 3318 722
rect 3352 704 3400 738
rect 3434 704 3482 738
rect 3516 704 3523 738
tri 3297 695 3306 704 ne
rect 3306 695 3523 704
rect 3000 652 3009 664
rect 3043 652 3052 664
rect 3000 577 3009 600
rect 3043 577 3052 600
rect 2847 575 2893 577
tri 2893 575 2895 577 sw
tri 2827 555 2847 575 se
rect 2847 555 2895 575
tri 2811 539 2827 555 se
rect 2827 539 2895 555
tri 2895 539 2931 575 sw
rect 3000 539 3052 577
rect 3159 683 3205 695
tri 3306 690 3311 695 ne
rect 3159 649 3165 683
rect 3199 649 3205 683
rect 3159 611 3205 649
rect 3159 577 3165 611
rect 3199 577 3205 611
rect 3159 557 3205 577
rect 3311 635 3523 695
rect 3311 601 3318 635
rect 3352 601 3400 635
rect 3434 601 3482 635
rect 3516 601 3523 635
tri 3205 557 3219 571 sw
tri 3141 539 3159 557 se
rect 3159 539 3219 557
rect 2226 535 2481 539
tri 2481 535 2485 539 sw
rect 2226 506 2485 535
rect 2186 505 2485 506
tri 2485 505 2515 535 sw
rect 2691 505 2697 539
rect 2731 505 2737 539
rect 2186 499 2515 505
tri 2515 499 2521 505 sw
rect 2186 494 2232 499
tri 2232 494 2237 499 nw
tri 2389 494 2394 499 ne
rect 2394 494 2521 499
tri 2521 494 2526 499 sw
tri 2394 450 2438 494 ne
rect 2438 483 2526 494
tri 2526 483 2537 494 sw
rect 2691 493 2737 505
tri 2807 535 2811 539 se
rect 2811 535 2853 539
rect 2887 535 2931 539
tri 2931 535 2935 539 sw
rect 2807 483 2813 535
rect 2865 483 2877 505
rect 2929 483 2935 535
rect 3000 505 3009 539
rect 3043 505 3052 539
rect 3000 493 3052 505
tri 3137 535 3141 539 se
rect 3141 535 3165 539
rect 3199 535 3219 539
tri 3219 535 3241 557 sw
rect 3137 483 3143 535
rect 3199 505 3207 535
rect 3195 483 3207 505
rect 3259 483 3265 535
rect 3311 533 3523 601
rect 3311 499 3318 533
rect 3352 499 3400 533
rect 3434 499 3482 533
rect 3516 499 3523 533
rect 3311 487 3523 499
tri 3587 487 3596 496 se
rect 3596 487 3642 1297
rect 3883 1689 3929 1714
rect 3883 1655 3889 1689
rect 3923 1655 3929 1689
tri 3829 1229 3883 1283 se
rect 3883 1229 3929 1655
rect 3801 1177 3807 1229
rect 3859 1177 3871 1229
rect 3923 1177 3929 1229
rect 3700 1082 3938 1094
rect 3700 1048 3706 1082
rect 3740 1072 3802 1082
rect 3836 1072 3898 1082
rect 3700 1020 3709 1048
rect 3761 1020 3793 1072
rect 3845 1020 3877 1072
rect 3932 1048 3938 1082
rect 3929 1020 3938 1048
rect 3700 1006 3938 1020
rect 3700 972 3706 1006
rect 3740 1000 3802 1006
rect 3836 1000 3898 1006
rect 3700 948 3709 972
rect 3761 948 3793 1000
rect 3845 948 3877 1000
rect 3932 972 3938 1006
rect 3929 948 3938 972
rect 3700 930 3938 948
rect 3700 896 3706 930
rect 3740 928 3802 930
rect 3836 928 3898 930
rect 3700 876 3709 896
rect 3761 876 3793 928
rect 3845 876 3877 928
rect 3932 896 3938 930
rect 3929 876 3938 896
rect 3700 856 3938 876
rect 3700 854 3709 856
rect 3700 820 3706 854
rect 3700 804 3709 820
rect 3761 804 3793 856
rect 3845 804 3877 856
rect 3929 854 3938 856
rect 3932 820 3938 854
rect 3929 804 3938 820
rect 3700 778 3938 804
rect 3700 744 3706 778
rect 3740 744 3802 778
rect 3836 744 3898 778
rect 3932 744 3938 778
rect 3700 732 3938 744
tri 3918 630 3996 708 se
rect 3996 688 4054 1885
tri 4119 1845 4141 1867 se
rect 4141 1845 4187 2208
tri 4187 2164 4231 2208 nw
tri 4330 1995 4394 2059 se
rect 4394 2039 4440 2579
rect 4522 3545 4528 3579
rect 4562 3545 4568 3579
rect 4522 3505 4568 3545
rect 4522 3471 4528 3505
rect 4562 3471 4568 3505
rect 4522 3431 4568 3471
rect 4522 3397 4528 3431
rect 4562 3397 4568 3431
rect 4522 3357 4568 3397
rect 4522 3323 4528 3357
rect 4562 3323 4568 3357
rect 4522 3283 4568 3323
rect 4522 3249 4528 3283
rect 4562 3249 4568 3283
rect 4522 3209 4568 3249
rect 4522 3175 4528 3209
rect 4562 3175 4568 3209
rect 4522 3135 4568 3175
rect 4522 3101 4528 3135
rect 4562 3101 4568 3135
rect 4522 3061 4568 3101
rect 4522 3027 4528 3061
rect 4562 3027 4568 3061
rect 4712 3644 4718 3678
rect 4752 3644 4802 3678
rect 4836 3644 4886 3678
rect 4920 3644 4926 3678
rect 4712 3603 4926 3644
rect 4712 3569 4718 3603
rect 4752 3569 4802 3603
rect 4836 3569 4886 3603
rect 4920 3569 4926 3603
rect 4712 3528 4926 3569
rect 4712 3494 4718 3528
rect 4752 3494 4802 3528
rect 4836 3494 4886 3528
rect 4920 3494 4926 3528
rect 4712 3453 4926 3494
rect 4712 3419 4718 3453
rect 4752 3419 4802 3453
rect 4836 3419 4886 3453
rect 4920 3419 4926 3453
rect 4712 3378 4926 3419
rect 4712 3344 4718 3378
rect 4752 3344 4802 3378
rect 4836 3344 4886 3378
rect 4920 3344 4926 3378
rect 4712 3303 4926 3344
rect 4712 3269 4718 3303
rect 4752 3269 4802 3303
rect 4836 3269 4886 3303
rect 4920 3269 4926 3303
rect 4712 3235 4926 3269
rect 4712 3183 4715 3235
rect 4767 3183 4793 3235
rect 4845 3183 4871 3235
rect 4923 3183 4926 3235
rect 4712 3153 4926 3183
rect 4712 3125 4718 3153
rect 4752 3125 4802 3153
rect 4836 3125 4886 3153
rect 4920 3125 4926 3153
rect 4712 3073 4715 3125
rect 4767 3073 4793 3125
rect 4845 3073 4871 3125
rect 4923 3073 4926 3125
rect 4712 3044 4718 3073
rect 4752 3044 4802 3073
rect 4836 3044 4886 3073
rect 4920 3044 4926 3073
rect 4522 2987 4568 3027
rect 4522 2953 4528 2987
rect 4562 2953 4568 2987
rect 4522 2912 4568 2953
rect 4522 2878 4528 2912
rect 4562 2878 4568 2912
rect 4522 2837 4568 2878
rect 4522 2803 4528 2837
rect 4562 2803 4568 2837
rect 4522 2762 4568 2803
rect 4522 2728 4528 2762
rect 4562 2728 4568 2762
rect 4522 2687 4568 2728
rect 4522 2653 4528 2687
rect 4562 2653 4568 2687
rect 4522 2612 4568 2653
rect 4522 2578 4528 2612
rect 4562 2578 4568 2612
rect 4522 2537 4568 2578
rect 4522 2503 4528 2537
rect 4562 2503 4568 2537
rect 4522 2462 4568 2503
rect 4522 2428 4528 2462
rect 4562 2428 4568 2462
rect 4522 2387 4568 2428
rect 4522 2353 4528 2387
rect 4562 2353 4568 2387
rect 4522 2341 4568 2353
rect 4620 3031 4672 3037
rect 4620 2967 4672 2979
tri 4613 2132 4620 2139 se
rect 4620 2132 4672 2915
rect 4712 3003 4926 3044
rect 4712 2969 4718 3003
rect 4752 2969 4802 3003
rect 4836 2969 4886 3003
rect 4920 2969 4926 3003
rect 4712 2928 4926 2969
rect 4712 2894 4718 2928
rect 4752 2894 4802 2928
rect 4836 2894 4886 2928
rect 4920 2894 4926 2928
rect 4712 2853 4926 2894
rect 4712 2819 4718 2853
rect 4752 2819 4802 2853
rect 4836 2819 4886 2853
rect 4920 2819 4926 2853
rect 4712 2778 4926 2819
rect 4712 2744 4718 2778
rect 4752 2744 4802 2778
rect 4836 2744 4886 2778
rect 4920 2744 4926 2778
rect 4712 2703 4926 2744
rect 4712 2669 4718 2703
rect 4752 2669 4802 2703
rect 4836 2669 4886 2703
rect 4920 2669 4926 2703
rect 4712 2628 4926 2669
rect 4712 2594 4718 2628
rect 4752 2594 4802 2628
rect 4836 2594 4886 2628
rect 4920 2594 4926 2628
rect 4712 2553 4926 2594
rect 4712 2519 4718 2553
rect 4752 2519 4802 2553
rect 4836 2519 4886 2553
rect 4920 2519 4926 2553
rect 4712 2478 4926 2519
rect 4712 2444 4718 2478
rect 4752 2444 4802 2478
rect 4836 2444 4886 2478
rect 4920 2444 4926 2478
rect 4712 2403 4926 2444
rect 5091 3653 5591 3705
rect 5091 3619 5173 3653
rect 5207 3619 5249 3653
rect 5283 3619 5325 3653
rect 5359 3619 5402 3653
rect 5436 3619 5479 3653
rect 5513 3619 5591 3653
rect 5091 3610 5591 3619
rect 5091 3594 5333 3610
tri 5333 3594 5349 3610 nw
tri 5452 3594 5468 3610 ne
rect 5468 3594 5591 3610
rect 5091 3581 5320 3594
tri 5320 3581 5333 3594 nw
tri 5468 3581 5481 3594 ne
rect 5481 3581 5591 3594
rect 5091 3547 5097 3581
rect 5131 3547 5286 3581
tri 5286 3547 5320 3581 nw
tri 5481 3547 5515 3581 ne
rect 5515 3547 5551 3581
rect 5585 3547 5591 3581
rect 5091 3505 5256 3547
tri 5256 3517 5286 3547 nw
tri 5515 3517 5545 3547 ne
rect 5091 3471 5097 3505
rect 5131 3471 5256 3505
rect 5545 3509 5591 3547
rect 5545 3475 5551 3509
rect 5585 3475 5591 3509
rect 5091 3462 5256 3471
rect 5091 3429 5216 3462
rect 5091 3395 5097 3429
rect 5131 3428 5216 3429
rect 5250 3428 5256 3462
rect 5131 3395 5256 3428
rect 5091 3390 5256 3395
rect 5091 3356 5216 3390
rect 5250 3356 5256 3390
rect 5091 3353 5256 3356
rect 5091 3319 5097 3353
rect 5131 3335 5256 3353
rect 5426 3462 5472 3474
rect 5426 3428 5432 3462
rect 5466 3428 5472 3462
rect 5426 3390 5472 3428
rect 5426 3356 5432 3390
rect 5466 3356 5472 3390
tri 5256 3335 5258 3337 sw
rect 5131 3331 5258 3335
tri 5258 3331 5262 3335 sw
tri 5422 3331 5426 3335 se
rect 5426 3331 5472 3356
rect 5131 3319 5262 3331
rect 5091 3318 5262 3319
tri 5262 3318 5275 3331 sw
tri 5409 3318 5422 3331 se
rect 5422 3318 5472 3331
rect 5091 3284 5216 3318
rect 5250 3292 5275 3318
tri 5275 3292 5301 3318 sw
tri 5383 3292 5409 3318 se
rect 5409 3292 5432 3318
rect 5250 3284 5432 3292
rect 5466 3284 5472 3318
rect 5091 3277 5472 3284
rect 5091 3243 5097 3277
rect 5131 3243 5472 3277
rect 5091 3217 5472 3243
rect 5091 3201 5327 3217
rect 5091 3167 5097 3201
rect 5131 3183 5327 3201
rect 5361 3183 5472 3217
rect 5131 3167 5472 3183
rect 5091 3145 5472 3167
rect 5091 3125 5327 3145
rect 5091 3091 5097 3125
rect 5131 3111 5327 3125
rect 5361 3111 5472 3145
rect 5131 3099 5472 3111
rect 5545 3437 5591 3475
rect 5545 3403 5551 3437
rect 5585 3403 5591 3437
rect 5545 3365 5591 3403
rect 5545 3331 5551 3365
rect 5585 3331 5591 3365
rect 5545 3293 5591 3331
rect 5545 3259 5551 3293
rect 5585 3259 5591 3293
rect 5545 3220 5591 3259
rect 5545 3186 5551 3220
rect 5585 3186 5591 3220
rect 5545 3147 5591 3186
rect 5545 3113 5551 3147
rect 5585 3113 5591 3147
rect 5131 3091 5301 3099
rect 5091 3075 5301 3091
tri 5301 3075 5325 3099 nw
rect 5091 3074 5300 3075
tri 5300 3074 5301 3075 nw
rect 5545 3074 5591 3113
rect 5091 3049 5266 3074
rect 5091 3015 5097 3049
rect 5131 3040 5266 3049
tri 5266 3040 5300 3074 nw
rect 5545 3040 5551 3074
rect 5585 3040 5591 3074
rect 5131 3035 5261 3040
tri 5261 3035 5266 3040 nw
rect 5131 3031 5257 3035
tri 5257 3031 5261 3035 nw
rect 5426 3031 5478 3037
rect 5131 3015 5256 3031
tri 5256 3030 5257 3031 nw
rect 5091 2973 5256 3015
rect 5091 2939 5097 2973
rect 5131 2956 5256 2973
rect 5131 2939 5216 2956
rect 5091 2922 5216 2939
rect 5250 2922 5256 2956
rect 5426 2967 5478 2979
rect 5091 2897 5256 2922
rect 5091 2863 5097 2897
rect 5131 2884 5256 2897
rect 5131 2863 5216 2884
rect 5091 2850 5216 2863
rect 5250 2850 5256 2884
rect 5091 2821 5256 2850
rect 5091 2787 5097 2821
rect 5131 2812 5256 2821
rect 5321 2942 5373 2948
rect 5321 2878 5373 2890
rect 5321 2814 5373 2826
rect 5426 2909 5478 2915
rect 5426 2884 5472 2909
tri 5472 2903 5478 2909 nw
rect 5545 3001 5591 3040
rect 5545 2967 5551 3001
rect 5585 2967 5591 3001
rect 5545 2928 5591 2967
rect 5426 2850 5432 2884
rect 5466 2850 5472 2884
rect 5131 2787 5216 2812
rect 5091 2778 5216 2787
rect 5250 2778 5256 2812
rect 5091 2757 5256 2778
rect 5426 2812 5472 2850
rect 5426 2778 5432 2812
rect 5466 2778 5472 2812
rect 5426 2766 5472 2778
rect 5545 2894 5551 2928
rect 5585 2894 5591 2928
rect 5545 2855 5591 2894
rect 5545 2821 5551 2855
rect 5585 2821 5591 2855
rect 5545 2782 5591 2821
rect 5091 2748 5192 2757
tri 5192 2748 5201 2757 nw
rect 5545 2748 5551 2782
rect 5585 2748 5591 2782
rect 5091 2745 5163 2748
rect 5091 2711 5097 2745
rect 5131 2719 5163 2745
tri 5163 2719 5192 2748 nw
rect 5545 2719 5591 2748
rect 5732 3676 5778 3724
rect 5732 3642 5738 3676
rect 5772 3642 5778 3676
rect 5732 3594 5778 3642
rect 5732 3560 5738 3594
rect 5772 3560 5778 3594
rect 5732 3512 5778 3560
rect 5732 3478 5738 3512
rect 5772 3478 5778 3512
rect 5732 3429 5778 3478
rect 5732 3395 5738 3429
rect 5772 3395 5778 3429
rect 5732 3383 5778 3395
tri 5778 3383 5931 3536 sw
rect 5732 3367 5931 3383
tri 5931 3367 5947 3383 sw
rect 5732 3342 5947 3367
rect 5732 3308 5738 3342
rect 5772 3317 5947 3342
rect 5772 3308 5829 3317
rect 5863 3308 5901 3317
rect 5935 3308 5947 3317
rect 5732 3256 5733 3308
rect 5785 3256 5811 3308
rect 5863 3256 5889 3308
rect 5941 3256 5947 3308
rect 6567 3358 6770 3366
rect 6567 3306 6568 3358
rect 6620 3306 6640 3358
rect 6692 3306 6712 3358
rect 5732 3231 5738 3256
rect 5772 3231 5947 3256
rect 5732 3220 5947 3231
rect 5732 3168 5733 3220
rect 5785 3168 5811 3220
rect 5863 3168 5889 3220
rect 5941 3168 5947 3220
rect 5732 3153 5738 3168
rect 5772 3153 5947 3168
rect 5732 3132 5947 3153
rect 5732 3080 5733 3132
rect 5785 3080 5811 3132
rect 5863 3080 5889 3132
rect 5941 3080 5947 3132
rect 5732 3075 5738 3080
rect 5772 3075 5947 3080
rect 5732 3031 5947 3075
rect 5732 2997 5738 3031
rect 5772 2997 5947 3031
rect 5732 2953 5947 2997
rect 5732 2919 5738 2953
rect 5772 2919 5947 2953
rect 5732 2875 5947 2919
rect 5732 2841 5738 2875
rect 5772 2841 5947 2875
rect 5732 2840 5947 2841
rect 5732 2806 5829 2840
rect 5863 2806 5901 2840
rect 5935 2806 5947 2840
rect 5732 2797 5947 2806
rect 5732 2763 5738 2797
rect 5772 2763 5947 2797
tri 5591 2719 5595 2723 sw
rect 5732 2719 5947 2763
rect 5131 2711 5153 2719
rect 5091 2709 5153 2711
tri 5153 2709 5163 2719 nw
rect 5545 2717 5595 2719
tri 5595 2717 5597 2719 sw
rect 5545 2711 5597 2717
rect 5091 2669 5137 2709
tri 5137 2693 5153 2709 nw
rect 5091 2635 5097 2669
rect 5131 2635 5137 2669
rect 5091 2593 5137 2635
rect 5206 2622 5212 2674
rect 5264 2622 5276 2674
rect 5328 2666 5363 2674
tri 5363 2666 5371 2674 sw
rect 5328 2664 5371 2666
tri 5371 2664 5373 2666 sw
rect 5328 2656 5373 2664
tri 5373 2656 5381 2664 sw
rect 5328 2641 5381 2656
tri 5381 2641 5396 2656 sw
rect 5545 2647 5597 2659
rect 5328 2622 5396 2641
tri 5396 2622 5415 2641 sw
tri 5349 2607 5364 2622 ne
rect 5364 2607 5415 2622
tri 5415 2607 5430 2622 sw
rect 5091 2559 5097 2593
rect 5131 2559 5137 2593
tri 5364 2590 5381 2607 ne
rect 5381 2590 5430 2607
tri 5430 2590 5447 2607 sw
tri 5381 2587 5384 2590 ne
rect 5384 2587 5447 2590
tri 5447 2587 5450 2590 sw
rect 5545 2589 5597 2595
rect 5732 2685 5738 2719
rect 5772 2685 5947 2719
rect 5732 2641 5947 2685
rect 5732 2607 5738 2641
rect 5772 2607 5947 2641
tri 5384 2573 5398 2587 ne
rect 5398 2573 5450 2587
tri 5450 2573 5464 2587 sw
rect 5732 2575 5947 2607
rect 6026 3282 6072 3294
rect 6026 3248 6032 3282
rect 6066 3248 6072 3282
rect 6026 3210 6072 3248
rect 6026 3176 6032 3210
rect 6066 3176 6072 3210
rect 5091 2517 5137 2559
rect 5204 2521 5210 2573
rect 5262 2521 5274 2573
rect 5326 2524 5332 2573
tri 5398 2564 5407 2573 ne
rect 5407 2567 5464 2573
tri 5464 2567 5470 2573 sw
rect 5407 2564 5470 2567
tri 5470 2564 5473 2567 sw
tri 6023 2564 6026 2567 se
rect 6026 2564 6072 3176
rect 6567 3283 6580 3306
rect 6614 3283 6652 3306
rect 6686 3299 6730 3306
rect 6764 3299 6770 3358
rect 6686 3283 6770 3299
rect 6567 3269 6770 3283
rect 6567 3217 6568 3269
rect 6620 3217 6640 3269
rect 6692 3217 6712 3269
rect 6764 3217 6770 3269
rect 6567 3181 6770 3217
rect 6248 3141 6378 3147
rect 6248 3107 6260 3141
rect 6294 3107 6332 3141
rect 6366 3107 6378 3141
rect 6248 3101 6378 3107
rect 6248 3095 6372 3101
tri 6372 3095 6378 3101 nw
rect 6567 3129 6568 3181
rect 6620 3129 6640 3181
rect 6692 3129 6712 3181
rect 6764 3129 6770 3181
rect 6567 3095 6770 3129
rect 6248 3081 6358 3095
tri 6358 3081 6372 3095 nw
tri 5332 2524 5372 2564 sw
tri 5407 2524 5447 2564 ne
rect 5447 2524 5473 2564
tri 5473 2524 5513 2564 sw
tri 5983 2524 6023 2564 se
rect 6023 2524 6072 2564
rect 5326 2521 5372 2524
rect 5091 2483 5097 2517
rect 5131 2483 5137 2517
tri 5309 2510 5320 2521 ne
rect 5320 2510 5372 2521
tri 5372 2510 5386 2524 sw
tri 5447 2510 5461 2524 ne
rect 5461 2510 6072 2524
tri 5320 2498 5332 2510 ne
rect 5332 2498 5386 2510
rect 5091 2444 5137 2483
tri 5332 2454 5376 2498 ne
rect 5376 2497 5386 2498
tri 5386 2497 5399 2510 sw
tri 5461 2497 5474 2510 ne
rect 5474 2507 6072 2510
rect 5474 2497 6062 2507
tri 6062 2497 6072 2507 nw
rect 6113 3069 6159 3081
rect 6113 3035 6119 3069
rect 6153 3035 6159 3069
rect 6113 2997 6159 3035
rect 6113 2963 6119 2997
rect 6153 2963 6159 2997
rect 5376 2478 5399 2497
tri 5399 2478 5418 2497 sw
tri 5474 2478 5493 2497 ne
rect 5493 2478 6043 2497
tri 6043 2478 6062 2497 nw
tri 6094 2478 6113 2497 se
rect 6113 2478 6159 2963
rect 6248 3061 6338 3081
tri 6338 3061 6358 3081 nw
rect 6567 3061 6730 3095
rect 6764 3061 6770 3095
tri 6221 2779 6248 2806 se
rect 6248 2779 6302 3061
tri 6302 3025 6338 3061 nw
rect 6567 3016 6770 3061
rect 6567 2982 6730 3016
rect 6764 2982 6770 3016
rect 6567 2965 6770 2982
rect 6567 2931 6580 2965
rect 6614 2931 6652 2965
rect 6686 2937 6770 2965
rect 6686 2931 6730 2937
rect 6567 2903 6730 2931
rect 6764 2903 6770 2937
rect 6567 2858 6770 2903
rect 6567 2840 6730 2858
rect 6567 2806 6580 2840
rect 6614 2806 6652 2840
rect 6686 2824 6730 2840
rect 6764 2824 6770 2858
rect 6686 2806 6770 2824
tri 6302 2779 6305 2782 sw
rect 6567 2779 6770 2806
tri 6198 2756 6221 2779 se
rect 6221 2756 6305 2779
tri 6305 2756 6328 2779 sw
rect 6198 2750 6328 2756
rect 6198 2716 6210 2750
rect 6244 2716 6282 2750
rect 6316 2716 6328 2750
rect 6198 2710 6328 2716
rect 6567 2745 6730 2779
rect 6764 2745 6770 2779
rect 6567 2700 6770 2745
rect 6247 2618 6253 2670
rect 6305 2618 6319 2670
rect 6371 2618 6377 2670
rect 6567 2666 6730 2700
rect 6764 2666 6770 2700
rect 6567 2621 6770 2666
rect 6567 2587 6730 2621
rect 6764 2587 6770 2621
rect 6567 2575 6770 2587
rect 5376 2454 5418 2478
tri 5137 2444 5147 2454 sw
tri 5376 2444 5386 2454 ne
rect 5386 2444 5418 2454
tri 5418 2444 5452 2478 sw
tri 6060 2444 6094 2478 se
rect 6094 2477 6159 2478
rect 6094 2444 6126 2477
tri 6126 2444 6159 2477 nw
rect 5091 2441 5147 2444
tri 5063 2407 5091 2435 se
rect 5091 2407 5097 2441
rect 5131 2407 5147 2441
rect 4712 2369 4718 2403
rect 4752 2369 4802 2403
rect 4836 2369 4886 2403
rect 4920 2369 4926 2403
rect 4712 2328 4926 2369
tri 5021 2365 5063 2407 se
rect 5063 2398 5147 2407
tri 5147 2398 5193 2444 sw
tri 5386 2398 5432 2444 ne
rect 5432 2398 6080 2444
tri 6080 2398 6126 2444 nw
rect 5063 2365 5193 2398
tri 4997 2341 5021 2365 se
rect 5021 2341 5097 2365
tri 4987 2331 4997 2341 se
rect 4997 2331 5097 2341
rect 5131 2341 5193 2365
tri 5193 2341 5250 2398 sw
rect 5131 2331 5250 2341
rect 4712 2294 4718 2328
rect 4752 2294 4802 2328
rect 4836 2294 4886 2328
rect 4920 2294 4926 2328
rect 4712 2254 4926 2294
rect 4712 2220 4718 2254
rect 4752 2220 4802 2254
rect 4836 2220 4886 2254
rect 4920 2220 4926 2254
rect 4712 2208 4926 2220
tri 4986 2330 4987 2331 se
rect 4987 2330 5250 2331
rect 4986 2301 5250 2330
tri 5250 2301 5290 2341 sw
rect 4986 2289 5509 2301
rect 5561 2289 5573 2301
rect 4986 2255 5169 2289
rect 5203 2255 5245 2289
rect 5279 2255 5320 2289
rect 5354 2255 5395 2289
rect 5429 2255 5470 2289
rect 5504 2255 5509 2289
rect 4986 2249 5509 2255
rect 5561 2249 5573 2255
rect 5625 2249 5631 2301
rect 4986 2218 5060 2249
tri 5060 2218 5091 2249 nw
tri 4547 2066 4613 2132 se
rect 4613 2117 4672 2132
rect 4613 2066 4621 2117
tri 4621 2066 4672 2117 nw
tri 4920 2066 4986 2132 se
rect 4986 2112 5032 2218
tri 5032 2190 5060 2218 nw
rect 5499 2166 5505 2218
rect 5557 2166 5569 2218
rect 5621 2166 6085 2218
rect 6137 2166 6149 2218
rect 6201 2166 6207 2218
tri 4986 2066 5032 2112 nw
tri 4546 2065 4547 2066 se
rect 4547 2065 4620 2066
tri 4620 2065 4621 2066 nw
tri 4919 2065 4920 2066 se
rect 4394 1995 4396 2039
tri 4396 1995 4440 2039 nw
tri 4481 2000 4546 2065 se
rect 4546 2000 4555 2065
tri 4555 2000 4620 2065 nw
tri 4854 2000 4919 2065 se
rect 4919 2000 4920 2065
tri 4920 2000 4986 2066 nw
tri 4476 1995 4481 2000 se
rect 4481 1995 4550 2000
tri 4550 1995 4555 2000 nw
tri 4849 1995 4854 2000 se
rect 4222 1943 4228 1995
rect 4280 1943 4292 1995
rect 4344 1989 4390 1995
tri 4390 1989 4396 1995 nw
tri 4472 1991 4476 1995 se
rect 4476 1991 4546 1995
tri 4546 1991 4550 1995 nw
tri 4845 1991 4849 1995 se
rect 4849 1991 4854 1995
tri 4470 1989 4472 1991 se
rect 4472 1989 4544 1991
tri 4544 1989 4546 1991 nw
tri 4843 1989 4845 1991 se
rect 4845 1989 4854 1991
rect 4344 1943 4350 1989
tri 4350 1949 4390 1989 nw
tri 4430 1949 4470 1989 se
rect 4470 1949 4498 1989
tri 4424 1943 4430 1949 se
rect 4430 1943 4498 1949
tri 4498 1943 4544 1989 nw
tri 4797 1943 4843 1989 se
rect 4843 1943 4854 1989
tri 4415 1934 4424 1943 se
rect 4424 1934 4489 1943
tri 4489 1934 4498 1943 nw
tri 4788 1934 4797 1943 se
rect 4797 1934 4854 1943
tri 4854 1934 4920 2000 nw
tri 4398 1917 4415 1934 se
rect 4415 1917 4472 1934
tri 4472 1917 4489 1934 nw
tri 4771 1917 4788 1934 se
tri 4387 1906 4398 1917 se
rect 4398 1906 4461 1917
tri 4461 1906 4472 1917 nw
tri 4760 1906 4771 1917 se
rect 4771 1906 4788 1917
tri 4349 1868 4387 1906 se
rect 4387 1868 4423 1906
tri 4423 1868 4461 1906 nw
tri 4722 1868 4760 1906 se
rect 4760 1868 4788 1906
tri 4788 1868 4854 1934 nw
rect 4119 1833 4187 1845
tri 4324 1843 4349 1868 se
rect 4349 1843 4398 1868
tri 4398 1843 4423 1868 nw
tri 4697 1843 4722 1868 se
rect 4119 1799 4125 1833
rect 4159 1799 4187 1833
rect 4119 1761 4187 1799
rect 4119 1727 4125 1761
rect 4159 1727 4187 1761
rect 4119 1689 4187 1727
rect 4119 1655 4125 1689
rect 4159 1655 4187 1689
rect 4119 1643 4187 1655
tri 4289 1808 4324 1843 se
rect 4324 1808 4363 1843
tri 4363 1808 4398 1843 nw
tri 4662 1808 4697 1843 se
rect 4697 1808 4722 1843
rect 4289 1802 4357 1808
tri 4357 1802 4363 1808 nw
tri 4656 1802 4662 1808 se
rect 4662 1802 4722 1808
tri 4722 1802 4788 1868 nw
rect 4289 1666 4341 1802
tri 4341 1786 4357 1802 nw
tri 4640 1786 4656 1802 se
tri 4590 1736 4640 1786 se
rect 4640 1736 4656 1786
tri 4656 1736 4722 1802 nw
tri 4524 1670 4590 1736 se
tri 4590 1670 4656 1736 nw
rect 4289 1602 4341 1614
tri 4458 1604 4524 1670 se
tri 4524 1604 4590 1670 nw
rect 4289 1544 4341 1550
tri 4398 1544 4458 1604 se
tri 4392 1538 4398 1544 se
rect 4398 1538 4458 1544
tri 4458 1538 4524 1604 nw
tri 4326 1472 4392 1538 se
tri 4392 1472 4458 1538 nw
tri 4260 1406 4326 1472 se
tri 4326 1406 4392 1472 nw
tri 4194 1340 4260 1406 se
tri 4260 1340 4326 1406 nw
tri 3996 630 4054 688 nw
tri 4149 1295 4194 1340 se
rect 4194 1295 4215 1340
tri 4215 1295 4260 1340 nw
tri 4111 630 4149 668 se
rect 4149 648 4195 1295
tri 4195 1275 4215 1295 nw
tri 3840 552 3918 630 se
tri 3918 552 3996 630 nw
tri 4083 602 4111 630 se
rect 4111 602 4149 630
tri 4149 602 4195 648 nw
tri 4033 552 4083 602 se
tri 3583 483 3587 487 se
rect 3587 483 3642 487
rect 2438 450 2537 483
tri 2537 450 2570 483 sw
tri 3550 450 3583 483 se
rect 3583 476 3642 483
rect 3583 450 3603 476
tri 2438 444 2444 450 ne
rect 2444 444 2570 450
rect 157 438 2229 444
rect 157 404 169 438
rect 203 404 241 438
rect 275 404 313 438
rect 347 404 385 438
rect 419 404 457 438
rect 491 404 529 438
rect 563 404 601 438
rect 635 404 673 438
rect 707 404 745 438
rect 779 404 817 438
rect 851 404 889 438
rect 923 404 961 438
rect 995 404 1033 438
rect 1067 404 1105 438
rect 1139 404 1177 438
rect 1211 404 1249 438
rect 1283 404 1321 438
rect 1355 404 1393 438
rect 1427 404 1465 438
rect 1499 404 1537 438
rect 1571 404 1609 438
rect 1643 404 1681 438
rect 1715 404 1753 438
rect 1787 404 1825 438
rect 1859 404 1897 438
rect 1931 404 1969 438
rect 2003 404 2041 438
rect 2075 404 2113 438
rect 2147 431 2229 438
tri 2229 431 2242 444 sw
tri 2444 431 2457 444 ne
rect 2457 437 2570 444
tri 2570 437 2583 450 sw
tri 3537 437 3550 450 se
rect 3550 437 3603 450
tri 3603 437 3642 476 nw
tri 3762 474 3840 552 se
tri 3840 474 3918 552 nw
tri 4017 536 4033 552 se
rect 4033 536 4083 552
tri 4083 536 4149 602 nw
tri 3955 474 4017 536 se
tri 3725 437 3762 474 se
rect 3762 437 3770 474
rect 2457 431 2583 437
tri 2583 431 2589 437 sw
rect 2753 431 3557 437
rect 2147 423 2242 431
tri 2242 423 2250 431 sw
tri 2457 423 2465 431 ne
rect 2465 423 2589 431
rect 2147 410 2250 423
tri 2250 410 2263 423 sw
tri 2465 410 2478 423 ne
rect 2478 410 2589 423
rect 2147 404 2263 410
rect 157 398 2263 404
tri 2209 397 2210 398 ne
rect 2210 397 2263 398
tri 2263 397 2276 410 sw
tri 2478 397 2491 410 ne
rect 2491 397 2589 410
tri 2589 397 2623 431 sw
rect 2753 397 2765 431
rect 2799 397 2847 431
rect 2881 397 2929 431
rect 2963 397 3010 431
rect 3044 397 3091 431
rect 3125 397 3557 431
tri 2210 344 2263 397 ne
rect 2263 344 2276 397
tri 2276 344 2329 397 sw
tri 2491 344 2544 397 ne
rect 2544 391 2623 397
tri 2623 391 2629 397 sw
rect 2753 391 3557 397
tri 3557 391 3603 437 nw
tri 3684 396 3725 437 se
rect 3725 404 3770 437
tri 3770 404 3840 474 nw
tri 3951 470 3955 474 se
rect 3955 470 4017 474
tri 4017 470 4083 536 nw
tri 3885 404 3951 470 se
tri 3951 404 4017 470 nw
rect 3725 396 3762 404
tri 3762 396 3770 404 nw
tri 3877 396 3885 404 se
tri 3679 391 3684 396 se
rect 3684 391 3704 396
rect 2544 344 2629 391
tri 2263 320 2287 344 ne
rect 2287 320 2329 344
tri 2329 320 2353 344 sw
tri 2544 320 2568 344 ne
rect 2568 320 2629 344
tri 2629 320 2700 391 sw
tri 3608 320 3679 391 se
rect 3679 338 3704 391
tri 3704 338 3762 396 nw
tri 3819 338 3877 396 se
rect 3877 338 3885 396
tri 3885 338 3951 404 nw
rect 3679 320 3684 338
tri 239 317 242 320 se
rect 242 317 248 320
rect 157 311 248 317
rect 300 311 328 320
rect 380 311 408 320
rect 460 311 488 320
rect 540 317 546 320
tri 546 317 549 320 sw
tri 2287 317 2290 320 ne
rect 2290 318 2353 320
tri 2353 318 2355 320 sw
tri 2568 318 2570 320 ne
rect 2570 318 2700 320
tri 2700 318 2702 320 sw
tri 3606 318 3608 320 se
rect 3608 318 3684 320
tri 3684 318 3704 338 nw
tri 3799 318 3819 338 se
rect 2290 317 2355 318
rect 540 311 2159 317
rect 157 277 169 311
rect 203 277 241 311
rect 300 277 313 311
rect 380 277 385 311
rect 563 277 601 311
rect 635 277 673 311
rect 707 277 745 311
rect 779 277 817 311
rect 851 277 889 311
rect 923 277 961 311
rect 995 277 1033 311
rect 1067 277 1105 311
rect 1139 277 1177 311
rect 1211 277 1249 311
rect 1283 277 1321 311
rect 1355 277 1393 311
rect 1427 277 1465 311
rect 1499 277 1537 311
rect 1571 277 1609 311
rect 1643 277 1681 311
rect 1715 277 1753 311
rect 1787 277 1825 311
rect 1859 277 1897 311
rect 1931 277 1969 311
rect 2003 277 2041 311
rect 2075 277 2113 311
rect 2147 277 2159 311
tri 2290 278 2329 317 ne
rect 2329 278 2355 317
tri 2355 278 2395 318 sw
tri 2570 278 2610 318 ne
rect 2610 278 3628 318
rect 157 271 248 277
tri 239 268 242 271 ne
rect 242 268 248 271
rect 300 268 328 277
rect 380 268 408 277
rect 460 268 488 277
rect 540 271 2159 277
tri 2329 271 2336 278 ne
rect 2336 271 2395 278
rect 540 268 546 271
tri 546 268 549 271 nw
tri 2336 268 2339 271 ne
rect 2339 268 2395 271
tri 2395 268 2405 278 sw
tri 2610 268 2620 278 ne
rect 2620 268 3628 278
tri 2339 220 2387 268 ne
rect 2387 262 2405 268
tri 2405 262 2411 268 sw
tri 2620 262 2626 268 ne
rect 2626 262 3628 268
tri 3628 262 3684 318 nw
tri 3753 272 3799 318 se
rect 3799 272 3819 318
tri 3819 272 3885 338 nw
tri 3743 262 3753 272 se
rect 3753 262 3759 272
rect 2387 220 2411 262
tri 2411 220 2453 262 sw
tri 3701 220 3743 262 se
rect 3743 220 3759 262
tri 2174 208 2186 220 se
rect 2186 208 2232 220
tri 2387 212 2395 220 ne
rect 2395 212 2453 220
tri 2453 212 2461 220 sw
tri 3693 212 3701 220 se
rect 3701 212 3759 220
tri 3759 212 3819 272 nw
tri 2157 191 2174 208 se
rect 2174 191 2192 208
rect 242 139 248 191
rect 300 139 328 191
rect 380 139 408 191
rect 460 139 488 191
rect 540 174 2192 191
rect 2226 174 2232 208
rect 540 139 2232 174
tri 2395 166 2441 212 ne
rect 2441 166 3713 212
tri 3713 166 3759 212 nw
tri 2156 136 2159 139 ne
rect 2159 136 2232 139
tri 2159 109 2186 136 ne
rect 2186 102 2192 136
rect 2226 102 2232 136
rect 2186 90 2232 102
tri 239 81 242 84 se
rect 242 81 248 84
rect 157 75 248 81
rect 300 75 328 84
rect 380 75 408 84
rect 460 75 488 84
rect 540 81 546 84
tri 546 81 549 84 sw
rect 540 75 2159 81
rect 157 41 169 75
rect 203 41 241 75
rect 300 41 313 75
rect 380 41 385 75
rect 563 41 601 75
rect 635 41 673 75
rect 707 41 745 75
rect 779 41 817 75
rect 851 41 889 75
rect 923 41 961 75
rect 995 41 1033 75
rect 1067 41 1105 75
rect 1139 41 1177 75
rect 1211 41 1249 75
rect 1283 41 1321 75
rect 1355 41 1393 75
rect 1427 41 1465 75
rect 1499 41 1537 75
rect 1571 41 1609 75
rect 1643 41 1681 75
rect 1715 41 1753 75
rect 1787 41 1825 75
rect 1859 41 1897 75
rect 1931 41 1969 75
rect 2003 41 2041 75
rect 2075 41 2113 75
rect 2147 41 2159 75
rect 157 35 248 41
tri 239 32 242 35 ne
rect 242 32 248 35
rect 300 32 328 41
rect 380 32 408 41
rect 460 32 488 41
rect 540 35 2159 41
rect 540 32 546 35
tri 546 32 549 35 nw
tri -1959 -625 -1893 -559 se
tri -1893 -625 -1827 -559 nw
tri -1693 -622 -1630 -559 se
rect -1630 -576 -1581 -559
rect -1630 -622 -1627 -576
tri -1627 -622 -1581 -576 nw
tri -1696 -625 -1693 -622 se
tri -2025 -691 -1959 -625 se
tri -1959 -691 -1893 -625 nw
tri -1759 -688 -1696 -625 se
rect -1696 -688 -1693 -625
tri -1693 -688 -1627 -622 nw
tri -1762 -691 -1759 -688 se
tri -2091 -757 -2025 -691 se
tri -2025 -757 -1959 -691 nw
tri -1825 -754 -1762 -691 se
rect -1762 -754 -1759 -691
tri -1759 -754 -1693 -688 nw
tri -1828 -757 -1825 -754 se
tri -2157 -823 -2091 -757 se
tri -2091 -823 -2025 -757 nw
tri -1891 -820 -1828 -757 se
rect -1828 -820 -1825 -757
tri -1825 -820 -1759 -754 nw
tri -1894 -823 -1891 -820 se
tri -2223 -889 -2157 -823 se
tri -2157 -889 -2091 -823 nw
tri -1957 -886 -1894 -823 se
rect -1894 -886 -1891 -823
tri -1891 -886 -1825 -820 nw
tri -1960 -889 -1957 -886 se
tri -2289 -955 -2223 -889 se
tri -2223 -955 -2157 -889 nw
tri -2023 -952 -1960 -889 se
rect -1960 -952 -1957 -889
tri -1957 -952 -1891 -886 nw
tri -2026 -955 -2023 -952 se
tri -2329 -995 -2289 -955 se
tri -9796 -1054 -9757 -1015 ne
rect -9757 -1021 -9750 -1015
tri -9750 -1021 -9724 -995 sw
tri -2355 -1021 -2329 -995 se
rect -2329 -1021 -2289 -995
tri -2289 -1021 -2223 -955 nw
tri -2089 -1018 -2026 -955 se
rect -2026 -1018 -2023 -955
tri -2023 -1018 -1957 -952 nw
tri -2092 -1021 -2089 -1018 se
rect -9757 -1054 -9724 -1021
tri -9724 -1054 -9691 -1021 sw
tri -2388 -1054 -2355 -1021 se
rect -28202 -1094 -28189 -1060
rect -28155 -1094 -28115 -1060
rect -28081 -1094 -28041 -1060
rect -28007 -1094 -27967 -1060
rect -27933 -1094 -27893 -1060
rect -27859 -1094 -27819 -1060
rect -27785 -1094 -27745 -1060
rect -27711 -1094 -27671 -1060
rect -27637 -1094 -27597 -1060
rect -27563 -1094 -27523 -1060
rect -27489 -1094 -27449 -1060
rect -27415 -1094 -27375 -1060
rect -27341 -1094 -27301 -1060
rect -27267 -1094 -27227 -1060
rect -27193 -1094 -27153 -1060
rect -27119 -1094 -27106 -1060
tri -9757 -1061 -9750 -1054 ne
rect -9750 -1061 -9691 -1054
rect -28202 -1132 -27106 -1094
tri -9750 -1120 -9691 -1061 ne
tri -9691 -1087 -9658 -1054 sw
tri -2421 -1087 -2388 -1054 se
rect -2388 -1087 -2355 -1054
tri -2355 -1087 -2289 -1021 nw
tri -2155 -1084 -2092 -1021 se
rect -2092 -1084 -2089 -1021
tri -2089 -1084 -2023 -1018 nw
tri -2158 -1087 -2155 -1084 se
rect -9691 -1120 -9658 -1087
tri -9658 -1120 -9625 -1087 sw
tri -2454 -1120 -2421 -1087 se
rect -28202 -1166 -28189 -1132
rect -28155 -1166 -28115 -1132
rect -28081 -1166 -28041 -1132
rect -28007 -1166 -27967 -1132
rect -27933 -1166 -27893 -1132
rect -27859 -1166 -27819 -1132
rect -27785 -1166 -27745 -1132
rect -27711 -1166 -27671 -1132
rect -27637 -1166 -27597 -1132
rect -27563 -1166 -27523 -1132
rect -27489 -1166 -27449 -1132
rect -27415 -1166 -27375 -1132
rect -27341 -1166 -27301 -1132
rect -27267 -1166 -27227 -1132
rect -27193 -1166 -27153 -1132
rect -27119 -1166 -27106 -1132
rect -28202 -1204 -27106 -1166
tri -9691 -1186 -9625 -1120 ne
tri -9625 -1153 -9592 -1120 sw
tri -2487 -1153 -2454 -1120 se
rect -2454 -1153 -2421 -1120
tri -2421 -1153 -2355 -1087 nw
tri -2221 -1150 -2158 -1087 se
rect -2158 -1150 -2155 -1087
tri -2155 -1150 -2089 -1084 nw
tri -2224 -1153 -2221 -1150 se
rect -9625 -1186 -9592 -1153
tri -9592 -1186 -9559 -1153 sw
tri -2520 -1186 -2487 -1153 se
rect -2487 -1186 -2454 -1153
tri -2454 -1186 -2421 -1153 nw
tri -2257 -1186 -2224 -1153 se
rect -2224 -1186 -2221 -1153
rect -28202 -1238 -28189 -1204
rect -28155 -1238 -28115 -1204
rect -28081 -1238 -28041 -1204
rect -28007 -1238 -27967 -1204
rect -27933 -1238 -27893 -1204
rect -27859 -1238 -27819 -1204
rect -27785 -1238 -27745 -1204
rect -27711 -1238 -27671 -1204
rect -27637 -1238 -27597 -1204
rect -27563 -1238 -27523 -1204
rect -27489 -1238 -27449 -1204
rect -27415 -1238 -27375 -1204
rect -27341 -1238 -27301 -1204
rect -27267 -1238 -27227 -1204
rect -27193 -1238 -27153 -1204
rect -27119 -1238 -27106 -1204
tri -9625 -1232 -9579 -1186 ne
rect -9579 -1232 -2500 -1186
tri -2500 -1232 -2454 -1186 nw
tri -2287 -1216 -2257 -1186 se
rect -2257 -1216 -2221 -1186
tri -2221 -1216 -2155 -1150 nw
tri -2303 -1232 -2287 -1216 se
rect -28202 -1276 -27106 -1238
rect -28202 -1310 -28189 -1276
rect -28155 -1310 -28115 -1276
rect -28081 -1310 -28041 -1276
rect -28007 -1310 -27967 -1276
rect -27933 -1310 -27893 -1276
rect -27859 -1310 -27819 -1276
rect -27785 -1310 -27745 -1276
rect -27711 -1310 -27671 -1276
rect -27637 -1310 -27597 -1276
rect -27563 -1310 -27523 -1276
rect -27489 -1310 -27449 -1276
rect -27415 -1310 -27375 -1276
rect -27341 -1310 -27301 -1276
rect -27267 -1310 -27227 -1276
rect -27193 -1310 -27153 -1276
rect -27119 -1310 -27106 -1276
tri -2353 -1282 -2303 -1232 se
rect -2303 -1282 -2287 -1232
tri -2287 -1282 -2221 -1216 nw
tri -2371 -1300 -2353 -1282 se
rect -2353 -1300 -2305 -1282
tri -2305 -1300 -2287 -1282 nw
rect -28202 -1348 -27106 -1310
rect -28202 -1382 -28189 -1348
rect -28155 -1382 -28115 -1348
rect -28081 -1382 -28041 -1348
rect -28007 -1382 -27967 -1348
rect -27933 -1382 -27893 -1348
rect -27859 -1382 -27819 -1348
rect -27785 -1382 -27745 -1348
rect -27711 -1382 -27671 -1348
rect -27637 -1382 -27597 -1348
rect -27563 -1382 -27523 -1348
rect -27489 -1382 -27449 -1348
rect -27415 -1382 -27375 -1348
rect -27341 -1382 -27301 -1348
rect -27267 -1382 -27227 -1348
rect -27193 -1382 -27153 -1348
rect -27119 -1382 -27106 -1348
tri -10781 -1366 -10715 -1300 se
rect -10715 -1346 -2351 -1300
tri -2351 -1346 -2305 -1300 nw
tri -10715 -1366 -10695 -1346 nw
rect -28202 -1420 -27106 -1382
rect -28202 -1454 -28189 -1420
rect -28155 -1454 -28115 -1420
rect -28081 -1454 -28041 -1420
rect -28007 -1454 -27967 -1420
rect -27933 -1454 -27893 -1420
rect -27859 -1454 -27819 -1420
rect -27785 -1454 -27745 -1420
rect -27711 -1454 -27671 -1420
rect -27637 -1454 -27597 -1420
rect -27563 -1454 -27523 -1420
rect -27489 -1454 -27449 -1420
rect -27415 -1454 -27375 -1420
rect -27341 -1454 -27301 -1420
rect -27267 -1454 -27227 -1420
rect -27193 -1454 -27153 -1420
rect -27119 -1454 -27106 -1420
tri -10847 -1432 -10781 -1366 se
tri -10781 -1432 -10715 -1366 nw
rect -28202 -1492 -27106 -1454
rect -28202 -1526 -28189 -1492
rect -28155 -1526 -28115 -1492
rect -28081 -1526 -28041 -1492
rect -28007 -1526 -27967 -1492
rect -27933 -1526 -27893 -1492
rect -27859 -1526 -27819 -1492
rect -27785 -1526 -27745 -1492
rect -27711 -1526 -27671 -1492
rect -27637 -1526 -27597 -1492
rect -27563 -1526 -27523 -1492
rect -27489 -1526 -27449 -1492
rect -27415 -1526 -27375 -1492
rect -27341 -1526 -27301 -1492
rect -27267 -1526 -27227 -1492
rect -27193 -1526 -27153 -1492
rect -27119 -1526 -27106 -1492
tri -10913 -1498 -10847 -1432 se
tri -10847 -1498 -10781 -1432 nw
rect -28202 -1564 -27106 -1526
tri -10979 -1564 -10913 -1498 se
tri -10913 -1564 -10847 -1498 nw
rect -28202 -1598 -28189 -1564
rect -28155 -1598 -28115 -1564
rect -28081 -1598 -28041 -1564
rect -28007 -1598 -27967 -1564
rect -27933 -1598 -27893 -1564
rect -27859 -1598 -27819 -1564
rect -27785 -1598 -27745 -1564
rect -27711 -1598 -27671 -1564
rect -27637 -1598 -27597 -1564
rect -27563 -1598 -27523 -1564
rect -27489 -1598 -27449 -1564
rect -27415 -1598 -27375 -1564
rect -27341 -1598 -27301 -1564
rect -27267 -1598 -27227 -1564
rect -27193 -1598 -27153 -1564
rect -27119 -1598 -27106 -1564
rect -28202 -1636 -27106 -1598
tri -11045 -1630 -10979 -1564 se
tri -10979 -1630 -10913 -1564 nw
rect -28202 -1670 -28189 -1636
rect -28155 -1670 -28115 -1636
rect -28081 -1670 -28041 -1636
rect -28007 -1670 -27967 -1636
rect -27933 -1670 -27893 -1636
rect -27859 -1670 -27819 -1636
rect -27785 -1670 -27745 -1636
rect -27711 -1670 -27671 -1636
rect -27637 -1670 -27597 -1636
rect -27563 -1670 -27523 -1636
rect -27489 -1670 -27449 -1636
rect -27415 -1670 -27375 -1636
rect -27341 -1670 -27301 -1636
rect -27267 -1670 -27227 -1636
rect -27193 -1670 -27153 -1636
rect -27119 -1670 -27106 -1636
rect -28202 -1708 -27106 -1670
tri -11111 -1696 -11045 -1630 se
tri -11045 -1696 -10979 -1630 nw
rect -28202 -1742 -28189 -1708
rect -28155 -1742 -28115 -1708
rect -28081 -1742 -28041 -1708
rect -28007 -1742 -27967 -1708
rect -27933 -1742 -27893 -1708
rect -27859 -1742 -27819 -1708
rect -27785 -1742 -27745 -1708
rect -27711 -1742 -27671 -1708
rect -27637 -1742 -27597 -1708
rect -27563 -1742 -27523 -1708
rect -27489 -1742 -27449 -1708
rect -27415 -1742 -27375 -1708
rect -27341 -1742 -27301 -1708
rect -27267 -1742 -27227 -1708
rect -27193 -1742 -27153 -1708
rect -27119 -1742 -27106 -1708
rect -28202 -1780 -27106 -1742
tri -11177 -1762 -11111 -1696 se
tri -11111 -1762 -11045 -1696 nw
rect -28202 -1814 -28189 -1780
rect -28155 -1814 -28115 -1780
rect -28081 -1814 -28041 -1780
rect -28007 -1814 -27967 -1780
rect -27933 -1814 -27893 -1780
rect -27859 -1814 -27819 -1780
rect -27785 -1814 -27745 -1780
rect -27711 -1814 -27671 -1780
rect -27637 -1814 -27597 -1780
rect -27563 -1814 -27523 -1780
rect -27489 -1814 -27449 -1780
rect -27415 -1814 -27375 -1780
rect -27341 -1814 -27301 -1780
rect -27267 -1814 -27227 -1780
rect -27193 -1814 -27153 -1780
rect -27119 -1814 -27106 -1780
rect -28202 -1852 -27106 -1814
tri -11243 -1828 -11177 -1762 se
tri -11177 -1828 -11111 -1762 nw
rect -28202 -1886 -28189 -1852
rect -28155 -1886 -28115 -1852
rect -28081 -1886 -28041 -1852
rect -28007 -1886 -27967 -1852
rect -27933 -1886 -27893 -1852
rect -27859 -1886 -27819 -1852
rect -27785 -1886 -27745 -1852
rect -27711 -1886 -27671 -1852
rect -27637 -1886 -27597 -1852
rect -27563 -1886 -27523 -1852
rect -27489 -1886 -27449 -1852
rect -27415 -1886 -27375 -1852
rect -27341 -1886 -27301 -1852
rect -27267 -1886 -27227 -1852
rect -27193 -1886 -27153 -1852
rect -27119 -1886 -27106 -1852
rect -28202 -1924 -27106 -1886
tri -11309 -1894 -11243 -1828 se
tri -11243 -1894 -11177 -1828 nw
rect -28202 -1958 -28189 -1924
rect -28155 -1958 -28115 -1924
rect -28081 -1958 -28041 -1924
rect -28007 -1958 -27967 -1924
rect -27933 -1958 -27893 -1924
rect -27859 -1958 -27819 -1924
rect -27785 -1958 -27745 -1924
rect -27711 -1958 -27671 -1924
rect -27637 -1958 -27597 -1924
rect -27563 -1958 -27523 -1924
rect -27489 -1958 -27449 -1924
rect -27415 -1958 -27375 -1924
rect -27341 -1958 -27301 -1924
rect -27267 -1958 -27227 -1924
rect -27193 -1958 -27153 -1924
rect -27119 -1958 -27106 -1924
rect -28202 -1996 -27106 -1958
tri -11375 -1960 -11309 -1894 se
tri -11309 -1960 -11243 -1894 nw
rect -28202 -2030 -28189 -1996
rect -28155 -2030 -28115 -1996
rect -28081 -2030 -28041 -1996
rect -28007 -2030 -27967 -1996
rect -27933 -2030 -27893 -1996
rect -27859 -2030 -27819 -1996
rect -27785 -2030 -27745 -1996
rect -27711 -2030 -27671 -1996
rect -27637 -2030 -27597 -1996
rect -27563 -2030 -27523 -1996
rect -27489 -2030 -27449 -1996
rect -27415 -2030 -27375 -1996
rect -27341 -2030 -27301 -1996
rect -27267 -2030 -27227 -1996
rect -27193 -2030 -27153 -1996
rect -27119 -2030 -27106 -1996
tri -11441 -2026 -11375 -1960 se
tri -11375 -2026 -11309 -1960 nw
rect -28202 -2068 -27106 -2030
rect -28202 -2102 -28189 -2068
rect -28155 -2102 -28115 -2068
rect -28081 -2102 -28041 -2068
rect -28007 -2102 -27967 -2068
rect -27933 -2102 -27893 -2068
rect -27859 -2102 -27819 -2068
rect -27785 -2102 -27745 -2068
rect -27711 -2102 -27671 -2068
rect -27637 -2102 -27597 -2068
rect -27563 -2102 -27523 -2068
rect -27489 -2102 -27449 -2068
rect -27415 -2102 -27375 -2068
rect -27341 -2102 -27301 -2068
rect -27267 -2102 -27227 -2068
rect -27193 -2102 -27153 -2068
rect -27119 -2102 -27106 -2068
tri -11507 -2092 -11441 -2026 se
tri -11441 -2092 -11375 -2026 nw
rect -28202 -2140 -27106 -2102
rect -28202 -2174 -28189 -2140
rect -28155 -2174 -28115 -2140
rect -28081 -2174 -28041 -2140
rect -28007 -2174 -27967 -2140
rect -27933 -2174 -27893 -2140
rect -27859 -2174 -27819 -2140
rect -27785 -2174 -27745 -2140
rect -27711 -2174 -27671 -2140
rect -27637 -2174 -27597 -2140
rect -27563 -2174 -27523 -2140
rect -27489 -2174 -27449 -2140
rect -27415 -2174 -27375 -2140
rect -27341 -2174 -27301 -2140
rect -27267 -2174 -27227 -2140
rect -27193 -2174 -27153 -2140
rect -27119 -2174 -27106 -2140
rect -28202 -2212 -27106 -2174
rect -28202 -2246 -28189 -2212
rect -28155 -2246 -28115 -2212
rect -28081 -2246 -28041 -2212
rect -28007 -2246 -27967 -2212
rect -27933 -2246 -27893 -2212
rect -27859 -2246 -27819 -2212
rect -27785 -2246 -27745 -2212
rect -27711 -2246 -27671 -2212
rect -27637 -2246 -27597 -2212
rect -27563 -2246 -27523 -2212
rect -27489 -2246 -27449 -2212
rect -27415 -2246 -27375 -2212
rect -27341 -2246 -27301 -2212
rect -27267 -2246 -27227 -2212
rect -27193 -2246 -27153 -2212
rect -27119 -2246 -27106 -2212
rect -28202 -2284 -27106 -2246
rect -28202 -2318 -28189 -2284
rect -28155 -2318 -28115 -2284
rect -28081 -2318 -28041 -2284
rect -28007 -2318 -27967 -2284
rect -27933 -2318 -27893 -2284
rect -27859 -2318 -27819 -2284
rect -27785 -2318 -27745 -2284
rect -27711 -2318 -27671 -2284
rect -27637 -2318 -27597 -2284
rect -27563 -2318 -27523 -2284
rect -27489 -2318 -27449 -2284
rect -27415 -2318 -27375 -2284
rect -27341 -2318 -27301 -2284
rect -27267 -2318 -27227 -2284
rect -27193 -2318 -27153 -2284
rect -27119 -2318 -27106 -2284
rect -28202 -2356 -27106 -2318
rect -28202 -2390 -28189 -2356
rect -28155 -2390 -28115 -2356
rect -28081 -2390 -28041 -2356
rect -28007 -2390 -27967 -2356
rect -27933 -2390 -27893 -2356
rect -27859 -2390 -27819 -2356
rect -27785 -2390 -27745 -2356
rect -27711 -2390 -27671 -2356
rect -27637 -2390 -27597 -2356
rect -27563 -2390 -27523 -2356
rect -27489 -2390 -27449 -2356
rect -27415 -2390 -27375 -2356
rect -27341 -2390 -27301 -2356
rect -27267 -2390 -27227 -2356
rect -27193 -2390 -27153 -2356
rect -27119 -2390 -27106 -2356
rect -28202 -2428 -27106 -2390
rect -28202 -2462 -28189 -2428
rect -28155 -2462 -28115 -2428
rect -28081 -2462 -28041 -2428
rect -28007 -2462 -27967 -2428
rect -27933 -2462 -27893 -2428
rect -27859 -2462 -27819 -2428
rect -27785 -2462 -27745 -2428
rect -27711 -2462 -27671 -2428
rect -27637 -2462 -27597 -2428
rect -27563 -2462 -27523 -2428
rect -27489 -2462 -27449 -2428
rect -27415 -2462 -27375 -2428
rect -27341 -2462 -27301 -2428
rect -27267 -2462 -27227 -2428
rect -27193 -2462 -27153 -2428
rect -27119 -2462 -27106 -2428
rect -28202 -2500 -27106 -2462
rect -28202 -2534 -28189 -2500
rect -28155 -2534 -28115 -2500
rect -28081 -2534 -28041 -2500
rect -28007 -2534 -27967 -2500
rect -27933 -2534 -27893 -2500
rect -27859 -2534 -27819 -2500
rect -27785 -2534 -27745 -2500
rect -27711 -2534 -27671 -2500
rect -27637 -2534 -27597 -2500
rect -27563 -2534 -27523 -2500
rect -27489 -2534 -27449 -2500
rect -27415 -2534 -27375 -2500
rect -27341 -2534 -27301 -2500
rect -27267 -2534 -27227 -2500
rect -27193 -2534 -27153 -2500
rect -27119 -2534 -27106 -2500
rect -28202 -2572 -27106 -2534
rect -28202 -2606 -28189 -2572
rect -28155 -2606 -28115 -2572
rect -28081 -2606 -28041 -2572
rect -28007 -2606 -27967 -2572
rect -27933 -2606 -27893 -2572
rect -27859 -2606 -27819 -2572
rect -27785 -2606 -27745 -2572
rect -27711 -2606 -27671 -2572
rect -27637 -2606 -27597 -2572
rect -27563 -2606 -27523 -2572
rect -27489 -2606 -27449 -2572
rect -27415 -2606 -27375 -2572
rect -27341 -2606 -27301 -2572
rect -27267 -2606 -27227 -2572
rect -27193 -2606 -27153 -2572
rect -27119 -2606 -27106 -2572
rect -28202 -2644 -27106 -2606
rect -28202 -2678 -28189 -2644
rect -28155 -2678 -28115 -2644
rect -28081 -2678 -28041 -2644
rect -28007 -2678 -27967 -2644
rect -27933 -2678 -27893 -2644
rect -27859 -2678 -27819 -2644
rect -27785 -2678 -27745 -2644
rect -27711 -2678 -27671 -2644
rect -27637 -2678 -27597 -2644
rect -27563 -2678 -27523 -2644
rect -27489 -2678 -27449 -2644
rect -27415 -2678 -27375 -2644
rect -27341 -2678 -27301 -2644
rect -27267 -2678 -27227 -2644
rect -27193 -2678 -27153 -2644
rect -27119 -2678 -27106 -2644
rect -28202 -2716 -27106 -2678
rect -28202 -2750 -28189 -2716
rect -28155 -2750 -28115 -2716
rect -28081 -2750 -28041 -2716
rect -28007 -2750 -27967 -2716
rect -27933 -2750 -27893 -2716
rect -27859 -2750 -27819 -2716
rect -27785 -2750 -27745 -2716
rect -27711 -2750 -27671 -2716
rect -27637 -2750 -27597 -2716
rect -27563 -2750 -27523 -2716
rect -27489 -2750 -27449 -2716
rect -27415 -2750 -27375 -2716
rect -27341 -2750 -27301 -2716
rect -27267 -2750 -27227 -2716
rect -27193 -2750 -27153 -2716
rect -27119 -2750 -27106 -2716
rect -28202 -2788 -27106 -2750
rect -28202 -2822 -28189 -2788
rect -28155 -2822 -28115 -2788
rect -28081 -2822 -28041 -2788
rect -28007 -2822 -27967 -2788
rect -27933 -2822 -27893 -2788
rect -27859 -2822 -27819 -2788
rect -27785 -2822 -27745 -2788
rect -27711 -2822 -27671 -2788
rect -27637 -2822 -27597 -2788
rect -27563 -2822 -27523 -2788
rect -27489 -2822 -27449 -2788
rect -27415 -2822 -27375 -2788
rect -27341 -2822 -27301 -2788
rect -27267 -2822 -27227 -2788
rect -27193 -2822 -27153 -2788
rect -27119 -2822 -27106 -2788
rect -28202 -2860 -27106 -2822
rect -28202 -2894 -28189 -2860
rect -28155 -2894 -28115 -2860
rect -28081 -2894 -28041 -2860
rect -28007 -2894 -27967 -2860
rect -27933 -2894 -27893 -2860
rect -27859 -2894 -27819 -2860
rect -27785 -2894 -27745 -2860
rect -27711 -2894 -27671 -2860
rect -27637 -2894 -27597 -2860
rect -27563 -2894 -27523 -2860
rect -27489 -2894 -27449 -2860
rect -27415 -2894 -27375 -2860
rect -27341 -2894 -27301 -2860
rect -27267 -2894 -27227 -2860
rect -27193 -2894 -27153 -2860
rect -27119 -2894 -27106 -2860
rect -28202 -2932 -27106 -2894
rect -28202 -2966 -28189 -2932
rect -28155 -2966 -28115 -2932
rect -28081 -2966 -28041 -2932
rect -28007 -2966 -27967 -2932
rect -27933 -2966 -27893 -2932
rect -27859 -2966 -27819 -2932
rect -27785 -2966 -27745 -2932
rect -27711 -2966 -27671 -2932
rect -27637 -2966 -27597 -2932
rect -27563 -2966 -27523 -2932
rect -27489 -2966 -27449 -2932
rect -27415 -2966 -27375 -2932
rect -27341 -2966 -27301 -2932
rect -27267 -2966 -27227 -2932
rect -27193 -2966 -27153 -2932
rect -27119 -2966 -27106 -2932
rect -28202 -3004 -27106 -2966
rect -28202 -3038 -28189 -3004
rect -28155 -3038 -28115 -3004
rect -28081 -3038 -28041 -3004
rect -28007 -3038 -27967 -3004
rect -27933 -3038 -27893 -3004
rect -27859 -3038 -27819 -3004
rect -27785 -3038 -27745 -3004
rect -27711 -3038 -27671 -3004
rect -27637 -3038 -27597 -3004
rect -27563 -3038 -27523 -3004
rect -27489 -3038 -27449 -3004
rect -27415 -3038 -27375 -3004
rect -27341 -3038 -27301 -3004
rect -27267 -3038 -27227 -3004
rect -27193 -3038 -27153 -3004
rect -27119 -3038 -27106 -3004
rect -28202 -3076 -27106 -3038
rect -28202 -3110 -28189 -3076
rect -28155 -3110 -28115 -3076
rect -28081 -3110 -28041 -3076
rect -28007 -3110 -27967 -3076
rect -27933 -3110 -27893 -3076
rect -27859 -3110 -27819 -3076
rect -27785 -3110 -27745 -3076
rect -27711 -3110 -27671 -3076
rect -27637 -3110 -27597 -3076
rect -27563 -3110 -27523 -3076
rect -27489 -3110 -27449 -3076
rect -27415 -3110 -27375 -3076
rect -27341 -3110 -27301 -3076
rect -27267 -3110 -27227 -3076
rect -27193 -3110 -27153 -3076
rect -27119 -3110 -27106 -3076
rect -28202 -3148 -27106 -3110
rect -28202 -3182 -28189 -3148
rect -28155 -3182 -28115 -3148
rect -28081 -3182 -28041 -3148
rect -28007 -3182 -27967 -3148
rect -27933 -3182 -27893 -3148
rect -27859 -3182 -27819 -3148
rect -27785 -3182 -27745 -3148
rect -27711 -3182 -27671 -3148
rect -27637 -3182 -27597 -3148
rect -27563 -3182 -27523 -3148
rect -27489 -3182 -27449 -3148
rect -27415 -3182 -27375 -3148
rect -27341 -3182 -27301 -3148
rect -27267 -3182 -27227 -3148
rect -27193 -3182 -27153 -3148
rect -27119 -3182 -27106 -3148
rect -28202 -3220 -27106 -3182
rect -28202 -3254 -28189 -3220
rect -28155 -3254 -28115 -3220
rect -28081 -3254 -28041 -3220
rect -28007 -3254 -27967 -3220
rect -27933 -3254 -27893 -3220
rect -27859 -3254 -27819 -3220
rect -27785 -3254 -27745 -3220
rect -27711 -3254 -27671 -3220
rect -27637 -3254 -27597 -3220
rect -27563 -3254 -27523 -3220
rect -27489 -3254 -27449 -3220
rect -27415 -3254 -27375 -3220
rect -27341 -3254 -27301 -3220
rect -27267 -3254 -27227 -3220
rect -27193 -3254 -27153 -3220
rect -27119 -3254 -27106 -3220
rect -28202 -3292 -27106 -3254
rect -28202 -3326 -28189 -3292
rect -28155 -3326 -28115 -3292
rect -28081 -3326 -28041 -3292
rect -28007 -3326 -27967 -3292
rect -27933 -3326 -27893 -3292
rect -27859 -3326 -27819 -3292
rect -27785 -3326 -27745 -3292
rect -27711 -3326 -27671 -3292
rect -27637 -3326 -27597 -3292
rect -27563 -3326 -27523 -3292
rect -27489 -3326 -27449 -3292
rect -27415 -3326 -27375 -3292
rect -27341 -3326 -27301 -3292
rect -27267 -3326 -27227 -3292
rect -27193 -3326 -27153 -3292
rect -27119 -3326 -27106 -3292
rect -28202 -3364 -27106 -3326
rect -28202 -3398 -28189 -3364
rect -28155 -3398 -28115 -3364
rect -28081 -3398 -28041 -3364
rect -28007 -3398 -27967 -3364
rect -27933 -3398 -27893 -3364
rect -27859 -3398 -27819 -3364
rect -27785 -3398 -27745 -3364
rect -27711 -3398 -27671 -3364
rect -27637 -3398 -27597 -3364
rect -27563 -3398 -27523 -3364
rect -27489 -3398 -27449 -3364
rect -27415 -3398 -27375 -3364
rect -27341 -3398 -27301 -3364
rect -27267 -3398 -27227 -3364
rect -27193 -3398 -27153 -3364
rect -27119 -3398 -27106 -3364
rect -28202 -3436 -27106 -3398
rect -28202 -3470 -28189 -3436
rect -28155 -3470 -28115 -3436
rect -28081 -3470 -28041 -3436
rect -28007 -3470 -27967 -3436
rect -27933 -3470 -27893 -3436
rect -27859 -3470 -27819 -3436
rect -27785 -3470 -27745 -3436
rect -27711 -3470 -27671 -3436
rect -27637 -3470 -27597 -3436
rect -27563 -3470 -27523 -3436
rect -27489 -3470 -27449 -3436
rect -27415 -3470 -27375 -3436
rect -27341 -3470 -27301 -3436
rect -27267 -3470 -27227 -3436
rect -27193 -3470 -27153 -3436
rect -27119 -3470 -27106 -3436
rect -28202 -3508 -27106 -3470
rect -28202 -3542 -28189 -3508
rect -28155 -3542 -28115 -3508
rect -28081 -3542 -28041 -3508
rect -28007 -3542 -27967 -3508
rect -27933 -3542 -27893 -3508
rect -27859 -3542 -27819 -3508
rect -27785 -3542 -27745 -3508
rect -27711 -3542 -27671 -3508
rect -27637 -3542 -27597 -3508
rect -27563 -3542 -27523 -3508
rect -27489 -3542 -27449 -3508
rect -27415 -3542 -27375 -3508
rect -27341 -3542 -27301 -3508
rect -27267 -3542 -27227 -3508
rect -27193 -3542 -27153 -3508
rect -27119 -3542 -27106 -3508
rect -28202 -3580 -27106 -3542
rect -28202 -3614 -28189 -3580
rect -28155 -3614 -28115 -3580
rect -28081 -3614 -28041 -3580
rect -28007 -3614 -27967 -3580
rect -27933 -3614 -27893 -3580
rect -27859 -3614 -27819 -3580
rect -27785 -3614 -27745 -3580
rect -27711 -3614 -27671 -3580
rect -27637 -3614 -27597 -3580
rect -27563 -3614 -27523 -3580
rect -27489 -3614 -27449 -3580
rect -27415 -3614 -27375 -3580
rect -27341 -3614 -27301 -3580
rect -27267 -3614 -27227 -3580
rect -27193 -3614 -27153 -3580
rect -27119 -3614 -27106 -3580
rect -28202 -3652 -27106 -3614
rect -28202 -3686 -28189 -3652
rect -28155 -3686 -28115 -3652
rect -28081 -3686 -28041 -3652
rect -28007 -3686 -27967 -3652
rect -27933 -3686 -27893 -3652
rect -27859 -3686 -27819 -3652
rect -27785 -3686 -27745 -3652
rect -27711 -3686 -27671 -3652
rect -27637 -3686 -27597 -3652
rect -27563 -3686 -27523 -3652
rect -27489 -3686 -27449 -3652
rect -27415 -3686 -27375 -3652
rect -27341 -3686 -27301 -3652
rect -27267 -3686 -27227 -3652
rect -27193 -3686 -27153 -3652
rect -27119 -3686 -27106 -3652
rect -28202 -3724 -27106 -3686
rect -28202 -3758 -28189 -3724
rect -28155 -3758 -28115 -3724
rect -28081 -3758 -28041 -3724
rect -28007 -3758 -27967 -3724
rect -27933 -3758 -27893 -3724
rect -27859 -3758 -27819 -3724
rect -27785 -3758 -27745 -3724
rect -27711 -3758 -27671 -3724
rect -27637 -3758 -27597 -3724
rect -27563 -3758 -27523 -3724
rect -27489 -3758 -27449 -3724
rect -27415 -3758 -27375 -3724
rect -27341 -3758 -27301 -3724
rect -27267 -3758 -27227 -3724
rect -27193 -3758 -27153 -3724
rect -27119 -3758 -27106 -3724
rect -28202 -3796 -27106 -3758
rect -28202 -3830 -28189 -3796
rect -28155 -3830 -28115 -3796
rect -28081 -3830 -28041 -3796
rect -28007 -3830 -27967 -3796
rect -27933 -3830 -27893 -3796
rect -27859 -3830 -27819 -3796
rect -27785 -3830 -27745 -3796
rect -27711 -3830 -27671 -3796
rect -27637 -3830 -27597 -3796
rect -27563 -3830 -27523 -3796
rect -27489 -3830 -27449 -3796
rect -27415 -3830 -27375 -3796
rect -27341 -3830 -27301 -3796
rect -27267 -3830 -27227 -3796
rect -27193 -3830 -27153 -3796
rect -27119 -3830 -27106 -3796
rect -28202 -3868 -27106 -3830
rect -28202 -3902 -28189 -3868
rect -28155 -3902 -28115 -3868
rect -28081 -3902 -28041 -3868
rect -28007 -3902 -27967 -3868
rect -27933 -3902 -27893 -3868
rect -27859 -3902 -27819 -3868
rect -27785 -3902 -27745 -3868
rect -27711 -3902 -27671 -3868
rect -27637 -3902 -27597 -3868
rect -27563 -3902 -27523 -3868
rect -27489 -3902 -27449 -3868
rect -27415 -3902 -27375 -3868
rect -27341 -3902 -27301 -3868
rect -27267 -3902 -27227 -3868
rect -27193 -3902 -27153 -3868
rect -27119 -3902 -27106 -3868
rect -28202 -3940 -27106 -3902
rect -28202 -3974 -28189 -3940
rect -28155 -3974 -28115 -3940
rect -28081 -3974 -28041 -3940
rect -28007 -3974 -27967 -3940
rect -27933 -3974 -27893 -3940
rect -27859 -3974 -27819 -3940
rect -27785 -3974 -27745 -3940
rect -27711 -3974 -27671 -3940
rect -27637 -3974 -27597 -3940
rect -27563 -3974 -27523 -3940
rect -27489 -3974 -27449 -3940
rect -27415 -3974 -27375 -3940
rect -27341 -3974 -27301 -3940
rect -27267 -3974 -27227 -3940
rect -27193 -3974 -27153 -3940
rect -27119 -3974 -27106 -3940
rect -28202 -4012 -27106 -3974
rect -28202 -4046 -28189 -4012
rect -28155 -4046 -28115 -4012
rect -28081 -4046 -28041 -4012
rect -28007 -4046 -27967 -4012
rect -27933 -4046 -27893 -4012
rect -27859 -4046 -27819 -4012
rect -27785 -4046 -27745 -4012
rect -27711 -4046 -27671 -4012
rect -27637 -4046 -27597 -4012
rect -27563 -4046 -27523 -4012
rect -27489 -4046 -27449 -4012
rect -27415 -4046 -27375 -4012
rect -27341 -4046 -27301 -4012
rect -27267 -4046 -27227 -4012
rect -27193 -4046 -27153 -4012
rect -27119 -4046 -27106 -4012
rect -28202 -4084 -27106 -4046
rect -28202 -4118 -28189 -4084
rect -28155 -4118 -28115 -4084
rect -28081 -4118 -28041 -4084
rect -28007 -4118 -27967 -4084
rect -27933 -4118 -27893 -4084
rect -27859 -4118 -27819 -4084
rect -27785 -4118 -27745 -4084
rect -27711 -4118 -27671 -4084
rect -27637 -4118 -27597 -4084
rect -27563 -4118 -27523 -4084
rect -27489 -4118 -27449 -4084
rect -27415 -4118 -27375 -4084
rect -27341 -4118 -27301 -4084
rect -27267 -4118 -27227 -4084
rect -27193 -4118 -27153 -4084
rect -27119 -4118 -27106 -4084
rect -28202 -4156 -27106 -4118
rect -28202 -4190 -28189 -4156
rect -28155 -4190 -28115 -4156
rect -28081 -4190 -28041 -4156
rect -28007 -4190 -27967 -4156
rect -27933 -4190 -27893 -4156
rect -27859 -4190 -27819 -4156
rect -27785 -4190 -27745 -4156
rect -27711 -4190 -27671 -4156
rect -27637 -4190 -27597 -4156
rect -27563 -4190 -27523 -4156
rect -27489 -4190 -27449 -4156
rect -27415 -4190 -27375 -4156
rect -27341 -4190 -27301 -4156
rect -27267 -4190 -27227 -4156
rect -27193 -4190 -27153 -4156
rect -27119 -4190 -27106 -4156
rect -28202 -4228 -27106 -4190
rect -28202 -4262 -28189 -4228
rect -28155 -4262 -28115 -4228
rect -28081 -4262 -28041 -4228
rect -28007 -4262 -27967 -4228
rect -27933 -4262 -27893 -4228
rect -27859 -4262 -27819 -4228
rect -27785 -4262 -27745 -4228
rect -27711 -4262 -27671 -4228
rect -27637 -4262 -27597 -4228
rect -27563 -4262 -27523 -4228
rect -27489 -4262 -27449 -4228
rect -27415 -4262 -27375 -4228
rect -27341 -4262 -27301 -4228
rect -27267 -4262 -27227 -4228
rect -27193 -4262 -27153 -4228
rect -27119 -4262 -27106 -4228
rect -28202 -4300 -27106 -4262
rect -28202 -4334 -28189 -4300
rect -28155 -4334 -28115 -4300
rect -28081 -4334 -28041 -4300
rect -28007 -4334 -27967 -4300
rect -27933 -4334 -27893 -4300
rect -27859 -4334 -27819 -4300
rect -27785 -4334 -27745 -4300
rect -27711 -4334 -27671 -4300
rect -27637 -4334 -27597 -4300
rect -27563 -4334 -27523 -4300
rect -27489 -4334 -27449 -4300
rect -27415 -4334 -27375 -4300
rect -27341 -4334 -27301 -4300
rect -27267 -4334 -27227 -4300
rect -27193 -4334 -27153 -4300
rect -27119 -4334 -27106 -4300
rect -28202 -4372 -27106 -4334
rect -28202 -4406 -28189 -4372
rect -28155 -4406 -28115 -4372
rect -28081 -4406 -28041 -4372
rect -28007 -4406 -27967 -4372
rect -27933 -4406 -27893 -4372
rect -27859 -4406 -27819 -4372
rect -27785 -4406 -27745 -4372
rect -27711 -4406 -27671 -4372
rect -27637 -4406 -27597 -4372
rect -27563 -4406 -27523 -4372
rect -27489 -4406 -27449 -4372
rect -27415 -4406 -27375 -4372
rect -27341 -4406 -27301 -4372
rect -27267 -4406 -27227 -4372
rect -27193 -4406 -27153 -4372
rect -27119 -4406 -27106 -4372
rect -28202 -4444 -27106 -4406
rect -28202 -4478 -28189 -4444
rect -28155 -4478 -28115 -4444
rect -28081 -4478 -28041 -4444
rect -28007 -4478 -27967 -4444
rect -27933 -4478 -27893 -4444
rect -27859 -4478 -27819 -4444
rect -27785 -4478 -27745 -4444
rect -27711 -4478 -27671 -4444
rect -27637 -4478 -27597 -4444
rect -27563 -4478 -27523 -4444
rect -27489 -4478 -27449 -4444
rect -27415 -4478 -27375 -4444
rect -27341 -4478 -27301 -4444
rect -27267 -4478 -27227 -4444
rect -27193 -4478 -27153 -4444
rect -27119 -4478 -27106 -4444
rect -28202 -4516 -27106 -4478
rect -28202 -4550 -28189 -4516
rect -28155 -4550 -28115 -4516
rect -28081 -4550 -28041 -4516
rect -28007 -4550 -27967 -4516
rect -27933 -4550 -27893 -4516
rect -27859 -4550 -27819 -4516
rect -27785 -4550 -27745 -4516
rect -27711 -4550 -27671 -4516
rect -27637 -4550 -27597 -4516
rect -27563 -4550 -27523 -4516
rect -27489 -4550 -27449 -4516
rect -27415 -4550 -27375 -4516
rect -27341 -4550 -27301 -4516
rect -27267 -4550 -27227 -4516
rect -27193 -4550 -27153 -4516
rect -27119 -4550 -27106 -4516
rect -28202 -4588 -27106 -4550
rect -28202 -4622 -28189 -4588
rect -28155 -4622 -28115 -4588
rect -28081 -4622 -28041 -4588
rect -28007 -4622 -27967 -4588
rect -27933 -4622 -27893 -4588
rect -27859 -4622 -27819 -4588
rect -27785 -4622 -27745 -4588
rect -27711 -4622 -27671 -4588
rect -27637 -4622 -27597 -4588
rect -27563 -4622 -27523 -4588
rect -27489 -4622 -27449 -4588
rect -27415 -4622 -27375 -4588
rect -27341 -4622 -27301 -4588
rect -27267 -4622 -27227 -4588
rect -27193 -4622 -27153 -4588
rect -27119 -4622 -27106 -4588
rect -28202 -4660 -27106 -4622
rect -28202 -4694 -28189 -4660
rect -28155 -4694 -28115 -4660
rect -28081 -4694 -28041 -4660
rect -28007 -4694 -27967 -4660
rect -27933 -4694 -27893 -4660
rect -27859 -4694 -27819 -4660
rect -27785 -4694 -27745 -4660
rect -27711 -4694 -27671 -4660
rect -27637 -4694 -27597 -4660
rect -27563 -4694 -27523 -4660
rect -27489 -4694 -27449 -4660
rect -27415 -4694 -27375 -4660
rect -27341 -4694 -27301 -4660
rect -27267 -4694 -27227 -4660
rect -27193 -4694 -27153 -4660
rect -27119 -4694 -27106 -4660
rect -28202 -4732 -27106 -4694
rect -28202 -4766 -28189 -4732
rect -28155 -4766 -28115 -4732
rect -28081 -4766 -28041 -4732
rect -28007 -4766 -27967 -4732
rect -27933 -4766 -27893 -4732
rect -27859 -4766 -27819 -4732
rect -27785 -4766 -27745 -4732
rect -27711 -4766 -27671 -4732
rect -27637 -4766 -27597 -4732
rect -27563 -4766 -27523 -4732
rect -27489 -4766 -27449 -4732
rect -27415 -4766 -27375 -4732
rect -27341 -4766 -27301 -4732
rect -27267 -4766 -27227 -4732
rect -27193 -4766 -27153 -4732
rect -27119 -4766 -27106 -4732
rect -28202 -4804 -27106 -4766
rect -28202 -4838 -28189 -4804
rect -28155 -4838 -28115 -4804
rect -28081 -4838 -28041 -4804
rect -28007 -4838 -27967 -4804
rect -27933 -4838 -27893 -4804
rect -27859 -4838 -27819 -4804
rect -27785 -4838 -27745 -4804
rect -27711 -4838 -27671 -4804
rect -27637 -4838 -27597 -4804
rect -27563 -4838 -27523 -4804
rect -27489 -4838 -27449 -4804
rect -27415 -4838 -27375 -4804
rect -27341 -4838 -27301 -4804
rect -27267 -4838 -27227 -4804
rect -27193 -4838 -27153 -4804
rect -27119 -4838 -27106 -4804
rect -28202 -4876 -27106 -4838
rect -28202 -4910 -28189 -4876
rect -28155 -4910 -28115 -4876
rect -28081 -4910 -28041 -4876
rect -28007 -4910 -27967 -4876
rect -27933 -4910 -27893 -4876
rect -27859 -4910 -27819 -4876
rect -27785 -4910 -27745 -4876
rect -27711 -4910 -27671 -4876
rect -27637 -4910 -27597 -4876
rect -27563 -4910 -27523 -4876
rect -27489 -4910 -27449 -4876
rect -27415 -4910 -27375 -4876
rect -27341 -4910 -27301 -4876
rect -27267 -4910 -27227 -4876
rect -27193 -4910 -27153 -4876
rect -27119 -4910 -27106 -4876
rect -28202 -4948 -27106 -4910
rect -28202 -4982 -28189 -4948
rect -28155 -4982 -28115 -4948
rect -28081 -4982 -28041 -4948
rect -28007 -4982 -27967 -4948
rect -27933 -4982 -27893 -4948
rect -27859 -4982 -27819 -4948
rect -27785 -4982 -27745 -4948
rect -27711 -4982 -27671 -4948
rect -27637 -4982 -27597 -4948
rect -27563 -4982 -27523 -4948
rect -27489 -4982 -27449 -4948
rect -27415 -4982 -27375 -4948
rect -27341 -4982 -27301 -4948
rect -27267 -4982 -27227 -4948
rect -27193 -4982 -27153 -4948
rect -27119 -4982 -27106 -4948
rect -28202 -5020 -27106 -4982
rect -28202 -5054 -28189 -5020
rect -28155 -5054 -28115 -5020
rect -28081 -5054 -28041 -5020
rect -28007 -5054 -27967 -5020
rect -27933 -5054 -27893 -5020
rect -27859 -5054 -27819 -5020
rect -27785 -5054 -27745 -5020
rect -27711 -5054 -27671 -5020
rect -27637 -5054 -27597 -5020
rect -27563 -5054 -27523 -5020
rect -27489 -5054 -27449 -5020
rect -27415 -5054 -27375 -5020
rect -27341 -5054 -27301 -5020
rect -27267 -5054 -27227 -5020
rect -27193 -5054 -27153 -5020
rect -27119 -5054 -27106 -5020
rect -28202 -5092 -27106 -5054
rect -28202 -5126 -28189 -5092
rect -28155 -5126 -28115 -5092
rect -28081 -5126 -28041 -5092
rect -28007 -5126 -27967 -5092
rect -27933 -5126 -27893 -5092
rect -27859 -5126 -27819 -5092
rect -27785 -5126 -27745 -5092
rect -27711 -5126 -27671 -5092
rect -27637 -5126 -27597 -5092
rect -27563 -5126 -27523 -5092
rect -27489 -5126 -27449 -5092
rect -27415 -5126 -27375 -5092
rect -27341 -5126 -27301 -5092
rect -27267 -5126 -27227 -5092
rect -27193 -5126 -27153 -5092
rect -27119 -5126 -27106 -5092
rect -28202 -5164 -27106 -5126
rect -28202 -5198 -28189 -5164
rect -28155 -5198 -28115 -5164
rect -28081 -5198 -28041 -5164
rect -28007 -5198 -27967 -5164
rect -27933 -5198 -27893 -5164
rect -27859 -5198 -27819 -5164
rect -27785 -5198 -27745 -5164
rect -27711 -5198 -27671 -5164
rect -27637 -5198 -27597 -5164
rect -27563 -5198 -27523 -5164
rect -27489 -5198 -27449 -5164
rect -27415 -5198 -27375 -5164
rect -27341 -5198 -27301 -5164
rect -27267 -5198 -27227 -5164
rect -27193 -5198 -27153 -5164
rect -27119 -5198 -27106 -5164
rect -28202 -5236 -27106 -5198
rect -28202 -5270 -28189 -5236
rect -28155 -5270 -28115 -5236
rect -28081 -5270 -28041 -5236
rect -28007 -5270 -27967 -5236
rect -27933 -5270 -27893 -5236
rect -27859 -5270 -27819 -5236
rect -27785 -5270 -27745 -5236
rect -27711 -5270 -27671 -5236
rect -27637 -5270 -27597 -5236
rect -27563 -5270 -27523 -5236
rect -27489 -5270 -27449 -5236
rect -27415 -5270 -27375 -5236
rect -27341 -5270 -27301 -5236
rect -27267 -5270 -27227 -5236
rect -27193 -5270 -27153 -5236
rect -27119 -5270 -27106 -5236
rect -28202 -5308 -27106 -5270
rect -28202 -5342 -28189 -5308
rect -28155 -5342 -28115 -5308
rect -28081 -5342 -28041 -5308
rect -28007 -5342 -27967 -5308
rect -27933 -5342 -27893 -5308
rect -27859 -5342 -27819 -5308
rect -27785 -5342 -27745 -5308
rect -27711 -5342 -27671 -5308
rect -27637 -5342 -27597 -5308
rect -27563 -5342 -27523 -5308
rect -27489 -5342 -27449 -5308
rect -27415 -5342 -27375 -5308
rect -27341 -5342 -27301 -5308
rect -27267 -5342 -27227 -5308
rect -27193 -5342 -27153 -5308
rect -27119 -5342 -27106 -5308
rect -28202 -5380 -27106 -5342
rect -28202 -5414 -28189 -5380
rect -28155 -5414 -28115 -5380
rect -28081 -5414 -28041 -5380
rect -28007 -5414 -27967 -5380
rect -27933 -5414 -27893 -5380
rect -27859 -5414 -27819 -5380
rect -27785 -5414 -27745 -5380
rect -27711 -5414 -27671 -5380
rect -27637 -5414 -27597 -5380
rect -27563 -5414 -27523 -5380
rect -27489 -5414 -27449 -5380
rect -27415 -5414 -27375 -5380
rect -27341 -5414 -27301 -5380
rect -27267 -5414 -27227 -5380
rect -27193 -5414 -27153 -5380
rect -27119 -5414 -27106 -5380
rect -28202 -5452 -27106 -5414
rect -28202 -5486 -28189 -5452
rect -28155 -5486 -28115 -5452
rect -28081 -5486 -28041 -5452
rect -28007 -5486 -27967 -5452
rect -27933 -5486 -27893 -5452
rect -27859 -5486 -27819 -5452
rect -27785 -5486 -27745 -5452
rect -27711 -5486 -27671 -5452
rect -27637 -5486 -27597 -5452
rect -27563 -5486 -27523 -5452
rect -27489 -5486 -27449 -5452
rect -27415 -5486 -27375 -5452
rect -27341 -5486 -27301 -5452
rect -27267 -5486 -27227 -5452
rect -27193 -5486 -27153 -5452
rect -27119 -5486 -27106 -5452
rect -28202 -5524 -27106 -5486
rect -28202 -5558 -28189 -5524
rect -28155 -5558 -28115 -5524
rect -28081 -5558 -28041 -5524
rect -28007 -5558 -27967 -5524
rect -27933 -5558 -27893 -5524
rect -27859 -5558 -27819 -5524
rect -27785 -5558 -27745 -5524
rect -27711 -5558 -27671 -5524
rect -27637 -5558 -27597 -5524
rect -27563 -5558 -27523 -5524
rect -27489 -5558 -27449 -5524
rect -27415 -5558 -27375 -5524
rect -27341 -5558 -27301 -5524
rect -27267 -5558 -27227 -5524
rect -27193 -5558 -27153 -5524
rect -27119 -5558 -27106 -5524
rect -28202 -5596 -27106 -5558
rect -28202 -5630 -28189 -5596
rect -28155 -5630 -28115 -5596
rect -28081 -5630 -28041 -5596
rect -28007 -5630 -27967 -5596
rect -27933 -5630 -27893 -5596
rect -27859 -5630 -27819 -5596
rect -27785 -5630 -27745 -5596
rect -27711 -5630 -27671 -5596
rect -27637 -5630 -27597 -5596
rect -27563 -5630 -27523 -5596
rect -27489 -5630 -27449 -5596
rect -27415 -5630 -27375 -5596
rect -27341 -5630 -27301 -5596
rect -27267 -5630 -27227 -5596
rect -27193 -5630 -27153 -5596
rect -27119 -5630 -27106 -5596
rect -28202 -5668 -27106 -5630
rect -28202 -5702 -28189 -5668
rect -28155 -5702 -28115 -5668
rect -28081 -5702 -28041 -5668
rect -28007 -5702 -27967 -5668
rect -27933 -5702 -27893 -5668
rect -27859 -5702 -27819 -5668
rect -27785 -5702 -27745 -5668
rect -27711 -5702 -27671 -5668
rect -27637 -5702 -27597 -5668
rect -27563 -5702 -27523 -5668
rect -27489 -5702 -27449 -5668
rect -27415 -5702 -27375 -5668
rect -27341 -5702 -27301 -5668
rect -27267 -5702 -27227 -5668
rect -27193 -5702 -27153 -5668
rect -27119 -5702 -27106 -5668
rect -28202 -5740 -27106 -5702
rect -28202 -5774 -28189 -5740
rect -28155 -5774 -28115 -5740
rect -28081 -5774 -28041 -5740
rect -28007 -5774 -27967 -5740
rect -27933 -5774 -27893 -5740
rect -27859 -5774 -27819 -5740
rect -27785 -5774 -27745 -5740
rect -27711 -5774 -27671 -5740
rect -27637 -5774 -27597 -5740
rect -27563 -5774 -27523 -5740
rect -27489 -5774 -27449 -5740
rect -27415 -5774 -27375 -5740
rect -27341 -5774 -27301 -5740
rect -27267 -5774 -27227 -5740
rect -27193 -5774 -27153 -5740
rect -27119 -5774 -27106 -5740
rect -28202 -5812 -27106 -5774
rect -28202 -5846 -28189 -5812
rect -28155 -5846 -28115 -5812
rect -28081 -5846 -28041 -5812
rect -28007 -5846 -27967 -5812
rect -27933 -5846 -27893 -5812
rect -27859 -5846 -27819 -5812
rect -27785 -5846 -27745 -5812
rect -27711 -5846 -27671 -5812
rect -27637 -5846 -27597 -5812
rect -27563 -5846 -27523 -5812
rect -27489 -5846 -27449 -5812
rect -27415 -5846 -27375 -5812
rect -27341 -5846 -27301 -5812
rect -27267 -5846 -27227 -5812
rect -27193 -5846 -27153 -5812
rect -27119 -5846 -27106 -5812
rect -28202 -5884 -27106 -5846
rect -28202 -5918 -28189 -5884
rect -28155 -5918 -28115 -5884
rect -28081 -5918 -28041 -5884
rect -28007 -5918 -27967 -5884
rect -27933 -5918 -27893 -5884
rect -27859 -5918 -27819 -5884
rect -27785 -5918 -27745 -5884
rect -27711 -5918 -27671 -5884
rect -27637 -5918 -27597 -5884
rect -27563 -5918 -27523 -5884
rect -27489 -5918 -27449 -5884
rect -27415 -5918 -27375 -5884
rect -27341 -5918 -27301 -5884
rect -27267 -5918 -27227 -5884
rect -27193 -5918 -27153 -5884
rect -27119 -5918 -27106 -5884
rect -28202 -5956 -27106 -5918
rect -28202 -5990 -28189 -5956
rect -28155 -5990 -28115 -5956
rect -28081 -5990 -28041 -5956
rect -28007 -5990 -27967 -5956
rect -27933 -5990 -27893 -5956
rect -27859 -5990 -27819 -5956
rect -27785 -5990 -27745 -5956
rect -27711 -5990 -27671 -5956
rect -27637 -5990 -27597 -5956
rect -27563 -5990 -27523 -5956
rect -27489 -5990 -27449 -5956
rect -27415 -5990 -27375 -5956
rect -27341 -5990 -27301 -5956
rect -27267 -5990 -27227 -5956
rect -27193 -5990 -27153 -5956
rect -27119 -5990 -27106 -5956
rect -28202 -6028 -27106 -5990
rect -28202 -6062 -28189 -6028
rect -28155 -6062 -28115 -6028
rect -28081 -6062 -28041 -6028
rect -28007 -6062 -27967 -6028
rect -27933 -6062 -27893 -6028
rect -27859 -6062 -27819 -6028
rect -27785 -6062 -27745 -6028
rect -27711 -6062 -27671 -6028
rect -27637 -6062 -27597 -6028
rect -27563 -6062 -27523 -6028
rect -27489 -6062 -27449 -6028
rect -27415 -6062 -27375 -6028
rect -27341 -6062 -27301 -6028
rect -27267 -6062 -27227 -6028
rect -27193 -6062 -27153 -6028
rect -27119 -6062 -27106 -6028
rect -28202 -6100 -27106 -6062
rect -28202 -6134 -28189 -6100
rect -28155 -6134 -28115 -6100
rect -28081 -6134 -28041 -6100
rect -28007 -6134 -27967 -6100
rect -27933 -6134 -27893 -6100
rect -27859 -6134 -27819 -6100
rect -27785 -6134 -27745 -6100
rect -27711 -6134 -27671 -6100
rect -27637 -6134 -27597 -6100
rect -27563 -6134 -27523 -6100
rect -27489 -6134 -27449 -6100
rect -27415 -6134 -27375 -6100
rect -27341 -6134 -27301 -6100
rect -27267 -6134 -27227 -6100
rect -27193 -6134 -27153 -6100
rect -27119 -6134 -27106 -6100
rect -28202 -6172 -27106 -6134
rect -28202 -6206 -28189 -6172
rect -28155 -6206 -28115 -6172
rect -28081 -6206 -28041 -6172
rect -28007 -6206 -27967 -6172
rect -27933 -6206 -27893 -6172
rect -27859 -6206 -27819 -6172
rect -27785 -6206 -27745 -6172
rect -27711 -6206 -27671 -6172
rect -27637 -6206 -27597 -6172
rect -27563 -6206 -27523 -6172
rect -27489 -6206 -27449 -6172
rect -27415 -6206 -27375 -6172
rect -27341 -6206 -27301 -6172
rect -27267 -6206 -27227 -6172
rect -27193 -6206 -27153 -6172
rect -27119 -6206 -27106 -6172
rect -28202 -6244 -27106 -6206
rect -28202 -6278 -28189 -6244
rect -28155 -6278 -28115 -6244
rect -28081 -6278 -28041 -6244
rect -28007 -6278 -27967 -6244
rect -27933 -6278 -27893 -6244
rect -27859 -6278 -27819 -6244
rect -27785 -6278 -27745 -6244
rect -27711 -6278 -27671 -6244
rect -27637 -6278 -27597 -6244
rect -27563 -6278 -27523 -6244
rect -27489 -6278 -27449 -6244
rect -27415 -6278 -27375 -6244
rect -27341 -6278 -27301 -6244
rect -27267 -6278 -27227 -6244
rect -27193 -6278 -27153 -6244
rect -27119 -6278 -27106 -6244
rect -28202 -6316 -27106 -6278
rect -28202 -6350 -28189 -6316
rect -28155 -6350 -28115 -6316
rect -28081 -6350 -28041 -6316
rect -28007 -6350 -27967 -6316
rect -27933 -6350 -27893 -6316
rect -27859 -6350 -27819 -6316
rect -27785 -6350 -27745 -6316
rect -27711 -6350 -27671 -6316
rect -27637 -6350 -27597 -6316
rect -27563 -6350 -27523 -6316
rect -27489 -6350 -27449 -6316
rect -27415 -6350 -27375 -6316
rect -27341 -6350 -27301 -6316
rect -27267 -6350 -27227 -6316
rect -27193 -6350 -27153 -6316
rect -27119 -6350 -27106 -6316
rect -28202 -6388 -27106 -6350
rect -28202 -6422 -28189 -6388
rect -28155 -6422 -28115 -6388
rect -28081 -6422 -28041 -6388
rect -28007 -6422 -27967 -6388
rect -27933 -6422 -27893 -6388
rect -27859 -6422 -27819 -6388
rect -27785 -6422 -27745 -6388
rect -27711 -6422 -27671 -6388
rect -27637 -6422 -27597 -6388
rect -27563 -6422 -27523 -6388
rect -27489 -6422 -27449 -6388
rect -27415 -6422 -27375 -6388
rect -27341 -6422 -27301 -6388
rect -27267 -6422 -27227 -6388
rect -27193 -6422 -27153 -6388
rect -27119 -6422 -27106 -6388
rect -28202 -6460 -27106 -6422
rect -28202 -6494 -28189 -6460
rect -28155 -6494 -28115 -6460
rect -28081 -6494 -28041 -6460
rect -28007 -6494 -27967 -6460
rect -27933 -6494 -27893 -6460
rect -27859 -6494 -27819 -6460
rect -27785 -6494 -27745 -6460
rect -27711 -6494 -27671 -6460
rect -27637 -6494 -27597 -6460
rect -27563 -6494 -27523 -6460
rect -27489 -6494 -27449 -6460
rect -27415 -6494 -27375 -6460
rect -27341 -6494 -27301 -6460
rect -27267 -6494 -27227 -6460
rect -27193 -6494 -27153 -6460
rect -27119 -6494 -27106 -6460
rect -28202 -6532 -27106 -6494
rect -28202 -6566 -28189 -6532
rect -28155 -6566 -28115 -6532
rect -28081 -6566 -28041 -6532
rect -28007 -6566 -27967 -6532
rect -27933 -6566 -27893 -6532
rect -27859 -6566 -27819 -6532
rect -27785 -6566 -27745 -6532
rect -27711 -6566 -27671 -6532
rect -27637 -6566 -27597 -6532
rect -27563 -6566 -27523 -6532
rect -27489 -6566 -27449 -6532
rect -27415 -6566 -27375 -6532
rect -27341 -6566 -27301 -6532
rect -27267 -6566 -27227 -6532
rect -27193 -6566 -27153 -6532
rect -27119 -6566 -27106 -6532
rect -28202 -6604 -27106 -6566
rect -28202 -6638 -28189 -6604
rect -28155 -6638 -28115 -6604
rect -28081 -6638 -28041 -6604
rect -28007 -6638 -27967 -6604
rect -27933 -6638 -27893 -6604
rect -27859 -6638 -27819 -6604
rect -27785 -6638 -27745 -6604
rect -27711 -6638 -27671 -6604
rect -27637 -6638 -27597 -6604
rect -27563 -6638 -27523 -6604
rect -27489 -6638 -27449 -6604
rect -27415 -6638 -27375 -6604
rect -27341 -6638 -27301 -6604
rect -27267 -6638 -27227 -6604
rect -27193 -6638 -27153 -6604
rect -27119 -6638 -27106 -6604
rect -28202 -6676 -27106 -6638
rect -28202 -6710 -28189 -6676
rect -28155 -6710 -28115 -6676
rect -28081 -6710 -28041 -6676
rect -28007 -6710 -27967 -6676
rect -27933 -6710 -27893 -6676
rect -27859 -6710 -27819 -6676
rect -27785 -6710 -27745 -6676
rect -27711 -6710 -27671 -6676
rect -27637 -6710 -27597 -6676
rect -27563 -6710 -27523 -6676
rect -27489 -6710 -27449 -6676
rect -27415 -6710 -27375 -6676
rect -27341 -6710 -27301 -6676
rect -27267 -6710 -27227 -6676
rect -27193 -6710 -27153 -6676
rect -27119 -6710 -27106 -6676
rect -28202 -6748 -27106 -6710
rect -28202 -6782 -28189 -6748
rect -28155 -6782 -28115 -6748
rect -28081 -6782 -28041 -6748
rect -28007 -6782 -27967 -6748
rect -27933 -6782 -27893 -6748
rect -27859 -6782 -27819 -6748
rect -27785 -6782 -27745 -6748
rect -27711 -6782 -27671 -6748
rect -27637 -6782 -27597 -6748
rect -27563 -6782 -27523 -6748
rect -27489 -6782 -27449 -6748
rect -27415 -6782 -27375 -6748
rect -27341 -6782 -27301 -6748
rect -27267 -6782 -27227 -6748
rect -27193 -6782 -27153 -6748
rect -27119 -6782 -27106 -6748
rect -28202 -6820 -27106 -6782
rect -28202 -6854 -28189 -6820
rect -28155 -6854 -28115 -6820
rect -28081 -6854 -28041 -6820
rect -28007 -6854 -27967 -6820
rect -27933 -6854 -27893 -6820
rect -27859 -6854 -27819 -6820
rect -27785 -6854 -27745 -6820
rect -27711 -6854 -27671 -6820
rect -27637 -6854 -27597 -6820
rect -27563 -6854 -27523 -6820
rect -27489 -6854 -27449 -6820
rect -27415 -6854 -27375 -6820
rect -27341 -6854 -27301 -6820
rect -27267 -6854 -27227 -6820
rect -27193 -6854 -27153 -6820
rect -27119 -6854 -27106 -6820
rect -28202 -6892 -27106 -6854
rect -28202 -6926 -28189 -6892
rect -28155 -6926 -28115 -6892
rect -28081 -6926 -28041 -6892
rect -28007 -6926 -27967 -6892
rect -27933 -6926 -27893 -6892
rect -27859 -6926 -27819 -6892
rect -27785 -6926 -27745 -6892
rect -27711 -6926 -27671 -6892
rect -27637 -6926 -27597 -6892
rect -27563 -6926 -27523 -6892
rect -27489 -6926 -27449 -6892
rect -27415 -6926 -27375 -6892
rect -27341 -6926 -27301 -6892
rect -27267 -6926 -27227 -6892
rect -27193 -6926 -27153 -6892
rect -27119 -6926 -27106 -6892
rect -28202 -6964 -27106 -6926
rect -28202 -6998 -28189 -6964
rect -28155 -6998 -28115 -6964
rect -28081 -6998 -28041 -6964
rect -28007 -6998 -27967 -6964
rect -27933 -6998 -27893 -6964
rect -27859 -6998 -27819 -6964
rect -27785 -6998 -27745 -6964
rect -27711 -6998 -27671 -6964
rect -27637 -6998 -27597 -6964
rect -27563 -6998 -27523 -6964
rect -27489 -6998 -27449 -6964
rect -27415 -6998 -27375 -6964
rect -27341 -6998 -27301 -6964
rect -27267 -6998 -27227 -6964
rect -27193 -6998 -27153 -6964
rect -27119 -6998 -27106 -6964
rect -28202 -7036 -27106 -6998
rect -28202 -7070 -28189 -7036
rect -28155 -7070 -28115 -7036
rect -28081 -7070 -28041 -7036
rect -28007 -7070 -27967 -7036
rect -27933 -7070 -27893 -7036
rect -27859 -7070 -27819 -7036
rect -27785 -7070 -27745 -7036
rect -27711 -7070 -27671 -7036
rect -27637 -7070 -27597 -7036
rect -27563 -7070 -27523 -7036
rect -27489 -7070 -27449 -7036
rect -27415 -7070 -27375 -7036
rect -27341 -7070 -27301 -7036
rect -27267 -7070 -27227 -7036
rect -27193 -7070 -27153 -7036
rect -27119 -7070 -27106 -7036
rect -28202 -7108 -27106 -7070
rect -28202 -7142 -28189 -7108
rect -28155 -7142 -28115 -7108
rect -28081 -7142 -28041 -7108
rect -28007 -7142 -27967 -7108
rect -27933 -7142 -27893 -7108
rect -27859 -7142 -27819 -7108
rect -27785 -7142 -27745 -7108
rect -27711 -7142 -27671 -7108
rect -27637 -7142 -27597 -7108
rect -27563 -7142 -27523 -7108
rect -27489 -7142 -27449 -7108
rect -27415 -7142 -27375 -7108
rect -27341 -7142 -27301 -7108
rect -27267 -7142 -27227 -7108
rect -27193 -7142 -27153 -7108
rect -27119 -7142 -27106 -7108
rect -28202 -7180 -27106 -7142
rect -28202 -7214 -28189 -7180
rect -28155 -7214 -28115 -7180
rect -28081 -7214 -28041 -7180
rect -28007 -7214 -27967 -7180
rect -27933 -7214 -27893 -7180
rect -27859 -7214 -27819 -7180
rect -27785 -7214 -27745 -7180
rect -27711 -7214 -27671 -7180
rect -27637 -7214 -27597 -7180
rect -27563 -7214 -27523 -7180
rect -27489 -7214 -27449 -7180
rect -27415 -7214 -27375 -7180
rect -27341 -7214 -27301 -7180
rect -27267 -7214 -27227 -7180
rect -27193 -7214 -27153 -7180
rect -27119 -7214 -27106 -7180
rect -28202 -7252 -27106 -7214
rect -28202 -7286 -28189 -7252
rect -28155 -7286 -28115 -7252
rect -28081 -7286 -28041 -7252
rect -28007 -7286 -27967 -7252
rect -27933 -7286 -27893 -7252
rect -27859 -7286 -27819 -7252
rect -27785 -7286 -27745 -7252
rect -27711 -7286 -27671 -7252
rect -27637 -7286 -27597 -7252
rect -27563 -7286 -27523 -7252
rect -27489 -7286 -27449 -7252
rect -27415 -7286 -27375 -7252
rect -27341 -7286 -27301 -7252
rect -27267 -7286 -27227 -7252
rect -27193 -7286 -27153 -7252
rect -27119 -7286 -27106 -7252
rect -28202 -7324 -27106 -7286
rect -28202 -7358 -28189 -7324
rect -28155 -7358 -28115 -7324
rect -28081 -7358 -28041 -7324
rect -28007 -7358 -27967 -7324
rect -27933 -7358 -27893 -7324
rect -27859 -7358 -27819 -7324
rect -27785 -7358 -27745 -7324
rect -27711 -7358 -27671 -7324
rect -27637 -7358 -27597 -7324
rect -27563 -7358 -27523 -7324
rect -27489 -7358 -27449 -7324
rect -27415 -7358 -27375 -7324
rect -27341 -7358 -27301 -7324
rect -27267 -7358 -27227 -7324
rect -27193 -7358 -27153 -7324
rect -27119 -7358 -27106 -7324
rect -28202 -7396 -27106 -7358
rect -28202 -7430 -28189 -7396
rect -28155 -7430 -28115 -7396
rect -28081 -7430 -28041 -7396
rect -28007 -7430 -27967 -7396
rect -27933 -7430 -27893 -7396
rect -27859 -7430 -27819 -7396
rect -27785 -7430 -27745 -7396
rect -27711 -7430 -27671 -7396
rect -27637 -7430 -27597 -7396
rect -27563 -7430 -27523 -7396
rect -27489 -7430 -27449 -7396
rect -27415 -7430 -27375 -7396
rect -27341 -7430 -27301 -7396
rect -27267 -7430 -27227 -7396
rect -27193 -7430 -27153 -7396
rect -27119 -7430 -27106 -7396
rect -28202 -7468 -27106 -7430
rect -28202 -7502 -28189 -7468
rect -28155 -7502 -28115 -7468
rect -28081 -7502 -28041 -7468
rect -28007 -7502 -27967 -7468
rect -27933 -7502 -27893 -7468
rect -27859 -7502 -27819 -7468
rect -27785 -7502 -27745 -7468
rect -27711 -7502 -27671 -7468
rect -27637 -7502 -27597 -7468
rect -27563 -7502 -27523 -7468
rect -27489 -7502 -27449 -7468
rect -27415 -7502 -27375 -7468
rect -27341 -7502 -27301 -7468
rect -27267 -7502 -27227 -7468
rect -27193 -7502 -27153 -7468
rect -27119 -7502 -27106 -7468
rect -28202 -7540 -27106 -7502
rect -28202 -7574 -28189 -7540
rect -28155 -7574 -28115 -7540
rect -28081 -7574 -28041 -7540
rect -28007 -7574 -27967 -7540
rect -27933 -7574 -27893 -7540
rect -27859 -7574 -27819 -7540
rect -27785 -7574 -27745 -7540
rect -27711 -7574 -27671 -7540
rect -27637 -7574 -27597 -7540
rect -27563 -7574 -27523 -7540
rect -27489 -7574 -27449 -7540
rect -27415 -7574 -27375 -7540
rect -27341 -7574 -27301 -7540
rect -27267 -7574 -27227 -7540
rect -27193 -7574 -27153 -7540
rect -27119 -7574 -27106 -7540
rect -28202 -7612 -27106 -7574
rect -28202 -7646 -28189 -7612
rect -28155 -7646 -28115 -7612
rect -28081 -7646 -28041 -7612
rect -28007 -7646 -27967 -7612
rect -27933 -7646 -27893 -7612
rect -27859 -7646 -27819 -7612
rect -27785 -7646 -27745 -7612
rect -27711 -7646 -27671 -7612
rect -27637 -7646 -27597 -7612
rect -27563 -7646 -27523 -7612
rect -27489 -7646 -27449 -7612
rect -27415 -7646 -27375 -7612
rect -27341 -7646 -27301 -7612
rect -27267 -7646 -27227 -7612
rect -27193 -7646 -27153 -7612
rect -27119 -7646 -27106 -7612
rect -28202 -7684 -27106 -7646
rect -28202 -7718 -28189 -7684
rect -28155 -7718 -28115 -7684
rect -28081 -7718 -28041 -7684
rect -28007 -7718 -27967 -7684
rect -27933 -7718 -27893 -7684
rect -27859 -7718 -27819 -7684
rect -27785 -7718 -27745 -7684
rect -27711 -7718 -27671 -7684
rect -27637 -7718 -27597 -7684
rect -27563 -7718 -27523 -7684
rect -27489 -7718 -27449 -7684
rect -27415 -7718 -27375 -7684
rect -27341 -7718 -27301 -7684
rect -27267 -7718 -27227 -7684
rect -27193 -7718 -27153 -7684
rect -27119 -7718 -27106 -7684
rect -28202 -7756 -27106 -7718
rect -28202 -7790 -28189 -7756
rect -28155 -7790 -28115 -7756
rect -28081 -7790 -28041 -7756
rect -28007 -7790 -27967 -7756
rect -27933 -7790 -27893 -7756
rect -27859 -7790 -27819 -7756
rect -27785 -7790 -27745 -7756
rect -27711 -7790 -27671 -7756
rect -27637 -7790 -27597 -7756
rect -27563 -7790 -27523 -7756
rect -27489 -7790 -27449 -7756
rect -27415 -7790 -27375 -7756
rect -27341 -7790 -27301 -7756
rect -27267 -7790 -27227 -7756
rect -27193 -7790 -27153 -7756
rect -27119 -7790 -27106 -7756
rect -28202 -7828 -27106 -7790
rect -28202 -7862 -28189 -7828
rect -28155 -7862 -28115 -7828
rect -28081 -7862 -28041 -7828
rect -28007 -7862 -27967 -7828
rect -27933 -7862 -27893 -7828
rect -27859 -7862 -27819 -7828
rect -27785 -7862 -27745 -7828
rect -27711 -7862 -27671 -7828
rect -27637 -7862 -27597 -7828
rect -27563 -7862 -27523 -7828
rect -27489 -7862 -27449 -7828
rect -27415 -7862 -27375 -7828
rect -27341 -7862 -27301 -7828
rect -27267 -7862 -27227 -7828
rect -27193 -7862 -27153 -7828
rect -27119 -7862 -27106 -7828
rect -28202 -7900 -27106 -7862
rect -28202 -7934 -28189 -7900
rect -28155 -7934 -28115 -7900
rect -28081 -7934 -28041 -7900
rect -28007 -7934 -27967 -7900
rect -27933 -7934 -27893 -7900
rect -27859 -7934 -27819 -7900
rect -27785 -7934 -27745 -7900
rect -27711 -7934 -27671 -7900
rect -27637 -7934 -27597 -7900
rect -27563 -7934 -27523 -7900
rect -27489 -7934 -27449 -7900
rect -27415 -7934 -27375 -7900
rect -27341 -7934 -27301 -7900
rect -27267 -7934 -27227 -7900
rect -27193 -7934 -27153 -7900
rect -27119 -7934 -27106 -7900
rect -28202 -7972 -27106 -7934
rect -28202 -8006 -28189 -7972
rect -28155 -8006 -28115 -7972
rect -28081 -8006 -28041 -7972
rect -28007 -8006 -27967 -7972
rect -27933 -8006 -27893 -7972
rect -27859 -8006 -27819 -7972
rect -27785 -8006 -27745 -7972
rect -27711 -8006 -27671 -7972
rect -27637 -8006 -27597 -7972
rect -27563 -8006 -27523 -7972
rect -27489 -8006 -27449 -7972
rect -27415 -8006 -27375 -7972
rect -27341 -8006 -27301 -7972
rect -27267 -8006 -27227 -7972
rect -27193 -8006 -27153 -7972
rect -27119 -8006 -27106 -7972
rect -28202 -8044 -27106 -8006
rect -28202 -8078 -28189 -8044
rect -28155 -8078 -28115 -8044
rect -28081 -8078 -28041 -8044
rect -28007 -8078 -27967 -8044
rect -27933 -8078 -27893 -8044
rect -27859 -8078 -27819 -8044
rect -27785 -8078 -27745 -8044
rect -27711 -8078 -27671 -8044
rect -27637 -8078 -27597 -8044
rect -27563 -8078 -27523 -8044
rect -27489 -8078 -27449 -8044
rect -27415 -8078 -27375 -8044
rect -27341 -8078 -27301 -8044
rect -27267 -8078 -27227 -8044
rect -27193 -8078 -27153 -8044
rect -27119 -8078 -27106 -8044
rect -28202 -8116 -27106 -8078
rect -28202 -8150 -28189 -8116
rect -28155 -8150 -28115 -8116
rect -28081 -8150 -28041 -8116
rect -28007 -8150 -27967 -8116
rect -27933 -8150 -27893 -8116
rect -27859 -8150 -27819 -8116
rect -27785 -8150 -27745 -8116
rect -27711 -8150 -27671 -8116
rect -27637 -8150 -27597 -8116
rect -27563 -8150 -27523 -8116
rect -27489 -8150 -27449 -8116
rect -27415 -8150 -27375 -8116
rect -27341 -8150 -27301 -8116
rect -27267 -8150 -27227 -8116
rect -27193 -8150 -27153 -8116
rect -27119 -8150 -27106 -8116
rect -28202 -8188 -27106 -8150
rect -28202 -8222 -28189 -8188
rect -28155 -8222 -28115 -8188
rect -28081 -8222 -28041 -8188
rect -28007 -8222 -27967 -8188
rect -27933 -8222 -27893 -8188
rect -27859 -8222 -27819 -8188
rect -27785 -8222 -27745 -8188
rect -27711 -8222 -27671 -8188
rect -27637 -8222 -27597 -8188
rect -27563 -8222 -27523 -8188
rect -27489 -8222 -27449 -8188
rect -27415 -8222 -27375 -8188
rect -27341 -8222 -27301 -8188
rect -27267 -8222 -27227 -8188
rect -27193 -8222 -27153 -8188
rect -27119 -8222 -27106 -8188
rect -28202 -8260 -27106 -8222
rect -28202 -8294 -28189 -8260
rect -28155 -8294 -28115 -8260
rect -28081 -8294 -28041 -8260
rect -28007 -8294 -27967 -8260
rect -27933 -8294 -27893 -8260
rect -27859 -8294 -27819 -8260
rect -27785 -8294 -27745 -8260
rect -27711 -8294 -27671 -8260
rect -27637 -8294 -27597 -8260
rect -27563 -8294 -27523 -8260
rect -27489 -8294 -27449 -8260
rect -27415 -8294 -27375 -8260
rect -27341 -8294 -27301 -8260
rect -27267 -8294 -27227 -8260
rect -27193 -8294 -27153 -8260
rect -27119 -8294 -27106 -8260
rect -28202 -8332 -27106 -8294
rect -28202 -8366 -28189 -8332
rect -28155 -8366 -28115 -8332
rect -28081 -8366 -28041 -8332
rect -28007 -8366 -27967 -8332
rect -27933 -8366 -27893 -8332
rect -27859 -8366 -27819 -8332
rect -27785 -8366 -27745 -8332
rect -27711 -8366 -27671 -8332
rect -27637 -8366 -27597 -8332
rect -27563 -8366 -27523 -8332
rect -27489 -8366 -27449 -8332
rect -27415 -8366 -27375 -8332
rect -27341 -8366 -27301 -8332
rect -27267 -8366 -27227 -8332
rect -27193 -8366 -27153 -8332
rect -27119 -8366 -27106 -8332
rect -28202 -8404 -27106 -8366
rect -28202 -8438 -28189 -8404
rect -28155 -8438 -28115 -8404
rect -28081 -8438 -28041 -8404
rect -28007 -8438 -27967 -8404
rect -27933 -8438 -27893 -8404
rect -27859 -8438 -27819 -8404
rect -27785 -8438 -27745 -8404
rect -27711 -8438 -27671 -8404
rect -27637 -8438 -27597 -8404
rect -27563 -8438 -27523 -8404
rect -27489 -8438 -27449 -8404
rect -27415 -8438 -27375 -8404
rect -27341 -8438 -27301 -8404
rect -27267 -8438 -27227 -8404
rect -27193 -8438 -27153 -8404
rect -27119 -8438 -27106 -8404
rect -28202 -8476 -27106 -8438
rect -28202 -8510 -28189 -8476
rect -28155 -8510 -28115 -8476
rect -28081 -8510 -28041 -8476
rect -28007 -8510 -27967 -8476
rect -27933 -8510 -27893 -8476
rect -27859 -8510 -27819 -8476
rect -27785 -8510 -27745 -8476
rect -27711 -8510 -27671 -8476
rect -27637 -8510 -27597 -8476
rect -27563 -8510 -27523 -8476
rect -27489 -8510 -27449 -8476
rect -27415 -8510 -27375 -8476
rect -27341 -8510 -27301 -8476
rect -27267 -8510 -27227 -8476
rect -27193 -8510 -27153 -8476
rect -27119 -8510 -27106 -8476
rect -28202 -8548 -27106 -8510
rect -28202 -8582 -28189 -8548
rect -28155 -8582 -28115 -8548
rect -28081 -8582 -28041 -8548
rect -28007 -8582 -27967 -8548
rect -27933 -8582 -27893 -8548
rect -27859 -8582 -27819 -8548
rect -27785 -8582 -27745 -8548
rect -27711 -8582 -27671 -8548
rect -27637 -8582 -27597 -8548
rect -27563 -8582 -27523 -8548
rect -27489 -8582 -27449 -8548
rect -27415 -8582 -27375 -8548
rect -27341 -8582 -27301 -8548
rect -27267 -8582 -27227 -8548
rect -27193 -8582 -27153 -8548
rect -27119 -8582 -27106 -8548
rect -28202 -8620 -27106 -8582
rect -28202 -8654 -28189 -8620
rect -28155 -8654 -28115 -8620
rect -28081 -8654 -28041 -8620
rect -28007 -8654 -27967 -8620
rect -27933 -8654 -27893 -8620
rect -27859 -8654 -27819 -8620
rect -27785 -8654 -27745 -8620
rect -27711 -8654 -27671 -8620
rect -27637 -8654 -27597 -8620
rect -27563 -8654 -27523 -8620
rect -27489 -8654 -27449 -8620
rect -27415 -8654 -27375 -8620
rect -27341 -8654 -27301 -8620
rect -27267 -8654 -27227 -8620
rect -27193 -8654 -27153 -8620
rect -27119 -8654 -27106 -8620
rect -28202 -8692 -27106 -8654
rect -28202 -8726 -28189 -8692
rect -28155 -8726 -28115 -8692
rect -28081 -8726 -28041 -8692
rect -28007 -8726 -27967 -8692
rect -27933 -8726 -27893 -8692
rect -27859 -8726 -27819 -8692
rect -27785 -8726 -27745 -8692
rect -27711 -8726 -27671 -8692
rect -27637 -8726 -27597 -8692
rect -27563 -8726 -27523 -8692
rect -27489 -8726 -27449 -8692
rect -27415 -8726 -27375 -8692
rect -27341 -8726 -27301 -8692
rect -27267 -8726 -27227 -8692
rect -27193 -8726 -27153 -8692
rect -27119 -8726 -27106 -8692
rect -28202 -8764 -27106 -8726
rect -28202 -8798 -28189 -8764
rect -28155 -8798 -28115 -8764
rect -28081 -8798 -28041 -8764
rect -28007 -8798 -27967 -8764
rect -27933 -8798 -27893 -8764
rect -27859 -8798 -27819 -8764
rect -27785 -8798 -27745 -8764
rect -27711 -8798 -27671 -8764
rect -27637 -8798 -27597 -8764
rect -27563 -8798 -27523 -8764
rect -27489 -8798 -27449 -8764
rect -27415 -8798 -27375 -8764
rect -27341 -8798 -27301 -8764
rect -27267 -8798 -27227 -8764
rect -27193 -8798 -27153 -8764
rect -27119 -8798 -27106 -8764
tri -11546 -2131 -11507 -2092 se
rect -11507 -2131 -11480 -2092
tri -11480 -2131 -11441 -2092 nw
rect -11546 -8658 -11500 -2131
tri -11500 -2151 -11480 -2131 nw
rect -11546 -8692 -11540 -8658
rect -11506 -8692 -11500 -8658
rect -11546 -8730 -11500 -8692
rect -11546 -8764 -11540 -8730
rect -11506 -8764 -11500 -8730
rect -11546 -8776 -11500 -8764
rect -28202 -8836 -27106 -8798
rect -28202 -8870 -28189 -8836
rect -28155 -8870 -28115 -8836
rect -28081 -8870 -28041 -8836
rect -28007 -8870 -27967 -8836
rect -27933 -8870 -27893 -8836
rect -27859 -8870 -27819 -8836
rect -27785 -8870 -27745 -8836
rect -27711 -8870 -27671 -8836
rect -27637 -8870 -27597 -8836
rect -27563 -8870 -27523 -8836
rect -27489 -8870 -27449 -8836
rect -27415 -8870 -27375 -8836
rect -27341 -8870 -27301 -8836
rect -27267 -8870 -27227 -8836
rect -27193 -8870 -27153 -8836
rect -27119 -8870 -27106 -8836
rect -28202 -8908 -27106 -8870
rect -28202 -8942 -28189 -8908
rect -28155 -8942 -28115 -8908
rect -28081 -8942 -28041 -8908
rect -28007 -8942 -27967 -8908
rect -27933 -8942 -27893 -8908
rect -27859 -8942 -27819 -8908
rect -27785 -8942 -27745 -8908
rect -27711 -8942 -27671 -8908
rect -27637 -8942 -27597 -8908
rect -27563 -8942 -27523 -8908
rect -27489 -8942 -27449 -8908
rect -27415 -8942 -27375 -8908
rect -27341 -8942 -27301 -8908
rect -27267 -8942 -27227 -8908
rect -27193 -8942 -27153 -8908
rect -27119 -8942 -27106 -8908
rect -28202 -8980 -27106 -8942
rect -28202 -9014 -28189 -8980
rect -28155 -9014 -28115 -8980
rect -28081 -9014 -28041 -8980
rect -28007 -9014 -27967 -8980
rect -27933 -9014 -27893 -8980
rect -27859 -9014 -27819 -8980
rect -27785 -9014 -27745 -8980
rect -27711 -9014 -27671 -8980
rect -27637 -9014 -27597 -8980
rect -27563 -9014 -27523 -8980
rect -27489 -9014 -27449 -8980
rect -27415 -9014 -27375 -8980
rect -27341 -9014 -27301 -8980
rect -27267 -9014 -27227 -8980
rect -27193 -9014 -27153 -8980
rect -27119 -9014 -27106 -8980
rect -28202 -9052 -27106 -9014
rect -28202 -9086 -28189 -9052
rect -28155 -9086 -28115 -9052
rect -28081 -9086 -28041 -9052
rect -28007 -9086 -27967 -9052
rect -27933 -9086 -27893 -9052
rect -27859 -9086 -27819 -9052
rect -27785 -9086 -27745 -9052
rect -27711 -9086 -27671 -9052
rect -27637 -9086 -27597 -9052
rect -27563 -9086 -27523 -9052
rect -27489 -9086 -27449 -9052
rect -27415 -9086 -27375 -9052
rect -27341 -9086 -27301 -9052
rect -27267 -9086 -27227 -9052
rect -27193 -9086 -27153 -9052
rect -27119 -9086 -27106 -9052
rect -28202 -9124 -27106 -9086
rect -28202 -9158 -28189 -9124
rect -28155 -9158 -28115 -9124
rect -28081 -9158 -28041 -9124
rect -28007 -9158 -27967 -9124
rect -27933 -9158 -27893 -9124
rect -27859 -9158 -27819 -9124
rect -27785 -9158 -27745 -9124
rect -27711 -9158 -27671 -9124
rect -27637 -9158 -27597 -9124
rect -27563 -9158 -27523 -9124
rect -27489 -9158 -27449 -9124
rect -27415 -9158 -27375 -9124
rect -27341 -9158 -27301 -9124
rect -27267 -9158 -27227 -9124
rect -27193 -9158 -27153 -9124
rect -27119 -9158 -27106 -9124
rect -28202 -9196 -27106 -9158
rect -28202 -9230 -28189 -9196
rect -28155 -9230 -28115 -9196
rect -28081 -9230 -28041 -9196
rect -28007 -9230 -27967 -9196
rect -27933 -9230 -27893 -9196
rect -27859 -9230 -27819 -9196
rect -27785 -9230 -27745 -9196
rect -27711 -9230 -27671 -9196
rect -27637 -9230 -27597 -9196
rect -27563 -9230 -27523 -9196
rect -27489 -9230 -27449 -9196
rect -27415 -9230 -27375 -9196
rect -27341 -9230 -27301 -9196
rect -27267 -9230 -27227 -9196
rect -27193 -9230 -27153 -9196
rect -27119 -9230 -27106 -9196
rect -28202 -9268 -27106 -9230
rect -28202 -9302 -28189 -9268
rect -28155 -9302 -28115 -9268
rect -28081 -9302 -28041 -9268
rect -28007 -9302 -27967 -9268
rect -27933 -9302 -27893 -9268
rect -27859 -9302 -27819 -9268
rect -27785 -9302 -27745 -9268
rect -27711 -9302 -27671 -9268
rect -27637 -9302 -27597 -9268
rect -27563 -9302 -27523 -9268
rect -27489 -9302 -27449 -9268
rect -27415 -9302 -27375 -9268
rect -27341 -9302 -27301 -9268
rect -27267 -9302 -27227 -9268
rect -27193 -9302 -27153 -9268
rect -27119 -9302 -27106 -9268
rect -28202 -9340 -27106 -9302
rect -28202 -9374 -28189 -9340
rect -28155 -9374 -28115 -9340
rect -28081 -9374 -28041 -9340
rect -28007 -9374 -27967 -9340
rect -27933 -9374 -27893 -9340
rect -27859 -9374 -27819 -9340
rect -27785 -9374 -27745 -9340
rect -27711 -9374 -27671 -9340
rect -27637 -9374 -27597 -9340
rect -27563 -9374 -27523 -9340
rect -27489 -9374 -27449 -9340
rect -27415 -9374 -27375 -9340
rect -27341 -9374 -27301 -9340
rect -27267 -9374 -27227 -9340
rect -27193 -9374 -27153 -9340
rect -27119 -9374 -27106 -9340
rect -28202 -9386 -27106 -9374
rect -30792 -9422 -29134 -9417
rect -30792 -9456 -30753 -9422
rect -30719 -9456 -30680 -9422
rect -30646 -9456 -30607 -9422
rect -30573 -9456 -30534 -9422
rect -30500 -9456 -30461 -9422
rect -30427 -9456 -30388 -9422
rect -30354 -9456 -30315 -9422
rect -30281 -9456 -30242 -9422
rect -30208 -9456 -30169 -9422
rect -30135 -9456 -30096 -9422
rect -30062 -9456 -30023 -9422
rect -29989 -9456 -29950 -9422
rect -29916 -9456 -29877 -9422
rect -29843 -9456 -29804 -9422
rect -29770 -9456 -29731 -9422
rect -29697 -9456 -29658 -9422
rect -29624 -9456 -29585 -9422
rect -29551 -9456 -29512 -9422
rect -29478 -9456 -29439 -9422
rect -29405 -9456 -29366 -9422
rect -29332 -9456 -29293 -9422
rect -29259 -9456 -29220 -9422
rect -29186 -9451 -29134 -9422
rect -29100 -9451 -29046 -9417
rect -29012 -9451 -28958 -9417
rect -28924 -9451 -28870 -9417
rect -28836 -9451 -28830 -9417
rect -29186 -9456 -28830 -9451
rect -30792 -9489 -28830 -9456
rect -30792 -9494 -29134 -9489
rect -30792 -9528 -30753 -9494
rect -30719 -9528 -30680 -9494
rect -30646 -9528 -30607 -9494
rect -30573 -9528 -30534 -9494
rect -30500 -9528 -30461 -9494
rect -30427 -9528 -30388 -9494
rect -30354 -9528 -30315 -9494
rect -30281 -9528 -30242 -9494
rect -30208 -9528 -30169 -9494
rect -30135 -9528 -30096 -9494
rect -30062 -9528 -30023 -9494
rect -29989 -9528 -29950 -9494
rect -29916 -9528 -29877 -9494
rect -29843 -9528 -29804 -9494
rect -29770 -9528 -29731 -9494
rect -29697 -9528 -29658 -9494
rect -29624 -9528 -29585 -9494
rect -29551 -9528 -29512 -9494
rect -29478 -9528 -29439 -9494
rect -29405 -9528 -29366 -9494
rect -29332 -9528 -29293 -9494
rect -29259 -9528 -29220 -9494
rect -29186 -9523 -29134 -9494
rect -29100 -9523 -29046 -9489
rect -29012 -9523 -28958 -9489
rect -28924 -9523 -28870 -9489
rect -28836 -9523 -28830 -9489
rect -29186 -9528 -28830 -9523
rect -30792 -9561 -28830 -9528
rect -30792 -9566 -29134 -9561
rect -30792 -9600 -30753 -9566
rect -30719 -9600 -30680 -9566
rect -30646 -9600 -30607 -9566
rect -30573 -9600 -30534 -9566
rect -30500 -9600 -30461 -9566
rect -30427 -9600 -30388 -9566
rect -30354 -9600 -30315 -9566
rect -30281 -9600 -30242 -9566
rect -30208 -9600 -30169 -9566
rect -30135 -9600 -30096 -9566
rect -30062 -9600 -30023 -9566
rect -29989 -9600 -29950 -9566
rect -29916 -9600 -29877 -9566
rect -29843 -9600 -29804 -9566
rect -29770 -9600 -29731 -9566
rect -29697 -9600 -29658 -9566
rect -29624 -9600 -29585 -9566
rect -29551 -9600 -29512 -9566
rect -29478 -9600 -29439 -9566
rect -29405 -9600 -29366 -9566
rect -29332 -9600 -29293 -9566
rect -29259 -9600 -29220 -9566
rect -29186 -9595 -29134 -9566
rect -29100 -9595 -29046 -9561
rect -29012 -9595 -28958 -9561
rect -28924 -9595 -28870 -9561
rect -28836 -9595 -28830 -9561
rect -29186 -9600 -28830 -9595
rect -32350 -9607 -28830 -9600
<< via1 >>
rect -28196 4843 -28144 4895
rect -28132 4843 -28080 4895
rect -28068 4843 -28016 4895
rect -28004 4843 -27952 4895
rect -27940 4843 -27888 4895
rect -27876 4843 -27824 4895
rect -27812 4843 -27760 4895
rect -27748 4843 -27696 4895
rect -27684 4843 -27632 4895
rect -27620 4843 -27568 4895
rect -27555 4843 -27503 4895
rect -27490 4843 -27438 4895
rect -27425 4843 -27373 4895
rect -27360 4843 -27308 4895
rect -27295 4843 -27243 4895
rect -27230 4843 -27178 4895
rect -27165 4843 -27113 4895
rect -28196 4721 -28144 4773
rect -28132 4721 -28080 4773
rect -28068 4721 -28016 4773
rect -28004 4721 -27952 4773
rect -27940 4721 -27888 4773
rect -27876 4721 -27824 4773
rect -27812 4721 -27760 4773
rect -27748 4721 -27696 4773
rect -27684 4721 -27632 4773
rect -27620 4721 -27568 4773
rect -27555 4721 -27503 4773
rect -27490 4721 -27438 4773
rect -27425 4721 -27373 4773
rect -27360 4721 -27308 4773
rect -27295 4721 -27243 4773
rect -27230 4721 -27178 4773
rect -27165 4721 -27113 4773
rect -32338 466 -32286 501
rect -32338 449 -32310 466
rect -32310 449 -32286 466
rect -32273 466 -32221 501
rect -32273 449 -32266 466
rect -32266 449 -32232 466
rect -32232 449 -32221 466
rect -32208 466 -32156 501
rect -32143 466 -32091 501
rect -32078 466 -32026 501
rect -32013 466 -31961 501
rect -31948 466 -31896 501
rect -32208 449 -32188 466
rect -32188 449 -32156 466
rect -32143 449 -32110 466
rect -32110 449 -32091 466
rect -32078 449 -32076 466
rect -32076 449 -32032 466
rect -32032 449 -32026 466
rect -32013 449 -31998 466
rect -31998 449 -31961 466
rect -31948 449 -31920 466
rect -31920 449 -31896 466
rect -31882 466 -31830 501
rect -31882 449 -31876 466
rect -31876 449 -31842 466
rect -31842 449 -31830 466
rect -31816 466 -31764 501
rect -31816 449 -31798 466
rect -31798 449 -31764 466
rect -32338 432 -32310 437
rect -32310 432 -32286 437
rect -32338 394 -32286 432
rect -32338 385 -32310 394
rect -32310 385 -32286 394
rect -32273 432 -32266 437
rect -32266 432 -32232 437
rect -32232 432 -32221 437
rect -32273 394 -32221 432
rect -32273 385 -32266 394
rect -32266 385 -32232 394
rect -32232 385 -32221 394
rect -32208 432 -32188 437
rect -32188 432 -32156 437
rect -32143 432 -32110 437
rect -32110 432 -32091 437
rect -32078 432 -32076 437
rect -32076 432 -32032 437
rect -32032 432 -32026 437
rect -32013 432 -31998 437
rect -31998 432 -31961 437
rect -31948 432 -31920 437
rect -31920 432 -31896 437
rect -32208 394 -32156 432
rect -32143 394 -32091 432
rect -32078 394 -32026 432
rect -32013 394 -31961 432
rect -31948 394 -31896 432
rect -32208 385 -32188 394
rect -32188 385 -32156 394
rect -32143 385 -32110 394
rect -32110 385 -32091 394
rect -32078 385 -32076 394
rect -32076 385 -32032 394
rect -32032 385 -32026 394
rect -32013 385 -31998 394
rect -31998 385 -31961 394
rect -31948 385 -31920 394
rect -31920 385 -31896 394
rect -31882 432 -31876 437
rect -31876 432 -31842 437
rect -31842 432 -31830 437
rect -31882 394 -31830 432
rect -31882 385 -31876 394
rect -31876 385 -31842 394
rect -31842 385 -31830 394
rect -31816 432 -31798 437
rect -31798 432 -31764 437
rect -31816 394 -31764 432
rect -31816 385 -31798 394
rect -31798 385 -31764 394
rect -32338 360 -32310 373
rect -32310 360 -32286 373
rect -32338 322 -32286 360
rect -32338 321 -32310 322
rect -32310 321 -32286 322
rect -32273 360 -32266 373
rect -32266 360 -32232 373
rect -32232 360 -32221 373
rect -32273 322 -32221 360
rect -32273 321 -32266 322
rect -32266 321 -32232 322
rect -32232 321 -32221 322
rect -32208 360 -32188 373
rect -32188 360 -32156 373
rect -32143 360 -32110 373
rect -32110 360 -32091 373
rect -32078 360 -32076 373
rect -32076 360 -32032 373
rect -32032 360 -32026 373
rect -32013 360 -31998 373
rect -31998 360 -31961 373
rect -31948 360 -31920 373
rect -31920 360 -31896 373
rect -32208 322 -32156 360
rect -32143 322 -32091 360
rect -32078 322 -32026 360
rect -32013 322 -31961 360
rect -31948 322 -31896 360
rect -32208 321 -32188 322
rect -32188 321 -32156 322
rect -32143 321 -32110 322
rect -32110 321 -32091 322
rect -32078 321 -32076 322
rect -32076 321 -32032 322
rect -32032 321 -32026 322
rect -32013 321 -31998 322
rect -31998 321 -31961 322
rect -31948 321 -31920 322
rect -31920 321 -31896 322
rect -31882 360 -31876 373
rect -31876 360 -31842 373
rect -31842 360 -31830 373
rect -31882 322 -31830 360
rect -31882 321 -31876 322
rect -31876 321 -31842 322
rect -31842 321 -31830 322
rect -31816 360 -31798 373
rect -31798 360 -31764 373
rect -31816 322 -31764 360
rect -31816 321 -31798 322
rect -31798 321 -31764 322
rect -32338 288 -32310 309
rect -32310 288 -32286 309
rect -32338 257 -32286 288
rect -32273 288 -32266 309
rect -32266 288 -32232 309
rect -32232 288 -32221 309
rect -32273 257 -32221 288
rect -32208 288 -32188 309
rect -32188 288 -32156 309
rect -32143 288 -32110 309
rect -32110 288 -32091 309
rect -32078 288 -32076 309
rect -32076 288 -32032 309
rect -32032 288 -32026 309
rect -32013 288 -31998 309
rect -31998 288 -31961 309
rect -31948 288 -31920 309
rect -31920 288 -31896 309
rect -32208 257 -32156 288
rect -32143 257 -32091 288
rect -32078 257 -32026 288
rect -32013 257 -31961 288
rect -31948 257 -31896 288
rect -31882 288 -31876 309
rect -31876 288 -31842 309
rect -31842 288 -31830 309
rect -31882 257 -31830 288
rect -31816 288 -31798 309
rect -31798 288 -31764 309
rect -31816 257 -31764 288
rect -32338 216 -32310 245
rect -32310 216 -32286 245
rect -32338 193 -32286 216
rect -32273 216 -32266 245
rect -32266 216 -32232 245
rect -32232 216 -32221 245
rect -32273 193 -32221 216
rect -32208 216 -32188 245
rect -32188 216 -32156 245
rect -32143 216 -32110 245
rect -32110 216 -32091 245
rect -32078 216 -32076 245
rect -32076 216 -32032 245
rect -32032 216 -32026 245
rect -32013 216 -31998 245
rect -31998 216 -31961 245
rect -31948 216 -31920 245
rect -31920 216 -31896 245
rect -32208 193 -32156 216
rect -32143 193 -32091 216
rect -32078 193 -32026 216
rect -32013 193 -31961 216
rect -31948 193 -31896 216
rect -31882 216 -31876 245
rect -31876 216 -31842 245
rect -31842 216 -31830 245
rect -31882 193 -31830 216
rect -31816 216 -31798 245
rect -31798 216 -31764 245
rect -31816 193 -31764 216
rect -32338 178 -32286 181
rect -32338 144 -32310 178
rect -32310 144 -32286 178
rect -32338 129 -32286 144
rect -32273 178 -32221 181
rect -32273 144 -32266 178
rect -32266 144 -32232 178
rect -32232 144 -32221 178
rect -32273 129 -32221 144
rect -32208 178 -32156 181
rect -32143 178 -32091 181
rect -32078 178 -32026 181
rect -32013 178 -31961 181
rect -31948 178 -31896 181
rect -32208 144 -32188 178
rect -32188 144 -32156 178
rect -32143 144 -32110 178
rect -32110 144 -32091 178
rect -32078 144 -32076 178
rect -32076 144 -32032 178
rect -32032 144 -32026 178
rect -32013 144 -31998 178
rect -31998 144 -31961 178
rect -31948 144 -31920 178
rect -31920 144 -31896 178
rect -32208 129 -32156 144
rect -32143 129 -32091 144
rect -32078 129 -32026 144
rect -32013 129 -31961 144
rect -31948 129 -31896 144
rect -31882 178 -31830 181
rect -31882 144 -31876 178
rect -31876 144 -31842 178
rect -31842 144 -31830 178
rect -31882 129 -31830 144
rect -31816 178 -31764 181
rect -31816 144 -31798 178
rect -31798 144 -31764 178
rect -31816 129 -31764 144
rect -32338 106 -32286 117
rect -32338 72 -32310 106
rect -32310 72 -32286 106
rect -32338 65 -32286 72
rect -32273 106 -32221 117
rect -32273 72 -32266 106
rect -32266 72 -32232 106
rect -32232 72 -32221 106
rect -32273 65 -32221 72
rect -32208 106 -32156 117
rect -32143 106 -32091 117
rect -32078 106 -32026 117
rect -32013 106 -31961 117
rect -31948 106 -31896 117
rect -32208 72 -32188 106
rect -32188 72 -32156 106
rect -32143 72 -32110 106
rect -32110 72 -32091 106
rect -32078 72 -32076 106
rect -32076 72 -32032 106
rect -32032 72 -32026 106
rect -32013 72 -31998 106
rect -31998 72 -31961 106
rect -31948 72 -31920 106
rect -31920 72 -31896 106
rect -32208 65 -32156 72
rect -32143 65 -32091 72
rect -32078 65 -32026 72
rect -32013 65 -31961 72
rect -31948 65 -31896 72
rect -31882 106 -31830 117
rect -31882 72 -31876 106
rect -31876 72 -31842 106
rect -31842 72 -31830 106
rect -31882 65 -31830 72
rect -31816 106 -31764 117
rect -31816 72 -31798 106
rect -31798 72 -31764 106
rect -31816 65 -31764 72
rect -32338 34 -32286 53
rect -32338 1 -32310 34
rect -32310 1 -32286 34
rect -32273 34 -32221 53
rect -32273 1 -32266 34
rect -32266 1 -32232 34
rect -32232 1 -32221 34
rect -32208 34 -32156 53
rect -32143 34 -32091 53
rect -32078 34 -32026 53
rect -32013 34 -31961 53
rect -31948 34 -31896 53
rect -32208 1 -32188 34
rect -32188 1 -32156 34
rect -32143 1 -32110 34
rect -32110 1 -32091 34
rect -32078 1 -32076 34
rect -32076 1 -32032 34
rect -32032 1 -32026 34
rect -32013 1 -31998 34
rect -31998 1 -31961 34
rect -31948 1 -31920 34
rect -31920 1 -31896 34
rect -31882 34 -31830 53
rect -31882 1 -31876 34
rect -31876 1 -31842 34
rect -31842 1 -31830 34
rect -31816 34 -31764 53
rect -31816 1 -31798 34
rect -31798 1 -31764 34
rect -32338 -38 -32286 -11
rect -32338 -63 -32310 -38
rect -32310 -63 -32286 -38
rect -32273 -38 -32221 -11
rect -32273 -63 -32266 -38
rect -32266 -63 -32232 -38
rect -32232 -63 -32221 -38
rect -32208 -38 -32156 -11
rect -32143 -38 -32091 -11
rect -32078 -38 -32026 -11
rect -32013 -38 -31961 -11
rect -31948 -38 -31896 -11
rect -32208 -63 -32188 -38
rect -32188 -63 -32156 -38
rect -32143 -63 -32110 -38
rect -32110 -63 -32091 -38
rect -32078 -63 -32076 -38
rect -32076 -63 -32032 -38
rect -32032 -63 -32026 -38
rect -32013 -63 -31998 -38
rect -31998 -63 -31961 -38
rect -31948 -63 -31920 -38
rect -31920 -63 -31896 -38
rect -31882 -38 -31830 -11
rect -31882 -63 -31876 -38
rect -31876 -63 -31842 -38
rect -31842 -63 -31830 -38
rect -31816 -38 -31764 -11
rect -31816 -63 -31798 -38
rect -31798 -63 -31764 -38
rect -32338 -110 -32286 -75
rect -32338 -127 -32310 -110
rect -32310 -127 -32286 -110
rect -32273 -110 -32221 -75
rect -32273 -127 -32266 -110
rect -32266 -127 -32232 -110
rect -32232 -127 -32221 -110
rect -32208 -110 -32156 -75
rect -32143 -110 -32091 -75
rect -32078 -110 -32026 -75
rect -32013 -110 -31961 -75
rect -31948 -110 -31896 -75
rect -32208 -127 -32188 -110
rect -32188 -127 -32156 -110
rect -32143 -127 -32110 -110
rect -32110 -127 -32091 -110
rect -32078 -127 -32076 -110
rect -32076 -127 -32032 -110
rect -32032 -127 -32026 -110
rect -32013 -127 -31998 -110
rect -31998 -127 -31961 -110
rect -31948 -127 -31920 -110
rect -31920 -127 -31896 -110
rect -31882 -110 -31830 -75
rect -31882 -127 -31876 -110
rect -31876 -127 -31842 -110
rect -31842 -127 -31830 -110
rect -31816 -110 -31764 -75
rect -31816 -127 -31798 -110
rect -31798 -127 -31764 -110
rect -32338 -144 -32310 -139
rect -32310 -144 -32286 -139
rect -32338 -182 -32286 -144
rect -32338 -191 -32310 -182
rect -32310 -191 -32286 -182
rect -32273 -144 -32266 -139
rect -32266 -144 -32232 -139
rect -32232 -144 -32221 -139
rect -32273 -182 -32221 -144
rect -32273 -191 -32266 -182
rect -32266 -191 -32232 -182
rect -32232 -191 -32221 -182
rect -32208 -144 -32188 -139
rect -32188 -144 -32156 -139
rect -32143 -144 -32110 -139
rect -32110 -144 -32091 -139
rect -32078 -144 -32076 -139
rect -32076 -144 -32032 -139
rect -32032 -144 -32026 -139
rect -32013 -144 -31998 -139
rect -31998 -144 -31961 -139
rect -31948 -144 -31920 -139
rect -31920 -144 -31896 -139
rect -32208 -182 -32156 -144
rect -32143 -182 -32091 -144
rect -32078 -182 -32026 -144
rect -32013 -182 -31961 -144
rect -31948 -182 -31896 -144
rect -32208 -191 -32188 -182
rect -32188 -191 -32156 -182
rect -32143 -191 -32110 -182
rect -32110 -191 -32091 -182
rect -32078 -191 -32076 -182
rect -32076 -191 -32032 -182
rect -32032 -191 -32026 -182
rect -32013 -191 -31998 -182
rect -31998 -191 -31961 -182
rect -31948 -191 -31920 -182
rect -31920 -191 -31896 -182
rect -31882 -144 -31876 -139
rect -31876 -144 -31842 -139
rect -31842 -144 -31830 -139
rect -31882 -182 -31830 -144
rect -31882 -191 -31876 -182
rect -31876 -191 -31842 -182
rect -31842 -191 -31830 -182
rect -31816 -144 -31798 -139
rect -31798 -144 -31764 -139
rect -31816 -182 -31764 -144
rect -31816 -191 -31798 -182
rect -31798 -191 -31764 -182
rect -32338 -216 -32310 -203
rect -32310 -216 -32286 -203
rect -32338 -254 -32286 -216
rect -32338 -255 -32310 -254
rect -32310 -255 -32286 -254
rect -32273 -216 -32266 -203
rect -32266 -216 -32232 -203
rect -32232 -216 -32221 -203
rect -32273 -254 -32221 -216
rect -32273 -255 -32266 -254
rect -32266 -255 -32232 -254
rect -32232 -255 -32221 -254
rect -32208 -216 -32188 -203
rect -32188 -216 -32156 -203
rect -32143 -216 -32110 -203
rect -32110 -216 -32091 -203
rect -32078 -216 -32076 -203
rect -32076 -216 -32032 -203
rect -32032 -216 -32026 -203
rect -32013 -216 -31998 -203
rect -31998 -216 -31961 -203
rect -31948 -216 -31920 -203
rect -31920 -216 -31896 -203
rect -32208 -254 -32156 -216
rect -32143 -254 -32091 -216
rect -32078 -254 -32026 -216
rect -32013 -254 -31961 -216
rect -31948 -254 -31896 -216
rect -32208 -255 -32188 -254
rect -32188 -255 -32156 -254
rect -32143 -255 -32110 -254
rect -32110 -255 -32091 -254
rect -32078 -255 -32076 -254
rect -32076 -255 -32032 -254
rect -32032 -255 -32026 -254
rect -32013 -255 -31998 -254
rect -31998 -255 -31961 -254
rect -31948 -255 -31920 -254
rect -31920 -255 -31896 -254
rect -31882 -216 -31876 -203
rect -31876 -216 -31842 -203
rect -31842 -216 -31830 -203
rect -31882 -254 -31830 -216
rect -31882 -255 -31876 -254
rect -31876 -255 -31842 -254
rect -31842 -255 -31830 -254
rect -31816 -216 -31798 -203
rect -31798 -216 -31764 -203
rect -31816 -254 -31764 -216
rect -31816 -255 -31798 -254
rect -31798 -255 -31764 -254
rect -32338 -288 -32310 -267
rect -32310 -288 -32286 -267
rect -32338 -319 -32286 -288
rect -32273 -288 -32266 -267
rect -32266 -288 -32232 -267
rect -32232 -288 -32221 -267
rect -32273 -319 -32221 -288
rect -32208 -288 -32188 -267
rect -32188 -288 -32156 -267
rect -32143 -288 -32110 -267
rect -32110 -288 -32091 -267
rect -32078 -288 -32076 -267
rect -32076 -288 -32032 -267
rect -32032 -288 -32026 -267
rect -32013 -288 -31998 -267
rect -31998 -288 -31961 -267
rect -31948 -288 -31920 -267
rect -31920 -288 -31896 -267
rect -32208 -319 -32156 -288
rect -32143 -319 -32091 -288
rect -32078 -319 -32026 -288
rect -32013 -319 -31961 -288
rect -31948 -319 -31896 -288
rect -31882 -288 -31876 -267
rect -31876 -288 -31842 -267
rect -31842 -288 -31830 -267
rect -31882 -319 -31830 -288
rect -31816 -288 -31798 -267
rect -31798 -288 -31764 -267
rect -31816 -319 -31764 -288
rect -32338 -360 -32310 -331
rect -32310 -360 -32286 -331
rect -32338 -383 -32286 -360
rect -32273 -360 -32266 -331
rect -32266 -360 -32232 -331
rect -32232 -360 -32221 -331
rect -32273 -383 -32221 -360
rect -32208 -360 -32188 -331
rect -32188 -360 -32156 -331
rect -32143 -360 -32110 -331
rect -32110 -360 -32091 -331
rect -32078 -360 -32076 -331
rect -32076 -360 -32032 -331
rect -32032 -360 -32026 -331
rect -32013 -360 -31998 -331
rect -31998 -360 -31961 -331
rect -31948 -360 -31920 -331
rect -31920 -360 -31896 -331
rect -32208 -383 -32156 -360
rect -32143 -383 -32091 -360
rect -32078 -383 -32026 -360
rect -32013 -383 -31961 -360
rect -31948 -383 -31896 -360
rect -31882 -360 -31876 -331
rect -31876 -360 -31842 -331
rect -31842 -360 -31830 -331
rect -31882 -383 -31830 -360
rect -31816 -360 -31798 -331
rect -31798 -360 -31764 -331
rect -31816 -383 -31764 -360
rect -29135 464 -29083 495
rect -29135 443 -29134 464
rect -29134 443 -29100 464
rect -29100 443 -29083 464
rect -29053 464 -29001 495
rect -29053 443 -29046 464
rect -29046 443 -29012 464
rect -29012 443 -29001 464
rect -28971 464 -28919 495
rect -28971 443 -28958 464
rect -28958 443 -28924 464
rect -28924 443 -28919 464
rect -28889 464 -28837 495
rect -28889 443 -28870 464
rect -28870 443 -28837 464
rect -29135 391 -29083 430
rect -29135 378 -29134 391
rect -29134 378 -29100 391
rect -29100 378 -29083 391
rect -29053 391 -29001 430
rect -29053 378 -29046 391
rect -29046 378 -29012 391
rect -29012 378 -29001 391
rect -28971 391 -28919 430
rect -28971 378 -28958 391
rect -28958 378 -28924 391
rect -28924 378 -28919 391
rect -28889 391 -28837 430
rect -28889 378 -28870 391
rect -28870 378 -28837 391
rect -29135 357 -29134 365
rect -29134 357 -29100 365
rect -29100 357 -29083 365
rect -29135 318 -29083 357
rect -29135 313 -29134 318
rect -29134 313 -29100 318
rect -29100 313 -29083 318
rect -29053 357 -29046 365
rect -29046 357 -29012 365
rect -29012 357 -29001 365
rect -29053 318 -29001 357
rect -29053 313 -29046 318
rect -29046 313 -29012 318
rect -29012 313 -29001 318
rect -28971 357 -28958 365
rect -28958 357 -28924 365
rect -28924 357 -28919 365
rect -28971 318 -28919 357
rect -28971 313 -28958 318
rect -28958 313 -28924 318
rect -28924 313 -28919 318
rect -28889 357 -28870 365
rect -28870 357 -28837 365
rect -28889 318 -28837 357
rect -28889 313 -28870 318
rect -28870 313 -28837 318
rect -29135 284 -29134 301
rect -29134 284 -29100 301
rect -29100 284 -29083 301
rect -29135 249 -29083 284
rect -29053 284 -29046 301
rect -29046 284 -29012 301
rect -29012 284 -29001 301
rect -29053 249 -29001 284
rect -28971 284 -28958 301
rect -28958 284 -28924 301
rect -28924 284 -28919 301
rect -28971 249 -28919 284
rect -28889 284 -28870 301
rect -28870 284 -28837 301
rect -28889 249 -28837 284
rect -29135 211 -29134 237
rect -29134 211 -29100 237
rect -29100 211 -29083 237
rect -29135 185 -29083 211
rect -29053 211 -29046 237
rect -29046 211 -29012 237
rect -29012 211 -29001 237
rect -29053 185 -29001 211
rect -28971 211 -28958 237
rect -28958 211 -28924 237
rect -28924 211 -28919 237
rect -28971 185 -28919 211
rect -28889 211 -28870 237
rect -28870 211 -28837 237
rect -28889 185 -28837 211
rect -29135 172 -29083 173
rect -29135 138 -29134 172
rect -29134 138 -29100 172
rect -29100 138 -29083 172
rect -29135 121 -29083 138
rect -29053 172 -29001 173
rect -29053 138 -29046 172
rect -29046 138 -29012 172
rect -29012 138 -29001 172
rect -29053 121 -29001 138
rect -28971 172 -28919 173
rect -28971 138 -28958 172
rect -28958 138 -28924 172
rect -28924 138 -28919 172
rect -28971 121 -28919 138
rect -28889 172 -28837 173
rect -28889 138 -28870 172
rect -28870 138 -28837 172
rect -28889 121 -28837 138
rect -29135 99 -29083 109
rect -29135 65 -29134 99
rect -29134 65 -29100 99
rect -29100 65 -29083 99
rect -29135 57 -29083 65
rect -29053 99 -29001 109
rect -29053 65 -29046 99
rect -29046 65 -29012 99
rect -29012 65 -29001 99
rect -29053 57 -29001 65
rect -28971 99 -28919 109
rect -28971 65 -28958 99
rect -28958 65 -28924 99
rect -28924 65 -28919 99
rect -28971 57 -28919 65
rect -28889 99 -28837 109
rect -28889 65 -28870 99
rect -28870 65 -28837 99
rect -28889 57 -28837 65
rect -29135 26 -29083 45
rect -29135 -7 -29134 26
rect -29134 -7 -29100 26
rect -29100 -7 -29083 26
rect -29053 26 -29001 45
rect -29053 -7 -29046 26
rect -29046 -7 -29012 26
rect -29012 -7 -29001 26
rect -28971 26 -28919 45
rect -28971 -7 -28958 26
rect -28958 -7 -28924 26
rect -28924 -7 -28919 26
rect -28889 26 -28837 45
rect -28889 -7 -28870 26
rect -28870 -7 -28837 26
rect -29135 -47 -29083 -19
rect -29135 -71 -29134 -47
rect -29134 -71 -29100 -47
rect -29100 -71 -29083 -47
rect -29053 -47 -29001 -19
rect -29053 -71 -29046 -47
rect -29046 -71 -29012 -47
rect -29012 -71 -29001 -47
rect -28971 -47 -28919 -19
rect -28971 -71 -28958 -47
rect -28958 -71 -28924 -47
rect -28924 -71 -28919 -47
rect -28889 -47 -28837 -19
rect -28889 -71 -28870 -47
rect -28870 -71 -28837 -47
rect -29135 -120 -29083 -83
rect -29135 -135 -29134 -120
rect -29134 -135 -29100 -120
rect -29100 -135 -29083 -120
rect -29053 -120 -29001 -83
rect -29053 -135 -29046 -120
rect -29046 -135 -29012 -120
rect -29012 -135 -29001 -120
rect -28971 -120 -28919 -83
rect -28971 -135 -28958 -120
rect -28958 -135 -28924 -120
rect -28924 -135 -28919 -120
rect -28889 -120 -28837 -83
rect -28889 -135 -28870 -120
rect -28870 -135 -28837 -120
rect -29135 -154 -29134 -147
rect -29134 -154 -29100 -147
rect -29100 -154 -29083 -147
rect -29135 -193 -29083 -154
rect -29135 -199 -29134 -193
rect -29134 -199 -29100 -193
rect -29100 -199 -29083 -193
rect -29053 -154 -29046 -147
rect -29046 -154 -29012 -147
rect -29012 -154 -29001 -147
rect -29053 -193 -29001 -154
rect -29053 -199 -29046 -193
rect -29046 -199 -29012 -193
rect -29012 -199 -29001 -193
rect -28971 -154 -28958 -147
rect -28958 -154 -28924 -147
rect -28924 -154 -28919 -147
rect -28971 -193 -28919 -154
rect -28971 -199 -28958 -193
rect -28958 -199 -28924 -193
rect -28924 -199 -28919 -193
rect -28889 -154 -28870 -147
rect -28870 -154 -28837 -147
rect -28889 -193 -28837 -154
rect -28889 -199 -28870 -193
rect -28870 -199 -28837 -193
rect -29135 -227 -29134 -211
rect -29134 -227 -29100 -211
rect -29100 -227 -29083 -211
rect -29135 -263 -29083 -227
rect -29053 -227 -29046 -211
rect -29046 -227 -29012 -211
rect -29012 -227 -29001 -211
rect -29053 -263 -29001 -227
rect -28971 -227 -28958 -211
rect -28958 -227 -28924 -211
rect -28924 -227 -28919 -211
rect -28971 -263 -28919 -227
rect -28889 -227 -28870 -211
rect -28870 -227 -28837 -211
rect -28889 -263 -28837 -227
rect -29135 -300 -29134 -275
rect -29134 -300 -29100 -275
rect -29100 -300 -29083 -275
rect -29135 -327 -29083 -300
rect -29053 -300 -29046 -275
rect -29046 -300 -29012 -275
rect -29012 -300 -29001 -275
rect -29053 -327 -29001 -300
rect -28971 -300 -28958 -275
rect -28958 -300 -28924 -275
rect -28924 -300 -28919 -275
rect -28971 -327 -28919 -300
rect -28889 -300 -28870 -275
rect -28870 -300 -28837 -275
rect -28889 -327 -28837 -300
rect -29135 -373 -29134 -339
rect -29134 -373 -29100 -339
rect -29100 -373 -29083 -339
rect -29135 -391 -29083 -373
rect -29053 -373 -29046 -339
rect -29046 -373 -29012 -339
rect -29012 -373 -29001 -339
rect -29053 -391 -29001 -373
rect -28971 -373 -28958 -339
rect -28958 -373 -28924 -339
rect -28924 -373 -28919 -339
rect -28971 -391 -28919 -373
rect -28889 -373 -28870 -339
rect -28870 -373 -28837 -339
rect -28889 -391 -28837 -373
rect -29280 -8593 -29228 -8589
rect -31521 -8659 -31512 -8625
rect -31512 -8659 -31478 -8625
rect -31478 -8659 -31469 -8625
rect -31521 -8677 -31469 -8659
rect -31521 -8697 -31469 -8689
rect -31521 -8731 -31512 -8697
rect -31512 -8731 -31478 -8697
rect -31478 -8731 -31469 -8697
rect -29280 -8627 -29268 -8593
rect -29268 -8627 -29234 -8593
rect -29234 -8627 -29228 -8593
rect -29280 -8641 -29228 -8627
rect -29280 -8665 -29228 -8653
rect -29280 -8699 -29268 -8665
rect -29268 -8699 -29234 -8665
rect -29234 -8699 -29228 -8665
rect -29280 -8705 -29228 -8699
rect -31521 -8741 -31469 -8731
rect -21221 4644 -21169 4696
rect -21145 4644 -21093 4696
rect -21069 4644 -21017 4696
rect -20993 4644 -20941 4696
rect -20917 4644 -20865 4696
rect -20841 4644 -20789 4696
rect -21221 4518 -21169 4570
rect -21145 4518 -21093 4570
rect -21069 4518 -21017 4570
rect -20993 4518 -20941 4570
rect -20917 4518 -20865 4570
rect -20841 4518 -20789 4570
rect -28188 452 -28136 488
rect -28188 436 -28155 452
rect -28155 436 -28136 452
rect -28122 452 -28070 488
rect -28122 436 -28115 452
rect -28115 436 -28081 452
rect -28081 436 -28070 452
rect -28056 452 -28004 488
rect -28056 436 -28041 452
rect -28041 436 -28007 452
rect -28007 436 -28004 452
rect -27990 452 -27938 488
rect -27924 452 -27872 488
rect -27858 452 -27806 488
rect -27792 452 -27740 488
rect -27726 452 -27674 488
rect -27659 452 -27607 488
rect -27592 452 -27540 488
rect -27990 436 -27967 452
rect -27967 436 -27938 452
rect -27924 436 -27893 452
rect -27893 436 -27872 452
rect -27858 436 -27819 452
rect -27819 436 -27806 452
rect -27792 436 -27785 452
rect -27785 436 -27745 452
rect -27745 436 -27740 452
rect -27726 436 -27711 452
rect -27711 436 -27674 452
rect -27659 436 -27637 452
rect -27637 436 -27607 452
rect -27592 436 -27563 452
rect -27563 436 -27540 452
rect -27525 452 -27473 488
rect -27525 436 -27523 452
rect -27523 436 -27489 452
rect -27489 436 -27473 452
rect -27458 452 -27406 488
rect -27458 436 -27449 452
rect -27449 436 -27415 452
rect -27415 436 -27406 452
rect -27391 452 -27339 488
rect -27391 436 -27375 452
rect -27375 436 -27341 452
rect -27341 436 -27339 452
rect -27324 452 -27272 488
rect -27257 452 -27205 488
rect -27190 452 -27138 488
rect -27324 436 -27301 452
rect -27301 436 -27272 452
rect -27257 436 -27227 452
rect -27227 436 -27205 452
rect -27190 436 -27153 452
rect -27153 436 -27138 452
rect -28188 418 -28155 420
rect -28155 418 -28136 420
rect -28188 380 -28136 418
rect -28188 368 -28155 380
rect -28155 368 -28136 380
rect -28122 418 -28115 420
rect -28115 418 -28081 420
rect -28081 418 -28070 420
rect -28122 380 -28070 418
rect -28122 368 -28115 380
rect -28115 368 -28081 380
rect -28081 368 -28070 380
rect -28056 418 -28041 420
rect -28041 418 -28007 420
rect -28007 418 -28004 420
rect -28056 380 -28004 418
rect -28056 368 -28041 380
rect -28041 368 -28007 380
rect -28007 368 -28004 380
rect -27990 418 -27967 420
rect -27967 418 -27938 420
rect -27924 418 -27893 420
rect -27893 418 -27872 420
rect -27858 418 -27819 420
rect -27819 418 -27806 420
rect -27792 418 -27785 420
rect -27785 418 -27745 420
rect -27745 418 -27740 420
rect -27726 418 -27711 420
rect -27711 418 -27674 420
rect -27659 418 -27637 420
rect -27637 418 -27607 420
rect -27592 418 -27563 420
rect -27563 418 -27540 420
rect -27990 380 -27938 418
rect -27924 380 -27872 418
rect -27858 380 -27806 418
rect -27792 380 -27740 418
rect -27726 380 -27674 418
rect -27659 380 -27607 418
rect -27592 380 -27540 418
rect -27990 368 -27967 380
rect -27967 368 -27938 380
rect -27924 368 -27893 380
rect -27893 368 -27872 380
rect -27858 368 -27819 380
rect -27819 368 -27806 380
rect -27792 368 -27785 380
rect -27785 368 -27745 380
rect -27745 368 -27740 380
rect -27726 368 -27711 380
rect -27711 368 -27674 380
rect -27659 368 -27637 380
rect -27637 368 -27607 380
rect -27592 368 -27563 380
rect -27563 368 -27540 380
rect -27525 418 -27523 420
rect -27523 418 -27489 420
rect -27489 418 -27473 420
rect -27525 380 -27473 418
rect -27525 368 -27523 380
rect -27523 368 -27489 380
rect -27489 368 -27473 380
rect -27458 418 -27449 420
rect -27449 418 -27415 420
rect -27415 418 -27406 420
rect -27458 380 -27406 418
rect -27458 368 -27449 380
rect -27449 368 -27415 380
rect -27415 368 -27406 380
rect -27391 418 -27375 420
rect -27375 418 -27341 420
rect -27341 418 -27339 420
rect -27391 380 -27339 418
rect -27391 368 -27375 380
rect -27375 368 -27341 380
rect -27341 368 -27339 380
rect -27324 418 -27301 420
rect -27301 418 -27272 420
rect -27257 418 -27227 420
rect -27227 418 -27205 420
rect -27190 418 -27153 420
rect -27153 418 -27138 420
rect -27324 380 -27272 418
rect -27257 380 -27205 418
rect -27190 380 -27138 418
rect -27324 368 -27301 380
rect -27301 368 -27272 380
rect -27257 368 -27227 380
rect -27227 368 -27205 380
rect -27190 368 -27153 380
rect -27153 368 -27138 380
rect -28188 346 -28155 352
rect -28155 346 -28136 352
rect -28188 308 -28136 346
rect -28188 300 -28155 308
rect -28155 300 -28136 308
rect -28122 346 -28115 352
rect -28115 346 -28081 352
rect -28081 346 -28070 352
rect -28122 308 -28070 346
rect -28122 300 -28115 308
rect -28115 300 -28081 308
rect -28081 300 -28070 308
rect -28056 346 -28041 352
rect -28041 346 -28007 352
rect -28007 346 -28004 352
rect -28056 308 -28004 346
rect -28056 300 -28041 308
rect -28041 300 -28007 308
rect -28007 300 -28004 308
rect -27990 346 -27967 352
rect -27967 346 -27938 352
rect -27924 346 -27893 352
rect -27893 346 -27872 352
rect -27858 346 -27819 352
rect -27819 346 -27806 352
rect -27792 346 -27785 352
rect -27785 346 -27745 352
rect -27745 346 -27740 352
rect -27726 346 -27711 352
rect -27711 346 -27674 352
rect -27659 346 -27637 352
rect -27637 346 -27607 352
rect -27592 346 -27563 352
rect -27563 346 -27540 352
rect -27990 308 -27938 346
rect -27924 308 -27872 346
rect -27858 308 -27806 346
rect -27792 308 -27740 346
rect -27726 308 -27674 346
rect -27659 308 -27607 346
rect -27592 308 -27540 346
rect -27990 300 -27967 308
rect -27967 300 -27938 308
rect -27924 300 -27893 308
rect -27893 300 -27872 308
rect -27858 300 -27819 308
rect -27819 300 -27806 308
rect -27792 300 -27785 308
rect -27785 300 -27745 308
rect -27745 300 -27740 308
rect -27726 300 -27711 308
rect -27711 300 -27674 308
rect -27659 300 -27637 308
rect -27637 300 -27607 308
rect -27592 300 -27563 308
rect -27563 300 -27540 308
rect -27525 346 -27523 352
rect -27523 346 -27489 352
rect -27489 346 -27473 352
rect -27525 308 -27473 346
rect -27525 300 -27523 308
rect -27523 300 -27489 308
rect -27489 300 -27473 308
rect -27458 346 -27449 352
rect -27449 346 -27415 352
rect -27415 346 -27406 352
rect -27458 308 -27406 346
rect -27458 300 -27449 308
rect -27449 300 -27415 308
rect -27415 300 -27406 308
rect -27391 346 -27375 352
rect -27375 346 -27341 352
rect -27341 346 -27339 352
rect -27391 308 -27339 346
rect -27391 300 -27375 308
rect -27375 300 -27341 308
rect -27341 300 -27339 308
rect -27324 346 -27301 352
rect -27301 346 -27272 352
rect -27257 346 -27227 352
rect -27227 346 -27205 352
rect -27190 346 -27153 352
rect -27153 346 -27138 352
rect -27324 308 -27272 346
rect -27257 308 -27205 346
rect -27190 308 -27138 346
rect -27324 300 -27301 308
rect -27301 300 -27272 308
rect -27257 300 -27227 308
rect -27227 300 -27205 308
rect -27190 300 -27153 308
rect -27153 300 -27138 308
rect -28188 274 -28155 284
rect -28155 274 -28136 284
rect -28188 236 -28136 274
rect -28188 232 -28155 236
rect -28155 232 -28136 236
rect -28122 274 -28115 284
rect -28115 274 -28081 284
rect -28081 274 -28070 284
rect -28122 236 -28070 274
rect -28122 232 -28115 236
rect -28115 232 -28081 236
rect -28081 232 -28070 236
rect -28056 274 -28041 284
rect -28041 274 -28007 284
rect -28007 274 -28004 284
rect -28056 236 -28004 274
rect -28056 232 -28041 236
rect -28041 232 -28007 236
rect -28007 232 -28004 236
rect -27990 274 -27967 284
rect -27967 274 -27938 284
rect -27924 274 -27893 284
rect -27893 274 -27872 284
rect -27858 274 -27819 284
rect -27819 274 -27806 284
rect -27792 274 -27785 284
rect -27785 274 -27745 284
rect -27745 274 -27740 284
rect -27726 274 -27711 284
rect -27711 274 -27674 284
rect -27659 274 -27637 284
rect -27637 274 -27607 284
rect -27592 274 -27563 284
rect -27563 274 -27540 284
rect -27990 236 -27938 274
rect -27924 236 -27872 274
rect -27858 236 -27806 274
rect -27792 236 -27740 274
rect -27726 236 -27674 274
rect -27659 236 -27607 274
rect -27592 236 -27540 274
rect -27990 232 -27967 236
rect -27967 232 -27938 236
rect -27924 232 -27893 236
rect -27893 232 -27872 236
rect -27858 232 -27819 236
rect -27819 232 -27806 236
rect -27792 232 -27785 236
rect -27785 232 -27745 236
rect -27745 232 -27740 236
rect -27726 232 -27711 236
rect -27711 232 -27674 236
rect -27659 232 -27637 236
rect -27637 232 -27607 236
rect -27592 232 -27563 236
rect -27563 232 -27540 236
rect -27525 274 -27523 284
rect -27523 274 -27489 284
rect -27489 274 -27473 284
rect -27525 236 -27473 274
rect -27525 232 -27523 236
rect -27523 232 -27489 236
rect -27489 232 -27473 236
rect -27458 274 -27449 284
rect -27449 274 -27415 284
rect -27415 274 -27406 284
rect -27458 236 -27406 274
rect -27458 232 -27449 236
rect -27449 232 -27415 236
rect -27415 232 -27406 236
rect -27391 274 -27375 284
rect -27375 274 -27341 284
rect -27341 274 -27339 284
rect -27391 236 -27339 274
rect -27391 232 -27375 236
rect -27375 232 -27341 236
rect -27341 232 -27339 236
rect -27324 274 -27301 284
rect -27301 274 -27272 284
rect -27257 274 -27227 284
rect -27227 274 -27205 284
rect -27190 274 -27153 284
rect -27153 274 -27138 284
rect -27324 236 -27272 274
rect -27257 236 -27205 274
rect -27190 236 -27138 274
rect -27324 232 -27301 236
rect -27301 232 -27272 236
rect -27257 232 -27227 236
rect -27227 232 -27205 236
rect -27190 232 -27153 236
rect -27153 232 -27138 236
rect -28188 202 -28155 216
rect -28155 202 -28136 216
rect -28188 164 -28136 202
rect -28122 202 -28115 216
rect -28115 202 -28081 216
rect -28081 202 -28070 216
rect -28122 164 -28070 202
rect -28056 202 -28041 216
rect -28041 202 -28007 216
rect -28007 202 -28004 216
rect -28056 164 -28004 202
rect -27990 202 -27967 216
rect -27967 202 -27938 216
rect -27924 202 -27893 216
rect -27893 202 -27872 216
rect -27858 202 -27819 216
rect -27819 202 -27806 216
rect -27792 202 -27785 216
rect -27785 202 -27745 216
rect -27745 202 -27740 216
rect -27726 202 -27711 216
rect -27711 202 -27674 216
rect -27659 202 -27637 216
rect -27637 202 -27607 216
rect -27592 202 -27563 216
rect -27563 202 -27540 216
rect -27990 164 -27938 202
rect -27924 164 -27872 202
rect -27858 164 -27806 202
rect -27792 164 -27740 202
rect -27726 164 -27674 202
rect -27659 164 -27607 202
rect -27592 164 -27540 202
rect -27525 202 -27523 216
rect -27523 202 -27489 216
rect -27489 202 -27473 216
rect -27525 164 -27473 202
rect -27458 202 -27449 216
rect -27449 202 -27415 216
rect -27415 202 -27406 216
rect -27458 164 -27406 202
rect -27391 202 -27375 216
rect -27375 202 -27341 216
rect -27341 202 -27339 216
rect -27391 164 -27339 202
rect -27324 202 -27301 216
rect -27301 202 -27272 216
rect -27257 202 -27227 216
rect -27227 202 -27205 216
rect -27190 202 -27153 216
rect -27153 202 -27138 216
rect -27324 164 -27272 202
rect -27257 164 -27205 202
rect -27190 164 -27138 202
rect -28188 130 -28155 148
rect -28155 130 -28136 148
rect -28188 96 -28136 130
rect -28122 130 -28115 148
rect -28115 130 -28081 148
rect -28081 130 -28070 148
rect -28122 96 -28070 130
rect -28056 130 -28041 148
rect -28041 130 -28007 148
rect -28007 130 -28004 148
rect -28056 96 -28004 130
rect -27990 130 -27967 148
rect -27967 130 -27938 148
rect -27924 130 -27893 148
rect -27893 130 -27872 148
rect -27858 130 -27819 148
rect -27819 130 -27806 148
rect -27792 130 -27785 148
rect -27785 130 -27745 148
rect -27745 130 -27740 148
rect -27726 130 -27711 148
rect -27711 130 -27674 148
rect -27659 130 -27637 148
rect -27637 130 -27607 148
rect -27592 130 -27563 148
rect -27563 130 -27540 148
rect -27990 96 -27938 130
rect -27924 96 -27872 130
rect -27858 96 -27806 130
rect -27792 96 -27740 130
rect -27726 96 -27674 130
rect -27659 96 -27607 130
rect -27592 96 -27540 130
rect -27525 130 -27523 148
rect -27523 130 -27489 148
rect -27489 130 -27473 148
rect -27525 96 -27473 130
rect -27458 130 -27449 148
rect -27449 130 -27415 148
rect -27415 130 -27406 148
rect -27458 96 -27406 130
rect -27391 130 -27375 148
rect -27375 130 -27341 148
rect -27341 130 -27339 148
rect -27391 96 -27339 130
rect -27324 130 -27301 148
rect -27301 130 -27272 148
rect -27257 130 -27227 148
rect -27227 130 -27205 148
rect -27190 130 -27153 148
rect -27153 130 -27138 148
rect -27324 96 -27272 130
rect -27257 96 -27205 130
rect -27190 96 -27138 130
rect -28188 58 -28155 80
rect -28155 58 -28136 80
rect -28188 28 -28136 58
rect -28122 58 -28115 80
rect -28115 58 -28081 80
rect -28081 58 -28070 80
rect -28122 28 -28070 58
rect -28056 58 -28041 80
rect -28041 58 -28007 80
rect -28007 58 -28004 80
rect -28056 28 -28004 58
rect -27990 58 -27967 80
rect -27967 58 -27938 80
rect -27924 58 -27893 80
rect -27893 58 -27872 80
rect -27858 58 -27819 80
rect -27819 58 -27806 80
rect -27792 58 -27785 80
rect -27785 58 -27745 80
rect -27745 58 -27740 80
rect -27726 58 -27711 80
rect -27711 58 -27674 80
rect -27659 58 -27637 80
rect -27637 58 -27607 80
rect -27592 58 -27563 80
rect -27563 58 -27540 80
rect -27990 28 -27938 58
rect -27924 28 -27872 58
rect -27858 28 -27806 58
rect -27792 28 -27740 58
rect -27726 28 -27674 58
rect -27659 28 -27607 58
rect -27592 28 -27540 58
rect -27525 58 -27523 80
rect -27523 58 -27489 80
rect -27489 58 -27473 80
rect -27525 28 -27473 58
rect -27458 58 -27449 80
rect -27449 58 -27415 80
rect -27415 58 -27406 80
rect -27458 28 -27406 58
rect -27391 58 -27375 80
rect -27375 58 -27341 80
rect -27341 58 -27339 80
rect -27391 28 -27339 58
rect -27324 58 -27301 80
rect -27301 58 -27272 80
rect -27257 58 -27227 80
rect -27227 58 -27205 80
rect -27190 58 -27153 80
rect -27153 58 -27138 80
rect -27324 28 -27272 58
rect -27257 28 -27205 58
rect -27190 28 -27138 58
rect -28188 -14 -28155 12
rect -28155 -14 -28136 12
rect -28188 -40 -28136 -14
rect -28122 -14 -28115 12
rect -28115 -14 -28081 12
rect -28081 -14 -28070 12
rect -28122 -40 -28070 -14
rect -28056 -14 -28041 12
rect -28041 -14 -28007 12
rect -28007 -14 -28004 12
rect -28056 -40 -28004 -14
rect -27990 -14 -27967 12
rect -27967 -14 -27938 12
rect -27924 -14 -27893 12
rect -27893 -14 -27872 12
rect -27858 -14 -27819 12
rect -27819 -14 -27806 12
rect -27792 -14 -27785 12
rect -27785 -14 -27745 12
rect -27745 -14 -27740 12
rect -27726 -14 -27711 12
rect -27711 -14 -27674 12
rect -27659 -14 -27637 12
rect -27637 -14 -27607 12
rect -27592 -14 -27563 12
rect -27563 -14 -27540 12
rect -27990 -40 -27938 -14
rect -27924 -40 -27872 -14
rect -27858 -40 -27806 -14
rect -27792 -40 -27740 -14
rect -27726 -40 -27674 -14
rect -27659 -40 -27607 -14
rect -27592 -40 -27540 -14
rect -27525 -14 -27523 12
rect -27523 -14 -27489 12
rect -27489 -14 -27473 12
rect -27525 -40 -27473 -14
rect -27458 -14 -27449 12
rect -27449 -14 -27415 12
rect -27415 -14 -27406 12
rect -27458 -40 -27406 -14
rect -27391 -14 -27375 12
rect -27375 -14 -27341 12
rect -27341 -14 -27339 12
rect -27391 -40 -27339 -14
rect -27324 -14 -27301 12
rect -27301 -14 -27272 12
rect -27257 -14 -27227 12
rect -27227 -14 -27205 12
rect -27190 -14 -27153 12
rect -27153 -14 -27138 12
rect -27324 -40 -27272 -14
rect -27257 -40 -27205 -14
rect -27190 -40 -27138 -14
rect -28188 -86 -28155 -56
rect -28155 -86 -28136 -56
rect -28188 -108 -28136 -86
rect -28122 -86 -28115 -56
rect -28115 -86 -28081 -56
rect -28081 -86 -28070 -56
rect -28122 -108 -28070 -86
rect -28056 -86 -28041 -56
rect -28041 -86 -28007 -56
rect -28007 -86 -28004 -56
rect -28056 -108 -28004 -86
rect -27990 -86 -27967 -56
rect -27967 -86 -27938 -56
rect -27924 -86 -27893 -56
rect -27893 -86 -27872 -56
rect -27858 -86 -27819 -56
rect -27819 -86 -27806 -56
rect -27792 -86 -27785 -56
rect -27785 -86 -27745 -56
rect -27745 -86 -27740 -56
rect -27726 -86 -27711 -56
rect -27711 -86 -27674 -56
rect -27659 -86 -27637 -56
rect -27637 -86 -27607 -56
rect -27592 -86 -27563 -56
rect -27563 -86 -27540 -56
rect -27990 -108 -27938 -86
rect -27924 -108 -27872 -86
rect -27858 -108 -27806 -86
rect -27792 -108 -27740 -86
rect -27726 -108 -27674 -86
rect -27659 -108 -27607 -86
rect -27592 -108 -27540 -86
rect -27525 -86 -27523 -56
rect -27523 -86 -27489 -56
rect -27489 -86 -27473 -56
rect -27525 -108 -27473 -86
rect -27458 -86 -27449 -56
rect -27449 -86 -27415 -56
rect -27415 -86 -27406 -56
rect -27458 -108 -27406 -86
rect -27391 -86 -27375 -56
rect -27375 -86 -27341 -56
rect -27341 -86 -27339 -56
rect -27391 -108 -27339 -86
rect -27324 -86 -27301 -56
rect -27301 -86 -27272 -56
rect -27257 -86 -27227 -56
rect -27227 -86 -27205 -56
rect -27190 -86 -27153 -56
rect -27153 -86 -27138 -56
rect -27324 -108 -27272 -86
rect -27257 -108 -27205 -86
rect -27190 -108 -27138 -86
rect -28188 -158 -28155 -124
rect -28155 -158 -28136 -124
rect -28188 -176 -28136 -158
rect -28122 -158 -28115 -124
rect -28115 -158 -28081 -124
rect -28081 -158 -28070 -124
rect -28122 -176 -28070 -158
rect -28056 -158 -28041 -124
rect -28041 -158 -28007 -124
rect -28007 -158 -28004 -124
rect -28056 -176 -28004 -158
rect -27990 -158 -27967 -124
rect -27967 -158 -27938 -124
rect -27924 -158 -27893 -124
rect -27893 -158 -27872 -124
rect -27858 -158 -27819 -124
rect -27819 -158 -27806 -124
rect -27792 -158 -27785 -124
rect -27785 -158 -27745 -124
rect -27745 -158 -27740 -124
rect -27726 -158 -27711 -124
rect -27711 -158 -27674 -124
rect -27659 -158 -27637 -124
rect -27637 -158 -27607 -124
rect -27592 -158 -27563 -124
rect -27563 -158 -27540 -124
rect -27990 -176 -27938 -158
rect -27924 -176 -27872 -158
rect -27858 -176 -27806 -158
rect -27792 -176 -27740 -158
rect -27726 -176 -27674 -158
rect -27659 -176 -27607 -158
rect -27592 -176 -27540 -158
rect -27525 -158 -27523 -124
rect -27523 -158 -27489 -124
rect -27489 -158 -27473 -124
rect -27525 -176 -27473 -158
rect -27458 -158 -27449 -124
rect -27449 -158 -27415 -124
rect -27415 -158 -27406 -124
rect -27458 -176 -27406 -158
rect -27391 -158 -27375 -124
rect -27375 -158 -27341 -124
rect -27341 -158 -27339 -124
rect -27391 -176 -27339 -158
rect -27324 -158 -27301 -124
rect -27301 -158 -27272 -124
rect -27257 -158 -27227 -124
rect -27227 -158 -27205 -124
rect -27190 -158 -27153 -124
rect -27153 -158 -27138 -124
rect -27324 -176 -27272 -158
rect -27257 -176 -27205 -158
rect -27190 -176 -27138 -158
rect -28188 -196 -28136 -192
rect -28188 -230 -28155 -196
rect -28155 -230 -28136 -196
rect -28188 -244 -28136 -230
rect -28122 -196 -28070 -192
rect -28122 -230 -28115 -196
rect -28115 -230 -28081 -196
rect -28081 -230 -28070 -196
rect -28122 -244 -28070 -230
rect -28056 -196 -28004 -192
rect -28056 -230 -28041 -196
rect -28041 -230 -28007 -196
rect -28007 -230 -28004 -196
rect -28056 -244 -28004 -230
rect -27990 -196 -27938 -192
rect -27924 -196 -27872 -192
rect -27858 -196 -27806 -192
rect -27792 -196 -27740 -192
rect -27726 -196 -27674 -192
rect -27659 -196 -27607 -192
rect -27592 -196 -27540 -192
rect -27990 -230 -27967 -196
rect -27967 -230 -27938 -196
rect -27924 -230 -27893 -196
rect -27893 -230 -27872 -196
rect -27858 -230 -27819 -196
rect -27819 -230 -27806 -196
rect -27792 -230 -27785 -196
rect -27785 -230 -27745 -196
rect -27745 -230 -27740 -196
rect -27726 -230 -27711 -196
rect -27711 -230 -27674 -196
rect -27659 -230 -27637 -196
rect -27637 -230 -27607 -196
rect -27592 -230 -27563 -196
rect -27563 -230 -27540 -196
rect -27990 -244 -27938 -230
rect -27924 -244 -27872 -230
rect -27858 -244 -27806 -230
rect -27792 -244 -27740 -230
rect -27726 -244 -27674 -230
rect -27659 -244 -27607 -230
rect -27592 -244 -27540 -230
rect -27525 -196 -27473 -192
rect -27525 -230 -27523 -196
rect -27523 -230 -27489 -196
rect -27489 -230 -27473 -196
rect -27525 -244 -27473 -230
rect -27458 -196 -27406 -192
rect -27458 -230 -27449 -196
rect -27449 -230 -27415 -196
rect -27415 -230 -27406 -196
rect -27458 -244 -27406 -230
rect -27391 -196 -27339 -192
rect -27391 -230 -27375 -196
rect -27375 -230 -27341 -196
rect -27341 -230 -27339 -196
rect -27391 -244 -27339 -230
rect -27324 -196 -27272 -192
rect -27257 -196 -27205 -192
rect -27190 -196 -27138 -192
rect -27324 -230 -27301 -196
rect -27301 -230 -27272 -196
rect -27257 -230 -27227 -196
rect -27227 -230 -27205 -196
rect -27190 -230 -27153 -196
rect -27153 -230 -27138 -196
rect -27324 -244 -27272 -230
rect -27257 -244 -27205 -230
rect -27190 -244 -27138 -230
rect -28188 -268 -28136 -260
rect -28188 -302 -28155 -268
rect -28155 -302 -28136 -268
rect -28188 -312 -28136 -302
rect -28122 -268 -28070 -260
rect -28122 -302 -28115 -268
rect -28115 -302 -28081 -268
rect -28081 -302 -28070 -268
rect -28122 -312 -28070 -302
rect -28056 -268 -28004 -260
rect -28056 -302 -28041 -268
rect -28041 -302 -28007 -268
rect -28007 -302 -28004 -268
rect -28056 -312 -28004 -302
rect -27990 -268 -27938 -260
rect -27924 -268 -27872 -260
rect -27858 -268 -27806 -260
rect -27792 -268 -27740 -260
rect -27726 -268 -27674 -260
rect -27659 -268 -27607 -260
rect -27592 -268 -27540 -260
rect -27990 -302 -27967 -268
rect -27967 -302 -27938 -268
rect -27924 -302 -27893 -268
rect -27893 -302 -27872 -268
rect -27858 -302 -27819 -268
rect -27819 -302 -27806 -268
rect -27792 -302 -27785 -268
rect -27785 -302 -27745 -268
rect -27745 -302 -27740 -268
rect -27726 -302 -27711 -268
rect -27711 -302 -27674 -268
rect -27659 -302 -27637 -268
rect -27637 -302 -27607 -268
rect -27592 -302 -27563 -268
rect -27563 -302 -27540 -268
rect -27990 -312 -27938 -302
rect -27924 -312 -27872 -302
rect -27858 -312 -27806 -302
rect -27792 -312 -27740 -302
rect -27726 -312 -27674 -302
rect -27659 -312 -27607 -302
rect -27592 -312 -27540 -302
rect -27525 -268 -27473 -260
rect -27525 -302 -27523 -268
rect -27523 -302 -27489 -268
rect -27489 -302 -27473 -268
rect -27525 -312 -27473 -302
rect -27458 -268 -27406 -260
rect -27458 -302 -27449 -268
rect -27449 -302 -27415 -268
rect -27415 -302 -27406 -268
rect -27458 -312 -27406 -302
rect -27391 -268 -27339 -260
rect -27391 -302 -27375 -268
rect -27375 -302 -27341 -268
rect -27341 -302 -27339 -268
rect -27391 -312 -27339 -302
rect -27324 -268 -27272 -260
rect -27257 -268 -27205 -260
rect -27190 -268 -27138 -260
rect -27324 -302 -27301 -268
rect -27301 -302 -27272 -268
rect -27257 -302 -27227 -268
rect -27227 -302 -27205 -268
rect -27190 -302 -27153 -268
rect -27153 -302 -27138 -268
rect -27324 -312 -27272 -302
rect -27257 -312 -27205 -302
rect -27190 -312 -27138 -302
rect -28188 -340 -28136 -328
rect -28188 -374 -28155 -340
rect -28155 -374 -28136 -340
rect -28188 -380 -28136 -374
rect -28122 -340 -28070 -328
rect -28122 -374 -28115 -340
rect -28115 -374 -28081 -340
rect -28081 -374 -28070 -340
rect -28122 -380 -28070 -374
rect -28056 -340 -28004 -328
rect -28056 -374 -28041 -340
rect -28041 -374 -28007 -340
rect -28007 -374 -28004 -340
rect -28056 -380 -28004 -374
rect -27990 -340 -27938 -328
rect -27924 -340 -27872 -328
rect -27858 -340 -27806 -328
rect -27792 -340 -27740 -328
rect -27726 -340 -27674 -328
rect -27659 -340 -27607 -328
rect -27592 -340 -27540 -328
rect -27990 -374 -27967 -340
rect -27967 -374 -27938 -340
rect -27924 -374 -27893 -340
rect -27893 -374 -27872 -340
rect -27858 -374 -27819 -340
rect -27819 -374 -27806 -340
rect -27792 -374 -27785 -340
rect -27785 -374 -27745 -340
rect -27745 -374 -27740 -340
rect -27726 -374 -27711 -340
rect -27711 -374 -27674 -340
rect -27659 -374 -27637 -340
rect -27637 -374 -27607 -340
rect -27592 -374 -27563 -340
rect -27563 -374 -27540 -340
rect -27990 -380 -27938 -374
rect -27924 -380 -27872 -374
rect -27858 -380 -27806 -374
rect -27792 -380 -27740 -374
rect -27726 -380 -27674 -374
rect -27659 -380 -27607 -374
rect -27592 -380 -27540 -374
rect -27525 -340 -27473 -328
rect -27525 -374 -27523 -340
rect -27523 -374 -27489 -340
rect -27489 -374 -27473 -340
rect -27525 -380 -27473 -374
rect -27458 -340 -27406 -328
rect -27458 -374 -27449 -340
rect -27449 -374 -27415 -340
rect -27415 -374 -27406 -340
rect -27458 -380 -27406 -374
rect -27391 -340 -27339 -328
rect -27391 -374 -27375 -340
rect -27375 -374 -27341 -340
rect -27341 -374 -27339 -340
rect -27391 -380 -27339 -374
rect -27324 -340 -27272 -328
rect -27257 -340 -27205 -328
rect -27190 -340 -27138 -328
rect -27324 -374 -27301 -340
rect -27301 -374 -27272 -340
rect -27257 -374 -27227 -340
rect -27227 -374 -27205 -340
rect -27190 -374 -27153 -340
rect -27153 -374 -27138 -340
rect -27324 -380 -27272 -374
rect -27257 -380 -27205 -374
rect -27190 -380 -27138 -374
rect -787 3688 -735 3700
rect -717 3688 -665 3700
rect -646 3688 -594 3700
rect -575 3688 -523 3700
rect -504 3688 -452 3700
rect -787 3654 -757 3688
rect -757 3654 -735 3688
rect -717 3654 -677 3688
rect -677 3654 -665 3688
rect -646 3654 -643 3688
rect -643 3654 -597 3688
rect -597 3654 -594 3688
rect -575 3654 -563 3688
rect -563 3654 -523 3688
rect -504 3654 -482 3688
rect -482 3654 -452 3688
rect -787 3648 -735 3654
rect -717 3648 -665 3654
rect -646 3648 -594 3654
rect -575 3648 -523 3654
rect -504 3648 -452 3654
rect 170 3688 222 3697
rect 170 3654 171 3688
rect 171 3654 205 3688
rect 205 3654 222 3688
rect 170 3645 222 3654
rect 235 3688 287 3697
rect 235 3654 244 3688
rect 244 3654 278 3688
rect 278 3654 287 3688
rect 235 3645 287 3654
rect 300 3688 352 3697
rect 300 3654 317 3688
rect 317 3654 351 3688
rect 351 3654 352 3688
rect 300 3645 352 3654
rect 365 3688 417 3697
rect 430 3688 482 3697
rect 495 3688 547 3697
rect 560 3688 612 3697
rect 625 3688 677 3697
rect 690 3688 742 3697
rect 365 3654 390 3688
rect 390 3654 417 3688
rect 430 3654 463 3688
rect 463 3654 482 3688
rect 495 3654 497 3688
rect 497 3654 536 3688
rect 536 3654 547 3688
rect 560 3654 570 3688
rect 570 3654 609 3688
rect 609 3654 612 3688
rect 625 3654 643 3688
rect 643 3654 677 3688
rect 690 3654 716 3688
rect 716 3654 742 3688
rect 365 3645 417 3654
rect 430 3645 482 3654
rect 495 3645 547 3654
rect 560 3645 612 3654
rect 625 3645 677 3654
rect 690 3645 742 3654
rect 755 3688 807 3697
rect 755 3654 789 3688
rect 789 3654 807 3688
rect 755 3645 807 3654
rect 820 3688 872 3697
rect 820 3654 828 3688
rect 828 3654 862 3688
rect 862 3654 872 3688
rect 820 3645 872 3654
rect 885 3688 937 3697
rect 885 3654 901 3688
rect 901 3654 935 3688
rect 935 3654 937 3688
rect 885 3645 937 3654
rect 950 3688 1002 3697
rect 1015 3688 1067 3697
rect 1080 3688 1132 3697
rect 1145 3688 1197 3697
rect 1210 3688 1262 3697
rect 1275 3688 1327 3697
rect 1340 3688 1392 3697
rect 950 3654 974 3688
rect 974 3654 1002 3688
rect 1015 3654 1047 3688
rect 1047 3654 1067 3688
rect 1080 3654 1081 3688
rect 1081 3654 1120 3688
rect 1120 3654 1132 3688
rect 1145 3654 1154 3688
rect 1154 3654 1193 3688
rect 1193 3654 1197 3688
rect 1210 3654 1227 3688
rect 1227 3654 1262 3688
rect 1275 3654 1300 3688
rect 1300 3654 1327 3688
rect 1340 3654 1373 3688
rect 1373 3654 1392 3688
rect 950 3645 1002 3654
rect 1015 3645 1067 3654
rect 1080 3645 1132 3654
rect 1145 3645 1197 3654
rect 1210 3645 1262 3654
rect 1275 3645 1327 3654
rect 1340 3645 1392 3654
rect 1405 3688 1457 3697
rect 1405 3654 1412 3688
rect 1412 3654 1446 3688
rect 1446 3654 1457 3688
rect 1405 3645 1457 3654
rect 1470 3688 1522 3697
rect 1470 3654 1485 3688
rect 1485 3654 1519 3688
rect 1519 3654 1522 3688
rect 1470 3645 1522 3654
rect 1535 3688 1587 3697
rect 1600 3688 1652 3697
rect 1665 3688 1717 3697
rect 1730 3688 1782 3697
rect 1795 3688 1847 3697
rect 1860 3688 1912 3697
rect 1925 3688 1977 3697
rect 1535 3654 1558 3688
rect 1558 3654 1587 3688
rect 1600 3654 1631 3688
rect 1631 3654 1652 3688
rect 1665 3654 1704 3688
rect 1704 3654 1717 3688
rect 1730 3654 1738 3688
rect 1738 3654 1777 3688
rect 1777 3654 1782 3688
rect 1795 3654 1811 3688
rect 1811 3654 1847 3688
rect 1860 3654 1884 3688
rect 1884 3654 1912 3688
rect 1925 3654 1957 3688
rect 1957 3654 1977 3688
rect 1535 3645 1587 3654
rect 1600 3645 1652 3654
rect 1665 3645 1717 3654
rect 1730 3645 1782 3654
rect 1795 3645 1847 3654
rect 1860 3645 1912 3654
rect 1925 3645 1977 3654
rect 1990 3688 2042 3697
rect 1990 3654 1995 3688
rect 1995 3654 2029 3688
rect 2029 3654 2042 3688
rect 1990 3645 2042 3654
rect 2055 3688 2107 3697
rect 2055 3654 2067 3688
rect 2067 3654 2101 3688
rect 2101 3654 2107 3688
rect 2055 3645 2107 3654
rect 2120 3688 2172 3697
rect 2185 3688 2237 3697
rect 2250 3688 2302 3697
rect 2315 3688 2367 3697
rect 2380 3688 2432 3697
rect 2445 3688 2497 3697
rect 2510 3688 2562 3697
rect 2575 3688 2627 3697
rect 2120 3654 2139 3688
rect 2139 3654 2172 3688
rect 2185 3654 2211 3688
rect 2211 3654 2237 3688
rect 2250 3654 2283 3688
rect 2283 3654 2302 3688
rect 2315 3654 2317 3688
rect 2317 3654 2355 3688
rect 2355 3654 2367 3688
rect 2380 3654 2389 3688
rect 2389 3654 2427 3688
rect 2427 3654 2432 3688
rect 2445 3654 2461 3688
rect 2461 3654 2497 3688
rect 2510 3654 2533 3688
rect 2533 3654 2562 3688
rect 2575 3654 2605 3688
rect 2605 3654 2627 3688
rect 2120 3645 2172 3654
rect 2185 3645 2237 3654
rect 2250 3645 2302 3654
rect 2315 3645 2367 3654
rect 2380 3645 2432 3654
rect 2445 3645 2497 3654
rect 2510 3645 2562 3654
rect 2575 3645 2627 3654
rect 2640 3688 2692 3697
rect 2640 3654 2643 3688
rect 2643 3654 2677 3688
rect 2677 3654 2692 3688
rect 2640 3645 2692 3654
rect 2705 3688 2757 3697
rect 2705 3654 2715 3688
rect 2715 3654 2749 3688
rect 2749 3654 2757 3688
rect 2705 3645 2757 3654
rect 2770 3688 2822 3697
rect 2770 3654 2787 3688
rect 2787 3654 2821 3688
rect 2821 3654 2822 3688
rect 2770 3645 2822 3654
rect 2835 3688 2887 3697
rect 2900 3688 2952 3697
rect 2965 3688 3017 3697
rect 3030 3688 3082 3697
rect 3095 3688 3147 3697
rect 3160 3688 3212 3697
rect 3224 3688 3276 3697
rect 2835 3654 2859 3688
rect 2859 3654 2887 3688
rect 2900 3654 2931 3688
rect 2931 3654 2952 3688
rect 2965 3654 3003 3688
rect 3003 3654 3017 3688
rect 3030 3654 3037 3688
rect 3037 3654 3075 3688
rect 3075 3654 3082 3688
rect 3095 3654 3109 3688
rect 3109 3654 3147 3688
rect 3160 3654 3181 3688
rect 3181 3654 3212 3688
rect 3224 3654 3253 3688
rect 3253 3654 3276 3688
rect 2835 3645 2887 3654
rect 2900 3645 2952 3654
rect 2965 3645 3017 3654
rect 3030 3645 3082 3654
rect 3095 3645 3147 3654
rect 3160 3645 3212 3654
rect 3224 3645 3276 3654
rect 3288 3688 3340 3697
rect 3288 3654 3291 3688
rect 3291 3654 3325 3688
rect 3325 3654 3340 3688
rect 3288 3645 3340 3654
rect 3352 3688 3404 3697
rect 3352 3654 3363 3688
rect 3363 3654 3397 3688
rect 3397 3654 3404 3688
rect 3352 3645 3404 3654
rect 3416 3688 3468 3697
rect 3480 3688 3532 3697
rect 3416 3654 3435 3688
rect 3435 3654 3468 3688
rect 3480 3654 3507 3688
rect 3507 3654 3532 3688
rect 3416 3645 3468 3654
rect 3480 3645 3532 3654
rect -597 3565 -545 3617
rect -597 3546 -545 3550
rect -597 3512 -590 3546
rect -590 3512 -556 3546
rect -556 3512 -545 3546
rect -597 3498 -545 3512
rect -597 3474 -545 3483
rect -597 3440 -590 3474
rect -590 3440 -556 3474
rect -556 3440 -545 3474
rect -597 3431 -545 3440
rect -597 3402 -545 3416
rect -597 3368 -590 3402
rect -590 3368 -556 3402
rect -556 3368 -545 3402
rect -597 3364 -545 3368
rect -597 3330 -545 3349
rect -597 3297 -590 3330
rect -590 3297 -556 3330
rect -556 3297 -545 3330
rect -597 3258 -545 3283
rect -597 3231 -590 3258
rect -590 3231 -556 3258
rect -556 3231 -545 3258
rect -597 3186 -545 3217
rect -597 3165 -590 3186
rect -590 3165 -556 3186
rect -556 3165 -545 3186
rect -597 3114 -545 3151
rect -597 3099 -590 3114
rect -590 3099 -556 3114
rect -556 3099 -545 3114
rect -597 3080 -590 3085
rect -590 3080 -556 3085
rect -556 3080 -545 3085
rect -597 3042 -545 3080
rect -597 3033 -590 3042
rect -590 3033 -556 3042
rect -556 3033 -545 3042
rect -597 3008 -590 3019
rect -590 3008 -556 3019
rect -556 3008 -545 3019
rect -597 2970 -545 3008
rect -597 2967 -590 2970
rect -590 2967 -556 2970
rect -556 2967 -545 2970
rect -597 2936 -590 2953
rect -590 2936 -556 2953
rect -556 2936 -545 2953
rect -597 2901 -545 2936
rect -597 2864 -590 2887
rect -590 2864 -556 2887
rect -556 2864 -545 2887
rect -597 2835 -545 2864
rect -597 2792 -590 2821
rect -590 2792 -556 2821
rect -556 2792 -545 2821
rect -597 2769 -545 2792
rect -597 2754 -545 2755
rect -597 2720 -590 2754
rect -590 2720 -556 2754
rect -556 2720 -545 2754
rect -597 2703 -545 2720
rect -597 2682 -545 2689
rect -597 2648 -590 2682
rect -590 2648 -556 2682
rect -556 2648 -545 2682
rect -597 2637 -545 2648
rect -597 2610 -545 2623
rect -597 2576 -590 2610
rect -590 2576 -556 2610
rect -556 2576 -545 2610
rect -597 2571 -545 2576
rect -1703 2213 -1651 2265
rect -1639 2213 -1587 2265
rect -1761 2120 -1709 2172
rect -1761 2056 -1709 2108
rect -805 2219 -753 2271
rect -739 2219 -687 2271
rect -673 2219 -621 2271
rect -606 2219 -554 2271
rect -539 2219 -487 2271
rect -805 2125 -753 2177
rect -739 2125 -687 2177
rect -673 2125 -621 2177
rect -606 2125 -554 2177
rect -539 2125 -487 2177
rect -716 1690 -664 1699
rect -716 1656 -710 1690
rect -710 1656 -676 1690
rect -676 1656 -664 1690
rect -716 1647 -664 1656
rect -650 1690 -598 1699
rect -650 1656 -638 1690
rect -638 1656 -604 1690
rect -604 1656 -598 1690
rect -650 1647 -598 1656
rect -725 1348 -673 1400
rect -650 1348 -598 1400
rect -574 1348 -522 1400
rect -498 1348 -446 1400
rect 315 3546 367 3557
rect 315 3512 324 3546
rect 324 3512 358 3546
rect 358 3512 367 3546
rect 315 3505 367 3512
rect 315 3474 367 3493
rect 315 3441 324 3474
rect 324 3441 358 3474
rect 358 3441 367 3474
rect 315 3402 367 3429
rect 315 3377 324 3402
rect 324 3377 358 3402
rect 358 3377 367 3402
rect -11 2380 41 2432
rect -11 2316 41 2368
rect -170 1982 -118 1994
rect -170 1948 -164 1982
rect -164 1948 -130 1982
rect -130 1948 -118 1982
rect -170 1942 -118 1948
rect -102 1982 -50 1994
rect -102 1948 -90 1982
rect -90 1948 -56 1982
rect -56 1948 -50 1982
rect -102 1942 -50 1948
rect 919 3546 971 3557
rect 919 3512 928 3546
rect 928 3512 962 3546
rect 962 3512 971 3546
rect 919 3505 971 3512
rect 919 3474 971 3493
rect 919 3441 928 3474
rect 928 3441 962 3474
rect 962 3441 971 3474
rect 919 3402 971 3429
rect 919 3377 928 3402
rect 928 3377 962 3402
rect 962 3377 971 3402
rect 607 3258 659 3275
rect 607 3224 616 3258
rect 616 3224 650 3258
rect 650 3224 659 3258
rect 607 3223 659 3224
rect 607 3186 659 3211
rect 607 3159 616 3186
rect 616 3159 650 3186
rect 650 3159 659 3186
rect 391 2516 443 2520
rect 391 2482 403 2516
rect 403 2482 437 2516
rect 437 2482 443 2516
rect 391 2468 443 2482
rect 391 2444 443 2456
rect 391 2410 403 2444
rect 403 2410 437 2444
rect 437 2410 443 2444
rect 391 2404 443 2410
rect 1406 3546 1458 3557
rect 1406 3512 1415 3546
rect 1415 3512 1449 3546
rect 1449 3512 1458 3546
rect 1406 3505 1458 3512
rect 1406 3474 1458 3493
rect 1406 3441 1415 3474
rect 1415 3441 1449 3474
rect 1449 3441 1458 3474
rect 1406 3402 1458 3429
rect 1406 3377 1415 3402
rect 1415 3377 1449 3402
rect 1449 3377 1458 3402
rect 1699 3511 1751 3557
rect 1699 3505 1708 3511
rect 1708 3505 1742 3511
rect 1742 3505 1751 3511
rect 1699 3477 1708 3493
rect 1708 3477 1742 3493
rect 1742 3477 1751 3493
rect 1699 3441 1751 3477
rect 1699 3405 1708 3429
rect 1708 3405 1742 3429
rect 1742 3405 1751 3429
rect 1699 3377 1751 3405
rect 1046 3258 1098 3275
rect 1046 3224 1055 3258
rect 1055 3224 1089 3258
rect 1089 3224 1098 3258
rect 1046 3223 1098 3224
rect 1046 3186 1098 3211
rect 1046 3159 1055 3186
rect 1055 3159 1089 3186
rect 1089 3159 1098 3186
rect 763 3080 772 3089
rect 772 3080 806 3089
rect 806 3080 815 3089
rect 763 3042 815 3080
rect 763 3037 772 3042
rect 772 3037 806 3042
rect 806 3037 815 3042
rect 763 3008 772 3025
rect 772 3008 806 3025
rect 806 3008 815 3025
rect 763 2973 815 3008
rect 1124 2831 1176 2883
rect 1124 2767 1176 2819
rect 613 2435 665 2487
rect 677 2482 695 2487
rect 695 2482 729 2487
rect 677 2444 729 2482
rect 677 2435 695 2444
rect 695 2435 729 2444
rect 480 2310 532 2362
rect 544 2310 596 2362
rect 851 2335 903 2387
rect 915 2335 967 2387
rect 446 2063 480 2092
rect 480 2063 498 2092
rect 510 2063 514 2092
rect 514 2063 562 2092
rect 446 2040 498 2063
rect 510 2040 562 2063
rect 771 2120 823 2129
rect 771 2086 778 2120
rect 778 2086 812 2120
rect 812 2086 823 2120
rect 771 2077 823 2086
rect 837 2120 889 2129
rect 904 2120 956 2129
rect 971 2120 1023 2129
rect 1038 2120 1090 2129
rect 837 2086 862 2120
rect 862 2086 889 2120
rect 904 2086 946 2120
rect 946 2086 956 2120
rect 971 2086 980 2120
rect 980 2086 1023 2120
rect 1038 2086 1064 2120
rect 1064 2086 1090 2120
rect 837 2077 889 2086
rect 904 2077 956 2086
rect 971 2077 1023 2086
rect 1038 2077 1090 2086
rect 1105 2120 1157 2129
rect 1105 2086 1114 2120
rect 1114 2086 1148 2120
rect 1148 2086 1157 2120
rect 1105 2077 1157 2086
rect 1412 2461 1464 2513
rect 1476 2482 1494 2513
rect 1494 2482 1528 2513
rect 1476 2461 1528 2482
rect 1299 2094 1351 2127
rect 1299 2075 1333 2094
rect 1333 2075 1351 2094
rect 1395 2094 1447 2127
rect 1395 2075 1413 2094
rect 1413 2075 1447 2094
rect 1688 2335 1740 2387
rect 1752 2375 1770 2387
rect 1770 2375 1804 2387
rect 1752 2335 1804 2375
rect 1933 2692 1985 2744
rect 1933 2628 1985 2680
rect 1782 2255 1834 2307
rect 1846 2255 1898 2307
rect 2458 3558 2510 3562
rect 2458 3524 2467 3558
rect 2467 3524 2501 3558
rect 2501 3524 2510 3558
rect 2458 3510 2510 3524
rect 2458 3486 2510 3498
rect 2458 3452 2467 3486
rect 2467 3452 2501 3486
rect 2501 3452 2510 3486
rect 2458 3446 2510 3452
rect 2299 2987 2351 3039
rect 2748 3549 2800 3561
rect 2748 3515 2757 3549
rect 2757 3515 2791 3549
rect 2791 3515 2800 3549
rect 2748 3509 2800 3515
rect 2748 3477 2800 3496
rect 2748 3444 2757 3477
rect 2757 3444 2791 3477
rect 2791 3444 2800 3477
rect 2748 3405 2800 3430
rect 2748 3378 2757 3405
rect 2757 3378 2791 3405
rect 2791 3378 2800 3405
rect 3031 3549 3083 3561
rect 3031 3515 3040 3549
rect 3040 3515 3074 3549
rect 3074 3515 3083 3549
rect 3031 3509 3083 3515
rect 3031 3477 3083 3496
rect 3031 3444 3040 3477
rect 3040 3444 3074 3477
rect 3074 3444 3083 3477
rect 3031 3405 3083 3430
rect 3031 3378 3040 3405
rect 3040 3378 3074 3405
rect 3074 3378 3083 3405
rect 3343 3549 3395 3561
rect 3343 3515 3352 3549
rect 3352 3515 3386 3549
rect 3386 3515 3395 3549
rect 3343 3509 3395 3515
rect 3343 3477 3395 3496
rect 3343 3444 3352 3477
rect 3352 3444 3386 3477
rect 3386 3444 3395 3477
rect 3343 3405 3395 3430
rect 3343 3378 3352 3405
rect 3352 3378 3386 3405
rect 3386 3378 3395 3405
rect 2299 2923 2351 2975
rect 2099 2481 2151 2487
rect 2099 2447 2133 2481
rect 2133 2447 2151 2481
rect 2099 2435 2151 2447
rect 2163 2435 2215 2487
rect 2740 2917 2792 2969
rect 2804 2917 2856 2969
rect 3187 3227 3196 3228
rect 3196 3227 3230 3228
rect 3230 3227 3239 3228
rect 3187 3189 3239 3227
rect 3187 3176 3196 3189
rect 3196 3176 3230 3189
rect 3230 3176 3239 3189
rect 3187 3155 3196 3164
rect 3196 3155 3230 3164
rect 3230 3155 3239 3164
rect 3187 3117 3239 3155
rect 3187 3112 3196 3117
rect 3196 3112 3230 3117
rect 3230 3112 3239 3117
rect 3500 3227 3508 3228
rect 3508 3227 3542 3228
rect 3542 3227 3552 3228
rect 3500 3189 3552 3227
rect 3500 3176 3508 3189
rect 3508 3176 3542 3189
rect 3542 3176 3552 3189
rect 3500 3155 3508 3164
rect 3508 3155 3542 3164
rect 3542 3155 3552 3164
rect 3500 3117 3552 3155
rect 3500 3112 3508 3117
rect 3508 3112 3542 3117
rect 3542 3112 3552 3117
rect 3929 3236 3981 3237
rect 3929 3202 3938 3236
rect 3938 3202 3972 3236
rect 3972 3202 3981 3236
rect 3929 3185 3981 3202
rect 3929 3084 3981 3125
rect 3929 3073 3938 3084
rect 3938 3073 3972 3084
rect 3972 3073 3981 3084
rect 4241 2435 4293 2487
rect 4305 2481 4357 2487
rect 4305 2447 4323 2481
rect 4323 2447 4357 2481
rect 4305 2435 4357 2447
rect 3953 2335 4005 2387
rect 4017 2335 4069 2387
rect 1938 2175 1990 2227
rect 2002 2175 2054 2227
rect 2146 2239 2198 2248
rect 2146 2205 2152 2239
rect 2152 2205 2186 2239
rect 2186 2205 2198 2239
rect 2146 2196 2198 2205
rect 2212 2239 2264 2248
rect 2212 2205 2224 2239
rect 2224 2205 2258 2239
rect 2258 2205 2264 2239
rect 2212 2196 2264 2205
rect 1754 1983 1806 1989
rect 1754 1949 1772 1983
rect 1772 1949 1806 1983
rect 1754 1937 1806 1949
rect 1821 1937 1873 1989
rect 1888 1937 1940 1989
rect 1955 1937 2007 1989
rect -230 1507 -178 1518
rect -230 1473 -221 1507
rect -221 1473 -187 1507
rect -187 1473 -178 1507
rect -230 1466 -178 1473
rect -230 1435 -178 1454
rect -230 1402 -221 1435
rect -221 1402 -187 1435
rect -187 1402 -178 1435
rect -310 1247 -258 1299
rect -310 1183 -258 1235
rect 333 1689 342 1693
rect 342 1689 376 1693
rect 376 1689 385 1693
rect 333 1651 385 1689
rect 333 1641 342 1651
rect 342 1641 376 1651
rect 376 1641 385 1651
rect 333 1617 342 1629
rect 342 1617 376 1629
rect 376 1617 385 1629
rect 333 1579 385 1617
rect 333 1577 342 1579
rect 342 1577 376 1579
rect 376 1577 385 1579
rect 117 1507 169 1518
rect 117 1473 126 1507
rect 126 1473 160 1507
rect 160 1473 169 1507
rect 117 1466 169 1473
rect 117 1435 169 1454
rect 117 1402 126 1435
rect 126 1402 160 1435
rect 160 1402 169 1435
rect 549 1507 601 1518
rect 549 1473 558 1507
rect 558 1473 592 1507
rect 592 1473 601 1507
rect 549 1466 601 1473
rect 549 1435 601 1454
rect 549 1402 558 1435
rect 558 1402 592 1435
rect 592 1402 601 1435
rect 1197 1833 1206 1863
rect 1206 1833 1240 1863
rect 1240 1833 1249 1863
rect 1197 1811 1249 1833
rect 1197 1795 1249 1799
rect 1197 1761 1206 1795
rect 1206 1761 1240 1795
rect 1240 1761 1249 1795
rect 1197 1747 1249 1761
rect 981 1507 1033 1518
rect 981 1473 990 1507
rect 990 1473 1024 1507
rect 1024 1473 1033 1507
rect 981 1466 1033 1473
rect 981 1435 1033 1454
rect 981 1402 990 1435
rect 990 1402 1024 1435
rect 1024 1402 1033 1435
rect 1629 1833 1638 1863
rect 1638 1833 1672 1863
rect 1672 1833 1681 1863
rect 1629 1811 1681 1833
rect 1629 1795 1681 1799
rect 1629 1761 1638 1795
rect 1638 1761 1672 1795
rect 1672 1761 1681 1795
rect 1629 1747 1681 1761
rect 765 1075 817 1077
rect 765 1041 774 1075
rect 774 1041 808 1075
rect 808 1041 817 1075
rect 765 1025 817 1041
rect 765 1003 817 1013
rect 765 969 774 1003
rect 774 969 808 1003
rect 808 969 817 1003
rect 765 961 817 969
rect 765 931 817 949
rect 765 897 774 931
rect 774 897 808 931
rect 808 897 817 931
rect 1413 1507 1465 1518
rect 1413 1473 1422 1507
rect 1422 1473 1456 1507
rect 1456 1473 1465 1507
rect 1413 1466 1465 1473
rect 1413 1435 1465 1454
rect 1413 1402 1422 1435
rect 1422 1402 1456 1435
rect 1456 1402 1465 1435
rect 1964 1641 2016 1693
rect 1964 1577 2016 1629
rect 1845 1507 1897 1518
rect 1845 1473 1854 1507
rect 1854 1473 1888 1507
rect 1888 1473 1897 1507
rect 1845 1466 1897 1473
rect 1845 1435 1897 1454
rect 1845 1402 1854 1435
rect 1854 1402 1888 1435
rect 1888 1402 1897 1435
rect 2476 2041 2528 2059
rect 2476 2007 2488 2041
rect 2488 2007 2522 2041
rect 2522 2007 2528 2041
rect 2476 1969 2528 1995
rect 2476 1943 2488 1969
rect 2488 1943 2522 1969
rect 2522 1943 2528 1969
rect 2803 2172 2855 2224
rect 2867 2172 2919 2224
rect 3116 2158 3168 2210
rect 3180 2158 3232 2210
rect 2691 1937 2743 1989
rect 2755 1983 2807 1989
rect 2755 1949 2785 1983
rect 2785 1949 2807 1983
rect 2755 1937 2807 1949
rect 3249 1983 3301 1995
rect 3249 1949 3267 1983
rect 3267 1949 3301 1983
rect 3249 1943 3301 1949
rect 3313 1943 3365 1995
rect 2844 1801 2896 1836
rect 2844 1784 2853 1801
rect 2853 1784 2887 1801
rect 2887 1784 2896 1801
rect 2844 1767 2853 1772
rect 2853 1767 2887 1772
rect 2887 1767 2896 1772
rect 2844 1729 2896 1767
rect 2844 1720 2853 1729
rect 2853 1720 2887 1729
rect 2887 1720 2896 1729
rect 2122 1025 2174 1077
rect 2122 961 2174 1013
rect 2122 897 2174 949
rect 2404 1025 2456 1077
rect 2404 961 2456 1013
rect 2404 897 2456 949
rect 2688 1047 2697 1077
rect 2697 1047 2731 1077
rect 2731 1047 2740 1077
rect 2688 1025 2740 1047
rect 2688 1009 2740 1013
rect 2688 975 2697 1009
rect 2697 975 2731 1009
rect 2731 975 2740 1009
rect 2688 961 2740 975
rect 2688 937 2740 949
rect 2688 903 2697 937
rect 2697 903 2731 937
rect 2731 903 2740 937
rect 2688 897 2740 903
rect 3156 1801 3208 1836
rect 3156 1784 3165 1801
rect 3165 1784 3199 1801
rect 3199 1784 3208 1801
rect 3156 1767 3165 1772
rect 3165 1767 3199 1772
rect 3199 1767 3208 1772
rect 3156 1729 3208 1767
rect 3156 1720 3165 1729
rect 3165 1720 3199 1729
rect 3199 1720 3208 1729
rect 3000 1047 3009 1077
rect 3009 1047 3043 1077
rect 3043 1047 3052 1077
rect 3000 1025 3052 1047
rect 3000 1009 3052 1013
rect 3000 975 3009 1009
rect 3009 975 3043 1009
rect 3043 975 3052 1009
rect 3000 961 3052 975
rect 3000 937 3052 949
rect 3000 903 3009 937
rect 3009 903 3043 937
rect 3043 903 3052 937
rect 3000 897 3052 903
rect 3315 1047 3321 1077
rect 3321 1047 3355 1077
rect 3355 1047 3367 1077
rect 3315 1025 3367 1047
rect 3436 1025 3488 1077
rect 3315 1009 3367 1013
rect 3315 975 3321 1009
rect 3321 975 3355 1009
rect 3355 975 3367 1009
rect 3315 961 3367 975
rect 3436 949 3488 1001
rect 3315 937 3367 949
rect 3315 903 3321 937
rect 3321 903 3355 937
rect 3355 903 3367 937
rect 3315 897 3367 903
rect 3436 872 3488 924
rect 169 832 221 841
rect 234 832 286 841
rect 299 832 351 841
rect 169 798 184 832
rect 184 798 221 832
rect 234 798 257 832
rect 257 798 286 832
rect 299 798 330 832
rect 330 798 351 832
rect 169 789 221 798
rect 234 789 286 798
rect 299 789 351 798
rect 363 832 415 841
rect 363 798 369 832
rect 369 798 403 832
rect 403 798 415 832
rect 363 789 415 798
rect 427 832 479 841
rect 427 798 441 832
rect 441 798 475 832
rect 475 798 479 832
rect 427 789 479 798
rect 491 832 543 841
rect 555 832 607 841
rect 619 832 671 841
rect 683 832 735 841
rect 747 832 799 841
rect 811 832 863 841
rect 875 832 927 841
rect 491 798 513 832
rect 513 798 543 832
rect 555 798 585 832
rect 585 798 607 832
rect 619 798 657 832
rect 657 798 671 832
rect 683 798 691 832
rect 691 798 729 832
rect 729 798 735 832
rect 747 798 763 832
rect 763 798 799 832
rect 811 798 835 832
rect 835 798 863 832
rect 875 798 907 832
rect 907 798 927 832
rect 491 789 543 798
rect 555 789 607 798
rect 619 789 671 798
rect 683 789 735 798
rect 747 789 799 798
rect 811 789 863 798
rect 875 789 927 798
rect 939 832 991 841
rect 939 798 945 832
rect 945 798 979 832
rect 979 798 991 832
rect 939 789 991 798
rect 1003 832 1055 841
rect 1003 798 1017 832
rect 1017 798 1051 832
rect 1051 798 1055 832
rect 1003 789 1055 798
rect 1067 832 1119 841
rect 1131 832 1183 841
rect 1195 832 1247 841
rect 1259 832 1311 841
rect 1323 832 1375 841
rect 1387 832 1439 841
rect 1451 832 1503 841
rect 1067 798 1089 832
rect 1089 798 1119 832
rect 1131 798 1161 832
rect 1161 798 1183 832
rect 1195 798 1233 832
rect 1233 798 1247 832
rect 1259 798 1267 832
rect 1267 798 1305 832
rect 1305 798 1311 832
rect 1323 798 1339 832
rect 1339 798 1375 832
rect 1387 798 1411 832
rect 1411 798 1439 832
rect 1451 798 1483 832
rect 1483 798 1503 832
rect 1067 789 1119 798
rect 1131 789 1183 798
rect 1195 789 1247 798
rect 1259 789 1311 798
rect 1323 789 1375 798
rect 1387 789 1439 798
rect 1451 789 1503 798
rect 1515 832 1567 841
rect 1515 798 1521 832
rect 1521 798 1555 832
rect 1555 798 1567 832
rect 1515 789 1567 798
rect 1579 832 1631 841
rect 1579 798 1593 832
rect 1593 798 1627 832
rect 1627 798 1631 832
rect 1579 789 1631 798
rect 1643 832 1695 841
rect 1707 832 1759 841
rect 1771 832 1823 841
rect 1835 832 1887 841
rect 1899 832 1951 841
rect 1963 832 2015 841
rect 2027 832 2079 841
rect 1643 798 1665 832
rect 1665 798 1695 832
rect 1707 798 1737 832
rect 1737 798 1759 832
rect 1771 798 1809 832
rect 1809 798 1823 832
rect 1835 798 1843 832
rect 1843 798 1881 832
rect 1881 798 1887 832
rect 1899 798 1915 832
rect 1915 798 1951 832
rect 1963 798 1987 832
rect 1987 798 2015 832
rect 2027 798 2059 832
rect 2059 798 2079 832
rect 1643 789 1695 798
rect 1707 789 1759 798
rect 1771 789 1823 798
rect 1835 789 1887 798
rect 1899 789 1951 798
rect 1963 789 2015 798
rect 2027 789 2079 798
rect 2091 832 2143 841
rect 2091 798 2097 832
rect 2097 798 2131 832
rect 2131 798 2143 832
rect 2091 789 2143 798
rect 2155 832 2207 841
rect 2155 798 2169 832
rect 2169 798 2203 832
rect 2203 798 2207 832
rect 2155 789 2207 798
rect 2219 832 2271 841
rect 2283 832 2335 841
rect 2347 832 2399 841
rect 2411 832 2463 841
rect 2475 832 2527 841
rect 2539 832 2591 841
rect 2603 832 2655 841
rect 2219 798 2241 832
rect 2241 798 2271 832
rect 2283 798 2313 832
rect 2313 798 2335 832
rect 2347 798 2385 832
rect 2385 798 2399 832
rect 2411 798 2419 832
rect 2419 798 2457 832
rect 2457 798 2463 832
rect 2475 798 2491 832
rect 2491 798 2527 832
rect 2539 798 2563 832
rect 2563 798 2591 832
rect 2603 798 2635 832
rect 2635 798 2655 832
rect 2219 789 2271 798
rect 2283 789 2335 798
rect 2347 789 2399 798
rect 2411 789 2463 798
rect 2475 789 2527 798
rect 2539 789 2591 798
rect 2603 789 2655 798
rect 2667 832 2719 841
rect 2667 798 2673 832
rect 2673 798 2707 832
rect 2707 798 2719 832
rect 2667 789 2719 798
rect 2731 832 2783 841
rect 2731 798 2745 832
rect 2745 798 2779 832
rect 2779 798 2783 832
rect 2731 789 2783 798
rect 2795 832 2847 841
rect 2859 832 2911 841
rect 2923 832 2975 841
rect 2987 832 3039 841
rect 3051 832 3103 841
rect 3115 832 3167 841
rect 3179 832 3231 841
rect 2795 798 2817 832
rect 2817 798 2847 832
rect 2859 798 2889 832
rect 2889 798 2911 832
rect 2923 798 2961 832
rect 2961 798 2975 832
rect 2987 798 2995 832
rect 2995 798 3033 832
rect 3033 798 3039 832
rect 3051 798 3067 832
rect 3067 798 3103 832
rect 3115 798 3139 832
rect 3139 798 3167 832
rect 3179 798 3211 832
rect 3211 798 3231 832
rect 2795 789 2847 798
rect 2859 789 2911 798
rect 2923 789 2975 798
rect 2987 789 3039 798
rect 3051 789 3103 798
rect 3115 789 3167 798
rect 3179 789 3231 798
rect 3243 832 3295 841
rect 3243 798 3249 832
rect 3249 798 3283 832
rect 3283 798 3295 832
rect 3243 789 3295 798
rect 3307 832 3359 841
rect 3307 798 3321 832
rect 3321 798 3355 832
rect 3355 798 3359 832
rect 3307 789 3359 798
rect 3436 795 3488 847
rect 3879 1833 3931 1836
rect 3879 1799 3889 1833
rect 3889 1799 3923 1833
rect 3923 1799 3931 1833
rect 3879 1784 3931 1799
rect 3879 1761 3931 1772
rect 3879 1727 3889 1761
rect 3889 1727 3923 1761
rect 3923 1727 3931 1761
rect 3879 1720 3931 1727
rect 2687 683 2739 716
rect 1291 674 1343 680
rect 1372 674 1424 680
rect 1291 640 1321 674
rect 1321 640 1343 674
rect 1372 640 1393 674
rect 1393 640 1424 674
rect 1291 628 1343 640
rect 1372 628 1424 640
rect 2687 664 2697 683
rect 2697 664 2731 683
rect 2731 664 2739 683
rect 2687 649 2697 652
rect 2697 649 2731 652
rect 2731 649 2739 652
rect 2687 611 2739 649
rect 2687 600 2697 611
rect 2697 600 2731 611
rect 2731 600 2739 611
rect 66 515 118 567
rect 130 515 182 567
rect 3000 683 3052 716
rect 3000 664 3009 683
rect 3009 664 3043 683
rect 3043 664 3052 683
rect 3000 649 3009 652
rect 3009 649 3043 652
rect 3043 649 3052 652
rect 3000 611 3052 649
rect 3000 600 3009 611
rect 3009 600 3043 611
rect 3043 600 3052 611
rect 2813 505 2853 535
rect 2853 505 2865 535
rect 2877 505 2887 535
rect 2887 505 2929 535
rect 2813 483 2865 505
rect 2877 483 2929 505
rect 3143 505 3165 535
rect 3165 505 3195 535
rect 3143 483 3195 505
rect 3207 483 3259 535
rect 3807 1177 3859 1229
rect 3871 1177 3923 1229
rect 3709 1048 3740 1072
rect 3740 1048 3761 1072
rect 3709 1020 3761 1048
rect 3793 1048 3802 1072
rect 3802 1048 3836 1072
rect 3836 1048 3845 1072
rect 3793 1020 3845 1048
rect 3877 1048 3898 1072
rect 3898 1048 3929 1072
rect 3877 1020 3929 1048
rect 3709 972 3740 1000
rect 3740 972 3761 1000
rect 3709 948 3761 972
rect 3793 972 3802 1000
rect 3802 972 3836 1000
rect 3836 972 3845 1000
rect 3793 948 3845 972
rect 3877 972 3898 1000
rect 3898 972 3929 1000
rect 3877 948 3929 972
rect 3709 896 3740 928
rect 3740 896 3761 928
rect 3709 876 3761 896
rect 3793 896 3802 928
rect 3802 896 3836 928
rect 3836 896 3845 928
rect 3793 876 3845 896
rect 3877 896 3898 928
rect 3898 896 3929 928
rect 3877 876 3929 896
rect 3709 854 3761 856
rect 3709 820 3740 854
rect 3740 820 3761 854
rect 3709 804 3761 820
rect 3793 854 3845 856
rect 3793 820 3802 854
rect 3802 820 3836 854
rect 3836 820 3845 854
rect 3793 804 3845 820
rect 3877 854 3929 856
rect 3877 820 3898 854
rect 3898 820 3929 854
rect 3877 804 3929 820
rect 4715 3228 4767 3235
rect 4715 3194 4718 3228
rect 4718 3194 4752 3228
rect 4752 3194 4767 3228
rect 4715 3183 4767 3194
rect 4793 3228 4845 3235
rect 4793 3194 4802 3228
rect 4802 3194 4836 3228
rect 4836 3194 4845 3228
rect 4793 3183 4845 3194
rect 4871 3228 4923 3235
rect 4871 3194 4886 3228
rect 4886 3194 4920 3228
rect 4920 3194 4923 3228
rect 4871 3183 4923 3194
rect 4715 3119 4718 3125
rect 4718 3119 4752 3125
rect 4752 3119 4767 3125
rect 4715 3078 4767 3119
rect 4715 3073 4718 3078
rect 4718 3073 4752 3078
rect 4752 3073 4767 3078
rect 4793 3119 4802 3125
rect 4802 3119 4836 3125
rect 4836 3119 4845 3125
rect 4793 3078 4845 3119
rect 4793 3073 4802 3078
rect 4802 3073 4836 3078
rect 4836 3073 4845 3078
rect 4871 3119 4886 3125
rect 4886 3119 4920 3125
rect 4920 3119 4923 3125
rect 4871 3078 4923 3119
rect 4871 3073 4886 3078
rect 4886 3073 4920 3078
rect 4920 3073 4923 3078
rect 4620 2979 4672 3031
rect 4620 2915 4672 2967
rect 5426 2979 5478 3031
rect 5426 2956 5478 2967
rect 5321 2936 5373 2942
rect 5321 2902 5329 2936
rect 5329 2902 5363 2936
rect 5363 2902 5373 2936
rect 5321 2890 5373 2902
rect 5321 2864 5373 2878
rect 5321 2830 5329 2864
rect 5329 2830 5363 2864
rect 5363 2830 5373 2864
rect 5321 2826 5373 2830
rect 5426 2922 5432 2956
rect 5432 2922 5466 2956
rect 5466 2922 5478 2956
rect 5426 2915 5478 2922
rect 5733 3265 5785 3308
rect 5733 3256 5738 3265
rect 5738 3256 5772 3265
rect 5772 3256 5785 3265
rect 5811 3283 5829 3308
rect 5829 3283 5863 3308
rect 5811 3256 5863 3283
rect 5889 3283 5901 3308
rect 5901 3283 5935 3308
rect 5935 3283 5941 3308
rect 5889 3256 5941 3283
rect 6568 3317 6620 3358
rect 6568 3306 6580 3317
rect 6580 3306 6614 3317
rect 6614 3306 6620 3317
rect 6640 3317 6692 3358
rect 6640 3306 6652 3317
rect 6652 3306 6686 3317
rect 6686 3306 6692 3317
rect 6712 3333 6764 3358
rect 6712 3306 6730 3333
rect 6730 3306 6764 3333
rect 5733 3187 5785 3220
rect 5733 3168 5738 3187
rect 5738 3168 5772 3187
rect 5772 3168 5785 3187
rect 5811 3168 5863 3220
rect 5889 3168 5941 3220
rect 5733 3109 5785 3132
rect 5733 3080 5738 3109
rect 5738 3080 5772 3109
rect 5772 3080 5785 3109
rect 5811 3080 5863 3132
rect 5889 3080 5941 3132
rect 5545 2709 5597 2711
rect 5545 2675 5551 2709
rect 5551 2675 5585 2709
rect 5585 2675 5597 2709
rect 5212 2622 5264 2674
rect 5276 2622 5328 2674
rect 5545 2659 5597 2675
rect 5545 2595 5597 2647
rect 5210 2521 5262 2573
rect 5274 2521 5326 2573
rect 6568 3217 6620 3269
rect 6640 3217 6692 3269
rect 6712 3253 6764 3269
rect 6712 3219 6730 3253
rect 6730 3219 6764 3253
rect 6712 3217 6764 3219
rect 6568 3129 6620 3181
rect 6640 3129 6692 3181
rect 6712 3174 6764 3181
rect 6712 3140 6730 3174
rect 6730 3140 6764 3174
rect 6712 3129 6764 3140
rect 6253 2664 6305 2670
rect 6253 2630 6259 2664
rect 6259 2630 6293 2664
rect 6293 2630 6305 2664
rect 6253 2618 6305 2630
rect 6319 2664 6371 2670
rect 6319 2630 6331 2664
rect 6331 2630 6365 2664
rect 6365 2630 6371 2664
rect 6319 2618 6371 2630
rect 5509 2289 5561 2301
rect 5573 2289 5625 2301
rect 5509 2255 5545 2289
rect 5545 2255 5561 2289
rect 5573 2255 5579 2289
rect 5579 2255 5625 2289
rect 5509 2249 5561 2255
rect 5573 2249 5625 2255
rect 5505 2166 5557 2218
rect 5569 2166 5621 2218
rect 6085 2166 6137 2218
rect 6149 2166 6201 2218
rect 4228 1943 4280 1995
rect 4292 1943 4344 1995
rect 4289 1614 4341 1666
rect 4289 1550 4341 1602
rect 248 311 300 320
rect 328 311 380 320
rect 408 311 460 320
rect 488 311 540 320
rect 248 277 275 311
rect 275 277 300 311
rect 328 277 347 311
rect 347 277 380 311
rect 408 277 419 311
rect 419 277 457 311
rect 457 277 460 311
rect 488 277 491 311
rect 491 277 529 311
rect 529 277 540 311
rect 248 268 300 277
rect 328 268 380 277
rect 408 268 460 277
rect 488 268 540 277
rect 248 139 300 191
rect 328 139 380 191
rect 408 139 460 191
rect 488 139 540 191
rect 248 75 300 84
rect 328 75 380 84
rect 408 75 460 84
rect 488 75 540 84
rect 248 41 275 75
rect 275 41 300 75
rect 328 41 347 75
rect 347 41 380 75
rect 408 41 419 75
rect 419 41 457 75
rect 457 41 460 75
rect 488 41 491 75
rect 491 41 529 75
rect 529 41 540 75
rect 248 32 300 41
rect 328 32 380 41
rect 408 32 460 41
rect 488 32 540 41
<< metal2 >>
rect -28256 4895 -22087 4896
tri -22087 4895 -22086 4896 sw
rect -28256 4843 -28196 4895
rect -28144 4843 -28132 4895
rect -28080 4843 -28068 4895
rect -28016 4843 -28004 4895
rect -27952 4843 -27940 4895
rect -27888 4843 -27876 4895
rect -27824 4843 -27812 4895
rect -27760 4843 -27748 4895
rect -27696 4843 -27684 4895
rect -27632 4843 -27620 4895
rect -27568 4843 -27555 4895
rect -27503 4843 -27490 4895
rect -27438 4843 -27425 4895
rect -27373 4843 -27360 4895
rect -27308 4843 -27295 4895
rect -27243 4843 -27230 4895
rect -27178 4843 -27165 4895
rect -27113 4843 -22086 4895
rect -28256 4773 -22086 4843
rect -28256 4721 -28196 4773
rect -28144 4721 -28132 4773
rect -28080 4721 -28068 4773
rect -28016 4721 -28004 4773
rect -27952 4721 -27940 4773
rect -27888 4721 -27876 4773
rect -27824 4721 -27812 4773
rect -27760 4721 -27748 4773
rect -27696 4721 -27684 4773
rect -27632 4721 -27620 4773
rect -27568 4721 -27555 4773
rect -27503 4721 -27490 4773
rect -27438 4721 -27425 4773
rect -27373 4721 -27360 4773
rect -27308 4721 -27295 4773
rect -27243 4721 -27230 4773
rect -27178 4721 -27165 4773
rect -27113 4721 -22086 4773
tri -22086 4721 -21912 4895 sw
rect -28256 4717 -21912 4721
tri -22160 4696 -22139 4717 ne
rect -22139 4696 -21912 4717
tri -21912 4696 -21887 4721 sw
tri -22139 4644 -22087 4696 ne
rect -22087 4644 -21221 4696
rect -21169 4644 -21145 4696
rect -21093 4644 -21069 4696
rect -21017 4644 -20993 4696
rect -20941 4644 -20917 4696
rect -20865 4644 -20841 4696
rect -20789 4644 -20783 4696
tri -22087 4570 -22013 4644 ne
rect -22013 4570 -20783 4644
tri -22013 4518 -21961 4570 ne
rect -21961 4518 -21221 4570
rect -21169 4518 -21145 4570
rect -21093 4518 -21069 4570
rect -21017 4518 -20993 4570
rect -20941 4518 -20917 4570
rect -20865 4518 -20841 4570
rect -20789 4518 -20783 4570
rect -812 3802 735 4150
tri 4028 3802 4100 3874 se
rect 4100 3802 6420 3874
rect -812 3705 -391 3802
tri -391 3705 -294 3802 nw
tri 3931 3705 4028 3802 se
rect 4028 3705 6420 3802
rect -812 3700 -396 3705
tri -396 3700 -391 3705 nw
rect -812 3648 -787 3700
rect -735 3648 -717 3700
rect -665 3648 -646 3700
rect -594 3648 -575 3700
rect -523 3648 -504 3700
rect -452 3697 -399 3700
tri -399 3697 -396 3700 nw
rect 94 3697 6420 3705
tri 6420 3697 6597 3874 sw
rect -452 3648 -446 3697
tri -446 3650 -399 3697 nw
rect -812 3617 -446 3648
rect -812 3565 -597 3617
rect -545 3565 -446 3617
rect -812 3550 -446 3565
rect -812 3498 -597 3550
rect -545 3498 -446 3550
rect -812 3483 -446 3498
rect -812 3431 -597 3483
rect -545 3431 -446 3483
rect -812 3416 -446 3431
rect -812 3364 -597 3416
rect -545 3364 -446 3416
rect 94 3645 170 3697
rect 222 3645 235 3697
rect 287 3645 300 3697
rect 352 3645 365 3697
rect 417 3645 430 3697
rect 482 3645 495 3697
rect 547 3645 560 3697
rect 612 3645 625 3697
rect 677 3645 690 3697
rect 742 3645 755 3697
rect 807 3645 820 3697
rect 872 3645 885 3697
rect 937 3645 950 3697
rect 1002 3645 1015 3697
rect 1067 3645 1080 3697
rect 1132 3645 1145 3697
rect 1197 3645 1210 3697
rect 1262 3645 1275 3697
rect 1327 3645 1340 3697
rect 1392 3645 1405 3697
rect 1457 3645 1470 3697
rect 1522 3645 1535 3697
rect 1587 3645 1600 3697
rect 1652 3645 1665 3697
rect 1717 3645 1730 3697
rect 1782 3645 1795 3697
rect 1847 3645 1860 3697
rect 1912 3645 1925 3697
rect 1977 3645 1990 3697
rect 2042 3645 2055 3697
rect 2107 3645 2120 3697
rect 2172 3645 2185 3697
rect 2237 3645 2250 3697
rect 2302 3645 2315 3697
rect 2367 3645 2380 3697
rect 2432 3645 2445 3697
rect 2497 3645 2510 3697
rect 2562 3645 2575 3697
rect 2627 3645 2640 3697
rect 2692 3645 2705 3697
rect 2757 3645 2770 3697
rect 2822 3645 2835 3697
rect 2887 3645 2900 3697
rect 2952 3645 2965 3697
rect 3017 3645 3030 3697
rect 3082 3645 3095 3697
rect 3147 3645 3160 3697
rect 3212 3645 3224 3697
rect 3276 3645 3288 3697
rect 3340 3645 3352 3697
rect 3404 3645 3416 3697
rect 3468 3645 3480 3697
rect 3532 3645 6597 3697
tri 6597 3645 6649 3697 sw
rect 94 3568 6649 3645
tri 6649 3568 6726 3645 sw
rect 94 3567 6726 3568
tri 6726 3567 6727 3568 sw
rect 94 3562 6727 3567
rect 94 3557 2458 3562
rect 94 3505 315 3557
rect 367 3505 919 3557
rect 971 3505 1406 3557
rect 1458 3505 1699 3557
rect 1751 3510 2458 3557
rect 2510 3561 6727 3562
rect 2510 3510 2748 3561
rect 1751 3509 2748 3510
rect 2800 3509 3031 3561
rect 3083 3509 3343 3561
rect 3395 3540 6727 3561
rect 3395 3526 4499 3540
tri 4499 3526 4513 3540 nw
tri 6282 3526 6296 3540 ne
rect 6296 3526 6727 3540
tri 6727 3526 6768 3567 sw
rect 3395 3509 4345 3526
rect 1751 3505 4345 3509
rect 94 3498 4345 3505
rect 94 3493 2458 3498
rect 94 3441 315 3493
rect 367 3441 919 3493
rect 971 3441 1406 3493
rect 1458 3441 1699 3493
rect 1751 3446 2458 3493
rect 2510 3496 4345 3498
rect 2510 3446 2748 3496
rect 1751 3444 2748 3446
rect 2800 3444 3031 3496
rect 3083 3444 3343 3496
rect 3395 3444 4345 3496
rect 1751 3441 4345 3444
rect 94 3430 4345 3441
rect 94 3429 2748 3430
rect 94 3377 315 3429
rect 367 3377 919 3429
rect 971 3377 1406 3429
rect 1458 3377 1699 3429
rect 1751 3378 2748 3429
rect 2800 3378 3031 3430
rect 3083 3378 3343 3430
rect 3395 3378 4345 3430
rect 1751 3377 4345 3378
rect 94 3372 4345 3377
tri 4345 3372 4499 3526 nw
tri 6296 3402 6420 3526 ne
rect 6420 3402 6768 3526
tri 6420 3372 6450 3402 ne
rect 6450 3372 6768 3402
rect 94 3371 4344 3372
tri 4344 3371 4345 3372 nw
tri 6450 3371 6451 3372 ne
rect 6451 3371 6768 3372
rect -812 3349 -446 3364
tri 6451 3358 6464 3371 ne
rect 6464 3358 6768 3371
rect -812 3297 -597 3349
rect -545 3297 -446 3349
tri 6464 3317 6505 3358 ne
rect 6505 3317 6568 3358
tri 5193 3314 5196 3317 se
rect 5196 3314 5947 3317
tri 5187 3308 5193 3314 se
rect 5193 3308 5947 3314
rect -812 3283 -446 3297
rect -812 3231 -597 3283
rect -545 3231 -446 3283
tri 5160 3281 5187 3308 se
rect 5187 3281 5733 3308
rect -812 3217 -446 3231
rect -812 3165 -597 3217
rect -545 3165 -446 3217
rect -812 3151 -446 3165
rect 607 3275 1899 3281
rect 659 3223 1046 3275
rect 1098 3245 1899 3275
tri 5135 3256 5160 3281 se
rect 5160 3256 5733 3281
rect 5785 3256 5811 3308
rect 5863 3256 5889 3308
rect 5941 3256 5947 3308
tri 6505 3306 6516 3317 ne
rect 6516 3306 6568 3317
rect 6620 3306 6640 3358
rect 6692 3306 6712 3358
rect 6764 3306 6768 3358
tri 6516 3281 6541 3306 ne
rect 6541 3281 6768 3306
tri 6541 3269 6553 3281 ne
rect 6553 3269 6768 3281
tri 6553 3257 6565 3269 ne
rect 1098 3223 1754 3245
rect 607 3211 1754 3223
rect 659 3159 1046 3211
rect 1098 3189 1754 3211
rect 1810 3189 1834 3245
rect 1890 3189 1899 3245
tri 5122 3243 5135 3256 se
rect 5135 3243 5947 3256
rect 3929 3237 5947 3243
rect 1098 3159 1899 3189
rect 607 3153 1899 3159
rect 2914 3228 3552 3234
rect 2914 3201 3187 3228
rect -812 3099 -597 3151
rect -545 3099 -446 3151
rect 2914 3145 2924 3201
rect 2980 3145 3004 3201
rect 3060 3176 3187 3201
rect 3239 3176 3500 3228
rect 3060 3164 3552 3176
rect 3060 3145 3187 3164
rect 2914 3112 3187 3145
rect 3239 3112 3500 3164
rect 2914 3106 3552 3112
rect 3981 3235 5947 3237
rect 3981 3185 4715 3235
rect 3929 3183 4715 3185
rect 4767 3183 4793 3235
rect 4845 3183 4871 3235
rect 4923 3220 5947 3235
rect 4923 3183 5733 3220
rect 3929 3168 5733 3183
rect 5785 3168 5811 3220
rect 5863 3168 5889 3220
rect 5941 3168 5947 3220
rect 3929 3132 5947 3168
rect 3929 3125 5733 3132
rect -812 3085 -446 3099
rect -812 3033 -597 3085
rect -545 3033 -446 3085
rect -812 3019 -446 3033
rect -812 2967 -597 3019
rect -545 2967 -446 3019
rect 763 3089 1653 3095
rect 815 3059 1653 3089
rect 3981 3073 4715 3125
rect 4767 3073 4793 3125
rect 4845 3073 4871 3125
rect 4923 3080 5733 3125
rect 5785 3080 5811 3132
rect 5863 3080 5889 3132
rect 5941 3080 5947 3132
rect 6565 3217 6568 3269
rect 6620 3217 6640 3269
rect 6692 3217 6712 3269
rect 6764 3217 6768 3269
rect 6565 3181 6768 3217
rect 6565 3129 6568 3181
rect 6620 3129 6640 3181
rect 6692 3129 6712 3181
rect 6764 3129 6768 3181
rect 6565 3123 6768 3129
rect 4923 3073 5947 3080
rect 3929 3067 5947 3073
rect 815 3037 1508 3059
rect 763 3025 1508 3037
rect 815 3003 1508 3025
rect 1564 3003 1588 3059
rect 1644 3003 1653 3059
rect 815 2973 1653 3003
rect 763 2967 1653 2973
rect 2299 3039 2351 3045
rect 4620 3031 5478 3037
rect 2299 2979 2351 2987
tri 2351 2979 2396 3024 sw
rect 4672 2979 5426 3031
rect 2299 2975 2396 2979
rect -812 2953 -446 2967
rect -812 2901 -597 2953
rect -545 2901 -446 2953
rect 2351 2969 2396 2975
tri 2396 2969 2406 2979 sw
rect 2351 2923 2740 2969
rect 2299 2917 2740 2923
rect 2792 2917 2804 2969
rect 2856 2917 2862 2969
rect 4620 2967 4730 2979
tri 4730 2967 4742 2979 nw
tri 5386 2967 5398 2979 ne
rect 5398 2967 5478 2979
tri 1727 2915 1729 2917 se
rect 1729 2915 2209 2917
tri 2209 2915 2211 2917 sw
rect 4672 2948 4711 2967
tri 4711 2948 4730 2967 nw
tri 5398 2948 5417 2967 ne
rect 5417 2948 5426 2967
rect 4672 2942 4705 2948
tri 4705 2942 4711 2948 nw
rect 5321 2942 5373 2948
rect -812 2887 -446 2901
tri 1702 2890 1727 2915 se
rect 1727 2909 2211 2915
tri 2211 2909 2217 2915 sw
rect 4620 2909 4672 2915
tri 4672 2909 4705 2942 nw
tri 5307 2909 5321 2923 se
rect 1727 2890 2217 2909
tri 2217 2890 2236 2909 sw
tri 5288 2890 5307 2909 se
rect 5307 2890 5321 2909
tri 5417 2939 5426 2948 ne
rect 5426 2909 5478 2915
tri 1701 2889 1702 2890 se
rect 1702 2889 2236 2890
tri 2236 2889 2237 2890 sw
tri 5287 2889 5288 2890 se
rect 5288 2889 5373 2890
rect -812 2835 -597 2887
rect -545 2835 -446 2887
rect 1124 2883 4478 2889
rect -812 2821 -446 2835
tri 1084 2831 1091 2838 ne
rect 1091 2831 1124 2838
rect 1176 2878 4478 2883
tri 4478 2878 4489 2889 sw
tri 4729 2878 4740 2889 se
rect 4740 2878 5373 2889
rect 1176 2873 4489 2878
tri 4489 2873 4494 2878 sw
tri 4724 2873 4729 2878 se
rect 4729 2873 5321 2878
rect 1176 2865 5321 2873
rect 1176 2837 1723 2865
tri 1723 2837 1751 2865 nw
tri 2187 2837 2215 2865 ne
rect 2215 2837 5321 2865
rect 1176 2831 1204 2837
tri 1091 2826 1096 2831 ne
rect 1096 2826 1204 2831
tri 1204 2826 1215 2837 nw
tri 4456 2826 4467 2837 ne
rect 4467 2826 4751 2837
tri 4751 2826 4762 2837 nw
tri 5304 2826 5315 2837 ne
rect 5315 2826 5321 2837
rect -812 2769 -597 2821
rect -545 2769 -446 2821
tri 1096 2819 1103 2826 ne
rect 1103 2820 1198 2826
tri 1198 2820 1204 2826 nw
tri 4467 2821 4472 2826 ne
rect 4472 2821 4746 2826
tri 4746 2821 4751 2826 nw
tri 5315 2821 5320 2826 ne
rect 5320 2821 5373 2826
tri 5320 2820 5321 2821 ne
rect 5321 2820 5373 2821
rect 1103 2819 1176 2820
tri 1103 2798 1124 2819 ne
rect -812 2755 -446 2769
tri 1176 2798 1198 2820 nw
rect 1124 2761 1176 2767
rect -812 2703 -597 2755
rect -545 2703 -446 2755
tri 1927 2744 1933 2750 se
rect 1933 2744 1985 2750
rect -812 2689 -446 2703
tri 1875 2692 1927 2744 se
rect 1927 2692 1933 2744
tri 1985 2711 2024 2750 sw
rect 5545 2711 5597 2717
rect 1985 2692 2024 2711
rect -812 2637 -597 2689
rect -545 2637 -446 2689
tri 1863 2680 1875 2692 se
rect 1875 2680 2024 2692
tri 1857 2674 1863 2680 se
rect 1863 2674 1933 2680
tri 1246 2664 1256 2674 se
rect 1256 2664 1933 2674
rect -812 2626 -446 2637
rect -812 2623 -450 2626
rect -812 2571 -597 2623
rect -545 2622 -450 2623
tri -450 2622 -446 2626 nw
rect 288 2628 341 2664
tri 341 2628 377 2664 nw
tri 1210 2628 1246 2664 se
rect 1246 2628 1933 2664
rect 1985 2674 2024 2680
tri 2024 2674 2061 2711 sw
rect 1985 2628 5212 2674
rect 288 2622 335 2628
tri 335 2622 341 2628 nw
tri 1204 2622 1210 2628 se
rect 1210 2622 5212 2628
rect 5264 2622 5276 2674
rect 5328 2622 5334 2674
rect 5545 2647 5597 2659
rect -545 2600 -472 2622
tri -472 2600 -450 2622 nw
rect 288 2600 313 2622
tri 313 2600 335 2622 nw
tri 1182 2600 1204 2622 se
rect 1204 2600 1256 2622
tri 1256 2600 1278 2622 nw
rect -545 2595 -477 2600
tri -477 2595 -472 2600 nw
rect 288 2595 308 2600
tri 308 2595 313 2600 nw
tri 1177 2595 1182 2600 se
rect 1182 2595 1251 2600
tri 1251 2595 1256 2600 nw
rect -545 2571 -479 2595
tri -479 2593 -477 2595 nw
rect 288 2593 306 2595
tri 306 2593 308 2595 nw
tri 1175 2593 1177 2595 se
rect 1177 2593 1229 2595
tri 288 2575 306 2593 nw
tri 1157 2575 1175 2593 se
rect 1175 2575 1229 2593
tri 1155 2573 1157 2575 se
rect 1157 2573 1229 2575
tri 1229 2573 1251 2595 nw
rect -812 2271 -479 2571
tri 1108 2526 1155 2573 se
rect 1155 2526 1182 2573
tri 1182 2526 1229 2573 nw
tri 1616 2526 1663 2573 se
rect 1663 2526 5210 2573
rect 391 2521 443 2526
tri 443 2521 448 2526 sw
tri 1103 2521 1108 2526 se
rect 1108 2521 1177 2526
tri 1177 2521 1182 2526 nw
tri 1611 2521 1616 2526 se
rect 1616 2521 5210 2526
rect 5262 2521 5274 2573
rect 5326 2521 5332 2573
rect 391 2520 448 2521
rect 443 2513 448 2520
tri 448 2513 456 2521 sw
tri 1095 2513 1103 2521 se
rect 1103 2513 1169 2521
tri 1169 2513 1177 2521 nw
tri 1603 2513 1611 2521 se
rect 1611 2513 1651 2521
rect 443 2487 456 2513
tri 456 2487 482 2513 sw
tri 1069 2487 1095 2513 se
rect 1095 2487 1143 2513
tri 1143 2487 1169 2513 nw
rect 443 2468 613 2487
rect 391 2456 613 2468
rect -11 2432 41 2438
tri 41 2404 75 2438 sw
rect 443 2435 613 2456
rect 665 2435 677 2487
rect 729 2461 1117 2487
tri 1117 2461 1143 2487 nw
rect 1406 2461 1412 2513
rect 1464 2461 1476 2513
rect 1528 2487 1651 2513
tri 1651 2487 1685 2521 nw
rect 1528 2461 1625 2487
tri 1625 2461 1651 2487 nw
rect 729 2435 1091 2461
tri 1091 2435 1117 2461 nw
rect 2093 2435 2099 2487
rect 2151 2435 2163 2487
rect 2215 2435 4241 2487
rect 4293 2435 4305 2487
rect 4357 2435 4364 2487
rect 41 2398 75 2404
tri 75 2398 81 2404 sw
rect 391 2398 443 2404
tri 443 2398 480 2435 nw
rect 41 2387 81 2398
tri 81 2387 92 2398 sw
rect 41 2380 92 2387
rect -11 2368 92 2380
rect 41 2362 92 2368
tri 92 2362 117 2387 sw
rect 41 2316 480 2362
rect -11 2310 480 2316
rect 532 2310 544 2362
rect 596 2310 602 2362
rect 845 2335 851 2387
rect 903 2335 915 2387
rect 967 2335 1688 2387
rect 1740 2335 1752 2387
rect 1804 2335 3953 2387
rect 4005 2335 4017 2387
rect 4069 2335 4699 2387
tri 4699 2335 4751 2387 sw
tri 5537 2335 5545 2343 se
rect 5545 2335 5597 2595
rect 6247 2618 6253 2670
rect 6305 2618 6319 2670
rect 6371 2618 6377 2670
rect 6247 2516 6377 2618
rect 6247 2487 6348 2516
tri 6348 2487 6377 2516 nw
rect 6247 2460 6321 2487
tri 6321 2460 6348 2487 nw
tri 6222 2435 6247 2460 se
tri 6185 2398 6222 2435 se
rect 6222 2398 6247 2435
tri 6174 2387 6185 2398 se
rect 6185 2387 6247 2398
tri 6173 2386 6174 2387 se
rect 6174 2386 6247 2387
tri 6247 2386 6321 2460 nw
tri 6122 2335 6173 2386 se
rect 6173 2335 6207 2386
tri 6207 2346 6247 2386 nw
tri 4677 2310 4702 2335 ne
rect 4702 2310 4751 2335
tri 4702 2307 4705 2310 ne
rect 4705 2307 4751 2310
rect -1709 2213 -1703 2265
rect -1651 2213 -1639 2265
rect -1587 2246 -1311 2265
tri -1311 2246 -1292 2265 sw
rect -1587 2219 -1292 2246
tri -1292 2219 -1265 2246 sw
rect -812 2219 -805 2271
rect -753 2219 -739 2271
rect -687 2219 -673 2271
rect -621 2219 -606 2271
rect -554 2219 -539 2271
rect -487 2219 -479 2271
tri 605 2265 647 2307 se
rect 647 2265 1782 2307
tri -242 2255 -232 2265 se
rect -232 2255 1782 2265
rect 1834 2255 1846 2307
rect 1898 2255 1904 2307
tri 4705 2301 4711 2307 ne
rect 4711 2301 4751 2307
tri 4751 2301 4785 2335 sw
tri 5503 2301 5537 2335 se
rect 5537 2301 5597 2335
tri 5597 2301 5631 2335 sw
tri 4711 2261 4751 2301 ne
rect 4751 2261 4785 2301
tri 4785 2261 4825 2301 sw
tri 4751 2255 4757 2261 ne
rect 4757 2255 4825 2261
tri -248 2249 -242 2255 se
rect -242 2249 663 2255
tri 663 2249 669 2255 nw
tri 4757 2249 4763 2255 ne
rect 4763 2249 4825 2255
tri 4825 2249 4837 2261 sw
rect 5503 2249 5509 2301
rect 5561 2249 5573 2301
rect 5625 2249 5631 2301
tri 6079 2292 6122 2335 se
rect 6122 2292 6207 2335
tri -249 2248 -248 2249 se
rect -248 2248 662 2249
tri 662 2248 663 2249 nw
tri 4763 2248 4764 2249 ne
rect 4764 2248 4837 2249
tri -270 2227 -249 2248 se
rect -249 2227 641 2248
tri 641 2227 662 2248 nw
rect -1587 2213 -1265 2219
tri -1333 2178 -1298 2213 ne
rect -1298 2191 -1265 2213
tri -1265 2191 -1237 2219 sw
rect -1298 2178 -1237 2191
rect -1761 2177 -1407 2178
tri -1407 2177 -1406 2178 sw
tri -1298 2177 -1297 2178 ne
rect -1297 2177 -1237 2178
tri -1237 2177 -1223 2191 sw
rect -812 2177 -479 2219
tri -306 2191 -270 2227 se
rect -270 2213 627 2227
tri 627 2213 641 2227 nw
tri 702 2224 705 2227 se
rect 705 2224 1938 2227
tri 691 2213 702 2224 se
rect 702 2213 1938 2224
rect -270 2191 -232 2213
tri -232 2191 -210 2213 nw
tri 669 2191 691 2213 se
rect 691 2191 1938 2213
rect -1761 2172 -1406 2177
tri -1406 2172 -1401 2177 sw
tri -1297 2172 -1292 2177 ne
rect -1292 2172 -1223 2177
tri -1223 2172 -1218 2177 sw
rect -1709 2164 -1401 2172
tri -1401 2164 -1393 2172 sw
tri -1292 2164 -1284 2172 ne
rect -1284 2164 -1218 2172
rect -1709 2150 -1393 2164
tri -1393 2150 -1379 2164 sw
tri -1284 2150 -1270 2164 ne
rect -1709 2126 -1379 2150
rect -1709 2125 -1634 2126
tri -1634 2125 -1633 2126 nw
tri -1429 2125 -1428 2126 ne
rect -1428 2125 -1379 2126
tri -1379 2125 -1354 2150 sw
rect -1709 2120 -1667 2125
rect -1761 2108 -1667 2120
rect -1709 2092 -1667 2108
tri -1667 2092 -1634 2125 nw
tri -1428 2092 -1395 2125 ne
rect -1395 2092 -1354 2125
tri -1354 2092 -1321 2125 sw
rect -1709 2090 -1669 2092
tri -1669 2090 -1667 2092 nw
tri -1395 2090 -1393 2092 ne
rect -1393 2090 -1321 2092
tri -1321 2090 -1319 2092 sw
rect -1761 2050 -1709 2056
tri -1709 2050 -1669 2090 nw
tri -1393 2068 -1371 2090 ne
rect -1371 1895 -1319 2090
rect -1270 1956 -1218 2164
rect -812 2125 -805 2177
rect -753 2125 -739 2177
rect -687 2125 -673 2177
rect -621 2125 -606 2177
rect -554 2125 -539 2177
rect -487 2125 -479 2177
tri -322 2175 -306 2191 se
rect -306 2175 -248 2191
tri -248 2175 -232 2191 nw
tri 656 2178 669 2191 se
rect 669 2178 1938 2191
tri -132 2175 -129 2178 se
rect -129 2175 1938 2178
rect 1990 2175 2002 2227
rect 2054 2175 2060 2227
rect 2140 2196 2146 2248
rect 2198 2196 2212 2248
rect 2264 2196 2270 2248
tri 4764 2224 4788 2248 ne
rect 4788 2224 4837 2248
tri -325 2172 -322 2175 se
rect -322 2172 -251 2175
tri -251 2172 -248 2175 nw
tri -135 2172 -132 2175 se
rect -132 2172 724 2175
tri 724 2172 727 2175 nw
rect 2797 2172 2803 2224
rect 2855 2172 2867 2224
rect 2919 2172 2925 2224
tri 4788 2218 4794 2224 ne
rect 4794 2218 4837 2224
tri 4837 2218 4868 2249 sw
rect 6079 2218 6207 2292
tri 4794 2210 4802 2218 ne
rect 4802 2210 5505 2218
tri -339 2158 -325 2172 se
rect -325 2158 -265 2172
tri -265 2158 -251 2172 nw
tri -149 2158 -135 2172 se
rect -135 2158 710 2172
tri 710 2158 724 2172 nw
tri 2797 2158 2811 2172 ne
rect 2811 2158 2911 2172
tri 2911 2158 2925 2172 nw
rect 3110 2158 3116 2210
rect 3168 2158 3180 2210
rect 3232 2158 3238 2210
tri 4802 2187 4825 2210 ne
rect 4825 2187 5505 2210
tri 4825 2166 4846 2187 ne
rect 4846 2166 5505 2187
rect 5557 2166 5569 2218
rect 5621 2166 5627 2218
rect 6079 2166 6085 2218
rect 6137 2166 6149 2218
rect 6201 2166 6207 2218
rect -812 2122 -479 2125
tri -355 2142 -339 2158 se
rect -339 2142 -281 2158
tri -281 2142 -265 2158 nw
tri -165 2142 -149 2158 se
rect -149 2142 694 2158
tri 694 2142 710 2158 nw
tri 2811 2142 2827 2158 ne
rect 2827 2142 2896 2158
tri 2896 2143 2911 2158 nw
tri 3110 2143 3125 2158 ne
rect 3125 2143 3208 2158
rect -355 2129 -294 2142
tri -294 2129 -281 2142 nw
tri -178 2129 -165 2142 se
rect -165 2129 681 2142
tri 681 2129 694 2142 nw
tri 2827 2129 2840 2142 ne
rect 2840 2129 2896 2142
tri -1218 1956 -1205 1969 sw
rect -1270 1947 -1205 1956
tri -1270 1942 -1265 1947 ne
rect -1265 1942 -1205 1947
tri -1205 1942 -1191 1956 sw
tri -369 1942 -355 1956 se
rect -355 1942 -303 2129
tri -303 2120 -294 2129 nw
tri -182 2125 -178 2129 se
rect -178 2126 678 2129
tri 678 2126 681 2129 nw
rect -178 2125 -108 2126
tri -108 2125 -107 2126 nw
tri -187 2120 -182 2125 se
rect -182 2120 -129 2125
tri -203 2104 -187 2120 se
rect -187 2104 -129 2120
tri -129 2104 -108 2125 nw
tri -215 2092 -203 2104 se
rect -203 2092 -141 2104
tri -141 2092 -129 2104 nw
tri -242 2065 -215 2092 se
rect -215 2065 -168 2092
tri -168 2065 -141 2092 nw
tri -267 2040 -242 2065 se
rect -242 2040 -193 2065
tri -193 2040 -168 2065 nw
rect 440 2040 446 2092
rect 498 2040 510 2092
rect 562 2040 568 2092
rect 765 2077 771 2129
rect 823 2077 837 2129
rect 889 2077 904 2129
rect 1090 2077 1098 2129
rect 1157 2127 1453 2129
rect 1157 2077 1299 2127
tri 916 2075 918 2077 ne
rect 918 2075 929 2077
tri 918 2073 920 2075 ne
rect 920 2073 929 2075
rect 985 2073 1013 2077
rect 1069 2073 1098 2077
rect 1154 2075 1299 2077
rect 1351 2075 1395 2127
rect 1447 2075 1453 2127
tri 2840 2125 2844 2129 ne
rect 1154 2073 1453 2075
tri -1265 1937 -1260 1942 ne
rect -1260 1937 -1191 1942
tri -1191 1937 -1186 1942 sw
tri -374 1937 -369 1942 se
rect -369 1937 -303 1942
tri -1260 1928 -1251 1937 ne
rect -1251 1928 -1186 1937
tri -1186 1928 -1177 1937 sw
tri -383 1928 -374 1937 se
rect -374 1934 -303 1937
rect -374 1928 -309 1934
tri -309 1928 -303 1934 nw
tri -268 2039 -267 2040 se
rect -267 2039 -194 2040
tri -194 2039 -193 2040 nw
tri -1251 1908 -1231 1928 ne
rect -1231 1912 -325 1928
tri -325 1912 -309 1928 nw
rect -1231 1908 -339 1912
tri -1319 1895 -1306 1908 sw
tri -1231 1895 -1218 1908 ne
rect -1218 1898 -339 1908
tri -339 1898 -325 1912 nw
tri -282 1898 -268 1912 se
rect -268 1898 -216 2039
tri -216 2017 -194 2039 nw
rect -1218 1895 -342 1898
tri -342 1895 -339 1898 nw
tri -285 1895 -282 1898 se
rect -282 1895 -216 1898
rect -1371 1886 -1306 1895
tri -1371 1863 -1348 1886 ne
rect -1348 1876 -1306 1886
tri -1306 1876 -1287 1895 sw
tri -1218 1876 -1199 1895 ne
rect -1199 1876 -361 1895
tri -361 1876 -342 1895 nw
tri -304 1876 -285 1895 se
rect -285 1890 -216 1895
rect -285 1876 -243 1890
rect -1348 1863 -1287 1876
tri -1287 1863 -1274 1876 sw
tri -317 1863 -304 1876 se
rect -304 1863 -243 1876
tri -243 1863 -216 1890 nw
rect -176 1942 -170 1994
rect -118 1942 -102 1994
rect -50 1942 -44 1994
tri -1348 1841 -1326 1863 ne
rect -1326 1841 -1274 1863
tri -1274 1841 -1252 1863 sw
tri -339 1841 -317 1863 se
rect -317 1841 -265 1863
tri -265 1841 -243 1863 nw
tri -1326 1834 -1319 1841 ne
rect -1319 1834 -272 1841
tri -272 1834 -265 1841 nw
tri -1319 1811 -1296 1834 ne
rect -1296 1811 -295 1834
tri -295 1811 -272 1834 nw
tri -1296 1799 -1284 1811 ne
rect -1284 1799 -307 1811
tri -307 1799 -295 1811 nw
rect -176 1799 -44 1942
rect 440 1937 568 2040
rect 2476 2059 2528 2065
tri 2455 2007 2476 2028 se
tri 2443 1995 2455 2007 se
rect 2455 1995 2528 2007
tri 2528 1995 2561 2028 sw
tri 2437 1989 2443 1995 se
rect 2443 1989 2476 1995
tri 568 1937 571 1940 sw
rect 1748 1937 1754 1989
rect 1806 1937 1821 1989
rect 1873 1937 1888 1989
rect 1940 1937 1955 1989
rect 2007 1943 2476 1989
rect 2528 1989 2561 1995
tri 2561 1989 2567 1995 sw
rect 2528 1943 2691 1989
rect 2007 1937 2691 1943
rect 2743 1937 2755 1989
rect 2807 1937 2813 1989
rect 440 1869 571 1937
tri 571 1869 639 1937 sw
rect 440 1863 1681 1869
rect 440 1811 1197 1863
rect 1249 1811 1629 1863
tri -44 1799 -38 1805 sw
rect 440 1799 1681 1811
tri -1284 1789 -1274 1799 ne
rect -1274 1789 -317 1799
tri -317 1789 -307 1799 nw
rect -176 1789 -38 1799
tri -38 1789 -28 1799 sw
rect -176 1747 -28 1789
tri -28 1747 14 1789 sw
rect 440 1747 1197 1799
rect 1249 1747 1629 1799
rect -176 1741 14 1747
tri 14 1741 20 1747 sw
rect 440 1741 1681 1747
rect 2844 1836 2896 2129
tri 3125 2112 3156 2143 ne
rect 2844 1772 2896 1784
rect -176 1720 20 1741
tri 20 1720 41 1741 sw
rect -176 1714 41 1720
tri 41 1714 47 1720 sw
rect 2844 1714 2896 1720
rect 3156 1836 3208 2143
tri 3208 2128 3238 2158 nw
rect 3243 1943 3249 1995
rect 3301 1943 3313 1995
rect 3365 1943 4228 1995
rect 4280 1943 4292 1995
rect 4344 1943 4350 1995
rect 3156 1772 3208 1784
rect 3156 1714 3208 1720
rect 3879 1836 3931 1842
rect 3879 1772 3931 1784
rect 3879 1714 3931 1720
rect -176 1699 47 1714
tri 47 1699 62 1714 sw
tri -837 1647 -785 1699 se
rect -785 1647 -716 1699
rect -664 1647 -650 1699
rect -598 1647 -592 1699
rect -176 1693 2441 1699
tri -843 1641 -837 1647 se
rect -837 1641 -769 1647
tri -769 1641 -763 1647 nw
rect -176 1641 333 1693
rect 385 1663 1964 1693
rect 385 1641 1294 1663
tri -855 1629 -843 1641 se
rect -843 1629 -781 1641
tri -781 1629 -769 1641 nw
rect -176 1629 1294 1641
tri -859 1625 -855 1629 se
rect -855 1625 -785 1629
tri -785 1625 -781 1629 nw
tri -876 1608 -859 1625 se
rect -859 1608 -802 1625
tri -802 1608 -785 1625 nw
rect -176 1618 333 1629
tri -176 1608 -166 1618 ne
rect -166 1608 333 1618
rect -876 971 -824 1608
tri -824 1586 -802 1608 nw
tri -166 1586 -144 1608 ne
rect -144 1586 333 1608
tri -144 1577 -135 1586 ne
rect -135 1577 333 1586
rect 385 1607 1294 1629
rect 1350 1607 1374 1663
rect 1430 1641 1964 1663
rect 2016 1672 2441 1693
tri 2441 1672 2468 1699 sw
rect 2016 1666 2468 1672
tri 2468 1666 2474 1672 sw
tri 3391 1666 3397 1672 se
rect 3397 1666 4341 1672
rect 2016 1641 2474 1666
rect 1430 1629 2474 1641
rect 1430 1607 1964 1629
rect 385 1577 1964 1607
rect 2016 1614 2474 1629
tri 2474 1614 2526 1666 sw
tri 3339 1614 3391 1666 se
rect 3391 1614 4289 1666
rect 2016 1602 4341 1614
rect 2016 1577 4289 1602
tri -135 1571 -129 1577 ne
rect -129 1571 4289 1577
tri 2387 1550 2408 1571 ne
rect 2408 1550 4289 1571
tri 2408 1544 2414 1550 ne
rect 2414 1544 4341 1550
tri 2414 1524 2434 1544 ne
rect 2434 1524 3393 1544
rect -230 1518 1897 1524
rect -178 1466 117 1518
rect 169 1466 549 1518
rect 601 1466 981 1518
rect 1033 1466 1413 1518
rect 1465 1466 1845 1518
tri 2434 1486 2472 1524 ne
rect 2472 1486 3393 1524
tri 3393 1486 3451 1544 nw
rect -230 1454 1897 1466
rect -734 1400 -440 1424
rect -734 1348 -725 1400
rect -673 1348 -650 1400
rect -598 1348 -574 1400
rect -522 1348 -498 1400
rect -446 1348 -440 1400
rect -178 1402 117 1454
rect 169 1402 549 1454
rect 601 1402 981 1454
rect 1033 1402 1413 1454
rect 1465 1402 1845 1454
rect -230 1396 1897 1402
rect -734 1235 -440 1348
rect -310 1299 -256 1305
rect -258 1247 -256 1299
tri -440 1235 -429 1246 sw
rect -310 1235 -256 1247
rect -734 1183 -429 1235
tri -429 1183 -377 1235 sw
rect -258 1229 -256 1235
tri -256 1229 -180 1305 sw
rect -258 1183 3807 1229
rect -734 1177 -377 1183
tri -377 1177 -371 1183 sw
rect -310 1177 3807 1183
rect 3859 1177 3871 1229
rect 3923 1177 3929 1229
rect -734 1083 -371 1177
tri -371 1083 -277 1177 sw
rect -734 1077 4200 1083
rect -734 1032 765 1077
tri -734 1025 -727 1032 ne
rect -727 1025 765 1032
rect 817 1068 2122 1077
rect 817 1025 930 1068
tri -727 1020 -722 1025 ne
rect -722 1020 930 1025
tri -722 1013 -715 1020 ne
rect -715 1013 930 1020
tri -715 993 -695 1013 ne
rect -695 993 765 1013
tri -824 971 -802 993 sw
tri -695 971 -673 993 ne
rect -673 971 765 993
tri -876 961 -866 971 ne
rect -866 961 -802 971
tri -802 961 -792 971 sw
tri -673 961 -663 971 ne
rect -663 961 765 971
rect 817 1012 930 1013
rect 986 1012 1014 1068
rect 1070 1012 1098 1068
rect 1154 1025 2122 1068
rect 2174 1025 2404 1077
rect 2456 1025 2688 1077
rect 2740 1025 3000 1077
rect 3052 1025 3315 1077
rect 3367 1025 3436 1077
rect 3488 1072 4200 1077
rect 3488 1025 3709 1072
rect 1154 1020 3709 1025
rect 3761 1020 3793 1072
rect 3845 1020 3877 1072
rect 3929 1020 4200 1072
rect 1154 1013 4200 1020
rect 1154 1012 2122 1013
rect 817 962 2122 1012
rect 817 961 930 962
tri -866 949 -854 961 ne
rect -854 949 -792 961
tri -792 949 -780 961 sw
tri -663 949 -651 961 ne
rect -651 949 930 961
tri -854 897 -802 949 ne
rect -802 897 -780 949
tri -780 897 -728 949 sw
tri -651 897 -599 949 ne
rect -599 897 765 949
rect 817 906 930 949
rect 986 906 1014 962
rect 1070 906 1098 962
rect 1154 961 2122 962
rect 2174 961 2404 1013
rect 2456 961 2688 1013
rect 2740 961 3000 1013
rect 3052 961 3315 1013
rect 3367 1001 4200 1013
rect 3367 961 3436 1001
rect 1154 949 3436 961
rect 3488 1000 4200 1001
rect 3488 949 3709 1000
rect 1154 906 2122 949
rect 817 897 2122 906
rect 2174 897 2404 949
rect 2456 897 2688 949
rect 2740 897 3000 949
rect 3052 897 3315 949
rect 3367 948 3709 949
rect 3761 948 3793 1000
rect 3845 948 3877 1000
rect 3929 948 4200 1000
rect 3367 928 4200 948
rect 3367 924 3709 928
rect 3367 897 3436 924
tri -802 891 -796 897 ne
rect -796 891 -728 897
tri -728 891 -722 897 sw
tri -599 891 -593 897 ne
rect -593 891 3436 897
tri -796 872 -777 891 ne
rect -777 872 -722 891
tri -722 872 -703 891 sw
tri -593 872 -574 891 ne
rect -574 872 3436 891
rect 3488 876 3709 924
rect 3761 876 3793 928
rect 3845 876 3877 928
rect 3929 876 4200 928
rect 3488 872 4200 876
tri -777 856 -761 872 ne
rect -761 856 -703 872
tri -703 856 -687 872 sw
tri -574 856 -558 872 ne
rect -558 857 4200 872
rect -558 856 930 857
tri -761 847 -752 856 ne
rect -752 847 -687 856
tri -687 847 -678 856 sw
tri -558 847 -549 856 ne
rect -549 847 930 856
tri -752 841 -746 847 ne
rect -746 841 -678 847
tri -678 841 -672 847 sw
tri -549 841 -543 847 ne
rect -543 841 930 847
rect 986 841 1014 857
rect 1070 841 1098 857
rect 1154 856 4200 857
rect 1154 847 3709 856
rect 1154 841 3436 847
tri -746 823 -728 841 ne
rect -728 823 -672 841
tri -672 823 -654 841 sw
tri -543 823 -525 841 ne
rect -525 823 169 841
tri -728 789 -694 823 ne
rect -694 789 -654 823
tri -654 789 -620 823 sw
tri -525 789 -491 823 ne
rect -491 789 169 823
rect 221 789 234 841
rect 286 789 299 841
rect 351 789 363 841
rect 415 789 427 841
rect 479 789 491 841
rect 543 789 555 841
rect 607 789 619 841
rect 671 789 683 841
rect 735 789 747 841
rect 799 789 811 841
rect 863 789 875 841
rect 927 801 930 841
rect 927 789 939 801
rect 991 789 1003 841
rect 1055 789 1067 801
rect 1119 789 1131 801
rect 1183 789 1195 841
rect 1247 789 1259 841
rect 1311 789 1323 841
rect 1375 789 1387 841
rect 1439 789 1451 841
rect 1503 789 1515 841
rect 1567 789 1579 841
rect 1631 789 1643 841
rect 1695 789 1707 841
rect 1759 789 1771 841
rect 1823 789 1835 841
rect 1887 789 1899 841
rect 1951 789 1963 841
rect 2015 789 2027 841
rect 2079 789 2091 841
rect 2143 789 2155 841
rect 2207 789 2219 841
rect 2271 789 2283 841
rect 2335 789 2347 841
rect 2399 789 2411 841
rect 2463 789 2475 841
rect 2527 789 2539 841
rect 2591 789 2603 841
rect 2655 789 2667 841
rect 2719 789 2731 841
rect 2783 789 2795 841
rect 2847 789 2859 841
rect 2911 789 2923 841
rect 2975 789 2987 841
rect 3039 789 3051 841
rect 3103 789 3115 841
rect 3167 789 3179 841
rect 3231 789 3243 841
rect 3295 789 3307 841
rect 3359 795 3436 841
rect 3488 804 3709 847
rect 3761 804 3793 856
rect 3845 804 3877 856
rect 3929 804 4200 856
rect 3488 795 4200 804
rect 3359 789 4200 795
tri -694 749 -654 789 ne
rect -654 749 -620 789
tri -620 749 -580 789 sw
tri 82 749 122 789 ne
rect 122 749 733 789
tri -654 722 -627 749 ne
rect -627 722 -580 749
tri -580 722 -553 749 sw
tri 122 722 149 749 ne
rect 149 722 733 749
tri 733 722 800 789 nw
tri -627 716 -621 722 ne
rect -621 716 -553 722
tri -553 716 -547 722 sw
tri 149 716 155 722 ne
rect 155 716 727 722
tri 727 716 733 722 nw
rect 2687 716 3052 789
tri -621 680 -585 716 ne
rect -585 680 -547 716
tri -547 680 -511 716 sw
tri 155 680 191 716 ne
rect 191 680 691 716
tri 691 680 727 716 nw
tri -585 675 -580 680 ne
rect -580 675 -511 680
tri -511 675 -506 680 sw
tri 191 675 196 680 ne
rect 196 675 640 680
tri -580 629 -534 675 ne
rect -534 629 -506 675
tri -506 629 -460 675 sw
tri 196 629 242 675 ne
rect 242 629 640 675
tri 640 629 691 680 nw
tri -534 628 -533 629 ne
rect -533 628 -460 629
tri -460 628 -459 629 sw
rect 242 628 639 629
tri 639 628 640 629 nw
rect 1285 628 1291 680
rect 1350 628 1372 680
tri -533 601 -506 628 ne
rect -506 601 -459 628
tri -459 601 -432 628 sw
tri -506 600 -505 601 ne
rect -505 600 -432 601
tri -432 600 -431 601 sw
rect 242 600 611 628
tri 611 600 639 628 nw
rect 1285 624 1294 628
rect 1350 624 1374 628
rect 1430 624 1439 680
rect 2739 664 3000 716
rect 2687 652 3052 664
rect 2739 600 3000 652
tri -505 567 -472 600 ne
rect -472 567 -431 600
tri -431 567 -398 600 sw
rect 242 594 605 600
tri 605 594 611 600 nw
rect 2687 594 3052 600
tri -472 527 -432 567 ne
rect -432 527 66 567
tri -432 515 -420 527 ne
rect -420 515 66 527
rect 118 515 130 567
rect 182 515 188 567
rect 242 543 554 594
tri 554 543 605 594 nw
rect -32350 501 -27106 504
rect -32350 449 -32338 501
rect -32286 449 -32273 501
rect -32221 449 -32208 501
rect -32156 449 -32143 501
rect -32091 449 -32078 501
rect -32026 449 -32013 501
rect -31961 449 -31948 501
rect -31896 449 -31882 501
rect -31830 449 -31816 501
rect -31764 495 -27106 501
rect -31764 449 -29135 495
rect -32350 443 -29135 449
rect -29083 443 -29053 495
rect -29001 443 -28971 495
rect -28919 443 -28889 495
rect -28837 488 -27106 495
rect -28837 443 -28188 488
rect -32350 437 -28188 443
rect -32350 385 -32338 437
rect -32286 385 -32273 437
rect -32221 385 -32208 437
rect -32156 385 -32143 437
rect -32091 385 -32078 437
rect -32026 385 -32013 437
rect -31961 385 -31948 437
rect -31896 385 -31882 437
rect -31830 385 -31816 437
rect -31764 436 -28188 437
rect -28136 436 -28122 488
rect -28070 436 -28056 488
rect -28004 436 -27990 488
rect -27938 436 -27924 488
rect -27872 436 -27858 488
rect -27806 436 -27792 488
rect -27740 436 -27726 488
rect -27674 436 -27659 488
rect -27607 436 -27592 488
rect -27540 436 -27525 488
rect -27473 436 -27458 488
rect -27406 436 -27391 488
rect -27339 436 -27324 488
rect -27272 436 -27257 488
rect -27205 436 -27190 488
rect -27138 436 -27106 488
rect -31764 430 -27106 436
rect -31764 385 -29135 430
rect -32350 378 -29135 385
rect -29083 378 -29053 430
rect -29001 378 -28971 430
rect -28919 378 -28889 430
rect -28837 420 -27106 430
rect -28837 378 -28188 420
rect -32350 373 -28188 378
rect -32350 321 -32338 373
rect -32286 321 -32273 373
rect -32221 321 -32208 373
rect -32156 321 -32143 373
rect -32091 321 -32078 373
rect -32026 321 -32013 373
rect -31961 321 -31948 373
rect -31896 321 -31882 373
rect -31830 321 -31816 373
rect -31764 368 -28188 373
rect -28136 368 -28122 420
rect -28070 368 -28056 420
rect -28004 368 -27990 420
rect -27938 368 -27924 420
rect -27872 368 -27858 420
rect -27806 368 -27792 420
rect -27740 368 -27726 420
rect -27674 368 -27659 420
rect -27607 368 -27592 420
rect -27540 368 -27525 420
rect -27473 368 -27458 420
rect -27406 368 -27391 420
rect -27339 368 -27324 420
rect -27272 368 -27257 420
rect -27205 368 -27190 420
rect -27138 368 -27106 420
rect -31764 365 -27106 368
rect -31764 321 -29135 365
rect -32350 313 -29135 321
rect -29083 313 -29053 365
rect -29001 313 -28971 365
rect -28919 313 -28889 365
rect -28837 352 -27106 365
rect -28837 313 -28188 352
rect -32350 309 -28188 313
rect -32350 257 -32338 309
rect -32286 257 -32273 309
rect -32221 257 -32208 309
rect -32156 257 -32143 309
rect -32091 257 -32078 309
rect -32026 257 -32013 309
rect -31961 257 -31948 309
rect -31896 257 -31882 309
rect -31830 257 -31816 309
rect -31764 301 -28188 309
rect -31764 257 -29135 301
rect -32350 249 -29135 257
rect -29083 249 -29053 301
rect -29001 249 -28971 301
rect -28919 249 -28889 301
rect -28837 300 -28188 301
rect -28136 300 -28122 352
rect -28070 300 -28056 352
rect -28004 300 -27990 352
rect -27938 300 -27924 352
rect -27872 300 -27858 352
rect -27806 300 -27792 352
rect -27740 300 -27726 352
rect -27674 300 -27659 352
rect -27607 300 -27592 352
rect -27540 300 -27525 352
rect -27473 300 -27458 352
rect -27406 300 -27391 352
rect -27339 300 -27324 352
rect -27272 300 -27257 352
rect -27205 300 -27190 352
rect -27138 300 -27106 352
rect -28837 284 -27106 300
rect -28837 249 -28188 284
rect -32350 245 -28188 249
rect -32350 193 -32338 245
rect -32286 193 -32273 245
rect -32221 193 -32208 245
rect -32156 193 -32143 245
rect -32091 193 -32078 245
rect -32026 193 -32013 245
rect -31961 193 -31948 245
rect -31896 193 -31882 245
rect -31830 193 -31816 245
rect -31764 237 -28188 245
rect -31764 193 -29135 237
rect -32350 185 -29135 193
rect -29083 185 -29053 237
rect -29001 185 -28971 237
rect -28919 185 -28889 237
rect -28837 232 -28188 237
rect -28136 232 -28122 284
rect -28070 232 -28056 284
rect -28004 232 -27990 284
rect -27938 232 -27924 284
rect -27872 232 -27858 284
rect -27806 232 -27792 284
rect -27740 232 -27726 284
rect -27674 232 -27659 284
rect -27607 232 -27592 284
rect -27540 232 -27525 284
rect -27473 232 -27458 284
rect -27406 232 -27391 284
rect -27339 232 -27324 284
rect -27272 232 -27257 284
rect -27205 232 -27190 284
rect -27138 232 -27106 284
rect -28837 216 -27106 232
rect -28837 185 -28188 216
rect -32350 181 -28188 185
rect -32350 129 -32338 181
rect -32286 129 -32273 181
rect -32221 129 -32208 181
rect -32156 129 -32143 181
rect -32091 129 -32078 181
rect -32026 129 -32013 181
rect -31961 129 -31948 181
rect -31896 129 -31882 181
rect -31830 129 -31816 181
rect -31764 173 -28188 181
rect -31764 129 -29135 173
rect -32350 121 -29135 129
rect -29083 121 -29053 173
rect -29001 121 -28971 173
rect -28919 121 -28889 173
rect -28837 164 -28188 173
rect -28136 164 -28122 216
rect -28070 164 -28056 216
rect -28004 164 -27990 216
rect -27938 164 -27924 216
rect -27872 164 -27858 216
rect -27806 164 -27792 216
rect -27740 164 -27726 216
rect -27674 164 -27659 216
rect -27607 164 -27592 216
rect -27540 164 -27525 216
rect -27473 164 -27458 216
rect -27406 164 -27391 216
rect -27339 164 -27324 216
rect -27272 164 -27257 216
rect -27205 164 -27190 216
rect -27138 164 -27106 216
rect -28837 148 -27106 164
rect -28837 121 -28188 148
rect -32350 117 -28188 121
rect -32350 65 -32338 117
rect -32286 65 -32273 117
rect -32221 65 -32208 117
rect -32156 65 -32143 117
rect -32091 65 -32078 117
rect -32026 65 -32013 117
rect -31961 65 -31948 117
rect -31896 65 -31882 117
rect -31830 65 -31816 117
rect -31764 109 -28188 117
rect -31764 65 -29135 109
rect -32350 57 -29135 65
rect -29083 57 -29053 109
rect -29001 57 -28971 109
rect -28919 57 -28889 109
rect -28837 96 -28188 109
rect -28136 96 -28122 148
rect -28070 96 -28056 148
rect -28004 96 -27990 148
rect -27938 96 -27924 148
rect -27872 96 -27858 148
rect -27806 96 -27792 148
rect -27740 96 -27726 148
rect -27674 96 -27659 148
rect -27607 96 -27592 148
rect -27540 96 -27525 148
rect -27473 96 -27458 148
rect -27406 96 -27391 148
rect -27339 96 -27324 148
rect -27272 96 -27257 148
rect -27205 96 -27190 148
rect -27138 96 -27106 148
rect -28837 80 -27106 96
rect -28837 57 -28188 80
rect -32350 53 -28188 57
rect -32350 1 -32338 53
rect -32286 1 -32273 53
rect -32221 1 -32208 53
rect -32156 1 -32143 53
rect -32091 1 -32078 53
rect -32026 1 -32013 53
rect -31961 1 -31948 53
rect -31896 1 -31882 53
rect -31830 1 -31816 53
rect -31764 45 -28188 53
rect -31764 1 -29135 45
rect -32350 -7 -29135 1
rect -29083 -7 -29053 45
rect -29001 -7 -28971 45
rect -28919 -7 -28889 45
rect -28837 28 -28188 45
rect -28136 28 -28122 80
rect -28070 28 -28056 80
rect -28004 28 -27990 80
rect -27938 28 -27924 80
rect -27872 28 -27858 80
rect -27806 28 -27792 80
rect -27740 28 -27726 80
rect -27674 28 -27659 80
rect -27607 28 -27592 80
rect -27540 28 -27525 80
rect -27473 28 -27458 80
rect -27406 28 -27391 80
rect -27339 28 -27324 80
rect -27272 28 -27257 80
rect -27205 28 -27190 80
rect -27138 28 -27106 80
rect 242 320 546 543
tri 546 535 554 543 nw
rect 2807 535 2924 543
rect 2807 483 2813 535
rect 2865 483 2877 535
rect 2980 487 3004 543
rect 3060 535 3265 543
rect 3060 487 3143 535
rect 2929 483 3143 487
rect 3195 483 3207 535
rect 3259 483 3265 535
rect 242 268 248 320
rect 300 268 328 320
rect 380 268 408 320
rect 460 268 488 320
rect 540 268 546 320
rect 242 191 546 268
rect 242 139 248 191
rect 300 139 328 191
rect 380 139 408 191
rect 460 139 488 191
rect 540 139 546 191
rect 242 84 546 139
rect 242 32 248 84
rect 300 32 328 84
rect 380 32 408 84
rect 460 32 488 84
rect 540 32 546 84
rect -28837 12 -27106 28
rect -28837 -7 -28188 12
rect -32350 -11 -28188 -7
rect -32350 -63 -32338 -11
rect -32286 -63 -32273 -11
rect -32221 -63 -32208 -11
rect -32156 -63 -32143 -11
rect -32091 -63 -32078 -11
rect -32026 -63 -32013 -11
rect -31961 -63 -31948 -11
rect -31896 -63 -31882 -11
rect -31830 -63 -31816 -11
rect -31764 -19 -28188 -11
rect -31764 -63 -29135 -19
rect -32350 -71 -29135 -63
rect -29083 -71 -29053 -19
rect -29001 -71 -28971 -19
rect -28919 -71 -28889 -19
rect -28837 -40 -28188 -19
rect -28136 -40 -28122 12
rect -28070 -40 -28056 12
rect -28004 -40 -27990 12
rect -27938 -40 -27924 12
rect -27872 -40 -27858 12
rect -27806 -40 -27792 12
rect -27740 -40 -27726 12
rect -27674 -40 -27659 12
rect -27607 -40 -27592 12
rect -27540 -40 -27525 12
rect -27473 -40 -27458 12
rect -27406 -40 -27391 12
rect -27339 -40 -27324 12
rect -27272 -40 -27257 12
rect -27205 -40 -27190 12
rect -27138 -40 -27106 12
rect -28837 -56 -27106 -40
rect -28837 -71 -28188 -56
rect -32350 -75 -28188 -71
rect -32350 -127 -32338 -75
rect -32286 -127 -32273 -75
rect -32221 -127 -32208 -75
rect -32156 -127 -32143 -75
rect -32091 -127 -32078 -75
rect -32026 -127 -32013 -75
rect -31961 -127 -31948 -75
rect -31896 -127 -31882 -75
rect -31830 -127 -31816 -75
rect -31764 -83 -28188 -75
rect -31764 -127 -29135 -83
rect -32350 -135 -29135 -127
rect -29083 -135 -29053 -83
rect -29001 -135 -28971 -83
rect -28919 -135 -28889 -83
rect -28837 -108 -28188 -83
rect -28136 -108 -28122 -56
rect -28070 -108 -28056 -56
rect -28004 -108 -27990 -56
rect -27938 -108 -27924 -56
rect -27872 -108 -27858 -56
rect -27806 -108 -27792 -56
rect -27740 -108 -27726 -56
rect -27674 -108 -27659 -56
rect -27607 -108 -27592 -56
rect -27540 -108 -27525 -56
rect -27473 -108 -27458 -56
rect -27406 -108 -27391 -56
rect -27339 -108 -27324 -56
rect -27272 -108 -27257 -56
rect -27205 -108 -27190 -56
rect -27138 -108 -27106 -56
rect -28837 -124 -27106 -108
rect -28837 -135 -28188 -124
rect -32350 -139 -28188 -135
rect -32350 -191 -32338 -139
rect -32286 -191 -32273 -139
rect -32221 -191 -32208 -139
rect -32156 -191 -32143 -139
rect -32091 -191 -32078 -139
rect -32026 -191 -32013 -139
rect -31961 -191 -31948 -139
rect -31896 -191 -31882 -139
rect -31830 -191 -31816 -139
rect -31764 -147 -28188 -139
rect -31764 -191 -29135 -147
rect -32350 -199 -29135 -191
rect -29083 -199 -29053 -147
rect -29001 -199 -28971 -147
rect -28919 -199 -28889 -147
rect -28837 -176 -28188 -147
rect -28136 -176 -28122 -124
rect -28070 -176 -28056 -124
rect -28004 -176 -27990 -124
rect -27938 -176 -27924 -124
rect -27872 -176 -27858 -124
rect -27806 -176 -27792 -124
rect -27740 -176 -27726 -124
rect -27674 -176 -27659 -124
rect -27607 -176 -27592 -124
rect -27540 -176 -27525 -124
rect -27473 -176 -27458 -124
rect -27406 -176 -27391 -124
rect -27339 -176 -27324 -124
rect -27272 -176 -27257 -124
rect -27205 -176 -27190 -124
rect -27138 -176 -27106 -124
rect -28837 -192 -27106 -176
rect -28837 -199 -28188 -192
rect -32350 -203 -28188 -199
rect -32350 -255 -32338 -203
rect -32286 -255 -32273 -203
rect -32221 -255 -32208 -203
rect -32156 -255 -32143 -203
rect -32091 -255 -32078 -203
rect -32026 -255 -32013 -203
rect -31961 -255 -31948 -203
rect -31896 -255 -31882 -203
rect -31830 -255 -31816 -203
rect -31764 -211 -28188 -203
rect -31764 -255 -29135 -211
rect -32350 -263 -29135 -255
rect -29083 -263 -29053 -211
rect -29001 -263 -28971 -211
rect -28919 -263 -28889 -211
rect -28837 -244 -28188 -211
rect -28136 -244 -28122 -192
rect -28070 -244 -28056 -192
rect -28004 -244 -27990 -192
rect -27938 -244 -27924 -192
rect -27872 -244 -27858 -192
rect -27806 -244 -27792 -192
rect -27740 -244 -27726 -192
rect -27674 -244 -27659 -192
rect -27607 -244 -27592 -192
rect -27540 -244 -27525 -192
rect -27473 -244 -27458 -192
rect -27406 -244 -27391 -192
rect -27339 -244 -27324 -192
rect -27272 -244 -27257 -192
rect -27205 -244 -27190 -192
rect -27138 -244 -27106 -192
rect -28837 -260 -27106 -244
rect -28837 -263 -28188 -260
rect -32350 -267 -28188 -263
rect -32350 -319 -32338 -267
rect -32286 -319 -32273 -267
rect -32221 -319 -32208 -267
rect -32156 -319 -32143 -267
rect -32091 -319 -32078 -267
rect -32026 -319 -32013 -267
rect -31961 -319 -31948 -267
rect -31896 -319 -31882 -267
rect -31830 -319 -31816 -267
rect -31764 -275 -28188 -267
rect -31764 -319 -29135 -275
rect -32350 -327 -29135 -319
rect -29083 -327 -29053 -275
rect -29001 -327 -28971 -275
rect -28919 -327 -28889 -275
rect -28837 -312 -28188 -275
rect -28136 -312 -28122 -260
rect -28070 -312 -28056 -260
rect -28004 -312 -27990 -260
rect -27938 -312 -27924 -260
rect -27872 -312 -27858 -260
rect -27806 -312 -27792 -260
rect -27740 -312 -27726 -260
rect -27674 -312 -27659 -260
rect -27607 -312 -27592 -260
rect -27540 -312 -27525 -260
rect -27473 -312 -27458 -260
rect -27406 -312 -27391 -260
rect -27339 -312 -27324 -260
rect -27272 -312 -27257 -260
rect -27205 -312 -27190 -260
rect -27138 -312 -27106 -260
rect -28837 -327 -27106 -312
rect -32350 -328 -27106 -327
rect -32350 -331 -28188 -328
rect -32350 -383 -32338 -331
rect -32286 -383 -32273 -331
rect -32221 -383 -32208 -331
rect -32156 -383 -32143 -331
rect -32091 -383 -32078 -331
rect -32026 -383 -32013 -331
rect -31961 -383 -31948 -331
rect -31896 -383 -31882 -331
rect -31830 -383 -31816 -331
rect -31764 -339 -28188 -331
rect -31764 -383 -29135 -339
rect -32350 -391 -29135 -383
rect -29083 -391 -29053 -339
rect -29001 -391 -28971 -339
rect -28919 -391 -28889 -339
rect -28837 -380 -28188 -339
rect -28136 -380 -28122 -328
rect -28070 -380 -28056 -328
rect -28004 -380 -27990 -328
rect -27938 -380 -27924 -328
rect -27872 -380 -27858 -328
rect -27806 -380 -27792 -328
rect -27740 -380 -27726 -328
rect -27674 -380 -27659 -328
rect -27607 -380 -27592 -328
rect -27540 -380 -27525 -328
rect -27473 -380 -27458 -328
rect -27406 -380 -27391 -328
rect -27339 -380 -27324 -328
rect -27272 -380 -27257 -328
rect -27205 -380 -27190 -328
rect -27138 -380 -27106 -328
rect -28837 -391 -27106 -380
rect -32350 -402 -27106 -391
tri 1495 -1856 1499 -1852 se
rect 1499 -1856 1508 -1852
rect -10881 -1908 1508 -1856
rect 1564 -1908 1588 -1852
rect 1644 -1908 1653 -1852
rect -29280 -8589 -29228 -8583
rect -31521 -8625 -31469 -8619
rect -31521 -8689 -31469 -8677
tri -31545 -9890 -31521 -9866 se
rect -31521 -9890 -31469 -8741
rect -29280 -8653 -29228 -8641
tri -29342 -9754 -29280 -9692 se
rect -29280 -9754 -29228 -8705
rect -10881 -9678 -10727 -1908
tri -10727 -1951 -10684 -1908 nw
tri 1741 -1945 1745 -1941 se
rect 1745 -1945 1754 -1941
tri -10596 -1951 -10590 -1945 se
rect -10590 -1951 1754 -1945
rect -10881 -9734 -10872 -9678
rect -10816 -9734 -10792 -9678
rect -10736 -9734 -10727 -9678
tri -10647 -2002 -10596 -1951 se
rect -10596 -1997 1754 -1951
rect 1810 -1997 1834 -1941
rect 1890 -1997 1899 -1941
rect -10596 -2002 -10403 -1997
tri -10403 -2002 -10398 -1997 nw
rect -10647 -9678 -10493 -2002
tri -10493 -2092 -10403 -2002 nw
rect -10647 -9734 -10638 -9678
rect -10582 -9734 -10558 -9678
rect -10502 -9734 -10493 -9678
tri -29358 -9770 -29342 -9754 se
rect -29342 -9770 -29228 -9754
tri -29228 -9770 -29212 -9754 sw
rect -29366 -9826 -29357 -9770
rect -29301 -9826 -29277 -9770
rect -29221 -9826 -29212 -9770
tri -31469 -9890 -31442 -9863 sw
rect -31545 -9946 -31536 -9890
rect -31480 -9946 -31456 -9890
rect -31400 -9946 -31391 -9890
<< via2 >>
rect 1754 3189 1810 3245
rect 1834 3189 1890 3245
rect 2924 3145 2980 3201
rect 3004 3145 3060 3201
rect 1508 3003 1564 3059
rect 1588 3003 1644 3059
rect 929 2077 956 2129
rect 956 2077 971 2129
rect 971 2077 985 2129
rect 1013 2077 1023 2129
rect 1023 2077 1038 2129
rect 1038 2077 1069 2129
rect 1098 2077 1105 2129
rect 1105 2077 1154 2129
rect 929 2073 985 2077
rect 1013 2073 1069 2077
rect 1098 2073 1154 2077
rect 1294 1607 1350 1663
rect 1374 1607 1430 1663
rect 930 1012 986 1068
rect 1014 1012 1070 1068
rect 1098 1012 1154 1068
rect 930 906 986 962
rect 1014 906 1070 962
rect 1098 906 1154 962
rect 930 841 986 857
rect 1014 841 1070 857
rect 1098 841 1154 857
rect 930 801 939 841
rect 939 801 986 841
rect 1014 801 1055 841
rect 1055 801 1067 841
rect 1067 801 1070 841
rect 1098 801 1119 841
rect 1119 801 1131 841
rect 1131 801 1154 841
rect 1294 628 1343 680
rect 1343 628 1350 680
rect 1374 628 1424 680
rect 1424 628 1430 680
rect 1294 624 1350 628
rect 1374 624 1430 628
rect 2924 535 2980 543
rect 2924 487 2929 535
rect 2929 487 2980 535
rect 3004 487 3060 543
rect 1508 -1908 1564 -1852
rect 1588 -1908 1644 -1852
rect -10872 -9734 -10816 -9678
rect -10792 -9734 -10736 -9678
rect 1754 -1997 1810 -1941
rect 1834 -1997 1890 -1941
rect -10638 -9734 -10582 -9678
rect -10558 -9734 -10502 -9678
rect -29357 -9826 -29301 -9770
rect -29277 -9826 -29221 -9770
rect -31536 -9946 -31480 -9890
rect -31456 -9946 -31400 -9890
<< metal3 >>
rect 1749 3245 1895 3286
rect 1749 3189 1754 3245
rect 1810 3189 1834 3245
rect 1890 3189 1895 3245
rect 1503 3059 1649 3100
rect 1503 3003 1508 3059
rect 1564 3003 1588 3059
rect 1644 3003 1649 3059
rect 924 2129 1159 2134
rect 924 2073 929 2129
rect 985 2073 1013 2129
rect 1069 2073 1098 2129
rect 1154 2073 1159 2129
rect 924 1068 1159 2073
rect 1289 1663 1435 1704
rect 1289 1607 1294 1663
rect 1350 1607 1374 1663
rect 1430 1607 1435 1663
rect 1289 1566 1435 1607
rect 924 1012 930 1068
rect 986 1012 1014 1068
rect 1070 1012 1098 1068
rect 1154 1012 1159 1068
rect 924 962 1159 1012
rect 924 906 930 962
rect 986 906 1014 962
rect 1070 906 1098 962
rect 1154 906 1159 962
rect 924 857 1159 906
rect 924 801 930 857
rect 986 801 1014 857
rect 1070 801 1098 857
rect 1154 801 1159 857
rect 924 795 1159 801
rect 1289 680 1435 751
rect 1289 624 1294 680
rect 1350 624 1374 680
rect 1430 624 1435 680
rect 1289 619 1435 624
rect 1503 -1852 1649 3003
rect 1503 -1908 1508 -1852
rect 1564 -1908 1588 -1852
rect 1644 -1908 1649 -1852
rect 1503 -1913 1649 -1908
rect 1749 -1941 1895 3189
rect 2919 3201 3065 3234
rect 2919 3145 2924 3201
rect 2980 3145 3004 3201
rect 3060 3145 3065 3201
rect 2919 543 3065 3145
rect 2919 487 2924 543
rect 2980 487 3004 543
rect 3060 487 3065 543
rect 2919 482 3065 487
rect 1749 -1997 1754 -1941
rect 1810 -1997 1834 -1941
rect 1890 -1997 1895 -1941
rect 1749 -2002 1895 -1997
tri -10882 -9678 -10877 -9673 se
rect -10877 -9678 -10731 -9673
tri -10938 -9734 -10882 -9678 se
rect -10882 -9734 -10872 -9678
rect -10816 -9734 -10792 -9678
rect -10736 -9734 -10731 -9678
tri -10969 -9765 -10938 -9734 se
rect -10938 -9765 -10731 -9734
rect -29362 -9770 -29216 -9765
rect -29362 -9826 -29357 -9770
rect -29301 -9826 -29277 -9770
rect -29221 -9771 -29216 -9770
tri -29216 -9771 -29210 -9765 sw
tri -10975 -9771 -10969 -9765 se
rect -10969 -9771 -10731 -9765
rect -29221 -9787 -10731 -9771
rect -29221 -9826 -10775 -9787
rect -29362 -9831 -10775 -9826
tri -10775 -9831 -10731 -9787 nw
rect -10643 -9678 -10497 -9673
rect -10643 -9734 -10638 -9678
rect -10582 -9734 -10558 -9678
rect -10502 -9734 -10497 -9678
tri -10663 -9831 -10643 -9811 se
rect -10643 -9831 -10497 -9734
tri -10717 -9885 -10663 -9831 se
rect -10663 -9885 -10497 -9831
rect -31541 -9890 -31395 -9885
rect -31541 -9946 -31536 -9890
rect -31480 -9946 -31456 -9890
rect -31400 -9891 -31395 -9890
tri -31395 -9891 -31389 -9885 sw
tri -10723 -9891 -10717 -9885 se
rect -10717 -9891 -10497 -9885
rect -31400 -9946 -10497 -9891
rect -31541 -9951 -10497 -9946
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_0
timestamp 1701704242
transform 0 1 5708 -1 0 2914
box 107 226 240 873
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_0
timestamp 1701704242
transform 0 1 5708 -1 0 3391
box 107 226 460 873
use sky130_fd_io__inv_1  sky130_fd_io__inv_1_0
timestamp 1701704242
transform 1 0 -745 0 1 1374
box -38 -49 326 715
use sky130_fd_io__tap_1  sky130_fd_io__tap_1_0
timestamp 1701704242
transform 1 0 -841 0 1 1374
box -38 -49 134 715
use sky130_fd_pr__nfet_01v8__example_55959141808770  sky130_fd_pr__nfet_01v8__example_55959141808770_0
timestamp 1701704242
transform -1 0 -16 0 1 901
box -1 0 161 1
use sky130_fd_pr__nfet_01v8__example_55959141808771  sky130_fd_pr__nfet_01v8__example_55959141808771_0
timestamp 1701704242
transform -1 0 979 0 1 901
box -1 0 377 1
use sky130_fd_pr__nfet_01v8__example_55959141808772  sky130_fd_pr__nfet_01v8__example_55959141808772_0
timestamp 1701704242
transform 0 -1 2143 -1 0 266
box -1 0 181 1
use sky130_fd_pr__nfet_01v8__example_55959141808773  sky130_fd_pr__nfet_01v8__example_55959141808773_0
timestamp 1701704242
transform 0 -1 2143 -1 0 629
box -1 0 181 1
use sky130_fd_pr__nfet_01v8__example_55959141808774  sky130_fd_pr__nfet_01v8__example_55959141808774_0
timestamp 1701704242
transform 1 0 2742 0 -1 679
box -1 0 413 1
use sky130_fd_pr__nfet_01v8__example_55959141808775  sky130_fd_pr__nfet_01v8__example_55959141808775_0
timestamp 1701704242
transform 1 0 1035 0 1 901
box -1 0 809 1
use sky130_fd_pr__nfet_01v8__example_55959141808776  sky130_fd_pr__nfet_01v8__example_55959141808776_0
timestamp 1701704242
transform -1 0 547 0 1 901
box -1 0 377 1
use sky130_fd_pr__nfet_01v8__example_55959141808777  sky130_fd_pr__nfet_01v8__example_55959141808777_0
timestamp 1701704242
transform 1 0 3491 0 1 1301
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808777  sky130_fd_pr__nfet_01v8__example_55959141808777_1
timestamp 1701704242
transform 1 0 2176 0 1 1286
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808777  sky130_fd_pr__nfet_01v8__example_55959141808777_2
timestamp 1701704242
transform 1 0 2459 0 1 1286
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808778  sky130_fd_pr__nfet_01v8__example_55959141808778_0
timestamp 1701704242
transform 1 0 2742 0 1 907
box -1 0 257 1
use sky130_fd_pr__nfet_01v8__example_55959141808778  sky130_fd_pr__nfet_01v8__example_55959141808778_1
timestamp 1701704242
transform 1 0 3054 0 1 907
box -1 0 257 1
use sky130_fd_pr__nfet_01v8__example_55959141808779  sky130_fd_pr__nfet_01v8__example_55959141808779_0
timestamp 1701704242
transform -1 0 469 0 -1 2237
box -1 0 181 1
use sky130_fd_pr__nfet_01v8__example_55959141808779  sky130_fd_pr__nfet_01v8__example_55959141808779_1
timestamp 1701704242
transform 1 0 3934 0 1 1659
box -1 0 181 1
use sky130_fd_pr__pfet_01v8__example_55959141808780  sky130_fd_pr__pfet_01v8__example_55959141808780_0
timestamp 1701704242
transform 1 0 1100 0 1 2580
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808781  sky130_fd_pr__pfet_01v8__example_55959141808781_0
timestamp 1701704242
transform 1 0 2802 0 -1 3545
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808783  sky130_fd_pr__pfet_01v8__example_55959141808783_0
timestamp 1701704242
transform -1 0 2456 0 -1 3482
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808783  sky130_fd_pr__pfet_01v8__example_55959141808783_1
timestamp 1701704242
transform 1 0 2512 0 -1 3482
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808784  sky130_fd_pr__pfet_01v8__example_55959141808784_0
timestamp 1701704242
transform 1 0 5261 0 1 3288
box -1 0 161 1
use sky130_fd_pr__pfet_01v8__example_55959141808784  sky130_fd_pr__pfet_01v8__example_55959141808784_1
timestamp 1701704242
transform -1 0 5421 0 1 2782
box -1 0 161 1
use sky130_fd_pr__pfet_01v8__example_55959141808785  sky130_fd_pr__pfet_01v8__example_55959141808785_0
timestamp 1701704242
transform 1 0 3085 0 -1 3545
box -1 0 413 1
use sky130_fd_pr__pfet_01v8__example_55959141808786  sky130_fd_pr__pfet_01v8__example_55959141808786_0
timestamp 1701704242
transform 1 0 -545 0 1 2580
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808786  sky130_fd_pr__pfet_01v8__example_55959141808786_1
timestamp 1701704242
transform -1 0 -601 0 1 2580
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808786  sky130_fd_pr__pfet_01v8__example_55959141808786_2
timestamp 1701704242
transform 1 0 369 0 1 2580
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808786  sky130_fd_pr__pfet_01v8__example_55959141808786_3
timestamp 1701704242
transform -1 0 917 0 1 2580
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808786  sky130_fd_pr__pfet_01v8__example_55959141808786_4
timestamp 1701704242
transform 1 0 1460 0 1 2580
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808786  sky130_fd_pr__pfet_01v8__example_55959141808786_5
timestamp 1701704242
transform 1 0 1753 0 1 2545
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808786  sky130_fd_pr__pfet_01v8__example_55959141808786_6
timestamp 1701704242
transform -1 0 313 0 1 2580
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808787  sky130_fd_pr__pfet_01v8__example_55959141808787_0
timestamp 1701704242
transform 1 0 1909 0 1 2545
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808787  sky130_fd_pr__pfet_01v8__example_55959141808787_1
timestamp 1701704242
transform -1 0 761 0 1 2580
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808787  sky130_fd_pr__pfet_01v8__example_55959141808787_2
timestamp 1701704242
transform -1 0 4389 0 -1 3545
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808787  sky130_fd_pr__pfet_01v8__example_55959141808787_3
timestamp 1701704242
transform 1 0 2065 0 1 2545
box -1 0 101 1
use sky130_fd_pr__res_bent_nd__example_55959141808769  sky130_fd_pr__res_bent_nd__example_55959141808769_0
timestamp 1701704242
transform 0 1 -29280 1 0 -8697
box -42 -2244 -29 1
use sky130_fd_pr__res_bent_po__example_55959141808768  sky130_fd_pr__res_bent_po__example_55959141808768_0
timestamp 1701704242
transform 0 1 -9813 -1 0 4210
box -50 -1753 12854 8
<< labels >>
flabel comment s 3904 1775 3904 1775 0 FreeSans 440 0 0 0 SWICH
flabel comment s 1375 707 1375 707 0 FreeSans 440 0 0 0 SWICH
flabel metal1 s 5763 2942 5815 2994 3 FreeSans 520 270 0 0 VGND
port 2 nsew
flabel metal1 s 318 789 370 841 3 FreeSans 520 0 0 0 VGND
port 2 nsew
flabel metal1 s 3187 3140 3239 3192 3 FreeSans 520 0 0 0 IN_H
port 3 nsew
flabel metal1 s 208 3645 260 3697 3 FreeSans 520 0 0 0 VDDIO
port 4 nsew
flabel metal1 s 241 2397 287 2449 3 FreeSans 520 0 0 0 VNORMAL
port 5 nsew
flabel metal1 s 675 2435 727 2487 3 FreeSans 520 0 0 0 VNORMAL_B
port 6 nsew
flabel metal1 s 5321 2837 5373 2889 3 FreeSans 520 0 0 0 PAD
port 7 nsew
flabel metal1 s 1493 2441 1534 2493 3 FreeSans 520 0 0 0 ENABLE_HV
port 8 nsew
flabel metal1 s 3133 2854 3185 2900 3 FreeSans 520 0 0 0 IN_H_N
port 9 nsew
flabel metal1 s -729 2135 -608 2224 3 FreeSans 520 0 0 0 VCCHIB
port 10 nsew
flabel metal1 s -663 1652 -628 1699 3 FreeSans 520 0 0 0 ENABLE_VDDIO_LV
port 11 nsew
<< properties >>
string GDS_END 56281106
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 55112898
<< end >>
