magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< pwell >>
rect -76 -26 724 226
<< mvnmos >>
rect 0 0 120 200
rect 176 0 296 200
rect 352 0 472 200
rect 528 0 648 200
<< mvndiff >>
rect -50 0 0 200
rect 648 0 698 200
<< poly >>
rect 0 200 120 226
rect 0 -26 120 0
rect 176 200 296 226
rect 176 -26 296 0
rect 352 200 472 226
rect 352 -26 472 0
rect 528 200 648 226
rect 528 -26 648 0
<< metal1 >>
rect -51 -16 -5 186
rect 125 -16 171 186
rect 301 -16 347 186
rect 477 -16 523 186
rect 653 -16 699 186
use hvDFM1sd2_CDNS_52468879185104  hvDFM1sd2_CDNS_52468879185104_0
timestamp 1701704242
transform 1 0 472 0 1 0
box -26 -26 82 226
use hvDFM1sd2_CDNS_52468879185104  hvDFM1sd2_CDNS_52468879185104_1
timestamp 1701704242
transform 1 0 296 0 1 0
box -26 -26 82 226
use hvDFM1sd2_CDNS_52468879185104  hvDFM1sd2_CDNS_52468879185104_2
timestamp 1701704242
transform 1 0 120 0 1 0
box -26 -26 82 226
use hvDFM1sd_CDNS_52468879185147  hvDFM1sd_CDNS_52468879185147_0
timestamp 1701704242
transform -1 0 0 0 1 0
box -26 -26 79 226
use hvDFM1sd_CDNS_52468879185147  hvDFM1sd_CDNS_52468879185147_1
timestamp 1701704242
transform 1 0 648 0 1 0
box -26 -26 79 226
<< labels >>
flabel comment s -28 85 -28 85 0 FreeSans 300 0 0 0 S
flabel comment s 148 85 148 85 0 FreeSans 300 0 0 0 D
flabel comment s 324 85 324 85 0 FreeSans 300 0 0 0 S
flabel comment s 500 85 500 85 0 FreeSans 300 0 0 0 D
flabel comment s 676 85 676 85 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 86868030
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86865640
<< end >>
