magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -85 1532 913 1568
rect -85 800 63 1532
rect 773 800 913 1532
<< pwell >>
rect -45 76 45 728
<< mvpsubdiff >>
rect -19 665 19 702
rect -19 631 -17 665
rect 17 631 19 665
rect -19 597 19 631
rect -19 563 -17 597
rect 17 563 19 597
rect -19 529 19 563
rect -19 495 -17 529
rect 17 495 19 529
rect -19 461 19 495
rect -19 427 -17 461
rect 17 427 19 461
rect -19 393 19 427
rect -19 359 -17 393
rect 17 359 19 393
rect -19 325 19 359
rect -19 291 -17 325
rect 17 291 19 325
rect -19 257 19 291
rect -19 223 -17 257
rect 17 223 19 257
rect -19 189 19 223
rect -19 155 -17 189
rect 17 155 19 189
rect -19 102 19 155
<< mvnsubdiff >>
rect -19 1413 19 1462
rect -19 1379 -17 1413
rect 17 1379 19 1413
rect -19 1345 19 1379
rect -19 1311 -17 1345
rect 17 1311 19 1345
rect -19 1277 19 1311
rect -19 1243 -17 1277
rect 17 1243 19 1277
rect -19 1209 19 1243
rect -19 1175 -17 1209
rect 17 1175 19 1209
rect -19 1134 19 1175
rect -19 1100 -17 1134
rect 17 1100 19 1134
rect -19 1066 19 1100
rect -19 1032 -17 1066
rect 17 1032 19 1066
rect -19 998 19 1032
rect -19 964 -17 998
rect 17 964 19 998
rect -19 930 19 964
rect -19 896 -17 930
rect 17 896 19 930
rect -19 866 19 896
rect 809 1413 847 1462
rect 809 1379 811 1413
rect 845 1379 847 1413
rect 809 1345 847 1379
rect 809 1311 811 1345
rect 845 1311 847 1345
rect 809 1277 847 1311
rect 809 1243 811 1277
rect 845 1243 847 1277
rect 809 1209 847 1243
rect 809 1175 811 1209
rect 845 1175 847 1209
rect 809 1134 847 1175
rect 809 1100 811 1134
rect 845 1100 847 1134
rect 809 1066 847 1100
rect 809 1032 811 1066
rect 845 1032 847 1066
rect 809 998 847 1032
rect 809 964 811 998
rect 845 964 847 998
rect 809 930 847 964
rect 809 896 811 930
rect 845 896 847 930
rect 809 866 847 896
<< mvpsubdiffcont >>
rect -17 631 17 665
rect -17 563 17 597
rect -17 495 17 529
rect -17 427 17 461
rect -17 359 17 393
rect -17 291 17 325
rect -17 223 17 257
rect -17 155 17 189
<< mvnsubdiffcont >>
rect -17 1379 17 1413
rect -17 1311 17 1345
rect -17 1243 17 1277
rect -17 1175 17 1209
rect -17 1100 17 1134
rect -17 1032 17 1066
rect -17 964 17 998
rect -17 896 17 930
rect 811 1379 845 1413
rect 811 1311 845 1345
rect 811 1243 845 1277
rect 811 1175 845 1209
rect 811 1100 845 1134
rect 811 1032 845 1066
rect 811 964 845 998
rect 811 896 845 930
<< poly >>
rect 290 1548 702 1568
rect 290 1514 342 1548
rect 376 1514 410 1548
rect 444 1514 478 1548
rect 512 1514 546 1548
rect 580 1514 614 1548
rect 648 1514 702 1548
rect 290 1492 702 1514
rect 92 782 234 840
rect 92 748 112 782
rect 146 748 180 782
rect 214 748 234 782
rect 92 728 234 748
rect 498 785 794 840
rect 498 751 527 785
rect 561 751 595 785
rect 629 751 663 785
rect 697 751 731 785
rect 765 751 794 785
rect 498 728 794 751
rect 146 54 442 76
rect 146 20 175 54
rect 209 20 243 54
rect 277 20 311 54
rect 345 20 379 54
rect 413 20 442 54
rect 146 0 442 20
rect 498 54 794 76
rect 498 20 527 54
rect 561 20 595 54
rect 629 20 663 54
rect 697 20 731 54
rect 765 20 794 54
rect 498 0 794 20
<< polycont >>
rect 342 1514 376 1548
rect 410 1514 444 1548
rect 478 1514 512 1548
rect 546 1514 580 1548
rect 614 1514 648 1548
rect 112 748 146 782
rect 180 748 214 782
rect 527 751 561 785
rect 595 751 629 785
rect 663 751 697 785
rect 731 751 765 785
rect 175 20 209 54
rect 243 20 277 54
rect 311 20 345 54
rect 379 20 413 54
rect 527 20 561 54
rect 595 20 629 54
rect 663 20 697 54
rect 731 20 765 54
<< locali >>
rect 326 1514 342 1548
rect 376 1514 410 1548
rect 444 1514 478 1548
rect 512 1514 546 1548
rect 580 1514 614 1548
rect 648 1514 664 1548
rect -17 1413 17 1454
rect -17 1345 17 1379
rect 811 1413 845 1454
rect 811 1345 845 1379
rect -17 1277 17 1311
rect 123 1298 161 1332
rect 409 1298 447 1332
rect 675 1298 713 1332
rect -17 1209 17 1243
rect -17 1134 17 1175
rect 811 1277 845 1311
rect 811 1209 845 1243
rect 811 1134 845 1175
rect -17 1066 17 1068
rect -17 1030 17 1032
rect -17 958 17 964
rect 245 1030 279 1068
rect 245 958 279 996
rect 557 1030 591 1068
rect 557 958 591 996
rect -17 874 17 896
rect 96 748 112 782
rect 146 748 180 782
rect 214 748 230 782
rect 401 717 435 928
rect 811 1066 845 1068
rect 811 1030 845 1032
rect 811 958 845 964
rect 811 874 845 896
rect 511 751 527 785
rect 561 751 595 785
rect 629 751 663 785
rect 697 751 731 785
rect 765 751 781 785
rect -17 665 17 694
rect 401 674 663 717
rect 629 640 663 674
rect -17 597 17 631
rect -17 529 17 542
rect -17 461 17 470
rect 277 504 311 542
rect 277 432 311 470
rect -17 393 17 398
rect -17 325 17 359
rect 169 295 207 329
rect 449 295 487 329
rect 733 295 771 329
rect -17 257 17 291
rect -17 189 17 223
rect -17 110 17 155
rect 159 20 175 54
rect 209 20 243 54
rect 277 20 311 54
rect 345 20 379 54
rect 413 20 429 54
rect 511 20 527 54
rect 561 20 595 54
rect 629 20 663 54
rect 697 20 731 54
rect 765 20 781 54
<< viali >>
rect 89 1298 123 1332
rect 161 1298 195 1332
rect 375 1298 409 1332
rect 447 1298 481 1332
rect 641 1298 675 1332
rect 713 1298 747 1332
rect -17 1100 17 1102
rect -17 1068 17 1100
rect -17 998 17 1030
rect -17 996 17 998
rect -17 930 17 958
rect -17 924 17 930
rect 245 1068 279 1102
rect 245 996 279 1030
rect 245 924 279 958
rect 557 1068 591 1102
rect 557 996 591 1030
rect 557 924 591 958
rect 811 1100 845 1102
rect 811 1068 845 1100
rect 811 998 845 1030
rect 811 996 845 998
rect 811 930 845 958
rect 811 924 845 930
rect -17 563 17 576
rect -17 542 17 563
rect -17 495 17 504
rect -17 470 17 495
rect -17 427 17 432
rect -17 398 17 427
rect 277 542 311 576
rect 277 470 311 504
rect 277 398 311 432
rect 135 295 169 329
rect 207 295 241 329
rect 415 295 449 329
rect 487 295 521 329
rect 699 295 733 329
rect 771 295 805 329
<< metal1 >>
rect 77 1332 759 1338
rect 77 1298 89 1332
rect 123 1298 161 1332
rect 195 1298 375 1332
rect 409 1298 447 1332
rect 481 1298 641 1332
rect 675 1298 713 1332
rect 747 1298 759 1332
rect 77 1292 759 1298
rect -29 1102 857 1108
rect -29 1068 -17 1102
rect 17 1068 245 1102
rect 279 1068 557 1102
rect 591 1068 811 1102
rect 845 1068 857 1102
rect -29 1030 857 1068
rect -29 996 -17 1030
rect 17 996 245 1030
rect 279 996 557 1030
rect 591 996 811 1030
rect 845 996 857 1030
rect -29 958 857 996
rect -29 924 -17 958
rect 17 924 245 958
rect 279 924 557 958
rect 591 924 811 958
rect 845 924 857 958
rect -29 906 857 924
rect -29 576 857 582
rect -29 542 -17 576
rect 17 542 277 576
rect 311 542 857 576
rect -29 504 857 542
rect -29 470 -17 504
rect 17 470 277 504
rect 311 470 857 504
rect -29 432 857 470
rect -29 398 -17 432
rect 17 398 277 432
rect 311 398 857 432
rect -29 380 857 398
rect 129 329 811 341
rect 129 295 135 329
rect 169 295 207 329
rect 241 295 415 329
rect 449 295 487 329
rect 521 295 699 329
rect 733 295 771 329
rect 805 295 811 329
rect 129 283 811 295
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_0
timestamp 1701704242
transform 0 -1 241 1 0 295
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_1
timestamp 1701704242
transform 0 -1 521 1 0 295
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_2
timestamp 1701704242
transform 0 -1 805 1 0 295
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1701704242
transform -1 0 195 0 -1 1332
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1701704242
transform -1 0 747 0 -1 1332
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1701704242
transform -1 0 481 0 -1 1332
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_0
timestamp 1701704242
transform 1 0 245 0 -1 1102
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_1
timestamp 1701704242
transform 1 0 557 0 -1 1102
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_2
timestamp 1701704242
transform 1 0 -17 0 -1 1102
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_3
timestamp 1701704242
transform 1 0 811 0 -1 1102
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_4
timestamp 1701704242
transform 1 0 277 0 1 398
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_5
timestamp 1701704242
transform 1 0 -17 0 1 398
box 0 0 1 1
use nfet_CDNS_52468879185365  nfet_CDNS_52468879185365_0
timestamp 1701704242
transform 1 0 146 0 1 102
box -79 -26 375 626
use nfet_CDNS_52468879185365  nfet_CDNS_52468879185365_1
timestamp 1701704242
transform 1 0 498 0 1 102
box -79 -26 375 626
use pfet_CDNS_52468879185366  pfet_CDNS_52468879185366_0
timestamp 1701704242
transform 1 0 290 0 -1 1466
box -119 -66 531 666
use pfet_CDNS_52468879185367  pfet_CDNS_52468879185367_0
timestamp 1701704242
transform -1 0 234 0 -1 1466
box -119 -66 219 666
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_0
timestamp 1701704242
transform 0 -1 230 -1 0 798
box 0 0 1 1
use PYL1_CDNS_52468879185289  PYL1_CDNS_52468879185289_0
timestamp 1701704242
transform 0 1 326 1 0 1498
box 0 0 1 1
use PYL1_CDNS_52468879185309  PYL1_CDNS_52468879185309_0
timestamp 1701704242
transform 0 -1 781 -1 0 801
box 0 0 1 1
use PYL1_CDNS_52468879185309  PYL1_CDNS_52468879185309_1
timestamp 1701704242
transform 0 1 159 1 0 4
box 0 0 1 1
use PYL1_CDNS_52468879185309  PYL1_CDNS_52468879185309_2
timestamp 1701704242
transform 0 1 511 1 0 4
box 0 0 1 1
<< labels >>
flabel comment s 389 312 389 312 0 FreeSans 200 0 0 0 int
flabel metal1 s 820 906 857 1108 6 FreeSans 300 180 0 0 vcc_io
port 1 nsew
flabel metal1 s 719 1292 759 1338 3 FreeSans 300 0 0 0 pu_h_n
port 2 nsew
flabel metal1 s 823 380 857 582 7 FreeSans 300 180 0 0 vgnd_io
port 3 nsew
flabel metal1 s -29 906 8 1108 7 FreeSans 300 0 0 0 vcc_io
port 1 nsew
flabel metal1 s -29 380 5 582 7 FreeSans 300 0 0 0 vgnd_io
port 3 nsew
flabel metal1 s 77 1292 117 1338 3 FreeSans 300 180 0 0 pu_h_n
port 2 nsew
flabel locali s 747 751 781 785 7 FreeSans 300 0 0 0 drvhi_h
port 5 nsew
flabel locali s 96 748 130 782 8 FreeSans 300 0 0 0 puen_h
port 6 nsew
<< properties >>
string GDS_END 87986800
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 87980940
<< end >>
