magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -38 261 2798 582
<< pwell >>
rect 1408 157 1769 201
rect 2201 157 2744 203
rect 1 21 2744 157
rect 29 -17 63 21
<< locali >>
rect 17 153 68 335
rect 210 153 267 335
rect 581 323 617 392
rect 581 211 713 323
rect 581 145 620 211
rect 2408 299 2474 490
rect 2429 265 2474 299
rect 2576 265 2642 493
rect 2429 211 2642 265
rect 2429 165 2474 211
rect 2408 55 2474 165
rect 2576 51 2642 211
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2760 561
rect 17 405 69 493
rect 103 439 157 527
rect 191 451 409 493
rect 191 405 225 451
rect 454 417 504 493
rect 538 428 597 527
rect 17 369 225 405
rect 259 369 339 417
rect 108 255 164 335
rect 108 221 121 255
rect 155 221 164 255
rect 108 153 164 221
rect 301 142 339 369
rect 373 354 504 417
rect 651 400 685 465
rect 719 455 785 527
rect 819 427 888 493
rect 651 398 797 400
rect 373 181 440 354
rect 651 366 799 398
rect 474 255 540 320
rect 474 221 489 255
rect 523 221 540 255
rect 474 215 540 221
rect 373 143 504 181
rect 747 177 799 366
rect 301 141 335 142
rect 299 133 335 141
rect 295 132 335 133
rect 295 129 334 132
rect 292 127 333 129
rect 289 126 333 127
rect 288 124 333 126
rect 286 123 332 124
rect 284 122 332 123
rect 281 121 332 122
rect 279 120 332 121
rect 276 119 332 120
rect 17 17 140 119
rect 174 115 330 119
rect 174 111 328 115
rect 174 51 325 111
rect 365 17 418 109
rect 452 51 504 143
rect 654 143 799 177
rect 833 284 888 427
rect 923 323 966 493
rect 1007 427 1151 493
rect 1189 455 1266 527
rect 923 318 983 323
rect 932 289 983 318
rect 1041 315 1083 391
rect 833 218 898 284
rect 538 17 620 111
rect 654 51 691 143
rect 833 117 867 218
rect 932 184 966 289
rect 1117 279 1151 427
rect 1321 421 1364 490
rect 1412 425 1603 527
rect 1637 425 1798 492
rect 1832 447 1898 527
rect 1185 387 1364 421
rect 1764 413 1798 425
rect 1932 413 1993 490
rect 2031 447 2097 527
rect 1185 315 1219 387
rect 1328 289 1413 353
rect 1447 334 1627 391
rect 1017 255 1295 279
rect 1471 255 1543 265
rect 725 17 791 109
rect 825 51 867 117
rect 901 51 966 184
rect 1000 245 1543 255
rect 1000 51 1088 245
rect 1129 161 1195 203
rect 1261 195 1543 245
rect 1577 181 1627 334
rect 1685 215 1730 381
rect 1764 379 2097 413
rect 1776 323 1989 345
rect 1776 289 1788 323
rect 1822 309 1989 323
rect 2031 321 2097 379
rect 1822 289 1827 309
rect 1776 285 1827 289
rect 2131 273 2183 493
rect 1764 181 1821 251
rect 1129 127 1307 161
rect 1122 17 1219 93
rect 1257 51 1307 127
rect 1341 17 1543 161
rect 1577 144 1821 181
rect 1864 239 2183 273
rect 1864 171 1906 239
rect 1942 157 2103 203
rect 1942 109 1982 157
rect 2137 117 2183 239
rect 1693 55 1982 109
rect 2023 17 2073 109
rect 2115 51 2183 117
rect 2217 265 2269 493
rect 2303 299 2374 527
rect 2508 299 2542 527
rect 2676 299 2743 527
rect 2217 199 2395 265
rect 2217 51 2269 199
rect 2303 17 2374 165
rect 2508 17 2542 177
rect 2676 17 2743 177
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2760 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 2605 527 2639 561
rect 2697 527 2731 561
rect 121 221 155 255
rect 489 221 523 255
rect 1788 289 1822 323
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
rect 2605 -17 2639 17
rect 2697 -17 2731 17
<< metal1 >>
rect 0 561 2760 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2760 561
rect 0 496 2760 527
rect 1316 320 1374 329
rect 1776 323 1834 329
rect 1776 320 1788 323
rect 1316 292 1788 320
rect 1316 283 1374 292
rect 1776 289 1788 292
rect 1822 289 1834 323
rect 1776 283 1834 289
rect 109 255 167 261
rect 109 221 121 255
rect 155 252 167 255
rect 477 255 535 261
rect 477 252 489 255
rect 155 224 489 252
rect 155 221 167 224
rect 109 215 167 221
rect 477 221 489 224
rect 523 221 535 255
rect 477 215 535 221
rect 0 17 2760 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2760 17
rect 0 -48 2760 -17
<< obsm1 >>
rect 753 388 811 397
rect 1029 388 1087 397
rect 1500 388 1558 397
rect 753 360 1558 388
rect 753 351 811 360
rect 1029 351 1087 360
rect 1500 351 1558 360
rect 293 320 351 329
rect 937 320 995 329
rect 293 292 995 320
rect 293 283 351 292
rect 937 283 995 292
rect 845 252 903 261
rect 1684 252 1742 261
rect 845 224 1742 252
rect 845 215 903 224
rect 1684 215 1742 224
<< labels >>
rlabel locali s 581 145 620 211 6 CLK
port 1 nsew clock input
rlabel locali s 581 211 713 323 6 CLK
port 1 nsew clock input
rlabel locali s 581 323 617 392 6 CLK
port 1 nsew clock input
rlabel locali s 210 153 267 335 6 D
port 2 nsew signal input
rlabel locali s 17 153 68 335 6 SCD
port 3 nsew signal input
rlabel metal1 s 477 215 535 224 6 SCE
port 4 nsew signal input
rlabel metal1 s 109 215 167 224 6 SCE
port 4 nsew signal input
rlabel metal1 s 109 224 535 252 6 SCE
port 4 nsew signal input
rlabel metal1 s 477 252 535 261 6 SCE
port 4 nsew signal input
rlabel metal1 s 109 252 167 261 6 SCE
port 4 nsew signal input
rlabel metal1 s 1776 283 1834 292 6 SET_B
port 5 nsew signal input
rlabel metal1 s 1316 283 1374 292 6 SET_B
port 5 nsew signal input
rlabel metal1 s 1316 292 1834 320 6 SET_B
port 5 nsew signal input
rlabel metal1 s 1776 320 1834 329 6 SET_B
port 5 nsew signal input
rlabel metal1 s 1316 320 1374 329 6 SET_B
port 5 nsew signal input
rlabel metal1 s 0 -48 2760 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 1 21 2744 157 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 2201 157 2744 203 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 1408 157 1769 201 6 VNB
port 7 nsew ground bidirectional
rlabel nwell s -38 261 2798 582 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 496 2760 592 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 2576 51 2642 211 6 Q
port 10 nsew signal output
rlabel locali s 2408 55 2474 165 6 Q
port 10 nsew signal output
rlabel locali s 2429 165 2474 211 6 Q
port 10 nsew signal output
rlabel locali s 2429 211 2642 265 6 Q
port 10 nsew signal output
rlabel locali s 2576 265 2642 493 6 Q
port 10 nsew signal output
rlabel locali s 2429 265 2474 299 6 Q
port 10 nsew signal output
rlabel locali s 2408 299 2474 490 6 Q
port 10 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 2760 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 326040
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 304594
<< end >>
