magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< pwell >>
rect -76 -26 276 226
<< mvnmos >>
rect 0 0 200 200
<< mvndiff >>
rect -50 0 0 200
rect 200 0 250 200
<< poly >>
rect 0 200 200 226
rect 0 -26 200 0
<< metal1 >>
rect -51 -16 -5 186
rect 205 -16 251 186
use hvDFM1sd_CDNS_52468879185147  hvDFM1sd_CDNS_52468879185147_0
timestamp 1701704242
transform -1 0 0 0 1 0
box -26 -26 79 226
use hvDFM1sd_CDNS_52468879185147  hvDFM1sd_CDNS_52468879185147_1
timestamp 1701704242
transform 1 0 200 0 1 0
box -26 -26 79 226
<< labels >>
flabel comment s -28 85 -28 85 0 FreeSans 300 0 0 0 S
flabel comment s 228 85 228 85 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 86001648
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86000758
<< end >>
