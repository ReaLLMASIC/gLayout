magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< pwell >>
rect -76 -26 176 626
<< mvnmos >>
rect 0 0 100 600
<< mvndiff >>
rect -50 0 0 600
rect 100 0 150 600
<< poly >>
rect 0 600 100 626
rect 0 -26 100 0
<< locali >>
rect -45 -4 -11 538
rect 111 -4 145 538
use hvDFL1sd_CDNS_52468879185311  hvDFL1sd_CDNS_52468879185311_0
timestamp 1701704242
transform -1 0 0 0 1 0
box -26 -26 79 626
use hvDFL1sd_CDNS_52468879185311  hvDFL1sd_CDNS_52468879185311_1
timestamp 1701704242
transform 1 0 100 0 1 0
box -26 -26 79 626
<< labels >>
flabel comment s -28 267 -28 267 0 FreeSans 300 0 0 0 S
flabel comment s 128 267 128 267 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 87767628
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 87766738
<< end >>
