magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -119 -66 927 266
<< mvpmos >>
rect 0 0 160 200
rect 216 0 376 200
rect 432 0 592 200
rect 648 0 808 200
<< mvpdiff >>
rect -53 182 0 200
rect -53 148 -45 182
rect -11 148 0 182
rect -53 114 0 148
rect -53 80 -45 114
rect -11 80 0 114
rect -53 46 0 80
rect -53 12 -45 46
rect -11 12 0 46
rect -53 0 0 12
rect 160 182 216 200
rect 160 148 171 182
rect 205 148 216 182
rect 160 114 216 148
rect 160 80 171 114
rect 205 80 216 114
rect 160 46 216 80
rect 160 12 171 46
rect 205 12 216 46
rect 160 0 216 12
rect 376 182 432 200
rect 376 148 387 182
rect 421 148 432 182
rect 376 114 432 148
rect 376 80 387 114
rect 421 80 432 114
rect 376 46 432 80
rect 376 12 387 46
rect 421 12 432 46
rect 376 0 432 12
rect 592 182 648 200
rect 592 148 603 182
rect 637 148 648 182
rect 592 114 648 148
rect 592 80 603 114
rect 637 80 648 114
rect 592 46 648 80
rect 592 12 603 46
rect 637 12 648 46
rect 592 0 648 12
rect 808 182 861 200
rect 808 148 819 182
rect 853 148 861 182
rect 808 114 861 148
rect 808 80 819 114
rect 853 80 861 114
rect 808 46 861 80
rect 808 12 819 46
rect 853 12 861 46
rect 808 0 861 12
<< mvpdiffc >>
rect -45 148 -11 182
rect -45 80 -11 114
rect -45 12 -11 46
rect 171 148 205 182
rect 171 80 205 114
rect 171 12 205 46
rect 387 148 421 182
rect 387 80 421 114
rect 387 12 421 46
rect 603 148 637 182
rect 603 80 637 114
rect 603 12 637 46
rect 819 148 853 182
rect 819 80 853 114
rect 819 12 853 46
<< poly >>
rect 0 200 160 226
rect 216 200 376 226
rect 432 200 592 226
rect 648 200 808 226
rect 0 -26 160 0
rect 216 -26 376 0
rect 432 -26 592 0
rect 648 -26 808 0
<< locali >>
rect -45 182 -11 198
rect -45 114 -11 148
rect -45 46 -11 80
rect -45 -4 -11 12
rect 171 182 205 198
rect 171 114 205 148
rect 171 46 205 80
rect 171 -4 205 12
rect 387 182 421 198
rect 387 114 421 148
rect 387 46 421 80
rect 387 -4 421 12
rect 603 182 637 198
rect 603 114 637 148
rect 603 46 637 80
rect 603 -4 637 12
rect 819 182 853 198
rect 819 114 853 148
rect 819 46 853 80
rect 819 -4 853 12
use hvDFL1sd2_CDNS_52468879185110  hvDFL1sd2_CDNS_52468879185110_0
timestamp 1701704242
transform 1 0 592 0 1 0
box 0 0 1 1
use hvDFL1sd2_CDNS_52468879185110  hvDFL1sd2_CDNS_52468879185110_1
timestamp 1701704242
transform 1 0 376 0 1 0
box 0 0 1 1
use hvDFL1sd2_CDNS_52468879185110  hvDFL1sd2_CDNS_52468879185110_2
timestamp 1701704242
transform 1 0 160 0 1 0
box 0 0 1 1
use hvDFL1sd_CDNS_5246887918589  hvDFL1sd_CDNS_5246887918589_0
timestamp 1701704242
transform -1 0 0 0 1 0
box 0 0 1 1
use hvDFL1sd_CDNS_5246887918589  hvDFL1sd_CDNS_5246887918589_1
timestamp 1701704242
transform 1 0 808 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s -28 97 -28 97 0 FreeSans 300 0 0 0 S
flabel comment s 188 97 188 97 0 FreeSans 300 0 0 0 D
flabel comment s 404 97 404 97 0 FreeSans 300 0 0 0 S
flabel comment s 620 97 620 97 0 FreeSans 300 0 0 0 D
flabel comment s 836 97 836 97 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 87754358
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 87751840
<< end >>
