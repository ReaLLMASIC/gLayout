magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -107 515 795 1337
<< pwell >>
rect -67 367 67 455
rect -51 345 67 367
rect 285 345 419 455
rect 637 367 771 455
rect 637 345 755 367
rect -51 93 755 345
<< mvnmos >>
rect 28 119 148 319
rect 204 119 324 319
rect 380 119 500 319
rect 556 119 676 319
<< mvpmos >>
rect 28 671 148 1271
rect 204 671 324 1271
rect 380 671 500 1271
rect 556 671 676 1271
<< mvndiff >>
rect -25 307 28 319
rect -25 273 -17 307
rect 17 273 28 307
rect -25 239 28 273
rect -25 205 -17 239
rect 17 205 28 239
rect -25 171 28 205
rect -25 137 -17 171
rect 17 137 28 171
rect -25 119 28 137
rect 148 307 204 319
rect 148 273 159 307
rect 193 273 204 307
rect 148 239 204 273
rect 148 205 159 239
rect 193 205 204 239
rect 148 171 204 205
rect 148 137 159 171
rect 193 137 204 171
rect 148 119 204 137
rect 324 307 380 319
rect 324 273 335 307
rect 369 273 380 307
rect 324 239 380 273
rect 324 205 335 239
rect 369 205 380 239
rect 324 171 380 205
rect 324 137 335 171
rect 369 137 380 171
rect 324 119 380 137
rect 500 307 556 319
rect 500 273 511 307
rect 545 273 556 307
rect 500 239 556 273
rect 500 205 511 239
rect 545 205 556 239
rect 500 171 556 205
rect 500 137 511 171
rect 545 137 556 171
rect 500 119 556 137
rect 676 307 729 319
rect 676 273 687 307
rect 721 273 729 307
rect 676 239 729 273
rect 676 205 687 239
rect 721 205 729 239
rect 676 171 729 205
rect 676 137 687 171
rect 721 137 729 171
rect 676 119 729 137
<< mvpdiff >>
rect -25 1193 28 1271
rect -25 1159 -17 1193
rect 17 1159 28 1193
rect -25 1125 28 1159
rect -25 1091 -17 1125
rect 17 1091 28 1125
rect -25 1057 28 1091
rect -25 1023 -17 1057
rect 17 1023 28 1057
rect -25 989 28 1023
rect -25 955 -17 989
rect 17 955 28 989
rect -25 921 28 955
rect -25 887 -17 921
rect 17 887 28 921
rect -25 853 28 887
rect -25 819 -17 853
rect 17 819 28 853
rect -25 785 28 819
rect -25 751 -17 785
rect 17 751 28 785
rect -25 717 28 751
rect -25 683 -17 717
rect 17 683 28 717
rect -25 671 28 683
rect 148 1193 204 1271
rect 148 1159 159 1193
rect 193 1159 204 1193
rect 148 1125 204 1159
rect 148 1091 159 1125
rect 193 1091 204 1125
rect 148 1057 204 1091
rect 148 1023 159 1057
rect 193 1023 204 1057
rect 148 989 204 1023
rect 148 955 159 989
rect 193 955 204 989
rect 148 921 204 955
rect 148 887 159 921
rect 193 887 204 921
rect 148 853 204 887
rect 148 819 159 853
rect 193 819 204 853
rect 148 785 204 819
rect 148 751 159 785
rect 193 751 204 785
rect 148 717 204 751
rect 148 683 159 717
rect 193 683 204 717
rect 148 671 204 683
rect 324 1193 380 1271
rect 324 1159 335 1193
rect 369 1159 380 1193
rect 324 1125 380 1159
rect 324 1091 335 1125
rect 369 1091 380 1125
rect 324 1057 380 1091
rect 324 1023 335 1057
rect 369 1023 380 1057
rect 324 989 380 1023
rect 324 955 335 989
rect 369 955 380 989
rect 324 921 380 955
rect 324 887 335 921
rect 369 887 380 921
rect 324 853 380 887
rect 324 819 335 853
rect 369 819 380 853
rect 324 785 380 819
rect 324 751 335 785
rect 369 751 380 785
rect 324 717 380 751
rect 324 683 335 717
rect 369 683 380 717
rect 324 671 380 683
rect 500 1193 556 1271
rect 500 1159 511 1193
rect 545 1159 556 1193
rect 500 1125 556 1159
rect 500 1091 511 1125
rect 545 1091 556 1125
rect 500 1057 556 1091
rect 500 1023 511 1057
rect 545 1023 556 1057
rect 500 989 556 1023
rect 500 955 511 989
rect 545 955 556 989
rect 500 921 556 955
rect 500 887 511 921
rect 545 887 556 921
rect 500 853 556 887
rect 500 819 511 853
rect 545 819 556 853
rect 500 785 556 819
rect 500 751 511 785
rect 545 751 556 785
rect 500 717 556 751
rect 500 683 511 717
rect 545 683 556 717
rect 500 671 556 683
rect 676 1193 729 1271
rect 676 1159 687 1193
rect 721 1159 729 1193
rect 676 1125 729 1159
rect 676 1091 687 1125
rect 721 1091 729 1125
rect 676 1057 729 1091
rect 676 1023 687 1057
rect 721 1023 729 1057
rect 676 989 729 1023
rect 676 955 687 989
rect 721 955 729 989
rect 676 921 729 955
rect 676 887 687 921
rect 721 887 729 921
rect 676 853 729 887
rect 676 819 687 853
rect 721 819 729 853
rect 676 785 729 819
rect 676 751 687 785
rect 721 751 729 785
rect 676 717 729 751
rect 676 683 687 717
rect 721 683 729 717
rect 676 671 729 683
<< mvndiffc >>
rect -17 273 17 307
rect -17 205 17 239
rect -17 137 17 171
rect 159 273 193 307
rect 159 205 193 239
rect 159 137 193 171
rect 335 273 369 307
rect 335 205 369 239
rect 335 137 369 171
rect 511 273 545 307
rect 511 205 545 239
rect 511 137 545 171
rect 687 273 721 307
rect 687 205 721 239
rect 687 137 721 171
<< mvpdiffc >>
rect -17 1159 17 1193
rect -17 1091 17 1125
rect -17 1023 17 1057
rect -17 955 17 989
rect -17 887 17 921
rect -17 819 17 853
rect -17 751 17 785
rect -17 683 17 717
rect 159 1159 193 1193
rect 159 1091 193 1125
rect 159 1023 193 1057
rect 159 955 193 989
rect 159 887 193 921
rect 159 819 193 853
rect 159 751 193 785
rect 159 683 193 717
rect 335 1159 369 1193
rect 335 1091 369 1125
rect 335 1023 369 1057
rect 335 955 369 989
rect 335 887 369 921
rect 335 819 369 853
rect 335 751 369 785
rect 335 683 369 717
rect 511 1159 545 1193
rect 511 1091 545 1125
rect 511 1023 545 1057
rect 511 955 545 989
rect 511 887 545 921
rect 511 819 545 853
rect 511 751 545 785
rect 511 683 545 717
rect 687 1159 721 1193
rect 687 1091 721 1125
rect 687 1023 721 1057
rect 687 955 721 989
rect 687 887 721 921
rect 687 819 721 853
rect 687 751 721 785
rect 687 683 721 717
<< mvpsubdiff >>
rect -41 427 41 429
rect -41 393 -17 427
rect 17 393 41 427
rect 311 427 393 429
rect 311 393 335 427
rect 369 393 393 427
rect 663 427 745 429
rect 663 393 687 427
rect 721 393 745 427
<< mvnsubdiff >>
rect -41 583 -17 617
rect 17 583 41 617
rect -41 581 41 583
rect 311 583 335 617
rect 369 583 393 617
rect 311 581 393 583
<< mvpsubdiffcont >>
rect -17 393 17 427
rect 335 393 369 427
rect 687 393 721 427
<< mvnsubdiffcont >>
rect -17 583 17 617
rect 335 583 369 617
<< poly >>
rect 21 1353 683 1369
rect 21 1319 37 1353
rect 71 1319 105 1353
rect 139 1319 213 1353
rect 247 1319 281 1353
rect 315 1319 389 1353
rect 423 1319 457 1353
rect 491 1319 565 1353
rect 599 1319 633 1353
rect 667 1319 683 1353
rect 21 1303 683 1319
rect 28 1297 676 1303
rect 28 1271 148 1297
rect 204 1271 324 1297
rect 380 1271 500 1297
rect 556 1271 676 1297
rect 28 645 148 671
rect 52 345 148 645
rect 28 319 148 345
rect 204 645 324 671
rect 380 645 500 671
rect 204 345 300 645
rect 404 345 500 645
rect 204 319 324 345
rect 380 319 500 345
rect 556 645 676 671
rect 556 345 652 645
rect 556 319 676 345
rect 28 93 148 119
rect 204 93 324 119
rect 380 93 500 119
rect 556 93 676 119
rect 21 71 683 93
rect 21 37 37 71
rect 71 37 105 71
rect 139 37 213 71
rect 247 37 281 71
rect 315 37 389 71
rect 423 37 457 71
rect 491 37 565 71
rect 599 37 633 71
rect 667 37 683 71
rect 21 21 683 37
<< polycont >>
rect 37 1319 71 1353
rect 105 1319 139 1353
rect 213 1319 247 1353
rect 281 1319 315 1353
rect 389 1319 423 1353
rect 457 1319 491 1353
rect 565 1319 599 1353
rect 633 1319 667 1353
rect 37 37 71 71
rect 105 37 139 71
rect 213 37 247 71
rect 281 37 315 71
rect 389 37 423 71
rect 457 37 491 71
rect 565 37 599 71
rect 633 37 667 71
<< locali >>
rect 37 1353 139 1369
rect 71 1319 105 1353
rect 37 1303 139 1319
rect 213 1353 491 1369
rect 247 1319 281 1353
rect 315 1319 389 1353
rect 423 1319 457 1353
rect 213 1303 491 1319
rect 565 1353 667 1369
rect 599 1319 633 1353
rect 565 1303 667 1319
rect -17 1193 17 1209
rect -17 1125 17 1159
rect -17 1057 17 1091
rect -17 989 17 1023
rect -17 921 17 955
rect -17 857 17 887
rect -17 785 17 819
rect -17 717 17 751
rect -17 667 17 679
rect -17 567 17 583
rect -17 427 17 443
rect -17 259 17 273
rect -17 187 17 205
rect -17 121 17 137
rect 51 87 125 1303
rect 159 1193 193 1270
rect 159 1125 193 1159
rect 159 1057 193 1091
rect 159 989 193 1023
rect 159 921 193 955
rect 159 853 193 887
rect 159 785 193 819
rect 159 717 193 751
rect 159 485 193 683
rect 159 307 193 451
rect 159 239 193 273
rect 159 171 193 205
rect 159 121 193 137
rect 227 87 301 1303
rect 335 1193 369 1209
rect 335 1125 369 1159
rect 335 1057 369 1091
rect 335 989 369 1023
rect 335 921 369 955
rect 335 857 369 887
rect 335 785 369 819
rect 335 717 369 751
rect 335 667 369 679
rect 335 567 369 583
rect 335 427 369 443
rect 335 259 369 273
rect 335 187 369 205
rect 335 121 369 137
rect 403 87 477 1303
rect 511 1193 545 1270
rect 511 1125 545 1159
rect 511 1057 545 1091
rect 511 989 545 1023
rect 511 921 545 955
rect 511 853 545 887
rect 511 785 545 819
rect 511 717 545 751
rect 511 485 545 683
rect 511 307 545 451
rect 511 239 545 273
rect 511 171 545 205
rect 511 121 545 137
rect 579 87 653 1303
rect 687 1193 721 1209
rect 687 1125 721 1159
rect 687 1057 721 1091
rect 687 989 721 1023
rect 687 921 721 955
rect 687 857 721 887
rect 687 785 721 819
rect 687 717 721 751
rect 687 667 721 679
rect 687 567 721 599
rect 687 427 721 443
rect 687 259 721 273
rect 687 187 721 205
rect 687 121 721 137
rect 37 71 139 87
rect 71 37 105 71
rect 37 21 139 37
rect 213 71 491 87
rect 247 37 281 71
rect 315 37 389 71
rect 423 37 457 71
rect 213 21 491 37
rect 565 71 667 87
rect 599 37 633 71
rect 565 21 667 37
<< viali >>
rect -17 853 17 857
rect -17 823 17 853
rect -17 751 17 785
rect -17 683 17 713
rect -17 679 17 683
rect -17 617 17 633
rect -17 599 17 617
rect -17 393 17 411
rect -17 377 17 393
rect -17 307 17 331
rect -17 297 17 307
rect -17 239 17 259
rect -17 225 17 239
rect -17 171 17 187
rect -17 153 17 171
rect 159 451 193 485
rect 335 853 369 857
rect 335 823 369 853
rect 335 751 369 785
rect 335 683 369 713
rect 335 679 369 683
rect 335 617 369 633
rect 335 599 369 617
rect 335 393 369 411
rect 335 377 369 393
rect 335 307 369 331
rect 335 297 369 307
rect 335 239 369 259
rect 335 225 369 239
rect 335 171 369 187
rect 335 153 369 171
rect 511 451 545 485
rect 687 853 721 857
rect 687 823 721 853
rect 687 751 721 785
rect 687 683 721 713
rect 687 679 721 683
rect 687 599 721 633
rect 687 393 721 411
rect 687 377 721 393
rect 687 307 721 331
rect 687 297 721 307
rect 687 239 721 259
rect 687 225 721 239
rect 687 171 721 187
rect 687 153 721 171
<< metal1 >>
rect -29 857 733 869
rect -29 823 -17 857
rect 17 823 335 857
rect 369 823 687 857
rect 721 823 733 857
rect -29 785 733 823
rect -29 751 -17 785
rect 17 751 335 785
rect 369 751 687 785
rect 721 751 733 785
rect -29 713 733 751
rect -29 679 -17 713
rect 17 679 335 713
rect 369 679 687 713
rect 721 679 733 713
rect -29 667 733 679
rect -29 633 733 639
rect -29 599 -17 633
rect 17 599 335 633
rect 369 599 687 633
rect 721 599 733 633
rect -29 593 733 599
rect 147 485 557 491
rect 147 451 159 485
rect 193 451 511 485
rect 545 451 557 485
rect 147 445 557 451
rect -29 411 733 417
rect -29 377 -17 411
rect 17 377 335 411
rect 369 377 687 411
rect 721 377 733 411
rect -29 371 733 377
rect -29 331 733 343
rect -29 297 -17 331
rect 17 297 335 331
rect 369 297 687 331
rect 721 297 733 331
rect -29 259 733 297
rect -29 225 -17 259
rect 17 225 335 259
rect 369 225 687 259
rect 721 225 733 259
rect -29 187 733 225
rect -29 153 -17 187
rect 17 153 335 187
rect 369 153 687 187
rect 721 153 733 187
rect -29 141 733 153
use sky130_fd_pr__model__nfet_highvoltage__example_55959141808145  sky130_fd_pr__model__nfet_highvoltage__example_55959141808145_0
timestamp 1701704242
transform 1 0 28 0 -1 319
box -1 0 649 1
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808146  sky130_fd_pr__model__pfet_highvoltage__example_55959141808146_0
timestamp 1701704242
transform 1 0 28 0 1 671
box -1 0 649 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_0
timestamp 1701704242
transform 0 -1 721 -1 0 331
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_1
timestamp 1701704242
transform 0 -1 369 -1 0 331
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_2
timestamp 1701704242
transform 0 -1 17 -1 0 331
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_3
timestamp 1701704242
transform 0 -1 369 1 0 679
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_4
timestamp 1701704242
transform 0 -1 721 1 0 679
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_5
timestamp 1701704242
transform 0 -1 17 1 0 679
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180898  sky130_fd_pr__via_l1m1__example_5595914180898_0
timestamp 1701704242
transform 1 0 511 0 1 451
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180898  sky130_fd_pr__via_l1m1__example_5595914180898_1
timestamp 1701704242
transform 1 0 159 0 1 451
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180898  sky130_fd_pr__via_l1m1__example_5595914180898_2
timestamp 1701704242
transform 1 0 -17 0 -1 633
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180898  sky130_fd_pr__via_l1m1__example_5595914180898_3
timestamp 1701704242
transform 1 0 335 0 -1 633
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180898  sky130_fd_pr__via_l1m1__example_5595914180898_4
timestamp 1701704242
transform 1 0 687 0 -1 633
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180898  sky130_fd_pr__via_l1m1__example_5595914180898_5
timestamp 1701704242
transform 1 0 335 0 -1 411
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180898  sky130_fd_pr__via_l1m1__example_5595914180898_6
timestamp 1701704242
transform 1 0 -17 0 -1 411
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180898  sky130_fd_pr__via_l1m1__example_5595914180898_7
timestamp 1701704242
transform 1 0 687 0 -1 411
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_0
timestamp 1701704242
transform -1 0 683 0 1 1303
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_1
timestamp 1701704242
transform -1 0 507 0 1 1303
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_2
timestamp 1701704242
transform -1 0 331 0 1 1303
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_3
timestamp 1701704242
transform -1 0 155 0 1 1303
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_4
timestamp 1701704242
transform -1 0 683 0 1 21
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_5
timestamp 1701704242
transform -1 0 507 0 1 21
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_6
timestamp 1701704242
transform -1 0 331 0 1 21
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_7
timestamp 1701704242
transform -1 0 155 0 1 21
box 0 0 1 1
<< labels >>
flabel metal1 s 0 667 12 869 3 FreeSans 200 0 0 0 VPWR
port 1 nsew
flabel metal1 s 0 593 12 639 3 FreeSans 200 0 0 0 VPB
port 2 nsew
flabel metal1 s 0 371 12 417 3 FreeSans 200 0 0 0 VNB
port 3 nsew
flabel metal1 s 0 141 12 343 3 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel metal1 s 692 141 704 343 3 FreeSans 200 180 0 0 VGND
port 4 nsew
flabel metal1 s 692 371 704 417 3 FreeSans 200 180 0 0 VNB
port 3 nsew
flabel metal1 s 692 593 704 639 3 FreeSans 200 180 0 0 VPB
port 2 nsew
flabel metal1 s 692 667 704 869 3 FreeSans 200 180 0 0 VPWR
port 1 nsew
flabel locali s 423 1319 457 1369 0 FreeSans 200 0 0 0 IN
port 5 nsew
flabel locali s 599 1319 633 1369 0 FreeSans 200 0 0 0 IN
port 5 nsew
flabel locali s 71 1319 105 1369 0 FreeSans 200 0 0 0 IN
port 5 nsew
flabel locali s 247 1319 281 1369 0 FreeSans 200 0 0 0 IN
port 5 nsew
flabel locali s 246 21 280 71 0 FreeSans 200 0 0 0 IN
port 5 nsew
flabel locali s 423 21 457 71 0 FreeSans 200 0 0 0 IN
port 5 nsew
flabel locali s 599 21 633 71 0 FreeSans 200 0 0 0 IN
port 5 nsew
flabel locali s 511 121 545 171 0 FreeSans 200 0 0 0 OUT
port 6 nsew
flabel locali s 159 121 193 171 0 FreeSans 200 0 0 0 OUT
port 6 nsew
flabel locali s 159 1221 193 1270 0 FreeSans 200 0 0 0 OUT
port 6 nsew
flabel locali s 511 1221 545 1270 0 FreeSans 200 0 0 0 OUT
port 6 nsew
flabel locali s 71 21 105 71 0 FreeSans 200 0 0 0 IN
port 5 nsew
<< properties >>
string GDS_END 70820006
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 70812028
<< end >>
