magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< dnwell >>
rect -336 1932 2037 4597
<< pwell >>
rect -88 4263 1789 4349
rect -88 2288 -2 4263
rect 1703 2288 1789 4263
rect -88 2202 1789 2288
<< psubdiff >>
rect -62 4289 29 4323
rect 63 4289 97 4323
rect 131 4289 165 4323
rect 199 4289 233 4323
rect 267 4289 301 4323
rect 335 4289 369 4323
rect 403 4289 437 4323
rect 471 4289 505 4323
rect 539 4289 573 4323
rect 607 4289 641 4323
rect 675 4289 709 4323
rect 743 4289 777 4323
rect 811 4289 845 4323
rect 879 4289 913 4323
rect 947 4289 981 4323
rect 1015 4289 1049 4323
rect 1083 4289 1117 4323
rect 1151 4289 1185 4323
rect 1219 4289 1253 4323
rect 1287 4289 1321 4323
rect 1355 4289 1389 4323
rect 1423 4289 1457 4323
rect 1491 4289 1525 4323
rect 1559 4289 1593 4323
rect 1627 4289 1661 4323
rect 1695 4289 1763 4323
rect -62 4255 -28 4289
rect -62 4187 -28 4221
rect 1729 4234 1763 4289
rect -62 4119 -28 4153
rect 1729 4166 1763 4200
rect -62 4051 -28 4085
rect -62 3983 -28 4017
rect -62 3915 -28 3949
rect -62 3847 -28 3881
rect 1729 4098 1763 4132
rect 1729 4030 1763 4064
rect 1729 3962 1763 3996
rect 1729 3894 1763 3928
rect 1729 3826 1763 3860
rect -62 3779 -28 3813
rect -62 3711 -28 3745
rect -62 3643 -28 3677
rect -62 3575 -28 3609
rect -62 3507 -28 3541
rect 1729 3758 1763 3792
rect 1729 3690 1763 3724
rect 1729 3622 1763 3656
rect 1729 3554 1763 3588
rect 1729 3486 1763 3520
rect -62 3439 -28 3473
rect 1729 3418 1763 3452
rect -62 3371 -28 3405
rect -62 3303 -28 3337
rect -62 3235 -28 3269
rect -62 3167 -28 3201
rect -62 3099 -28 3133
rect -62 3031 -28 3065
rect 1729 3350 1763 3384
rect 1729 3282 1763 3316
rect 1729 3214 1763 3248
rect 1729 3146 1763 3180
rect 1729 3078 1763 3112
rect -62 2963 -28 2997
rect 1729 3010 1763 3044
rect -62 2895 -28 2929
rect -62 2827 -28 2861
rect -62 2759 -28 2793
rect 1729 2942 1763 2976
rect 1729 2874 1763 2908
rect 1729 2806 1763 2840
rect 1729 2738 1763 2772
rect -62 2691 -28 2725
rect -62 2623 -28 2657
rect 1729 2670 1763 2704
rect -62 2555 -28 2589
rect -62 2487 -28 2521
rect -62 2419 -28 2453
rect -62 2351 -28 2385
rect -62 2262 -28 2317
rect 1729 2602 1763 2636
rect 1729 2534 1763 2568
rect 1729 2466 1763 2500
rect 1729 2398 1763 2432
rect 1729 2330 1763 2364
rect 1729 2262 1763 2296
rect -62 2228 6 2262
rect 40 2228 74 2262
rect 108 2228 142 2262
rect 176 2228 210 2262
rect 244 2228 278 2262
rect 312 2228 346 2262
rect 380 2228 414 2262
rect 448 2228 482 2262
rect 516 2228 550 2262
rect 584 2228 618 2262
rect 652 2228 686 2262
rect 720 2228 754 2262
rect 788 2228 822 2262
rect 856 2228 890 2262
rect 924 2228 1021 2262
rect 1055 2228 1089 2262
rect 1123 2228 1157 2262
rect 1191 2228 1225 2262
rect 1259 2228 1293 2262
rect 1327 2228 1361 2262
rect 1395 2228 1429 2262
rect 1463 2228 1497 2262
rect 1531 2228 1565 2262
rect 1599 2228 1633 2262
rect 1667 2228 1763 2262
<< psubdiffcont >>
rect 29 4289 63 4323
rect 97 4289 131 4323
rect 165 4289 199 4323
rect 233 4289 267 4323
rect 301 4289 335 4323
rect 369 4289 403 4323
rect 437 4289 471 4323
rect 505 4289 539 4323
rect 573 4289 607 4323
rect 641 4289 675 4323
rect 709 4289 743 4323
rect 777 4289 811 4323
rect 845 4289 879 4323
rect 913 4289 947 4323
rect 981 4289 1015 4323
rect 1049 4289 1083 4323
rect 1117 4289 1151 4323
rect 1185 4289 1219 4323
rect 1253 4289 1287 4323
rect 1321 4289 1355 4323
rect 1389 4289 1423 4323
rect 1457 4289 1491 4323
rect 1525 4289 1559 4323
rect 1593 4289 1627 4323
rect 1661 4289 1695 4323
rect -62 4221 -28 4255
rect -62 4153 -28 4187
rect 1729 4200 1763 4234
rect -62 4085 -28 4119
rect -62 4017 -28 4051
rect -62 3949 -28 3983
rect -62 3881 -28 3915
rect -62 3813 -28 3847
rect 1729 4132 1763 4166
rect 1729 4064 1763 4098
rect 1729 3996 1763 4030
rect 1729 3928 1763 3962
rect 1729 3860 1763 3894
rect -62 3745 -28 3779
rect 1729 3792 1763 3826
rect -62 3677 -28 3711
rect -62 3609 -28 3643
rect -62 3541 -28 3575
rect -62 3473 -28 3507
rect 1729 3724 1763 3758
rect 1729 3656 1763 3690
rect 1729 3588 1763 3622
rect 1729 3520 1763 3554
rect -62 3405 -28 3439
rect 1729 3452 1763 3486
rect -62 3337 -28 3371
rect -62 3269 -28 3303
rect -62 3201 -28 3235
rect -62 3133 -28 3167
rect -62 3065 -28 3099
rect 1729 3384 1763 3418
rect 1729 3316 1763 3350
rect 1729 3248 1763 3282
rect 1729 3180 1763 3214
rect 1729 3112 1763 3146
rect 1729 3044 1763 3078
rect -62 2997 -28 3031
rect 1729 2976 1763 3010
rect -62 2929 -28 2963
rect -62 2861 -28 2895
rect -62 2793 -28 2827
rect -62 2725 -28 2759
rect 1729 2908 1763 2942
rect 1729 2840 1763 2874
rect 1729 2772 1763 2806
rect -62 2657 -28 2691
rect 1729 2704 1763 2738
rect -62 2589 -28 2623
rect 1729 2636 1763 2670
rect -62 2521 -28 2555
rect -62 2453 -28 2487
rect -62 2385 -28 2419
rect -62 2317 -28 2351
rect 1729 2568 1763 2602
rect 1729 2500 1763 2534
rect 1729 2432 1763 2466
rect 1729 2364 1763 2398
rect 1729 2296 1763 2330
rect 6 2228 40 2262
rect 74 2228 108 2262
rect 142 2228 176 2262
rect 210 2228 244 2262
rect 278 2228 312 2262
rect 346 2228 380 2262
rect 414 2228 448 2262
rect 482 2228 516 2262
rect 550 2228 584 2262
rect 618 2228 652 2262
rect 686 2228 720 2262
rect 754 2228 788 2262
rect 822 2228 856 2262
rect 890 2228 924 2262
rect 1021 2228 1055 2262
rect 1089 2228 1123 2262
rect 1157 2228 1191 2262
rect 1225 2228 1259 2262
rect 1293 2228 1327 2262
rect 1361 2228 1395 2262
rect 1429 2228 1463 2262
rect 1497 2228 1531 2262
rect 1565 2228 1599 2262
rect 1633 2228 1667 2262
<< poly >>
rect 247 4194 535 4210
rect 247 4160 263 4194
rect 297 4160 337 4194
rect 371 4160 411 4194
rect 445 4160 485 4194
rect 519 4160 535 4194
rect 247 4144 535 4160
rect 1016 4194 1304 4210
rect 1016 4160 1032 4194
rect 1066 4160 1106 4194
rect 1140 4160 1180 4194
rect 1214 4160 1254 4194
rect 1288 4160 1304 4194
rect 1016 4144 1304 4160
rect 1134 3810 1562 3826
rect 1134 3776 1150 3810
rect 1184 3776 1222 3810
rect 1256 3776 1294 3810
rect 1328 3776 1366 3810
rect 1400 3776 1439 3810
rect 1473 3776 1512 3810
rect 1546 3776 1562 3810
rect 1134 3760 1562 3776
rect 141 3458 793 3474
rect 141 3424 157 3458
rect 191 3424 231 3458
rect 265 3424 305 3458
rect 339 3424 378 3458
rect 412 3424 451 3458
rect 485 3424 524 3458
rect 558 3424 597 3458
rect 631 3424 670 3458
rect 704 3424 743 3458
rect 777 3424 793 3458
rect 141 3408 793 3424
rect 328 3022 462 3038
rect 328 2988 344 3022
rect 378 2988 412 3022
rect 446 2988 462 3022
rect 328 2972 462 2988
rect 795 2722 929 2738
rect 795 2688 811 2722
rect 845 2688 879 2722
rect 913 2688 929 2722
rect 795 2672 929 2688
rect 1167 2672 1367 2688
rect 1167 2638 1183 2672
rect 1217 2638 1317 2672
rect 1351 2638 1367 2672
rect 1167 2622 1367 2638
rect 854 748 988 764
rect 854 714 870 748
rect 904 714 938 748
rect 972 714 988 748
rect 854 698 988 714
rect 1346 615 1412 631
rect 1346 581 1362 615
rect 1396 581 1412 615
rect 1346 547 1412 581
rect 1346 513 1362 547
rect 1396 513 1412 547
rect 1346 497 1412 513
rect 1346 229 1412 245
rect 1346 195 1362 229
rect 1396 195 1412 229
rect 1346 161 1412 195
rect 1346 127 1362 161
rect 1396 127 1412 161
rect 1346 111 1412 127
rect 447 18 581 34
rect 447 -16 463 18
rect 497 -16 531 18
rect 565 -16 581 18
rect 447 -32 581 -16
<< polycont >>
rect 263 4160 297 4194
rect 337 4160 371 4194
rect 411 4160 445 4194
rect 485 4160 519 4194
rect 1032 4160 1066 4194
rect 1106 4160 1140 4194
rect 1180 4160 1214 4194
rect 1254 4160 1288 4194
rect 1150 3776 1184 3810
rect 1222 3776 1256 3810
rect 1294 3776 1328 3810
rect 1366 3776 1400 3810
rect 1439 3776 1473 3810
rect 1512 3776 1546 3810
rect 157 3424 191 3458
rect 231 3424 265 3458
rect 305 3424 339 3458
rect 378 3424 412 3458
rect 451 3424 485 3458
rect 524 3424 558 3458
rect 597 3424 631 3458
rect 670 3424 704 3458
rect 743 3424 777 3458
rect 344 2988 378 3022
rect 412 2988 446 3022
rect 811 2688 845 2722
rect 879 2688 913 2722
rect 1183 2638 1217 2672
rect 1317 2638 1351 2672
rect 870 714 904 748
rect 938 714 972 748
rect 1362 581 1396 615
rect 1362 513 1396 547
rect 1362 195 1396 229
rect 1362 127 1396 161
rect 463 -16 497 18
rect 531 -16 565 18
<< locali >>
rect -62 4289 29 4323
rect 63 4289 97 4323
rect 131 4289 165 4323
rect 199 4289 233 4323
rect 267 4289 301 4323
rect 335 4289 369 4323
rect 403 4289 437 4323
rect 471 4289 505 4323
rect 539 4289 573 4323
rect 607 4289 641 4323
rect 675 4289 709 4323
rect 743 4289 777 4323
rect 811 4289 845 4323
rect 879 4289 913 4323
rect 947 4289 981 4323
rect 1015 4289 1049 4323
rect 1083 4289 1117 4323
rect 1151 4289 1185 4323
rect 1219 4289 1253 4323
rect 1287 4289 1321 4323
rect 1355 4289 1389 4323
rect 1423 4289 1457 4323
rect 1491 4289 1525 4323
rect 1559 4289 1593 4323
rect 1627 4289 1661 4323
rect 1695 4289 1763 4323
rect -62 4255 -28 4289
rect -62 4187 -28 4221
rect 1729 4234 1763 4289
rect 247 4160 263 4194
rect 297 4160 326 4194
rect 371 4160 398 4194
rect 445 4160 485 4194
rect 519 4160 535 4194
rect 1016 4160 1032 4194
rect 1066 4160 1106 4194
rect 1158 4160 1180 4194
rect 1230 4160 1254 4194
rect 1288 4160 1304 4194
rect 1729 4166 1763 4200
rect -62 4119 -28 4153
rect -62 4051 -28 4076
rect -62 3983 -28 4002
rect -62 3915 -28 3928
rect 134 4076 168 4110
rect 202 4076 236 4110
rect 134 4026 236 4076
rect 134 3992 168 4026
rect 202 3992 236 4026
rect 134 3942 236 3992
rect 134 3908 168 3942
rect 202 3908 236 3942
rect -62 3847 -28 3854
rect 277 3798 333 4112
rect 374 4038 408 4076
rect 449 3798 505 4112
rect 546 4076 580 4110
rect 614 4076 648 4110
rect 546 4026 648 4076
rect 546 3992 580 4026
rect 614 3992 648 4026
rect 546 3942 648 3992
rect 546 3908 580 3942
rect 614 3908 648 3942
rect 903 4076 937 4110
rect 971 4076 1005 4110
rect 903 4026 1005 4076
rect 903 3992 937 4026
rect 971 3992 1005 4026
rect 1729 4110 1763 4132
rect 1143 4042 1177 4080
rect 1315 4076 1349 4110
rect 1383 4076 1417 4110
rect 1315 4026 1417 4076
rect 903 3942 1005 3992
rect 1315 3992 1349 4026
rect 1383 3992 1417 4026
rect 903 3908 937 3942
rect 971 3908 1005 3942
rect 1057 3882 1091 3920
rect 1229 3882 1263 3920
rect 1315 3942 1417 3992
rect 1315 3908 1349 3942
rect 1383 3908 1417 3942
rect 1729 4036 1763 4064
rect 1729 3962 1763 3996
rect 1729 3894 1763 3928
rect 1729 3826 1763 3854
rect -62 3779 -28 3780
rect -62 3740 -28 3745
rect -62 3666 -28 3677
rect -62 3592 -28 3609
rect -62 3518 -28 3541
rect 88 3748 613 3798
rect 1134 3776 1150 3810
rect 1184 3776 1222 3810
rect 1256 3776 1294 3810
rect 1328 3776 1366 3810
rect 1417 3776 1439 3810
rect 1489 3776 1512 3810
rect 1546 3776 1562 3810
rect 88 3506 141 3748
rect 299 3579 405 3710
rect 333 3545 371 3579
rect 299 3508 405 3545
rect 557 3506 613 3748
rect 1729 3758 1763 3780
rect 768 3579 874 3710
rect 1729 3690 1763 3706
rect 802 3545 840 3579
rect 1089 3585 1123 3623
rect 1729 3622 1763 3632
rect 1729 3554 1763 3558
rect 768 3508 874 3545
rect 1729 3518 1763 3520
rect -62 3444 -28 3473
rect 141 3424 157 3458
rect 191 3424 231 3458
rect 265 3424 305 3458
rect 339 3424 378 3458
rect 412 3424 451 3458
rect 485 3424 523 3458
rect 558 3424 595 3458
rect 631 3424 670 3458
rect 704 3424 743 3458
rect 777 3424 793 3458
rect 1729 3444 1763 3452
rect -62 3371 -28 3405
rect -62 3303 -28 3336
rect -62 3235 -28 3262
rect -62 3167 -28 3188
rect 60 3340 231 3374
rect 60 3306 191 3340
rect 225 3306 231 3340
rect 60 3268 231 3306
rect 60 3234 191 3268
rect 225 3234 231 3268
rect 60 3172 231 3234
rect 299 3243 405 3374
rect 333 3209 371 3243
rect 299 3172 405 3209
rect 532 3346 638 3374
rect 566 3312 604 3346
rect 532 3172 638 3312
rect 768 3243 874 3374
rect 1729 3370 1763 3384
rect 1729 3296 1763 3316
rect 802 3209 840 3243
rect 768 3172 874 3209
rect 1397 3174 1431 3212
rect 1227 3120 1265 3154
rect 1573 3174 1607 3212
rect 1729 3222 1763 3248
rect 1729 3148 1763 3180
rect -62 3099 -28 3114
rect -62 3031 -28 3040
rect 1729 3078 1763 3112
rect 436 3022 474 3028
rect 328 2988 344 3022
rect 378 2994 402 3022
rect 446 2994 474 3022
rect 1729 3010 1763 3040
rect 378 2988 412 2994
rect 446 2988 462 2994
rect -62 2963 -28 2966
rect -62 2925 -28 2929
rect 717 2896 751 2934
rect 1729 2942 1763 2966
rect -62 2850 -28 2861
rect 973 2828 1007 2866
rect -62 2775 -28 2793
rect -62 2700 -28 2725
rect 464 2726 498 2764
rect 1058 2752 1168 2924
rect 1344 2812 1378 2850
rect 1729 2874 1763 2891
rect 1729 2806 1763 2816
rect 795 2688 807 2722
rect 845 2688 879 2722
rect 913 2688 929 2722
rect 1007 2710 1202 2752
rect 1729 2738 1763 2741
rect -62 2625 -28 2657
rect -62 2555 -28 2589
rect -62 2487 -28 2516
rect -62 2419 -28 2441
rect 288 2400 322 2438
rect 685 2453 791 2638
rect 719 2419 757 2453
rect -62 2351 -28 2366
rect 858 2332 967 2638
rect -62 2262 -28 2317
rect 883 2298 921 2332
rect 955 2298 967 2332
rect 1007 2610 1129 2710
rect 1729 2700 1763 2704
rect 1167 2638 1183 2672
rect 1217 2638 1253 2672
rect 1287 2638 1317 2672
rect 1359 2638 1367 2672
rect 1729 2625 1763 2636
rect 1007 2332 1082 2610
rect 1122 2465 1228 2570
rect 1156 2431 1194 2465
rect 1361 2564 1653 2570
rect 1361 2530 1364 2564
rect 1398 2530 1436 2564
rect 1470 2558 1653 2564
rect 1470 2530 1613 2558
rect 1361 2524 1613 2530
rect 1647 2524 1653 2558
rect 1361 2486 1653 2524
rect 1361 2452 1613 2486
rect 1647 2452 1653 2486
rect 1361 2436 1653 2452
rect 1729 2550 1763 2568
rect 1729 2475 1763 2500
rect 1729 2400 1763 2432
rect 1007 2298 1019 2332
rect 1053 2298 1091 2332
rect 1729 2330 1763 2364
rect 1729 2262 1763 2296
rect -62 2228 6 2262
rect 40 2228 74 2262
rect 108 2228 142 2262
rect 176 2228 210 2262
rect 244 2228 278 2262
rect 312 2228 346 2262
rect 380 2228 414 2262
rect 448 2228 482 2262
rect 516 2228 550 2262
rect 584 2228 618 2262
rect 652 2228 686 2262
rect 720 2228 754 2262
rect 788 2228 822 2262
rect 856 2228 890 2262
rect 924 2228 1021 2262
rect 1055 2228 1089 2262
rect 1123 2228 1157 2262
rect 1191 2228 1225 2262
rect 1259 2228 1293 2262
rect 1327 2228 1361 2262
rect 1395 2228 1429 2262
rect 1463 2228 1497 2262
rect 1531 2228 1565 2262
rect 1599 2228 1633 2262
rect 1667 2228 1763 2262
rect 854 748 1294 793
rect 854 714 870 748
rect 904 714 938 748
rect 972 714 1294 748
rect 854 659 1294 714
rect 408 523 442 561
rect 686 423 746 616
rect 643 389 709 423
rect 743 389 809 423
rect 609 339 843 389
rect 643 305 709 339
rect 743 305 809 339
rect 686 62 746 305
rect 889 222 950 659
rect 1160 658 1294 659
rect 1160 636 1168 658
rect 1202 624 1240 658
rect 1274 636 1294 658
rect 1362 615 1396 631
rect 990 523 1024 561
rect 1362 564 1396 581
rect 1362 547 1365 564
rect 1399 530 1449 564
rect 1483 530 1532 564
rect 1362 497 1396 513
rect 1160 389 1184 400
rect 1218 389 1256 423
rect 1290 389 1306 400
rect 1160 340 1306 389
rect 1184 339 1290 340
rect 1218 305 1256 339
rect 889 188 905 222
rect 939 188 950 222
rect 1362 229 1396 245
rect 889 150 950 188
rect 1310 165 1348 199
rect 1382 165 1396 195
rect 889 116 905 150
rect 939 116 950 150
rect 1362 161 1396 165
rect 889 102 950 116
rect 1202 82 1240 116
rect 1362 111 1396 127
rect 1436 116 1566 530
rect 1436 82 1448 116
rect 1482 82 1520 116
rect 1554 82 1566 116
rect 1436 76 1566 82
rect 447 -16 460 18
rect 497 -16 531 18
rect 566 -16 581 18
<< viali >>
rect 326 4160 337 4194
rect 337 4160 360 4194
rect 398 4160 411 4194
rect 411 4160 432 4194
rect 1124 4160 1140 4194
rect 1140 4160 1158 4194
rect 1196 4160 1214 4194
rect 1214 4160 1230 4194
rect -62 4085 -28 4110
rect -62 4076 -28 4085
rect -62 4017 -28 4036
rect -62 4002 -28 4017
rect -62 3949 -28 3962
rect -62 3928 -28 3949
rect 168 4076 202 4110
rect 168 3992 202 4026
rect 168 3908 202 3942
rect -62 3881 -28 3888
rect -62 3854 -28 3881
rect -62 3813 -28 3814
rect -62 3780 -28 3813
rect 374 4076 408 4110
rect 374 4004 408 4038
rect 580 4076 614 4110
rect 580 3992 614 4026
rect 580 3908 614 3942
rect 937 4076 971 4110
rect 937 3992 971 4026
rect 1143 4080 1177 4114
rect 1143 4008 1177 4042
rect 1349 4076 1383 4110
rect 1349 3992 1383 4026
rect 937 3908 971 3942
rect 1057 3920 1091 3954
rect 1057 3848 1091 3882
rect 1229 3920 1263 3954
rect 1349 3908 1383 3942
rect 1729 4098 1763 4110
rect 1729 4076 1763 4098
rect 1729 4030 1763 4036
rect 1729 4002 1763 4030
rect 1729 3928 1763 3962
rect 1229 3848 1263 3882
rect 1729 3860 1763 3888
rect 1729 3854 1763 3860
rect -62 3711 -28 3740
rect -62 3706 -28 3711
rect -62 3643 -28 3666
rect -62 3632 -28 3643
rect -62 3575 -28 3592
rect -62 3558 -28 3575
rect -62 3507 -28 3518
rect -62 3484 -28 3507
rect 1383 3776 1400 3810
rect 1400 3776 1417 3810
rect 1455 3776 1473 3810
rect 1473 3776 1489 3810
rect 1729 3792 1763 3814
rect 1729 3780 1763 3792
rect 299 3545 333 3579
rect 371 3545 405 3579
rect 1729 3724 1763 3740
rect 1729 3706 1763 3724
rect 768 3545 802 3579
rect 840 3545 874 3579
rect 1089 3623 1123 3657
rect 1089 3551 1123 3585
rect 1729 3656 1763 3666
rect 1729 3632 1763 3656
rect 1729 3588 1763 3592
rect 1729 3558 1763 3588
rect 1729 3486 1763 3518
rect 1729 3484 1763 3486
rect -62 3439 -28 3444
rect -62 3410 -28 3439
rect 523 3424 524 3458
rect 524 3424 557 3458
rect 595 3424 597 3458
rect 597 3424 629 3458
rect 1729 3418 1763 3444
rect 1729 3410 1763 3418
rect -62 3337 -28 3370
rect -62 3336 -28 3337
rect -62 3269 -28 3296
rect -62 3262 -28 3269
rect -62 3201 -28 3222
rect -62 3188 -28 3201
rect 191 3306 225 3340
rect 191 3234 225 3268
rect 299 3209 333 3243
rect 371 3209 405 3243
rect 532 3312 566 3346
rect 604 3312 638 3346
rect 1729 3350 1763 3370
rect 1729 3336 1763 3350
rect 1729 3282 1763 3296
rect 1729 3262 1763 3282
rect 768 3209 802 3243
rect 840 3209 874 3243
rect 1397 3212 1431 3246
rect -62 3133 -28 3148
rect -62 3114 -28 3133
rect 1193 3120 1227 3154
rect 1265 3120 1299 3154
rect 1397 3140 1431 3174
rect 1573 3212 1607 3246
rect 1573 3140 1607 3174
rect 1729 3214 1763 3222
rect 1729 3188 1763 3214
rect 1729 3146 1763 3148
rect -62 3065 -28 3074
rect -62 3040 -28 3065
rect 1729 3114 1763 3146
rect 1729 3044 1763 3074
rect 1729 3040 1763 3044
rect 402 3022 436 3028
rect -62 2997 -28 3000
rect -62 2966 -28 2997
rect 402 2994 412 3022
rect 412 2994 436 3022
rect 474 2994 508 3028
rect 1729 2976 1763 3000
rect -62 2895 -28 2925
rect -62 2891 -28 2895
rect 717 2934 751 2968
rect 1729 2966 1763 2976
rect 717 2862 751 2896
rect 973 2866 1007 2900
rect -62 2827 -28 2850
rect -62 2816 -28 2827
rect -62 2759 -28 2775
rect -62 2741 -28 2759
rect -62 2691 -28 2700
rect 464 2764 498 2798
rect 973 2794 1007 2828
rect 1729 2908 1763 2925
rect 1729 2891 1763 2908
rect 1344 2850 1378 2884
rect 1344 2778 1378 2812
rect 1729 2840 1763 2850
rect 1729 2816 1763 2840
rect 1729 2772 1763 2775
rect 464 2692 498 2726
rect -62 2666 -28 2691
rect 807 2688 811 2722
rect 811 2688 841 2722
rect 879 2688 913 2722
rect 1729 2741 1763 2772
rect -62 2623 -28 2625
rect -62 2591 -28 2623
rect -62 2521 -28 2550
rect -62 2516 -28 2521
rect -62 2453 -28 2475
rect -62 2441 -28 2453
rect -62 2385 -28 2400
rect -62 2366 -28 2385
rect 288 2438 322 2472
rect 685 2419 719 2453
rect 757 2419 791 2453
rect 288 2366 322 2400
rect 849 2298 883 2332
rect 921 2298 955 2332
rect 1253 2638 1287 2672
rect 1325 2638 1351 2672
rect 1351 2638 1359 2672
rect 1729 2670 1763 2700
rect 1729 2666 1763 2670
rect 1729 2602 1763 2625
rect 1729 2591 1763 2602
rect 1122 2431 1156 2465
rect 1194 2431 1228 2465
rect 1364 2530 1398 2564
rect 1436 2530 1470 2564
rect 1613 2524 1647 2558
rect 1613 2452 1647 2486
rect 1729 2534 1763 2550
rect 1729 2516 1763 2534
rect 1729 2466 1763 2475
rect 1729 2441 1763 2466
rect 1729 2398 1763 2400
rect 1729 2366 1763 2398
rect 1019 2298 1053 2332
rect 1091 2298 1125 2332
rect 408 561 442 595
rect 408 489 442 523
rect 609 389 643 423
rect 709 389 743 423
rect 809 389 843 423
rect 609 305 643 339
rect 709 305 743 339
rect 809 305 843 339
rect 1168 624 1202 658
rect 1240 624 1274 658
rect 990 561 1024 595
rect 990 489 1024 523
rect 1365 547 1399 564
rect 1365 530 1396 547
rect 1396 530 1399 547
rect 1449 530 1483 564
rect 1532 530 1566 564
rect 1184 389 1218 423
rect 1256 389 1290 423
rect 1184 305 1218 339
rect 1256 305 1290 339
rect 905 188 939 222
rect 1276 165 1310 199
rect 1348 195 1362 199
rect 1362 195 1382 199
rect 1348 165 1382 195
rect 905 116 939 150
rect 1168 82 1202 116
rect 1240 82 1274 116
rect 1448 82 1482 116
rect 1520 82 1554 116
rect 460 -16 463 18
rect 463 -16 494 18
rect 532 -16 565 18
rect 565 -16 566 18
<< metal1 >>
rect 314 4194 444 4200
rect 314 4160 326 4194
rect 360 4160 398 4194
rect 432 4160 444 4194
rect 314 4154 444 4160
rect 1112 4194 1242 4200
rect 1112 4160 1124 4194
rect 1158 4160 1196 4194
rect 1230 4160 1242 4194
rect 1112 4154 1242 4160
tri 1133 4122 1137 4126 se
rect 1137 4122 1183 4126
tri 1183 4122 1187 4126 sw
rect -68 4114 1769 4122
rect -68 4110 1143 4114
rect -68 4076 -62 4110
rect -28 4076 168 4110
rect 202 4076 374 4110
rect 408 4076 580 4110
rect 614 4076 937 4110
rect 971 4080 1143 4110
rect 1177 4110 1769 4114
rect 1177 4080 1349 4110
rect 971 4076 1349 4080
rect 1383 4076 1729 4110
rect 1763 4076 1769 4110
rect -68 4042 1769 4076
rect -68 4038 1143 4042
rect -68 4036 374 4038
rect -68 4002 -62 4036
rect -28 4026 374 4036
rect -28 4002 168 4026
rect -68 3992 168 4002
rect 202 4004 374 4026
rect 408 4026 1143 4038
rect 408 4004 580 4026
rect 202 3996 580 4004
rect 202 3992 300 3996
tri 300 3992 304 3996 nw
tri 364 3992 368 3996 ne
rect 368 3992 414 3996
tri 414 3992 418 3996 nw
tri 503 3992 507 3996 ne
rect 507 3992 580 3996
rect 614 3996 937 4026
rect 614 3992 687 3996
tri 687 3992 691 3996 nw
tri 860 3992 864 3996 ne
rect 864 3992 937 3996
rect 971 4008 1143 4026
rect 1177 4036 1769 4042
rect 1177 4026 1729 4036
rect 1177 4008 1349 4026
rect 971 3996 1349 4008
rect 971 3992 1036 3996
tri 1036 3992 1040 3996 nw
tri 1280 3992 1284 3996 ne
rect 1284 3992 1349 3996
rect 1383 4002 1729 4026
rect 1763 4002 1769 4036
rect 1383 3996 1769 4002
rect 1383 3992 1423 3996
rect -68 3962 270 3992
tri 270 3962 300 3992 nw
tri 507 3962 537 3992 ne
rect 537 3962 657 3992
tri 657 3962 687 3992 nw
tri 864 3967 889 3992 ne
rect 889 3967 1011 3992
tri 1011 3967 1036 3992 nw
tri 1284 3967 1309 3992 ne
tri 889 3962 894 3967 ne
rect 894 3962 1011 3967
rect -68 3928 -62 3962
rect -28 3954 262 3962
tri 262 3954 270 3962 nw
tri 537 3959 540 3962 ne
rect -28 3942 250 3954
tri 250 3942 262 3954 nw
rect 540 3942 654 3962
tri 654 3959 657 3962 nw
tri 894 3959 897 3962 ne
rect -28 3928 168 3942
rect -68 3908 168 3928
rect 202 3908 242 3942
tri 242 3934 250 3942 nw
rect -68 3896 242 3908
rect 540 3908 580 3942
rect 614 3908 654 3942
rect 540 3896 654 3908
rect 897 3942 1011 3962
rect 897 3908 937 3942
rect 971 3908 1011 3942
rect 897 3896 1011 3908
rect 1051 3954 1269 3966
rect 1051 3920 1057 3954
rect 1091 3920 1229 3954
rect 1263 3920 1269 3954
rect -68 3888 234 3896
tri 234 3888 242 3896 nw
rect -68 3854 -62 3888
rect -28 3882 228 3888
tri 228 3882 234 3888 nw
rect 1051 3882 1269 3920
rect 1309 3942 1423 3992
tri 1423 3967 1452 3996 nw
tri 1680 3967 1709 3996 ne
rect 1709 3967 1769 3996
tri 1709 3962 1714 3967 ne
rect 1714 3962 1769 3967
tri 1714 3959 1717 3962 ne
rect 1717 3959 1729 3962
tri 1717 3953 1723 3959 ne
rect 1309 3908 1349 3942
rect 1383 3908 1423 3942
rect 1309 3896 1423 3908
rect 1723 3928 1729 3959
rect 1763 3928 1769 3962
rect -28 3854 194 3882
rect -68 3848 194 3854
tri 194 3848 228 3882 nw
rect 1051 3848 1057 3882
rect 1091 3848 1229 3882
rect 1263 3848 1269 3882
rect -68 3814 160 3848
tri 160 3814 194 3848 nw
rect 1051 3836 1269 3848
tri 1168 3816 1188 3836 ne
rect 1188 3816 1269 3836
rect 1723 3888 1769 3928
rect 1723 3854 1729 3888
rect 1763 3854 1769 3888
tri 1188 3814 1190 3816 ne
rect 1190 3814 1269 3816
rect -68 3780 -62 3814
rect -28 3810 156 3814
tri 156 3810 160 3814 nw
tri 1190 3810 1194 3814 ne
rect 1194 3810 1269 3814
rect -28 3780 122 3810
rect -68 3776 122 3780
tri 122 3776 156 3810 nw
tri 1194 3781 1223 3810 ne
rect -68 3740 95 3776
tri 95 3749 122 3776 nw
rect -68 3706 -62 3740
rect -28 3706 95 3740
rect -68 3666 95 3706
rect -68 3632 -62 3666
rect -28 3632 95 3666
rect -68 3592 95 3632
rect 1083 3657 1129 3669
rect 1083 3623 1089 3657
rect 1123 3623 1129 3657
tri 1053 3592 1083 3622 se
rect 1083 3592 1129 3623
rect -68 3558 -62 3592
rect -28 3558 95 3592
tri 1046 3585 1053 3592 se
rect 1053 3585 1129 3592
rect -68 3518 95 3558
rect 287 3579 1089 3585
rect 287 3545 299 3579
rect 333 3545 371 3579
rect 405 3545 768 3579
rect 802 3545 840 3579
rect 874 3551 1089 3579
rect 1123 3551 1129 3585
rect 874 3545 1129 3551
rect 287 3539 1129 3545
rect -68 3484 -62 3518
rect -28 3484 95 3518
rect -68 3444 95 3484
rect -68 3410 -62 3444
rect -28 3410 95 3444
rect 511 3458 641 3464
rect 511 3424 523 3458
rect 557 3424 595 3458
rect 629 3424 641 3458
rect 511 3418 641 3424
rect -68 3370 95 3410
tri 1201 3370 1223 3392 se
rect 1223 3370 1269 3810
rect 1371 3810 1501 3816
rect 1371 3776 1383 3810
rect 1417 3776 1455 3810
rect 1489 3776 1501 3810
rect 1371 3770 1501 3776
rect 1723 3814 1769 3854
rect 1723 3780 1729 3814
rect 1763 3780 1769 3814
rect -68 3336 -62 3370
rect -28 3336 95 3370
tri 1183 3352 1201 3370 se
rect 1201 3352 1269 3370
rect -68 3296 95 3336
rect -68 3262 -62 3296
rect -28 3262 95 3296
rect -68 3222 95 3262
rect 185 3346 1269 3352
rect 185 3340 532 3346
rect 185 3306 191 3340
rect 225 3312 532 3340
rect 566 3312 604 3346
rect 638 3312 1269 3346
rect 225 3306 1269 3312
rect 1723 3740 1769 3780
rect 1723 3706 1729 3740
rect 1763 3706 1769 3740
rect 1723 3666 1769 3706
rect 1723 3632 1729 3666
rect 1763 3632 1769 3666
rect 1723 3592 1769 3632
rect 1723 3558 1729 3592
rect 1763 3558 1769 3592
rect 1723 3518 1769 3558
rect 1723 3484 1729 3518
rect 1763 3484 1769 3518
rect 1723 3444 1769 3484
rect 1723 3410 1729 3444
rect 1763 3410 1769 3444
rect 1723 3370 1769 3410
rect 1723 3336 1729 3370
rect 1763 3336 1769 3370
rect 185 3296 258 3306
tri 258 3296 268 3306 nw
rect 1723 3296 1769 3336
rect 185 3268 231 3296
tri 231 3269 258 3296 nw
rect 185 3234 191 3268
rect 225 3234 231 3268
rect 1723 3262 1729 3296
rect 1763 3262 1769 3296
tri 1382 3249 1391 3258 se
rect 1391 3249 1437 3258
rect 185 3222 231 3234
rect 287 3246 1437 3249
rect 287 3243 1397 3246
rect -68 3188 -62 3222
rect -28 3188 95 3222
rect 287 3209 299 3243
rect 333 3209 371 3243
rect 405 3209 768 3243
rect 802 3209 840 3243
rect 874 3212 1397 3243
rect 1431 3212 1437 3246
rect 874 3209 1437 3212
rect 287 3203 1437 3209
tri 1357 3188 1372 3203 ne
rect 1372 3188 1437 3203
rect -68 3148 95 3188
tri 1372 3174 1386 3188 ne
rect 1386 3174 1437 3188
tri 1386 3169 1391 3174 ne
rect -68 3114 -62 3148
rect -28 3114 95 3148
rect 1181 3154 1311 3160
rect 1181 3120 1193 3154
rect 1227 3120 1265 3154
rect 1299 3140 1311 3154
tri 1311 3140 1328 3157 sw
rect 1391 3140 1397 3174
rect 1431 3140 1437 3174
rect 1299 3128 1328 3140
tri 1328 3128 1340 3140 sw
rect 1391 3128 1437 3140
rect 1567 3246 1613 3258
rect 1567 3212 1573 3246
rect 1607 3212 1613 3246
rect 1567 3174 1613 3212
rect 1567 3140 1573 3174
rect 1607 3140 1613 3174
rect 1299 3120 1340 3128
rect 1181 3114 1340 3120
tri 1340 3114 1354 3128 sw
rect -68 3074 95 3114
tri 1288 3104 1298 3114 ne
rect 1298 3104 1354 3114
tri 1354 3104 1364 3114 sw
tri 1298 3094 1308 3104 ne
rect 1308 3094 1364 3104
tri 1308 3074 1328 3094 ne
rect 1328 3074 1364 3094
tri 1364 3074 1394 3104 sw
rect -68 3040 -62 3074
rect -28 3040 95 3074
tri 1328 3061 1341 3074 ne
rect 1341 3061 1394 3074
tri 1394 3061 1407 3074 sw
rect 1567 3061 1613 3140
rect 1723 3222 1769 3262
rect 1723 3188 1729 3222
rect 1763 3188 1769 3222
rect 1723 3148 1769 3188
rect 1723 3114 1729 3148
rect 1763 3114 1769 3148
rect 1723 3074 1769 3114
tri 1613 3061 1625 3073 sw
rect -68 3000 95 3040
rect 675 3060 1255 3061
tri 1255 3060 1256 3061 sw
tri 1341 3060 1342 3061 ne
rect 1342 3060 1407 3061
tri 1407 3060 1408 3061 sw
rect 1567 3060 1625 3061
tri 1625 3060 1626 3061 sw
rect 675 3040 1256 3060
tri 1256 3040 1276 3060 sw
tri 1342 3040 1362 3060 ne
rect 1362 3040 1408 3060
tri 1408 3040 1428 3060 sw
rect 1567 3053 1626 3060
tri 1567 3040 1580 3053 ne
rect 1580 3040 1626 3053
tri 1626 3040 1646 3060 sw
rect 1723 3040 1729 3074
rect 1763 3040 1769 3074
rect 675 3038 1276 3040
tri 1276 3038 1278 3040 sw
tri 1362 3038 1364 3040 ne
rect 1364 3038 1428 3040
tri 1428 3038 1430 3040 sw
tri 1580 3038 1582 3040 ne
rect 1582 3038 1646 3040
rect -68 2966 -62 3000
rect -28 2994 95 3000
rect 390 3028 520 3034
tri 95 2994 100 2999 sw
rect 390 2994 402 3028
rect 436 2994 474 3028
rect 508 2994 520 3028
tri 662 3000 675 3013 se
rect 675 3000 1278 3038
tri 1278 3000 1316 3038 sw
tri 1364 3000 1402 3038 ne
rect 1402 3033 1430 3038
tri 1430 3033 1435 3038 sw
tri 1582 3033 1587 3038 ne
rect 1587 3033 1646 3038
tri 1646 3033 1653 3040 sw
rect 1402 3013 1435 3033
tri 1435 3013 1455 3033 sw
tri 1587 3013 1607 3033 ne
rect 1402 3000 1455 3013
tri 1455 3000 1468 3013 sw
rect -28 2968 100 2994
tri 100 2968 126 2994 sw
rect 390 2988 520 2994
tri 650 2988 662 3000 se
rect 662 2988 1316 3000
tri 630 2968 650 2988 se
rect 650 2972 1316 2988
tri 1316 2972 1344 3000 sw
tri 1402 2972 1430 3000 ne
rect 1430 2972 1468 3000
tri 1468 2972 1496 3000 sw
rect 650 2968 1344 2972
rect -28 2966 126 2968
rect -68 2952 126 2966
tri 126 2952 142 2968 sw
tri 614 2952 630 2968 se
rect 630 2952 717 2968
rect -68 2934 717 2952
rect 751 2966 1344 2968
tri 1344 2966 1350 2972 sw
tri 1430 2966 1436 2972 ne
rect 1436 2966 1496 2972
tri 1496 2966 1502 2972 sw
rect 751 2959 1350 2966
rect 751 2952 840 2959
tri 840 2952 847 2959 nw
tri 1213 2952 1220 2959 ne
rect 1220 2952 1350 2959
rect 751 2934 813 2952
rect -68 2925 813 2934
tri 813 2925 840 2952 nw
tri 1220 2925 1247 2952 ne
rect 1247 2925 1350 2952
tri 1350 2925 1391 2966 sw
tri 1436 2925 1477 2966 ne
rect 1477 2925 1502 2966
tri 1502 2925 1543 2966 sw
rect -68 2891 -62 2925
rect -28 2916 804 2925
tri 804 2916 813 2925 nw
tri 1247 2916 1256 2925 ne
rect 1256 2916 1391 2925
tri 1391 2916 1400 2925 sw
rect -28 2900 788 2916
tri 788 2900 804 2916 nw
tri 1256 2912 1260 2916 ne
rect 1260 2912 1400 2916
rect 967 2900 1013 2912
rect -28 2896 786 2900
tri 786 2898 788 2900 nw
rect -28 2891 717 2896
rect -68 2862 717 2891
rect 751 2862 786 2896
rect -68 2850 786 2862
rect 967 2866 973 2900
rect 1007 2866 1013 2900
tri 1260 2898 1274 2912 ne
rect 1274 2898 1400 2912
tri 1477 2906 1496 2925 ne
rect 1496 2906 1543 2925
tri 1543 2906 1562 2925 sw
tri 1274 2891 1281 2898 ne
rect 1281 2891 1400 2898
tri 1496 2891 1511 2906 ne
rect 1511 2891 1562 2906
tri 1281 2884 1288 2891 ne
rect 1288 2884 1400 2891
tri 1511 2886 1516 2891 ne
rect -68 2816 -62 2850
rect -28 2828 120 2850
tri 120 2828 142 2850 nw
tri 954 2828 967 2841 se
rect 967 2828 1013 2866
tri 1288 2860 1312 2884 ne
rect -28 2816 95 2828
rect -68 2775 95 2816
tri 95 2803 120 2828 nw
tri 936 2810 954 2828 se
rect 954 2810 973 2828
rect -68 2741 -62 2775
rect -28 2741 95 2775
rect -68 2700 95 2741
rect -68 2666 -62 2700
rect -28 2666 95 2700
rect 458 2798 973 2810
rect 458 2764 464 2798
rect 498 2794 973 2798
rect 1007 2794 1013 2828
rect 498 2764 1013 2794
rect 1312 2850 1344 2884
rect 1378 2850 1400 2884
rect 1312 2812 1400 2850
rect 1312 2778 1344 2812
rect 1378 2778 1400 2812
rect 1312 2766 1400 2778
rect 458 2741 512 2764
tri 512 2741 535 2764 nw
tri 936 2741 959 2764 ne
rect 959 2741 1013 2764
rect 458 2726 504 2741
tri 504 2733 512 2741 nw
tri 959 2733 967 2741 ne
rect 458 2692 464 2726
rect 498 2692 504 2726
rect 458 2680 504 2692
rect 795 2722 925 2728
rect 795 2688 807 2722
rect 841 2688 879 2722
rect 913 2688 925 2722
rect 795 2682 925 2688
rect 967 2707 1013 2741
tri 1013 2707 1024 2718 sw
rect 967 2700 1024 2707
tri 1024 2700 1031 2707 sw
tri 1509 2700 1516 2707 se
rect 1516 2700 1562 2891
rect 967 2698 1031 2700
tri 1031 2698 1033 2700 sw
tri 1507 2698 1509 2700 se
rect 1509 2698 1562 2700
tri 967 2682 983 2698 ne
rect 983 2682 1033 2698
tri 1033 2682 1049 2698 sw
tri 1491 2682 1507 2698 se
rect 1507 2682 1562 2698
tri 806 2680 808 2682 ne
rect 808 2680 904 2682
tri 808 2672 816 2680 ne
rect 816 2672 904 2680
tri 904 2672 914 2682 nw
tri 983 2678 987 2682 ne
rect 987 2678 1049 2682
tri 1049 2678 1053 2682 sw
tri 1487 2678 1491 2682 se
rect 1491 2678 1562 2682
tri 987 2672 993 2678 ne
rect 993 2672 1562 2678
rect -68 2625 95 2666
tri 816 2651 837 2672 ne
rect -68 2591 -62 2625
rect -28 2591 95 2625
rect -68 2550 95 2591
rect -68 2516 -62 2550
rect -28 2516 95 2550
rect 837 2591 883 2672
tri 883 2651 904 2672 nw
tri 993 2651 1014 2672 ne
rect 1014 2651 1253 2672
tri 1014 2638 1027 2651 ne
rect 1027 2638 1253 2651
rect 1287 2638 1325 2672
rect 1359 2638 1562 2672
tri 1027 2632 1033 2638 ne
rect 1033 2632 1562 2638
tri 1487 2625 1494 2632 ne
rect 1494 2625 1562 2632
tri 1494 2603 1516 2625 ne
tri 883 2591 893 2601 sw
rect 837 2570 893 2591
tri 893 2570 914 2591 sw
rect 837 2564 1482 2570
rect 837 2530 1364 2564
rect 1398 2530 1436 2564
rect 1470 2530 1482 2564
rect 837 2524 1482 2530
rect -68 2484 95 2516
rect -68 2475 1240 2484
rect -68 2441 -62 2475
rect -28 2472 1240 2475
rect -28 2441 288 2472
rect -68 2438 288 2441
rect 322 2465 1240 2472
rect 322 2453 1122 2465
rect 322 2438 685 2453
rect -68 2419 685 2438
rect 719 2419 757 2453
rect 791 2431 1122 2453
rect 1156 2431 1194 2465
rect 1228 2431 1240 2465
rect 791 2419 1240 2431
rect -68 2400 1240 2419
rect -68 2366 -62 2400
rect -28 2370 288 2400
rect -28 2366 107 2370
tri 107 2366 111 2370 nw
tri 266 2366 270 2370 ne
rect 270 2366 288 2370
rect 322 2370 1240 2400
rect 322 2366 340 2370
tri 340 2366 344 2370 nw
rect -68 2354 95 2366
tri 95 2354 107 2366 nw
tri 270 2354 282 2366 ne
rect 282 2354 328 2366
tri 328 2354 340 2366 nw
rect 837 2332 967 2338
rect 837 2298 849 2332
rect 883 2298 921 2332
rect 955 2298 967 2332
rect 837 2292 967 2298
rect 1007 2332 1137 2338
rect 1007 2298 1019 2332
rect 1053 2298 1091 2332
rect 1125 2298 1137 2332
rect 1007 2292 1137 2298
tri 842 2262 872 2292 ne
rect 872 2287 938 2292
tri 938 2287 943 2292 nw
tri 1029 2287 1034 2292 ne
rect 1034 2287 1100 2292
rect 872 2282 933 2287
tri 933 2282 938 2287 nw
tri 1034 2282 1039 2287 ne
rect 1039 2282 1100 2287
rect 872 2277 928 2282
tri 928 2277 933 2282 nw
tri 1039 2277 1044 2282 ne
rect 1044 2277 1100 2282
rect 872 2272 923 2277
tri 923 2272 928 2277 nw
tri 1044 2272 1049 2277 ne
rect 1049 2272 1100 2277
tri 869 624 872 627 se
rect 872 624 918 2272
tri 918 2267 923 2272 nw
tri 1049 2267 1054 2272 ne
tri 1034 2044 1054 2064 se
rect 1054 2044 1100 2272
tri 1100 2267 1125 2292 nw
tri 1030 2040 1034 2044 se
rect 1034 2040 1096 2044
tri 1096 2040 1100 2044 nw
tri 852 607 869 624 se
rect 869 607 918 624
rect 402 595 448 607
tri 840 595 852 607 se
rect 852 595 906 607
tri 906 595 918 607 nw
tri 984 1994 1030 2040 se
rect 984 595 1030 1994
tri 1030 1974 1096 2040 nw
tri 1460 664 1516 720 se
rect 1516 700 1562 2625
rect 1516 664 1526 700
tri 1526 664 1562 700 nw
rect 1607 2558 1653 3033
rect 1607 2524 1613 2558
rect 1647 2524 1653 2558
rect 1607 2486 1653 2524
rect 1607 2452 1613 2486
rect 1647 2452 1653 2486
rect 1156 658 1480 664
rect 1156 624 1168 658
rect 1202 624 1240 658
rect 1274 624 1480 658
rect 1156 618 1480 624
tri 1480 618 1526 664 nw
rect 402 561 408 595
rect 442 585 448 595
tri 837 592 840 595 se
rect 840 592 896 595
tri 448 585 455 592 sw
tri 830 585 837 592 se
rect 837 585 896 592
tri 896 585 906 595 nw
rect 442 565 455 585
tri 455 565 475 585 sw
tri 810 565 830 585 se
rect 830 565 872 585
rect 442 561 872 565
tri 872 561 896 585 nw
rect 984 561 990 595
rect 1024 561 1030 595
tri 1578 570 1607 599 se
rect 1607 571 1653 2452
rect 1723 3000 1769 3040
rect 1723 2966 1729 3000
rect 1763 2966 1769 3000
rect 1723 2925 1769 2966
rect 1723 2891 1729 2925
rect 1763 2891 1769 2925
rect 1723 2850 1769 2891
rect 1723 2816 1729 2850
rect 1763 2816 1769 2850
rect 1723 2775 1769 2816
rect 1723 2741 1729 2775
rect 1763 2741 1769 2775
rect 1723 2700 1769 2741
rect 1723 2666 1729 2700
rect 1763 2666 1769 2700
rect 1723 2625 1769 2666
rect 1723 2591 1729 2625
rect 1763 2591 1769 2625
rect 1723 2550 1769 2591
rect 1723 2516 1729 2550
rect 1763 2516 1769 2550
rect 1723 2475 1769 2516
rect 1723 2441 1729 2475
rect 1763 2441 1769 2475
rect 1723 2400 1769 2441
rect 1723 2366 1729 2400
rect 1763 2366 1769 2400
rect 1723 2354 1769 2366
rect 1607 570 1652 571
tri 1652 570 1653 571 nw
rect 402 530 841 561
tri 841 530 872 561 nw
rect 402 523 834 530
tri 834 523 841 530 nw
rect 984 523 1030 561
rect 1353 564 1606 570
rect 1353 530 1365 564
rect 1399 530 1449 564
rect 1483 530 1532 564
rect 1566 530 1606 564
rect 1353 524 1606 530
tri 1606 524 1652 570 nw
rect 402 489 408 523
rect 442 519 830 523
tri 830 519 834 523 nw
rect 442 489 448 519
tri 448 492 475 519 nw
rect 402 477 448 489
rect 984 489 990 523
rect 1024 489 1030 523
rect 984 477 1030 489
rect 264 423 1652 429
rect 264 389 609 423
rect 643 389 709 423
rect 743 389 809 423
rect 843 389 1184 423
rect 1218 389 1256 423
rect 1290 389 1652 423
rect 264 339 1652 389
rect 264 305 609 339
rect 643 305 709 339
rect 743 305 809 339
rect 843 305 1184 339
rect 1218 305 1256 339
rect 1290 305 1652 339
rect 264 299 1652 305
rect 899 222 945 234
rect 899 188 905 222
rect 939 205 945 222
tri 945 205 972 232 sw
rect 939 199 1394 205
rect 939 188 1276 199
rect 899 165 1276 188
rect 1310 165 1348 199
rect 1382 165 1394 199
rect 899 159 1394 165
rect 899 150 945 159
rect 899 116 905 150
rect 939 116 945 150
tri 945 132 972 159 nw
tri 1078 116 1084 122 se
rect 1084 116 1566 122
rect 899 104 945 116
tri 1066 104 1078 116 se
rect 1078 104 1168 116
tri 1044 82 1066 104 se
rect 1066 82 1168 104
rect 1202 82 1240 116
rect 1274 82 1448 116
rect 1482 82 1520 116
rect 1554 82 1566 116
tri 1038 76 1044 82 se
rect 1044 76 1566 82
tri 1006 44 1038 76 se
rect 1038 44 1072 76
tri 1072 44 1104 76 nw
tri 986 24 1006 44 se
rect 1006 24 1052 44
tri 1052 24 1072 44 nw
rect 448 18 1006 24
rect 448 -16 460 18
rect 494 -16 532 18
rect 566 -16 1006 18
rect 448 -22 1006 -16
tri 1006 -22 1052 24 nw
use nfet_CDNS_52468879185512  nfet_CDNS_52468879185512_0
timestamp 1701704242
transform -1 0 1562 0 1 3128
box -79 -32 199 632
use nfet_CDNS_52468879185512  nfet_CDNS_52468879185512_1
timestamp 1701704242
transform -1 0 1254 0 1 3128
box -79 -32 199 632
use nfet_CDNS_52468879185512  nfet_CDNS_52468879185512_2
timestamp 1701704242
transform 1 0 333 0 1 2340
box -79 -32 199 632
use nfet_CDNS_52468879185793  nfet_CDNS_52468879185793_0
timestamp 1701704242
transform 1 0 141 0 -1 3706
box -79 -32 731 232
use nfet_CDNS_52468879185793  nfet_CDNS_52468879185793_1
timestamp 1701704242
transform 1 0 141 0 1 3176
box -79 -32 731 232
use nfet_CDNS_52468879185796  nfet_CDNS_52468879185796_0
timestamp 1701704242
transform 1 0 762 0 -1 2920
box -79 -32 279 182
use nfet_CDNS_52468879185796  nfet_CDNS_52468879185796_1
timestamp 1701704242
transform 1 0 1167 0 1 2440
box -79 -32 279 182
use nfet_CDNS_52468879185797  nfet_CDNS_52468879185797_0
timestamp 1701704242
transform -1 0 1333 0 -1 2920
box -79 -32 199 232
use nfet_CDNS_52468879185797  nfet_CDNS_52468879185797_1
timestamp 1701704242
transform 1 0 802 0 1 2440
box -79 -32 199 232
use nfet_CDNS_52468879185915  nfet_CDNS_52468879185915_0
timestamp 1701704242
transform 1 0 1016 0 1 3912
box -151 -32 439 232
use nfet_CDNS_52468879185915  nfet_CDNS_52468879185915_1
timestamp 1701704242
transform 1 0 247 0 1 3912
box -151 -32 439 232
use pfet_CDNS_52468879185911  pfet_CDNS_52468879185911_0
timestamp 1701704242
transform 0 1 1164 -1 0 227
box -266 -66 219 216
use pfet_CDNS_52468879185911  pfet_CDNS_52468879185911_1
timestamp 1701704242
transform 0 1 1164 1 0 513
box -266 -66 219 216
use pfet_CDNS_52468879185913  pfet_CDNS_52468879185913_0
timestamp 1701704242
transform -1 0 573 0 1 66
box -266 -66 239 666
use pfet_CDNS_52468879185913  pfet_CDNS_52468879185913_1
timestamp 1701704242
transform 1 0 859 0 1 66
box -266 -66 239 666
<< labels >>
flabel metal1 s 1409 3770 1477 3816 0 FreeSans 500 0 0 0 hld_h_n
port 1 nsew
flabel metal1 s 1152 4154 1211 4200 0 FreeSans 500 0 0 0 in
port 2 nsew
flabel metal1 s 359 4154 411 4200 0 FreeSans 500 0 0 0 in_n
port 3 nsew
flabel metal1 s 432 2988 489 3034 0 FreeSans 500 0 0 0 rst_h
port 4 nsew
flabel metal1 s 976 300 1090 428 0 FreeSans 500 0 0 0 vdda
port 5 nsew
flabel metal1 s 553 3418 603 3464 0 FreeSans 500 0 0 0 vpwr
port 6 nsew
flabel metal1 s 713 4016 820 4111 0 FreeSans 500 0 0 0 vssa
port 7 nsew
flabel metal1 s 872 1429 918 1486 0 FreeSans 500 90 0 0 out_h
port 8 nsew
flabel metal1 s 984 1433 1030 1486 0 FreeSans 500 90 0 0 out_h_n
port 9 nsew
flabel metal1 s 1539 1436 1539 1436 0 FreeSans 500 90 0 0 fbk
flabel metal1 s 1629 1435 1629 1435 0 FreeSans 500 90 0 0 fbk_n
<< properties >>
string GDS_END 80732718
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 80698482
string path 24.675 56.125 43.650 56.125 43.650 107.650 -1.125 107.650 -1.125 56.125 24.675 56.125 
<< end >>
