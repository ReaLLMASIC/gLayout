magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< poly >>
rect -50 50 0 66
rect -50 16 -34 50
rect -50 0 0 16
rect 800 50 850 66
rect 834 16 850 50
rect 800 0 850 16
<< polycont >>
rect -34 16 0 50
rect 800 16 834 50
<< npolyres >>
rect 0 0 800 66
<< locali >>
rect -34 50 0 66
rect -34 0 0 16
rect 800 50 834 66
rect 800 0 834 16
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_0
timestamp 1701704242
transform -1 0 16 0 1 0
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_1
timestamp 1701704242
transform 1 0 784 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 87732146
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 87731712
<< end >>
