magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< obsli1 >>
rect -1208 6870 1508 7182
rect -1208 -894 -896 6870
rect 0 0 300 6000
rect -189 -651 489 -649
rect -190 -894 489 -651
rect 1196 -894 1508 6870
rect -1208 -1182 1508 -894
<< obsm1 >>
rect -1208 6683 1508 7182
rect -1208 6450 -623 6683
tri -623 6450 -390 6683 nw
tri 689 6450 922 6683 ne
rect 922 6450 1508 6683
rect -1208 -450 -710 6450
tri -710 6363 -623 6450 nw
tri -449 6374 -373 6450 se
rect -373 6374 674 6450
tri 674 6374 750 6450 sw
tri -710 -450 -623 -363 sw
rect -449 -374 750 6374
tri 922 6362 1010 6450 ne
tri -449 -386 -437 -374 ne
rect -437 -386 738 -374
tri 738 -386 750 -374 nw
tri -437 -450 -373 -386 ne
rect -373 -450 674 -386
tri 674 -450 738 -386 nw
tri 924 -450 1010 -364 se
rect 1010 -450 1508 6450
rect -1208 -684 -623 -450
tri -623 -684 -389 -450 sw
tri 690 -684 924 -450 se
rect 924 -684 1508 -450
rect -1208 -1182 1508 -684
<< obsm2 >>
rect -1208 6683 1508 7182
rect -1208 6433 -640 6683
tri -640 6433 -390 6683 nw
tri 689 6450 922 6683 ne
rect 922 6450 1508 6683
tri -390 6433 -373 6450 se
rect -373 6433 674 6450
rect -1208 -450 -710 6433
tri -710 6363 -640 6433 nw
tri -449 6374 -390 6433 se
rect -390 6374 674 6433
tri 674 6374 750 6450 sw
tri -710 -450 -623 -363 sw
rect -449 -374 750 6374
tri 922 6362 1010 6450 ne
tri -449 -388 -435 -374 ne
rect -435 -388 736 -374
tri 736 -388 750 -374 nw
tri -435 -450 -373 -388 ne
rect -373 -450 674 -388
tri 674 -450 736 -388 nw
tri 924 -450 1010 -364 se
rect 1010 -450 1508 6450
rect -1208 -684 -623 -450
tri -623 -684 -389 -450 sw
tri 690 -684 924 -450 se
rect 924 -684 1508 -450
rect -1208 -1182 1508 -684
<< obsm3 >>
rect -1208 6683 1508 7182
rect -1208 6433 -640 6683
tri -640 6433 -390 6683 nw
tri 689 6450 922 6683 ne
rect 922 6450 1508 6683
tri -390 6433 -373 6450 se
rect -373 6433 674 6450
rect -1208 -450 -710 6433
tri -710 6363 -640 6433 nw
tri -449 6374 -390 6433 se
rect -390 6374 674 6433
tri 674 6374 750 6450 sw
tri -710 -450 -623 -363 sw
rect -449 -374 750 6374
tri 922 6362 1010 6450 ne
tri -449 -392 -431 -374 ne
rect -431 -392 732 -374
tri 732 -392 750 -374 nw
tri -431 -450 -373 -392 ne
rect -373 -450 674 -392
tri 674 -450 732 -392 nw
tri 924 -450 1010 -364 se
rect 1010 -450 1508 6450
rect -1208 -684 -623 -450
tri -623 -684 -389 -450 sw
tri 690 -684 924 -450 se
rect 924 -684 1508 -450
rect -1208 -1182 1508 -684
<< obsm4 >>
rect -1208 6683 1508 7182
rect -1208 6433 -640 6683
tri -640 6433 -390 6683 nw
tri 689 6450 922 6683 ne
rect 922 6450 1508 6683
tri -390 6433 -373 6450 se
rect -373 6433 674 6450
rect -1208 -450 -710 6433
tri -710 6363 -640 6433 nw
tri -449 6374 -390 6433 se
rect -390 6374 674 6433
tri 674 6374 750 6450 sw
tri -710 -450 -623 -363 sw
rect -449 -374 750 6374
tri 922 6362 1010 6450 ne
tri -449 -450 -373 -374 ne
rect -373 -450 674 -374
tri 674 -450 750 -374 nw
tri 924 -450 1010 -364 se
rect 1010 -450 1508 6450
rect -1208 -684 -623 -450
tri -623 -684 -389 -450 sw
tri 690 -684 924 -450 se
rect 924 -684 1508 -450
rect -1208 -1182 1508 -684
<< obsm5 >>
rect -1208 5182 1508 7182
rect -958 818 1258 5182
rect -1208 -1182 1508 818
<< properties >>
string FIXED_BBOX -1208 -1182 1508 7182
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 3906134
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 3132498
<< end >>
