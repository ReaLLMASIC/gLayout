magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< metal3 >>
rect 0 470 224 476
rect 0 0 224 6
<< via3 >>
rect 0 6 224 470
<< metal4 >>
rect -1 470 225 471
rect -1 6 0 470
rect 224 6 225 470
rect -1 5 225 6
<< properties >>
string GDS_END 88494566
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 88493282
<< end >>
