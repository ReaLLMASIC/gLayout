magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< nwell >>
rect 6326 18415 7817 19733
rect 6910 17883 7817 18415
rect 7565 14183 7817 17883
rect 6818 2410 7046 3057
rect 7517 2410 7817 7960
<< pwell >>
rect 2564 27439 8028 27933
rect 3706 24321 6218 24543
rect 7057 23272 7211 27439
rect 6029 22472 8028 23272
rect 2803 13289 6140 13393
rect 6338 12516 6424 14090
rect 7278 12516 7364 13952
rect 6338 12430 7654 12516
rect 3089 10752 4618 10838
rect 4962 10654 6261 10740
rect 3196 9743 6465 9852
rect 6691 8411 6777 11087
rect 7045 14 8028 2336
<< mvpsubdiff >>
rect 2590 27873 2624 27907
rect 2658 27873 2693 27907
rect 2727 27873 2762 27907
rect 2796 27873 2831 27907
rect 2865 27873 2900 27907
rect 2934 27873 2969 27907
rect 3003 27873 3038 27907
rect 2590 27839 3038 27873
rect 2590 27805 2624 27839
rect 2658 27805 2693 27839
rect 2727 27805 2762 27839
rect 2796 27805 2831 27839
rect 2865 27805 2900 27839
rect 2934 27805 2969 27839
rect 3003 27805 3038 27839
rect 2590 27771 3038 27805
rect 2590 27737 2624 27771
rect 2658 27737 2693 27771
rect 2727 27737 2762 27771
rect 2796 27737 2831 27771
rect 2865 27737 2900 27771
rect 2934 27737 2969 27771
rect 3003 27737 3038 27771
rect 2590 27703 3038 27737
rect 2590 27669 2624 27703
rect 2658 27669 2693 27703
rect 2727 27669 2762 27703
rect 2796 27669 2831 27703
rect 2865 27669 2900 27703
rect 2934 27669 2969 27703
rect 3003 27669 3038 27703
rect 2590 27635 3038 27669
rect 2590 27601 2624 27635
rect 2658 27601 2693 27635
rect 2727 27601 2762 27635
rect 2796 27601 2831 27635
rect 2865 27601 2900 27635
rect 2934 27601 2969 27635
rect 3003 27601 3038 27635
rect 2590 27567 3038 27601
rect 2590 27533 2624 27567
rect 2658 27533 2693 27567
rect 2727 27533 2762 27567
rect 2796 27533 2831 27567
rect 2865 27533 2900 27567
rect 2934 27533 2969 27567
rect 3003 27533 3038 27567
rect 2590 27499 3038 27533
rect 2590 27465 2624 27499
rect 2658 27465 2693 27499
rect 2727 27465 2762 27499
rect 2796 27465 2831 27499
rect 2865 27465 2900 27499
rect 2934 27465 2969 27499
rect 3003 27465 3038 27499
rect 7968 27465 8002 27907
rect 7083 27291 7185 27397
rect 7117 27257 7151 27291
rect 7083 27151 7185 27257
rect 7117 27117 7151 27151
rect 7083 27011 7185 27117
rect 7117 26977 7151 27011
rect 7083 26871 7185 26977
rect 7117 26837 7151 26871
rect 7083 26731 7185 26837
rect 7117 26697 7151 26731
rect 7083 26591 7185 26697
rect 7117 26557 7151 26591
rect 7083 26451 7185 26557
rect 7117 26417 7151 26451
rect 7083 26311 7185 26417
rect 7117 26277 7151 26311
rect 7083 26171 7185 26277
rect 7117 26137 7151 26171
rect 7083 26031 7185 26137
rect 7117 25997 7151 26031
rect 7083 25891 7185 25997
rect 7117 25857 7151 25891
rect 7083 25751 7185 25857
rect 7117 25717 7151 25751
rect 7083 25611 7185 25717
rect 7117 25577 7151 25611
rect 7083 25471 7185 25577
rect 7117 25437 7151 25471
rect 7083 25330 7185 25437
rect 7117 25296 7151 25330
rect 7083 25189 7185 25296
rect 7117 25155 7151 25189
rect 7083 25048 7185 25155
rect 7117 25014 7151 25048
rect 7083 24907 7185 25014
rect 7117 24873 7151 24907
rect 7083 24766 7185 24873
rect 7117 24732 7151 24766
rect 7083 24625 7185 24732
rect 7117 24591 7151 24625
rect 3732 24483 3766 24517
rect 3800 24483 3836 24517
rect 3870 24483 3906 24517
rect 3940 24483 3976 24517
rect 4010 24483 4046 24517
rect 4080 24483 4116 24517
rect 4150 24483 4186 24517
rect 4220 24483 4256 24517
rect 4290 24483 4326 24517
rect 4360 24483 4396 24517
rect 4430 24483 4466 24517
rect 4500 24483 4536 24517
rect 4570 24483 4606 24517
rect 4640 24483 4675 24517
rect 4709 24483 4744 24517
rect 4778 24483 4813 24517
rect 4847 24483 4882 24517
rect 4916 24483 4951 24517
rect 4985 24483 5020 24517
rect 5054 24483 5089 24517
rect 5123 24483 5158 24517
rect 5192 24483 5227 24517
rect 5261 24483 5296 24517
rect 5330 24483 5365 24517
rect 5399 24483 5434 24517
rect 5468 24483 5503 24517
rect 5537 24483 5572 24517
rect 5606 24483 5641 24517
rect 5675 24483 5710 24517
rect 5744 24483 5779 24517
rect 5813 24483 5848 24517
rect 5882 24483 5917 24517
rect 5951 24483 5986 24517
rect 6020 24483 6055 24517
rect 6089 24483 6124 24517
rect 6158 24483 6192 24517
rect 3732 24449 6192 24483
rect 3732 24415 3766 24449
rect 3800 24415 3836 24449
rect 3870 24415 3906 24449
rect 3940 24415 3976 24449
rect 4010 24415 4046 24449
rect 4080 24415 4116 24449
rect 4150 24415 4186 24449
rect 4220 24415 4256 24449
rect 4290 24415 4326 24449
rect 4360 24415 4396 24449
rect 4430 24415 4466 24449
rect 4500 24415 4536 24449
rect 4570 24415 4606 24449
rect 4640 24415 4675 24449
rect 4709 24415 4744 24449
rect 4778 24415 4813 24449
rect 4847 24415 4882 24449
rect 4916 24415 4951 24449
rect 4985 24415 5020 24449
rect 5054 24415 5089 24449
rect 5123 24415 5158 24449
rect 5192 24415 5227 24449
rect 5261 24415 5296 24449
rect 5330 24415 5365 24449
rect 5399 24415 5434 24449
rect 5468 24415 5503 24449
rect 5537 24415 5572 24449
rect 5606 24415 5641 24449
rect 5675 24415 5710 24449
rect 5744 24415 5779 24449
rect 5813 24415 5848 24449
rect 5882 24415 5917 24449
rect 5951 24415 5986 24449
rect 6020 24415 6055 24449
rect 6089 24415 6124 24449
rect 6158 24415 6192 24449
rect 3732 24381 6192 24415
rect 3732 24347 3766 24381
rect 3800 24347 3836 24381
rect 3870 24347 3906 24381
rect 3940 24347 3976 24381
rect 4010 24347 4046 24381
rect 4080 24347 4116 24381
rect 4150 24347 4186 24381
rect 4220 24347 4256 24381
rect 4290 24347 4326 24381
rect 4360 24347 4396 24381
rect 4430 24347 4466 24381
rect 4500 24347 4536 24381
rect 4570 24347 4606 24381
rect 4640 24347 4675 24381
rect 4709 24347 4744 24381
rect 4778 24347 4813 24381
rect 4847 24347 4882 24381
rect 4916 24347 4951 24381
rect 4985 24347 5020 24381
rect 5054 24347 5089 24381
rect 5123 24347 5158 24381
rect 5192 24347 5227 24381
rect 5261 24347 5296 24381
rect 5330 24347 5365 24381
rect 5399 24347 5434 24381
rect 5468 24347 5503 24381
rect 5537 24347 5572 24381
rect 5606 24347 5641 24381
rect 5675 24347 5710 24381
rect 5744 24347 5779 24381
rect 5813 24347 5848 24381
rect 5882 24347 5917 24381
rect 5951 24347 5986 24381
rect 6020 24347 6055 24381
rect 6089 24347 6124 24381
rect 6158 24347 6192 24381
rect 7083 24484 7185 24591
rect 7117 24450 7151 24484
rect 7083 24343 7185 24450
rect 7117 24309 7151 24343
rect 7083 24202 7185 24309
rect 7117 24168 7151 24202
rect 7083 24061 7185 24168
rect 7117 24027 7151 24061
rect 7083 23920 7185 24027
rect 7117 23886 7151 23920
rect 7083 23779 7185 23886
rect 7117 23745 7151 23779
rect 7083 23638 7185 23745
rect 7117 23604 7151 23638
rect 7083 23497 7185 23604
rect 7117 23463 7151 23497
rect 7083 23356 7185 23463
rect 7117 23322 7151 23356
rect 7083 23246 7185 23322
rect 6055 23212 6089 23246
rect 6123 23212 6230 23246
rect 6264 23212 6372 23246
rect 6406 23212 6514 23246
rect 6548 23212 6656 23246
rect 6690 23212 6798 23246
rect 6832 23212 6940 23246
rect 6974 23212 7082 23246
rect 7116 23212 7224 23246
rect 7258 23212 7366 23246
rect 7400 23212 7508 23246
rect 7542 23212 7650 23246
rect 7684 23212 7792 23246
rect 7826 23212 7934 23246
rect 7968 23212 8002 23246
rect 6055 23144 8002 23212
rect 6055 23110 6089 23144
rect 6123 23110 6230 23144
rect 6264 23110 6372 23144
rect 6406 23110 6514 23144
rect 6548 23110 6656 23144
rect 6690 23110 6798 23144
rect 6832 23110 6940 23144
rect 6974 23110 7082 23144
rect 7116 23110 7224 23144
rect 7258 23110 7366 23144
rect 7400 23110 7508 23144
rect 7542 23110 7650 23144
rect 7684 23110 7792 23144
rect 7826 23110 7934 23144
rect 7968 23110 8002 23144
rect 6055 23042 8002 23110
rect 6055 23008 6089 23042
rect 6123 23008 6230 23042
rect 6264 23008 6372 23042
rect 6406 23008 6514 23042
rect 6548 23008 6656 23042
rect 6690 23008 6798 23042
rect 6832 23008 6940 23042
rect 6974 23008 7082 23042
rect 7116 23008 7224 23042
rect 7258 23008 7366 23042
rect 7400 23008 7508 23042
rect 7542 23008 7650 23042
rect 7684 23008 7792 23042
rect 7826 23008 7934 23042
rect 7968 23008 8002 23042
rect 6055 22940 8002 23008
rect 6055 22906 6089 22940
rect 6123 22906 6230 22940
rect 6264 22906 6372 22940
rect 6406 22906 6514 22940
rect 6548 22906 6656 22940
rect 6690 22906 6798 22940
rect 6832 22906 6940 22940
rect 6974 22906 7082 22940
rect 7116 22906 7224 22940
rect 7258 22906 7366 22940
rect 7400 22906 7508 22940
rect 7542 22906 7650 22940
rect 7684 22906 7792 22940
rect 7826 22906 7934 22940
rect 7968 22906 8002 22940
rect 6055 22838 8002 22906
rect 6055 22804 6089 22838
rect 6123 22804 6230 22838
rect 6264 22804 6372 22838
rect 6406 22804 6514 22838
rect 6548 22804 6656 22838
rect 6690 22804 6798 22838
rect 6832 22804 6940 22838
rect 6974 22804 7082 22838
rect 7116 22804 7224 22838
rect 7258 22804 7366 22838
rect 7400 22804 7508 22838
rect 7542 22804 7650 22838
rect 7684 22804 7792 22838
rect 7826 22804 7934 22838
rect 7968 22804 8002 22838
rect 6055 22736 8002 22804
rect 6055 22702 6089 22736
rect 6123 22702 6230 22736
rect 6264 22702 6372 22736
rect 6406 22702 6514 22736
rect 6548 22702 6656 22736
rect 6690 22702 6798 22736
rect 6832 22702 6940 22736
rect 6974 22702 7082 22736
rect 7116 22702 7224 22736
rect 7258 22702 7366 22736
rect 7400 22702 7508 22736
rect 7542 22702 7650 22736
rect 7684 22702 7792 22736
rect 7826 22702 7934 22736
rect 7968 22702 8002 22736
rect 6055 22634 8002 22702
rect 6055 22600 6089 22634
rect 6123 22600 6230 22634
rect 6264 22600 6372 22634
rect 6406 22600 6514 22634
rect 6548 22600 6656 22634
rect 6690 22600 6798 22634
rect 6832 22600 6940 22634
rect 6974 22600 7082 22634
rect 7116 22600 7224 22634
rect 7258 22600 7366 22634
rect 7400 22600 7508 22634
rect 7542 22600 7650 22634
rect 7684 22600 7792 22634
rect 7826 22600 7934 22634
rect 7968 22600 8002 22634
rect 6055 22532 8002 22600
rect 6055 22498 6089 22532
rect 6123 22498 6230 22532
rect 6264 22498 6372 22532
rect 6406 22498 6514 22532
rect 6548 22498 6656 22532
rect 6690 22498 6798 22532
rect 6832 22498 6940 22532
rect 6974 22498 7082 22532
rect 7116 22498 7224 22532
rect 7258 22498 7366 22532
rect 7400 22498 7508 22532
rect 7542 22498 7650 22532
rect 7684 22498 7792 22532
rect 7826 22498 7934 22532
rect 7968 22498 8002 22532
rect 6364 14040 6398 14064
rect 6364 13971 6398 14006
rect 6364 13902 6398 13937
rect 6364 13833 6398 13868
rect 6364 13764 6398 13799
rect 6364 13695 6398 13730
rect 6364 13625 6398 13661
rect 6364 13555 6398 13591
rect 6364 13485 6398 13521
rect 6364 13415 6398 13451
rect 7304 13902 7338 13926
rect 7304 13834 7338 13868
rect 7304 13766 7338 13800
rect 7304 13698 7338 13732
rect 7304 13630 7338 13664
rect 6364 13345 6398 13381
rect 6364 13275 6398 13311
rect 6364 13205 6398 13241
rect 6364 13135 6398 13171
rect 6364 13065 6398 13101
rect 6364 12995 6398 13031
rect 6364 12925 6398 12961
rect 6364 12855 6398 12891
rect 6364 12785 6398 12821
rect 7304 13562 7338 13596
rect 7304 13494 7338 13528
rect 7304 13426 7338 13460
rect 7304 13358 7338 13392
rect 7304 13289 7338 13324
rect 7304 13220 7338 13255
rect 7304 13151 7338 13186
rect 7304 13082 7338 13117
rect 7304 13013 7338 13048
rect 7304 12944 7338 12979
rect 7304 12875 7338 12910
rect 6364 12715 6398 12751
rect 6364 12645 6398 12681
rect 7304 12806 7338 12841
rect 7304 12737 7338 12772
rect 7304 12679 7338 12703
rect 6364 12587 6398 12611
rect 6364 12456 6388 12490
rect 6422 12456 6458 12490
rect 6492 12456 6528 12490
rect 6562 12456 6598 12490
rect 6632 12456 6668 12490
rect 6702 12456 6738 12490
rect 6772 12456 6808 12490
rect 6842 12456 6878 12490
rect 6912 12456 6948 12490
rect 6982 12456 7018 12490
rect 7052 12456 7087 12490
rect 7121 12456 7156 12490
rect 7190 12456 7225 12490
rect 7259 12456 7294 12490
rect 7328 12456 7363 12490
rect 7397 12456 7432 12490
rect 7466 12456 7501 12490
rect 7535 12456 7570 12490
rect 7604 12456 7628 12490
rect 6717 11037 6751 11061
rect 6717 10968 6751 11003
rect 6717 10899 6751 10934
rect 6717 10830 6751 10865
rect 3115 10778 3139 10812
rect 3173 10778 3209 10812
rect 3243 10778 3279 10812
rect 3313 10778 3349 10812
rect 3383 10778 3419 10812
rect 3453 10778 3489 10812
rect 3523 10778 3559 10812
rect 3593 10778 3629 10812
rect 3663 10778 3699 10812
rect 3733 10778 3769 10812
rect 3803 10778 3839 10812
rect 3873 10778 3909 10812
rect 3943 10778 3979 10812
rect 4013 10778 4049 10812
rect 4083 10778 4119 10812
rect 4153 10778 4189 10812
rect 4223 10778 4258 10812
rect 4292 10778 4327 10812
rect 4361 10778 4396 10812
rect 4430 10778 4465 10812
rect 4499 10778 4534 10812
rect 4568 10778 4592 10812
rect 6717 10761 6751 10796
rect 4988 10680 5012 10714
rect 5046 10680 5081 10714
rect 5115 10680 5150 10714
rect 5184 10680 5219 10714
rect 5253 10680 5288 10714
rect 5322 10680 5357 10714
rect 5391 10680 5426 10714
rect 5460 10680 5495 10714
rect 5529 10680 5564 10714
rect 5598 10680 5633 10714
rect 5667 10680 5701 10714
rect 5735 10680 5769 10714
rect 5803 10680 5837 10714
rect 5871 10680 5905 10714
rect 5939 10680 5973 10714
rect 6007 10680 6041 10714
rect 6075 10680 6109 10714
rect 6143 10680 6177 10714
rect 6211 10680 6235 10714
rect 6717 10692 6751 10727
rect 6717 10623 6751 10658
rect 6717 10554 6751 10589
rect 6717 10485 6751 10520
rect 6717 10416 6751 10451
rect 6717 10347 6751 10382
rect 6717 10278 6751 10313
rect 6717 10209 6751 10244
rect 6717 10140 6751 10175
rect 6717 10071 6751 10106
rect 6717 10002 6751 10037
rect 6717 9933 6751 9968
rect 6717 9864 6751 9899
rect 6717 9795 6751 9830
rect 6717 9726 6751 9761
rect 6717 9657 6751 9692
rect 6717 9588 6751 9623
rect 6717 9519 6751 9554
rect 6717 9450 6751 9485
rect 6717 9381 6751 9416
rect 6717 9312 6751 9347
rect 6717 9243 6751 9278
rect 6717 9175 6751 9209
rect 6717 9107 6751 9141
rect 6717 9039 6751 9073
rect 6717 8971 6751 9005
rect 6717 8903 6751 8937
rect 6717 8835 6751 8869
rect 6717 8767 6751 8801
rect 6717 8699 6751 8733
rect 6717 8631 6751 8665
rect 6717 8563 6751 8597
rect 6717 8495 6751 8529
rect 6717 8437 6751 8461
rect 7071 2276 8002 2310
rect 7105 2242 7139 2276
rect 7173 2242 7207 2276
rect 7241 2242 7275 2276
rect 7309 2242 7343 2276
rect 7377 2242 7411 2276
rect 7445 2242 7479 2276
rect 7513 2242 7547 2276
rect 7581 2242 7615 2276
rect 7649 2242 7683 2276
rect 7717 2242 7751 2276
rect 7785 2242 7819 2276
rect 7853 2242 7887 2276
rect 7921 2242 8002 2276
rect 7071 2207 8002 2242
rect 7105 2173 7139 2207
rect 7173 2173 7207 2207
rect 7241 2173 7275 2207
rect 7309 2173 7343 2207
rect 7377 2173 7411 2207
rect 7445 2173 7479 2207
rect 7513 2173 7547 2207
rect 7581 2173 7615 2207
rect 7649 2173 7683 2207
rect 7717 2173 7751 2207
rect 7785 2173 7819 2207
rect 7853 2173 7887 2207
rect 7921 2173 8002 2207
rect 7071 2138 8002 2173
rect 7105 2104 7139 2138
rect 7173 2104 7207 2138
rect 7241 2104 7275 2138
rect 7309 2104 7343 2138
rect 7377 2104 7411 2138
rect 7445 2104 7479 2138
rect 7513 2104 7547 2138
rect 7581 2104 7615 2138
rect 7649 2104 7683 2138
rect 7717 2104 7751 2138
rect 7785 2104 7819 2138
rect 7853 2104 7887 2138
rect 7921 2104 8002 2138
rect 7071 2068 8002 2104
rect 7105 2034 7139 2068
rect 7173 2034 7207 2068
rect 7241 2034 7275 2068
rect 7309 2034 7343 2068
rect 7377 2034 7411 2068
rect 7445 2034 7479 2068
rect 7513 2034 7547 2068
rect 7581 2034 7615 2068
rect 7649 2034 7683 2068
rect 7717 2034 7751 2068
rect 7785 2034 7819 2068
rect 7853 2034 7887 2068
rect 7921 2034 8002 2068
rect 7071 1998 8002 2034
rect 7105 1964 7139 1998
rect 7173 1964 7207 1998
rect 7241 1964 7275 1998
rect 7309 1964 7343 1998
rect 7377 1964 7411 1998
rect 7445 1964 7479 1998
rect 7513 1964 7547 1998
rect 7581 1964 7615 1998
rect 7649 1964 7683 1998
rect 7717 1964 7751 1998
rect 7785 1964 7819 1998
rect 7853 1964 7887 1998
rect 7921 1964 8002 1998
rect 7071 1928 8002 1964
rect 7105 1894 7139 1928
rect 7173 1894 7207 1928
rect 7241 1894 7275 1928
rect 7309 1894 7343 1928
rect 7377 1894 7411 1928
rect 7445 1894 7479 1928
rect 7513 1894 7547 1928
rect 7581 1894 7615 1928
rect 7649 1894 7683 1928
rect 7717 1894 7751 1928
rect 7785 1894 7819 1928
rect 7853 1894 7887 1928
rect 7921 1894 8002 1928
rect 7071 1858 8002 1894
rect 7105 1824 7139 1858
rect 7173 1824 7207 1858
rect 7241 1824 7275 1858
rect 7309 1824 7343 1858
rect 7377 1824 7411 1858
rect 7445 1824 7479 1858
rect 7513 1824 7547 1858
rect 7581 1824 7615 1858
rect 7649 1824 7683 1858
rect 7717 1824 7751 1858
rect 7785 1824 7819 1858
rect 7853 1824 7887 1858
rect 7921 1824 8002 1858
rect 7071 1788 8002 1824
rect 7105 1754 7139 1788
rect 7173 1754 7207 1788
rect 7241 1754 7275 1788
rect 7309 1754 7343 1788
rect 7377 1754 7411 1788
rect 7445 1754 7479 1788
rect 7513 1754 7547 1788
rect 7581 1754 7615 1788
rect 7649 1754 7683 1788
rect 7717 1754 7751 1788
rect 7785 1754 7819 1788
rect 7853 1754 7887 1788
rect 7921 1754 8002 1788
rect 7071 1718 8002 1754
rect 7105 1684 7139 1718
rect 7173 1684 7207 1718
rect 7241 1684 7275 1718
rect 7309 1684 7343 1718
rect 7377 1684 7411 1718
rect 7445 1684 7479 1718
rect 7513 1684 7547 1718
rect 7581 1684 7615 1718
rect 7649 1684 7683 1718
rect 7717 1684 7751 1718
rect 7785 1684 7819 1718
rect 7853 1684 7887 1718
rect 7921 1684 8002 1718
rect 7071 1648 8002 1684
rect 7105 1614 7139 1648
rect 7173 1614 7207 1648
rect 7241 1614 7275 1648
rect 7309 1614 7343 1648
rect 7377 1614 7411 1648
rect 7445 1614 7479 1648
rect 7513 1614 7547 1648
rect 7581 1614 7615 1648
rect 7649 1614 7683 1648
rect 7717 1614 7751 1648
rect 7785 1614 7819 1648
rect 7853 1614 7887 1648
rect 7921 1614 8002 1648
rect 7071 1578 8002 1614
rect 7105 1544 7139 1578
rect 7173 1544 7207 1578
rect 7241 1544 7275 1578
rect 7309 1544 7343 1578
rect 7377 1544 7411 1578
rect 7445 1544 7479 1578
rect 7513 1544 7547 1578
rect 7581 1544 7615 1578
rect 7649 1544 7683 1578
rect 7717 1544 7751 1578
rect 7785 1544 7819 1578
rect 7853 1544 7887 1578
rect 7921 1544 8002 1578
rect 7071 1508 8002 1544
rect 7105 1474 7139 1508
rect 7173 1474 7207 1508
rect 7241 1474 7275 1508
rect 7309 1474 7343 1508
rect 7377 1474 7411 1508
rect 7445 1474 7479 1508
rect 7513 1474 7547 1508
rect 7581 1474 7615 1508
rect 7649 1474 7683 1508
rect 7717 1474 7751 1508
rect 7785 1474 7819 1508
rect 7853 1474 7887 1508
rect 7921 1474 8002 1508
rect 7071 1438 8002 1474
rect 7105 1404 7139 1438
rect 7173 1404 7207 1438
rect 7241 1404 7275 1438
rect 7309 1404 7343 1438
rect 7377 1404 7411 1438
rect 7445 1404 7479 1438
rect 7513 1404 7547 1438
rect 7581 1404 7615 1438
rect 7649 1404 7683 1438
rect 7717 1404 7751 1438
rect 7785 1404 7819 1438
rect 7853 1404 7887 1438
rect 7921 1404 8002 1438
rect 7071 1368 8002 1404
rect 7105 1334 7139 1368
rect 7173 1334 7207 1368
rect 7241 1334 7275 1368
rect 7309 1334 7343 1368
rect 7377 1334 7411 1368
rect 7445 1334 7479 1368
rect 7513 1334 7547 1368
rect 7581 1334 7615 1368
rect 7649 1334 7683 1368
rect 7717 1334 7751 1368
rect 7785 1334 7819 1368
rect 7853 1334 7887 1368
rect 7921 1334 8002 1368
rect 7071 1298 8002 1334
rect 7105 1264 7139 1298
rect 7173 1264 7207 1298
rect 7241 1264 7275 1298
rect 7309 1264 7343 1298
rect 7377 1264 7411 1298
rect 7445 1264 7479 1298
rect 7513 1264 7547 1298
rect 7581 1264 7615 1298
rect 7649 1264 7683 1298
rect 7717 1264 7751 1298
rect 7785 1264 7819 1298
rect 7853 1264 7887 1298
rect 7921 1264 8002 1298
rect 7071 1228 8002 1264
rect 7105 1194 7139 1228
rect 7173 1194 7207 1228
rect 7241 1194 7275 1228
rect 7309 1194 7343 1228
rect 7377 1194 7411 1228
rect 7445 1194 7479 1228
rect 7513 1194 7547 1228
rect 7581 1194 7615 1228
rect 7649 1194 7683 1228
rect 7717 1194 7751 1228
rect 7785 1194 7819 1228
rect 7853 1194 7887 1228
rect 7921 1194 8002 1228
rect 7071 1158 8002 1194
rect 7105 1124 7139 1158
rect 7173 1124 7207 1158
rect 7241 1124 7275 1158
rect 7309 1124 7343 1158
rect 7377 1124 7411 1158
rect 7445 1124 7479 1158
rect 7513 1124 7547 1158
rect 7581 1124 7615 1158
rect 7649 1124 7683 1158
rect 7717 1124 7751 1158
rect 7785 1124 7819 1158
rect 7853 1124 7887 1158
rect 7921 1124 8002 1158
rect 7071 1088 8002 1124
rect 7105 1054 7139 1088
rect 7173 1054 7207 1088
rect 7241 1054 7275 1088
rect 7309 1054 7343 1088
rect 7377 1054 7411 1088
rect 7445 1054 7479 1088
rect 7513 1054 7547 1088
rect 7581 1054 7615 1088
rect 7649 1054 7683 1088
rect 7717 1054 7751 1088
rect 7785 1054 7819 1088
rect 7853 1054 7887 1088
rect 7921 1054 8002 1088
rect 7071 1018 8002 1054
rect 7105 984 7139 1018
rect 7173 984 7207 1018
rect 7241 984 7275 1018
rect 7309 984 7343 1018
rect 7377 984 7411 1018
rect 7445 984 7479 1018
rect 7513 984 7547 1018
rect 7581 984 7615 1018
rect 7649 984 7683 1018
rect 7717 984 7751 1018
rect 7785 984 7819 1018
rect 7853 984 7887 1018
rect 7921 984 8002 1018
rect 7071 948 8002 984
rect 7105 914 7139 948
rect 7173 914 7207 948
rect 7241 914 7275 948
rect 7309 914 7343 948
rect 7377 914 7411 948
rect 7445 914 7479 948
rect 7513 914 7547 948
rect 7581 914 7615 948
rect 7649 914 7683 948
rect 7717 914 7751 948
rect 7785 914 7819 948
rect 7853 914 7887 948
rect 7921 914 8002 948
rect 7071 878 8002 914
rect 7105 844 7139 878
rect 7173 844 7207 878
rect 7241 844 7275 878
rect 7309 844 7343 878
rect 7377 844 7411 878
rect 7445 844 7479 878
rect 7513 844 7547 878
rect 7581 844 7615 878
rect 7649 844 7683 878
rect 7717 844 7751 878
rect 7785 844 7819 878
rect 7853 844 7887 878
rect 7921 844 8002 878
rect 7071 808 8002 844
rect 7105 774 7139 808
rect 7173 774 7207 808
rect 7241 774 7275 808
rect 7309 774 7343 808
rect 7377 774 7411 808
rect 7445 774 7479 808
rect 7513 774 7547 808
rect 7581 774 7615 808
rect 7649 774 7683 808
rect 7717 774 7751 808
rect 7785 774 7819 808
rect 7853 774 7887 808
rect 7921 774 8002 808
rect 7071 738 8002 774
rect 7105 704 7139 738
rect 7173 704 7207 738
rect 7241 704 7275 738
rect 7309 704 7343 738
rect 7377 704 7411 738
rect 7445 704 7479 738
rect 7513 704 7547 738
rect 7581 704 7615 738
rect 7649 704 7683 738
rect 7717 704 7751 738
rect 7785 704 7819 738
rect 7853 704 7887 738
rect 7921 704 8002 738
rect 7071 668 8002 704
rect 7105 634 7139 668
rect 7173 634 7207 668
rect 7241 634 7275 668
rect 7309 634 7343 668
rect 7377 634 7411 668
rect 7445 634 7479 668
rect 7513 634 7547 668
rect 7581 634 7615 668
rect 7649 634 7683 668
rect 7717 634 7751 668
rect 7785 634 7819 668
rect 7853 634 7887 668
rect 7921 634 8002 668
rect 7071 598 8002 634
rect 7105 564 7139 598
rect 7173 564 7207 598
rect 7241 564 7275 598
rect 7309 564 7343 598
rect 7377 564 7411 598
rect 7445 564 7479 598
rect 7513 564 7547 598
rect 7581 564 7615 598
rect 7649 564 7683 598
rect 7717 564 7751 598
rect 7785 564 7819 598
rect 7853 564 7887 598
rect 7921 564 8002 598
rect 7071 528 8002 564
rect 7105 494 7139 528
rect 7173 494 7207 528
rect 7241 494 7275 528
rect 7309 494 7343 528
rect 7377 494 7411 528
rect 7445 494 7479 528
rect 7513 494 7547 528
rect 7581 494 7615 528
rect 7649 494 7683 528
rect 7717 494 7751 528
rect 7785 494 7819 528
rect 7853 494 7887 528
rect 7921 494 8002 528
rect 7071 458 8002 494
rect 7105 424 7139 458
rect 7173 424 7207 458
rect 7241 424 7275 458
rect 7309 424 7343 458
rect 7377 424 7411 458
rect 7445 424 7479 458
rect 7513 424 7547 458
rect 7581 424 7615 458
rect 7649 424 7683 458
rect 7717 424 7751 458
rect 7785 424 7819 458
rect 7853 424 7887 458
rect 7921 424 8002 458
rect 7071 388 8002 424
rect 7105 354 7139 388
rect 7173 354 7207 388
rect 7241 354 7275 388
rect 7309 354 7343 388
rect 7377 354 7411 388
rect 7445 354 7479 388
rect 7513 354 7547 388
rect 7581 354 7615 388
rect 7649 354 7683 388
rect 7717 354 7751 388
rect 7785 354 7819 388
rect 7853 354 7887 388
rect 7921 354 8002 388
rect 7071 318 8002 354
rect 7105 284 7139 318
rect 7173 284 7207 318
rect 7241 284 7275 318
rect 7309 284 7343 318
rect 7377 284 7411 318
rect 7445 284 7479 318
rect 7513 284 7547 318
rect 7581 284 7615 318
rect 7649 284 7683 318
rect 7717 284 7751 318
rect 7785 284 7819 318
rect 7853 284 7887 318
rect 7921 284 8002 318
rect 7071 248 8002 284
rect 7105 214 7139 248
rect 7173 214 7207 248
rect 7241 214 7275 248
rect 7309 214 7343 248
rect 7377 214 7411 248
rect 7445 214 7479 248
rect 7513 214 7547 248
rect 7581 214 7615 248
rect 7649 214 7683 248
rect 7717 214 7751 248
rect 7785 214 7819 248
rect 7853 214 7887 248
rect 7921 214 8002 248
rect 7071 178 8002 214
rect 7105 144 7139 178
rect 7173 144 7207 178
rect 7241 144 7275 178
rect 7309 144 7343 178
rect 7377 144 7411 178
rect 7445 144 7479 178
rect 7513 144 7547 178
rect 7581 144 7615 178
rect 7649 144 7683 178
rect 7717 144 7751 178
rect 7785 144 7819 178
rect 7853 144 7887 178
rect 7921 144 8002 178
rect 7071 108 8002 144
rect 7105 74 7139 108
rect 7173 74 7207 108
rect 7241 74 7275 108
rect 7309 74 7343 108
rect 7377 74 7411 108
rect 7445 74 7479 108
rect 7513 74 7547 108
rect 7581 74 7615 108
rect 7649 74 7683 108
rect 7717 74 7751 108
rect 7785 74 7819 108
rect 7853 74 7887 108
rect 7921 74 8002 108
rect 7071 40 8002 74
<< mvnsubdiff >>
rect 7716 19622 7750 19666
rect 7716 19554 7750 19588
rect 7716 19486 7750 19520
rect 7716 19418 7750 19452
rect 7716 19350 7750 19384
rect 7716 19282 7750 19316
rect 7716 19214 7750 19248
rect 7716 19146 7750 19180
rect 7716 19078 7750 19112
rect 7716 19010 7750 19044
rect 7716 18942 7750 18976
rect 7716 18874 7750 18908
rect 7716 18806 7750 18840
rect 7716 18738 7750 18772
rect 7716 18670 7750 18704
rect 7716 18602 7750 18636
rect 7716 18534 7750 18568
rect 7716 18466 7750 18500
rect 7716 18398 7750 18432
rect 7716 18330 7750 18364
rect 7716 18262 7750 18296
rect 7716 18194 7750 18228
rect 7716 18126 7750 18160
rect 7716 18058 7750 18092
rect 7716 17990 7750 18024
rect 7716 17922 7750 17956
rect 7716 17854 7750 17888
rect 7716 17786 7750 17820
rect 7716 17718 7750 17752
rect 7716 17650 7750 17684
rect 7716 17582 7750 17616
rect 7716 17514 7750 17548
rect 7716 17446 7750 17480
rect 7716 17378 7750 17412
rect 7716 17310 7750 17344
rect 7716 17242 7750 17276
rect 7716 17174 7750 17208
rect 7716 17106 7750 17140
rect 7716 17038 7750 17072
rect 7716 16970 7750 17004
rect 7716 16902 7750 16936
rect 7716 16834 7750 16868
rect 7716 16766 7750 16800
rect 7716 16698 7750 16732
rect 7716 16630 7750 16664
rect 7716 16562 7750 16596
rect 7716 16494 7750 16528
rect 7716 16426 7750 16460
rect 7716 16358 7750 16392
rect 7716 16290 7750 16324
rect 7716 16222 7750 16256
rect 7716 16154 7750 16188
rect 7716 16086 7750 16120
rect 7716 16018 7750 16052
rect 7716 15950 7750 15984
rect 7716 15882 7750 15916
rect 7716 15814 7750 15848
rect 7716 15746 7750 15780
rect 7716 15678 7750 15712
rect 7716 15610 7750 15644
rect 7716 15542 7750 15576
rect 7716 15474 7750 15508
rect 7716 15406 7750 15440
rect 7716 15338 7750 15372
rect 7716 15270 7750 15304
rect 7716 15202 7750 15236
rect 7716 15134 7750 15168
rect 7716 15066 7750 15100
rect 7716 14998 7750 15032
rect 7716 14930 7750 14964
rect 7716 14862 7750 14896
rect 7716 14794 7750 14828
rect 7716 14726 7750 14760
rect 7716 14658 7750 14692
rect 7716 14590 7750 14624
rect 7716 14522 7750 14556
rect 7716 14454 7750 14488
rect 7716 14386 7750 14420
rect 7716 14318 7750 14352
rect 7716 14250 7750 14284
rect 7716 7849 7750 7893
rect 7716 7781 7750 7815
rect 7716 7713 7750 7747
rect 7716 7645 7750 7679
rect 7716 7577 7750 7611
rect 7716 7509 7750 7543
rect 7716 7441 7750 7475
rect 7716 7373 7750 7407
rect 7716 7305 7750 7339
rect 7716 7237 7750 7271
rect 7716 7169 7750 7203
rect 7716 7101 7750 7135
rect 7716 7033 7750 7067
rect 7716 6965 7750 6999
rect 7716 6897 7750 6931
rect 7716 6829 7750 6863
rect 7716 6761 7750 6795
rect 7716 6693 7750 6727
rect 7716 6625 7750 6659
rect 7716 6557 7750 6591
rect 7716 6489 7750 6523
rect 7716 6421 7750 6455
rect 7716 6353 7750 6387
rect 7716 6285 7750 6319
rect 7716 6217 7750 6251
rect 7716 6149 7750 6183
rect 7716 6081 7750 6115
rect 7716 6013 7750 6047
rect 7716 5945 7750 5979
rect 7716 5877 7750 5911
rect 7716 5809 7750 5843
rect 7716 5741 7750 5775
rect 7716 5673 7750 5707
rect 7716 5605 7750 5639
rect 7716 5537 7750 5571
rect 7716 5469 7750 5503
rect 7716 5401 7750 5435
rect 7716 5333 7750 5367
rect 7716 5265 7750 5299
rect 7716 5197 7750 5231
rect 7716 5129 7750 5163
rect 7716 5061 7750 5095
rect 7716 4993 7750 5027
rect 7716 4925 7750 4959
rect 7716 4857 7750 4891
rect 7716 4789 7750 4823
rect 7716 4721 7750 4755
rect 7716 4653 7750 4687
rect 7716 4585 7750 4619
rect 7716 4517 7750 4551
rect 7716 4449 7750 4483
rect 7716 4381 7750 4415
rect 7716 4313 7750 4347
rect 7716 4245 7750 4279
rect 7716 4177 7750 4211
rect 7716 4109 7750 4143
rect 7716 4041 7750 4075
rect 7716 3973 7750 4007
rect 7716 3905 7750 3939
rect 7716 3837 7750 3871
rect 7716 3769 7750 3803
rect 7716 3701 7750 3735
rect 7716 3633 7750 3667
rect 7716 3565 7750 3599
rect 7716 3497 7750 3531
rect 7716 3429 7750 3463
rect 7716 3361 7750 3395
rect 7716 3293 7750 3327
rect 7716 3225 7750 3259
rect 7716 3157 7750 3191
rect 7716 3089 7750 3123
rect 7716 3021 7750 3055
rect 7716 2953 7750 2987
rect 7716 2885 7750 2919
rect 7716 2817 7750 2851
rect 7716 2749 7750 2783
rect 7716 2681 7750 2715
rect 7716 2613 7750 2647
rect 7716 2545 7750 2579
rect 7716 2477 7750 2511
<< mvpsubdiffcont >>
rect 2624 27873 2658 27907
rect 2693 27873 2727 27907
rect 2762 27873 2796 27907
rect 2831 27873 2865 27907
rect 2900 27873 2934 27907
rect 2969 27873 3003 27907
rect 2624 27805 2658 27839
rect 2693 27805 2727 27839
rect 2762 27805 2796 27839
rect 2831 27805 2865 27839
rect 2900 27805 2934 27839
rect 2969 27805 3003 27839
rect 2624 27737 2658 27771
rect 2693 27737 2727 27771
rect 2762 27737 2796 27771
rect 2831 27737 2865 27771
rect 2900 27737 2934 27771
rect 2969 27737 3003 27771
rect 2624 27669 2658 27703
rect 2693 27669 2727 27703
rect 2762 27669 2796 27703
rect 2831 27669 2865 27703
rect 2900 27669 2934 27703
rect 2969 27669 3003 27703
rect 2624 27601 2658 27635
rect 2693 27601 2727 27635
rect 2762 27601 2796 27635
rect 2831 27601 2865 27635
rect 2900 27601 2934 27635
rect 2969 27601 3003 27635
rect 2624 27533 2658 27567
rect 2693 27533 2727 27567
rect 2762 27533 2796 27567
rect 2831 27533 2865 27567
rect 2900 27533 2934 27567
rect 2969 27533 3003 27567
rect 2624 27465 2658 27499
rect 2693 27465 2727 27499
rect 2762 27465 2796 27499
rect 2831 27465 2865 27499
rect 2900 27465 2934 27499
rect 2969 27465 3003 27499
rect 3038 27465 7968 27907
rect 7083 27397 7185 27465
rect 7083 27257 7117 27291
rect 7151 27257 7185 27291
rect 7083 27117 7117 27151
rect 7151 27117 7185 27151
rect 7083 26977 7117 27011
rect 7151 26977 7185 27011
rect 7083 26837 7117 26871
rect 7151 26837 7185 26871
rect 7083 26697 7117 26731
rect 7151 26697 7185 26731
rect 7083 26557 7117 26591
rect 7151 26557 7185 26591
rect 7083 26417 7117 26451
rect 7151 26417 7185 26451
rect 7083 26277 7117 26311
rect 7151 26277 7185 26311
rect 7083 26137 7117 26171
rect 7151 26137 7185 26171
rect 7083 25997 7117 26031
rect 7151 25997 7185 26031
rect 7083 25857 7117 25891
rect 7151 25857 7185 25891
rect 7083 25717 7117 25751
rect 7151 25717 7185 25751
rect 7083 25577 7117 25611
rect 7151 25577 7185 25611
rect 7083 25437 7117 25471
rect 7151 25437 7185 25471
rect 7083 25296 7117 25330
rect 7151 25296 7185 25330
rect 7083 25155 7117 25189
rect 7151 25155 7185 25189
rect 7083 25014 7117 25048
rect 7151 25014 7185 25048
rect 7083 24873 7117 24907
rect 7151 24873 7185 24907
rect 7083 24732 7117 24766
rect 7151 24732 7185 24766
rect 7083 24591 7117 24625
rect 7151 24591 7185 24625
rect 3766 24483 3800 24517
rect 3836 24483 3870 24517
rect 3906 24483 3940 24517
rect 3976 24483 4010 24517
rect 4046 24483 4080 24517
rect 4116 24483 4150 24517
rect 4186 24483 4220 24517
rect 4256 24483 4290 24517
rect 4326 24483 4360 24517
rect 4396 24483 4430 24517
rect 4466 24483 4500 24517
rect 4536 24483 4570 24517
rect 4606 24483 4640 24517
rect 4675 24483 4709 24517
rect 4744 24483 4778 24517
rect 4813 24483 4847 24517
rect 4882 24483 4916 24517
rect 4951 24483 4985 24517
rect 5020 24483 5054 24517
rect 5089 24483 5123 24517
rect 5158 24483 5192 24517
rect 5227 24483 5261 24517
rect 5296 24483 5330 24517
rect 5365 24483 5399 24517
rect 5434 24483 5468 24517
rect 5503 24483 5537 24517
rect 5572 24483 5606 24517
rect 5641 24483 5675 24517
rect 5710 24483 5744 24517
rect 5779 24483 5813 24517
rect 5848 24483 5882 24517
rect 5917 24483 5951 24517
rect 5986 24483 6020 24517
rect 6055 24483 6089 24517
rect 6124 24483 6158 24517
rect 3766 24415 3800 24449
rect 3836 24415 3870 24449
rect 3906 24415 3940 24449
rect 3976 24415 4010 24449
rect 4046 24415 4080 24449
rect 4116 24415 4150 24449
rect 4186 24415 4220 24449
rect 4256 24415 4290 24449
rect 4326 24415 4360 24449
rect 4396 24415 4430 24449
rect 4466 24415 4500 24449
rect 4536 24415 4570 24449
rect 4606 24415 4640 24449
rect 4675 24415 4709 24449
rect 4744 24415 4778 24449
rect 4813 24415 4847 24449
rect 4882 24415 4916 24449
rect 4951 24415 4985 24449
rect 5020 24415 5054 24449
rect 5089 24415 5123 24449
rect 5158 24415 5192 24449
rect 5227 24415 5261 24449
rect 5296 24415 5330 24449
rect 5365 24415 5399 24449
rect 5434 24415 5468 24449
rect 5503 24415 5537 24449
rect 5572 24415 5606 24449
rect 5641 24415 5675 24449
rect 5710 24415 5744 24449
rect 5779 24415 5813 24449
rect 5848 24415 5882 24449
rect 5917 24415 5951 24449
rect 5986 24415 6020 24449
rect 6055 24415 6089 24449
rect 6124 24415 6158 24449
rect 3766 24347 3800 24381
rect 3836 24347 3870 24381
rect 3906 24347 3940 24381
rect 3976 24347 4010 24381
rect 4046 24347 4080 24381
rect 4116 24347 4150 24381
rect 4186 24347 4220 24381
rect 4256 24347 4290 24381
rect 4326 24347 4360 24381
rect 4396 24347 4430 24381
rect 4466 24347 4500 24381
rect 4536 24347 4570 24381
rect 4606 24347 4640 24381
rect 4675 24347 4709 24381
rect 4744 24347 4778 24381
rect 4813 24347 4847 24381
rect 4882 24347 4916 24381
rect 4951 24347 4985 24381
rect 5020 24347 5054 24381
rect 5089 24347 5123 24381
rect 5158 24347 5192 24381
rect 5227 24347 5261 24381
rect 5296 24347 5330 24381
rect 5365 24347 5399 24381
rect 5434 24347 5468 24381
rect 5503 24347 5537 24381
rect 5572 24347 5606 24381
rect 5641 24347 5675 24381
rect 5710 24347 5744 24381
rect 5779 24347 5813 24381
rect 5848 24347 5882 24381
rect 5917 24347 5951 24381
rect 5986 24347 6020 24381
rect 6055 24347 6089 24381
rect 6124 24347 6158 24381
rect 7083 24450 7117 24484
rect 7151 24450 7185 24484
rect 7083 24309 7117 24343
rect 7151 24309 7185 24343
rect 7083 24168 7117 24202
rect 7151 24168 7185 24202
rect 7083 24027 7117 24061
rect 7151 24027 7185 24061
rect 7083 23886 7117 23920
rect 7151 23886 7185 23920
rect 7083 23745 7117 23779
rect 7151 23745 7185 23779
rect 7083 23604 7117 23638
rect 7151 23604 7185 23638
rect 7083 23463 7117 23497
rect 7151 23463 7185 23497
rect 7083 23322 7117 23356
rect 7151 23322 7185 23356
rect 6089 23212 6123 23246
rect 6230 23212 6264 23246
rect 6372 23212 6406 23246
rect 6514 23212 6548 23246
rect 6656 23212 6690 23246
rect 6798 23212 6832 23246
rect 6940 23212 6974 23246
rect 7082 23212 7116 23246
rect 7224 23212 7258 23246
rect 7366 23212 7400 23246
rect 7508 23212 7542 23246
rect 7650 23212 7684 23246
rect 7792 23212 7826 23246
rect 7934 23212 7968 23246
rect 6089 23110 6123 23144
rect 6230 23110 6264 23144
rect 6372 23110 6406 23144
rect 6514 23110 6548 23144
rect 6656 23110 6690 23144
rect 6798 23110 6832 23144
rect 6940 23110 6974 23144
rect 7082 23110 7116 23144
rect 7224 23110 7258 23144
rect 7366 23110 7400 23144
rect 7508 23110 7542 23144
rect 7650 23110 7684 23144
rect 7792 23110 7826 23144
rect 7934 23110 7968 23144
rect 6089 23008 6123 23042
rect 6230 23008 6264 23042
rect 6372 23008 6406 23042
rect 6514 23008 6548 23042
rect 6656 23008 6690 23042
rect 6798 23008 6832 23042
rect 6940 23008 6974 23042
rect 7082 23008 7116 23042
rect 7224 23008 7258 23042
rect 7366 23008 7400 23042
rect 7508 23008 7542 23042
rect 7650 23008 7684 23042
rect 7792 23008 7826 23042
rect 7934 23008 7968 23042
rect 6089 22906 6123 22940
rect 6230 22906 6264 22940
rect 6372 22906 6406 22940
rect 6514 22906 6548 22940
rect 6656 22906 6690 22940
rect 6798 22906 6832 22940
rect 6940 22906 6974 22940
rect 7082 22906 7116 22940
rect 7224 22906 7258 22940
rect 7366 22906 7400 22940
rect 7508 22906 7542 22940
rect 7650 22906 7684 22940
rect 7792 22906 7826 22940
rect 7934 22906 7968 22940
rect 6089 22804 6123 22838
rect 6230 22804 6264 22838
rect 6372 22804 6406 22838
rect 6514 22804 6548 22838
rect 6656 22804 6690 22838
rect 6798 22804 6832 22838
rect 6940 22804 6974 22838
rect 7082 22804 7116 22838
rect 7224 22804 7258 22838
rect 7366 22804 7400 22838
rect 7508 22804 7542 22838
rect 7650 22804 7684 22838
rect 7792 22804 7826 22838
rect 7934 22804 7968 22838
rect 6089 22702 6123 22736
rect 6230 22702 6264 22736
rect 6372 22702 6406 22736
rect 6514 22702 6548 22736
rect 6656 22702 6690 22736
rect 6798 22702 6832 22736
rect 6940 22702 6974 22736
rect 7082 22702 7116 22736
rect 7224 22702 7258 22736
rect 7366 22702 7400 22736
rect 7508 22702 7542 22736
rect 7650 22702 7684 22736
rect 7792 22702 7826 22736
rect 7934 22702 7968 22736
rect 6089 22600 6123 22634
rect 6230 22600 6264 22634
rect 6372 22600 6406 22634
rect 6514 22600 6548 22634
rect 6656 22600 6690 22634
rect 6798 22600 6832 22634
rect 6940 22600 6974 22634
rect 7082 22600 7116 22634
rect 7224 22600 7258 22634
rect 7366 22600 7400 22634
rect 7508 22600 7542 22634
rect 7650 22600 7684 22634
rect 7792 22600 7826 22634
rect 7934 22600 7968 22634
rect 6089 22498 6123 22532
rect 6230 22498 6264 22532
rect 6372 22498 6406 22532
rect 6514 22498 6548 22532
rect 6656 22498 6690 22532
rect 6798 22498 6832 22532
rect 6940 22498 6974 22532
rect 7082 22498 7116 22532
rect 7224 22498 7258 22532
rect 7366 22498 7400 22532
rect 7508 22498 7542 22532
rect 7650 22498 7684 22532
rect 7792 22498 7826 22532
rect 7934 22498 7968 22532
rect 6364 14006 6398 14040
rect 6364 13937 6398 13971
rect 6364 13868 6398 13902
rect 6364 13799 6398 13833
rect 6364 13730 6398 13764
rect 6364 13661 6398 13695
rect 6364 13591 6398 13625
rect 6364 13521 6398 13555
rect 6364 13451 6398 13485
rect 7304 13868 7338 13902
rect 7304 13800 7338 13834
rect 7304 13732 7338 13766
rect 7304 13664 7338 13698
rect 7304 13596 7338 13630
rect 6364 13381 6398 13415
rect 6364 13311 6398 13345
rect 6364 13241 6398 13275
rect 6364 13171 6398 13205
rect 6364 13101 6398 13135
rect 6364 13031 6398 13065
rect 6364 12961 6398 12995
rect 6364 12891 6398 12925
rect 6364 12821 6398 12855
rect 7304 13528 7338 13562
rect 7304 13460 7338 13494
rect 7304 13392 7338 13426
rect 7304 13324 7338 13358
rect 7304 13255 7338 13289
rect 7304 13186 7338 13220
rect 7304 13117 7338 13151
rect 7304 13048 7338 13082
rect 7304 12979 7338 13013
rect 7304 12910 7338 12944
rect 7304 12841 7338 12875
rect 6364 12751 6398 12785
rect 6364 12681 6398 12715
rect 6364 12611 6398 12645
rect 7304 12772 7338 12806
rect 7304 12703 7338 12737
rect 6388 12456 6422 12490
rect 6458 12456 6492 12490
rect 6528 12456 6562 12490
rect 6598 12456 6632 12490
rect 6668 12456 6702 12490
rect 6738 12456 6772 12490
rect 6808 12456 6842 12490
rect 6878 12456 6912 12490
rect 6948 12456 6982 12490
rect 7018 12456 7052 12490
rect 7087 12456 7121 12490
rect 7156 12456 7190 12490
rect 7225 12456 7259 12490
rect 7294 12456 7328 12490
rect 7363 12456 7397 12490
rect 7432 12456 7466 12490
rect 7501 12456 7535 12490
rect 7570 12456 7604 12490
rect 6717 11003 6751 11037
rect 6717 10934 6751 10968
rect 6717 10865 6751 10899
rect 3139 10778 3173 10812
rect 3209 10778 3243 10812
rect 3279 10778 3313 10812
rect 3349 10778 3383 10812
rect 3419 10778 3453 10812
rect 3489 10778 3523 10812
rect 3559 10778 3593 10812
rect 3629 10778 3663 10812
rect 3699 10778 3733 10812
rect 3769 10778 3803 10812
rect 3839 10778 3873 10812
rect 3909 10778 3943 10812
rect 3979 10778 4013 10812
rect 4049 10778 4083 10812
rect 4119 10778 4153 10812
rect 4189 10778 4223 10812
rect 4258 10778 4292 10812
rect 4327 10778 4361 10812
rect 4396 10778 4430 10812
rect 4465 10778 4499 10812
rect 4534 10778 4568 10812
rect 6717 10796 6751 10830
rect 6717 10727 6751 10761
rect 5012 10680 5046 10714
rect 5081 10680 5115 10714
rect 5150 10680 5184 10714
rect 5219 10680 5253 10714
rect 5288 10680 5322 10714
rect 5357 10680 5391 10714
rect 5426 10680 5460 10714
rect 5495 10680 5529 10714
rect 5564 10680 5598 10714
rect 5633 10680 5667 10714
rect 5701 10680 5735 10714
rect 5769 10680 5803 10714
rect 5837 10680 5871 10714
rect 5905 10680 5939 10714
rect 5973 10680 6007 10714
rect 6041 10680 6075 10714
rect 6109 10680 6143 10714
rect 6177 10680 6211 10714
rect 6717 10658 6751 10692
rect 6717 10589 6751 10623
rect 6717 10520 6751 10554
rect 6717 10451 6751 10485
rect 6717 10382 6751 10416
rect 6717 10313 6751 10347
rect 6717 10244 6751 10278
rect 6717 10175 6751 10209
rect 6717 10106 6751 10140
rect 6717 10037 6751 10071
rect 6717 9968 6751 10002
rect 6717 9899 6751 9933
rect 6717 9830 6751 9864
rect 6717 9761 6751 9795
rect 6717 9692 6751 9726
rect 6717 9623 6751 9657
rect 6717 9554 6751 9588
rect 6717 9485 6751 9519
rect 6717 9416 6751 9450
rect 6717 9347 6751 9381
rect 6717 9278 6751 9312
rect 6717 9209 6751 9243
rect 6717 9141 6751 9175
rect 6717 9073 6751 9107
rect 6717 9005 6751 9039
rect 6717 8937 6751 8971
rect 6717 8869 6751 8903
rect 6717 8801 6751 8835
rect 6717 8733 6751 8767
rect 6717 8665 6751 8699
rect 6717 8597 6751 8631
rect 6717 8529 6751 8563
rect 6717 8461 6751 8495
rect 7071 2242 7105 2276
rect 7139 2242 7173 2276
rect 7207 2242 7241 2276
rect 7275 2242 7309 2276
rect 7343 2242 7377 2276
rect 7411 2242 7445 2276
rect 7479 2242 7513 2276
rect 7547 2242 7581 2276
rect 7615 2242 7649 2276
rect 7683 2242 7717 2276
rect 7751 2242 7785 2276
rect 7819 2242 7853 2276
rect 7887 2242 7921 2276
rect 7071 2173 7105 2207
rect 7139 2173 7173 2207
rect 7207 2173 7241 2207
rect 7275 2173 7309 2207
rect 7343 2173 7377 2207
rect 7411 2173 7445 2207
rect 7479 2173 7513 2207
rect 7547 2173 7581 2207
rect 7615 2173 7649 2207
rect 7683 2173 7717 2207
rect 7751 2173 7785 2207
rect 7819 2173 7853 2207
rect 7887 2173 7921 2207
rect 7071 2104 7105 2138
rect 7139 2104 7173 2138
rect 7207 2104 7241 2138
rect 7275 2104 7309 2138
rect 7343 2104 7377 2138
rect 7411 2104 7445 2138
rect 7479 2104 7513 2138
rect 7547 2104 7581 2138
rect 7615 2104 7649 2138
rect 7683 2104 7717 2138
rect 7751 2104 7785 2138
rect 7819 2104 7853 2138
rect 7887 2104 7921 2138
rect 7071 2034 7105 2068
rect 7139 2034 7173 2068
rect 7207 2034 7241 2068
rect 7275 2034 7309 2068
rect 7343 2034 7377 2068
rect 7411 2034 7445 2068
rect 7479 2034 7513 2068
rect 7547 2034 7581 2068
rect 7615 2034 7649 2068
rect 7683 2034 7717 2068
rect 7751 2034 7785 2068
rect 7819 2034 7853 2068
rect 7887 2034 7921 2068
rect 7071 1964 7105 1998
rect 7139 1964 7173 1998
rect 7207 1964 7241 1998
rect 7275 1964 7309 1998
rect 7343 1964 7377 1998
rect 7411 1964 7445 1998
rect 7479 1964 7513 1998
rect 7547 1964 7581 1998
rect 7615 1964 7649 1998
rect 7683 1964 7717 1998
rect 7751 1964 7785 1998
rect 7819 1964 7853 1998
rect 7887 1964 7921 1998
rect 7071 1894 7105 1928
rect 7139 1894 7173 1928
rect 7207 1894 7241 1928
rect 7275 1894 7309 1928
rect 7343 1894 7377 1928
rect 7411 1894 7445 1928
rect 7479 1894 7513 1928
rect 7547 1894 7581 1928
rect 7615 1894 7649 1928
rect 7683 1894 7717 1928
rect 7751 1894 7785 1928
rect 7819 1894 7853 1928
rect 7887 1894 7921 1928
rect 7071 1824 7105 1858
rect 7139 1824 7173 1858
rect 7207 1824 7241 1858
rect 7275 1824 7309 1858
rect 7343 1824 7377 1858
rect 7411 1824 7445 1858
rect 7479 1824 7513 1858
rect 7547 1824 7581 1858
rect 7615 1824 7649 1858
rect 7683 1824 7717 1858
rect 7751 1824 7785 1858
rect 7819 1824 7853 1858
rect 7887 1824 7921 1858
rect 7071 1754 7105 1788
rect 7139 1754 7173 1788
rect 7207 1754 7241 1788
rect 7275 1754 7309 1788
rect 7343 1754 7377 1788
rect 7411 1754 7445 1788
rect 7479 1754 7513 1788
rect 7547 1754 7581 1788
rect 7615 1754 7649 1788
rect 7683 1754 7717 1788
rect 7751 1754 7785 1788
rect 7819 1754 7853 1788
rect 7887 1754 7921 1788
rect 7071 1684 7105 1718
rect 7139 1684 7173 1718
rect 7207 1684 7241 1718
rect 7275 1684 7309 1718
rect 7343 1684 7377 1718
rect 7411 1684 7445 1718
rect 7479 1684 7513 1718
rect 7547 1684 7581 1718
rect 7615 1684 7649 1718
rect 7683 1684 7717 1718
rect 7751 1684 7785 1718
rect 7819 1684 7853 1718
rect 7887 1684 7921 1718
rect 7071 1614 7105 1648
rect 7139 1614 7173 1648
rect 7207 1614 7241 1648
rect 7275 1614 7309 1648
rect 7343 1614 7377 1648
rect 7411 1614 7445 1648
rect 7479 1614 7513 1648
rect 7547 1614 7581 1648
rect 7615 1614 7649 1648
rect 7683 1614 7717 1648
rect 7751 1614 7785 1648
rect 7819 1614 7853 1648
rect 7887 1614 7921 1648
rect 7071 1544 7105 1578
rect 7139 1544 7173 1578
rect 7207 1544 7241 1578
rect 7275 1544 7309 1578
rect 7343 1544 7377 1578
rect 7411 1544 7445 1578
rect 7479 1544 7513 1578
rect 7547 1544 7581 1578
rect 7615 1544 7649 1578
rect 7683 1544 7717 1578
rect 7751 1544 7785 1578
rect 7819 1544 7853 1578
rect 7887 1544 7921 1578
rect 7071 1474 7105 1508
rect 7139 1474 7173 1508
rect 7207 1474 7241 1508
rect 7275 1474 7309 1508
rect 7343 1474 7377 1508
rect 7411 1474 7445 1508
rect 7479 1474 7513 1508
rect 7547 1474 7581 1508
rect 7615 1474 7649 1508
rect 7683 1474 7717 1508
rect 7751 1474 7785 1508
rect 7819 1474 7853 1508
rect 7887 1474 7921 1508
rect 7071 1404 7105 1438
rect 7139 1404 7173 1438
rect 7207 1404 7241 1438
rect 7275 1404 7309 1438
rect 7343 1404 7377 1438
rect 7411 1404 7445 1438
rect 7479 1404 7513 1438
rect 7547 1404 7581 1438
rect 7615 1404 7649 1438
rect 7683 1404 7717 1438
rect 7751 1404 7785 1438
rect 7819 1404 7853 1438
rect 7887 1404 7921 1438
rect 7071 1334 7105 1368
rect 7139 1334 7173 1368
rect 7207 1334 7241 1368
rect 7275 1334 7309 1368
rect 7343 1334 7377 1368
rect 7411 1334 7445 1368
rect 7479 1334 7513 1368
rect 7547 1334 7581 1368
rect 7615 1334 7649 1368
rect 7683 1334 7717 1368
rect 7751 1334 7785 1368
rect 7819 1334 7853 1368
rect 7887 1334 7921 1368
rect 7071 1264 7105 1298
rect 7139 1264 7173 1298
rect 7207 1264 7241 1298
rect 7275 1264 7309 1298
rect 7343 1264 7377 1298
rect 7411 1264 7445 1298
rect 7479 1264 7513 1298
rect 7547 1264 7581 1298
rect 7615 1264 7649 1298
rect 7683 1264 7717 1298
rect 7751 1264 7785 1298
rect 7819 1264 7853 1298
rect 7887 1264 7921 1298
rect 7071 1194 7105 1228
rect 7139 1194 7173 1228
rect 7207 1194 7241 1228
rect 7275 1194 7309 1228
rect 7343 1194 7377 1228
rect 7411 1194 7445 1228
rect 7479 1194 7513 1228
rect 7547 1194 7581 1228
rect 7615 1194 7649 1228
rect 7683 1194 7717 1228
rect 7751 1194 7785 1228
rect 7819 1194 7853 1228
rect 7887 1194 7921 1228
rect 7071 1124 7105 1158
rect 7139 1124 7173 1158
rect 7207 1124 7241 1158
rect 7275 1124 7309 1158
rect 7343 1124 7377 1158
rect 7411 1124 7445 1158
rect 7479 1124 7513 1158
rect 7547 1124 7581 1158
rect 7615 1124 7649 1158
rect 7683 1124 7717 1158
rect 7751 1124 7785 1158
rect 7819 1124 7853 1158
rect 7887 1124 7921 1158
rect 7071 1054 7105 1088
rect 7139 1054 7173 1088
rect 7207 1054 7241 1088
rect 7275 1054 7309 1088
rect 7343 1054 7377 1088
rect 7411 1054 7445 1088
rect 7479 1054 7513 1088
rect 7547 1054 7581 1088
rect 7615 1054 7649 1088
rect 7683 1054 7717 1088
rect 7751 1054 7785 1088
rect 7819 1054 7853 1088
rect 7887 1054 7921 1088
rect 7071 984 7105 1018
rect 7139 984 7173 1018
rect 7207 984 7241 1018
rect 7275 984 7309 1018
rect 7343 984 7377 1018
rect 7411 984 7445 1018
rect 7479 984 7513 1018
rect 7547 984 7581 1018
rect 7615 984 7649 1018
rect 7683 984 7717 1018
rect 7751 984 7785 1018
rect 7819 984 7853 1018
rect 7887 984 7921 1018
rect 7071 914 7105 948
rect 7139 914 7173 948
rect 7207 914 7241 948
rect 7275 914 7309 948
rect 7343 914 7377 948
rect 7411 914 7445 948
rect 7479 914 7513 948
rect 7547 914 7581 948
rect 7615 914 7649 948
rect 7683 914 7717 948
rect 7751 914 7785 948
rect 7819 914 7853 948
rect 7887 914 7921 948
rect 7071 844 7105 878
rect 7139 844 7173 878
rect 7207 844 7241 878
rect 7275 844 7309 878
rect 7343 844 7377 878
rect 7411 844 7445 878
rect 7479 844 7513 878
rect 7547 844 7581 878
rect 7615 844 7649 878
rect 7683 844 7717 878
rect 7751 844 7785 878
rect 7819 844 7853 878
rect 7887 844 7921 878
rect 7071 774 7105 808
rect 7139 774 7173 808
rect 7207 774 7241 808
rect 7275 774 7309 808
rect 7343 774 7377 808
rect 7411 774 7445 808
rect 7479 774 7513 808
rect 7547 774 7581 808
rect 7615 774 7649 808
rect 7683 774 7717 808
rect 7751 774 7785 808
rect 7819 774 7853 808
rect 7887 774 7921 808
rect 7071 704 7105 738
rect 7139 704 7173 738
rect 7207 704 7241 738
rect 7275 704 7309 738
rect 7343 704 7377 738
rect 7411 704 7445 738
rect 7479 704 7513 738
rect 7547 704 7581 738
rect 7615 704 7649 738
rect 7683 704 7717 738
rect 7751 704 7785 738
rect 7819 704 7853 738
rect 7887 704 7921 738
rect 7071 634 7105 668
rect 7139 634 7173 668
rect 7207 634 7241 668
rect 7275 634 7309 668
rect 7343 634 7377 668
rect 7411 634 7445 668
rect 7479 634 7513 668
rect 7547 634 7581 668
rect 7615 634 7649 668
rect 7683 634 7717 668
rect 7751 634 7785 668
rect 7819 634 7853 668
rect 7887 634 7921 668
rect 7071 564 7105 598
rect 7139 564 7173 598
rect 7207 564 7241 598
rect 7275 564 7309 598
rect 7343 564 7377 598
rect 7411 564 7445 598
rect 7479 564 7513 598
rect 7547 564 7581 598
rect 7615 564 7649 598
rect 7683 564 7717 598
rect 7751 564 7785 598
rect 7819 564 7853 598
rect 7887 564 7921 598
rect 7071 494 7105 528
rect 7139 494 7173 528
rect 7207 494 7241 528
rect 7275 494 7309 528
rect 7343 494 7377 528
rect 7411 494 7445 528
rect 7479 494 7513 528
rect 7547 494 7581 528
rect 7615 494 7649 528
rect 7683 494 7717 528
rect 7751 494 7785 528
rect 7819 494 7853 528
rect 7887 494 7921 528
rect 7071 424 7105 458
rect 7139 424 7173 458
rect 7207 424 7241 458
rect 7275 424 7309 458
rect 7343 424 7377 458
rect 7411 424 7445 458
rect 7479 424 7513 458
rect 7547 424 7581 458
rect 7615 424 7649 458
rect 7683 424 7717 458
rect 7751 424 7785 458
rect 7819 424 7853 458
rect 7887 424 7921 458
rect 7071 354 7105 388
rect 7139 354 7173 388
rect 7207 354 7241 388
rect 7275 354 7309 388
rect 7343 354 7377 388
rect 7411 354 7445 388
rect 7479 354 7513 388
rect 7547 354 7581 388
rect 7615 354 7649 388
rect 7683 354 7717 388
rect 7751 354 7785 388
rect 7819 354 7853 388
rect 7887 354 7921 388
rect 7071 284 7105 318
rect 7139 284 7173 318
rect 7207 284 7241 318
rect 7275 284 7309 318
rect 7343 284 7377 318
rect 7411 284 7445 318
rect 7479 284 7513 318
rect 7547 284 7581 318
rect 7615 284 7649 318
rect 7683 284 7717 318
rect 7751 284 7785 318
rect 7819 284 7853 318
rect 7887 284 7921 318
rect 7071 214 7105 248
rect 7139 214 7173 248
rect 7207 214 7241 248
rect 7275 214 7309 248
rect 7343 214 7377 248
rect 7411 214 7445 248
rect 7479 214 7513 248
rect 7547 214 7581 248
rect 7615 214 7649 248
rect 7683 214 7717 248
rect 7751 214 7785 248
rect 7819 214 7853 248
rect 7887 214 7921 248
rect 7071 144 7105 178
rect 7139 144 7173 178
rect 7207 144 7241 178
rect 7275 144 7309 178
rect 7343 144 7377 178
rect 7411 144 7445 178
rect 7479 144 7513 178
rect 7547 144 7581 178
rect 7615 144 7649 178
rect 7683 144 7717 178
rect 7751 144 7785 178
rect 7819 144 7853 178
rect 7887 144 7921 178
rect 7071 74 7105 108
rect 7139 74 7173 108
rect 7207 74 7241 108
rect 7275 74 7309 108
rect 7343 74 7377 108
rect 7411 74 7445 108
rect 7479 74 7513 108
rect 7547 74 7581 108
rect 7615 74 7649 108
rect 7683 74 7717 108
rect 7751 74 7785 108
rect 7819 74 7853 108
rect 7887 74 7921 108
<< mvnsubdiffcont >>
rect 7716 19588 7750 19622
rect 7716 19520 7750 19554
rect 7716 19452 7750 19486
rect 7716 19384 7750 19418
rect 7716 19316 7750 19350
rect 7716 19248 7750 19282
rect 7716 19180 7750 19214
rect 7716 19112 7750 19146
rect 7716 19044 7750 19078
rect 7716 18976 7750 19010
rect 7716 18908 7750 18942
rect 7716 18840 7750 18874
rect 7716 18772 7750 18806
rect 7716 18704 7750 18738
rect 7716 18636 7750 18670
rect 7716 18568 7750 18602
rect 7716 18500 7750 18534
rect 7716 18432 7750 18466
rect 7716 18364 7750 18398
rect 7716 18296 7750 18330
rect 7716 18228 7750 18262
rect 7716 18160 7750 18194
rect 7716 18092 7750 18126
rect 7716 18024 7750 18058
rect 7716 17956 7750 17990
rect 7716 17888 7750 17922
rect 7716 17820 7750 17854
rect 7716 17752 7750 17786
rect 7716 17684 7750 17718
rect 7716 17616 7750 17650
rect 7716 17548 7750 17582
rect 7716 17480 7750 17514
rect 7716 17412 7750 17446
rect 7716 17344 7750 17378
rect 7716 17276 7750 17310
rect 7716 17208 7750 17242
rect 7716 17140 7750 17174
rect 7716 17072 7750 17106
rect 7716 17004 7750 17038
rect 7716 16936 7750 16970
rect 7716 16868 7750 16902
rect 7716 16800 7750 16834
rect 7716 16732 7750 16766
rect 7716 16664 7750 16698
rect 7716 16596 7750 16630
rect 7716 16528 7750 16562
rect 7716 16460 7750 16494
rect 7716 16392 7750 16426
rect 7716 16324 7750 16358
rect 7716 16256 7750 16290
rect 7716 16188 7750 16222
rect 7716 16120 7750 16154
rect 7716 16052 7750 16086
rect 7716 15984 7750 16018
rect 7716 15916 7750 15950
rect 7716 15848 7750 15882
rect 7716 15780 7750 15814
rect 7716 15712 7750 15746
rect 7716 15644 7750 15678
rect 7716 15576 7750 15610
rect 7716 15508 7750 15542
rect 7716 15440 7750 15474
rect 7716 15372 7750 15406
rect 7716 15304 7750 15338
rect 7716 15236 7750 15270
rect 7716 15168 7750 15202
rect 7716 15100 7750 15134
rect 7716 15032 7750 15066
rect 7716 14964 7750 14998
rect 7716 14896 7750 14930
rect 7716 14828 7750 14862
rect 7716 14760 7750 14794
rect 7716 14692 7750 14726
rect 7716 14624 7750 14658
rect 7716 14556 7750 14590
rect 7716 14488 7750 14522
rect 7716 14420 7750 14454
rect 7716 14352 7750 14386
rect 7716 14284 7750 14318
rect 7716 7815 7750 7849
rect 7716 7747 7750 7781
rect 7716 7679 7750 7713
rect 7716 7611 7750 7645
rect 7716 7543 7750 7577
rect 7716 7475 7750 7509
rect 7716 7407 7750 7441
rect 7716 7339 7750 7373
rect 7716 7271 7750 7305
rect 7716 7203 7750 7237
rect 7716 7135 7750 7169
rect 7716 7067 7750 7101
rect 7716 6999 7750 7033
rect 7716 6931 7750 6965
rect 7716 6863 7750 6897
rect 7716 6795 7750 6829
rect 7716 6727 7750 6761
rect 7716 6659 7750 6693
rect 7716 6591 7750 6625
rect 7716 6523 7750 6557
rect 7716 6455 7750 6489
rect 7716 6387 7750 6421
rect 7716 6319 7750 6353
rect 7716 6251 7750 6285
rect 7716 6183 7750 6217
rect 7716 6115 7750 6149
rect 7716 6047 7750 6081
rect 7716 5979 7750 6013
rect 7716 5911 7750 5945
rect 7716 5843 7750 5877
rect 7716 5775 7750 5809
rect 7716 5707 7750 5741
rect 7716 5639 7750 5673
rect 7716 5571 7750 5605
rect 7716 5503 7750 5537
rect 7716 5435 7750 5469
rect 7716 5367 7750 5401
rect 7716 5299 7750 5333
rect 7716 5231 7750 5265
rect 7716 5163 7750 5197
rect 7716 5095 7750 5129
rect 7716 5027 7750 5061
rect 7716 4959 7750 4993
rect 7716 4891 7750 4925
rect 7716 4823 7750 4857
rect 7716 4755 7750 4789
rect 7716 4687 7750 4721
rect 7716 4619 7750 4653
rect 7716 4551 7750 4585
rect 7716 4483 7750 4517
rect 7716 4415 7750 4449
rect 7716 4347 7750 4381
rect 7716 4279 7750 4313
rect 7716 4211 7750 4245
rect 7716 4143 7750 4177
rect 7716 4075 7750 4109
rect 7716 4007 7750 4041
rect 7716 3939 7750 3973
rect 7716 3871 7750 3905
rect 7716 3803 7750 3837
rect 7716 3735 7750 3769
rect 7716 3667 7750 3701
rect 7716 3599 7750 3633
rect 7716 3531 7750 3565
rect 7716 3463 7750 3497
rect 7716 3395 7750 3429
rect 7716 3327 7750 3361
rect 7716 3259 7750 3293
rect 7716 3191 7750 3225
rect 7716 3123 7750 3157
rect 7716 3055 7750 3089
rect 7716 2987 7750 3021
rect 7716 2919 7750 2953
rect 7716 2851 7750 2885
rect 7716 2783 7750 2817
rect 7716 2715 7750 2749
rect 7716 2647 7750 2681
rect 7716 2579 7750 2613
rect 7716 2511 7750 2545
<< poly >>
rect 3268 27296 3340 27330
rect 3268 27262 3284 27296
rect 3318 27262 3340 27296
rect 3268 27230 3340 27262
rect 5472 27296 5544 27330
rect 5472 27262 5494 27296
rect 5528 27262 5544 27296
rect 5472 27230 5544 27262
rect 6357 19869 6423 19885
rect 6357 19835 6373 19869
rect 6407 19835 6423 19869
rect 6357 19798 6423 19835
rect 6357 19764 6373 19798
rect 6407 19764 6423 19798
rect 6357 19727 6423 19764
rect 6357 19693 6373 19727
rect 6407 19693 6423 19727
rect 6357 19655 6423 19693
rect 6357 19621 6373 19655
rect 6407 19621 6423 19655
rect 6357 19583 6423 19621
rect 6357 19549 6373 19583
rect 6407 19549 6423 19583
rect 6357 19511 6423 19549
rect 6357 19477 6373 19511
rect 6407 19477 6423 19511
rect 6357 19439 6423 19477
rect 6357 19405 6373 19439
rect 6407 19405 6423 19439
rect 6357 19367 6423 19405
rect 6357 19333 6373 19367
rect 6407 19333 6423 19367
rect 7608 19598 7674 19614
rect 7608 19564 7624 19598
rect 7658 19564 7674 19598
rect 7608 19503 7674 19564
rect 7608 19469 7624 19503
rect 7658 19469 7674 19503
rect 7608 19408 7674 19469
rect 7608 19374 7624 19408
rect 7658 19374 7674 19408
rect 7608 19358 7674 19374
rect 6357 19317 6423 19333
rect 7608 19286 7674 19302
rect 6357 19245 6423 19261
rect 6357 19211 6373 19245
rect 6407 19211 6423 19245
rect 6357 19174 6423 19211
rect 6357 19140 6373 19174
rect 6407 19140 6423 19174
rect 6357 19103 6423 19140
rect 6357 19069 6373 19103
rect 6407 19069 6423 19103
rect 6357 19031 6423 19069
rect 6357 18997 6373 19031
rect 6407 18997 6423 19031
rect 6357 18959 6423 18997
rect 6357 18925 6373 18959
rect 6407 18925 6423 18959
rect 6357 18887 6423 18925
rect 6357 18853 6373 18887
rect 6407 18853 6423 18887
rect 6357 18815 6423 18853
rect 6357 18781 6373 18815
rect 6407 18781 6423 18815
rect 6357 18743 6423 18781
rect 6357 18709 6373 18743
rect 6407 18709 6423 18743
rect 6357 18693 6423 18709
rect 7608 19252 7624 19286
rect 7658 19252 7674 19286
rect 7608 19216 7674 19252
rect 7608 19182 7624 19216
rect 7658 19182 7674 19216
rect 7608 19146 7674 19182
rect 7608 19112 7624 19146
rect 7658 19112 7674 19146
rect 7608 19076 7674 19112
rect 7608 19042 7624 19076
rect 7658 19042 7674 19076
rect 7608 19006 7674 19042
rect 7608 18972 7624 19006
rect 7658 18972 7674 19006
rect 7608 18936 7674 18972
rect 7608 18902 7624 18936
rect 7658 18902 7674 18936
rect 7608 18866 7674 18902
rect 7608 18832 7624 18866
rect 7658 18832 7674 18866
rect 7608 18796 7674 18832
rect 7608 18762 7624 18796
rect 7658 18762 7674 18796
rect 7608 18726 7674 18762
rect 7608 18692 7624 18726
rect 7658 18692 7674 18726
rect 7608 18656 7674 18692
rect 6357 18621 6423 18637
rect 6357 18587 6373 18621
rect 6407 18587 6423 18621
rect 6357 18553 6423 18587
rect 6357 18519 6373 18553
rect 6407 18519 6423 18553
rect 6357 18503 6423 18519
rect 7608 18622 7624 18656
rect 7658 18622 7674 18656
rect 7608 18586 7674 18622
rect 7608 18552 7624 18586
rect 7658 18552 7674 18586
rect 7608 18515 7674 18552
rect 7608 18481 7624 18515
rect 7658 18481 7674 18515
rect 7608 18444 7674 18481
rect 7608 18410 7624 18444
rect 7658 18410 7674 18444
rect 7608 18373 7674 18410
rect 7608 18339 7624 18373
rect 7658 18339 7674 18373
rect 7608 18302 7674 18339
rect 7608 18268 7624 18302
rect 7658 18268 7674 18302
rect 7608 18231 7674 18268
rect 7608 18197 7624 18231
rect 7658 18197 7674 18231
rect 7608 18160 7674 18197
rect 7608 18126 7624 18160
rect 7658 18126 7674 18160
rect 7608 18110 7674 18126
rect 7608 18038 7674 18054
rect 7608 18004 7624 18038
rect 7658 18004 7674 18038
rect 7608 17969 7674 18004
rect 7608 17935 7624 17969
rect 7658 17935 7674 17969
rect 7608 17919 7674 17935
rect 7608 17772 7674 17788
rect 7608 17738 7624 17772
rect 7658 17738 7674 17772
rect 7608 17677 7674 17738
rect 7608 17643 7624 17677
rect 7658 17643 7674 17677
rect 7608 17582 7674 17643
rect 7608 17548 7624 17582
rect 7658 17548 7674 17582
rect 7608 17532 7674 17548
rect 7608 17460 7674 17476
rect 7608 17426 7624 17460
rect 7658 17426 7674 17460
rect 7608 17390 7674 17426
rect 7608 17356 7624 17390
rect 7658 17356 7674 17390
rect 7608 17320 7674 17356
rect 7608 17286 7624 17320
rect 7658 17286 7674 17320
rect 7608 17250 7674 17286
rect 7608 17216 7624 17250
rect 7658 17216 7674 17250
rect 7608 17180 7674 17216
rect 7608 17146 7624 17180
rect 7658 17146 7674 17180
rect 7608 17110 7674 17146
rect 7608 17076 7624 17110
rect 7658 17076 7674 17110
rect 7608 17040 7674 17076
rect 7608 17006 7624 17040
rect 7658 17006 7674 17040
rect 7608 16970 7674 17006
rect 7608 16936 7624 16970
rect 7658 16936 7674 16970
rect 7608 16900 7674 16936
rect 7608 16866 7624 16900
rect 7658 16866 7674 16900
rect 7608 16830 7674 16866
rect 7608 16796 7624 16830
rect 7658 16796 7674 16830
rect 7608 16760 7674 16796
rect 7608 16726 7624 16760
rect 7658 16726 7674 16760
rect 7608 16689 7674 16726
rect 7608 16655 7624 16689
rect 7658 16655 7674 16689
rect 7608 16618 7674 16655
rect 7608 16584 7624 16618
rect 7658 16584 7674 16618
rect 7608 16547 7674 16584
rect 7608 16513 7624 16547
rect 7658 16513 7674 16547
rect 7608 16476 7674 16513
rect 7608 16442 7624 16476
rect 7658 16442 7674 16476
rect 7608 16405 7674 16442
rect 7608 16371 7624 16405
rect 7658 16371 7674 16405
rect 7608 16334 7674 16371
rect 7608 16300 7624 16334
rect 7658 16300 7674 16334
rect 7608 16284 7674 16300
rect 7608 16212 7674 16228
rect 7608 16178 7624 16212
rect 7658 16178 7674 16212
rect 7608 16142 7674 16178
rect 7608 16108 7624 16142
rect 7658 16108 7674 16142
rect 7608 16092 7674 16108
rect 7608 15946 7674 15962
rect 7608 15912 7624 15946
rect 7658 15912 7674 15946
rect 7608 15851 7674 15912
rect 7608 15817 7624 15851
rect 7658 15817 7674 15851
rect 7608 15756 7674 15817
rect 7608 15722 7624 15756
rect 7658 15722 7674 15756
rect 7608 15706 7674 15722
rect 7608 15634 7674 15650
rect 7608 15600 7624 15634
rect 7658 15600 7674 15634
rect 7608 15564 7674 15600
rect 7608 15530 7624 15564
rect 7658 15530 7674 15564
rect 7608 15494 7674 15530
rect 7608 15460 7624 15494
rect 7658 15460 7674 15494
rect 7608 15424 7674 15460
rect 7608 15390 7624 15424
rect 7658 15390 7674 15424
rect 7608 15354 7674 15390
rect 7608 15320 7624 15354
rect 7658 15320 7674 15354
rect 7608 15284 7674 15320
rect 7608 15250 7624 15284
rect 7658 15250 7674 15284
rect 7608 15214 7674 15250
rect 7608 15180 7624 15214
rect 7658 15180 7674 15214
rect 7608 15144 7674 15180
rect 7608 15110 7624 15144
rect 7658 15110 7674 15144
rect 7608 15074 7674 15110
rect 7608 15040 7624 15074
rect 7658 15040 7674 15074
rect 7608 15004 7674 15040
rect 7608 14970 7624 15004
rect 7658 14970 7674 15004
rect 7608 14934 7674 14970
rect 7608 14900 7624 14934
rect 7658 14900 7674 14934
rect 7608 14863 7674 14900
rect 7608 14829 7624 14863
rect 7658 14829 7674 14863
rect 7608 14792 7674 14829
rect 7608 14758 7624 14792
rect 7658 14758 7674 14792
rect 7608 14721 7674 14758
rect 7608 14687 7624 14721
rect 7658 14687 7674 14721
rect 7608 14650 7674 14687
rect 7608 14616 7624 14650
rect 7658 14616 7674 14650
rect 7608 14579 7674 14616
rect 7608 14545 7624 14579
rect 7658 14545 7674 14579
rect 7608 14508 7674 14545
rect 7608 14474 7624 14508
rect 7658 14474 7674 14508
rect 7608 14458 7674 14474
rect 7608 14386 7674 14402
rect 7608 14352 7624 14386
rect 7658 14352 7674 14386
rect 7608 14317 7674 14352
rect 7608 14283 7624 14317
rect 7658 14283 7674 14317
rect 7608 14267 7674 14283
rect 6817 14015 6883 14031
rect 6654 13982 6720 13998
rect 6654 13948 6670 13982
rect 6704 13948 6720 13982
rect 6654 13911 6720 13948
rect 6654 13877 6670 13911
rect 6704 13877 6720 13911
rect 6654 13840 6720 13877
rect 6654 13806 6670 13840
rect 6704 13806 6720 13840
rect 6654 13768 6720 13806
rect 6654 13734 6670 13768
rect 6704 13734 6720 13768
rect 6654 13696 6720 13734
rect 6654 13662 6670 13696
rect 6704 13662 6720 13696
rect 6654 13624 6720 13662
rect 6654 13590 6670 13624
rect 6704 13590 6720 13624
rect 6817 13981 6833 14015
rect 6867 13981 6883 14015
rect 6817 13945 6883 13981
rect 6817 13911 6833 13945
rect 6867 13911 6883 13945
rect 7799 14015 7865 14031
rect 7799 13981 7815 14015
rect 7849 13981 7865 14015
rect 7799 13945 7865 13981
rect 6817 13876 6883 13911
rect 6817 13842 6833 13876
rect 6867 13842 6883 13876
rect 6817 13807 6883 13842
rect 6817 13773 6833 13807
rect 6867 13773 6883 13807
rect 6817 13738 6883 13773
rect 6817 13704 6833 13738
rect 6867 13704 6883 13738
rect 6817 13669 6883 13704
rect 6817 13635 6833 13669
rect 6867 13635 6883 13669
rect 6817 13619 6883 13635
rect 6654 13552 6720 13590
rect 7799 13911 7815 13945
rect 7849 13911 7865 13945
rect 7799 13876 7865 13911
rect 7799 13842 7815 13876
rect 7849 13842 7865 13876
rect 7799 13807 7865 13842
rect 7799 13773 7815 13807
rect 7849 13773 7865 13807
rect 7799 13738 7865 13773
rect 7799 13704 7815 13738
rect 7849 13704 7865 13738
rect 7799 13669 7865 13704
rect 7799 13635 7815 13669
rect 7849 13635 7865 13669
rect 7799 13619 7865 13635
rect 6654 13518 6670 13552
rect 6704 13518 6720 13552
rect 6654 13480 6720 13518
rect 6654 13446 6670 13480
rect 6704 13446 6720 13480
rect 6654 13430 6720 13446
rect 6817 13547 6883 13563
rect 6817 13513 6833 13547
rect 6867 13513 6883 13547
rect 6817 13475 6883 13513
rect 6817 13441 6833 13475
rect 6867 13441 6883 13475
rect 6817 13403 6883 13441
rect 6654 13358 6720 13374
rect 6654 13324 6670 13358
rect 6704 13324 6720 13358
rect 6654 13287 6720 13324
rect 6654 13253 6670 13287
rect 6704 13253 6720 13287
rect 6654 13216 6720 13253
rect 6654 13182 6670 13216
rect 6704 13182 6720 13216
rect 6654 13144 6720 13182
rect 6654 13110 6670 13144
rect 6704 13110 6720 13144
rect 6654 13072 6720 13110
rect 6654 13038 6670 13072
rect 6704 13038 6720 13072
rect 6654 13000 6720 13038
rect 6654 12966 6670 13000
rect 6704 12966 6720 13000
rect 6817 13369 6833 13403
rect 6867 13369 6883 13403
rect 6817 13331 6883 13369
rect 6817 13297 6833 13331
rect 6867 13297 6883 13331
rect 6817 13259 6883 13297
rect 6817 13225 6833 13259
rect 6867 13225 6883 13259
rect 6817 13187 6883 13225
rect 6817 13153 6833 13187
rect 6867 13153 6883 13187
rect 6817 13116 6883 13153
rect 6817 13082 6833 13116
rect 6867 13082 6883 13116
rect 6817 13045 6883 13082
rect 6817 13011 6833 13045
rect 6867 13011 6883 13045
rect 6817 12995 6883 13011
rect 6654 12928 6720 12966
rect 6654 12894 6670 12928
rect 6704 12894 6720 12928
rect 6654 12856 6720 12894
rect 6654 12822 6670 12856
rect 6704 12822 6720 12856
rect 7799 13547 7865 13563
rect 7799 13513 7815 13547
rect 7849 13513 7865 13547
rect 7799 13475 7865 13513
rect 7799 13441 7815 13475
rect 7849 13441 7865 13475
rect 7799 13403 7865 13441
rect 7799 13369 7815 13403
rect 7849 13369 7865 13403
rect 7799 13331 7865 13369
rect 7799 13297 7815 13331
rect 7849 13297 7865 13331
rect 7799 13259 7865 13297
rect 7799 13225 7815 13259
rect 7849 13225 7865 13259
rect 7799 13187 7865 13225
rect 7799 13153 7815 13187
rect 7849 13153 7865 13187
rect 7799 13116 7865 13153
rect 7799 13082 7815 13116
rect 7849 13082 7865 13116
rect 7799 13045 7865 13082
rect 7799 13011 7815 13045
rect 7849 13011 7865 13045
rect 7799 12995 7865 13011
rect 6654 12806 6720 12822
rect 6927 12813 6993 12829
rect 6927 12779 6943 12813
rect 6977 12779 6993 12813
rect 6654 12734 6720 12750
rect 6654 12700 6670 12734
rect 6704 12700 6720 12734
rect 6654 12666 6720 12700
rect 6927 12745 6993 12779
rect 6927 12711 6943 12745
rect 6977 12711 6993 12745
rect 6927 12695 6993 12711
rect 7649 12813 7715 12829
rect 7649 12779 7665 12813
rect 7699 12779 7715 12813
rect 7649 12745 7715 12779
rect 7649 12711 7665 12745
rect 7699 12711 7715 12745
rect 7649 12695 7715 12711
rect 6654 12632 6670 12666
rect 6704 12632 6720 12666
rect 6654 12616 6720 12632
rect 6397 12129 6531 12145
rect 6397 12095 6413 12129
rect 6447 12095 6481 12129
rect 6515 12095 6531 12129
rect 6397 12079 6531 12095
rect 6697 11979 7109 11995
rect 6697 11945 6713 11979
rect 6747 11945 6782 11979
rect 6816 11945 6851 11979
rect 6885 11945 6920 11979
rect 6954 11945 6989 11979
rect 7023 11945 7059 11979
rect 7093 11945 7109 11979
rect 6697 11929 7109 11945
rect 7165 11979 7733 11995
rect 7165 11945 7181 11979
rect 7215 11945 7252 11979
rect 7286 11945 7323 11979
rect 7357 11945 7395 11979
rect 7429 11945 7467 11979
rect 7501 11945 7539 11979
rect 7573 11945 7611 11979
rect 7645 11945 7683 11979
rect 7717 11945 7733 11979
rect 7165 11929 7733 11945
rect 5004 11172 5138 11188
rect 5004 11138 5020 11172
rect 5054 11138 5088 11172
rect 5122 11138 5138 11172
rect 3144 11118 3278 11134
rect 3144 11084 3160 11118
rect 3194 11084 3228 11118
rect 3262 11084 3278 11118
rect 3144 11068 3278 11084
rect 3334 11118 3902 11134
rect 3334 11084 3350 11118
rect 3384 11084 3422 11118
rect 3456 11084 3494 11118
rect 3528 11084 3566 11118
rect 3600 11084 3638 11118
rect 3672 11084 3710 11118
rect 3744 11084 3781 11118
rect 3815 11084 3852 11118
rect 3886 11084 3902 11118
rect 3334 11068 3902 11084
rect 3958 11118 4526 11134
rect 5004 11122 5138 11138
rect 5304 11172 5716 11188
rect 5304 11138 5320 11172
rect 5354 11138 5389 11172
rect 5423 11138 5458 11172
rect 5492 11138 5527 11172
rect 5561 11138 5596 11172
rect 5630 11138 5666 11172
rect 5700 11138 5716 11172
rect 5304 11122 5716 11138
rect 5772 11172 6340 11188
rect 5772 11138 5788 11172
rect 5822 11138 5859 11172
rect 5893 11138 5930 11172
rect 5964 11138 6002 11172
rect 6036 11138 6074 11172
rect 6108 11138 6146 11172
rect 6180 11138 6218 11172
rect 6252 11138 6290 11172
rect 6324 11138 6340 11172
rect 5772 11122 6340 11138
rect 3958 11084 3974 11118
rect 4008 11084 4046 11118
rect 4080 11084 4118 11118
rect 4152 11084 4190 11118
rect 4224 11084 4262 11118
rect 4296 11084 4334 11118
rect 4368 11084 4405 11118
rect 4439 11084 4476 11118
rect 4510 11084 4526 11118
rect 3958 11068 4526 11084
rect 7062 11055 7128 11071
rect 7062 11021 7078 11055
rect 7112 11021 7128 11055
rect 7062 10987 7128 11021
rect 7062 10953 7078 10987
rect 7112 10953 7128 10987
rect 7062 10937 7128 10953
rect 7212 10755 7278 10771
rect 7212 10721 7228 10755
rect 7262 10721 7278 10755
rect 7212 10686 7278 10721
rect 7212 10652 7228 10686
rect 7262 10652 7278 10686
rect 7212 10617 7278 10652
rect 7212 10583 7228 10617
rect 7262 10583 7278 10617
rect 7212 10548 7278 10583
rect 7212 10514 7228 10548
rect 7262 10514 7278 10548
rect 7212 10479 7278 10514
rect 7212 10445 7228 10479
rect 7262 10445 7278 10479
rect 7212 10409 7278 10445
rect 7212 10375 7228 10409
rect 7262 10375 7278 10409
rect 7212 10359 7278 10375
rect 7212 10287 7278 10303
rect 7212 10253 7228 10287
rect 7262 10253 7278 10287
rect 7212 10216 7278 10253
rect 7212 10182 7228 10216
rect 7262 10182 7278 10216
rect 7212 10145 7278 10182
rect 7212 10111 7228 10145
rect 7262 10111 7278 10145
rect 7212 10073 7278 10111
rect 7212 10039 7228 10073
rect 7262 10039 7278 10073
rect 7212 10001 7278 10039
rect 7212 9967 7228 10001
rect 7262 9967 7278 10001
rect 7212 9929 7278 9967
rect 7212 9895 7228 9929
rect 7262 9895 7278 9929
rect 7212 9857 7278 9895
rect 7212 9823 7228 9857
rect 7262 9823 7278 9857
rect 7212 9785 7278 9823
rect 7212 9751 7228 9785
rect 7262 9751 7278 9785
rect 7212 9735 7278 9751
rect 7212 9663 7278 9679
rect 7212 9629 7228 9663
rect 7262 9629 7278 9663
rect 7212 9592 7278 9629
rect 7212 9558 7228 9592
rect 7262 9558 7278 9592
rect 7212 9521 7278 9558
rect 7212 9487 7228 9521
rect 7262 9487 7278 9521
rect 7212 9449 7278 9487
rect 7212 9415 7228 9449
rect 7262 9415 7278 9449
rect 7212 9377 7278 9415
rect 7212 9343 7228 9377
rect 7262 9343 7278 9377
rect 7212 9305 7278 9343
rect 7212 9271 7228 9305
rect 7262 9271 7278 9305
rect 7212 9233 7278 9271
rect 7212 9199 7228 9233
rect 7262 9199 7278 9233
rect 7212 9161 7278 9199
rect 7212 9127 7228 9161
rect 7262 9127 7278 9161
rect 7212 9111 7278 9127
rect 7212 9039 7278 9055
rect 7212 9005 7228 9039
rect 7262 9005 7278 9039
rect 7212 8970 7278 9005
rect 7212 8936 7228 8970
rect 7262 8936 7278 8970
rect 7212 8901 7278 8936
rect 7212 8867 7228 8901
rect 7262 8867 7278 8901
rect 7212 8832 7278 8867
rect 7212 8798 7228 8832
rect 7262 8798 7278 8832
rect 7212 8763 7278 8798
rect 7212 8729 7228 8763
rect 7262 8729 7278 8763
rect 7212 8694 7278 8729
rect 7212 8660 7228 8694
rect 7262 8660 7278 8694
rect 7212 8644 7278 8660
rect 7062 8461 7128 8477
rect 7062 8427 7078 8461
rect 7112 8427 7128 8461
rect 7062 8393 7128 8427
rect 7062 8359 7078 8393
rect 7112 8359 7128 8393
rect 7062 8343 7128 8359
rect 7608 7825 7674 7841
rect 7608 7791 7624 7825
rect 7658 7791 7674 7825
rect 7608 7730 7674 7791
rect 7608 7696 7624 7730
rect 7658 7696 7674 7730
rect 7608 7635 7674 7696
rect 7608 7601 7624 7635
rect 7658 7601 7674 7635
rect 7608 7585 7674 7601
rect 7608 7513 7674 7529
rect 7608 7479 7624 7513
rect 7658 7479 7674 7513
rect 7608 7443 7674 7479
rect 7608 7409 7624 7443
rect 7658 7409 7674 7443
rect 7608 7373 7674 7409
rect 7608 7339 7624 7373
rect 7658 7339 7674 7373
rect 7608 7303 7674 7339
rect 7608 7269 7624 7303
rect 7658 7269 7674 7303
rect 7608 7233 7674 7269
rect 7608 7199 7624 7233
rect 7658 7199 7674 7233
rect 7608 7163 7674 7199
rect 7608 7129 7624 7163
rect 7658 7129 7674 7163
rect 7608 7093 7674 7129
rect 7608 7059 7624 7093
rect 7658 7059 7674 7093
rect 7608 7023 7674 7059
rect 7608 6989 7624 7023
rect 7658 6989 7674 7023
rect 7608 6953 7674 6989
rect 7608 6919 7624 6953
rect 7658 6919 7674 6953
rect 7608 6883 7674 6919
rect 7608 6849 7624 6883
rect 7658 6849 7674 6883
rect 7608 6813 7674 6849
rect 7608 6779 7624 6813
rect 7658 6779 7674 6813
rect 7608 6742 7674 6779
rect 7608 6708 7624 6742
rect 7658 6708 7674 6742
rect 7608 6671 7674 6708
rect 7608 6637 7624 6671
rect 7658 6637 7674 6671
rect 7608 6600 7674 6637
rect 7608 6566 7624 6600
rect 7658 6566 7674 6600
rect 7608 6529 7674 6566
rect 7608 6495 7624 6529
rect 7658 6495 7674 6529
rect 7608 6458 7674 6495
rect 7608 6424 7624 6458
rect 7658 6424 7674 6458
rect 7608 6387 7674 6424
rect 7608 6353 7624 6387
rect 7658 6353 7674 6387
rect 7608 6337 7674 6353
rect 7608 6265 7674 6281
rect 7608 6231 7624 6265
rect 7658 6231 7674 6265
rect 7608 6196 7674 6231
rect 7608 6162 7624 6196
rect 7658 6162 7674 6196
rect 7608 6146 7674 6162
rect 7608 5999 7674 6015
rect 7608 5965 7624 5999
rect 7658 5965 7674 5999
rect 7608 5904 7674 5965
rect 7608 5870 7624 5904
rect 7658 5870 7674 5904
rect 7608 5809 7674 5870
rect 7608 5775 7624 5809
rect 7658 5775 7674 5809
rect 7608 5759 7674 5775
rect 7608 5687 7674 5703
rect 7608 5653 7624 5687
rect 7658 5653 7674 5687
rect 7608 5617 7674 5653
rect 7608 5583 7624 5617
rect 7658 5583 7674 5617
rect 7608 5547 7674 5583
rect 7608 5513 7624 5547
rect 7658 5513 7674 5547
rect 7608 5477 7674 5513
rect 7608 5443 7624 5477
rect 7658 5443 7674 5477
rect 7608 5407 7674 5443
rect 7608 5373 7624 5407
rect 7658 5373 7674 5407
rect 7608 5337 7674 5373
rect 7608 5303 7624 5337
rect 7658 5303 7674 5337
rect 7608 5267 7674 5303
rect 7608 5233 7624 5267
rect 7658 5233 7674 5267
rect 7608 5197 7674 5233
rect 7608 5163 7624 5197
rect 7658 5163 7674 5197
rect 7608 5127 7674 5163
rect 7608 5093 7624 5127
rect 7658 5093 7674 5127
rect 7608 5057 7674 5093
rect 7608 5023 7624 5057
rect 7658 5023 7674 5057
rect 7608 4987 7674 5023
rect 7608 4953 7624 4987
rect 7658 4953 7674 4987
rect 7608 4916 7674 4953
rect 7608 4882 7624 4916
rect 7658 4882 7674 4916
rect 7608 4845 7674 4882
rect 7608 4811 7624 4845
rect 7658 4811 7674 4845
rect 7608 4774 7674 4811
rect 7608 4740 7624 4774
rect 7658 4740 7674 4774
rect 7608 4703 7674 4740
rect 7608 4669 7624 4703
rect 7658 4669 7674 4703
rect 7608 4632 7674 4669
rect 7608 4598 7624 4632
rect 7658 4598 7674 4632
rect 7608 4561 7674 4598
rect 7608 4527 7624 4561
rect 7658 4527 7674 4561
rect 7608 4511 7674 4527
rect 7608 4439 7674 4455
rect 7608 4405 7624 4439
rect 7658 4405 7674 4439
rect 7608 4370 7674 4405
rect 7608 4336 7624 4370
rect 7658 4336 7674 4370
rect 7608 4320 7674 4336
rect 7608 4173 7674 4189
rect 7608 4139 7624 4173
rect 7658 4139 7674 4173
rect 7608 4078 7674 4139
rect 7608 4044 7624 4078
rect 7658 4044 7674 4078
rect 7608 3983 7674 4044
rect 7608 3949 7624 3983
rect 7658 3949 7674 3983
rect 7608 3933 7674 3949
rect 7608 3861 7674 3877
rect 7608 3827 7624 3861
rect 7658 3827 7674 3861
rect 7608 3791 7674 3827
rect 7608 3757 7624 3791
rect 7658 3757 7674 3791
rect 7608 3721 7674 3757
rect 7608 3687 7624 3721
rect 7658 3687 7674 3721
rect 7608 3651 7674 3687
rect 7608 3617 7624 3651
rect 7658 3617 7674 3651
rect 4363 3591 4497 3607
rect 4363 3557 4379 3591
rect 4413 3557 4447 3591
rect 4481 3557 4497 3591
rect 4363 3541 4497 3557
rect 4553 3591 5121 3607
rect 4553 3557 4569 3591
rect 4603 3557 4641 3591
rect 4675 3557 4713 3591
rect 4747 3557 4785 3591
rect 4819 3557 4857 3591
rect 4891 3557 4929 3591
rect 4963 3557 5000 3591
rect 5034 3557 5071 3591
rect 5105 3557 5121 3591
rect 4553 3541 5121 3557
rect 5177 3591 5745 3607
rect 5177 3557 5193 3591
rect 5227 3557 5265 3591
rect 5299 3557 5337 3591
rect 5371 3557 5409 3591
rect 5443 3557 5481 3591
rect 5515 3557 5553 3591
rect 5587 3557 5624 3591
rect 5658 3557 5695 3591
rect 5729 3557 5745 3591
rect 5177 3541 5745 3557
rect 7608 3581 7674 3617
rect 7608 3547 7624 3581
rect 7658 3547 7674 3581
rect 7608 3511 7674 3547
rect 7608 3477 7624 3511
rect 7658 3477 7674 3511
rect 7608 3441 7674 3477
rect 7608 3407 7624 3441
rect 7658 3407 7674 3441
rect 7608 3371 7674 3407
rect 7608 3337 7624 3371
rect 7658 3337 7674 3371
rect 7608 3301 7674 3337
rect 7608 3267 7624 3301
rect 7658 3267 7674 3301
rect 7608 3231 7674 3267
rect 7608 3197 7624 3231
rect 7658 3197 7674 3231
rect 7608 3161 7674 3197
rect 7608 3127 7624 3161
rect 7658 3127 7674 3161
rect 7608 3090 7674 3127
rect 7608 3056 7624 3090
rect 7658 3056 7674 3090
rect 7608 3019 7674 3056
rect 7608 2985 7624 3019
rect 7658 2985 7674 3019
rect 7608 2948 7674 2985
rect 7608 2914 7624 2948
rect 7658 2914 7674 2948
rect 7608 2877 7674 2914
rect 7608 2843 7624 2877
rect 7658 2843 7674 2877
rect 7608 2806 7674 2843
rect 7608 2772 7624 2806
rect 7658 2772 7674 2806
rect 7608 2735 7674 2772
rect 7608 2701 7624 2735
rect 7658 2701 7674 2735
rect 7608 2685 7674 2701
rect 7608 2613 7674 2629
rect 7608 2579 7624 2613
rect 7658 2579 7674 2613
rect 7608 2545 7674 2579
rect 7608 2511 7624 2545
rect 7658 2511 7674 2545
rect 7608 2495 7674 2511
<< polycont >>
rect 3284 27262 3318 27296
rect 5494 27262 5528 27296
rect 6373 19835 6407 19869
rect 6373 19764 6407 19798
rect 6373 19693 6407 19727
rect 6373 19621 6407 19655
rect 6373 19549 6407 19583
rect 6373 19477 6407 19511
rect 6373 19405 6407 19439
rect 6373 19333 6407 19367
rect 7624 19564 7658 19598
rect 7624 19469 7658 19503
rect 7624 19374 7658 19408
rect 6373 19211 6407 19245
rect 6373 19140 6407 19174
rect 6373 19069 6407 19103
rect 6373 18997 6407 19031
rect 6373 18925 6407 18959
rect 6373 18853 6407 18887
rect 6373 18781 6407 18815
rect 6373 18709 6407 18743
rect 7624 19252 7658 19286
rect 7624 19182 7658 19216
rect 7624 19112 7658 19146
rect 7624 19042 7658 19076
rect 7624 18972 7658 19006
rect 7624 18902 7658 18936
rect 7624 18832 7658 18866
rect 7624 18762 7658 18796
rect 7624 18692 7658 18726
rect 6373 18587 6407 18621
rect 6373 18519 6407 18553
rect 7624 18622 7658 18656
rect 7624 18552 7658 18586
rect 7624 18481 7658 18515
rect 7624 18410 7658 18444
rect 7624 18339 7658 18373
rect 7624 18268 7658 18302
rect 7624 18197 7658 18231
rect 7624 18126 7658 18160
rect 7624 18004 7658 18038
rect 7624 17935 7658 17969
rect 7624 17738 7658 17772
rect 7624 17643 7658 17677
rect 7624 17548 7658 17582
rect 7624 17426 7658 17460
rect 7624 17356 7658 17390
rect 7624 17286 7658 17320
rect 7624 17216 7658 17250
rect 7624 17146 7658 17180
rect 7624 17076 7658 17110
rect 7624 17006 7658 17040
rect 7624 16936 7658 16970
rect 7624 16866 7658 16900
rect 7624 16796 7658 16830
rect 7624 16726 7658 16760
rect 7624 16655 7658 16689
rect 7624 16584 7658 16618
rect 7624 16513 7658 16547
rect 7624 16442 7658 16476
rect 7624 16371 7658 16405
rect 7624 16300 7658 16334
rect 7624 16178 7658 16212
rect 7624 16108 7658 16142
rect 7624 15912 7658 15946
rect 7624 15817 7658 15851
rect 7624 15722 7658 15756
rect 7624 15600 7658 15634
rect 7624 15530 7658 15564
rect 7624 15460 7658 15494
rect 7624 15390 7658 15424
rect 7624 15320 7658 15354
rect 7624 15250 7658 15284
rect 7624 15180 7658 15214
rect 7624 15110 7658 15144
rect 7624 15040 7658 15074
rect 7624 14970 7658 15004
rect 7624 14900 7658 14934
rect 7624 14829 7658 14863
rect 7624 14758 7658 14792
rect 7624 14687 7658 14721
rect 7624 14616 7658 14650
rect 7624 14545 7658 14579
rect 7624 14474 7658 14508
rect 7624 14352 7658 14386
rect 7624 14283 7658 14317
rect 6670 13948 6704 13982
rect 6670 13877 6704 13911
rect 6670 13806 6704 13840
rect 6670 13734 6704 13768
rect 6670 13662 6704 13696
rect 6670 13590 6704 13624
rect 6833 13981 6867 14015
rect 6833 13911 6867 13945
rect 7815 13981 7849 14015
rect 6833 13842 6867 13876
rect 6833 13773 6867 13807
rect 6833 13704 6867 13738
rect 6833 13635 6867 13669
rect 7815 13911 7849 13945
rect 7815 13842 7849 13876
rect 7815 13773 7849 13807
rect 7815 13704 7849 13738
rect 7815 13635 7849 13669
rect 6670 13518 6704 13552
rect 6670 13446 6704 13480
rect 6833 13513 6867 13547
rect 6833 13441 6867 13475
rect 6670 13324 6704 13358
rect 6670 13253 6704 13287
rect 6670 13182 6704 13216
rect 6670 13110 6704 13144
rect 6670 13038 6704 13072
rect 6670 12966 6704 13000
rect 6833 13369 6867 13403
rect 6833 13297 6867 13331
rect 6833 13225 6867 13259
rect 6833 13153 6867 13187
rect 6833 13082 6867 13116
rect 6833 13011 6867 13045
rect 6670 12894 6704 12928
rect 6670 12822 6704 12856
rect 7815 13513 7849 13547
rect 7815 13441 7849 13475
rect 7815 13369 7849 13403
rect 7815 13297 7849 13331
rect 7815 13225 7849 13259
rect 7815 13153 7849 13187
rect 7815 13082 7849 13116
rect 7815 13011 7849 13045
rect 6943 12779 6977 12813
rect 6670 12700 6704 12734
rect 6943 12711 6977 12745
rect 7665 12779 7699 12813
rect 7665 12711 7699 12745
rect 6670 12632 6704 12666
rect 6413 12095 6447 12129
rect 6481 12095 6515 12129
rect 6713 11945 6747 11979
rect 6782 11945 6816 11979
rect 6851 11945 6885 11979
rect 6920 11945 6954 11979
rect 6989 11945 7023 11979
rect 7059 11945 7093 11979
rect 7181 11945 7215 11979
rect 7252 11945 7286 11979
rect 7323 11945 7357 11979
rect 7395 11945 7429 11979
rect 7467 11945 7501 11979
rect 7539 11945 7573 11979
rect 7611 11945 7645 11979
rect 7683 11945 7717 11979
rect 5020 11138 5054 11172
rect 5088 11138 5122 11172
rect 3160 11084 3194 11118
rect 3228 11084 3262 11118
rect 3350 11084 3384 11118
rect 3422 11084 3456 11118
rect 3494 11084 3528 11118
rect 3566 11084 3600 11118
rect 3638 11084 3672 11118
rect 3710 11084 3744 11118
rect 3781 11084 3815 11118
rect 3852 11084 3886 11118
rect 5320 11138 5354 11172
rect 5389 11138 5423 11172
rect 5458 11138 5492 11172
rect 5527 11138 5561 11172
rect 5596 11138 5630 11172
rect 5666 11138 5700 11172
rect 5788 11138 5822 11172
rect 5859 11138 5893 11172
rect 5930 11138 5964 11172
rect 6002 11138 6036 11172
rect 6074 11138 6108 11172
rect 6146 11138 6180 11172
rect 6218 11138 6252 11172
rect 6290 11138 6324 11172
rect 3974 11084 4008 11118
rect 4046 11084 4080 11118
rect 4118 11084 4152 11118
rect 4190 11084 4224 11118
rect 4262 11084 4296 11118
rect 4334 11084 4368 11118
rect 4405 11084 4439 11118
rect 4476 11084 4510 11118
rect 7078 11021 7112 11055
rect 7078 10953 7112 10987
rect 7228 10721 7262 10755
rect 7228 10652 7262 10686
rect 7228 10583 7262 10617
rect 7228 10514 7262 10548
rect 7228 10445 7262 10479
rect 7228 10375 7262 10409
rect 7228 10253 7262 10287
rect 7228 10182 7262 10216
rect 7228 10111 7262 10145
rect 7228 10039 7262 10073
rect 7228 9967 7262 10001
rect 7228 9895 7262 9929
rect 7228 9823 7262 9857
rect 7228 9751 7262 9785
rect 7228 9629 7262 9663
rect 7228 9558 7262 9592
rect 7228 9487 7262 9521
rect 7228 9415 7262 9449
rect 7228 9343 7262 9377
rect 7228 9271 7262 9305
rect 7228 9199 7262 9233
rect 7228 9127 7262 9161
rect 7228 9005 7262 9039
rect 7228 8936 7262 8970
rect 7228 8867 7262 8901
rect 7228 8798 7262 8832
rect 7228 8729 7262 8763
rect 7228 8660 7262 8694
rect 7078 8427 7112 8461
rect 7078 8359 7112 8393
rect 7624 7791 7658 7825
rect 7624 7696 7658 7730
rect 7624 7601 7658 7635
rect 7624 7479 7658 7513
rect 7624 7409 7658 7443
rect 7624 7339 7658 7373
rect 7624 7269 7658 7303
rect 7624 7199 7658 7233
rect 7624 7129 7658 7163
rect 7624 7059 7658 7093
rect 7624 6989 7658 7023
rect 7624 6919 7658 6953
rect 7624 6849 7658 6883
rect 7624 6779 7658 6813
rect 7624 6708 7658 6742
rect 7624 6637 7658 6671
rect 7624 6566 7658 6600
rect 7624 6495 7658 6529
rect 7624 6424 7658 6458
rect 7624 6353 7658 6387
rect 7624 6231 7658 6265
rect 7624 6162 7658 6196
rect 7624 5965 7658 5999
rect 7624 5870 7658 5904
rect 7624 5775 7658 5809
rect 7624 5653 7658 5687
rect 7624 5583 7658 5617
rect 7624 5513 7658 5547
rect 7624 5443 7658 5477
rect 7624 5373 7658 5407
rect 7624 5303 7658 5337
rect 7624 5233 7658 5267
rect 7624 5163 7658 5197
rect 7624 5093 7658 5127
rect 7624 5023 7658 5057
rect 7624 4953 7658 4987
rect 7624 4882 7658 4916
rect 7624 4811 7658 4845
rect 7624 4740 7658 4774
rect 7624 4669 7658 4703
rect 7624 4598 7658 4632
rect 7624 4527 7658 4561
rect 7624 4405 7658 4439
rect 7624 4336 7658 4370
rect 7624 4139 7658 4173
rect 7624 4044 7658 4078
rect 7624 3949 7658 3983
rect 7624 3827 7658 3861
rect 7624 3757 7658 3791
rect 7624 3687 7658 3721
rect 7624 3617 7658 3651
rect 4379 3557 4413 3591
rect 4447 3557 4481 3591
rect 4569 3557 4603 3591
rect 4641 3557 4675 3591
rect 4713 3557 4747 3591
rect 4785 3557 4819 3591
rect 4857 3557 4891 3591
rect 4929 3557 4963 3591
rect 5000 3557 5034 3591
rect 5071 3557 5105 3591
rect 5193 3557 5227 3591
rect 5265 3557 5299 3591
rect 5337 3557 5371 3591
rect 5409 3557 5443 3591
rect 5481 3557 5515 3591
rect 5553 3557 5587 3591
rect 5624 3557 5658 3591
rect 5695 3557 5729 3591
rect 7624 3547 7658 3581
rect 7624 3477 7658 3511
rect 7624 3407 7658 3441
rect 7624 3337 7658 3371
rect 7624 3267 7658 3301
rect 7624 3197 7658 3231
rect 7624 3127 7658 3161
rect 7624 3056 7658 3090
rect 7624 2985 7658 3019
rect 7624 2914 7658 2948
rect 7624 2843 7658 2877
rect 7624 2772 7658 2806
rect 7624 2701 7658 2735
rect 7624 2579 7658 2613
rect 7624 2511 7658 2545
<< locali >>
rect 2590 27873 2624 27907
rect 2658 27873 2693 27907
rect 2727 27873 2762 27907
rect 2796 27873 2831 27907
rect 2865 27903 2900 27907
rect 2934 27903 2969 27907
rect 3003 27903 3038 27907
rect 2865 27873 2884 27903
rect 2934 27873 2957 27903
rect 3003 27873 3030 27903
rect 2590 27869 2884 27873
rect 2918 27869 2957 27873
rect 2991 27869 3030 27873
rect 2590 27839 3038 27869
rect 2590 27805 2624 27839
rect 2658 27805 2693 27839
rect 2727 27805 2762 27839
rect 2796 27805 2831 27839
rect 2865 27823 2900 27839
rect 2934 27823 2969 27839
rect 3003 27823 3038 27839
rect 2865 27805 2884 27823
rect 2934 27805 2957 27823
rect 3003 27805 3030 27823
rect 2590 27789 2884 27805
rect 2918 27789 2957 27805
rect 2991 27789 3030 27805
rect 2590 27771 3038 27789
rect 2590 27737 2624 27771
rect 2658 27737 2693 27771
rect 2727 27737 2762 27771
rect 2796 27737 2831 27771
rect 2865 27743 2900 27771
rect 2934 27743 2969 27771
rect 3003 27743 3038 27771
rect 2865 27737 2884 27743
rect 2934 27737 2957 27743
rect 3003 27737 3030 27743
rect 2590 27709 2884 27737
rect 2918 27709 2957 27737
rect 2991 27709 3030 27737
rect 2590 27703 3038 27709
rect 2590 27669 2624 27703
rect 2658 27669 2693 27703
rect 2727 27669 2762 27703
rect 2796 27669 2831 27703
rect 2865 27669 2900 27703
rect 2934 27669 2969 27703
rect 3003 27669 3038 27703
rect 2590 27663 3038 27669
rect 2590 27635 2884 27663
rect 2918 27635 2957 27663
rect 2991 27635 3030 27663
rect 2590 27601 2624 27635
rect 2658 27601 2693 27635
rect 2727 27601 2762 27635
rect 2796 27601 2831 27635
rect 2865 27629 2884 27635
rect 2934 27629 2957 27635
rect 3003 27629 3030 27635
rect 2865 27601 2900 27629
rect 2934 27601 2969 27629
rect 3003 27601 3038 27629
rect 2590 27583 3038 27601
rect 2590 27567 2884 27583
rect 2918 27567 2957 27583
rect 2991 27567 3030 27583
rect 2590 27533 2624 27567
rect 2658 27533 2693 27567
rect 2727 27533 2762 27567
rect 2796 27533 2831 27567
rect 2865 27549 2884 27567
rect 2934 27549 2957 27567
rect 3003 27549 3030 27567
rect 2865 27533 2900 27549
rect 2934 27533 2969 27549
rect 3003 27533 3038 27549
rect 2590 27503 3038 27533
rect 2590 27499 2884 27503
rect 2918 27499 2957 27503
rect 2991 27499 3030 27503
rect 2590 27465 2624 27499
rect 2658 27465 2693 27499
rect 2727 27465 2762 27499
rect 2796 27465 2831 27499
rect 2865 27469 2884 27499
rect 2934 27469 2957 27499
rect 3003 27469 3030 27499
rect 2865 27465 2900 27469
rect 2934 27465 2969 27469
rect 3003 27465 3038 27469
rect 7968 27465 8002 27907
rect 3268 27296 3316 27330
rect 3268 27262 3284 27296
rect 3268 27224 3316 27262
rect 5501 27296 5544 27329
rect 5528 27262 5544 27296
rect 5501 27223 5544 27262
rect 7083 27291 7185 27397
rect 7117 27257 7151 27291
rect 7083 27151 7185 27257
rect 7117 27117 7151 27151
rect 7083 27011 7185 27117
rect 7117 26977 7151 27011
rect 7083 26954 7185 26977
rect 7074 26922 7192 26954
rect 7074 26888 7080 26922
rect 7114 26888 7152 26922
rect 7186 26888 7192 26922
rect 7074 26871 7192 26888
rect 7074 26849 7083 26871
rect 7074 26815 7080 26849
rect 7117 26837 7151 26871
rect 7185 26849 7192 26871
rect 7114 26815 7152 26837
rect 7186 26815 7192 26849
rect 7074 26776 7192 26815
rect 7074 26742 7080 26776
rect 7114 26742 7152 26776
rect 7186 26742 7192 26776
rect 7074 26731 7192 26742
rect 7074 26703 7083 26731
rect 7074 26669 7080 26703
rect 7117 26697 7151 26731
rect 7185 26703 7192 26731
rect 7114 26669 7152 26697
rect 7186 26669 7192 26703
rect 7074 26630 7192 26669
rect 7074 26596 7080 26630
rect 7114 26596 7152 26630
rect 7186 26596 7192 26630
rect 7074 26591 7192 26596
rect 7074 26557 7083 26591
rect 7117 26557 7151 26591
rect 7185 26557 7192 26591
rect 7074 26523 7080 26557
rect 7114 26523 7152 26557
rect 7186 26523 7192 26557
rect 7074 26484 7192 26523
rect 7074 26450 7080 26484
rect 7114 26451 7152 26484
rect 7074 26417 7083 26450
rect 7117 26417 7151 26451
rect 7186 26450 7192 26484
rect 7185 26417 7192 26450
rect 7074 26411 7192 26417
rect 7074 26377 7080 26411
rect 7114 26377 7152 26411
rect 7186 26377 7192 26411
rect 7074 26338 7192 26377
rect 7074 26304 7080 26338
rect 7114 26311 7152 26338
rect 7074 26277 7083 26304
rect 7117 26277 7151 26311
rect 7186 26304 7192 26338
rect 7185 26277 7192 26304
rect 7074 26265 7192 26277
rect 7074 26231 7080 26265
rect 7114 26231 7152 26265
rect 7186 26231 7192 26265
rect 7074 26192 7192 26231
rect 7074 26158 7080 26192
rect 7114 26171 7152 26192
rect 7074 26137 7083 26158
rect 7117 26137 7151 26171
rect 7186 26158 7192 26192
rect 7185 26137 7192 26158
rect 7074 26119 7192 26137
rect 7074 26085 7080 26119
rect 7114 26085 7152 26119
rect 7186 26085 7192 26119
rect 7074 26046 7192 26085
rect 7074 26012 7080 26046
rect 7114 26031 7152 26046
rect 7074 25997 7083 26012
rect 7117 25997 7151 26031
rect 7186 26012 7192 26046
rect 7185 25997 7192 26012
rect 7074 25973 7192 25997
rect 7074 25939 7080 25973
rect 7114 25939 7152 25973
rect 7186 25939 7192 25973
rect 7074 25900 7192 25939
rect 7074 25866 7080 25900
rect 7114 25891 7152 25900
rect 7074 25857 7083 25866
rect 7117 25857 7151 25891
rect 7186 25866 7192 25900
rect 7185 25857 7192 25866
rect 7074 25827 7192 25857
rect 7074 25793 7080 25827
rect 7114 25793 7152 25827
rect 7186 25793 7192 25827
rect 7074 25754 7192 25793
rect 7074 25720 7080 25754
rect 7114 25751 7152 25754
rect 7074 25717 7083 25720
rect 7117 25717 7151 25751
rect 7186 25720 7192 25754
rect 7185 25717 7192 25720
rect 7074 25681 7192 25717
rect 7074 25647 7080 25681
rect 7114 25647 7152 25681
rect 7186 25647 7192 25681
rect 7074 25611 7192 25647
rect 7074 25608 7083 25611
rect 7074 25574 7080 25608
rect 7117 25577 7151 25611
rect 7185 25608 7192 25611
rect 7114 25574 7152 25577
rect 7186 25574 7192 25608
rect 7074 25535 7192 25574
rect 7074 25501 7080 25535
rect 7114 25501 7152 25535
rect 7186 25501 7192 25535
rect 7074 25471 7192 25501
rect 7074 25462 7083 25471
rect 7074 25428 7080 25462
rect 7117 25437 7151 25471
rect 7185 25462 7192 25471
rect 7114 25428 7152 25437
rect 7186 25428 7192 25462
rect 7074 25389 7192 25428
rect 7074 25355 7080 25389
rect 7114 25355 7152 25389
rect 7186 25355 7192 25389
rect 7074 25330 7192 25355
rect 7074 25316 7083 25330
rect 7074 25282 7080 25316
rect 7117 25296 7151 25330
rect 7185 25316 7192 25330
rect 7114 25282 7152 25296
rect 7186 25282 7192 25316
rect 7074 25243 7192 25282
rect 7074 25209 7080 25243
rect 7114 25209 7152 25243
rect 7186 25209 7192 25243
rect 7074 25189 7192 25209
rect 7074 25170 7083 25189
rect 7074 25136 7080 25170
rect 7117 25155 7151 25189
rect 7185 25170 7192 25189
rect 7114 25136 7152 25155
rect 7186 25136 7192 25170
rect 7074 25097 7192 25136
rect 7074 25063 7080 25097
rect 7114 25063 7152 25097
rect 7186 25063 7192 25097
rect 7074 25048 7192 25063
rect 7074 25024 7083 25048
rect 7074 24990 7080 25024
rect 7117 25014 7151 25048
rect 7185 25024 7192 25048
rect 7114 24990 7152 25014
rect 7186 24990 7192 25024
rect 7074 24951 7192 24990
rect 7074 24917 7080 24951
rect 7114 24917 7152 24951
rect 7186 24917 7192 24951
rect 7074 24907 7192 24917
rect 7074 24878 7083 24907
rect 7074 24844 7080 24878
rect 7117 24873 7151 24907
rect 7185 24878 7192 24907
rect 7114 24844 7152 24873
rect 7186 24844 7192 24878
rect 7074 24805 7192 24844
rect 7074 24771 7080 24805
rect 7114 24771 7152 24805
rect 7186 24771 7192 24805
rect 7074 24766 7192 24771
rect 7074 24732 7083 24766
rect 7117 24732 7151 24766
rect 7185 24732 7192 24766
rect 7074 24698 7080 24732
rect 7114 24698 7152 24732
rect 7186 24698 7192 24732
rect 7074 24659 7192 24698
rect 7074 24625 7080 24659
rect 7114 24625 7152 24659
rect 7186 24625 7192 24659
rect 7074 24591 7083 24625
rect 7117 24591 7151 24625
rect 7185 24591 7192 24625
rect 7074 24586 7192 24591
rect 7074 24552 7080 24586
rect 7114 24552 7152 24586
rect 7186 24552 7192 24586
rect 3732 24483 3766 24517
rect 3800 24483 3836 24517
rect 3870 24483 3906 24517
rect 3940 24483 3976 24517
rect 4010 24483 4046 24517
rect 4096 24483 4116 24517
rect 4169 24483 4186 24517
rect 4242 24483 4256 24517
rect 4315 24483 4326 24517
rect 4388 24483 4396 24517
rect 4461 24483 4466 24517
rect 4534 24483 4536 24517
rect 4570 24483 4573 24517
rect 4640 24483 4646 24517
rect 4709 24483 4719 24517
rect 4778 24483 4792 24517
rect 4847 24483 4865 24517
rect 4916 24483 4938 24517
rect 4985 24483 5011 24517
rect 5054 24483 5084 24517
rect 5123 24483 5157 24517
rect 5192 24483 5227 24517
rect 5264 24483 5296 24517
rect 5337 24483 5365 24517
rect 5410 24483 5434 24517
rect 5483 24483 5503 24517
rect 5556 24483 5572 24517
rect 5629 24483 5641 24517
rect 5701 24483 5710 24517
rect 5773 24483 5779 24517
rect 5845 24483 5848 24517
rect 5882 24483 5883 24517
rect 5951 24483 5955 24517
rect 6020 24483 6027 24517
rect 6089 24483 6124 24517
rect 6158 24483 6192 24517
rect 3732 24449 6192 24483
rect 3732 24415 3766 24449
rect 3800 24415 3836 24449
rect 3870 24415 3906 24449
rect 3940 24415 3976 24449
rect 4010 24415 4046 24449
rect 4080 24415 4116 24449
rect 4150 24415 4186 24449
rect 4220 24415 4256 24449
rect 4290 24415 4326 24449
rect 4360 24415 4396 24449
rect 4430 24415 4466 24449
rect 4500 24415 4536 24449
rect 4570 24415 4606 24449
rect 4640 24415 4675 24449
rect 4709 24415 4744 24449
rect 4778 24415 4813 24449
rect 4847 24415 4882 24449
rect 4916 24415 4951 24449
rect 4985 24415 5020 24449
rect 5054 24415 5089 24449
rect 5123 24415 5158 24449
rect 5192 24415 5227 24449
rect 5261 24415 5296 24449
rect 5330 24415 5365 24449
rect 5399 24415 5434 24449
rect 5468 24415 5503 24449
rect 5537 24415 5572 24449
rect 5606 24415 5641 24449
rect 5675 24415 5710 24449
rect 5744 24415 5779 24449
rect 5813 24415 5848 24449
rect 5882 24415 5917 24449
rect 5951 24415 5986 24449
rect 6020 24415 6055 24449
rect 6089 24415 6124 24449
rect 6158 24415 6192 24449
rect 3732 24381 6192 24415
rect 3732 24347 3766 24381
rect 3800 24347 3836 24381
rect 3870 24347 3906 24381
rect 3940 24347 3976 24381
rect 4010 24347 4046 24381
rect 4096 24347 4116 24381
rect 4169 24347 4186 24381
rect 4242 24347 4256 24381
rect 4315 24347 4326 24381
rect 4388 24347 4396 24381
rect 4461 24347 4466 24381
rect 4534 24347 4536 24381
rect 4570 24347 4573 24381
rect 4640 24347 4646 24381
rect 4709 24347 4719 24381
rect 4778 24347 4792 24381
rect 4847 24347 4865 24381
rect 4916 24347 4938 24381
rect 4985 24347 5011 24381
rect 5054 24347 5084 24381
rect 5123 24347 5157 24381
rect 5192 24347 5227 24381
rect 5264 24347 5296 24381
rect 5337 24347 5365 24381
rect 5410 24347 5434 24381
rect 5483 24347 5503 24381
rect 5556 24347 5572 24381
rect 5629 24347 5641 24381
rect 5701 24347 5710 24381
rect 5773 24347 5779 24381
rect 5845 24347 5848 24381
rect 5882 24347 5883 24381
rect 5951 24347 5955 24381
rect 6020 24347 6027 24381
rect 6089 24347 6124 24381
rect 6158 24347 6192 24381
rect 7074 24513 7192 24552
rect 7074 24479 7080 24513
rect 7114 24484 7152 24513
rect 7074 24450 7083 24479
rect 7117 24450 7151 24484
rect 7186 24479 7192 24513
rect 7185 24450 7192 24479
rect 7074 24440 7192 24450
rect 7074 24406 7080 24440
rect 7114 24406 7152 24440
rect 7186 24406 7192 24440
rect 7074 24367 7192 24406
rect 7074 24333 7080 24367
rect 7114 24343 7152 24367
rect 7074 24309 7083 24333
rect 7117 24309 7151 24343
rect 7186 24333 7192 24367
rect 7185 24309 7192 24333
rect 7074 24294 7192 24309
rect 7074 24260 7080 24294
rect 7114 24260 7152 24294
rect 7186 24260 7192 24294
rect 7074 24221 7192 24260
rect 7074 24187 7080 24221
rect 7114 24202 7152 24221
rect 7074 24168 7083 24187
rect 7117 24168 7151 24202
rect 7186 24187 7192 24221
rect 7185 24168 7192 24187
rect 7074 24148 7192 24168
rect 7074 24114 7080 24148
rect 7114 24114 7152 24148
rect 7186 24114 7192 24148
rect 7074 24075 7192 24114
rect 7074 24041 7080 24075
rect 7114 24061 7152 24075
rect 7074 24027 7083 24041
rect 7117 24027 7151 24061
rect 7186 24041 7192 24075
rect 7185 24027 7192 24041
rect 7074 24002 7192 24027
rect 7074 23968 7080 24002
rect 7114 23968 7152 24002
rect 7186 23968 7192 24002
rect 7074 23929 7192 23968
rect 7074 23895 7080 23929
rect 7114 23920 7152 23929
rect 7074 23886 7083 23895
rect 7117 23886 7151 23920
rect 7186 23895 7192 23929
rect 7185 23886 7192 23895
rect 7074 23856 7192 23886
rect 7074 23822 7080 23856
rect 7114 23822 7152 23856
rect 7186 23822 7192 23856
rect 7074 23782 7192 23822
rect 7074 23748 7080 23782
rect 7114 23779 7152 23782
rect 7074 23745 7083 23748
rect 7117 23745 7151 23779
rect 7186 23748 7192 23782
rect 7185 23745 7192 23748
rect 7074 23708 7192 23745
rect 7074 23674 7080 23708
rect 7114 23674 7152 23708
rect 7186 23674 7192 23708
rect 7074 23638 7192 23674
rect 7074 23634 7083 23638
rect 7074 23600 7080 23634
rect 7117 23604 7151 23638
rect 7185 23634 7192 23638
rect 7114 23600 7152 23604
rect 7186 23600 7192 23634
rect 7074 23560 7192 23600
rect 7074 23526 7080 23560
rect 7114 23526 7152 23560
rect 7186 23526 7192 23560
rect 7074 23497 7192 23526
rect 7074 23486 7083 23497
rect 7074 23452 7080 23486
rect 7117 23463 7151 23497
rect 7185 23486 7192 23497
rect 7114 23452 7152 23463
rect 7186 23452 7192 23486
rect 7074 23412 7192 23452
rect 7074 23378 7080 23412
rect 7114 23378 7152 23412
rect 7186 23378 7192 23412
rect 7074 23356 7192 23378
rect 7074 23322 7083 23356
rect 7117 23322 7151 23356
rect 7185 23322 7192 23356
rect 7074 23256 7192 23322
rect 6056 23246 6067 23256
rect 7757 23246 7768 23256
rect 6055 22790 6067 23246
rect 7757 23212 7792 23246
rect 7826 23212 7934 23246
rect 7968 23212 8002 23246
rect 7757 23144 8002 23212
rect 7757 23110 7792 23144
rect 7826 23110 7934 23144
rect 7968 23110 8002 23144
rect 7757 23042 8002 23110
rect 7757 23008 7792 23042
rect 7826 23008 7934 23042
rect 7968 23008 8002 23042
rect 7757 22940 8002 23008
rect 7757 22906 7792 22940
rect 7826 22906 7934 22940
rect 7968 22906 8002 22940
rect 7757 22838 8002 22906
rect 7757 22804 7792 22838
rect 7826 22804 7934 22838
rect 7968 22804 8002 22838
rect 7757 22790 8002 22804
rect 6055 22751 8002 22790
rect 6055 22717 6067 22751
rect 6101 22736 6139 22751
rect 6123 22717 6139 22736
rect 6173 22717 6211 22751
rect 6245 22736 6283 22751
rect 6264 22717 6283 22736
rect 6317 22717 6355 22751
rect 6389 22736 6427 22751
rect 6406 22717 6427 22736
rect 6461 22717 6499 22751
rect 6533 22736 6571 22751
rect 6548 22717 6571 22736
rect 6605 22717 6643 22751
rect 6677 22736 6715 22751
rect 6690 22717 6715 22736
rect 6749 22717 6787 22751
rect 6821 22736 6859 22751
rect 6832 22717 6859 22736
rect 6893 22717 6931 22751
rect 6965 22736 7003 22751
rect 6974 22717 7003 22736
rect 7037 22717 7075 22751
rect 7109 22736 7147 22751
rect 7116 22717 7147 22736
rect 7181 22717 7219 22751
rect 7253 22736 7291 22751
rect 7258 22717 7291 22736
rect 7325 22717 7363 22751
rect 7397 22736 7435 22751
rect 7400 22717 7435 22736
rect 7469 22717 7507 22751
rect 7541 22736 7579 22751
rect 7542 22717 7579 22736
rect 7613 22736 7651 22751
rect 7613 22717 7650 22736
rect 7685 22717 7723 22751
rect 7757 22736 8002 22751
rect 7757 22717 7792 22736
rect 6055 22702 6089 22717
rect 6123 22702 6230 22717
rect 6264 22702 6372 22717
rect 6406 22702 6514 22717
rect 6548 22702 6656 22717
rect 6690 22702 6798 22717
rect 6832 22702 6940 22717
rect 6974 22702 7082 22717
rect 7116 22702 7224 22717
rect 7258 22702 7366 22717
rect 7400 22702 7508 22717
rect 7542 22702 7650 22717
rect 7684 22702 7792 22717
rect 7826 22702 7934 22736
rect 7968 22702 8002 22736
rect 6055 22678 8002 22702
rect 6055 22644 6067 22678
rect 6101 22644 6139 22678
rect 6173 22644 6211 22678
rect 6245 22644 6283 22678
rect 6317 22644 6355 22678
rect 6389 22644 6427 22678
rect 6461 22644 6499 22678
rect 6533 22644 6571 22678
rect 6605 22644 6643 22678
rect 6677 22644 6715 22678
rect 6749 22644 6787 22678
rect 6821 22644 6859 22678
rect 6893 22644 6931 22678
rect 6965 22644 7003 22678
rect 7037 22644 7075 22678
rect 7109 22644 7147 22678
rect 7181 22644 7219 22678
rect 7253 22644 7291 22678
rect 7325 22644 7363 22678
rect 7397 22644 7435 22678
rect 7469 22644 7507 22678
rect 7541 22644 7579 22678
rect 7613 22644 7651 22678
rect 7685 22644 7723 22678
rect 7757 22644 8002 22678
rect 6055 22634 8002 22644
rect 6055 22605 6089 22634
rect 6123 22605 6230 22634
rect 6264 22605 6372 22634
rect 6406 22605 6514 22634
rect 6548 22605 6656 22634
rect 6690 22605 6798 22634
rect 6832 22605 6940 22634
rect 6974 22605 7082 22634
rect 7116 22605 7224 22634
rect 7258 22605 7366 22634
rect 7400 22605 7508 22634
rect 7542 22605 7650 22634
rect 7684 22605 7792 22634
rect 6055 22571 6067 22605
rect 6123 22600 6139 22605
rect 6101 22571 6139 22600
rect 6173 22571 6211 22605
rect 6264 22600 6283 22605
rect 6245 22571 6283 22600
rect 6317 22571 6355 22605
rect 6406 22600 6427 22605
rect 6389 22571 6427 22600
rect 6461 22571 6499 22605
rect 6548 22600 6571 22605
rect 6533 22571 6571 22600
rect 6605 22571 6643 22605
rect 6690 22600 6715 22605
rect 6677 22571 6715 22600
rect 6749 22571 6787 22605
rect 6832 22600 6859 22605
rect 6821 22571 6859 22600
rect 6893 22571 6931 22605
rect 6974 22600 7003 22605
rect 6965 22571 7003 22600
rect 7037 22571 7075 22605
rect 7116 22600 7147 22605
rect 7109 22571 7147 22600
rect 7181 22571 7219 22605
rect 7258 22600 7291 22605
rect 7253 22571 7291 22600
rect 7325 22571 7363 22605
rect 7400 22600 7435 22605
rect 7397 22571 7435 22600
rect 7469 22571 7507 22605
rect 7542 22600 7579 22605
rect 7541 22571 7579 22600
rect 7613 22600 7650 22605
rect 7613 22571 7651 22600
rect 7685 22571 7723 22605
rect 7757 22600 7792 22605
rect 7826 22600 7934 22634
rect 7968 22600 8002 22634
rect 7757 22571 8002 22600
rect 6055 22532 8002 22571
rect 6055 22498 6067 22532
rect 6123 22498 6139 22532
rect 6173 22498 6211 22532
rect 6264 22498 6283 22532
rect 6317 22498 6355 22532
rect 6406 22498 6427 22532
rect 6461 22498 6499 22532
rect 6548 22498 6571 22532
rect 6605 22498 6643 22532
rect 6690 22498 6715 22532
rect 6749 22498 6787 22532
rect 6832 22498 6859 22532
rect 6893 22498 6931 22532
rect 6974 22498 7003 22532
rect 7037 22498 7075 22532
rect 7116 22498 7147 22532
rect 7181 22498 7219 22532
rect 7258 22498 7291 22532
rect 7325 22498 7363 22532
rect 7400 22498 7435 22532
rect 7469 22498 7507 22532
rect 7542 22498 7579 22532
rect 7613 22498 7650 22532
rect 7685 22498 7723 22532
rect 7757 22498 7792 22532
rect 7826 22498 7934 22532
rect 7968 22498 8002 22532
rect 6373 19869 6407 19885
rect 6373 19798 6407 19835
rect 6373 19727 6407 19764
rect 6373 19655 6407 19660
rect 7006 19625 7052 19659
rect 7086 19625 7132 19659
rect 7166 19625 7212 19659
rect 7246 19625 7292 19659
rect 7326 19625 7372 19659
rect 7406 19625 7451 19659
rect 7485 19625 7530 19659
rect 7716 19622 7750 19632
rect 6373 19583 6407 19588
rect 6373 19511 6407 19516
rect 7624 19602 7658 19614
rect 7624 19508 7658 19564
rect 7150 19469 7199 19503
rect 7233 19469 7282 19503
rect 7316 19469 7365 19503
rect 7399 19469 7448 19503
rect 7482 19469 7530 19503
rect 6373 19439 6407 19444
rect 6373 19367 6407 19371
rect 7624 19414 7658 19469
rect 7624 19358 7658 19374
rect 7716 19554 7750 19560
rect 7716 19486 7750 19488
rect 7716 19450 7750 19452
rect 7716 19378 7750 19384
rect 6373 19317 6407 19333
rect 7006 19313 7058 19347
rect 7092 19313 7144 19347
rect 7178 19313 7230 19347
rect 7264 19313 7316 19347
rect 7350 19313 7402 19347
rect 7716 19306 7750 19316
rect 7624 19286 7658 19302
rect 6373 19245 6407 19261
rect 6373 19174 6407 19197
rect 7624 19216 7658 19246
rect 7178 19157 7222 19191
rect 7256 19157 7299 19191
rect 7333 19157 7376 19191
rect 7410 19157 7453 19191
rect 7487 19157 7530 19191
rect 6373 19103 6407 19122
rect 6373 19031 6407 19047
rect 7624 19146 7658 19172
rect 7624 19076 7658 19098
rect 7006 19001 7058 19035
rect 7092 19001 7144 19035
rect 7178 19001 7230 19035
rect 7264 19001 7316 19035
rect 7350 19001 7402 19035
rect 7624 19006 7658 19024
rect 6373 18959 6407 18972
rect 6373 18887 6407 18897
rect 7624 18936 7658 18950
rect 7178 18845 7222 18879
rect 7256 18845 7299 18879
rect 7333 18845 7376 18879
rect 7410 18845 7453 18879
rect 7487 18845 7530 18879
rect 7624 18866 7658 18876
rect 6373 18815 6407 18822
rect 6373 18743 6407 18747
rect 7624 18796 7658 18802
rect 7624 18726 7658 18728
rect 6373 18693 6407 18709
rect 7006 18689 7058 18723
rect 7092 18689 7144 18723
rect 7178 18689 7230 18723
rect 7264 18689 7316 18723
rect 7350 18689 7402 18723
rect 7624 18688 7658 18692
rect 6373 18621 6407 18637
rect 6373 18553 6407 18580
rect 7624 18614 7658 18622
rect 7178 18533 7222 18567
rect 7256 18533 7299 18567
rect 7333 18533 7376 18567
rect 7410 18533 7453 18567
rect 7487 18533 7530 18567
rect 7624 18540 7658 18552
rect 6373 18503 6407 18508
rect 7624 18466 7658 18481
rect 7006 18377 7058 18411
rect 7092 18377 7144 18411
rect 7178 18377 7230 18411
rect 7264 18377 7316 18411
rect 7350 18377 7402 18411
rect 7624 18392 7658 18410
rect 7624 18318 7658 18339
rect 7178 18221 7222 18255
rect 7256 18221 7299 18255
rect 7333 18221 7376 18255
rect 7410 18221 7453 18255
rect 7487 18221 7530 18255
rect 7624 18244 7658 18268
rect 7624 18170 7658 18197
rect 7624 18110 7658 18126
rect 7716 19234 7750 19248
rect 7716 19162 7750 19180
rect 7716 19090 7750 19112
rect 7716 19018 7750 19044
rect 7716 18946 7750 18976
rect 7716 18874 7750 18908
rect 7716 18806 7750 18840
rect 7716 18738 7750 18768
rect 7716 18670 7750 18696
rect 7716 18602 7750 18624
rect 7716 18534 7750 18552
rect 7716 18466 7750 18480
rect 7716 18398 7750 18407
rect 7716 18330 7750 18334
rect 7716 18295 7750 18296
rect 7716 18222 7750 18228
rect 7716 18149 7750 18160
rect 7006 18065 7058 18099
rect 7092 18065 7144 18099
rect 7178 18065 7230 18099
rect 7264 18065 7316 18099
rect 7350 18065 7402 18099
rect 7716 18076 7750 18092
rect 7624 18040 7658 18054
rect 7624 17969 7658 18004
rect 7178 17909 7222 17943
rect 7256 17909 7299 17943
rect 7333 17909 7376 17943
rect 7410 17909 7453 17943
rect 7487 17909 7530 17943
rect 7624 17919 7658 17934
rect 7716 18003 7750 18024
rect 7716 17930 7750 17956
rect 7716 17857 7750 17888
rect 7006 17799 7052 17833
rect 7086 17799 7132 17833
rect 7166 17799 7212 17833
rect 7246 17799 7292 17833
rect 7326 17799 7372 17833
rect 7406 17799 7451 17833
rect 7485 17799 7530 17833
rect 7624 17776 7658 17788
rect 7624 17680 7658 17738
rect 7150 17643 7194 17677
rect 7228 17643 7271 17677
rect 7305 17643 7348 17677
rect 7382 17643 7425 17677
rect 7459 17643 7502 17677
rect 7624 17583 7658 17643
rect 7624 17532 7658 17548
rect 7716 17786 7750 17820
rect 7716 17718 7750 17750
rect 7716 17650 7750 17677
rect 7716 17582 7750 17604
rect 7006 17487 7058 17521
rect 7092 17487 7144 17521
rect 7178 17487 7230 17521
rect 7264 17487 7316 17521
rect 7350 17487 7402 17521
rect 7716 17514 7750 17531
rect 7624 17468 7658 17476
rect 7624 17394 7658 17426
rect 7178 17331 7222 17365
rect 7256 17331 7299 17365
rect 7333 17331 7376 17365
rect 7410 17331 7453 17365
rect 7487 17331 7530 17365
rect 7624 17320 7658 17356
rect 7624 17250 7658 17285
rect 7006 17175 7058 17209
rect 7092 17175 7144 17209
rect 7178 17175 7230 17209
rect 7264 17175 7316 17209
rect 7350 17175 7402 17209
rect 7624 17180 7658 17210
rect 7624 17110 7658 17135
rect 7178 17019 7222 17053
rect 7256 17019 7299 17053
rect 7333 17019 7376 17053
rect 7410 17019 7453 17053
rect 7487 17019 7530 17053
rect 7624 17040 7658 17060
rect 7624 16970 7658 16985
rect 7624 16900 7658 16910
rect 7006 16863 7058 16897
rect 7092 16863 7144 16897
rect 7178 16863 7230 16897
rect 7264 16863 7316 16897
rect 7350 16863 7402 16897
rect 7624 16830 7658 16835
rect 7624 16794 7658 16796
rect 7178 16707 7222 16741
rect 7256 16707 7299 16741
rect 7333 16707 7376 16741
rect 7410 16707 7453 16741
rect 7487 16707 7530 16741
rect 7624 16719 7658 16726
rect 7624 16644 7658 16655
rect 7006 16551 7058 16585
rect 7092 16551 7144 16585
rect 7178 16551 7230 16585
rect 7264 16551 7316 16585
rect 7350 16551 7402 16585
rect 7624 16569 7658 16584
rect 7624 16494 7658 16513
rect 7178 16395 7222 16429
rect 7256 16395 7299 16429
rect 7333 16395 7376 16429
rect 7410 16395 7453 16429
rect 7487 16395 7530 16429
rect 7624 16419 7658 16442
rect 7624 16344 7658 16371
rect 7624 16284 7658 16300
rect 7716 17446 7750 17458
rect 7716 17378 7750 17385
rect 7716 17310 7750 17312
rect 7716 17273 7750 17276
rect 7716 17200 7750 17208
rect 7716 17127 7750 17140
rect 7716 17054 7750 17072
rect 7716 16981 7750 17004
rect 7716 16908 7750 16936
rect 7716 16835 7750 16868
rect 7716 16766 7750 16800
rect 7716 16698 7750 16728
rect 7716 16630 7750 16655
rect 7716 16562 7750 16582
rect 7716 16494 7750 16509
rect 7716 16426 7750 16436
rect 7716 16358 7750 16363
rect 7006 16239 7058 16273
rect 7092 16239 7144 16273
rect 7178 16239 7230 16273
rect 7264 16239 7316 16273
rect 7350 16239 7402 16273
rect 7716 16251 7750 16256
rect 7624 16216 7658 16228
rect 7624 16144 7658 16178
rect 7178 16083 7222 16117
rect 7256 16083 7299 16117
rect 7333 16083 7376 16117
rect 7410 16083 7453 16117
rect 7487 16083 7530 16117
rect 7624 16092 7658 16108
rect 7716 16178 7750 16188
rect 7716 16105 7750 16120
rect 7716 16032 7750 16052
rect 7006 15973 7052 16007
rect 7086 15973 7132 16007
rect 7166 15973 7212 16007
rect 7246 15973 7292 16007
rect 7326 15973 7372 16007
rect 7406 15973 7451 16007
rect 7485 15973 7530 16007
rect 7624 15950 7658 15962
rect 7624 15861 7658 15912
rect 7150 15817 7194 15851
rect 7228 15817 7271 15851
rect 7305 15817 7348 15851
rect 7382 15817 7425 15851
rect 7459 15817 7502 15851
rect 7624 15772 7658 15817
rect 7624 15706 7658 15722
rect 7716 15959 7750 15984
rect 7716 15886 7750 15916
rect 7716 15814 7750 15848
rect 7716 15746 7750 15779
rect 7006 15661 7058 15695
rect 7092 15661 7144 15695
rect 7178 15661 7230 15695
rect 7264 15661 7316 15695
rect 7350 15661 7402 15695
rect 7716 15678 7750 15706
rect 7624 15634 7658 15650
rect 7624 15564 7658 15596
rect 7178 15505 7222 15539
rect 7256 15505 7299 15539
rect 7333 15505 7376 15539
rect 7410 15505 7453 15539
rect 7487 15505 7530 15539
rect 7624 15494 7658 15522
rect 7624 15424 7658 15448
rect 7006 15349 7058 15383
rect 7092 15349 7144 15383
rect 7178 15349 7230 15383
rect 7264 15349 7316 15383
rect 7350 15349 7402 15383
rect 7624 15354 7658 15374
rect 7624 15284 7658 15300
rect 7178 15193 7222 15227
rect 7256 15193 7299 15227
rect 7333 15193 7376 15227
rect 7410 15193 7453 15227
rect 7487 15193 7530 15227
rect 7624 15214 7658 15226
rect 7624 15144 7658 15152
rect 7624 15074 7658 15078
rect 7006 15037 7058 15071
rect 7092 15037 7144 15071
rect 7178 15037 7230 15071
rect 7264 15037 7316 15071
rect 7350 15037 7402 15071
rect 7624 15038 7658 15040
rect 7624 14964 7658 14970
rect 7178 14881 7222 14915
rect 7256 14881 7299 14915
rect 7333 14881 7376 14915
rect 7410 14881 7453 14915
rect 7487 14881 7530 14915
rect 7624 14890 7658 14900
rect 7624 14816 7658 14829
rect 7006 14725 7058 14759
rect 7092 14725 7144 14759
rect 7178 14725 7230 14759
rect 7264 14725 7316 14759
rect 7350 14725 7402 14759
rect 7624 14742 7658 14758
rect 7624 14668 7658 14687
rect 7178 14569 7222 14603
rect 7256 14569 7299 14603
rect 7333 14569 7376 14603
rect 7410 14569 7453 14603
rect 7487 14569 7530 14603
rect 7624 14593 7658 14616
rect 7624 14518 7658 14545
rect 7624 14458 7658 14474
rect 7716 15610 7750 15633
rect 7716 15542 7750 15560
rect 7716 15474 7750 15487
rect 7716 15406 7750 15414
rect 7716 15338 7750 15341
rect 7716 15302 7750 15304
rect 7716 15229 7750 15236
rect 7716 15156 7750 15168
rect 7716 15083 7750 15100
rect 7716 15010 7750 15032
rect 7716 14937 7750 14964
rect 7716 14864 7750 14896
rect 7716 14794 7750 14828
rect 7716 14726 7750 14757
rect 7716 14658 7750 14684
rect 7716 14590 7750 14611
rect 7716 14522 7750 14538
rect 7716 14454 7750 14465
rect 7006 14413 7058 14447
rect 7092 14413 7144 14447
rect 7178 14413 7230 14447
rect 7264 14413 7316 14447
rect 7350 14413 7402 14447
rect 7624 14390 7658 14402
rect 7624 14318 7658 14352
rect 7178 14257 7222 14291
rect 7256 14257 7299 14291
rect 7333 14257 7376 14291
rect 7410 14257 7453 14291
rect 7487 14257 7530 14291
rect 7624 14267 7658 14283
rect 7716 14386 7750 14392
rect 7716 14318 7750 14319
rect 7716 14280 7750 14284
rect 6364 14040 6398 14064
rect 7061 14042 7106 14076
rect 7140 14042 7185 14076
rect 7564 14042 7629 14076
rect 6364 13971 6398 14003
rect 6833 14015 6867 14031
rect 6364 13902 6398 13930
rect 6364 13833 6398 13857
rect 6364 13764 6398 13783
rect 6364 13695 6398 13709
rect 6364 13625 6398 13635
rect 6364 13555 6398 13561
rect 6364 13485 6398 13487
rect 6364 13447 6398 13451
rect 6670 13982 6704 13998
rect 6670 13911 6704 13945
rect 6670 13840 6704 13864
rect 6670 13768 6704 13783
rect 6670 13696 6704 13701
rect 6670 13653 6704 13662
rect 6833 13945 6867 13981
rect 7815 14019 7849 14031
rect 7815 13945 7849 13981
rect 6833 13880 6867 13911
rect 7061 13886 7169 13920
rect 7304 13902 7338 13911
rect 6833 13807 6867 13842
rect 7457 13886 7526 13920
rect 7560 13886 7629 13920
rect 7304 13834 7338 13839
rect 7304 13766 7338 13767
rect 6833 13738 6867 13739
rect 6993 13730 7035 13764
rect 7069 13730 7110 13764
rect 7144 13730 7185 13764
rect 7815 13876 7849 13897
rect 7815 13807 7849 13809
rect 6833 13669 6867 13704
rect 6833 13619 6867 13631
rect 7304 13729 7338 13732
rect 7555 13730 7629 13764
rect 7815 13754 7849 13773
rect 7304 13657 7338 13664
rect 6670 13571 6704 13590
rect 7061 13574 7169 13608
rect 7815 13669 7849 13704
rect 7815 13619 7849 13631
rect 7304 13585 7338 13596
rect 6670 13489 6704 13518
rect 6670 13430 6704 13446
rect 6833 13554 6867 13563
rect 6833 13482 6867 13513
rect 7457 13574 7526 13608
rect 7560 13574 7629 13608
rect 7304 13513 7338 13528
rect 6364 13373 6398 13381
rect 6833 13410 6867 13441
rect 6971 13418 7016 13452
rect 7050 13418 7095 13452
rect 7304 13441 7338 13460
rect 7815 13490 7849 13513
rect 2829 13315 6114 13371
rect 6364 13299 6398 13311
rect 6364 13225 6398 13241
rect 6364 13151 6398 13171
rect 6364 13077 6398 13101
rect 6364 13003 6398 13031
rect 6364 12929 6398 12961
rect 6364 12855 6398 12891
rect 6364 12785 6398 12821
rect 6670 13358 6704 13374
rect 6670 13287 6704 13314
rect 6670 13216 6704 13233
rect 6670 13144 6704 13152
rect 6670 13105 6704 13110
rect 6670 13024 6704 13038
rect 6833 13338 6867 13369
rect 6833 13266 6867 13297
rect 7541 13418 7608 13452
rect 7642 13418 7709 13452
rect 7304 13369 7338 13392
rect 7304 13297 7338 13324
rect 7061 13262 7100 13296
rect 7134 13262 7173 13296
rect 7815 13417 7849 13441
rect 7815 13344 7849 13369
rect 6833 13194 6867 13225
rect 6833 13121 6867 13153
rect 7457 13262 7526 13296
rect 7560 13262 7629 13296
rect 7815 13270 7849 13297
rect 7304 13225 7338 13255
rect 7304 13152 7338 13186
rect 6971 13106 7016 13140
rect 7050 13106 7095 13140
rect 7815 13196 7849 13225
rect 6833 13048 6867 13082
rect 6833 12995 6867 13011
rect 7304 13082 7338 13117
rect 7539 13106 7607 13140
rect 7641 13106 7709 13140
rect 7815 13122 7849 13153
rect 7304 13013 7338 13045
rect 6670 12943 6704 12966
rect 7061 12950 7100 12984
rect 7134 12950 7173 12984
rect 7815 13048 7849 13082
rect 7815 12995 7849 13011
rect 6670 12861 6704 12894
rect 7304 12944 7338 12972
rect 7473 12950 7522 12984
rect 7556 12950 7605 12984
rect 7639 12950 7687 12984
rect 7304 12875 7338 12899
rect 7147 12840 7185 12874
rect 6670 12806 6704 12822
rect 6943 12813 6977 12829
rect 6943 12754 6977 12779
rect 6364 12715 6398 12747
rect 6364 12645 6398 12673
rect 6670 12734 6704 12750
rect 6670 12666 6704 12698
rect 7457 12840 7495 12874
rect 7304 12806 7338 12826
rect 7304 12737 7338 12753
rect 6943 12682 6977 12711
rect 7057 12690 7095 12724
rect 7665 12813 7699 12829
rect 7665 12760 7699 12779
rect 7533 12690 7571 12724
rect 7304 12679 7338 12680
rect 7665 12688 7699 12711
rect 6670 12616 6704 12626
rect 6364 12587 6398 12599
rect 6364 12456 6388 12490
rect 6422 12456 6458 12490
rect 6492 12456 6528 12490
rect 6582 12456 6598 12490
rect 6659 12456 6668 12490
rect 6735 12456 6738 12490
rect 6772 12456 6777 12490
rect 6842 12456 6853 12490
rect 6912 12456 6929 12490
rect 6982 12456 7005 12490
rect 7052 12456 7081 12490
rect 7121 12456 7156 12490
rect 7191 12456 7225 12490
rect 7267 12456 7294 12490
rect 7343 12456 7363 12490
rect 7419 12456 7432 12490
rect 7495 12456 7501 12490
rect 7535 12456 7537 12490
rect 7604 12456 7613 12490
rect 6392 12299 6426 12337
rect 6542 12299 6576 12337
rect 6672 12167 6706 12265
rect 6798 12263 6832 12325
rect 6798 12167 6832 12229
rect 6964 12167 6998 12265
rect 7120 12263 7154 12325
rect 7120 12167 7154 12229
rect 7276 12203 7310 12265
rect 6397 12095 6413 12129
rect 6447 12095 6472 12129
rect 6515 12095 6544 12129
rect 7276 12107 7310 12169
rect 7432 12263 7466 12325
rect 7432 12167 7466 12229
rect 7588 12203 7622 12265
rect 7588 12107 7622 12169
rect 7744 12203 7778 12265
rect 7744 12107 7778 12169
rect 6697 11945 6713 11979
rect 6758 11945 6782 11979
rect 6842 11945 6851 11979
rect 6885 11945 6892 11979
rect 6954 11945 6975 11979
rect 7023 11945 7058 11979
rect 7093 11945 7109 11979
rect 7165 11945 7181 11979
rect 7238 11945 7252 11979
rect 7286 11945 7289 11979
rect 7357 11945 7373 11979
rect 7429 11945 7457 11979
rect 7501 11945 7539 11979
rect 7575 11945 7611 11979
rect 7645 11945 7683 11979
rect 7717 11945 7733 11979
rect 5004 11138 5018 11172
rect 5054 11138 5088 11172
rect 5124 11138 5138 11172
rect 5304 11138 5320 11172
rect 5361 11138 5389 11172
rect 5438 11138 5458 11172
rect 5515 11138 5527 11172
rect 5592 11138 5596 11172
rect 5630 11138 5634 11172
rect 5700 11138 5716 11172
rect 5772 11138 5788 11172
rect 5837 11138 5859 11172
rect 5925 11138 5930 11172
rect 5964 11138 5979 11172
rect 6036 11138 6067 11172
rect 6108 11138 6146 11172
rect 6189 11138 6218 11172
rect 6252 11138 6290 11172
rect 6324 11138 6340 11172
rect 3144 11084 3154 11118
rect 3194 11084 3226 11118
rect 3262 11084 3278 11118
rect 3334 11084 3350 11118
rect 3389 11084 3422 11118
rect 3471 11084 3494 11118
rect 3552 11084 3566 11118
rect 3633 11084 3638 11118
rect 3672 11084 3680 11118
rect 3744 11084 3761 11118
rect 3815 11084 3842 11118
rect 3886 11084 3902 11118
rect 3958 11084 3974 11118
rect 4017 11084 4046 11118
rect 4099 11084 4118 11118
rect 4181 11084 4190 11118
rect 4224 11084 4229 11118
rect 4296 11084 4311 11118
rect 4368 11084 4392 11118
rect 4439 11084 4473 11118
rect 4510 11084 4526 11118
rect 4999 10930 5033 10968
rect 5149 10930 5183 10968
rect 5272 10970 5306 11016
rect 5415 10993 5449 11044
rect 5415 10908 5449 10959
rect 5571 10970 5605 11044
rect 5727 10917 5761 10968
rect 5883 10998 5917 11044
rect 5727 10832 5761 10883
rect 3115 10778 3127 10812
rect 3173 10778 3202 10812
rect 3243 10778 3276 10812
rect 3313 10778 3349 10812
rect 3384 10778 3419 10812
rect 3458 10778 3489 10812
rect 3532 10778 3559 10812
rect 3606 10778 3629 10812
rect 3680 10778 3699 10812
rect 3754 10778 3769 10812
rect 3828 10778 3839 10812
rect 3902 10778 3909 10812
rect 3976 10778 3979 10812
rect 4013 10778 4016 10812
rect 4083 10778 4090 10812
rect 4153 10778 4164 10812
rect 4223 10778 4238 10812
rect 4292 10778 4312 10812
rect 4361 10778 4386 10812
rect 4430 10778 4460 10812
rect 4499 10778 4534 10812
rect 4568 10778 4592 10812
rect 6039 10916 6073 10968
rect 6195 10998 6229 11044
rect 6717 11060 6751 11061
rect 6870 11042 6908 11076
rect 7078 11057 7112 11071
rect 6039 10831 6073 10882
rect 6351 10926 6385 10968
rect 6351 10850 6385 10892
rect 6717 10987 6751 11003
rect 7078 10987 7112 11021
rect 7078 10937 7112 10951
rect 6717 10914 6751 10934
rect 6870 10892 6908 10926
rect 6717 10841 6751 10865
rect 6717 10768 6751 10796
rect 6957 10784 7022 10818
rect 7056 10784 7122 10818
rect 4988 10680 4989 10714
rect 5046 10680 5062 10714
rect 5115 10680 5135 10714
rect 5184 10680 5208 10714
rect 5253 10680 5281 10714
rect 5322 10680 5354 10714
rect 5391 10680 5426 10714
rect 5461 10680 5495 10714
rect 5534 10680 5564 10714
rect 5606 10680 5633 10714
rect 5678 10680 5701 10714
rect 5750 10680 5769 10714
rect 5822 10680 5837 10714
rect 5894 10680 5905 10714
rect 5966 10680 5973 10714
rect 6038 10680 6041 10714
rect 6075 10680 6076 10714
rect 6143 10680 6148 10714
rect 6211 10680 6220 10714
rect 6717 10695 6751 10727
rect 7228 10755 7262 10771
rect 7228 10686 7262 10692
rect 6717 10623 6751 10658
rect 6870 10626 6938 10660
rect 6972 10626 7040 10660
rect 7228 10651 7262 10652
rect 6717 10554 6751 10588
rect 6717 10485 6751 10515
rect 7228 10576 7262 10583
rect 6956 10470 7040 10504
rect 7228 10501 7262 10514
rect 6717 10416 6751 10443
rect 6717 10347 6751 10371
rect 7228 10426 7262 10445
rect 7228 10359 7262 10375
rect 6870 10314 6938 10348
rect 6972 10314 7040 10348
rect 6717 10278 6751 10299
rect 6717 10209 6751 10227
rect 7228 10287 7262 10303
rect 7228 10216 7262 10247
rect 6955 10158 7021 10192
rect 7055 10158 7122 10192
rect 6717 10140 6751 10155
rect 6717 10071 6751 10083
rect 7228 10145 7262 10169
rect 7228 10073 7262 10091
rect 6717 10002 6751 10011
rect 6870 10002 6938 10036
rect 6972 10002 7040 10036
rect 6717 9933 6751 9939
rect 7228 10001 7262 10014
rect 7228 9929 7262 9937
rect 7228 9894 7262 9895
rect 6717 9864 6751 9867
rect 6958 9846 7023 9880
rect 7057 9846 7122 9880
rect 7228 9857 7262 9860
rect 6717 9829 6751 9830
rect 3105 9769 6439 9827
rect 6717 9726 6751 9761
rect 7228 9785 7262 9823
rect 7228 9735 7262 9751
rect 6870 9690 6938 9724
rect 6972 9690 7040 9724
rect 6717 9657 6751 9668
rect 6717 9588 6751 9595
rect 7228 9663 7262 9679
rect 7228 9592 7262 9614
rect 6958 9534 7023 9568
rect 7057 9534 7122 9568
rect 6717 9519 6751 9522
rect 6717 9483 6751 9485
rect 6717 9410 6751 9416
rect 7228 9521 7262 9537
rect 7228 9449 7262 9459
rect 6870 9378 6938 9412
rect 6972 9378 7040 9412
rect 6717 9337 6751 9347
rect 6717 9264 6751 9278
rect 7228 9377 7262 9381
rect 7228 9337 7262 9343
rect 7228 9259 7262 9271
rect 6958 9222 7023 9256
rect 7057 9222 7122 9256
rect 6717 9191 6751 9209
rect 6717 9119 6751 9141
rect 7228 9181 7262 9199
rect 7228 9111 7262 9127
rect 6717 9047 6751 9073
rect 6870 9066 6938 9100
rect 6972 9066 7040 9100
rect 6717 8975 6751 9005
rect 7228 9039 7262 9055
rect 7228 8970 7262 8999
rect 6717 8903 6751 8937
rect 6958 8910 7023 8944
rect 7057 8910 7122 8944
rect 6717 8835 6751 8869
rect 6717 8767 6751 8797
rect 7228 8901 7262 8912
rect 7228 8859 7262 8867
rect 6870 8754 6938 8788
rect 6972 8754 7040 8788
rect 7228 8772 7262 8798
rect 6717 8699 6751 8725
rect 6717 8631 6751 8653
rect 7228 8694 7262 8729
rect 7228 8644 7262 8651
rect 6958 8598 7023 8632
rect 7057 8598 7122 8632
rect 6717 8563 6751 8581
rect 6717 8495 6751 8509
rect 6945 8488 6983 8522
rect 7078 8461 7112 8477
rect 7078 8393 7112 8400
rect 6870 8332 6908 8366
rect 7078 8327 7112 8359
rect 2842 7920 6744 7926
rect 2842 7886 2874 7920
rect 2908 7886 2948 7920
rect 2982 7886 3022 7920
rect 3056 7886 3096 7920
rect 3130 7886 3170 7920
rect 3204 7886 3244 7920
rect 3278 7886 3318 7920
rect 3352 7886 3392 7920
rect 3426 7886 3466 7920
rect 3500 7886 3539 7920
rect 3573 7886 3612 7920
rect 3646 7886 3685 7920
rect 3719 7886 3758 7920
rect 3792 7886 3831 7920
rect 3865 7886 3904 7920
rect 3938 7886 3977 7920
rect 4011 7886 4050 7920
rect 4084 7886 4123 7920
rect 4157 7886 4196 7920
rect 4230 7886 4269 7920
rect 4303 7886 4342 7920
rect 4376 7886 4415 7920
rect 4449 7886 4488 7920
rect 4522 7886 4561 7920
rect 4595 7886 4634 7920
rect 4668 7886 4707 7920
rect 4741 7886 4780 7920
rect 4814 7886 4853 7920
rect 4887 7886 4926 7920
rect 4960 7886 4999 7920
rect 5033 7886 5072 7920
rect 5106 7886 5145 7920
rect 5179 7886 5218 7920
rect 5252 7886 5291 7920
rect 5325 7886 5364 7920
rect 5398 7886 5437 7920
rect 5471 7886 5510 7920
rect 5544 7886 5583 7920
rect 5617 7886 5656 7920
rect 5690 7886 5729 7920
rect 5763 7886 5802 7920
rect 5836 7886 5875 7920
rect 5909 7886 5948 7920
rect 5982 7886 6021 7920
rect 6055 7886 6094 7920
rect 6128 7886 6167 7920
rect 6201 7886 6240 7920
rect 6274 7886 6313 7920
rect 6347 7886 6386 7920
rect 6420 7886 6459 7920
rect 6493 7886 6532 7920
rect 6566 7886 6605 7920
rect 6639 7886 6678 7920
rect 6712 7886 6744 7920
rect 2842 7880 6744 7886
rect 7006 7852 7052 7886
rect 7086 7852 7132 7886
rect 7166 7852 7212 7886
rect 7246 7852 7292 7886
rect 7326 7852 7372 7886
rect 7406 7852 7451 7886
rect 7485 7852 7530 7886
rect 7716 7881 7750 7893
rect 7624 7829 7658 7841
rect 7624 7738 7658 7791
rect 7178 7696 7222 7730
rect 7256 7696 7299 7730
rect 7333 7696 7376 7730
rect 7410 7696 7453 7730
rect 7487 7696 7530 7730
rect 7624 7646 7658 7696
rect 7624 7585 7658 7601
rect 7716 7809 7750 7815
rect 7716 7737 7750 7747
rect 7716 7665 7750 7679
rect 7716 7593 7750 7611
rect 7006 7540 7058 7574
rect 7092 7540 7144 7574
rect 7178 7540 7230 7574
rect 7264 7540 7316 7574
rect 7350 7540 7402 7574
rect 7624 7513 7658 7529
rect 7624 7443 7658 7470
rect 7178 7384 7222 7418
rect 7256 7384 7299 7418
rect 7333 7384 7376 7418
rect 7410 7384 7453 7418
rect 7487 7384 7530 7418
rect 7624 7373 7658 7397
rect 7624 7303 7658 7324
rect 7006 7228 7058 7262
rect 7092 7228 7144 7262
rect 7178 7228 7230 7262
rect 7264 7228 7316 7262
rect 7350 7228 7402 7262
rect 7624 7233 7658 7251
rect 7624 7163 7658 7177
rect 7178 7072 7222 7106
rect 7256 7072 7299 7106
rect 7333 7072 7376 7106
rect 7410 7072 7453 7106
rect 7487 7072 7530 7106
rect 7624 7093 7658 7103
rect 7624 7023 7658 7029
rect 7624 6953 7658 6955
rect 7006 6916 7058 6950
rect 7092 6916 7144 6950
rect 7178 6916 7230 6950
rect 7264 6916 7316 6950
rect 7350 6916 7402 6950
rect 7624 6915 7658 6919
rect 7624 6841 7658 6849
rect 7178 6760 7222 6794
rect 7256 6760 7299 6794
rect 7333 6760 7376 6794
rect 7410 6760 7453 6794
rect 7487 6760 7530 6794
rect 7624 6767 7658 6779
rect 7624 6693 7658 6708
rect 7006 6604 7058 6638
rect 7092 6604 7144 6638
rect 7178 6604 7230 6638
rect 7264 6604 7316 6638
rect 7350 6604 7402 6638
rect 7624 6619 7658 6637
rect 7624 6545 7658 6566
rect 7178 6448 7222 6482
rect 7256 6448 7299 6482
rect 7333 6448 7376 6482
rect 7410 6448 7453 6482
rect 7487 6448 7530 6482
rect 7624 6471 7658 6495
rect 7624 6397 7658 6424
rect 7624 6337 7658 6353
rect 7716 7521 7750 7543
rect 7716 7449 7750 7475
rect 7716 7377 7750 7407
rect 7716 7305 7750 7339
rect 7716 7237 7750 7271
rect 7716 7169 7750 7199
rect 7716 7101 7750 7127
rect 7716 7033 7750 7055
rect 7716 6965 7750 6983
rect 7716 6897 7750 6911
rect 7716 6829 7750 6839
rect 7716 6761 7750 6767
rect 7716 6693 7750 6695
rect 7716 6657 7750 6659
rect 7716 6585 7750 6591
rect 7716 6513 7750 6523
rect 7716 6441 7750 6455
rect 7716 6369 7750 6387
rect 7006 6292 7058 6326
rect 7092 6292 7144 6326
rect 7178 6292 7230 6326
rect 7264 6292 7316 6326
rect 7350 6292 7402 6326
rect 7716 6297 7750 6319
rect 7624 6267 7658 6281
rect 7624 6196 7658 6231
rect 7178 6136 7222 6170
rect 7256 6136 7299 6170
rect 7333 6136 7376 6170
rect 7410 6136 7453 6170
rect 7487 6136 7530 6170
rect 7624 6146 7658 6161
rect 7716 6225 7750 6251
rect 7716 6153 7750 6183
rect 7716 6081 7750 6115
rect 7006 6026 7052 6060
rect 7086 6026 7132 6060
rect 7166 6026 7212 6060
rect 7246 6026 7292 6060
rect 7326 6026 7372 6060
rect 7406 6026 7451 6060
rect 7485 6026 7530 6060
rect 7624 6003 7658 6015
rect 7624 5916 7658 5965
rect 7178 5870 7222 5904
rect 7256 5870 7299 5904
rect 7333 5870 7376 5904
rect 7410 5870 7453 5904
rect 7487 5870 7530 5904
rect 7624 5828 7658 5870
rect 7624 5759 7658 5775
rect 7716 6013 7750 6047
rect 7716 5945 7750 5975
rect 7716 5877 7750 5903
rect 7716 5809 7750 5831
rect 7006 5714 7058 5748
rect 7092 5714 7144 5748
rect 7178 5714 7230 5748
rect 7264 5714 7316 5748
rect 7350 5714 7402 5748
rect 7716 5741 7750 5759
rect 7624 5687 7658 5703
rect 7624 5617 7658 5636
rect 7178 5558 7222 5592
rect 7256 5558 7299 5592
rect 7333 5558 7376 5592
rect 7410 5558 7453 5592
rect 7487 5558 7530 5592
rect 7624 5547 7658 5563
rect 7624 5477 7658 5490
rect 7006 5402 7058 5436
rect 7092 5402 7144 5436
rect 7178 5402 7230 5436
rect 7264 5402 7316 5436
rect 7350 5402 7402 5436
rect 7624 5407 7658 5417
rect 7624 5337 7658 5344
rect 7178 5246 7222 5280
rect 7256 5246 7299 5280
rect 7333 5246 7376 5280
rect 7410 5246 7453 5280
rect 7487 5246 7530 5280
rect 7624 5267 7658 5271
rect 7624 5232 7658 5233
rect 7624 5197 7658 5198
rect 7624 5159 7658 5163
rect 7006 5090 7058 5124
rect 7092 5090 7144 5124
rect 7178 5090 7230 5124
rect 7264 5090 7316 5124
rect 7350 5090 7402 5124
rect 7624 5086 7658 5093
rect 7624 5013 7658 5023
rect 7178 4934 7222 4968
rect 7256 4934 7299 4968
rect 7333 4934 7376 4968
rect 7410 4934 7453 4968
rect 7487 4934 7530 4968
rect 7624 4940 7658 4953
rect 7624 4867 7658 4882
rect 7006 4778 7058 4812
rect 7092 4778 7144 4812
rect 7178 4778 7230 4812
rect 7264 4778 7316 4812
rect 7350 4778 7402 4812
rect 7624 4793 7658 4811
rect 7624 4719 7658 4740
rect 7178 4622 7222 4656
rect 7256 4622 7299 4656
rect 7333 4622 7376 4656
rect 7410 4622 7453 4656
rect 7487 4622 7530 4656
rect 7624 4645 7658 4669
rect 7624 4571 7658 4598
rect 7624 4511 7658 4527
rect 7716 5673 7750 5687
rect 7716 5605 7750 5615
rect 7716 5537 7750 5543
rect 7716 5469 7750 5471
rect 7716 5432 7750 5435
rect 7716 5359 7750 5367
rect 7716 5286 7750 5299
rect 7716 5213 7750 5231
rect 7716 5140 7750 5163
rect 7716 5067 7750 5095
rect 7716 4994 7750 5027
rect 7716 4925 7750 4959
rect 7716 4857 7750 4887
rect 7716 4789 7750 4814
rect 7716 4721 7750 4741
rect 7716 4653 7750 4668
rect 7716 4585 7750 4595
rect 7716 4517 7750 4522
rect 7006 4466 7058 4500
rect 7092 4466 7144 4500
rect 7178 4466 7230 4500
rect 7264 4466 7316 4500
rect 7350 4466 7402 4500
rect 7624 4439 7658 4455
rect 7624 4370 7658 4405
rect 7178 4310 7222 4344
rect 7256 4310 7299 4344
rect 7333 4310 7376 4344
rect 7410 4310 7453 4344
rect 7487 4310 7530 4344
rect 7624 4320 7658 4333
rect 7716 4410 7750 4415
rect 7716 4337 7750 4347
rect 7716 4264 7750 4279
rect 7006 4200 7052 4234
rect 7086 4200 7132 4234
rect 7166 4200 7212 4234
rect 7246 4200 7292 4234
rect 7326 4200 7372 4234
rect 7406 4200 7451 4234
rect 7485 4200 7530 4234
rect 7716 4191 7750 4211
rect 7624 4177 7658 4189
rect 7624 4099 7658 4139
rect 7178 4044 7222 4078
rect 7256 4044 7299 4078
rect 7333 4044 7376 4078
rect 7410 4044 7453 4078
rect 7487 4044 7530 4078
rect 7624 4020 7658 4044
rect 7624 3983 7658 3986
rect 7624 3933 7658 3949
rect 7716 4118 7750 4143
rect 7716 4045 7750 4075
rect 7716 3973 7750 4007
rect 7006 3888 7058 3922
rect 7092 3888 7144 3922
rect 7178 3888 7230 3922
rect 7264 3888 7316 3922
rect 7350 3888 7402 3922
rect 7716 3905 7750 3938
rect 7624 3861 7658 3877
rect 7624 3791 7658 3816
rect 7178 3732 7222 3766
rect 7256 3732 7299 3766
rect 7333 3732 7376 3766
rect 7410 3732 7453 3766
rect 7487 3732 7530 3766
rect 7624 3721 7658 3741
rect 7624 3651 7658 3666
rect 4363 3557 4368 3591
rect 4413 3557 4440 3591
rect 4481 3557 4497 3591
rect 4553 3557 4569 3591
rect 4603 3557 4607 3591
rect 4675 3557 4682 3591
rect 4747 3557 4757 3591
rect 4819 3557 4832 3591
rect 4891 3557 4907 3591
rect 4963 3557 4982 3591
rect 5034 3557 5057 3591
rect 5105 3557 5121 3591
rect 5177 3557 5193 3591
rect 5227 3557 5228 3591
rect 5262 3557 5265 3591
rect 5299 3557 5320 3591
rect 5371 3557 5409 3591
rect 5446 3557 5481 3591
rect 5537 3557 5553 3591
rect 5587 3557 5624 3591
rect 5658 3557 5695 3591
rect 5729 3557 5745 3591
rect 7006 3576 7058 3610
rect 7092 3576 7144 3610
rect 7178 3576 7230 3610
rect 7264 3576 7316 3610
rect 7350 3576 7402 3610
rect 7624 3581 7658 3591
rect 7624 3511 7658 3516
rect 7624 3475 7658 3477
rect 7178 3420 7222 3454
rect 7256 3420 7299 3454
rect 7333 3420 7376 3454
rect 7410 3420 7453 3454
rect 7487 3420 7530 3454
rect 7624 3399 7658 3407
rect 7624 3323 7658 3337
rect 7006 3264 7058 3298
rect 7092 3264 7144 3298
rect 7178 3264 7230 3298
rect 7264 3264 7316 3298
rect 7350 3264 7402 3298
rect 7624 3247 7658 3267
rect 7624 3171 7658 3197
rect 7178 3108 7222 3142
rect 7256 3108 7299 3142
rect 7333 3108 7376 3142
rect 7410 3108 7453 3142
rect 7487 3108 7530 3142
rect 7624 3095 7658 3127
rect 7624 3019 7658 3056
rect 7006 2952 7058 2986
rect 7092 2952 7144 2986
rect 7178 2952 7230 2986
rect 7264 2952 7316 2986
rect 7350 2952 7402 2986
rect 7624 2948 7658 2985
rect 7624 2877 7658 2909
rect 7178 2796 7227 2830
rect 7261 2796 7310 2830
rect 7344 2796 7392 2830
rect 7426 2796 7474 2830
rect 7624 2806 7658 2833
rect 7624 2735 7658 2757
rect 7624 2685 7658 2701
rect 7716 3837 7750 3865
rect 7716 3769 7750 3792
rect 7716 3701 7750 3719
rect 7716 3633 7750 3646
rect 7716 3565 7750 3573
rect 7716 3497 7750 3500
rect 7716 3461 7750 3463
rect 7716 3388 7750 3395
rect 7716 3315 7750 3327
rect 7716 3242 7750 3259
rect 7716 3169 7750 3191
rect 7716 3096 7750 3123
rect 7716 3023 7750 3055
rect 7716 2953 7750 2987
rect 7716 2885 7750 2916
rect 7716 2817 7750 2843
rect 7716 2749 7750 2770
rect 7716 2681 7750 2715
rect 7006 2640 7058 2674
rect 7092 2640 7144 2674
rect 7178 2640 7230 2674
rect 7264 2640 7316 2674
rect 7350 2640 7402 2674
rect 7624 2617 7658 2629
rect 7624 2613 7625 2617
rect 7658 2579 7659 2583
rect 7624 2545 7659 2579
rect 7658 2523 7659 2545
rect 7178 2484 7222 2518
rect 7256 2484 7299 2518
rect 7333 2484 7376 2518
rect 7410 2484 7453 2518
rect 7487 2484 7530 2518
rect 7624 2495 7625 2511
rect 7716 2613 7750 2647
rect 7716 2545 7750 2579
rect 7716 2477 7750 2511
rect 7044 2310 7926 2316
rect 7044 2309 8002 2310
rect 7044 2276 7076 2309
rect 7110 2276 7155 2309
rect 7189 2276 7234 2309
rect 7268 2276 7313 2309
rect 7347 2276 7392 2309
rect 7426 2276 7470 2309
rect 7504 2276 7548 2309
rect 7582 2276 7626 2309
rect 7660 2276 7704 2309
rect 7738 2276 7782 2309
rect 7816 2276 7860 2309
rect 7894 2276 8002 2309
rect 7044 2242 7071 2276
rect 7110 2275 7139 2276
rect 7189 2275 7207 2276
rect 7268 2275 7275 2276
rect 7105 2242 7139 2275
rect 7173 2242 7207 2275
rect 7241 2242 7275 2275
rect 7309 2275 7313 2276
rect 7377 2275 7392 2276
rect 7445 2275 7470 2276
rect 7309 2242 7343 2275
rect 7377 2242 7411 2275
rect 7445 2242 7479 2275
rect 7513 2242 7547 2276
rect 7582 2275 7615 2276
rect 7660 2275 7683 2276
rect 7738 2275 7751 2276
rect 7816 2275 7819 2276
rect 7581 2242 7615 2275
rect 7649 2242 7683 2275
rect 7717 2242 7751 2275
rect 7785 2242 7819 2275
rect 7853 2275 7860 2276
rect 7853 2242 7887 2275
rect 7921 2242 8002 2276
rect 7044 2231 8002 2242
rect 7044 2207 7076 2231
rect 7110 2207 7155 2231
rect 7189 2207 7234 2231
rect 7268 2207 7313 2231
rect 7347 2207 7392 2231
rect 7426 2207 7470 2231
rect 7504 2207 7548 2231
rect 7582 2207 7626 2231
rect 7660 2207 7704 2231
rect 7738 2207 7782 2231
rect 7816 2207 7860 2231
rect 7894 2207 8002 2231
rect 7044 2173 7071 2207
rect 7110 2197 7139 2207
rect 7189 2197 7207 2207
rect 7268 2197 7275 2207
rect 7105 2173 7139 2197
rect 7173 2173 7207 2197
rect 7241 2173 7275 2197
rect 7309 2197 7313 2207
rect 7377 2197 7392 2207
rect 7445 2197 7470 2207
rect 7309 2173 7343 2197
rect 7377 2173 7411 2197
rect 7445 2173 7479 2197
rect 7513 2173 7547 2207
rect 7582 2197 7615 2207
rect 7660 2197 7683 2207
rect 7738 2197 7751 2207
rect 7816 2197 7819 2207
rect 7581 2173 7615 2197
rect 7649 2173 7683 2197
rect 7717 2173 7751 2197
rect 7785 2173 7819 2197
rect 7853 2197 7860 2207
rect 7853 2173 7887 2197
rect 7921 2173 8002 2207
rect 7044 2153 8002 2173
rect 7044 2138 7076 2153
rect 7110 2138 7155 2153
rect 7189 2138 7234 2153
rect 7268 2138 7313 2153
rect 7347 2138 7392 2153
rect 7426 2138 7470 2153
rect 7504 2138 7548 2153
rect 7582 2138 7626 2153
rect 7660 2138 7704 2153
rect 7738 2138 7782 2153
rect 7816 2138 7860 2153
rect 7894 2138 8002 2153
rect 7044 2104 7071 2138
rect 7110 2119 7139 2138
rect 7189 2119 7207 2138
rect 7268 2119 7275 2138
rect 7105 2104 7139 2119
rect 7173 2104 7207 2119
rect 7241 2104 7275 2119
rect 7309 2119 7313 2138
rect 7377 2119 7392 2138
rect 7445 2119 7470 2138
rect 7309 2104 7343 2119
rect 7377 2104 7411 2119
rect 7445 2104 7479 2119
rect 7513 2104 7547 2138
rect 7582 2119 7615 2138
rect 7660 2119 7683 2138
rect 7738 2119 7751 2138
rect 7816 2119 7819 2138
rect 7581 2104 7615 2119
rect 7649 2104 7683 2119
rect 7717 2104 7751 2119
rect 7785 2104 7819 2119
rect 7853 2119 7860 2138
rect 7853 2104 7887 2119
rect 7921 2104 8002 2138
rect 7044 2075 8002 2104
rect 7044 2068 7076 2075
rect 7110 2068 7155 2075
rect 7189 2068 7234 2075
rect 7268 2068 7313 2075
rect 7347 2068 7392 2075
rect 7426 2068 7470 2075
rect 7504 2068 7548 2075
rect 7582 2068 7626 2075
rect 7660 2068 7704 2075
rect 7738 2068 7782 2075
rect 7816 2068 7860 2075
rect 7894 2068 8002 2075
rect 7044 2034 7071 2068
rect 7110 2041 7139 2068
rect 7189 2041 7207 2068
rect 7268 2041 7275 2068
rect 7105 2034 7139 2041
rect 7173 2034 7207 2041
rect 7241 2034 7275 2041
rect 7309 2041 7313 2068
rect 7377 2041 7392 2068
rect 7445 2041 7470 2068
rect 7309 2034 7343 2041
rect 7377 2034 7411 2041
rect 7445 2034 7479 2041
rect 7513 2034 7547 2068
rect 7582 2041 7615 2068
rect 7660 2041 7683 2068
rect 7738 2041 7751 2068
rect 7816 2041 7819 2068
rect 7581 2034 7615 2041
rect 7649 2034 7683 2041
rect 7717 2034 7751 2041
rect 7785 2034 7819 2041
rect 7853 2041 7860 2068
rect 7853 2034 7887 2041
rect 7921 2034 8002 2068
rect 7044 1998 8002 2034
rect 7044 1964 7071 1998
rect 7105 1997 7139 1998
rect 7173 1997 7207 1998
rect 7241 1997 7275 1998
rect 7110 1964 7139 1997
rect 7189 1964 7207 1997
rect 7268 1964 7275 1997
rect 7309 1997 7343 1998
rect 7377 1997 7411 1998
rect 7445 1997 7479 1998
rect 7309 1964 7313 1997
rect 7377 1964 7392 1997
rect 7445 1964 7470 1997
rect 7513 1964 7547 1998
rect 7581 1997 7615 1998
rect 7649 1997 7683 1998
rect 7717 1997 7751 1998
rect 7785 1997 7819 1998
rect 7582 1964 7615 1997
rect 7660 1964 7683 1997
rect 7738 1964 7751 1997
rect 7816 1964 7819 1997
rect 7853 1997 7887 1998
rect 7853 1964 7860 1997
rect 7921 1964 8002 1998
rect 7044 1963 7076 1964
rect 7110 1963 7155 1964
rect 7189 1963 7234 1964
rect 7268 1963 7313 1964
rect 7347 1963 7392 1964
rect 7426 1963 7470 1964
rect 7504 1963 7548 1964
rect 7582 1963 7626 1964
rect 7660 1963 7704 1964
rect 7738 1963 7782 1964
rect 7816 1963 7860 1964
rect 7894 1963 8002 1964
rect 7044 1928 8002 1963
rect 7044 1894 7071 1928
rect 7105 1919 7139 1928
rect 7173 1919 7207 1928
rect 7241 1919 7275 1928
rect 7110 1894 7139 1919
rect 7189 1894 7207 1919
rect 7268 1894 7275 1919
rect 7309 1919 7343 1928
rect 7377 1919 7411 1928
rect 7445 1919 7479 1928
rect 7309 1894 7313 1919
rect 7377 1894 7392 1919
rect 7445 1894 7470 1919
rect 7513 1894 7547 1928
rect 7581 1919 7615 1928
rect 7649 1919 7683 1928
rect 7717 1919 7751 1928
rect 7785 1919 7819 1928
rect 7582 1894 7615 1919
rect 7660 1894 7683 1919
rect 7738 1894 7751 1919
rect 7816 1894 7819 1919
rect 7853 1919 7887 1928
rect 7853 1894 7860 1919
rect 7921 1894 8002 1928
rect 7044 1885 7076 1894
rect 7110 1885 7155 1894
rect 7189 1885 7234 1894
rect 7268 1885 7313 1894
rect 7347 1885 7392 1894
rect 7426 1885 7470 1894
rect 7504 1885 7548 1894
rect 7582 1885 7626 1894
rect 7660 1885 7704 1894
rect 7738 1885 7782 1894
rect 7816 1885 7860 1894
rect 7894 1885 8002 1894
rect 7044 1858 8002 1885
rect 7044 1824 7071 1858
rect 7105 1841 7139 1858
rect 7173 1841 7207 1858
rect 7241 1841 7275 1858
rect 7110 1824 7139 1841
rect 7189 1824 7207 1841
rect 7268 1824 7275 1841
rect 7309 1841 7343 1858
rect 7377 1841 7411 1858
rect 7445 1841 7479 1858
rect 7309 1824 7313 1841
rect 7377 1824 7392 1841
rect 7445 1824 7470 1841
rect 7513 1824 7547 1858
rect 7581 1841 7615 1858
rect 7649 1841 7683 1858
rect 7717 1841 7751 1858
rect 7785 1841 7819 1858
rect 7582 1824 7615 1841
rect 7660 1824 7683 1841
rect 7738 1824 7751 1841
rect 7816 1824 7819 1841
rect 7853 1841 7887 1858
rect 7853 1824 7860 1841
rect 7921 1824 8002 1858
rect 7044 1807 7076 1824
rect 7110 1807 7155 1824
rect 7189 1807 7234 1824
rect 7268 1807 7313 1824
rect 7347 1807 7392 1824
rect 7426 1807 7470 1824
rect 7504 1807 7548 1824
rect 7582 1807 7626 1824
rect 7660 1807 7704 1824
rect 7738 1807 7782 1824
rect 7816 1807 7860 1824
rect 7894 1807 8002 1824
rect 7044 1800 8002 1807
rect 7071 1788 8002 1800
rect 7105 1754 7139 1788
rect 7173 1754 7207 1788
rect 7241 1754 7275 1788
rect 7309 1754 7343 1788
rect 7377 1754 7411 1788
rect 7445 1754 7479 1788
rect 7513 1754 7547 1788
rect 7581 1754 7615 1788
rect 7649 1754 7683 1788
rect 7717 1754 7751 1788
rect 7785 1754 7819 1788
rect 7853 1754 7887 1788
rect 7921 1754 8002 1788
rect 7071 1718 8002 1754
rect 2843 1622 3506 1688
rect 7105 1684 7139 1718
rect 7173 1684 7207 1718
rect 7241 1684 7275 1718
rect 7309 1684 7343 1718
rect 7377 1684 7411 1718
rect 7445 1684 7479 1718
rect 7513 1684 7547 1718
rect 7581 1684 7615 1718
rect 7649 1684 7683 1718
rect 7717 1684 7751 1718
rect 7785 1684 7819 1718
rect 7853 1684 7887 1718
rect 7921 1684 8002 1718
rect 7071 1648 8002 1684
rect 7105 1614 7139 1648
rect 7173 1614 7207 1648
rect 7241 1614 7275 1648
rect 7309 1614 7343 1648
rect 7377 1614 7411 1648
rect 7445 1614 7479 1648
rect 7513 1614 7547 1648
rect 7581 1614 7615 1648
rect 7649 1614 7683 1648
rect 7717 1614 7751 1648
rect 7785 1614 7819 1648
rect 7853 1614 7887 1648
rect 7921 1614 8002 1648
rect 7071 1578 8002 1614
rect 7105 1545 7139 1578
rect 7173 1545 7207 1578
rect 7241 1545 7275 1578
rect 7309 1545 7343 1578
rect 7377 1545 7411 1578
rect 7044 1511 7049 1545
rect 7105 1544 7121 1545
rect 7173 1544 7193 1545
rect 7241 1544 7265 1545
rect 7309 1544 7337 1545
rect 7377 1544 7409 1545
rect 7445 1544 7479 1578
rect 7513 1545 7547 1578
rect 7581 1545 7615 1578
rect 7649 1545 7683 1578
rect 7717 1545 7751 1578
rect 7785 1545 7819 1578
rect 7853 1545 7887 1578
rect 7515 1544 7547 1545
rect 7587 1544 7615 1545
rect 7659 1544 7683 1545
rect 7731 1544 7751 1545
rect 7803 1544 7819 1545
rect 7875 1544 7887 1545
rect 7921 1544 8002 1578
rect 7083 1511 7121 1544
rect 7155 1511 7193 1544
rect 7227 1511 7265 1544
rect 7299 1511 7337 1544
rect 7371 1511 7409 1544
rect 7443 1511 7481 1544
rect 7515 1511 7553 1544
rect 7587 1511 7625 1544
rect 7659 1511 7697 1544
rect 7731 1511 7769 1544
rect 7803 1511 7841 1544
rect 7875 1511 8002 1544
rect 7044 1508 8002 1511
rect 7044 1474 7071 1508
rect 7105 1474 7139 1508
rect 7173 1474 7207 1508
rect 7241 1474 7275 1508
rect 7309 1474 7343 1508
rect 7377 1474 7411 1508
rect 7445 1474 7479 1508
rect 7513 1474 7547 1508
rect 7581 1474 7615 1508
rect 7649 1474 7683 1508
rect 7717 1474 7751 1508
rect 7785 1474 7819 1508
rect 7853 1474 7887 1508
rect 7921 1474 8002 1508
rect 7044 1472 8002 1474
rect 7044 1438 7049 1472
rect 7083 1438 7121 1472
rect 7155 1438 7193 1472
rect 7227 1438 7265 1472
rect 7299 1438 7337 1472
rect 7371 1438 7409 1472
rect 7443 1438 7481 1472
rect 7515 1438 7553 1472
rect 7587 1438 7625 1472
rect 7659 1438 7697 1472
rect 7731 1438 7769 1472
rect 7803 1438 7841 1472
rect 7875 1438 8002 1472
rect 7044 1404 7071 1438
rect 7105 1404 7139 1438
rect 7173 1404 7207 1438
rect 7241 1404 7275 1438
rect 7309 1404 7343 1438
rect 7377 1404 7411 1438
rect 7445 1404 7479 1438
rect 7513 1404 7547 1438
rect 7581 1404 7615 1438
rect 7649 1404 7683 1438
rect 7717 1404 7751 1438
rect 7785 1404 7819 1438
rect 7853 1404 7887 1438
rect 7921 1404 8002 1438
rect 7044 1399 8002 1404
rect 7044 1365 7049 1399
rect 7083 1368 7121 1399
rect 7155 1368 7193 1399
rect 7227 1368 7265 1399
rect 7299 1368 7337 1399
rect 7371 1368 7409 1399
rect 7443 1368 7481 1399
rect 7515 1368 7553 1399
rect 7587 1368 7625 1399
rect 7659 1368 7697 1399
rect 7731 1368 7769 1399
rect 7803 1368 7841 1399
rect 7875 1368 8002 1399
rect 7105 1365 7121 1368
rect 7173 1365 7193 1368
rect 7241 1365 7265 1368
rect 7309 1365 7337 1368
rect 7377 1365 7409 1368
rect 7044 1334 7071 1365
rect 7105 1334 7139 1365
rect 7173 1334 7207 1365
rect 7241 1334 7275 1365
rect 7309 1334 7343 1365
rect 7377 1334 7411 1365
rect 7445 1334 7479 1368
rect 7515 1365 7547 1368
rect 7587 1365 7615 1368
rect 7659 1365 7683 1368
rect 7731 1365 7751 1368
rect 7803 1365 7819 1368
rect 7875 1365 7887 1368
rect 7513 1334 7547 1365
rect 7581 1334 7615 1365
rect 7649 1334 7683 1365
rect 7717 1334 7751 1365
rect 7785 1334 7819 1365
rect 7853 1334 7887 1365
rect 7921 1334 8002 1368
rect 7044 1326 8002 1334
rect 7044 1292 7049 1326
rect 7083 1298 7121 1326
rect 7155 1298 7193 1326
rect 7227 1298 7265 1326
rect 7299 1298 7337 1326
rect 7371 1298 7409 1326
rect 7443 1298 7481 1326
rect 7515 1298 7553 1326
rect 7587 1298 7625 1326
rect 7659 1298 7697 1326
rect 7731 1298 7769 1326
rect 7803 1298 7841 1326
rect 7875 1298 8002 1326
rect 7105 1292 7121 1298
rect 7173 1292 7193 1298
rect 7241 1292 7265 1298
rect 7309 1292 7337 1298
rect 7377 1292 7409 1298
rect 7044 1264 7071 1292
rect 7105 1264 7139 1292
rect 7173 1264 7207 1292
rect 7241 1264 7275 1292
rect 7309 1264 7343 1292
rect 7377 1264 7411 1292
rect 7445 1264 7479 1298
rect 7515 1292 7547 1298
rect 7587 1292 7615 1298
rect 7659 1292 7683 1298
rect 7731 1292 7751 1298
rect 7803 1292 7819 1298
rect 7875 1292 7887 1298
rect 7513 1264 7547 1292
rect 7581 1264 7615 1292
rect 7649 1264 7683 1292
rect 7717 1264 7751 1292
rect 7785 1264 7819 1292
rect 7853 1264 7887 1292
rect 7921 1264 8002 1298
rect 7044 1253 8002 1264
rect 7044 1219 7049 1253
rect 7083 1228 7121 1253
rect 7155 1228 7193 1253
rect 7227 1228 7265 1253
rect 7299 1228 7337 1253
rect 7371 1228 7409 1253
rect 7443 1228 7481 1253
rect 7515 1228 7553 1253
rect 7587 1228 7625 1253
rect 7659 1228 7697 1253
rect 7731 1228 7769 1253
rect 7803 1228 7841 1253
rect 7875 1228 8002 1253
rect 7105 1219 7121 1228
rect 7173 1219 7193 1228
rect 7241 1219 7265 1228
rect 7309 1219 7337 1228
rect 7377 1219 7409 1228
rect 7044 1194 7071 1219
rect 7105 1194 7139 1219
rect 7173 1194 7207 1219
rect 7241 1194 7275 1219
rect 7309 1194 7343 1219
rect 7377 1194 7411 1219
rect 7445 1194 7479 1228
rect 7515 1219 7547 1228
rect 7587 1219 7615 1228
rect 7659 1219 7683 1228
rect 7731 1219 7751 1228
rect 7803 1219 7819 1228
rect 7875 1219 7887 1228
rect 7513 1194 7547 1219
rect 7581 1194 7615 1219
rect 7649 1194 7683 1219
rect 7717 1194 7751 1219
rect 7785 1194 7819 1219
rect 7853 1194 7887 1219
rect 7921 1194 8002 1228
rect 7044 1180 8002 1194
rect 7044 1146 7049 1180
rect 7083 1158 7121 1180
rect 7155 1158 7193 1180
rect 7227 1158 7265 1180
rect 7299 1158 7337 1180
rect 7371 1158 7409 1180
rect 7443 1158 7481 1180
rect 7515 1158 7553 1180
rect 7587 1158 7625 1180
rect 7659 1158 7697 1180
rect 7731 1158 7769 1180
rect 7803 1158 7841 1180
rect 7875 1158 8002 1180
rect 7105 1146 7121 1158
rect 7173 1146 7193 1158
rect 7241 1146 7265 1158
rect 7309 1146 7337 1158
rect 7377 1146 7409 1158
rect 7044 1124 7071 1146
rect 7105 1124 7139 1146
rect 7173 1124 7207 1146
rect 7241 1124 7275 1146
rect 7309 1124 7343 1146
rect 7377 1124 7411 1146
rect 7445 1124 7479 1158
rect 7515 1146 7547 1158
rect 7587 1146 7615 1158
rect 7659 1146 7683 1158
rect 7731 1146 7751 1158
rect 7803 1146 7819 1158
rect 7875 1146 7887 1158
rect 7513 1124 7547 1146
rect 7581 1124 7615 1146
rect 7649 1124 7683 1146
rect 7717 1124 7751 1146
rect 7785 1124 7819 1146
rect 7853 1124 7887 1146
rect 7921 1124 8002 1158
rect 7044 1107 8002 1124
rect 7044 1073 7049 1107
rect 7083 1088 7121 1107
rect 7155 1088 7193 1107
rect 7227 1088 7265 1107
rect 7299 1088 7337 1107
rect 7371 1088 7409 1107
rect 7443 1088 7481 1107
rect 7515 1088 7553 1107
rect 7587 1088 7625 1107
rect 7659 1088 7697 1107
rect 7731 1088 7769 1107
rect 7803 1088 7841 1107
rect 7875 1088 8002 1107
rect 7105 1073 7121 1088
rect 7173 1073 7193 1088
rect 7241 1073 7265 1088
rect 7309 1073 7337 1088
rect 7377 1073 7409 1088
rect 7044 1054 7071 1073
rect 7105 1054 7139 1073
rect 7173 1054 7207 1073
rect 7241 1054 7275 1073
rect 7309 1054 7343 1073
rect 7377 1054 7411 1073
rect 7445 1054 7479 1088
rect 7515 1073 7547 1088
rect 7587 1073 7615 1088
rect 7659 1073 7683 1088
rect 7731 1073 7751 1088
rect 7803 1073 7819 1088
rect 7875 1073 7887 1088
rect 7513 1054 7547 1073
rect 7581 1054 7615 1073
rect 7649 1054 7683 1073
rect 7717 1054 7751 1073
rect 7785 1054 7819 1073
rect 7853 1054 7887 1073
rect 7921 1054 8002 1088
rect 7044 1034 8002 1054
rect 7044 1000 7049 1034
rect 7083 1018 7121 1034
rect 7155 1018 7193 1034
rect 7227 1018 7265 1034
rect 7299 1018 7337 1034
rect 7371 1018 7409 1034
rect 7443 1018 7481 1034
rect 7515 1018 7553 1034
rect 7587 1018 7625 1034
rect 7659 1018 7697 1034
rect 7731 1018 7769 1034
rect 7803 1018 7841 1034
rect 7875 1018 8002 1034
rect 7105 1000 7121 1018
rect 7173 1000 7193 1018
rect 7241 1000 7265 1018
rect 7309 1000 7337 1018
rect 7377 1000 7409 1018
rect 7044 984 7071 1000
rect 7105 984 7139 1000
rect 7173 984 7207 1000
rect 7241 984 7275 1000
rect 7309 984 7343 1000
rect 7377 984 7411 1000
rect 7445 984 7479 1018
rect 7515 1000 7547 1018
rect 7587 1000 7615 1018
rect 7659 1000 7683 1018
rect 7731 1000 7751 1018
rect 7803 1000 7819 1018
rect 7875 1000 7887 1018
rect 7513 984 7547 1000
rect 7581 984 7615 1000
rect 7649 984 7683 1000
rect 7717 984 7751 1000
rect 7785 984 7819 1000
rect 7853 984 7887 1000
rect 7921 984 8002 1018
rect 7044 961 8002 984
rect 7044 927 7049 961
rect 7083 948 7121 961
rect 7155 948 7193 961
rect 7227 948 7265 961
rect 7299 948 7337 961
rect 7371 948 7409 961
rect 7443 948 7481 961
rect 7515 948 7553 961
rect 7587 948 7625 961
rect 7659 948 7697 961
rect 7731 948 7769 961
rect 7803 948 7841 961
rect 7875 948 8002 961
rect 7105 927 7121 948
rect 7173 927 7193 948
rect 7241 927 7265 948
rect 7309 927 7337 948
rect 7377 927 7409 948
rect 7044 914 7071 927
rect 7105 914 7139 927
rect 7173 914 7207 927
rect 7241 914 7275 927
rect 7309 914 7343 927
rect 7377 914 7411 927
rect 7445 914 7479 948
rect 7515 927 7547 948
rect 7587 927 7615 948
rect 7659 927 7683 948
rect 7731 927 7751 948
rect 7803 927 7819 948
rect 7875 927 7887 948
rect 7513 914 7547 927
rect 7581 914 7615 927
rect 7649 914 7683 927
rect 7717 914 7751 927
rect 7785 914 7819 927
rect 7853 914 7887 927
rect 7921 914 8002 948
rect 7044 888 8002 914
rect 7044 854 7049 888
rect 7083 878 7121 888
rect 7155 878 7193 888
rect 7227 878 7265 888
rect 7299 878 7337 888
rect 7371 878 7409 888
rect 7443 878 7481 888
rect 7515 878 7553 888
rect 7587 878 7625 888
rect 7659 878 7697 888
rect 7731 878 7769 888
rect 7803 878 7841 888
rect 7875 878 8002 888
rect 7105 854 7121 878
rect 7173 854 7193 878
rect 7241 854 7265 878
rect 7309 854 7337 878
rect 7377 854 7409 878
rect 7044 844 7071 854
rect 7105 844 7139 854
rect 7173 844 7207 854
rect 7241 844 7275 854
rect 7309 844 7343 854
rect 7377 844 7411 854
rect 7445 844 7479 878
rect 7515 854 7547 878
rect 7587 854 7615 878
rect 7659 854 7683 878
rect 7731 854 7751 878
rect 7803 854 7819 878
rect 7875 854 7887 878
rect 7513 844 7547 854
rect 7581 844 7615 854
rect 7649 844 7683 854
rect 7717 844 7751 854
rect 7785 844 7819 854
rect 7853 844 7887 854
rect 7921 844 8002 878
rect 7044 814 8002 844
rect 7044 780 7049 814
rect 7083 808 7121 814
rect 7155 808 7193 814
rect 7227 808 7265 814
rect 7299 808 7337 814
rect 7371 808 7409 814
rect 7443 808 7481 814
rect 7515 808 7553 814
rect 7587 808 7625 814
rect 7659 808 7697 814
rect 7731 808 7769 814
rect 7803 808 7841 814
rect 7875 808 8002 814
rect 7105 780 7121 808
rect 7173 780 7193 808
rect 7241 780 7265 808
rect 7309 780 7337 808
rect 7377 780 7409 808
rect 7044 774 7071 780
rect 7105 774 7139 780
rect 7173 774 7207 780
rect 7241 774 7275 780
rect 7309 774 7343 780
rect 7377 774 7411 780
rect 7445 774 7479 808
rect 7515 780 7547 808
rect 7587 780 7615 808
rect 7659 780 7683 808
rect 7731 780 7751 808
rect 7803 780 7819 808
rect 7875 780 7887 808
rect 7513 774 7547 780
rect 7581 774 7615 780
rect 7649 774 7683 780
rect 7717 774 7751 780
rect 7785 774 7819 780
rect 7853 774 7887 780
rect 7921 774 8002 808
rect 7044 740 8002 774
rect 7044 706 7049 740
rect 7083 738 7121 740
rect 7155 738 7193 740
rect 7227 738 7265 740
rect 7299 738 7337 740
rect 7371 738 7409 740
rect 7443 738 7481 740
rect 7515 738 7553 740
rect 7587 738 7625 740
rect 7659 738 7697 740
rect 7731 738 7769 740
rect 7803 738 7841 740
rect 7875 738 8002 740
rect 7105 706 7121 738
rect 7173 706 7193 738
rect 7241 706 7265 738
rect 7309 706 7337 738
rect 7377 706 7409 738
rect 7044 704 7071 706
rect 7105 704 7139 706
rect 7173 704 7207 706
rect 7241 704 7275 706
rect 7309 704 7343 706
rect 7377 704 7411 706
rect 7445 704 7479 738
rect 7515 706 7547 738
rect 7587 706 7615 738
rect 7659 706 7683 738
rect 7731 706 7751 738
rect 7803 706 7819 738
rect 7875 706 7887 738
rect 7513 704 7547 706
rect 7581 704 7615 706
rect 7649 704 7683 706
rect 7717 704 7751 706
rect 7785 704 7819 706
rect 7853 704 7887 706
rect 7921 704 8002 738
rect 7044 668 8002 704
rect 7044 666 7071 668
rect 7105 666 7139 668
rect 7173 666 7207 668
rect 7241 666 7275 668
rect 7309 666 7343 668
rect 7377 666 7411 668
rect 7044 632 7049 666
rect 7105 634 7121 666
rect 7173 634 7193 666
rect 7241 634 7265 666
rect 7309 634 7337 666
rect 7377 634 7409 666
rect 7445 634 7479 668
rect 7513 666 7547 668
rect 7581 666 7615 668
rect 7649 666 7683 668
rect 7717 666 7751 668
rect 7785 666 7819 668
rect 7853 666 7887 668
rect 7515 634 7547 666
rect 7587 634 7615 666
rect 7659 634 7683 666
rect 7731 634 7751 666
rect 7803 634 7819 666
rect 7875 634 7887 666
rect 7921 634 8002 668
rect 7083 632 7121 634
rect 7155 632 7193 634
rect 7227 632 7265 634
rect 7299 632 7337 634
rect 7371 632 7409 634
rect 7443 632 7481 634
rect 7515 632 7553 634
rect 7587 632 7625 634
rect 7659 632 7697 634
rect 7731 632 7769 634
rect 7803 632 7841 634
rect 7875 632 8002 634
rect 7044 598 8002 632
rect 7044 592 7071 598
rect 7105 592 7139 598
rect 7173 592 7207 598
rect 7241 592 7275 598
rect 7309 592 7343 598
rect 7377 592 7411 598
rect 7044 558 7049 592
rect 7105 564 7121 592
rect 7173 564 7193 592
rect 7241 564 7265 592
rect 7309 564 7337 592
rect 7377 564 7409 592
rect 7445 564 7479 598
rect 7513 592 7547 598
rect 7581 592 7615 598
rect 7649 592 7683 598
rect 7717 592 7751 598
rect 7785 592 7819 598
rect 7853 592 7887 598
rect 7515 564 7547 592
rect 7587 564 7615 592
rect 7659 564 7683 592
rect 7731 564 7751 592
rect 7803 564 7819 592
rect 7875 564 7887 592
rect 7921 564 8002 598
rect 7083 558 7121 564
rect 7155 558 7193 564
rect 7227 558 7265 564
rect 7299 558 7337 564
rect 7371 558 7409 564
rect 7443 558 7481 564
rect 7515 558 7553 564
rect 7587 558 7625 564
rect 7659 558 7697 564
rect 7731 558 7769 564
rect 7803 558 7841 564
rect 7875 558 8002 564
rect 7044 528 8002 558
rect 7044 518 7071 528
rect 7105 518 7139 528
rect 7173 518 7207 528
rect 7241 518 7275 528
rect 7309 518 7343 528
rect 7377 518 7411 528
rect 7044 484 7049 518
rect 7105 494 7121 518
rect 7173 494 7193 518
rect 7241 494 7265 518
rect 7309 494 7337 518
rect 7377 494 7409 518
rect 7445 494 7479 528
rect 7513 518 7547 528
rect 7581 518 7615 528
rect 7649 518 7683 528
rect 7717 518 7751 528
rect 7785 518 7819 528
rect 7853 518 7887 528
rect 7515 494 7547 518
rect 7587 494 7615 518
rect 7659 494 7683 518
rect 7731 494 7751 518
rect 7803 494 7819 518
rect 7875 494 7887 518
rect 7921 494 8002 528
rect 7083 484 7121 494
rect 7155 484 7193 494
rect 7227 484 7265 494
rect 7299 484 7337 494
rect 7371 484 7409 494
rect 7443 484 7481 494
rect 7515 484 7553 494
rect 7587 484 7625 494
rect 7659 484 7697 494
rect 7731 484 7769 494
rect 7803 484 7841 494
rect 7875 484 8002 494
rect 7044 458 8002 484
rect 7044 444 7071 458
rect 7105 444 7139 458
rect 7173 444 7207 458
rect 7241 444 7275 458
rect 7309 444 7343 458
rect 7377 444 7411 458
rect 7044 410 7049 444
rect 7105 424 7121 444
rect 7173 424 7193 444
rect 7241 424 7265 444
rect 7309 424 7337 444
rect 7377 424 7409 444
rect 7445 424 7479 458
rect 7513 444 7547 458
rect 7581 444 7615 458
rect 7649 444 7683 458
rect 7717 444 7751 458
rect 7785 444 7819 458
rect 7853 444 7887 458
rect 7515 424 7547 444
rect 7587 424 7615 444
rect 7659 424 7683 444
rect 7731 424 7751 444
rect 7803 424 7819 444
rect 7875 424 7887 444
rect 7921 424 8002 458
rect 7083 410 7121 424
rect 7155 410 7193 424
rect 7227 410 7265 424
rect 7299 410 7337 424
rect 7371 410 7409 424
rect 7443 410 7481 424
rect 7515 410 7553 424
rect 7587 410 7625 424
rect 7659 410 7697 424
rect 7731 410 7769 424
rect 7803 410 7841 424
rect 7875 410 8002 424
rect 7044 388 8002 410
rect 7044 370 7071 388
rect 7105 370 7139 388
rect 7173 370 7207 388
rect 7241 370 7275 388
rect 7309 370 7343 388
rect 7377 370 7411 388
rect 7044 336 7049 370
rect 7105 354 7121 370
rect 7173 354 7193 370
rect 7241 354 7265 370
rect 7309 354 7337 370
rect 7377 354 7409 370
rect 7445 354 7479 388
rect 7513 370 7547 388
rect 7581 370 7615 388
rect 7649 370 7683 388
rect 7717 370 7751 388
rect 7785 370 7819 388
rect 7853 370 7887 388
rect 7515 354 7547 370
rect 7587 354 7615 370
rect 7659 354 7683 370
rect 7731 354 7751 370
rect 7803 354 7819 370
rect 7875 354 7887 370
rect 7921 354 8002 388
rect 7083 336 7121 354
rect 7155 336 7193 354
rect 7227 336 7265 354
rect 7299 336 7337 354
rect 7371 336 7409 354
rect 7443 336 7481 354
rect 7515 336 7553 354
rect 7587 336 7625 354
rect 7659 336 7697 354
rect 7731 336 7769 354
rect 7803 336 7841 354
rect 7875 336 8002 354
rect 7044 318 8002 336
rect 7044 296 7071 318
rect 7105 296 7139 318
rect 7173 296 7207 318
rect 7241 296 7275 318
rect 7309 296 7343 318
rect 7377 296 7411 318
rect 7044 262 7049 296
rect 7105 284 7121 296
rect 7173 284 7193 296
rect 7241 284 7265 296
rect 7309 284 7337 296
rect 7377 284 7409 296
rect 7445 284 7479 318
rect 7513 296 7547 318
rect 7581 296 7615 318
rect 7649 296 7683 318
rect 7717 296 7751 318
rect 7785 296 7819 318
rect 7853 296 7887 318
rect 7515 284 7547 296
rect 7587 284 7615 296
rect 7659 284 7683 296
rect 7731 284 7751 296
rect 7803 284 7819 296
rect 7875 284 7887 296
rect 7921 284 8002 318
rect 7083 262 7121 284
rect 7155 262 7193 284
rect 7227 262 7265 284
rect 7299 262 7337 284
rect 7371 262 7409 284
rect 7443 262 7481 284
rect 7515 262 7553 284
rect 7587 262 7625 284
rect 7659 262 7697 284
rect 7731 262 7769 284
rect 7803 262 7841 284
rect 7875 262 8002 284
rect 7044 248 8002 262
rect 7044 222 7071 248
rect 7105 222 7139 248
rect 7173 222 7207 248
rect 7241 222 7275 248
rect 7309 222 7343 248
rect 7377 222 7411 248
rect 7044 188 7049 222
rect 7105 214 7121 222
rect 7173 214 7193 222
rect 7241 214 7265 222
rect 7309 214 7337 222
rect 7377 214 7409 222
rect 7445 214 7479 248
rect 7513 222 7547 248
rect 7581 222 7615 248
rect 7649 222 7683 248
rect 7717 222 7751 248
rect 7785 222 7819 248
rect 7853 222 7887 248
rect 7515 214 7547 222
rect 7587 214 7615 222
rect 7659 214 7683 222
rect 7731 214 7751 222
rect 7803 214 7819 222
rect 7875 214 7887 222
rect 7921 214 8002 248
rect 7083 188 7121 214
rect 7155 188 7193 214
rect 7227 188 7265 214
rect 7299 188 7337 214
rect 7371 188 7409 214
rect 7443 188 7481 214
rect 7515 188 7553 214
rect 7587 188 7625 214
rect 7659 188 7697 214
rect 7731 188 7769 214
rect 7803 188 7841 214
rect 7875 188 8002 214
rect 7044 178 8002 188
rect 7044 148 7071 178
rect 7105 148 7139 178
rect 7173 148 7207 178
rect 7241 148 7275 178
rect 7309 148 7343 178
rect 7377 148 7411 178
rect 7044 114 7049 148
rect 7105 144 7121 148
rect 7173 144 7193 148
rect 7241 144 7265 148
rect 7309 144 7337 148
rect 7377 144 7409 148
rect 7445 144 7479 178
rect 7513 148 7547 178
rect 7581 148 7615 178
rect 7649 148 7683 178
rect 7717 148 7751 178
rect 7785 148 7819 178
rect 7853 148 7887 178
rect 7515 144 7547 148
rect 7587 144 7615 148
rect 7659 144 7683 148
rect 7731 144 7751 148
rect 7803 144 7819 148
rect 7875 144 7887 148
rect 7921 144 8002 178
rect 7083 114 7121 144
rect 7155 114 7193 144
rect 7227 114 7265 144
rect 7299 114 7337 144
rect 7371 114 7409 144
rect 7443 114 7481 144
rect 7515 114 7553 144
rect 7587 114 7625 144
rect 7659 114 7697 144
rect 7731 114 7769 144
rect 7803 114 7841 144
rect 7875 114 8002 144
rect 7044 108 8002 114
rect 7044 74 7071 108
rect 7105 74 7139 108
rect 7173 74 7207 108
rect 7241 74 7275 108
rect 7309 74 7343 108
rect 7377 74 7411 108
rect 7445 74 7479 108
rect 7513 74 7547 108
rect 7581 74 7615 108
rect 7649 74 7683 108
rect 7717 74 7751 108
rect 7785 74 7819 108
rect 7853 74 7887 108
rect 7921 74 8002 108
rect 7044 40 7049 74
rect 7083 40 7121 74
rect 7155 40 7193 74
rect 7227 40 7265 74
rect 7299 40 7337 74
rect 7371 40 7409 74
rect 7443 40 7481 74
rect 7515 40 7553 74
rect 7587 40 7625 74
rect 7659 40 7697 74
rect 7731 40 7769 74
rect 7803 40 7841 74
rect 7875 40 8002 74
<< viali >>
rect 2884 27873 2900 27903
rect 2900 27873 2918 27903
rect 2957 27873 2969 27903
rect 2969 27873 2991 27903
rect 2884 27869 2918 27873
rect 2957 27869 2991 27873
rect 3030 27869 3038 27903
rect 3038 27869 3064 27903
rect 3103 27869 3137 27903
rect 3176 27869 3210 27903
rect 3249 27869 3283 27903
rect 3322 27869 3356 27903
rect 3395 27869 3429 27903
rect 3468 27869 3502 27903
rect 3541 27869 3575 27903
rect 3614 27869 3648 27903
rect 3687 27869 3721 27903
rect 3760 27869 3794 27903
rect 3833 27869 3867 27903
rect 3906 27869 3940 27903
rect 3979 27869 4013 27903
rect 4052 27869 4086 27903
rect 4125 27869 4159 27903
rect 4198 27869 4232 27903
rect 4271 27869 4305 27903
rect 4344 27869 4378 27903
rect 4417 27869 4451 27903
rect 4490 27869 4524 27903
rect 4563 27869 4597 27903
rect 4636 27869 4670 27903
rect 4709 27869 4743 27903
rect 4782 27869 4816 27903
rect 4855 27869 4889 27903
rect 4928 27869 4962 27903
rect 5001 27869 5035 27903
rect 5074 27869 5108 27903
rect 5147 27869 5181 27903
rect 5220 27869 5254 27903
rect 5293 27869 5327 27903
rect 5366 27869 5400 27903
rect 5439 27869 5473 27903
rect 5512 27869 5546 27903
rect 5585 27869 5619 27903
rect 5658 27869 5692 27903
rect 5731 27869 5765 27903
rect 5804 27869 5838 27903
rect 5877 27869 5911 27903
rect 5950 27869 5984 27903
rect 6023 27869 6057 27903
rect 2884 27805 2900 27823
rect 2900 27805 2918 27823
rect 2957 27805 2969 27823
rect 2969 27805 2991 27823
rect 2884 27789 2918 27805
rect 2957 27789 2991 27805
rect 3030 27789 3038 27823
rect 3038 27789 3064 27823
rect 3103 27789 3137 27823
rect 3176 27789 3210 27823
rect 3249 27789 3283 27823
rect 3322 27789 3356 27823
rect 3395 27789 3429 27823
rect 3468 27789 3502 27823
rect 3541 27789 3575 27823
rect 3614 27789 3648 27823
rect 3687 27789 3721 27823
rect 3760 27789 3794 27823
rect 3833 27789 3867 27823
rect 3906 27789 3940 27823
rect 3979 27789 4013 27823
rect 4052 27789 4086 27823
rect 4125 27789 4159 27823
rect 4198 27789 4232 27823
rect 4271 27789 4305 27823
rect 4344 27789 4378 27823
rect 4417 27789 4451 27823
rect 4490 27789 4524 27823
rect 4563 27789 4597 27823
rect 4636 27789 4670 27823
rect 4709 27789 4743 27823
rect 4782 27789 4816 27823
rect 4855 27789 4889 27823
rect 4928 27789 4962 27823
rect 5001 27789 5035 27823
rect 5074 27789 5108 27823
rect 5147 27789 5181 27823
rect 5220 27789 5254 27823
rect 5293 27789 5327 27823
rect 5366 27789 5400 27823
rect 5439 27789 5473 27823
rect 5512 27789 5546 27823
rect 5585 27789 5619 27823
rect 5658 27789 5692 27823
rect 5731 27789 5765 27823
rect 5804 27789 5838 27823
rect 5877 27789 5911 27823
rect 5950 27789 5984 27823
rect 6023 27789 6057 27823
rect 2884 27737 2900 27743
rect 2900 27737 2918 27743
rect 2957 27737 2969 27743
rect 2969 27737 2991 27743
rect 2884 27709 2918 27737
rect 2957 27709 2991 27737
rect 3030 27709 3038 27743
rect 3038 27709 3064 27743
rect 3103 27709 3137 27743
rect 3176 27709 3210 27743
rect 3249 27709 3283 27743
rect 3322 27709 3356 27743
rect 3395 27709 3429 27743
rect 3468 27709 3502 27743
rect 3541 27709 3575 27743
rect 3614 27709 3648 27743
rect 3687 27709 3721 27743
rect 3760 27709 3794 27743
rect 3833 27709 3867 27743
rect 3906 27709 3940 27743
rect 3979 27709 4013 27743
rect 4052 27709 4086 27743
rect 4125 27709 4159 27743
rect 4198 27709 4232 27743
rect 4271 27709 4305 27743
rect 4344 27709 4378 27743
rect 4417 27709 4451 27743
rect 4490 27709 4524 27743
rect 4563 27709 4597 27743
rect 4636 27709 4670 27743
rect 4709 27709 4743 27743
rect 4782 27709 4816 27743
rect 4855 27709 4889 27743
rect 4928 27709 4962 27743
rect 5001 27709 5035 27743
rect 5074 27709 5108 27743
rect 5147 27709 5181 27743
rect 5220 27709 5254 27743
rect 5293 27709 5327 27743
rect 5366 27709 5400 27743
rect 5439 27709 5473 27743
rect 5512 27709 5546 27743
rect 5585 27709 5619 27743
rect 5658 27709 5692 27743
rect 5731 27709 5765 27743
rect 5804 27709 5838 27743
rect 5877 27709 5911 27743
rect 5950 27709 5984 27743
rect 6023 27709 6057 27743
rect 2884 27635 2918 27663
rect 2957 27635 2991 27663
rect 2884 27629 2900 27635
rect 2900 27629 2918 27635
rect 2957 27629 2969 27635
rect 2969 27629 2991 27635
rect 3030 27629 3038 27663
rect 3038 27629 3064 27663
rect 3103 27629 3137 27663
rect 3176 27629 3210 27663
rect 3249 27629 3283 27663
rect 3322 27629 3356 27663
rect 3395 27629 3429 27663
rect 3468 27629 3502 27663
rect 3541 27629 3575 27663
rect 3614 27629 3648 27663
rect 3687 27629 3721 27663
rect 3760 27629 3794 27663
rect 3833 27629 3867 27663
rect 3906 27629 3940 27663
rect 3979 27629 4013 27663
rect 4052 27629 4086 27663
rect 4125 27629 4159 27663
rect 4198 27629 4232 27663
rect 4271 27629 4305 27663
rect 4344 27629 4378 27663
rect 4417 27629 4451 27663
rect 4490 27629 4524 27663
rect 4563 27629 4597 27663
rect 4636 27629 4670 27663
rect 4709 27629 4743 27663
rect 4782 27629 4816 27663
rect 4855 27629 4889 27663
rect 4928 27629 4962 27663
rect 5001 27629 5035 27663
rect 5074 27629 5108 27663
rect 5147 27629 5181 27663
rect 5220 27629 5254 27663
rect 5293 27629 5327 27663
rect 5366 27629 5400 27663
rect 5439 27629 5473 27663
rect 5512 27629 5546 27663
rect 5585 27629 5619 27663
rect 5658 27629 5692 27663
rect 5731 27629 5765 27663
rect 5804 27629 5838 27663
rect 5877 27629 5911 27663
rect 5950 27629 5984 27663
rect 6023 27629 6057 27663
rect 2884 27567 2918 27583
rect 2957 27567 2991 27583
rect 2884 27549 2900 27567
rect 2900 27549 2918 27567
rect 2957 27549 2969 27567
rect 2969 27549 2991 27567
rect 3030 27549 3038 27583
rect 3038 27549 3064 27583
rect 3103 27549 3137 27583
rect 3176 27549 3210 27583
rect 3249 27549 3283 27583
rect 3322 27549 3356 27583
rect 3395 27549 3429 27583
rect 3468 27549 3502 27583
rect 3541 27549 3575 27583
rect 3614 27549 3648 27583
rect 3687 27549 3721 27583
rect 3760 27549 3794 27583
rect 3833 27549 3867 27583
rect 3906 27549 3940 27583
rect 3979 27549 4013 27583
rect 4052 27549 4086 27583
rect 4125 27549 4159 27583
rect 4198 27549 4232 27583
rect 4271 27549 4305 27583
rect 4344 27549 4378 27583
rect 4417 27549 4451 27583
rect 4490 27549 4524 27583
rect 4563 27549 4597 27583
rect 4636 27549 4670 27583
rect 4709 27549 4743 27583
rect 4782 27549 4816 27583
rect 4855 27549 4889 27583
rect 4928 27549 4962 27583
rect 5001 27549 5035 27583
rect 5074 27549 5108 27583
rect 5147 27549 5181 27583
rect 5220 27549 5254 27583
rect 5293 27549 5327 27583
rect 5366 27549 5400 27583
rect 5439 27549 5473 27583
rect 5512 27549 5546 27583
rect 5585 27549 5619 27583
rect 5658 27549 5692 27583
rect 5731 27549 5765 27583
rect 5804 27549 5838 27583
rect 5877 27549 5911 27583
rect 5950 27549 5984 27583
rect 6023 27549 6057 27583
rect 2884 27499 2918 27503
rect 2957 27499 2991 27503
rect 2884 27469 2900 27499
rect 2900 27469 2918 27499
rect 2957 27469 2969 27499
rect 2969 27469 2991 27499
rect 3030 27469 3038 27503
rect 3038 27469 3064 27503
rect 3103 27469 3137 27503
rect 3176 27469 3210 27503
rect 3249 27469 3283 27503
rect 3322 27469 3356 27503
rect 3395 27469 3429 27503
rect 3468 27469 3502 27503
rect 3541 27469 3575 27503
rect 3614 27469 3648 27503
rect 3687 27469 3721 27503
rect 3760 27469 3794 27503
rect 3833 27469 3867 27503
rect 3906 27469 3940 27503
rect 3979 27469 4013 27503
rect 4052 27469 4086 27503
rect 4125 27469 4159 27503
rect 4198 27469 4232 27503
rect 4271 27469 4305 27503
rect 4344 27469 4378 27503
rect 4417 27469 4451 27503
rect 4490 27469 4524 27503
rect 4563 27469 4597 27503
rect 4636 27469 4670 27503
rect 4709 27469 4743 27503
rect 4782 27469 4816 27503
rect 4855 27469 4889 27503
rect 4928 27469 4962 27503
rect 5001 27469 5035 27503
rect 5074 27469 5108 27503
rect 5147 27469 5181 27503
rect 5220 27469 5254 27503
rect 5293 27469 5327 27503
rect 5366 27469 5400 27503
rect 5439 27469 5473 27503
rect 5512 27469 5546 27503
rect 5585 27469 5619 27503
rect 5658 27469 5692 27503
rect 5731 27469 5765 27503
rect 5804 27469 5838 27503
rect 5877 27469 5911 27503
rect 5950 27469 5984 27503
rect 6023 27469 6057 27503
rect 3316 27296 3422 27330
rect 3316 27262 3318 27296
rect 3318 27262 3422 27296
rect 3316 27224 3422 27262
rect 5395 27296 5501 27329
rect 5395 27262 5494 27296
rect 5494 27262 5501 27296
rect 5395 27223 5501 27262
rect 7080 26888 7114 26922
rect 7152 26888 7186 26922
rect 7080 26837 7083 26849
rect 7083 26837 7114 26849
rect 7152 26837 7185 26849
rect 7185 26837 7186 26849
rect 7080 26815 7114 26837
rect 7152 26815 7186 26837
rect 7080 26742 7114 26776
rect 7152 26742 7186 26776
rect 7080 26697 7083 26703
rect 7083 26697 7114 26703
rect 7152 26697 7185 26703
rect 7185 26697 7186 26703
rect 7080 26669 7114 26697
rect 7152 26669 7186 26697
rect 7080 26596 7114 26630
rect 7152 26596 7186 26630
rect 7080 26523 7114 26557
rect 7152 26523 7186 26557
rect 7080 26451 7114 26484
rect 7152 26451 7186 26484
rect 7080 26450 7083 26451
rect 7083 26450 7114 26451
rect 7152 26450 7185 26451
rect 7185 26450 7186 26451
rect 7080 26377 7114 26411
rect 7152 26377 7186 26411
rect 7080 26311 7114 26338
rect 7152 26311 7186 26338
rect 7080 26304 7083 26311
rect 7083 26304 7114 26311
rect 7152 26304 7185 26311
rect 7185 26304 7186 26311
rect 7080 26231 7114 26265
rect 7152 26231 7186 26265
rect 7080 26171 7114 26192
rect 7152 26171 7186 26192
rect 7080 26158 7083 26171
rect 7083 26158 7114 26171
rect 7152 26158 7185 26171
rect 7185 26158 7186 26171
rect 7080 26085 7114 26119
rect 7152 26085 7186 26119
rect 7080 26031 7114 26046
rect 7152 26031 7186 26046
rect 7080 26012 7083 26031
rect 7083 26012 7114 26031
rect 7152 26012 7185 26031
rect 7185 26012 7186 26031
rect 7080 25939 7114 25973
rect 7152 25939 7186 25973
rect 7080 25891 7114 25900
rect 7152 25891 7186 25900
rect 7080 25866 7083 25891
rect 7083 25866 7114 25891
rect 7152 25866 7185 25891
rect 7185 25866 7186 25891
rect 7080 25793 7114 25827
rect 7152 25793 7186 25827
rect 7080 25751 7114 25754
rect 7152 25751 7186 25754
rect 7080 25720 7083 25751
rect 7083 25720 7114 25751
rect 7152 25720 7185 25751
rect 7185 25720 7186 25751
rect 7080 25647 7114 25681
rect 7152 25647 7186 25681
rect 7080 25577 7083 25608
rect 7083 25577 7114 25608
rect 7152 25577 7185 25608
rect 7185 25577 7186 25608
rect 7080 25574 7114 25577
rect 7152 25574 7186 25577
rect 7080 25501 7114 25535
rect 7152 25501 7186 25535
rect 7080 25437 7083 25462
rect 7083 25437 7114 25462
rect 7152 25437 7185 25462
rect 7185 25437 7186 25462
rect 7080 25428 7114 25437
rect 7152 25428 7186 25437
rect 7080 25355 7114 25389
rect 7152 25355 7186 25389
rect 7080 25296 7083 25316
rect 7083 25296 7114 25316
rect 7152 25296 7185 25316
rect 7185 25296 7186 25316
rect 7080 25282 7114 25296
rect 7152 25282 7186 25296
rect 7080 25209 7114 25243
rect 7152 25209 7186 25243
rect 7080 25155 7083 25170
rect 7083 25155 7114 25170
rect 7152 25155 7185 25170
rect 7185 25155 7186 25170
rect 7080 25136 7114 25155
rect 7152 25136 7186 25155
rect 7080 25063 7114 25097
rect 7152 25063 7186 25097
rect 7080 25014 7083 25024
rect 7083 25014 7114 25024
rect 7152 25014 7185 25024
rect 7185 25014 7186 25024
rect 7080 24990 7114 25014
rect 7152 24990 7186 25014
rect 7080 24917 7114 24951
rect 7152 24917 7186 24951
rect 7080 24873 7083 24878
rect 7083 24873 7114 24878
rect 7152 24873 7185 24878
rect 7185 24873 7186 24878
rect 7080 24844 7114 24873
rect 7152 24844 7186 24873
rect 7080 24771 7114 24805
rect 7152 24771 7186 24805
rect 7080 24698 7114 24732
rect 7152 24698 7186 24732
rect 7080 24625 7114 24659
rect 7152 24625 7186 24659
rect 7080 24552 7114 24586
rect 7152 24552 7186 24586
rect 4062 24483 4080 24517
rect 4080 24483 4096 24517
rect 4135 24483 4150 24517
rect 4150 24483 4169 24517
rect 4208 24483 4220 24517
rect 4220 24483 4242 24517
rect 4281 24483 4290 24517
rect 4290 24483 4315 24517
rect 4354 24483 4360 24517
rect 4360 24483 4388 24517
rect 4427 24483 4430 24517
rect 4430 24483 4461 24517
rect 4500 24483 4534 24517
rect 4573 24483 4606 24517
rect 4606 24483 4607 24517
rect 4646 24483 4675 24517
rect 4675 24483 4680 24517
rect 4719 24483 4744 24517
rect 4744 24483 4753 24517
rect 4792 24483 4813 24517
rect 4813 24483 4826 24517
rect 4865 24483 4882 24517
rect 4882 24483 4899 24517
rect 4938 24483 4951 24517
rect 4951 24483 4972 24517
rect 5011 24483 5020 24517
rect 5020 24483 5045 24517
rect 5084 24483 5089 24517
rect 5089 24483 5118 24517
rect 5157 24483 5158 24517
rect 5158 24483 5191 24517
rect 5230 24483 5261 24517
rect 5261 24483 5264 24517
rect 5303 24483 5330 24517
rect 5330 24483 5337 24517
rect 5376 24483 5399 24517
rect 5399 24483 5410 24517
rect 5449 24483 5468 24517
rect 5468 24483 5483 24517
rect 5522 24483 5537 24517
rect 5537 24483 5556 24517
rect 5595 24483 5606 24517
rect 5606 24483 5629 24517
rect 5667 24483 5675 24517
rect 5675 24483 5701 24517
rect 5739 24483 5744 24517
rect 5744 24483 5773 24517
rect 5811 24483 5813 24517
rect 5813 24483 5845 24517
rect 5883 24483 5917 24517
rect 5955 24483 5986 24517
rect 5986 24483 5989 24517
rect 6027 24483 6055 24517
rect 6055 24483 6061 24517
rect 4062 24347 4080 24381
rect 4080 24347 4096 24381
rect 4135 24347 4150 24381
rect 4150 24347 4169 24381
rect 4208 24347 4220 24381
rect 4220 24347 4242 24381
rect 4281 24347 4290 24381
rect 4290 24347 4315 24381
rect 4354 24347 4360 24381
rect 4360 24347 4388 24381
rect 4427 24347 4430 24381
rect 4430 24347 4461 24381
rect 4500 24347 4534 24381
rect 4573 24347 4606 24381
rect 4606 24347 4607 24381
rect 4646 24347 4675 24381
rect 4675 24347 4680 24381
rect 4719 24347 4744 24381
rect 4744 24347 4753 24381
rect 4792 24347 4813 24381
rect 4813 24347 4826 24381
rect 4865 24347 4882 24381
rect 4882 24347 4899 24381
rect 4938 24347 4951 24381
rect 4951 24347 4972 24381
rect 5011 24347 5020 24381
rect 5020 24347 5045 24381
rect 5084 24347 5089 24381
rect 5089 24347 5118 24381
rect 5157 24347 5158 24381
rect 5158 24347 5191 24381
rect 5230 24347 5261 24381
rect 5261 24347 5264 24381
rect 5303 24347 5330 24381
rect 5330 24347 5337 24381
rect 5376 24347 5399 24381
rect 5399 24347 5410 24381
rect 5449 24347 5468 24381
rect 5468 24347 5483 24381
rect 5522 24347 5537 24381
rect 5537 24347 5556 24381
rect 5595 24347 5606 24381
rect 5606 24347 5629 24381
rect 5667 24347 5675 24381
rect 5675 24347 5701 24381
rect 5739 24347 5744 24381
rect 5744 24347 5773 24381
rect 5811 24347 5813 24381
rect 5813 24347 5845 24381
rect 5883 24347 5917 24381
rect 5955 24347 5986 24381
rect 5986 24347 5989 24381
rect 6027 24347 6055 24381
rect 6055 24347 6061 24381
rect 7080 24484 7114 24513
rect 7152 24484 7186 24513
rect 7080 24479 7083 24484
rect 7083 24479 7114 24484
rect 7152 24479 7185 24484
rect 7185 24479 7186 24484
rect 7080 24406 7114 24440
rect 7152 24406 7186 24440
rect 7080 24343 7114 24367
rect 7152 24343 7186 24367
rect 7080 24333 7083 24343
rect 7083 24333 7114 24343
rect 7152 24333 7185 24343
rect 7185 24333 7186 24343
rect 7080 24260 7114 24294
rect 7152 24260 7186 24294
rect 7080 24202 7114 24221
rect 7152 24202 7186 24221
rect 7080 24187 7083 24202
rect 7083 24187 7114 24202
rect 7152 24187 7185 24202
rect 7185 24187 7186 24202
rect 7080 24114 7114 24148
rect 7152 24114 7186 24148
rect 7080 24061 7114 24075
rect 7152 24061 7186 24075
rect 7080 24041 7083 24061
rect 7083 24041 7114 24061
rect 7152 24041 7185 24061
rect 7185 24041 7186 24061
rect 7080 23968 7114 24002
rect 7152 23968 7186 24002
rect 7080 23920 7114 23929
rect 7152 23920 7186 23929
rect 7080 23895 7083 23920
rect 7083 23895 7114 23920
rect 7152 23895 7185 23920
rect 7185 23895 7186 23920
rect 7080 23822 7114 23856
rect 7152 23822 7186 23856
rect 7080 23779 7114 23782
rect 7152 23779 7186 23782
rect 7080 23748 7083 23779
rect 7083 23748 7114 23779
rect 7152 23748 7185 23779
rect 7185 23748 7186 23779
rect 7080 23674 7114 23708
rect 7152 23674 7186 23708
rect 7080 23604 7083 23634
rect 7083 23604 7114 23634
rect 7152 23604 7185 23634
rect 7185 23604 7186 23634
rect 7080 23600 7114 23604
rect 7152 23600 7186 23604
rect 7080 23526 7114 23560
rect 7152 23526 7186 23560
rect 7080 23463 7083 23486
rect 7083 23463 7114 23486
rect 7152 23463 7185 23486
rect 7185 23463 7186 23486
rect 7080 23452 7114 23463
rect 7152 23452 7186 23463
rect 7080 23378 7114 23412
rect 7152 23378 7186 23412
rect 6067 23246 7757 23256
rect 6067 23212 6089 23246
rect 6089 23212 6123 23246
rect 6123 23212 6230 23246
rect 6230 23212 6264 23246
rect 6264 23212 6372 23246
rect 6372 23212 6406 23246
rect 6406 23212 6514 23246
rect 6514 23212 6548 23246
rect 6548 23212 6656 23246
rect 6656 23212 6690 23246
rect 6690 23212 6798 23246
rect 6798 23212 6832 23246
rect 6832 23212 6940 23246
rect 6940 23212 6974 23246
rect 6974 23212 7082 23246
rect 7082 23212 7116 23246
rect 7116 23212 7224 23246
rect 7224 23212 7258 23246
rect 7258 23212 7366 23246
rect 7366 23212 7400 23246
rect 7400 23212 7508 23246
rect 7508 23212 7542 23246
rect 7542 23212 7650 23246
rect 7650 23212 7684 23246
rect 7684 23212 7757 23246
rect 6067 23144 7757 23212
rect 6067 23110 6089 23144
rect 6089 23110 6123 23144
rect 6123 23110 6230 23144
rect 6230 23110 6264 23144
rect 6264 23110 6372 23144
rect 6372 23110 6406 23144
rect 6406 23110 6514 23144
rect 6514 23110 6548 23144
rect 6548 23110 6656 23144
rect 6656 23110 6690 23144
rect 6690 23110 6798 23144
rect 6798 23110 6832 23144
rect 6832 23110 6940 23144
rect 6940 23110 6974 23144
rect 6974 23110 7082 23144
rect 7082 23110 7116 23144
rect 7116 23110 7224 23144
rect 7224 23110 7258 23144
rect 7258 23110 7366 23144
rect 7366 23110 7400 23144
rect 7400 23110 7508 23144
rect 7508 23110 7542 23144
rect 7542 23110 7650 23144
rect 7650 23110 7684 23144
rect 7684 23110 7757 23144
rect 6067 23042 7757 23110
rect 6067 23008 6089 23042
rect 6089 23008 6123 23042
rect 6123 23008 6230 23042
rect 6230 23008 6264 23042
rect 6264 23008 6372 23042
rect 6372 23008 6406 23042
rect 6406 23008 6514 23042
rect 6514 23008 6548 23042
rect 6548 23008 6656 23042
rect 6656 23008 6690 23042
rect 6690 23008 6798 23042
rect 6798 23008 6832 23042
rect 6832 23008 6940 23042
rect 6940 23008 6974 23042
rect 6974 23008 7082 23042
rect 7082 23008 7116 23042
rect 7116 23008 7224 23042
rect 7224 23008 7258 23042
rect 7258 23008 7366 23042
rect 7366 23008 7400 23042
rect 7400 23008 7508 23042
rect 7508 23008 7542 23042
rect 7542 23008 7650 23042
rect 7650 23008 7684 23042
rect 7684 23008 7757 23042
rect 6067 22940 7757 23008
rect 6067 22906 6089 22940
rect 6089 22906 6123 22940
rect 6123 22906 6230 22940
rect 6230 22906 6264 22940
rect 6264 22906 6372 22940
rect 6372 22906 6406 22940
rect 6406 22906 6514 22940
rect 6514 22906 6548 22940
rect 6548 22906 6656 22940
rect 6656 22906 6690 22940
rect 6690 22906 6798 22940
rect 6798 22906 6832 22940
rect 6832 22906 6940 22940
rect 6940 22906 6974 22940
rect 6974 22906 7082 22940
rect 7082 22906 7116 22940
rect 7116 22906 7224 22940
rect 7224 22906 7258 22940
rect 7258 22906 7366 22940
rect 7366 22906 7400 22940
rect 7400 22906 7508 22940
rect 7508 22906 7542 22940
rect 7542 22906 7650 22940
rect 7650 22906 7684 22940
rect 7684 22906 7757 22940
rect 6067 22838 7757 22906
rect 6067 22804 6089 22838
rect 6089 22804 6123 22838
rect 6123 22804 6230 22838
rect 6230 22804 6264 22838
rect 6264 22804 6372 22838
rect 6372 22804 6406 22838
rect 6406 22804 6514 22838
rect 6514 22804 6548 22838
rect 6548 22804 6656 22838
rect 6656 22804 6690 22838
rect 6690 22804 6798 22838
rect 6798 22804 6832 22838
rect 6832 22804 6940 22838
rect 6940 22804 6974 22838
rect 6974 22804 7082 22838
rect 7082 22804 7116 22838
rect 7116 22804 7224 22838
rect 7224 22804 7258 22838
rect 7258 22804 7366 22838
rect 7366 22804 7400 22838
rect 7400 22804 7508 22838
rect 7508 22804 7542 22838
rect 7542 22804 7650 22838
rect 7650 22804 7684 22838
rect 7684 22804 7757 22838
rect 6067 22790 7757 22804
rect 6067 22736 6101 22751
rect 6067 22717 6089 22736
rect 6089 22717 6101 22736
rect 6139 22717 6173 22751
rect 6211 22736 6245 22751
rect 6211 22717 6230 22736
rect 6230 22717 6245 22736
rect 6283 22717 6317 22751
rect 6355 22736 6389 22751
rect 6355 22717 6372 22736
rect 6372 22717 6389 22736
rect 6427 22717 6461 22751
rect 6499 22736 6533 22751
rect 6499 22717 6514 22736
rect 6514 22717 6533 22736
rect 6571 22717 6605 22751
rect 6643 22736 6677 22751
rect 6643 22717 6656 22736
rect 6656 22717 6677 22736
rect 6715 22717 6749 22751
rect 6787 22736 6821 22751
rect 6787 22717 6798 22736
rect 6798 22717 6821 22736
rect 6859 22717 6893 22751
rect 6931 22736 6965 22751
rect 6931 22717 6940 22736
rect 6940 22717 6965 22736
rect 7003 22717 7037 22751
rect 7075 22736 7109 22751
rect 7075 22717 7082 22736
rect 7082 22717 7109 22736
rect 7147 22717 7181 22751
rect 7219 22736 7253 22751
rect 7219 22717 7224 22736
rect 7224 22717 7253 22736
rect 7291 22717 7325 22751
rect 7363 22736 7397 22751
rect 7363 22717 7366 22736
rect 7366 22717 7397 22736
rect 7435 22717 7469 22751
rect 7507 22736 7541 22751
rect 7507 22717 7508 22736
rect 7508 22717 7541 22736
rect 7579 22717 7613 22751
rect 7651 22736 7685 22751
rect 7651 22717 7684 22736
rect 7684 22717 7685 22736
rect 7723 22717 7757 22751
rect 6067 22644 6101 22678
rect 6139 22644 6173 22678
rect 6211 22644 6245 22678
rect 6283 22644 6317 22678
rect 6355 22644 6389 22678
rect 6427 22644 6461 22678
rect 6499 22644 6533 22678
rect 6571 22644 6605 22678
rect 6643 22644 6677 22678
rect 6715 22644 6749 22678
rect 6787 22644 6821 22678
rect 6859 22644 6893 22678
rect 6931 22644 6965 22678
rect 7003 22644 7037 22678
rect 7075 22644 7109 22678
rect 7147 22644 7181 22678
rect 7219 22644 7253 22678
rect 7291 22644 7325 22678
rect 7363 22644 7397 22678
rect 7435 22644 7469 22678
rect 7507 22644 7541 22678
rect 7579 22644 7613 22678
rect 7651 22644 7685 22678
rect 7723 22644 7757 22678
rect 6067 22600 6089 22605
rect 6089 22600 6101 22605
rect 6067 22571 6101 22600
rect 6139 22571 6173 22605
rect 6211 22600 6230 22605
rect 6230 22600 6245 22605
rect 6211 22571 6245 22600
rect 6283 22571 6317 22605
rect 6355 22600 6372 22605
rect 6372 22600 6389 22605
rect 6355 22571 6389 22600
rect 6427 22571 6461 22605
rect 6499 22600 6514 22605
rect 6514 22600 6533 22605
rect 6499 22571 6533 22600
rect 6571 22571 6605 22605
rect 6643 22600 6656 22605
rect 6656 22600 6677 22605
rect 6643 22571 6677 22600
rect 6715 22571 6749 22605
rect 6787 22600 6798 22605
rect 6798 22600 6821 22605
rect 6787 22571 6821 22600
rect 6859 22571 6893 22605
rect 6931 22600 6940 22605
rect 6940 22600 6965 22605
rect 6931 22571 6965 22600
rect 7003 22571 7037 22605
rect 7075 22600 7082 22605
rect 7082 22600 7109 22605
rect 7075 22571 7109 22600
rect 7147 22571 7181 22605
rect 7219 22600 7224 22605
rect 7224 22600 7253 22605
rect 7219 22571 7253 22600
rect 7291 22571 7325 22605
rect 7363 22600 7366 22605
rect 7366 22600 7397 22605
rect 7363 22571 7397 22600
rect 7435 22571 7469 22605
rect 7507 22600 7508 22605
rect 7508 22600 7541 22605
rect 7507 22571 7541 22600
rect 7579 22571 7613 22605
rect 7651 22600 7684 22605
rect 7684 22600 7685 22605
rect 7651 22571 7685 22600
rect 7723 22571 7757 22605
rect 6067 22498 6089 22532
rect 6089 22498 6101 22532
rect 6139 22498 6173 22532
rect 6211 22498 6230 22532
rect 6230 22498 6245 22532
rect 6283 22498 6317 22532
rect 6355 22498 6372 22532
rect 6372 22498 6389 22532
rect 6427 22498 6461 22532
rect 6499 22498 6514 22532
rect 6514 22498 6533 22532
rect 6571 22498 6605 22532
rect 6643 22498 6656 22532
rect 6656 22498 6677 22532
rect 6715 22498 6749 22532
rect 6787 22498 6798 22532
rect 6798 22498 6821 22532
rect 6859 22498 6893 22532
rect 6931 22498 6940 22532
rect 6940 22498 6965 22532
rect 7003 22498 7037 22532
rect 7075 22498 7082 22532
rect 7082 22498 7109 22532
rect 7147 22498 7181 22532
rect 7219 22498 7224 22532
rect 7224 22498 7253 22532
rect 7291 22498 7325 22532
rect 7363 22498 7366 22532
rect 7366 22498 7397 22532
rect 7435 22498 7469 22532
rect 7507 22498 7508 22532
rect 7508 22498 7541 22532
rect 7579 22498 7613 22532
rect 7651 22498 7684 22532
rect 7684 22498 7685 22532
rect 7723 22498 7757 22532
rect 6373 19693 6407 19694
rect 6373 19660 6407 19693
rect 6972 19625 7006 19659
rect 7052 19625 7086 19659
rect 7132 19625 7166 19659
rect 7212 19625 7246 19659
rect 7292 19625 7326 19659
rect 7372 19625 7406 19659
rect 7451 19625 7485 19659
rect 7530 19625 7564 19659
rect 7716 19632 7750 19666
rect 6373 19621 6407 19622
rect 6373 19588 6407 19621
rect 6373 19549 6407 19550
rect 6373 19516 6407 19549
rect 7624 19598 7658 19602
rect 7624 19568 7658 19598
rect 7624 19503 7658 19508
rect 6373 19477 6407 19478
rect 6373 19444 6407 19477
rect 7116 19469 7150 19503
rect 7199 19469 7233 19503
rect 7282 19469 7316 19503
rect 7365 19469 7399 19503
rect 7448 19469 7482 19503
rect 7530 19469 7564 19503
rect 7624 19474 7658 19503
rect 6373 19371 6407 19405
rect 7624 19408 7658 19414
rect 7624 19380 7658 19408
rect 7716 19588 7750 19594
rect 7716 19560 7750 19588
rect 7716 19520 7750 19522
rect 7716 19488 7750 19520
rect 7716 19418 7750 19450
rect 7716 19416 7750 19418
rect 7716 19350 7750 19378
rect 6972 19313 7006 19347
rect 7058 19313 7092 19347
rect 7144 19313 7178 19347
rect 7230 19313 7264 19347
rect 7316 19313 7350 19347
rect 7402 19313 7436 19347
rect 7716 19344 7750 19350
rect 6373 19211 6407 19231
rect 6373 19197 6407 19211
rect 7624 19252 7658 19280
rect 7624 19246 7658 19252
rect 7144 19157 7178 19191
rect 7222 19157 7256 19191
rect 7299 19157 7333 19191
rect 7376 19157 7410 19191
rect 7453 19157 7487 19191
rect 7530 19157 7564 19191
rect 7624 19182 7658 19206
rect 7624 19172 7658 19182
rect 6373 19140 6407 19156
rect 6373 19122 6407 19140
rect 6373 19069 6407 19081
rect 6373 19047 6407 19069
rect 7624 19112 7658 19132
rect 7624 19098 7658 19112
rect 7624 19042 7658 19058
rect 6373 18997 6407 19006
rect 6972 19001 7006 19035
rect 7058 19001 7092 19035
rect 7144 19001 7178 19035
rect 7230 19001 7264 19035
rect 7316 19001 7350 19035
rect 7402 19001 7436 19035
rect 7624 19024 7658 19042
rect 6373 18972 6407 18997
rect 6373 18925 6407 18931
rect 6373 18897 6407 18925
rect 7624 18972 7658 18984
rect 7624 18950 7658 18972
rect 7624 18902 7658 18910
rect 6373 18853 6407 18856
rect 6373 18822 6407 18853
rect 7144 18845 7178 18879
rect 7222 18845 7256 18879
rect 7299 18845 7333 18879
rect 7376 18845 7410 18879
rect 7453 18845 7487 18879
rect 7530 18845 7564 18879
rect 7624 18876 7658 18902
rect 6373 18747 6407 18781
rect 7624 18832 7658 18836
rect 7624 18802 7658 18832
rect 7624 18728 7658 18762
rect 6972 18689 7006 18723
rect 7058 18689 7092 18723
rect 7144 18689 7178 18723
rect 7230 18689 7264 18723
rect 7316 18689 7350 18723
rect 7402 18689 7436 18723
rect 7624 18656 7658 18688
rect 7624 18654 7658 18656
rect 6373 18587 6407 18614
rect 6373 18580 6407 18587
rect 7624 18586 7658 18614
rect 7624 18580 7658 18586
rect 6373 18519 6407 18542
rect 7144 18533 7178 18567
rect 7222 18533 7256 18567
rect 7299 18533 7333 18567
rect 7376 18533 7410 18567
rect 7453 18533 7487 18567
rect 7530 18533 7564 18567
rect 6373 18508 6407 18519
rect 7624 18515 7658 18540
rect 7624 18506 7658 18515
rect 7624 18444 7658 18466
rect 7624 18432 7658 18444
rect 6972 18377 7006 18411
rect 7058 18377 7092 18411
rect 7144 18377 7178 18411
rect 7230 18377 7264 18411
rect 7316 18377 7350 18411
rect 7402 18377 7436 18411
rect 7624 18373 7658 18392
rect 7624 18358 7658 18373
rect 7624 18302 7658 18318
rect 7624 18284 7658 18302
rect 7144 18221 7178 18255
rect 7222 18221 7256 18255
rect 7299 18221 7333 18255
rect 7376 18221 7410 18255
rect 7453 18221 7487 18255
rect 7530 18221 7564 18255
rect 7624 18231 7658 18244
rect 7624 18210 7658 18231
rect 7624 18160 7658 18170
rect 7624 18136 7658 18160
rect 7716 19282 7750 19306
rect 7716 19272 7750 19282
rect 7716 19214 7750 19234
rect 7716 19200 7750 19214
rect 7716 19146 7750 19162
rect 7716 19128 7750 19146
rect 7716 19078 7750 19090
rect 7716 19056 7750 19078
rect 7716 19010 7750 19018
rect 7716 18984 7750 19010
rect 7716 18942 7750 18946
rect 7716 18912 7750 18942
rect 7716 18840 7750 18874
rect 7716 18772 7750 18802
rect 7716 18768 7750 18772
rect 7716 18704 7750 18730
rect 7716 18696 7750 18704
rect 7716 18636 7750 18658
rect 7716 18624 7750 18636
rect 7716 18568 7750 18586
rect 7716 18552 7750 18568
rect 7716 18500 7750 18514
rect 7716 18480 7750 18500
rect 7716 18432 7750 18441
rect 7716 18407 7750 18432
rect 7716 18364 7750 18368
rect 7716 18334 7750 18364
rect 7716 18262 7750 18295
rect 7716 18261 7750 18262
rect 7716 18194 7750 18222
rect 7716 18188 7750 18194
rect 7716 18126 7750 18149
rect 7716 18115 7750 18126
rect 6972 18065 7006 18099
rect 7058 18065 7092 18099
rect 7144 18065 7178 18099
rect 7230 18065 7264 18099
rect 7316 18065 7350 18099
rect 7402 18065 7436 18099
rect 7716 18058 7750 18076
rect 7624 18038 7658 18040
rect 7624 18006 7658 18038
rect 7144 17909 7178 17943
rect 7222 17909 7256 17943
rect 7299 17909 7333 17943
rect 7376 17909 7410 17943
rect 7453 17909 7487 17943
rect 7530 17909 7564 17943
rect 7624 17935 7658 17968
rect 7624 17934 7658 17935
rect 7716 18042 7750 18058
rect 7716 17990 7750 18003
rect 7716 17969 7750 17990
rect 7716 17922 7750 17930
rect 7716 17896 7750 17922
rect 7716 17854 7750 17857
rect 6972 17799 7006 17833
rect 7052 17799 7086 17833
rect 7132 17799 7166 17833
rect 7212 17799 7246 17833
rect 7292 17799 7326 17833
rect 7372 17799 7406 17833
rect 7451 17799 7485 17833
rect 7530 17799 7564 17833
rect 7716 17823 7750 17854
rect 7624 17772 7658 17776
rect 7624 17742 7658 17772
rect 7624 17677 7658 17680
rect 7116 17643 7150 17677
rect 7194 17643 7228 17677
rect 7271 17643 7305 17677
rect 7348 17643 7382 17677
rect 7425 17643 7459 17677
rect 7502 17643 7536 17677
rect 7624 17646 7658 17677
rect 7624 17582 7658 17583
rect 7624 17549 7658 17582
rect 7716 17752 7750 17784
rect 7716 17750 7750 17752
rect 7716 17684 7750 17711
rect 7716 17677 7750 17684
rect 7716 17616 7750 17638
rect 7716 17604 7750 17616
rect 7716 17548 7750 17565
rect 7716 17531 7750 17548
rect 6972 17487 7006 17521
rect 7058 17487 7092 17521
rect 7144 17487 7178 17521
rect 7230 17487 7264 17521
rect 7316 17487 7350 17521
rect 7402 17487 7436 17521
rect 7716 17480 7750 17492
rect 7624 17460 7658 17468
rect 7624 17434 7658 17460
rect 7624 17390 7658 17394
rect 7144 17331 7178 17365
rect 7222 17331 7256 17365
rect 7299 17331 7333 17365
rect 7376 17331 7410 17365
rect 7453 17331 7487 17365
rect 7530 17331 7564 17365
rect 7624 17360 7658 17390
rect 7624 17286 7658 17319
rect 7624 17285 7658 17286
rect 7624 17216 7658 17244
rect 7624 17210 7658 17216
rect 6972 17175 7006 17209
rect 7058 17175 7092 17209
rect 7144 17175 7178 17209
rect 7230 17175 7264 17209
rect 7316 17175 7350 17209
rect 7402 17175 7436 17209
rect 7624 17146 7658 17169
rect 7624 17135 7658 17146
rect 7624 17076 7658 17094
rect 7624 17060 7658 17076
rect 7144 17019 7178 17053
rect 7222 17019 7256 17053
rect 7299 17019 7333 17053
rect 7376 17019 7410 17053
rect 7453 17019 7487 17053
rect 7530 17019 7564 17053
rect 7624 17006 7658 17019
rect 7624 16985 7658 17006
rect 7624 16936 7658 16944
rect 7624 16910 7658 16936
rect 6972 16863 7006 16897
rect 7058 16863 7092 16897
rect 7144 16863 7178 16897
rect 7230 16863 7264 16897
rect 7316 16863 7350 16897
rect 7402 16863 7436 16897
rect 7624 16866 7658 16869
rect 7624 16835 7658 16866
rect 7624 16760 7658 16794
rect 7144 16707 7178 16741
rect 7222 16707 7256 16741
rect 7299 16707 7333 16741
rect 7376 16707 7410 16741
rect 7453 16707 7487 16741
rect 7530 16707 7564 16741
rect 7624 16689 7658 16719
rect 7624 16685 7658 16689
rect 7624 16618 7658 16644
rect 7624 16610 7658 16618
rect 6972 16551 7006 16585
rect 7058 16551 7092 16585
rect 7144 16551 7178 16585
rect 7230 16551 7264 16585
rect 7316 16551 7350 16585
rect 7402 16551 7436 16585
rect 7624 16547 7658 16569
rect 7624 16535 7658 16547
rect 7624 16476 7658 16494
rect 7624 16460 7658 16476
rect 7144 16395 7178 16429
rect 7222 16395 7256 16429
rect 7299 16395 7333 16429
rect 7376 16395 7410 16429
rect 7453 16395 7487 16429
rect 7530 16395 7564 16429
rect 7624 16405 7658 16419
rect 7624 16385 7658 16405
rect 7624 16334 7658 16344
rect 7624 16310 7658 16334
rect 7716 17458 7750 17480
rect 7716 17412 7750 17419
rect 7716 17385 7750 17412
rect 7716 17344 7750 17346
rect 7716 17312 7750 17344
rect 7716 17242 7750 17273
rect 7716 17239 7750 17242
rect 7716 17174 7750 17200
rect 7716 17166 7750 17174
rect 7716 17106 7750 17127
rect 7716 17093 7750 17106
rect 7716 17038 7750 17054
rect 7716 17020 7750 17038
rect 7716 16970 7750 16981
rect 7716 16947 7750 16970
rect 7716 16902 7750 16908
rect 7716 16874 7750 16902
rect 7716 16834 7750 16835
rect 7716 16801 7750 16834
rect 7716 16732 7750 16762
rect 7716 16728 7750 16732
rect 7716 16664 7750 16689
rect 7716 16655 7750 16664
rect 7716 16596 7750 16616
rect 7716 16582 7750 16596
rect 7716 16528 7750 16543
rect 7716 16509 7750 16528
rect 7716 16460 7750 16470
rect 7716 16436 7750 16460
rect 7716 16392 7750 16397
rect 7716 16363 7750 16392
rect 7716 16290 7750 16324
rect 6972 16239 7006 16273
rect 7058 16239 7092 16273
rect 7144 16239 7178 16273
rect 7230 16239 7264 16273
rect 7316 16239 7350 16273
rect 7402 16239 7436 16273
rect 7624 16212 7658 16216
rect 7624 16182 7658 16212
rect 7624 16142 7658 16144
rect 7144 16083 7178 16117
rect 7222 16083 7256 16117
rect 7299 16083 7333 16117
rect 7376 16083 7410 16117
rect 7453 16083 7487 16117
rect 7530 16083 7564 16117
rect 7624 16110 7658 16142
rect 7716 16222 7750 16251
rect 7716 16217 7750 16222
rect 7716 16154 7750 16178
rect 7716 16144 7750 16154
rect 7716 16086 7750 16105
rect 7716 16071 7750 16086
rect 7716 16018 7750 16032
rect 6972 15973 7006 16007
rect 7052 15973 7086 16007
rect 7132 15973 7166 16007
rect 7212 15973 7246 16007
rect 7292 15973 7326 16007
rect 7372 15973 7406 16007
rect 7451 15973 7485 16007
rect 7530 15973 7564 16007
rect 7716 15998 7750 16018
rect 7624 15946 7658 15950
rect 7624 15916 7658 15946
rect 7624 15851 7658 15861
rect 7116 15817 7150 15851
rect 7194 15817 7228 15851
rect 7271 15817 7305 15851
rect 7348 15817 7382 15851
rect 7425 15817 7459 15851
rect 7502 15817 7536 15851
rect 7624 15827 7658 15851
rect 7624 15756 7658 15772
rect 7624 15738 7658 15756
rect 7716 15950 7750 15959
rect 7716 15925 7750 15950
rect 7716 15882 7750 15886
rect 7716 15852 7750 15882
rect 7716 15780 7750 15813
rect 7716 15779 7750 15780
rect 7716 15712 7750 15740
rect 7716 15706 7750 15712
rect 6972 15661 7006 15695
rect 7058 15661 7092 15695
rect 7144 15661 7178 15695
rect 7230 15661 7264 15695
rect 7316 15661 7350 15695
rect 7402 15661 7436 15695
rect 7624 15600 7658 15630
rect 7624 15596 7658 15600
rect 7144 15505 7178 15539
rect 7222 15505 7256 15539
rect 7299 15505 7333 15539
rect 7376 15505 7410 15539
rect 7453 15505 7487 15539
rect 7530 15505 7564 15539
rect 7624 15530 7658 15556
rect 7624 15522 7658 15530
rect 7624 15460 7658 15482
rect 7624 15448 7658 15460
rect 7624 15390 7658 15408
rect 6972 15349 7006 15383
rect 7058 15349 7092 15383
rect 7144 15349 7178 15383
rect 7230 15349 7264 15383
rect 7316 15349 7350 15383
rect 7402 15349 7436 15383
rect 7624 15374 7658 15390
rect 7624 15320 7658 15334
rect 7624 15300 7658 15320
rect 7624 15250 7658 15260
rect 7144 15193 7178 15227
rect 7222 15193 7256 15227
rect 7299 15193 7333 15227
rect 7376 15193 7410 15227
rect 7453 15193 7487 15227
rect 7530 15193 7564 15227
rect 7624 15226 7658 15250
rect 7624 15180 7658 15186
rect 7624 15152 7658 15180
rect 7624 15110 7658 15112
rect 7624 15078 7658 15110
rect 6972 15037 7006 15071
rect 7058 15037 7092 15071
rect 7144 15037 7178 15071
rect 7230 15037 7264 15071
rect 7316 15037 7350 15071
rect 7402 15037 7436 15071
rect 7624 15004 7658 15038
rect 7624 14934 7658 14964
rect 7624 14930 7658 14934
rect 7144 14881 7178 14915
rect 7222 14881 7256 14915
rect 7299 14881 7333 14915
rect 7376 14881 7410 14915
rect 7453 14881 7487 14915
rect 7530 14881 7564 14915
rect 7624 14863 7658 14890
rect 7624 14856 7658 14863
rect 7624 14792 7658 14816
rect 7624 14782 7658 14792
rect 6972 14725 7006 14759
rect 7058 14725 7092 14759
rect 7144 14725 7178 14759
rect 7230 14725 7264 14759
rect 7316 14725 7350 14759
rect 7402 14725 7436 14759
rect 7624 14721 7658 14742
rect 7624 14708 7658 14721
rect 7624 14650 7658 14668
rect 7624 14634 7658 14650
rect 7144 14569 7178 14603
rect 7222 14569 7256 14603
rect 7299 14569 7333 14603
rect 7376 14569 7410 14603
rect 7453 14569 7487 14603
rect 7530 14569 7564 14603
rect 7624 14579 7658 14593
rect 7624 14559 7658 14579
rect 7624 14508 7658 14518
rect 7624 14484 7658 14508
rect 7716 15644 7750 15667
rect 7716 15633 7750 15644
rect 7716 15576 7750 15594
rect 7716 15560 7750 15576
rect 7716 15508 7750 15521
rect 7716 15487 7750 15508
rect 7716 15440 7750 15448
rect 7716 15414 7750 15440
rect 7716 15372 7750 15375
rect 7716 15341 7750 15372
rect 7716 15270 7750 15302
rect 7716 15268 7750 15270
rect 7716 15202 7750 15229
rect 7716 15195 7750 15202
rect 7716 15134 7750 15156
rect 7716 15122 7750 15134
rect 7716 15066 7750 15083
rect 7716 15049 7750 15066
rect 7716 14998 7750 15010
rect 7716 14976 7750 14998
rect 7716 14930 7750 14937
rect 7716 14903 7750 14930
rect 7716 14862 7750 14864
rect 7716 14830 7750 14862
rect 7716 14760 7750 14791
rect 7716 14757 7750 14760
rect 7716 14692 7750 14718
rect 7716 14684 7750 14692
rect 7716 14624 7750 14645
rect 7716 14611 7750 14624
rect 7716 14556 7750 14572
rect 7716 14538 7750 14556
rect 7716 14488 7750 14499
rect 7716 14465 7750 14488
rect 6972 14413 7006 14447
rect 7058 14413 7092 14447
rect 7144 14413 7178 14447
rect 7230 14413 7264 14447
rect 7316 14413 7350 14447
rect 7402 14413 7436 14447
rect 7716 14420 7750 14426
rect 7624 14386 7658 14390
rect 7624 14356 7658 14386
rect 7624 14317 7658 14318
rect 7144 14257 7178 14291
rect 7222 14257 7256 14291
rect 7299 14257 7333 14291
rect 7376 14257 7410 14291
rect 7453 14257 7487 14291
rect 7530 14257 7564 14291
rect 7624 14284 7658 14317
rect 7716 14392 7750 14420
rect 7716 14352 7750 14353
rect 7716 14319 7750 14352
rect 7716 14246 7750 14280
rect 7027 14042 7061 14076
rect 7106 14042 7140 14076
rect 7185 14042 7219 14076
rect 7530 14042 7564 14076
rect 7629 14042 7663 14076
rect 6364 14006 6398 14037
rect 6364 14003 6398 14006
rect 6364 13937 6398 13964
rect 6364 13930 6398 13937
rect 6364 13868 6398 13891
rect 6364 13857 6398 13868
rect 6364 13799 6398 13817
rect 6364 13783 6398 13799
rect 6364 13730 6398 13743
rect 6364 13709 6398 13730
rect 6364 13661 6398 13669
rect 6364 13635 6398 13661
rect 6364 13591 6398 13595
rect 6364 13561 6398 13591
rect 6364 13487 6398 13521
rect 6364 13415 6398 13447
rect 6670 13948 6704 13979
rect 6670 13945 6704 13948
rect 6670 13877 6704 13898
rect 6670 13864 6704 13877
rect 6670 13806 6704 13817
rect 6670 13783 6704 13806
rect 6670 13734 6704 13735
rect 6670 13701 6704 13734
rect 6670 13624 6704 13653
rect 6670 13619 6704 13624
rect 7815 14015 7849 14019
rect 7815 13985 7849 14015
rect 7027 13886 7061 13920
rect 7169 13886 7203 13920
rect 7304 13911 7338 13945
rect 6833 13876 6867 13880
rect 6833 13846 6867 13876
rect 6833 13739 6867 13773
rect 7423 13886 7457 13920
rect 7526 13886 7560 13920
rect 7629 13886 7663 13920
rect 7815 13911 7849 13931
rect 7815 13897 7849 13911
rect 7304 13868 7338 13873
rect 7304 13839 7338 13868
rect 7304 13800 7338 13801
rect 7304 13767 7338 13800
rect 6959 13730 6993 13764
rect 7035 13730 7069 13764
rect 7110 13730 7144 13764
rect 7185 13730 7219 13764
rect 7815 13842 7849 13843
rect 7815 13809 7849 13842
rect 6833 13635 6867 13665
rect 6833 13631 6867 13635
rect 7521 13730 7555 13764
rect 7629 13730 7663 13764
rect 7815 13738 7849 13754
rect 7304 13698 7338 13729
rect 7304 13695 7338 13698
rect 7304 13630 7338 13657
rect 7304 13623 7338 13630
rect 7027 13574 7061 13608
rect 7169 13574 7203 13608
rect 7815 13720 7849 13738
rect 7815 13635 7849 13665
rect 7815 13631 7849 13635
rect 6670 13552 6704 13571
rect 6670 13537 6704 13552
rect 6670 13480 6704 13489
rect 6670 13455 6704 13480
rect 6833 13547 6867 13554
rect 6833 13520 6867 13547
rect 6833 13475 6867 13482
rect 6833 13448 6867 13475
rect 7304 13562 7338 13585
rect 7423 13574 7457 13608
rect 7526 13574 7560 13608
rect 7629 13574 7663 13608
rect 7304 13551 7338 13562
rect 7304 13494 7338 13513
rect 7304 13479 7338 13494
rect 6364 13413 6398 13415
rect 6937 13418 6971 13452
rect 7016 13418 7050 13452
rect 7095 13418 7129 13452
rect 7815 13547 7849 13563
rect 7815 13529 7849 13547
rect 7815 13475 7849 13490
rect 7815 13456 7849 13475
rect 7304 13426 7338 13441
rect 6833 13403 6867 13410
rect 6833 13376 6867 13403
rect 6364 13345 6398 13373
rect 6364 13339 6398 13345
rect 6364 13275 6398 13299
rect 6364 13265 6398 13275
rect 6364 13205 6398 13225
rect 6364 13191 6398 13205
rect 6364 13135 6398 13151
rect 6364 13117 6398 13135
rect 6364 13065 6398 13077
rect 6364 13043 6398 13065
rect 6364 12995 6398 13003
rect 6364 12969 6398 12995
rect 6364 12925 6398 12929
rect 6364 12895 6398 12925
rect 6364 12821 6398 12855
rect 6670 13324 6704 13348
rect 6670 13314 6704 13324
rect 6670 13253 6704 13267
rect 6670 13233 6704 13253
rect 6670 13182 6704 13186
rect 6670 13152 6704 13182
rect 6670 13072 6704 13105
rect 6670 13071 6704 13072
rect 6670 13000 6704 13024
rect 6670 12990 6704 13000
rect 6833 13331 6867 13338
rect 6833 13304 6867 13331
rect 7304 13407 7338 13426
rect 7507 13418 7541 13452
rect 7608 13418 7642 13452
rect 7709 13418 7743 13452
rect 7304 13358 7338 13369
rect 7304 13335 7338 13358
rect 6833 13259 6867 13266
rect 7027 13262 7061 13296
rect 7100 13262 7134 13296
rect 7173 13262 7207 13296
rect 7304 13289 7338 13297
rect 7815 13403 7849 13417
rect 7815 13383 7849 13403
rect 7815 13331 7849 13344
rect 7815 13310 7849 13331
rect 7304 13263 7338 13289
rect 6833 13232 6867 13259
rect 6833 13187 6867 13194
rect 6833 13160 6867 13187
rect 7423 13262 7457 13296
rect 7526 13262 7560 13296
rect 7629 13262 7663 13296
rect 7304 13220 7338 13225
rect 7304 13191 7338 13220
rect 7304 13151 7338 13152
rect 6833 13116 6867 13121
rect 6833 13087 6867 13116
rect 6937 13106 6971 13140
rect 7016 13106 7050 13140
rect 7095 13106 7129 13140
rect 7304 13118 7338 13151
rect 7815 13259 7849 13270
rect 7815 13236 7849 13259
rect 7815 13187 7849 13196
rect 7815 13162 7849 13187
rect 6833 13045 6867 13048
rect 6833 13014 6867 13045
rect 7505 13106 7539 13140
rect 7607 13106 7641 13140
rect 7709 13106 7743 13140
rect 7815 13116 7849 13122
rect 7304 13048 7338 13079
rect 7304 13045 7338 13048
rect 7027 12950 7061 12984
rect 7100 12950 7134 12984
rect 7173 12950 7207 12984
rect 7304 12979 7338 13006
rect 7815 13088 7849 13116
rect 7815 13045 7849 13048
rect 7815 13014 7849 13045
rect 7304 12972 7338 12979
rect 6670 12928 6704 12943
rect 6670 12909 6704 12928
rect 7439 12950 7473 12984
rect 7522 12950 7556 12984
rect 7605 12950 7639 12984
rect 7687 12950 7721 12984
rect 7304 12910 7338 12933
rect 7304 12899 7338 12910
rect 6670 12856 6704 12861
rect 6670 12827 6704 12856
rect 7113 12840 7147 12874
rect 7185 12840 7219 12874
rect 7304 12841 7338 12860
rect 6364 12751 6398 12781
rect 6364 12747 6398 12751
rect 6364 12681 6398 12707
rect 6364 12673 6398 12681
rect 6364 12611 6398 12633
rect 6670 12700 6704 12732
rect 6670 12698 6704 12700
rect 6670 12632 6704 12660
rect 6943 12745 6977 12754
rect 6943 12720 6977 12745
rect 7304 12826 7338 12841
rect 7423 12840 7457 12874
rect 7495 12840 7529 12874
rect 7304 12772 7338 12787
rect 7304 12753 7338 12772
rect 7023 12690 7057 12724
rect 7095 12690 7129 12724
rect 7665 12745 7699 12760
rect 7665 12726 7699 12745
rect 7304 12703 7338 12714
rect 6943 12648 6977 12682
rect 7304 12680 7338 12703
rect 7499 12690 7533 12724
rect 7571 12690 7605 12724
rect 7665 12654 7699 12688
rect 6670 12626 6704 12632
rect 6364 12599 6398 12611
rect 6548 12456 6562 12490
rect 6562 12456 6582 12490
rect 6625 12456 6632 12490
rect 6632 12456 6659 12490
rect 6701 12456 6702 12490
rect 6702 12456 6735 12490
rect 6777 12456 6808 12490
rect 6808 12456 6811 12490
rect 6853 12456 6878 12490
rect 6878 12456 6887 12490
rect 6929 12456 6948 12490
rect 6948 12456 6963 12490
rect 7005 12456 7018 12490
rect 7018 12456 7039 12490
rect 7081 12456 7087 12490
rect 7087 12456 7115 12490
rect 7157 12456 7190 12490
rect 7190 12456 7191 12490
rect 7233 12456 7259 12490
rect 7259 12456 7267 12490
rect 7309 12456 7328 12490
rect 7328 12456 7343 12490
rect 7385 12456 7397 12490
rect 7397 12456 7419 12490
rect 7461 12456 7466 12490
rect 7466 12456 7495 12490
rect 7537 12456 7570 12490
rect 7570 12456 7571 12490
rect 7613 12456 7647 12490
rect 6392 12337 6426 12371
rect 6392 12265 6426 12299
rect 6542 12337 6576 12371
rect 6798 12325 6832 12359
rect 6542 12265 6576 12299
rect 6672 12265 6706 12299
rect 6672 12133 6706 12167
rect 7120 12325 7154 12359
rect 6798 12229 6832 12263
rect 6798 12133 6832 12167
rect 6964 12265 6998 12299
rect 6964 12133 6998 12167
rect 7432 12325 7466 12359
rect 7120 12229 7154 12263
rect 7120 12133 7154 12167
rect 7276 12265 7310 12299
rect 7276 12169 7310 12203
rect 6472 12095 6481 12129
rect 6481 12095 6506 12129
rect 6544 12095 6578 12129
rect 7432 12229 7466 12263
rect 7432 12133 7466 12167
rect 7588 12265 7622 12299
rect 7588 12169 7622 12203
rect 7276 12073 7310 12107
rect 7588 12073 7622 12107
rect 7744 12265 7778 12299
rect 7744 12169 7778 12203
rect 7744 12073 7778 12107
rect 6724 11945 6747 11979
rect 6747 11945 6758 11979
rect 6808 11945 6816 11979
rect 6816 11945 6842 11979
rect 6892 11945 6920 11979
rect 6920 11945 6926 11979
rect 6975 11945 6989 11979
rect 6989 11945 7009 11979
rect 7058 11945 7059 11979
rect 7059 11945 7092 11979
rect 7204 11945 7215 11979
rect 7215 11945 7238 11979
rect 7289 11945 7323 11979
rect 7373 11945 7395 11979
rect 7395 11945 7407 11979
rect 7457 11945 7467 11979
rect 7467 11945 7491 11979
rect 7541 11945 7573 11979
rect 7573 11945 7575 11979
rect 5018 11138 5020 11172
rect 5020 11138 5052 11172
rect 5090 11138 5122 11172
rect 5122 11138 5124 11172
rect 5327 11138 5354 11172
rect 5354 11138 5361 11172
rect 5404 11138 5423 11172
rect 5423 11138 5438 11172
rect 5481 11138 5492 11172
rect 5492 11138 5515 11172
rect 5558 11138 5561 11172
rect 5561 11138 5592 11172
rect 5634 11138 5666 11172
rect 5666 11138 5668 11172
rect 5803 11138 5822 11172
rect 5822 11138 5837 11172
rect 5891 11138 5893 11172
rect 5893 11138 5925 11172
rect 5979 11138 6002 11172
rect 6002 11138 6013 11172
rect 6067 11138 6074 11172
rect 6074 11138 6101 11172
rect 6155 11138 6180 11172
rect 6180 11138 6189 11172
rect 3154 11084 3160 11118
rect 3160 11084 3188 11118
rect 3226 11084 3228 11118
rect 3228 11084 3260 11118
rect 3355 11084 3384 11118
rect 3384 11084 3389 11118
rect 3437 11084 3456 11118
rect 3456 11084 3471 11118
rect 3518 11084 3528 11118
rect 3528 11084 3552 11118
rect 3599 11084 3600 11118
rect 3600 11084 3633 11118
rect 3680 11084 3710 11118
rect 3710 11084 3714 11118
rect 3761 11084 3781 11118
rect 3781 11084 3795 11118
rect 3842 11084 3852 11118
rect 3852 11084 3876 11118
rect 3983 11084 4008 11118
rect 4008 11084 4017 11118
rect 4065 11084 4080 11118
rect 4080 11084 4099 11118
rect 4147 11084 4152 11118
rect 4152 11084 4181 11118
rect 4229 11084 4262 11118
rect 4262 11084 4263 11118
rect 4311 11084 4334 11118
rect 4334 11084 4345 11118
rect 4392 11084 4405 11118
rect 4405 11084 4426 11118
rect 4473 11084 4476 11118
rect 4476 11084 4507 11118
rect 5272 11016 5306 11050
rect 4999 10968 5033 11002
rect 4999 10896 5033 10930
rect 5149 10968 5183 11002
rect 5272 10936 5306 10970
rect 5415 11044 5449 11078
rect 5415 10959 5449 10993
rect 5149 10896 5183 10930
rect 5571 11044 5605 11078
rect 5883 11044 5917 11078
rect 5571 10936 5605 10970
rect 5727 10968 5761 11002
rect 5415 10874 5449 10908
rect 6195 11044 6229 11078
rect 5883 10964 5917 10998
rect 6039 10968 6073 11002
rect 5727 10883 5761 10917
rect 3127 10778 3139 10812
rect 3139 10778 3161 10812
rect 3202 10778 3209 10812
rect 3209 10778 3236 10812
rect 3276 10778 3279 10812
rect 3279 10778 3310 10812
rect 3350 10778 3383 10812
rect 3383 10778 3384 10812
rect 3424 10778 3453 10812
rect 3453 10778 3458 10812
rect 3498 10778 3523 10812
rect 3523 10778 3532 10812
rect 3572 10778 3593 10812
rect 3593 10778 3606 10812
rect 3646 10778 3663 10812
rect 3663 10778 3680 10812
rect 3720 10778 3733 10812
rect 3733 10778 3754 10812
rect 3794 10778 3803 10812
rect 3803 10778 3828 10812
rect 3868 10778 3873 10812
rect 3873 10778 3902 10812
rect 3942 10778 3943 10812
rect 3943 10778 3976 10812
rect 4016 10778 4049 10812
rect 4049 10778 4050 10812
rect 4090 10778 4119 10812
rect 4119 10778 4124 10812
rect 4164 10778 4189 10812
rect 4189 10778 4198 10812
rect 4238 10778 4258 10812
rect 4258 10778 4272 10812
rect 4312 10778 4327 10812
rect 4327 10778 4346 10812
rect 4386 10778 4396 10812
rect 4396 10778 4420 10812
rect 4460 10778 4465 10812
rect 4465 10778 4494 10812
rect 4534 10778 4568 10812
rect 5727 10798 5761 10832
rect 6717 11037 6751 11060
rect 6836 11042 6870 11076
rect 6908 11042 6942 11076
rect 7078 11055 7112 11057
rect 6717 11026 6751 11037
rect 6195 10964 6229 10998
rect 6351 10968 6385 11002
rect 6039 10882 6073 10916
rect 6039 10797 6073 10831
rect 6351 10892 6385 10926
rect 6351 10816 6385 10850
rect 6717 10968 6751 10987
rect 6717 10953 6751 10968
rect 7078 11023 7112 11055
rect 7078 10953 7112 10985
rect 7078 10951 7112 10953
rect 6717 10899 6751 10914
rect 6717 10880 6751 10899
rect 6836 10892 6870 10926
rect 6908 10892 6942 10926
rect 6717 10830 6751 10841
rect 6717 10807 6751 10830
rect 6923 10784 6957 10818
rect 7022 10784 7056 10818
rect 7122 10784 7156 10818
rect 6717 10761 6751 10768
rect 6717 10734 6751 10761
rect 4989 10680 5012 10714
rect 5012 10680 5023 10714
rect 5062 10680 5081 10714
rect 5081 10680 5096 10714
rect 5135 10680 5150 10714
rect 5150 10680 5169 10714
rect 5208 10680 5219 10714
rect 5219 10680 5242 10714
rect 5281 10680 5288 10714
rect 5288 10680 5315 10714
rect 5354 10680 5357 10714
rect 5357 10680 5388 10714
rect 5427 10680 5460 10714
rect 5460 10680 5461 10714
rect 5500 10680 5529 10714
rect 5529 10680 5534 10714
rect 5572 10680 5598 10714
rect 5598 10680 5606 10714
rect 5644 10680 5667 10714
rect 5667 10680 5678 10714
rect 5716 10680 5735 10714
rect 5735 10680 5750 10714
rect 5788 10680 5803 10714
rect 5803 10680 5822 10714
rect 5860 10680 5871 10714
rect 5871 10680 5894 10714
rect 5932 10680 5939 10714
rect 5939 10680 5966 10714
rect 6004 10680 6007 10714
rect 6007 10680 6038 10714
rect 6076 10680 6109 10714
rect 6109 10680 6110 10714
rect 6148 10680 6177 10714
rect 6177 10680 6182 10714
rect 6220 10680 6254 10714
rect 6717 10692 6751 10695
rect 6717 10661 6751 10692
rect 7228 10721 7262 10726
rect 7228 10692 7262 10721
rect 6836 10626 6870 10660
rect 6938 10626 6972 10660
rect 7040 10626 7074 10660
rect 6717 10589 6751 10622
rect 6717 10588 6751 10589
rect 6717 10520 6751 10549
rect 6717 10515 6751 10520
rect 7228 10617 7262 10651
rect 7228 10548 7262 10576
rect 7228 10542 7262 10548
rect 6717 10451 6751 10477
rect 6922 10470 6956 10504
rect 7040 10470 7074 10504
rect 7228 10479 7262 10501
rect 6717 10443 6751 10451
rect 6717 10382 6751 10405
rect 6717 10371 6751 10382
rect 7228 10467 7262 10479
rect 7228 10409 7262 10426
rect 7228 10392 7262 10409
rect 6717 10313 6751 10333
rect 6836 10314 6870 10348
rect 6938 10314 6972 10348
rect 7040 10314 7074 10348
rect 6717 10299 6751 10313
rect 6717 10244 6751 10261
rect 6717 10227 6751 10244
rect 7228 10253 7262 10281
rect 7228 10247 7262 10253
rect 6717 10175 6751 10189
rect 6717 10155 6751 10175
rect 6921 10158 6955 10192
rect 7021 10158 7055 10192
rect 7122 10158 7156 10192
rect 7228 10182 7262 10203
rect 7228 10169 7262 10182
rect 6717 10106 6751 10117
rect 6717 10083 6751 10106
rect 6717 10037 6751 10045
rect 6717 10011 6751 10037
rect 7228 10111 7262 10125
rect 7228 10091 7262 10111
rect 7228 10039 7262 10048
rect 6836 10002 6870 10036
rect 6938 10002 6972 10036
rect 7040 10002 7074 10036
rect 7228 10014 7262 10039
rect 6717 9968 6751 9973
rect 6717 9939 6751 9968
rect 6717 9899 6751 9901
rect 6717 9867 6751 9899
rect 7228 9967 7262 9971
rect 7228 9937 7262 9967
rect 6924 9846 6958 9880
rect 7023 9846 7057 9880
rect 7122 9846 7156 9880
rect 7228 9860 7262 9894
rect 6717 9795 6751 9829
rect 6717 9692 6751 9702
rect 6717 9668 6751 9692
rect 6836 9690 6870 9724
rect 6938 9690 6972 9724
rect 7040 9690 7074 9724
rect 6717 9623 6751 9629
rect 6717 9595 6751 9623
rect 7228 9629 7262 9648
rect 7228 9614 7262 9629
rect 6717 9554 6751 9556
rect 6717 9522 6751 9554
rect 6924 9534 6958 9568
rect 7023 9534 7057 9568
rect 7122 9534 7156 9568
rect 7228 9558 7262 9571
rect 7228 9537 7262 9558
rect 6717 9450 6751 9483
rect 6717 9449 6751 9450
rect 7228 9487 7262 9493
rect 7228 9459 7262 9487
rect 6717 9381 6751 9410
rect 6717 9376 6751 9381
rect 6836 9378 6870 9412
rect 6938 9378 6972 9412
rect 7040 9378 7074 9412
rect 7228 9381 7262 9415
rect 6717 9312 6751 9337
rect 6717 9303 6751 9312
rect 6717 9243 6751 9264
rect 7228 9305 7262 9337
rect 7228 9303 7262 9305
rect 6717 9230 6751 9243
rect 6924 9222 6958 9256
rect 7023 9222 7057 9256
rect 7122 9222 7156 9256
rect 7228 9233 7262 9259
rect 7228 9225 7262 9233
rect 6717 9175 6751 9191
rect 6717 9157 6751 9175
rect 6717 9107 6751 9119
rect 7228 9161 7262 9181
rect 7228 9147 7262 9161
rect 6717 9085 6751 9107
rect 6836 9066 6870 9100
rect 6938 9066 6972 9100
rect 7040 9066 7074 9100
rect 6717 9039 6751 9047
rect 6717 9013 6751 9039
rect 6717 8971 6751 8975
rect 6717 8941 6751 8971
rect 7228 9005 7262 9033
rect 7228 8999 7262 9005
rect 6924 8910 6958 8944
rect 7023 8910 7057 8944
rect 7122 8910 7156 8944
rect 7228 8936 7262 8946
rect 7228 8912 7262 8936
rect 6717 8869 6751 8903
rect 6717 8801 6751 8831
rect 6717 8797 6751 8801
rect 7228 8832 7262 8859
rect 7228 8825 7262 8832
rect 6717 8733 6751 8759
rect 6836 8754 6870 8788
rect 6938 8754 6972 8788
rect 7040 8754 7074 8788
rect 7228 8763 7262 8772
rect 6717 8725 6751 8733
rect 6717 8665 6751 8687
rect 6717 8653 6751 8665
rect 7228 8738 7262 8763
rect 7228 8660 7262 8685
rect 7228 8651 7262 8660
rect 6717 8597 6751 8615
rect 6924 8598 6958 8632
rect 7023 8598 7057 8632
rect 7122 8598 7156 8632
rect 6717 8581 6751 8597
rect 6717 8529 6751 8543
rect 6717 8509 6751 8529
rect 6911 8488 6945 8522
rect 6983 8488 7017 8522
rect 6717 8461 6751 8471
rect 6717 8437 6751 8461
rect 7078 8427 7112 8434
rect 7078 8400 7112 8427
rect 6836 8332 6870 8366
rect 6908 8332 6942 8366
rect 7078 8293 7112 8327
rect 2874 7886 2908 7920
rect 2948 7886 2982 7920
rect 3022 7886 3056 7920
rect 3096 7886 3130 7920
rect 3170 7886 3204 7920
rect 3244 7886 3278 7920
rect 3318 7886 3352 7920
rect 3392 7886 3426 7920
rect 3466 7886 3500 7920
rect 3539 7886 3573 7920
rect 3612 7886 3646 7920
rect 3685 7886 3719 7920
rect 3758 7886 3792 7920
rect 3831 7886 3865 7920
rect 3904 7886 3938 7920
rect 3977 7886 4011 7920
rect 4050 7886 4084 7920
rect 4123 7886 4157 7920
rect 4196 7886 4230 7920
rect 4269 7886 4303 7920
rect 4342 7886 4376 7920
rect 4415 7886 4449 7920
rect 4488 7886 4522 7920
rect 4561 7886 4595 7920
rect 4634 7886 4668 7920
rect 4707 7886 4741 7920
rect 4780 7886 4814 7920
rect 4853 7886 4887 7920
rect 4926 7886 4960 7920
rect 4999 7886 5033 7920
rect 5072 7886 5106 7920
rect 5145 7886 5179 7920
rect 5218 7886 5252 7920
rect 5291 7886 5325 7920
rect 5364 7886 5398 7920
rect 5437 7886 5471 7920
rect 5510 7886 5544 7920
rect 5583 7886 5617 7920
rect 5656 7886 5690 7920
rect 5729 7886 5763 7920
rect 5802 7886 5836 7920
rect 5875 7886 5909 7920
rect 5948 7886 5982 7920
rect 6021 7886 6055 7920
rect 6094 7886 6128 7920
rect 6167 7886 6201 7920
rect 6240 7886 6274 7920
rect 6313 7886 6347 7920
rect 6386 7886 6420 7920
rect 6459 7886 6493 7920
rect 6532 7886 6566 7920
rect 6605 7886 6639 7920
rect 6678 7886 6712 7920
rect 6972 7852 7006 7886
rect 7052 7852 7086 7886
rect 7132 7852 7166 7886
rect 7212 7852 7246 7886
rect 7292 7852 7326 7886
rect 7372 7852 7406 7886
rect 7451 7852 7485 7886
rect 7530 7852 7564 7886
rect 7716 7849 7750 7881
rect 7716 7847 7750 7849
rect 7624 7825 7658 7829
rect 7624 7795 7658 7825
rect 7624 7730 7658 7738
rect 7144 7696 7178 7730
rect 7222 7696 7256 7730
rect 7299 7696 7333 7730
rect 7376 7696 7410 7730
rect 7453 7696 7487 7730
rect 7530 7696 7564 7730
rect 7624 7704 7658 7730
rect 7624 7635 7658 7646
rect 7624 7612 7658 7635
rect 7716 7781 7750 7809
rect 7716 7775 7750 7781
rect 7716 7713 7750 7737
rect 7716 7703 7750 7713
rect 7716 7645 7750 7665
rect 7716 7631 7750 7645
rect 7716 7577 7750 7593
rect 6972 7540 7006 7574
rect 7058 7540 7092 7574
rect 7144 7540 7178 7574
rect 7230 7540 7264 7574
rect 7316 7540 7350 7574
rect 7402 7540 7436 7574
rect 7716 7559 7750 7577
rect 7624 7479 7658 7504
rect 7624 7470 7658 7479
rect 7144 7384 7178 7418
rect 7222 7384 7256 7418
rect 7299 7384 7333 7418
rect 7376 7384 7410 7418
rect 7453 7384 7487 7418
rect 7530 7384 7564 7418
rect 7624 7409 7658 7431
rect 7624 7397 7658 7409
rect 7624 7339 7658 7358
rect 7624 7324 7658 7339
rect 7624 7269 7658 7285
rect 6972 7228 7006 7262
rect 7058 7228 7092 7262
rect 7144 7228 7178 7262
rect 7230 7228 7264 7262
rect 7316 7228 7350 7262
rect 7402 7228 7436 7262
rect 7624 7251 7658 7269
rect 7624 7199 7658 7211
rect 7624 7177 7658 7199
rect 7624 7129 7658 7137
rect 7144 7072 7178 7106
rect 7222 7072 7256 7106
rect 7299 7072 7333 7106
rect 7376 7072 7410 7106
rect 7453 7072 7487 7106
rect 7530 7072 7564 7106
rect 7624 7103 7658 7129
rect 7624 7059 7658 7063
rect 7624 7029 7658 7059
rect 7624 6955 7658 6989
rect 6972 6916 7006 6950
rect 7058 6916 7092 6950
rect 7144 6916 7178 6950
rect 7230 6916 7264 6950
rect 7316 6916 7350 6950
rect 7402 6916 7436 6950
rect 7624 6883 7658 6915
rect 7624 6881 7658 6883
rect 7624 6813 7658 6841
rect 7624 6807 7658 6813
rect 7144 6760 7178 6794
rect 7222 6760 7256 6794
rect 7299 6760 7333 6794
rect 7376 6760 7410 6794
rect 7453 6760 7487 6794
rect 7530 6760 7564 6794
rect 7624 6742 7658 6767
rect 7624 6733 7658 6742
rect 7624 6671 7658 6693
rect 7624 6659 7658 6671
rect 6972 6604 7006 6638
rect 7058 6604 7092 6638
rect 7144 6604 7178 6638
rect 7230 6604 7264 6638
rect 7316 6604 7350 6638
rect 7402 6604 7436 6638
rect 7624 6600 7658 6619
rect 7624 6585 7658 6600
rect 7624 6529 7658 6545
rect 7624 6511 7658 6529
rect 7144 6448 7178 6482
rect 7222 6448 7256 6482
rect 7299 6448 7333 6482
rect 7376 6448 7410 6482
rect 7453 6448 7487 6482
rect 7530 6448 7564 6482
rect 7624 6458 7658 6471
rect 7624 6437 7658 6458
rect 7624 6387 7658 6397
rect 7624 6363 7658 6387
rect 7716 7509 7750 7521
rect 7716 7487 7750 7509
rect 7716 7441 7750 7449
rect 7716 7415 7750 7441
rect 7716 7373 7750 7377
rect 7716 7343 7750 7373
rect 7716 7271 7750 7305
rect 7716 7203 7750 7233
rect 7716 7199 7750 7203
rect 7716 7135 7750 7161
rect 7716 7127 7750 7135
rect 7716 7067 7750 7089
rect 7716 7055 7750 7067
rect 7716 6999 7750 7017
rect 7716 6983 7750 6999
rect 7716 6931 7750 6945
rect 7716 6911 7750 6931
rect 7716 6863 7750 6873
rect 7716 6839 7750 6863
rect 7716 6795 7750 6801
rect 7716 6767 7750 6795
rect 7716 6727 7750 6729
rect 7716 6695 7750 6727
rect 7716 6625 7750 6657
rect 7716 6623 7750 6625
rect 7716 6557 7750 6585
rect 7716 6551 7750 6557
rect 7716 6489 7750 6513
rect 7716 6479 7750 6489
rect 7716 6421 7750 6441
rect 7716 6407 7750 6421
rect 7716 6353 7750 6369
rect 7716 6335 7750 6353
rect 6972 6292 7006 6326
rect 7058 6292 7092 6326
rect 7144 6292 7178 6326
rect 7230 6292 7264 6326
rect 7316 6292 7350 6326
rect 7402 6292 7436 6326
rect 7716 6285 7750 6297
rect 7624 6265 7658 6267
rect 7624 6233 7658 6265
rect 7144 6136 7178 6170
rect 7222 6136 7256 6170
rect 7299 6136 7333 6170
rect 7376 6136 7410 6170
rect 7453 6136 7487 6170
rect 7530 6136 7564 6170
rect 7624 6162 7658 6195
rect 7624 6161 7658 6162
rect 7716 6263 7750 6285
rect 7716 6217 7750 6225
rect 7716 6191 7750 6217
rect 7716 6149 7750 6153
rect 7716 6119 7750 6149
rect 6972 6026 7006 6060
rect 7052 6026 7086 6060
rect 7132 6026 7166 6060
rect 7212 6026 7246 6060
rect 7292 6026 7326 6060
rect 7372 6026 7406 6060
rect 7451 6026 7485 6060
rect 7530 6026 7564 6060
rect 7716 6047 7750 6081
rect 7624 5999 7658 6003
rect 7624 5969 7658 5999
rect 7624 5904 7658 5916
rect 7144 5870 7178 5904
rect 7222 5870 7256 5904
rect 7299 5870 7333 5904
rect 7376 5870 7410 5904
rect 7453 5870 7487 5904
rect 7530 5870 7564 5904
rect 7624 5882 7658 5904
rect 7624 5809 7658 5828
rect 7624 5794 7658 5809
rect 7716 5979 7750 6009
rect 7716 5975 7750 5979
rect 7716 5911 7750 5937
rect 7716 5903 7750 5911
rect 7716 5843 7750 5865
rect 7716 5831 7750 5843
rect 7716 5775 7750 5793
rect 7716 5759 7750 5775
rect 6972 5714 7006 5748
rect 7058 5714 7092 5748
rect 7144 5714 7178 5748
rect 7230 5714 7264 5748
rect 7316 5714 7350 5748
rect 7402 5714 7436 5748
rect 7716 5707 7750 5721
rect 7624 5653 7658 5670
rect 7624 5636 7658 5653
rect 7144 5558 7178 5592
rect 7222 5558 7256 5592
rect 7299 5558 7333 5592
rect 7376 5558 7410 5592
rect 7453 5558 7487 5592
rect 7530 5558 7564 5592
rect 7624 5583 7658 5597
rect 7624 5563 7658 5583
rect 7624 5513 7658 5524
rect 7624 5490 7658 5513
rect 7624 5443 7658 5451
rect 6972 5402 7006 5436
rect 7058 5402 7092 5436
rect 7144 5402 7178 5436
rect 7230 5402 7264 5436
rect 7316 5402 7350 5436
rect 7402 5402 7436 5436
rect 7624 5417 7658 5443
rect 7624 5373 7658 5378
rect 7624 5344 7658 5373
rect 7624 5303 7658 5305
rect 7144 5246 7178 5280
rect 7222 5246 7256 5280
rect 7299 5246 7333 5280
rect 7376 5246 7410 5280
rect 7453 5246 7487 5280
rect 7530 5246 7564 5280
rect 7624 5271 7658 5303
rect 7624 5198 7658 5232
rect 7624 5127 7658 5159
rect 7624 5125 7658 5127
rect 6972 5090 7006 5124
rect 7058 5090 7092 5124
rect 7144 5090 7178 5124
rect 7230 5090 7264 5124
rect 7316 5090 7350 5124
rect 7402 5090 7436 5124
rect 7624 5057 7658 5086
rect 7624 5052 7658 5057
rect 7624 4987 7658 5013
rect 7624 4979 7658 4987
rect 7144 4934 7178 4968
rect 7222 4934 7256 4968
rect 7299 4934 7333 4968
rect 7376 4934 7410 4968
rect 7453 4934 7487 4968
rect 7530 4934 7564 4968
rect 7624 4916 7658 4940
rect 7624 4906 7658 4916
rect 7624 4845 7658 4867
rect 7624 4833 7658 4845
rect 6972 4778 7006 4812
rect 7058 4778 7092 4812
rect 7144 4778 7178 4812
rect 7230 4778 7264 4812
rect 7316 4778 7350 4812
rect 7402 4778 7436 4812
rect 7624 4774 7658 4793
rect 7624 4759 7658 4774
rect 7624 4703 7658 4719
rect 7624 4685 7658 4703
rect 7144 4622 7178 4656
rect 7222 4622 7256 4656
rect 7299 4622 7333 4656
rect 7376 4622 7410 4656
rect 7453 4622 7487 4656
rect 7530 4622 7564 4656
rect 7624 4632 7658 4645
rect 7624 4611 7658 4632
rect 7624 4561 7658 4571
rect 7624 4537 7658 4561
rect 7716 5687 7750 5707
rect 7716 5639 7750 5649
rect 7716 5615 7750 5639
rect 7716 5571 7750 5577
rect 7716 5543 7750 5571
rect 7716 5503 7750 5505
rect 7716 5471 7750 5503
rect 7716 5401 7750 5432
rect 7716 5398 7750 5401
rect 7716 5333 7750 5359
rect 7716 5325 7750 5333
rect 7716 5265 7750 5286
rect 7716 5252 7750 5265
rect 7716 5197 7750 5213
rect 7716 5179 7750 5197
rect 7716 5129 7750 5140
rect 7716 5106 7750 5129
rect 7716 5061 7750 5067
rect 7716 5033 7750 5061
rect 7716 4993 7750 4994
rect 7716 4960 7750 4993
rect 7716 4891 7750 4921
rect 7716 4887 7750 4891
rect 7716 4823 7750 4848
rect 7716 4814 7750 4823
rect 7716 4755 7750 4775
rect 7716 4741 7750 4755
rect 7716 4687 7750 4702
rect 7716 4668 7750 4687
rect 7716 4619 7750 4629
rect 7716 4595 7750 4619
rect 7716 4551 7750 4556
rect 7716 4522 7750 4551
rect 6972 4466 7006 4500
rect 7058 4466 7092 4500
rect 7144 4466 7178 4500
rect 7230 4466 7264 4500
rect 7316 4466 7350 4500
rect 7402 4466 7436 4500
rect 7624 4405 7658 4439
rect 7144 4310 7178 4344
rect 7222 4310 7256 4344
rect 7299 4310 7333 4344
rect 7376 4310 7410 4344
rect 7453 4310 7487 4344
rect 7530 4310 7564 4344
rect 7624 4336 7658 4367
rect 7624 4333 7658 4336
rect 7716 4449 7750 4483
rect 7716 4381 7750 4410
rect 7716 4376 7750 4381
rect 7716 4313 7750 4337
rect 7716 4303 7750 4313
rect 7716 4245 7750 4264
rect 6972 4200 7006 4234
rect 7052 4200 7086 4234
rect 7132 4200 7166 4234
rect 7212 4200 7246 4234
rect 7292 4200 7326 4234
rect 7372 4200 7406 4234
rect 7451 4200 7485 4234
rect 7530 4200 7564 4234
rect 7716 4230 7750 4245
rect 7624 4173 7658 4177
rect 7624 4143 7658 4173
rect 7624 4078 7658 4099
rect 7144 4044 7178 4078
rect 7222 4044 7256 4078
rect 7299 4044 7333 4078
rect 7376 4044 7410 4078
rect 7453 4044 7487 4078
rect 7530 4044 7564 4078
rect 7624 4065 7658 4078
rect 7624 3986 7658 4020
rect 7716 4177 7750 4191
rect 7716 4157 7750 4177
rect 7716 4109 7750 4118
rect 7716 4084 7750 4109
rect 7716 4041 7750 4045
rect 7716 4011 7750 4041
rect 7716 3939 7750 3972
rect 7716 3938 7750 3939
rect 6972 3888 7006 3922
rect 7058 3888 7092 3922
rect 7144 3888 7178 3922
rect 7230 3888 7264 3922
rect 7316 3888 7350 3922
rect 7402 3888 7436 3922
rect 7624 3827 7658 3850
rect 7624 3816 7658 3827
rect 7144 3732 7178 3766
rect 7222 3732 7256 3766
rect 7299 3732 7333 3766
rect 7376 3732 7410 3766
rect 7453 3732 7487 3766
rect 7530 3732 7564 3766
rect 7624 3757 7658 3775
rect 7624 3741 7658 3757
rect 7624 3687 7658 3700
rect 7624 3666 7658 3687
rect 7624 3617 7658 3625
rect 4368 3557 4379 3591
rect 4379 3557 4402 3591
rect 4440 3557 4447 3591
rect 4447 3557 4474 3591
rect 4607 3557 4641 3591
rect 4682 3557 4713 3591
rect 4713 3557 4716 3591
rect 4757 3557 4785 3591
rect 4785 3557 4791 3591
rect 4832 3557 4857 3591
rect 4857 3557 4866 3591
rect 4907 3557 4929 3591
rect 4929 3557 4941 3591
rect 4982 3557 5000 3591
rect 5000 3557 5016 3591
rect 5057 3557 5071 3591
rect 5071 3557 5091 3591
rect 5228 3557 5262 3591
rect 5320 3557 5337 3591
rect 5337 3557 5354 3591
rect 5412 3557 5443 3591
rect 5443 3557 5446 3591
rect 5503 3557 5515 3591
rect 5515 3557 5537 3591
rect 6972 3576 7006 3610
rect 7058 3576 7092 3610
rect 7144 3576 7178 3610
rect 7230 3576 7264 3610
rect 7316 3576 7350 3610
rect 7402 3576 7436 3610
rect 7624 3591 7658 3617
rect 7624 3547 7658 3550
rect 7624 3516 7658 3547
rect 7144 3420 7178 3454
rect 7222 3420 7256 3454
rect 7299 3420 7333 3454
rect 7376 3420 7410 3454
rect 7453 3420 7487 3454
rect 7530 3420 7564 3454
rect 7624 3441 7658 3475
rect 7624 3371 7658 3399
rect 7624 3365 7658 3371
rect 7624 3301 7658 3323
rect 6972 3264 7006 3298
rect 7058 3264 7092 3298
rect 7144 3264 7178 3298
rect 7230 3264 7264 3298
rect 7316 3264 7350 3298
rect 7402 3264 7436 3298
rect 7624 3289 7658 3301
rect 7624 3231 7658 3247
rect 7624 3213 7658 3231
rect 7624 3161 7658 3171
rect 7144 3108 7178 3142
rect 7222 3108 7256 3142
rect 7299 3108 7333 3142
rect 7376 3108 7410 3142
rect 7453 3108 7487 3142
rect 7530 3108 7564 3142
rect 7624 3137 7658 3161
rect 7624 3090 7658 3095
rect 7624 3061 7658 3090
rect 6972 2952 7006 2986
rect 7058 2952 7092 2986
rect 7144 2952 7178 2986
rect 7230 2952 7264 2986
rect 7316 2952 7350 2986
rect 7402 2952 7436 2986
rect 7624 2985 7658 3019
rect 7624 2914 7658 2943
rect 7624 2909 7658 2914
rect 7624 2843 7658 2867
rect 7624 2833 7658 2843
rect 7144 2796 7178 2830
rect 7227 2796 7261 2830
rect 7310 2796 7344 2830
rect 7392 2796 7426 2830
rect 7474 2796 7508 2830
rect 7624 2772 7658 2791
rect 7624 2757 7658 2772
rect 7716 3871 7750 3899
rect 7716 3865 7750 3871
rect 7716 3803 7750 3826
rect 7716 3792 7750 3803
rect 7716 3735 7750 3753
rect 7716 3719 7750 3735
rect 7716 3667 7750 3680
rect 7716 3646 7750 3667
rect 7716 3599 7750 3607
rect 7716 3573 7750 3599
rect 7716 3531 7750 3534
rect 7716 3500 7750 3531
rect 7716 3429 7750 3461
rect 7716 3427 7750 3429
rect 7716 3361 7750 3388
rect 7716 3354 7750 3361
rect 7716 3293 7750 3315
rect 7716 3281 7750 3293
rect 7716 3225 7750 3242
rect 7716 3208 7750 3225
rect 7716 3157 7750 3169
rect 7716 3135 7750 3157
rect 7716 3089 7750 3096
rect 7716 3062 7750 3089
rect 7716 3021 7750 3023
rect 7716 2989 7750 3021
rect 7716 2919 7750 2950
rect 7716 2916 7750 2919
rect 7716 2851 7750 2877
rect 7716 2843 7750 2851
rect 7716 2783 7750 2804
rect 7716 2770 7750 2783
rect 6972 2640 7006 2674
rect 7058 2640 7092 2674
rect 7144 2640 7178 2674
rect 7230 2640 7264 2674
rect 7316 2640 7350 2674
rect 7402 2640 7436 2674
rect 7625 2613 7659 2617
rect 7625 2583 7658 2613
rect 7658 2583 7659 2613
rect 7144 2484 7178 2518
rect 7222 2484 7256 2518
rect 7299 2484 7333 2518
rect 7376 2484 7410 2518
rect 7453 2484 7487 2518
rect 7530 2484 7564 2518
rect 7625 2511 7658 2523
rect 7658 2511 7659 2523
rect 7625 2489 7659 2511
rect 7076 2276 7110 2309
rect 7155 2276 7189 2309
rect 7234 2276 7268 2309
rect 7313 2276 7347 2309
rect 7392 2276 7426 2309
rect 7470 2276 7504 2309
rect 7548 2276 7582 2309
rect 7626 2276 7660 2309
rect 7704 2276 7738 2309
rect 7782 2276 7816 2309
rect 7860 2276 7894 2309
rect 7076 2275 7105 2276
rect 7105 2275 7110 2276
rect 7155 2275 7173 2276
rect 7173 2275 7189 2276
rect 7234 2275 7241 2276
rect 7241 2275 7268 2276
rect 7313 2275 7343 2276
rect 7343 2275 7347 2276
rect 7392 2275 7411 2276
rect 7411 2275 7426 2276
rect 7470 2275 7479 2276
rect 7479 2275 7504 2276
rect 7548 2275 7581 2276
rect 7581 2275 7582 2276
rect 7626 2275 7649 2276
rect 7649 2275 7660 2276
rect 7704 2275 7717 2276
rect 7717 2275 7738 2276
rect 7782 2275 7785 2276
rect 7785 2275 7816 2276
rect 7860 2275 7887 2276
rect 7887 2275 7894 2276
rect 7076 2207 7110 2231
rect 7155 2207 7189 2231
rect 7234 2207 7268 2231
rect 7313 2207 7347 2231
rect 7392 2207 7426 2231
rect 7470 2207 7504 2231
rect 7548 2207 7582 2231
rect 7626 2207 7660 2231
rect 7704 2207 7738 2231
rect 7782 2207 7816 2231
rect 7860 2207 7894 2231
rect 7076 2197 7105 2207
rect 7105 2197 7110 2207
rect 7155 2197 7173 2207
rect 7173 2197 7189 2207
rect 7234 2197 7241 2207
rect 7241 2197 7268 2207
rect 7313 2197 7343 2207
rect 7343 2197 7347 2207
rect 7392 2197 7411 2207
rect 7411 2197 7426 2207
rect 7470 2197 7479 2207
rect 7479 2197 7504 2207
rect 7548 2197 7581 2207
rect 7581 2197 7582 2207
rect 7626 2197 7649 2207
rect 7649 2197 7660 2207
rect 7704 2197 7717 2207
rect 7717 2197 7738 2207
rect 7782 2197 7785 2207
rect 7785 2197 7816 2207
rect 7860 2197 7887 2207
rect 7887 2197 7894 2207
rect 7076 2138 7110 2153
rect 7155 2138 7189 2153
rect 7234 2138 7268 2153
rect 7313 2138 7347 2153
rect 7392 2138 7426 2153
rect 7470 2138 7504 2153
rect 7548 2138 7582 2153
rect 7626 2138 7660 2153
rect 7704 2138 7738 2153
rect 7782 2138 7816 2153
rect 7860 2138 7894 2153
rect 7076 2119 7105 2138
rect 7105 2119 7110 2138
rect 7155 2119 7173 2138
rect 7173 2119 7189 2138
rect 7234 2119 7241 2138
rect 7241 2119 7268 2138
rect 7313 2119 7343 2138
rect 7343 2119 7347 2138
rect 7392 2119 7411 2138
rect 7411 2119 7426 2138
rect 7470 2119 7479 2138
rect 7479 2119 7504 2138
rect 7548 2119 7581 2138
rect 7581 2119 7582 2138
rect 7626 2119 7649 2138
rect 7649 2119 7660 2138
rect 7704 2119 7717 2138
rect 7717 2119 7738 2138
rect 7782 2119 7785 2138
rect 7785 2119 7816 2138
rect 7860 2119 7887 2138
rect 7887 2119 7894 2138
rect 7076 2068 7110 2075
rect 7155 2068 7189 2075
rect 7234 2068 7268 2075
rect 7313 2068 7347 2075
rect 7392 2068 7426 2075
rect 7470 2068 7504 2075
rect 7548 2068 7582 2075
rect 7626 2068 7660 2075
rect 7704 2068 7738 2075
rect 7782 2068 7816 2075
rect 7860 2068 7894 2075
rect 7076 2041 7105 2068
rect 7105 2041 7110 2068
rect 7155 2041 7173 2068
rect 7173 2041 7189 2068
rect 7234 2041 7241 2068
rect 7241 2041 7268 2068
rect 7313 2041 7343 2068
rect 7343 2041 7347 2068
rect 7392 2041 7411 2068
rect 7411 2041 7426 2068
rect 7470 2041 7479 2068
rect 7479 2041 7504 2068
rect 7548 2041 7581 2068
rect 7581 2041 7582 2068
rect 7626 2041 7649 2068
rect 7649 2041 7660 2068
rect 7704 2041 7717 2068
rect 7717 2041 7738 2068
rect 7782 2041 7785 2068
rect 7785 2041 7816 2068
rect 7860 2041 7887 2068
rect 7887 2041 7894 2068
rect 7076 1964 7105 1997
rect 7105 1964 7110 1997
rect 7155 1964 7173 1997
rect 7173 1964 7189 1997
rect 7234 1964 7241 1997
rect 7241 1964 7268 1997
rect 7313 1964 7343 1997
rect 7343 1964 7347 1997
rect 7392 1964 7411 1997
rect 7411 1964 7426 1997
rect 7470 1964 7479 1997
rect 7479 1964 7504 1997
rect 7548 1964 7581 1997
rect 7581 1964 7582 1997
rect 7626 1964 7649 1997
rect 7649 1964 7660 1997
rect 7704 1964 7717 1997
rect 7717 1964 7738 1997
rect 7782 1964 7785 1997
rect 7785 1964 7816 1997
rect 7860 1964 7887 1997
rect 7887 1964 7894 1997
rect 7076 1963 7110 1964
rect 7155 1963 7189 1964
rect 7234 1963 7268 1964
rect 7313 1963 7347 1964
rect 7392 1963 7426 1964
rect 7470 1963 7504 1964
rect 7548 1963 7582 1964
rect 7626 1963 7660 1964
rect 7704 1963 7738 1964
rect 7782 1963 7816 1964
rect 7860 1963 7894 1964
rect 7076 1894 7105 1919
rect 7105 1894 7110 1919
rect 7155 1894 7173 1919
rect 7173 1894 7189 1919
rect 7234 1894 7241 1919
rect 7241 1894 7268 1919
rect 7313 1894 7343 1919
rect 7343 1894 7347 1919
rect 7392 1894 7411 1919
rect 7411 1894 7426 1919
rect 7470 1894 7479 1919
rect 7479 1894 7504 1919
rect 7548 1894 7581 1919
rect 7581 1894 7582 1919
rect 7626 1894 7649 1919
rect 7649 1894 7660 1919
rect 7704 1894 7717 1919
rect 7717 1894 7738 1919
rect 7782 1894 7785 1919
rect 7785 1894 7816 1919
rect 7860 1894 7887 1919
rect 7887 1894 7894 1919
rect 7076 1885 7110 1894
rect 7155 1885 7189 1894
rect 7234 1885 7268 1894
rect 7313 1885 7347 1894
rect 7392 1885 7426 1894
rect 7470 1885 7504 1894
rect 7548 1885 7582 1894
rect 7626 1885 7660 1894
rect 7704 1885 7738 1894
rect 7782 1885 7816 1894
rect 7860 1885 7894 1894
rect 7076 1824 7105 1841
rect 7105 1824 7110 1841
rect 7155 1824 7173 1841
rect 7173 1824 7189 1841
rect 7234 1824 7241 1841
rect 7241 1824 7268 1841
rect 7313 1824 7343 1841
rect 7343 1824 7347 1841
rect 7392 1824 7411 1841
rect 7411 1824 7426 1841
rect 7470 1824 7479 1841
rect 7479 1824 7504 1841
rect 7548 1824 7581 1841
rect 7581 1824 7582 1841
rect 7626 1824 7649 1841
rect 7649 1824 7660 1841
rect 7704 1824 7717 1841
rect 7717 1824 7738 1841
rect 7782 1824 7785 1841
rect 7785 1824 7816 1841
rect 7860 1824 7887 1841
rect 7887 1824 7894 1841
rect 7076 1807 7110 1824
rect 7155 1807 7189 1824
rect 7234 1807 7268 1824
rect 7313 1807 7347 1824
rect 7392 1807 7426 1824
rect 7470 1807 7504 1824
rect 7548 1807 7582 1824
rect 7626 1807 7660 1824
rect 7704 1807 7738 1824
rect 7782 1807 7816 1824
rect 7860 1807 7894 1824
rect 7049 1544 7071 1545
rect 7071 1544 7083 1545
rect 7121 1544 7139 1545
rect 7139 1544 7155 1545
rect 7193 1544 7207 1545
rect 7207 1544 7227 1545
rect 7265 1544 7275 1545
rect 7275 1544 7299 1545
rect 7337 1544 7343 1545
rect 7343 1544 7371 1545
rect 7409 1544 7411 1545
rect 7411 1544 7443 1545
rect 7481 1544 7513 1545
rect 7513 1544 7515 1545
rect 7553 1544 7581 1545
rect 7581 1544 7587 1545
rect 7625 1544 7649 1545
rect 7649 1544 7659 1545
rect 7697 1544 7717 1545
rect 7717 1544 7731 1545
rect 7769 1544 7785 1545
rect 7785 1544 7803 1545
rect 7841 1544 7853 1545
rect 7853 1544 7875 1545
rect 7049 1511 7083 1544
rect 7121 1511 7155 1544
rect 7193 1511 7227 1544
rect 7265 1511 7299 1544
rect 7337 1511 7371 1544
rect 7409 1511 7443 1544
rect 7481 1511 7515 1544
rect 7553 1511 7587 1544
rect 7625 1511 7659 1544
rect 7697 1511 7731 1544
rect 7769 1511 7803 1544
rect 7841 1511 7875 1544
rect 7049 1438 7083 1472
rect 7121 1438 7155 1472
rect 7193 1438 7227 1472
rect 7265 1438 7299 1472
rect 7337 1438 7371 1472
rect 7409 1438 7443 1472
rect 7481 1438 7515 1472
rect 7553 1438 7587 1472
rect 7625 1438 7659 1472
rect 7697 1438 7731 1472
rect 7769 1438 7803 1472
rect 7841 1438 7875 1472
rect 7049 1368 7083 1399
rect 7121 1368 7155 1399
rect 7193 1368 7227 1399
rect 7265 1368 7299 1399
rect 7337 1368 7371 1399
rect 7409 1368 7443 1399
rect 7481 1368 7515 1399
rect 7553 1368 7587 1399
rect 7625 1368 7659 1399
rect 7697 1368 7731 1399
rect 7769 1368 7803 1399
rect 7841 1368 7875 1399
rect 7049 1365 7071 1368
rect 7071 1365 7083 1368
rect 7121 1365 7139 1368
rect 7139 1365 7155 1368
rect 7193 1365 7207 1368
rect 7207 1365 7227 1368
rect 7265 1365 7275 1368
rect 7275 1365 7299 1368
rect 7337 1365 7343 1368
rect 7343 1365 7371 1368
rect 7409 1365 7411 1368
rect 7411 1365 7443 1368
rect 7481 1365 7513 1368
rect 7513 1365 7515 1368
rect 7553 1365 7581 1368
rect 7581 1365 7587 1368
rect 7625 1365 7649 1368
rect 7649 1365 7659 1368
rect 7697 1365 7717 1368
rect 7717 1365 7731 1368
rect 7769 1365 7785 1368
rect 7785 1365 7803 1368
rect 7841 1365 7853 1368
rect 7853 1365 7875 1368
rect 7049 1298 7083 1326
rect 7121 1298 7155 1326
rect 7193 1298 7227 1326
rect 7265 1298 7299 1326
rect 7337 1298 7371 1326
rect 7409 1298 7443 1326
rect 7481 1298 7515 1326
rect 7553 1298 7587 1326
rect 7625 1298 7659 1326
rect 7697 1298 7731 1326
rect 7769 1298 7803 1326
rect 7841 1298 7875 1326
rect 7049 1292 7071 1298
rect 7071 1292 7083 1298
rect 7121 1292 7139 1298
rect 7139 1292 7155 1298
rect 7193 1292 7207 1298
rect 7207 1292 7227 1298
rect 7265 1292 7275 1298
rect 7275 1292 7299 1298
rect 7337 1292 7343 1298
rect 7343 1292 7371 1298
rect 7409 1292 7411 1298
rect 7411 1292 7443 1298
rect 7481 1292 7513 1298
rect 7513 1292 7515 1298
rect 7553 1292 7581 1298
rect 7581 1292 7587 1298
rect 7625 1292 7649 1298
rect 7649 1292 7659 1298
rect 7697 1292 7717 1298
rect 7717 1292 7731 1298
rect 7769 1292 7785 1298
rect 7785 1292 7803 1298
rect 7841 1292 7853 1298
rect 7853 1292 7875 1298
rect 7049 1228 7083 1253
rect 7121 1228 7155 1253
rect 7193 1228 7227 1253
rect 7265 1228 7299 1253
rect 7337 1228 7371 1253
rect 7409 1228 7443 1253
rect 7481 1228 7515 1253
rect 7553 1228 7587 1253
rect 7625 1228 7659 1253
rect 7697 1228 7731 1253
rect 7769 1228 7803 1253
rect 7841 1228 7875 1253
rect 7049 1219 7071 1228
rect 7071 1219 7083 1228
rect 7121 1219 7139 1228
rect 7139 1219 7155 1228
rect 7193 1219 7207 1228
rect 7207 1219 7227 1228
rect 7265 1219 7275 1228
rect 7275 1219 7299 1228
rect 7337 1219 7343 1228
rect 7343 1219 7371 1228
rect 7409 1219 7411 1228
rect 7411 1219 7443 1228
rect 7481 1219 7513 1228
rect 7513 1219 7515 1228
rect 7553 1219 7581 1228
rect 7581 1219 7587 1228
rect 7625 1219 7649 1228
rect 7649 1219 7659 1228
rect 7697 1219 7717 1228
rect 7717 1219 7731 1228
rect 7769 1219 7785 1228
rect 7785 1219 7803 1228
rect 7841 1219 7853 1228
rect 7853 1219 7875 1228
rect 7049 1158 7083 1180
rect 7121 1158 7155 1180
rect 7193 1158 7227 1180
rect 7265 1158 7299 1180
rect 7337 1158 7371 1180
rect 7409 1158 7443 1180
rect 7481 1158 7515 1180
rect 7553 1158 7587 1180
rect 7625 1158 7659 1180
rect 7697 1158 7731 1180
rect 7769 1158 7803 1180
rect 7841 1158 7875 1180
rect 7049 1146 7071 1158
rect 7071 1146 7083 1158
rect 7121 1146 7139 1158
rect 7139 1146 7155 1158
rect 7193 1146 7207 1158
rect 7207 1146 7227 1158
rect 7265 1146 7275 1158
rect 7275 1146 7299 1158
rect 7337 1146 7343 1158
rect 7343 1146 7371 1158
rect 7409 1146 7411 1158
rect 7411 1146 7443 1158
rect 7481 1146 7513 1158
rect 7513 1146 7515 1158
rect 7553 1146 7581 1158
rect 7581 1146 7587 1158
rect 7625 1146 7649 1158
rect 7649 1146 7659 1158
rect 7697 1146 7717 1158
rect 7717 1146 7731 1158
rect 7769 1146 7785 1158
rect 7785 1146 7803 1158
rect 7841 1146 7853 1158
rect 7853 1146 7875 1158
rect 7049 1088 7083 1107
rect 7121 1088 7155 1107
rect 7193 1088 7227 1107
rect 7265 1088 7299 1107
rect 7337 1088 7371 1107
rect 7409 1088 7443 1107
rect 7481 1088 7515 1107
rect 7553 1088 7587 1107
rect 7625 1088 7659 1107
rect 7697 1088 7731 1107
rect 7769 1088 7803 1107
rect 7841 1088 7875 1107
rect 7049 1073 7071 1088
rect 7071 1073 7083 1088
rect 7121 1073 7139 1088
rect 7139 1073 7155 1088
rect 7193 1073 7207 1088
rect 7207 1073 7227 1088
rect 7265 1073 7275 1088
rect 7275 1073 7299 1088
rect 7337 1073 7343 1088
rect 7343 1073 7371 1088
rect 7409 1073 7411 1088
rect 7411 1073 7443 1088
rect 7481 1073 7513 1088
rect 7513 1073 7515 1088
rect 7553 1073 7581 1088
rect 7581 1073 7587 1088
rect 7625 1073 7649 1088
rect 7649 1073 7659 1088
rect 7697 1073 7717 1088
rect 7717 1073 7731 1088
rect 7769 1073 7785 1088
rect 7785 1073 7803 1088
rect 7841 1073 7853 1088
rect 7853 1073 7875 1088
rect 7049 1018 7083 1034
rect 7121 1018 7155 1034
rect 7193 1018 7227 1034
rect 7265 1018 7299 1034
rect 7337 1018 7371 1034
rect 7409 1018 7443 1034
rect 7481 1018 7515 1034
rect 7553 1018 7587 1034
rect 7625 1018 7659 1034
rect 7697 1018 7731 1034
rect 7769 1018 7803 1034
rect 7841 1018 7875 1034
rect 7049 1000 7071 1018
rect 7071 1000 7083 1018
rect 7121 1000 7139 1018
rect 7139 1000 7155 1018
rect 7193 1000 7207 1018
rect 7207 1000 7227 1018
rect 7265 1000 7275 1018
rect 7275 1000 7299 1018
rect 7337 1000 7343 1018
rect 7343 1000 7371 1018
rect 7409 1000 7411 1018
rect 7411 1000 7443 1018
rect 7481 1000 7513 1018
rect 7513 1000 7515 1018
rect 7553 1000 7581 1018
rect 7581 1000 7587 1018
rect 7625 1000 7649 1018
rect 7649 1000 7659 1018
rect 7697 1000 7717 1018
rect 7717 1000 7731 1018
rect 7769 1000 7785 1018
rect 7785 1000 7803 1018
rect 7841 1000 7853 1018
rect 7853 1000 7875 1018
rect 7049 948 7083 961
rect 7121 948 7155 961
rect 7193 948 7227 961
rect 7265 948 7299 961
rect 7337 948 7371 961
rect 7409 948 7443 961
rect 7481 948 7515 961
rect 7553 948 7587 961
rect 7625 948 7659 961
rect 7697 948 7731 961
rect 7769 948 7803 961
rect 7841 948 7875 961
rect 7049 927 7071 948
rect 7071 927 7083 948
rect 7121 927 7139 948
rect 7139 927 7155 948
rect 7193 927 7207 948
rect 7207 927 7227 948
rect 7265 927 7275 948
rect 7275 927 7299 948
rect 7337 927 7343 948
rect 7343 927 7371 948
rect 7409 927 7411 948
rect 7411 927 7443 948
rect 7481 927 7513 948
rect 7513 927 7515 948
rect 7553 927 7581 948
rect 7581 927 7587 948
rect 7625 927 7649 948
rect 7649 927 7659 948
rect 7697 927 7717 948
rect 7717 927 7731 948
rect 7769 927 7785 948
rect 7785 927 7803 948
rect 7841 927 7853 948
rect 7853 927 7875 948
rect 7049 878 7083 888
rect 7121 878 7155 888
rect 7193 878 7227 888
rect 7265 878 7299 888
rect 7337 878 7371 888
rect 7409 878 7443 888
rect 7481 878 7515 888
rect 7553 878 7587 888
rect 7625 878 7659 888
rect 7697 878 7731 888
rect 7769 878 7803 888
rect 7841 878 7875 888
rect 7049 854 7071 878
rect 7071 854 7083 878
rect 7121 854 7139 878
rect 7139 854 7155 878
rect 7193 854 7207 878
rect 7207 854 7227 878
rect 7265 854 7275 878
rect 7275 854 7299 878
rect 7337 854 7343 878
rect 7343 854 7371 878
rect 7409 854 7411 878
rect 7411 854 7443 878
rect 7481 854 7513 878
rect 7513 854 7515 878
rect 7553 854 7581 878
rect 7581 854 7587 878
rect 7625 854 7649 878
rect 7649 854 7659 878
rect 7697 854 7717 878
rect 7717 854 7731 878
rect 7769 854 7785 878
rect 7785 854 7803 878
rect 7841 854 7853 878
rect 7853 854 7875 878
rect 7049 808 7083 814
rect 7121 808 7155 814
rect 7193 808 7227 814
rect 7265 808 7299 814
rect 7337 808 7371 814
rect 7409 808 7443 814
rect 7481 808 7515 814
rect 7553 808 7587 814
rect 7625 808 7659 814
rect 7697 808 7731 814
rect 7769 808 7803 814
rect 7841 808 7875 814
rect 7049 780 7071 808
rect 7071 780 7083 808
rect 7121 780 7139 808
rect 7139 780 7155 808
rect 7193 780 7207 808
rect 7207 780 7227 808
rect 7265 780 7275 808
rect 7275 780 7299 808
rect 7337 780 7343 808
rect 7343 780 7371 808
rect 7409 780 7411 808
rect 7411 780 7443 808
rect 7481 780 7513 808
rect 7513 780 7515 808
rect 7553 780 7581 808
rect 7581 780 7587 808
rect 7625 780 7649 808
rect 7649 780 7659 808
rect 7697 780 7717 808
rect 7717 780 7731 808
rect 7769 780 7785 808
rect 7785 780 7803 808
rect 7841 780 7853 808
rect 7853 780 7875 808
rect 7049 738 7083 740
rect 7121 738 7155 740
rect 7193 738 7227 740
rect 7265 738 7299 740
rect 7337 738 7371 740
rect 7409 738 7443 740
rect 7481 738 7515 740
rect 7553 738 7587 740
rect 7625 738 7659 740
rect 7697 738 7731 740
rect 7769 738 7803 740
rect 7841 738 7875 740
rect 7049 706 7071 738
rect 7071 706 7083 738
rect 7121 706 7139 738
rect 7139 706 7155 738
rect 7193 706 7207 738
rect 7207 706 7227 738
rect 7265 706 7275 738
rect 7275 706 7299 738
rect 7337 706 7343 738
rect 7343 706 7371 738
rect 7409 706 7411 738
rect 7411 706 7443 738
rect 7481 706 7513 738
rect 7513 706 7515 738
rect 7553 706 7581 738
rect 7581 706 7587 738
rect 7625 706 7649 738
rect 7649 706 7659 738
rect 7697 706 7717 738
rect 7717 706 7731 738
rect 7769 706 7785 738
rect 7785 706 7803 738
rect 7841 706 7853 738
rect 7853 706 7875 738
rect 7049 634 7071 666
rect 7071 634 7083 666
rect 7121 634 7139 666
rect 7139 634 7155 666
rect 7193 634 7207 666
rect 7207 634 7227 666
rect 7265 634 7275 666
rect 7275 634 7299 666
rect 7337 634 7343 666
rect 7343 634 7371 666
rect 7409 634 7411 666
rect 7411 634 7443 666
rect 7481 634 7513 666
rect 7513 634 7515 666
rect 7553 634 7581 666
rect 7581 634 7587 666
rect 7625 634 7649 666
rect 7649 634 7659 666
rect 7697 634 7717 666
rect 7717 634 7731 666
rect 7769 634 7785 666
rect 7785 634 7803 666
rect 7841 634 7853 666
rect 7853 634 7875 666
rect 7049 632 7083 634
rect 7121 632 7155 634
rect 7193 632 7227 634
rect 7265 632 7299 634
rect 7337 632 7371 634
rect 7409 632 7443 634
rect 7481 632 7515 634
rect 7553 632 7587 634
rect 7625 632 7659 634
rect 7697 632 7731 634
rect 7769 632 7803 634
rect 7841 632 7875 634
rect 7049 564 7071 592
rect 7071 564 7083 592
rect 7121 564 7139 592
rect 7139 564 7155 592
rect 7193 564 7207 592
rect 7207 564 7227 592
rect 7265 564 7275 592
rect 7275 564 7299 592
rect 7337 564 7343 592
rect 7343 564 7371 592
rect 7409 564 7411 592
rect 7411 564 7443 592
rect 7481 564 7513 592
rect 7513 564 7515 592
rect 7553 564 7581 592
rect 7581 564 7587 592
rect 7625 564 7649 592
rect 7649 564 7659 592
rect 7697 564 7717 592
rect 7717 564 7731 592
rect 7769 564 7785 592
rect 7785 564 7803 592
rect 7841 564 7853 592
rect 7853 564 7875 592
rect 7049 558 7083 564
rect 7121 558 7155 564
rect 7193 558 7227 564
rect 7265 558 7299 564
rect 7337 558 7371 564
rect 7409 558 7443 564
rect 7481 558 7515 564
rect 7553 558 7587 564
rect 7625 558 7659 564
rect 7697 558 7731 564
rect 7769 558 7803 564
rect 7841 558 7875 564
rect 7049 494 7071 518
rect 7071 494 7083 518
rect 7121 494 7139 518
rect 7139 494 7155 518
rect 7193 494 7207 518
rect 7207 494 7227 518
rect 7265 494 7275 518
rect 7275 494 7299 518
rect 7337 494 7343 518
rect 7343 494 7371 518
rect 7409 494 7411 518
rect 7411 494 7443 518
rect 7481 494 7513 518
rect 7513 494 7515 518
rect 7553 494 7581 518
rect 7581 494 7587 518
rect 7625 494 7649 518
rect 7649 494 7659 518
rect 7697 494 7717 518
rect 7717 494 7731 518
rect 7769 494 7785 518
rect 7785 494 7803 518
rect 7841 494 7853 518
rect 7853 494 7875 518
rect 7049 484 7083 494
rect 7121 484 7155 494
rect 7193 484 7227 494
rect 7265 484 7299 494
rect 7337 484 7371 494
rect 7409 484 7443 494
rect 7481 484 7515 494
rect 7553 484 7587 494
rect 7625 484 7659 494
rect 7697 484 7731 494
rect 7769 484 7803 494
rect 7841 484 7875 494
rect 7049 424 7071 444
rect 7071 424 7083 444
rect 7121 424 7139 444
rect 7139 424 7155 444
rect 7193 424 7207 444
rect 7207 424 7227 444
rect 7265 424 7275 444
rect 7275 424 7299 444
rect 7337 424 7343 444
rect 7343 424 7371 444
rect 7409 424 7411 444
rect 7411 424 7443 444
rect 7481 424 7513 444
rect 7513 424 7515 444
rect 7553 424 7581 444
rect 7581 424 7587 444
rect 7625 424 7649 444
rect 7649 424 7659 444
rect 7697 424 7717 444
rect 7717 424 7731 444
rect 7769 424 7785 444
rect 7785 424 7803 444
rect 7841 424 7853 444
rect 7853 424 7875 444
rect 7049 410 7083 424
rect 7121 410 7155 424
rect 7193 410 7227 424
rect 7265 410 7299 424
rect 7337 410 7371 424
rect 7409 410 7443 424
rect 7481 410 7515 424
rect 7553 410 7587 424
rect 7625 410 7659 424
rect 7697 410 7731 424
rect 7769 410 7803 424
rect 7841 410 7875 424
rect 7049 354 7071 370
rect 7071 354 7083 370
rect 7121 354 7139 370
rect 7139 354 7155 370
rect 7193 354 7207 370
rect 7207 354 7227 370
rect 7265 354 7275 370
rect 7275 354 7299 370
rect 7337 354 7343 370
rect 7343 354 7371 370
rect 7409 354 7411 370
rect 7411 354 7443 370
rect 7481 354 7513 370
rect 7513 354 7515 370
rect 7553 354 7581 370
rect 7581 354 7587 370
rect 7625 354 7649 370
rect 7649 354 7659 370
rect 7697 354 7717 370
rect 7717 354 7731 370
rect 7769 354 7785 370
rect 7785 354 7803 370
rect 7841 354 7853 370
rect 7853 354 7875 370
rect 7049 336 7083 354
rect 7121 336 7155 354
rect 7193 336 7227 354
rect 7265 336 7299 354
rect 7337 336 7371 354
rect 7409 336 7443 354
rect 7481 336 7515 354
rect 7553 336 7587 354
rect 7625 336 7659 354
rect 7697 336 7731 354
rect 7769 336 7803 354
rect 7841 336 7875 354
rect 7049 284 7071 296
rect 7071 284 7083 296
rect 7121 284 7139 296
rect 7139 284 7155 296
rect 7193 284 7207 296
rect 7207 284 7227 296
rect 7265 284 7275 296
rect 7275 284 7299 296
rect 7337 284 7343 296
rect 7343 284 7371 296
rect 7409 284 7411 296
rect 7411 284 7443 296
rect 7481 284 7513 296
rect 7513 284 7515 296
rect 7553 284 7581 296
rect 7581 284 7587 296
rect 7625 284 7649 296
rect 7649 284 7659 296
rect 7697 284 7717 296
rect 7717 284 7731 296
rect 7769 284 7785 296
rect 7785 284 7803 296
rect 7841 284 7853 296
rect 7853 284 7875 296
rect 7049 262 7083 284
rect 7121 262 7155 284
rect 7193 262 7227 284
rect 7265 262 7299 284
rect 7337 262 7371 284
rect 7409 262 7443 284
rect 7481 262 7515 284
rect 7553 262 7587 284
rect 7625 262 7659 284
rect 7697 262 7731 284
rect 7769 262 7803 284
rect 7841 262 7875 284
rect 7049 214 7071 222
rect 7071 214 7083 222
rect 7121 214 7139 222
rect 7139 214 7155 222
rect 7193 214 7207 222
rect 7207 214 7227 222
rect 7265 214 7275 222
rect 7275 214 7299 222
rect 7337 214 7343 222
rect 7343 214 7371 222
rect 7409 214 7411 222
rect 7411 214 7443 222
rect 7481 214 7513 222
rect 7513 214 7515 222
rect 7553 214 7581 222
rect 7581 214 7587 222
rect 7625 214 7649 222
rect 7649 214 7659 222
rect 7697 214 7717 222
rect 7717 214 7731 222
rect 7769 214 7785 222
rect 7785 214 7803 222
rect 7841 214 7853 222
rect 7853 214 7875 222
rect 7049 188 7083 214
rect 7121 188 7155 214
rect 7193 188 7227 214
rect 7265 188 7299 214
rect 7337 188 7371 214
rect 7409 188 7443 214
rect 7481 188 7515 214
rect 7553 188 7587 214
rect 7625 188 7659 214
rect 7697 188 7731 214
rect 7769 188 7803 214
rect 7841 188 7875 214
rect 7049 144 7071 148
rect 7071 144 7083 148
rect 7121 144 7139 148
rect 7139 144 7155 148
rect 7193 144 7207 148
rect 7207 144 7227 148
rect 7265 144 7275 148
rect 7275 144 7299 148
rect 7337 144 7343 148
rect 7343 144 7371 148
rect 7409 144 7411 148
rect 7411 144 7443 148
rect 7481 144 7513 148
rect 7513 144 7515 148
rect 7553 144 7581 148
rect 7581 144 7587 148
rect 7625 144 7649 148
rect 7649 144 7659 148
rect 7697 144 7717 148
rect 7717 144 7731 148
rect 7769 144 7785 148
rect 7785 144 7803 148
rect 7841 144 7853 148
rect 7853 144 7875 148
rect 7049 114 7083 144
rect 7121 114 7155 144
rect 7193 114 7227 144
rect 7265 114 7299 144
rect 7337 114 7371 144
rect 7409 114 7443 144
rect 7481 114 7515 144
rect 7553 114 7587 144
rect 7625 114 7659 144
rect 7697 114 7731 144
rect 7769 114 7803 144
rect 7841 114 7875 144
rect 7049 40 7083 74
rect 7121 40 7155 74
rect 7193 40 7227 74
rect 7265 40 7299 74
rect 7337 40 7371 74
rect 7409 40 7443 74
rect 7481 40 7515 74
rect 7553 40 7587 74
rect 7625 40 7659 74
rect 7697 40 7731 74
rect 7769 40 7803 74
rect 7841 40 7875 74
<< metal1 >>
tri 2862 39800 2896 39834 nw
tri 7706 39800 7740 39834 ne
tri 9712 39776 9713 39777 ne
rect 9713 39776 9746 39777
rect 484 39743 485 39776
tri 485 39743 518 39776 nw
tri 2447 39743 2480 39776 ne
rect 2480 39743 2481 39776
tri 9713 39743 9746 39776 ne
tri 9792 39743 9826 39777 nw
tri 484 39742 485 39743 nw
tri 2480 39742 2481 39743 ne
tri 628 39475 662 39509 nw
rect 3122 39452 5447 39574
tri 5447 39540 5481 39574 nw
tri 5600 39540 5634 39574 ne
tri 3122 39418 3156 39452 nw
tri 4289 39418 4323 39452 ne
rect 3165 30425 3217 39365
tri 4289 39042 4323 39076 se
tri 4289 38962 4323 38996 ne
tri 4289 38586 4323 38620 se
tri 4289 38506 4323 38540 ne
tri 4289 38130 4323 38164 se
tri 4289 38050 4323 38084 ne
tri 4289 37674 4323 37708 se
tri 4289 37594 4323 37628 ne
tri 4289 37218 4323 37252 se
tri 4289 37138 4323 37172 ne
tri 4289 36762 4323 36796 se
tri 4289 36682 4323 36716 ne
tri 4289 36306 4323 36340 se
tri 4289 36226 4323 36260 ne
tri 4289 35850 4323 35884 se
tri 4289 35770 4323 35804 ne
tri 4289 35394 4323 35428 se
tri 4289 35314 4323 35348 ne
tri 4289 34938 4323 34972 se
tri 4289 34858 4323 34892 ne
tri 4289 34482 4323 34516 se
tri 4289 34402 4323 34436 ne
tri 4289 34026 4323 34060 se
tri 4289 33946 4323 33980 ne
tri 4289 33570 4323 33604 se
tri 4289 33490 4323 33524 ne
tri 4289 33114 4323 33148 se
tri 4289 33034 4323 33068 ne
tri 4289 32658 4323 32692 se
tri 4289 32578 4323 32612 ne
tri 4289 32202 4323 32236 se
tri 4289 32122 4323 32156 ne
tri 4289 31746 4323 31780 se
tri 4289 31666 4323 31700 ne
tri 4289 31290 4323 31324 se
tri 4289 31210 4323 31244 ne
tri 4289 30834 4323 30868 se
tri 4289 30754 4323 30788 ne
tri 4289 30378 4323 30412 se
rect 4323 30332 5447 39452
rect 8481 30284 8488 30336
rect 8540 30284 8552 30336
rect 8604 30284 8610 30336
rect 8481 30134 8610 30284
tri 4860 30131 4863 30134 se
tri 4860 30082 4863 30085 ne
rect 8481 30082 8487 30134
rect 8539 30082 8551 30134
rect 8603 30082 8610 30134
rect 3550 29896 3602 30057
rect 5261 29899 5313 30057
rect 8481 30054 8610 30082
rect 8481 30002 8487 30054
rect 8539 30002 8551 30054
rect 8603 30002 8610 30054
rect 8481 29974 8610 30002
rect 8481 29922 8487 29974
rect 8539 29922 8551 29974
rect 8603 29922 8610 29974
rect 8481 29894 8610 29922
rect 8481 29842 8487 29894
rect 8539 29842 8551 29894
rect 8603 29842 8610 29894
rect 8481 29814 8610 29842
rect 8481 29762 8487 29814
rect 8539 29762 8551 29814
rect 8603 29762 8610 29814
rect 8481 29699 8610 29762
rect 8481 29647 8487 29699
rect 8539 29647 8551 29699
rect 8603 29647 8610 29699
rect 3550 29481 3602 29633
rect 5261 29465 5313 29633
rect 8481 29460 8610 29647
rect 8481 29408 8488 29460
rect 8540 29408 8552 29460
rect 8604 29408 8610 29460
rect 8481 29406 8610 29408
tri 4375 29195 4409 29229 ne
tri 4455 29195 4489 29229 nw
rect 3703 29095 4376 29147
rect 4503 29095 5235 29147
rect 3550 28913 3602 29073
tri 4374 29009 4409 29044 se
tri 4455 29009 4489 29043 sw
tri 4374 28923 4408 28957 ne
rect 4408 28923 4409 28957
tri 4455 28923 4489 28957 nw
tri 4408 28922 4409 28923 ne
rect 5261 28913 5313 29073
tri 3122 28443 3156 28477 sw
tri 5600 28443 5634 28477 se
rect 3076 28391 5680 28443
tri 2862 28183 2896 28217 sw
rect 2816 28131 5940 28183
tri 9792 28008 9812 28028 sw
tri 9732 27994 9746 28008 se
rect 9792 27994 9812 28008
tri 9812 27994 9826 28008 sw
rect 366 27988 484 27994
rect 418 27936 432 27988
rect 366 27921 484 27936
rect 418 27869 432 27921
rect 366 27854 484 27869
rect 418 27802 432 27854
rect 366 27787 484 27802
rect 418 27735 432 27787
rect 366 27720 484 27735
rect 418 27668 432 27720
rect 366 27653 484 27668
rect 418 27601 432 27653
rect 366 27586 484 27601
rect 418 27534 432 27586
rect 366 27519 484 27534
rect 418 27467 432 27519
rect 366 27452 484 27467
rect 418 27400 432 27452
rect 366 27394 484 27400
rect 2481 27988 2599 27994
rect 2533 27936 2547 27988
rect 9732 27988 9862 27994
rect 2481 27921 2599 27936
rect 2533 27869 2547 27921
tri 7960 27913 7994 27947 se
rect 2481 27854 2599 27869
rect 2533 27802 2547 27854
rect 2481 27787 2599 27802
rect 2533 27735 2547 27787
rect 2481 27720 2599 27735
rect 2533 27668 2547 27720
rect 2481 27653 2599 27668
rect 2533 27601 2547 27653
rect 2481 27586 2599 27601
rect 2533 27534 2547 27586
rect 2481 27519 2599 27534
rect 2533 27467 2547 27519
rect 2481 27452 2599 27467
rect 2872 27912 7994 27913
rect 2872 27860 2878 27912
rect 2930 27903 3008 27912
rect 3060 27903 3138 27912
rect 3190 27903 3268 27912
rect 3320 27903 3398 27912
rect 3450 27903 3528 27912
rect 3580 27903 3658 27912
rect 3710 27903 3788 27912
rect 3840 27903 3918 27912
rect 3970 27903 4048 27912
rect 4100 27903 4178 27912
rect 4230 27903 4308 27912
rect 4360 27903 4438 27912
rect 4490 27903 4568 27912
rect 4620 27903 4698 27912
rect 4750 27903 4828 27912
rect 4880 27903 4958 27912
rect 5010 27903 5088 27912
rect 5140 27903 5218 27912
rect 5270 27903 5348 27912
rect 5400 27903 5478 27912
rect 5530 27903 5608 27912
rect 5660 27903 5738 27912
rect 5790 27903 5868 27912
rect 5920 27903 5998 27912
rect 6050 27903 6128 27912
rect 2930 27869 2957 27903
rect 2991 27869 3008 27903
rect 3064 27869 3103 27903
rect 3137 27869 3138 27903
rect 3210 27869 3249 27903
rect 3320 27869 3322 27903
rect 3356 27869 3395 27903
rect 3450 27869 3468 27903
rect 3502 27869 3528 27903
rect 3580 27869 3614 27903
rect 3648 27869 3658 27903
rect 3721 27869 3760 27903
rect 3867 27869 3906 27903
rect 3970 27869 3979 27903
rect 4013 27869 4048 27903
rect 4100 27869 4125 27903
rect 4159 27869 4178 27903
rect 4232 27869 4271 27903
rect 4305 27869 4308 27903
rect 4378 27869 4417 27903
rect 4524 27869 4563 27903
rect 4620 27869 4636 27903
rect 4670 27869 4698 27903
rect 4750 27869 4782 27903
rect 4816 27869 4828 27903
rect 4889 27869 4928 27903
rect 5035 27869 5074 27903
rect 5140 27869 5147 27903
rect 5181 27869 5218 27903
rect 5270 27869 5293 27903
rect 5327 27869 5348 27903
rect 5400 27869 5439 27903
rect 5473 27869 5478 27903
rect 5546 27869 5585 27903
rect 5692 27869 5731 27903
rect 5790 27869 5804 27903
rect 5838 27869 5868 27903
rect 5920 27869 5950 27903
rect 5984 27869 5998 27903
rect 6057 27869 6128 27903
rect 2930 27860 3008 27869
rect 3060 27860 3138 27869
rect 3190 27860 3268 27869
rect 3320 27860 3398 27869
rect 3450 27860 3528 27869
rect 3580 27860 3658 27869
rect 3710 27860 3788 27869
rect 3840 27860 3918 27869
rect 3970 27860 4048 27869
rect 4100 27860 4178 27869
rect 4230 27860 4308 27869
rect 4360 27860 4438 27869
rect 4490 27860 4568 27869
rect 4620 27860 4698 27869
rect 4750 27860 4828 27869
rect 4880 27860 4958 27869
rect 5010 27860 5088 27869
rect 5140 27860 5218 27869
rect 5270 27860 5348 27869
rect 5400 27860 5478 27869
rect 5530 27860 5608 27869
rect 5660 27860 5738 27869
rect 5790 27860 5868 27869
rect 5920 27860 5998 27869
rect 6050 27860 6128 27869
rect 6180 27860 6258 27912
rect 6310 27860 6388 27912
rect 6440 27860 6517 27912
rect 6569 27860 6646 27912
rect 6698 27860 6775 27912
rect 6827 27860 6904 27912
rect 6956 27860 7033 27912
rect 7085 27860 7162 27912
rect 7214 27860 7291 27912
rect 7343 27860 7420 27912
rect 7472 27860 7549 27912
rect 7601 27860 7678 27912
rect 7730 27860 7807 27912
rect 7859 27860 7936 27912
rect 7988 27860 7994 27912
rect 2872 27832 7994 27860
rect 2872 27780 2878 27832
rect 2930 27823 3008 27832
rect 3060 27823 3138 27832
rect 3190 27823 3268 27832
rect 3320 27823 3398 27832
rect 3450 27823 3528 27832
rect 3580 27823 3658 27832
rect 3710 27823 3788 27832
rect 3840 27823 3918 27832
rect 3970 27823 4048 27832
rect 4100 27823 4178 27832
rect 4230 27823 4308 27832
rect 4360 27823 4438 27832
rect 4490 27823 4568 27832
rect 4620 27823 4698 27832
rect 4750 27823 4828 27832
rect 4880 27823 4958 27832
rect 5010 27823 5088 27832
rect 5140 27823 5218 27832
rect 5270 27823 5348 27832
rect 5400 27823 5478 27832
rect 5530 27823 5608 27832
rect 5660 27823 5738 27832
rect 5790 27823 5868 27832
rect 5920 27823 5998 27832
rect 6050 27823 6128 27832
rect 2930 27789 2957 27823
rect 2991 27789 3008 27823
rect 3064 27789 3103 27823
rect 3137 27789 3138 27823
rect 3210 27789 3249 27823
rect 3320 27789 3322 27823
rect 3356 27789 3395 27823
rect 3450 27789 3468 27823
rect 3502 27789 3528 27823
rect 3580 27789 3614 27823
rect 3648 27789 3658 27823
rect 3721 27789 3760 27823
rect 3867 27789 3906 27823
rect 3970 27789 3979 27823
rect 4013 27789 4048 27823
rect 4100 27789 4125 27823
rect 4159 27789 4178 27823
rect 4232 27789 4271 27823
rect 4305 27789 4308 27823
rect 4378 27789 4417 27823
rect 4524 27789 4563 27823
rect 4620 27789 4636 27823
rect 4670 27789 4698 27823
rect 4750 27789 4782 27823
rect 4816 27789 4828 27823
rect 4889 27789 4928 27823
rect 5035 27789 5074 27823
rect 5140 27789 5147 27823
rect 5181 27789 5218 27823
rect 5270 27789 5293 27823
rect 5327 27789 5348 27823
rect 5400 27789 5439 27823
rect 5473 27789 5478 27823
rect 5546 27789 5585 27823
rect 5692 27789 5731 27823
rect 5790 27789 5804 27823
rect 5838 27789 5868 27823
rect 5920 27789 5950 27823
rect 5984 27789 5998 27823
rect 6057 27789 6128 27823
rect 2930 27780 3008 27789
rect 3060 27780 3138 27789
rect 3190 27780 3268 27789
rect 3320 27780 3398 27789
rect 3450 27780 3528 27789
rect 3580 27780 3658 27789
rect 3710 27780 3788 27789
rect 3840 27780 3918 27789
rect 3970 27780 4048 27789
rect 4100 27780 4178 27789
rect 4230 27780 4308 27789
rect 4360 27780 4438 27789
rect 4490 27780 4568 27789
rect 4620 27780 4698 27789
rect 4750 27780 4828 27789
rect 4880 27780 4958 27789
rect 5010 27780 5088 27789
rect 5140 27780 5218 27789
rect 5270 27780 5348 27789
rect 5400 27780 5478 27789
rect 5530 27780 5608 27789
rect 5660 27780 5738 27789
rect 5790 27780 5868 27789
rect 5920 27780 5998 27789
rect 6050 27780 6128 27789
rect 6180 27780 6258 27832
rect 6310 27780 6388 27832
rect 6440 27780 6517 27832
rect 6569 27780 6646 27832
rect 6698 27780 6775 27832
rect 6827 27780 6904 27832
rect 6956 27780 7033 27832
rect 7085 27780 7162 27832
rect 7214 27780 7291 27832
rect 7343 27780 7420 27832
rect 7472 27780 7549 27832
rect 7601 27780 7678 27832
rect 7730 27780 7807 27832
rect 7859 27780 7936 27832
rect 7988 27780 7994 27832
rect 2872 27752 7994 27780
rect 2872 27700 2878 27752
rect 2930 27743 3008 27752
rect 3060 27743 3138 27752
rect 3190 27743 3268 27752
rect 3320 27743 3398 27752
rect 3450 27743 3528 27752
rect 3580 27743 3658 27752
rect 3710 27743 3788 27752
rect 3840 27743 3918 27752
rect 3970 27743 4048 27752
rect 4100 27743 4178 27752
rect 4230 27743 4308 27752
rect 4360 27743 4438 27752
rect 4490 27743 4568 27752
rect 4620 27743 4698 27752
rect 4750 27743 4828 27752
rect 4880 27743 4958 27752
rect 5010 27743 5088 27752
rect 5140 27743 5218 27752
rect 5270 27743 5348 27752
rect 5400 27743 5478 27752
rect 5530 27743 5608 27752
rect 5660 27743 5738 27752
rect 5790 27743 5868 27752
rect 5920 27743 5998 27752
rect 6050 27743 6128 27752
rect 2930 27709 2957 27743
rect 2991 27709 3008 27743
rect 3064 27709 3103 27743
rect 3137 27709 3138 27743
rect 3210 27709 3249 27743
rect 3320 27709 3322 27743
rect 3356 27709 3395 27743
rect 3450 27709 3468 27743
rect 3502 27709 3528 27743
rect 3580 27709 3614 27743
rect 3648 27709 3658 27743
rect 3721 27709 3760 27743
rect 3867 27709 3906 27743
rect 3970 27709 3979 27743
rect 4013 27709 4048 27743
rect 4100 27709 4125 27743
rect 4159 27709 4178 27743
rect 4232 27709 4271 27743
rect 4305 27709 4308 27743
rect 4378 27709 4417 27743
rect 4524 27709 4563 27743
rect 4620 27709 4636 27743
rect 4670 27709 4698 27743
rect 4750 27709 4782 27743
rect 4816 27709 4828 27743
rect 4889 27709 4928 27743
rect 5035 27709 5074 27743
rect 5140 27709 5147 27743
rect 5181 27709 5218 27743
rect 5270 27709 5293 27743
rect 5327 27709 5348 27743
rect 5400 27709 5439 27743
rect 5473 27709 5478 27743
rect 5546 27709 5585 27743
rect 5692 27709 5731 27743
rect 5790 27709 5804 27743
rect 5838 27709 5868 27743
rect 5920 27709 5950 27743
rect 5984 27709 5998 27743
rect 6057 27709 6128 27743
rect 2930 27700 3008 27709
rect 3060 27700 3138 27709
rect 3190 27700 3268 27709
rect 3320 27700 3398 27709
rect 3450 27700 3528 27709
rect 3580 27700 3658 27709
rect 3710 27700 3788 27709
rect 3840 27700 3918 27709
rect 3970 27700 4048 27709
rect 4100 27700 4178 27709
rect 4230 27700 4308 27709
rect 4360 27700 4438 27709
rect 4490 27700 4568 27709
rect 4620 27700 4698 27709
rect 4750 27700 4828 27709
rect 4880 27700 4958 27709
rect 5010 27700 5088 27709
rect 5140 27700 5218 27709
rect 5270 27700 5348 27709
rect 5400 27700 5478 27709
rect 5530 27700 5608 27709
rect 5660 27700 5738 27709
rect 5790 27700 5868 27709
rect 5920 27700 5998 27709
rect 6050 27700 6128 27709
rect 6180 27700 6258 27752
rect 6310 27700 6388 27752
rect 6440 27700 6517 27752
rect 6569 27700 6646 27752
rect 6698 27700 6775 27752
rect 6827 27700 6904 27752
rect 6956 27700 7033 27752
rect 7085 27700 7162 27752
rect 7214 27700 7291 27752
rect 7343 27700 7420 27752
rect 7472 27700 7549 27752
rect 7601 27700 7678 27752
rect 7730 27700 7807 27752
rect 7859 27700 7936 27752
rect 7988 27700 7994 27752
rect 2872 27672 7994 27700
rect 2872 27620 2878 27672
rect 2930 27663 3008 27672
rect 3060 27663 3138 27672
rect 3190 27663 3268 27672
rect 3320 27663 3398 27672
rect 3450 27663 3528 27672
rect 3580 27663 3658 27672
rect 3710 27663 3788 27672
rect 3840 27663 3918 27672
rect 3970 27663 4048 27672
rect 4100 27663 4178 27672
rect 4230 27663 4308 27672
rect 4360 27663 4438 27672
rect 4490 27663 4568 27672
rect 4620 27663 4698 27672
rect 4750 27663 4828 27672
rect 4880 27663 4958 27672
rect 5010 27663 5088 27672
rect 5140 27663 5218 27672
rect 5270 27663 5348 27672
rect 5400 27663 5478 27672
rect 5530 27663 5608 27672
rect 5660 27663 5738 27672
rect 5790 27663 5868 27672
rect 5920 27663 5998 27672
rect 6050 27663 6128 27672
rect 2930 27629 2957 27663
rect 2991 27629 3008 27663
rect 3064 27629 3103 27663
rect 3137 27629 3138 27663
rect 3210 27629 3249 27663
rect 3320 27629 3322 27663
rect 3356 27629 3395 27663
rect 3450 27629 3468 27663
rect 3502 27629 3528 27663
rect 3580 27629 3614 27663
rect 3648 27629 3658 27663
rect 3721 27629 3760 27663
rect 3867 27629 3906 27663
rect 3970 27629 3979 27663
rect 4013 27629 4048 27663
rect 4100 27629 4125 27663
rect 4159 27629 4178 27663
rect 4232 27629 4271 27663
rect 4305 27629 4308 27663
rect 4378 27629 4417 27663
rect 4524 27629 4563 27663
rect 4620 27629 4636 27663
rect 4670 27629 4698 27663
rect 4750 27629 4782 27663
rect 4816 27629 4828 27663
rect 4889 27629 4928 27663
rect 5035 27629 5074 27663
rect 5140 27629 5147 27663
rect 5181 27629 5218 27663
rect 5270 27629 5293 27663
rect 5327 27629 5348 27663
rect 5400 27629 5439 27663
rect 5473 27629 5478 27663
rect 5546 27629 5585 27663
rect 5692 27629 5731 27663
rect 5790 27629 5804 27663
rect 5838 27629 5868 27663
rect 5920 27629 5950 27663
rect 5984 27629 5998 27663
rect 6057 27629 6128 27663
rect 2930 27620 3008 27629
rect 3060 27620 3138 27629
rect 3190 27620 3268 27629
rect 3320 27620 3398 27629
rect 3450 27620 3528 27629
rect 3580 27620 3658 27629
rect 3710 27620 3788 27629
rect 3840 27620 3918 27629
rect 3970 27620 4048 27629
rect 4100 27620 4178 27629
rect 4230 27620 4308 27629
rect 4360 27620 4438 27629
rect 4490 27620 4568 27629
rect 4620 27620 4698 27629
rect 4750 27620 4828 27629
rect 4880 27620 4958 27629
rect 5010 27620 5088 27629
rect 5140 27620 5218 27629
rect 5270 27620 5348 27629
rect 5400 27620 5478 27629
rect 5530 27620 5608 27629
rect 5660 27620 5738 27629
rect 5790 27620 5868 27629
rect 5920 27620 5998 27629
rect 6050 27620 6128 27629
rect 6180 27620 6258 27672
rect 6310 27620 6388 27672
rect 6440 27620 6517 27672
rect 6569 27620 6646 27672
rect 6698 27620 6775 27672
rect 6827 27620 6904 27672
rect 6956 27620 7033 27672
rect 7085 27620 7162 27672
rect 7214 27620 7291 27672
rect 7343 27620 7420 27672
rect 7472 27620 7549 27672
rect 7601 27620 7678 27672
rect 7730 27620 7807 27672
rect 7859 27620 7936 27672
rect 7988 27620 7994 27672
rect 2872 27592 7994 27620
rect 2872 27540 2878 27592
rect 2930 27583 3008 27592
rect 3060 27583 3138 27592
rect 3190 27583 3268 27592
rect 3320 27583 3398 27592
rect 3450 27583 3528 27592
rect 3580 27583 3658 27592
rect 3710 27583 3788 27592
rect 3840 27583 3918 27592
rect 3970 27583 4048 27592
rect 4100 27583 4178 27592
rect 4230 27583 4308 27592
rect 4360 27583 4438 27592
rect 4490 27583 4568 27592
rect 4620 27583 4698 27592
rect 4750 27583 4828 27592
rect 4880 27583 4958 27592
rect 5010 27583 5088 27592
rect 5140 27583 5218 27592
rect 5270 27583 5348 27592
rect 5400 27583 5478 27592
rect 5530 27583 5608 27592
rect 5660 27583 5738 27592
rect 5790 27583 5868 27592
rect 5920 27583 5998 27592
rect 6050 27583 6128 27592
rect 2930 27549 2957 27583
rect 2991 27549 3008 27583
rect 3064 27549 3103 27583
rect 3137 27549 3138 27583
rect 3210 27549 3249 27583
rect 3320 27549 3322 27583
rect 3356 27549 3395 27583
rect 3450 27549 3468 27583
rect 3502 27549 3528 27583
rect 3580 27549 3614 27583
rect 3648 27549 3658 27583
rect 3721 27549 3760 27583
rect 3867 27549 3906 27583
rect 3970 27549 3979 27583
rect 4013 27549 4048 27583
rect 4100 27549 4125 27583
rect 4159 27549 4178 27583
rect 4232 27549 4271 27583
rect 4305 27549 4308 27583
rect 4378 27549 4417 27583
rect 4524 27549 4563 27583
rect 4620 27549 4636 27583
rect 4670 27549 4698 27583
rect 4750 27549 4782 27583
rect 4816 27549 4828 27583
rect 4889 27549 4928 27583
rect 5035 27549 5074 27583
rect 5140 27549 5147 27583
rect 5181 27549 5218 27583
rect 5270 27549 5293 27583
rect 5327 27549 5348 27583
rect 5400 27549 5439 27583
rect 5473 27549 5478 27583
rect 5546 27549 5585 27583
rect 5692 27549 5731 27583
rect 5790 27549 5804 27583
rect 5838 27549 5868 27583
rect 5920 27549 5950 27583
rect 5984 27549 5998 27583
rect 6057 27549 6128 27583
rect 2930 27540 3008 27549
rect 3060 27540 3138 27549
rect 3190 27540 3268 27549
rect 3320 27540 3398 27549
rect 3450 27540 3528 27549
rect 3580 27540 3658 27549
rect 3710 27540 3788 27549
rect 3840 27540 3918 27549
rect 3970 27540 4048 27549
rect 4100 27540 4178 27549
rect 4230 27540 4308 27549
rect 4360 27540 4438 27549
rect 4490 27540 4568 27549
rect 4620 27540 4698 27549
rect 4750 27540 4828 27549
rect 4880 27540 4958 27549
rect 5010 27540 5088 27549
rect 5140 27540 5218 27549
rect 5270 27540 5348 27549
rect 5400 27540 5478 27549
rect 5530 27540 5608 27549
rect 5660 27540 5738 27549
rect 5790 27540 5868 27549
rect 5920 27540 5998 27549
rect 6050 27540 6128 27549
rect 6180 27540 6258 27592
rect 6310 27540 6388 27592
rect 6440 27540 6517 27592
rect 6569 27540 6646 27592
rect 6698 27540 6775 27592
rect 6827 27540 6904 27592
rect 6956 27540 7033 27592
rect 7085 27540 7162 27592
rect 7214 27540 7291 27592
rect 7343 27540 7420 27592
rect 7472 27540 7549 27592
rect 7601 27540 7678 27592
rect 7730 27540 7807 27592
rect 7859 27540 7936 27592
rect 7988 27540 7994 27592
rect 2872 27512 7994 27540
rect 2872 27460 2878 27512
rect 2930 27503 3008 27512
rect 3060 27503 3138 27512
rect 3190 27503 3268 27512
rect 3320 27503 3398 27512
rect 3450 27503 3528 27512
rect 3580 27503 3658 27512
rect 3710 27503 3788 27512
rect 3840 27503 3918 27512
rect 3970 27503 4048 27512
rect 4100 27503 4178 27512
rect 4230 27503 4308 27512
rect 4360 27503 4438 27512
rect 4490 27503 4568 27512
rect 4620 27503 4698 27512
rect 4750 27503 4828 27512
rect 4880 27503 4958 27512
rect 5010 27503 5088 27512
rect 5140 27503 5218 27512
rect 5270 27503 5348 27512
rect 5400 27503 5478 27512
rect 5530 27503 5608 27512
rect 5660 27503 5738 27512
rect 5790 27503 5868 27512
rect 5920 27503 5998 27512
rect 6050 27503 6128 27512
rect 2930 27469 2957 27503
rect 2991 27469 3008 27503
rect 3064 27469 3103 27503
rect 3137 27469 3138 27503
rect 3210 27469 3249 27503
rect 3320 27469 3322 27503
rect 3356 27469 3395 27503
rect 3450 27469 3468 27503
rect 3502 27469 3528 27503
rect 3580 27469 3614 27503
rect 3648 27469 3658 27503
rect 3721 27469 3760 27503
rect 3867 27469 3906 27503
rect 3970 27469 3979 27503
rect 4013 27469 4048 27503
rect 4100 27469 4125 27503
rect 4159 27469 4178 27503
rect 4232 27469 4271 27503
rect 4305 27469 4308 27503
rect 4378 27469 4417 27503
rect 4524 27469 4563 27503
rect 4620 27469 4636 27503
rect 4670 27469 4698 27503
rect 4750 27469 4782 27503
rect 4816 27469 4828 27503
rect 4889 27469 4928 27503
rect 5035 27469 5074 27503
rect 5140 27469 5147 27503
rect 5181 27469 5218 27503
rect 5270 27469 5293 27503
rect 5327 27469 5348 27503
rect 5400 27469 5439 27503
rect 5473 27469 5478 27503
rect 5546 27469 5585 27503
rect 5692 27469 5731 27503
rect 5790 27469 5804 27503
rect 5838 27469 5868 27503
rect 5920 27469 5950 27503
rect 5984 27469 5998 27503
rect 6057 27469 6128 27503
rect 2930 27460 3008 27469
rect 3060 27460 3138 27469
rect 3190 27460 3268 27469
rect 3320 27460 3398 27469
rect 3450 27460 3528 27469
rect 3580 27460 3658 27469
rect 3710 27460 3788 27469
rect 3840 27460 3918 27469
rect 3970 27460 4048 27469
rect 4100 27460 4178 27469
rect 4230 27460 4308 27469
rect 4360 27460 4438 27469
rect 4490 27460 4568 27469
rect 4620 27460 4698 27469
rect 4750 27460 4828 27469
rect 4880 27460 4958 27469
rect 5010 27460 5088 27469
rect 5140 27460 5218 27469
rect 5270 27460 5348 27469
rect 5400 27460 5478 27469
rect 5530 27460 5608 27469
rect 5660 27460 5738 27469
rect 5790 27460 5868 27469
rect 5920 27460 5998 27469
rect 6050 27460 6128 27469
rect 6180 27460 6258 27512
rect 6310 27460 6388 27512
rect 6440 27460 6517 27512
rect 6569 27460 6646 27512
rect 6698 27460 6775 27512
rect 6827 27460 6904 27512
rect 6956 27460 7033 27512
rect 7085 27460 7162 27512
rect 7214 27460 7291 27512
rect 7343 27460 7420 27512
rect 7472 27460 7549 27512
rect 7601 27460 7678 27512
rect 7730 27460 7807 27512
rect 7859 27460 7936 27512
rect 7988 27460 7994 27512
rect 2872 27459 7994 27460
rect 2533 27400 2547 27452
tri 7960 27425 7994 27459 ne
rect 9784 27936 9810 27988
rect 9732 27921 9862 27936
rect 9784 27869 9810 27921
rect 9732 27854 9862 27869
rect 9784 27802 9810 27854
rect 9732 27787 9862 27802
rect 9784 27735 9810 27787
rect 9732 27720 9862 27735
rect 9784 27668 9810 27720
rect 9732 27653 9862 27668
rect 9784 27601 9810 27653
rect 9732 27586 9862 27601
rect 9784 27534 9810 27586
rect 9732 27519 9862 27534
rect 9784 27467 9810 27519
rect 9732 27452 9862 27467
rect 2481 27394 2599 27400
rect 9784 27400 9810 27452
rect 9732 27394 9862 27400
tri 9732 27380 9746 27394 ne
rect 9792 27380 9812 27394
tri 9812 27380 9826 27394 nw
tri 9792 27360 9812 27380 nw
rect 3304 27284 3310 27336
rect 3362 27330 3376 27336
rect 3428 27284 3441 27336
rect 3304 27270 3316 27284
rect 3422 27270 3441 27284
rect 3304 27218 3310 27270
rect 3362 27218 3376 27224
rect 3428 27218 3441 27270
rect 5383 27334 5513 27335
rect 5383 27218 5389 27334
rect 5505 27218 5513 27334
rect 5383 27217 5513 27218
tri 7271 27163 7305 27197 ne
tri 7436 27163 7470 27197 nw
tri 7635 27163 7669 27197 ne
rect 2816 27008 2868 27138
rect 7305 26968 7318 26998
rect 7669 26968 7679 26996
rect 7074 26922 7192 26954
rect 7074 26888 7080 26922
rect 7114 26888 7152 26922
rect 7186 26888 7192 26922
tri 6797 26853 6831 26887 se
rect 3268 26847 3458 26853
rect 3268 26795 3269 26847
rect 3321 26795 3337 26847
rect 3389 26795 3405 26847
rect 3457 26795 3458 26847
rect 3268 26763 3458 26795
rect 3268 26711 3269 26763
rect 3321 26711 3337 26763
rect 3389 26711 3405 26763
rect 3457 26711 3458 26763
rect 3268 26679 3458 26711
rect 3268 26627 3269 26679
rect 3321 26627 3337 26679
rect 3389 26627 3405 26679
rect 3457 26627 3458 26679
rect 3268 26594 3458 26627
rect 3268 26542 3269 26594
rect 3321 26542 3337 26594
rect 3389 26542 3405 26594
rect 3457 26542 3458 26594
rect 3268 26509 3458 26542
rect 3268 26457 3269 26509
rect 3321 26457 3337 26509
rect 3389 26457 3405 26509
rect 3457 26457 3458 26509
rect 3268 26451 3458 26457
rect 7074 26849 7192 26888
rect 7074 26815 7080 26849
rect 7114 26815 7152 26849
rect 7186 26815 7192 26849
rect 7074 26776 7192 26815
rect 7074 26742 7080 26776
rect 7114 26742 7152 26776
rect 7186 26742 7192 26776
rect 7074 26703 7192 26742
rect 7074 26669 7080 26703
rect 7114 26669 7152 26703
rect 7186 26669 7192 26703
rect 7074 26630 7192 26669
rect 7074 26596 7080 26630
rect 7114 26596 7152 26630
rect 7186 26596 7192 26630
rect 7074 26557 7192 26596
rect 7074 26523 7080 26557
rect 7114 26523 7152 26557
rect 7186 26523 7192 26557
rect 7074 26484 7192 26523
rect 7074 26450 7080 26484
rect 7114 26450 7152 26484
rect 7186 26450 7192 26484
rect 7074 26411 7192 26450
rect 7074 26377 7080 26411
rect 7114 26377 7152 26411
rect 7186 26377 7192 26411
rect 7074 26338 7192 26377
rect 7074 26304 7080 26338
rect 7114 26304 7152 26338
rect 7186 26304 7192 26338
rect 7074 26265 7192 26304
rect 7074 26231 7080 26265
rect 7114 26231 7152 26265
rect 7186 26231 7192 26265
rect 5091 26156 5575 26208
rect 7074 26192 7192 26231
rect 7074 26158 7080 26192
rect 7114 26158 7152 26192
rect 7186 26158 7192 26192
rect 2820 25466 2950 25531
rect 3999 24701 4051 26128
rect 7074 26119 7192 26158
rect 7074 26085 7080 26119
rect 7114 26085 7152 26119
rect 7186 26085 7192 26119
rect 4344 24701 4396 26083
rect 4500 24701 4552 26083
rect 4656 24701 4708 26083
rect 4812 24701 4864 26083
rect 4968 24701 5020 26083
rect 5124 24701 5176 26083
rect 5280 24701 5332 26083
rect 5436 24701 5488 26083
rect 5592 24701 5644 26083
rect 5937 24701 5989 26083
rect 7074 26046 7192 26085
rect 7074 26012 7080 26046
rect 7114 26012 7152 26046
rect 7186 26012 7192 26046
rect 7074 25973 7192 26012
rect 7074 25939 7080 25973
rect 7114 25939 7152 25973
rect 7186 25939 7192 25973
rect 7074 25900 7192 25939
rect 7074 25866 7080 25900
rect 7114 25866 7152 25900
rect 7186 25866 7192 25900
rect 7074 25827 7192 25866
rect 7074 25793 7080 25827
rect 7114 25793 7152 25827
rect 7186 25793 7192 25827
rect 7074 25754 7192 25793
rect 7074 25720 7080 25754
rect 7114 25720 7152 25754
rect 7186 25720 7192 25754
rect 7074 25681 7192 25720
rect 7074 25647 7080 25681
rect 7114 25647 7152 25681
rect 7186 25647 7192 25681
rect 7074 25608 7192 25647
rect 7074 25574 7080 25608
rect 7114 25574 7152 25608
rect 7186 25574 7192 25608
rect 7074 25535 7192 25574
rect 7074 25501 7080 25535
rect 7114 25501 7152 25535
rect 7186 25501 7192 25535
rect 7074 25462 7192 25501
rect 7074 25428 7080 25462
rect 7114 25428 7152 25462
rect 7186 25428 7192 25462
rect 7074 25389 7192 25428
rect 7074 25355 7080 25389
rect 7114 25355 7152 25389
rect 7186 25355 7192 25389
rect 7074 25316 7192 25355
rect 7074 25282 7080 25316
rect 7114 25282 7152 25316
rect 7186 25282 7192 25316
rect 7074 25243 7192 25282
rect 7074 25209 7080 25243
rect 7114 25209 7152 25243
rect 7186 25209 7192 25243
rect 7074 25170 7192 25209
rect 7074 25136 7080 25170
rect 7114 25136 7152 25170
rect 7186 25136 7192 25170
rect 7074 25097 7192 25136
rect 7074 25063 7080 25097
rect 7114 25063 7152 25097
rect 7186 25063 7192 25097
rect 7074 25024 7192 25063
rect 7074 24990 7080 25024
rect 7114 24990 7152 25024
rect 7186 24990 7192 25024
rect 7074 24951 7192 24990
rect 7074 24917 7080 24951
rect 7114 24917 7152 24951
rect 7186 24917 7192 24951
rect 7074 24878 7192 24917
rect 7074 24844 7080 24878
rect 7114 24844 7152 24878
rect 7186 24844 7192 24878
rect 7074 24805 7192 24844
rect 7074 24771 7080 24805
rect 7114 24771 7152 24805
rect 7186 24771 7192 24805
rect 7074 24732 7192 24771
rect 7074 24698 7080 24732
rect 7114 24698 7152 24732
rect 7186 24698 7192 24732
rect 7074 24659 7192 24698
rect 7074 24625 7080 24659
rect 7114 24625 7152 24659
rect 7186 24625 7192 24659
rect 7074 24586 7192 24625
rect 7074 24552 7080 24586
rect 7114 24552 7152 24586
rect 7186 24552 7192 24586
rect 4050 24522 6218 24523
rect 4050 24470 4056 24522
rect 4108 24517 4187 24522
rect 4239 24517 4318 24522
rect 4370 24517 4449 24522
rect 4501 24517 4580 24522
rect 4632 24517 4711 24522
rect 4763 24517 4842 24522
rect 4894 24517 4973 24522
rect 5025 24517 5104 24522
rect 5156 24517 5235 24522
rect 5287 24517 5365 24522
rect 5417 24517 5495 24522
rect 5547 24517 5625 24522
rect 5677 24517 5755 24522
rect 5807 24517 5885 24522
rect 5937 24517 6015 24522
rect 4108 24483 4135 24517
rect 4169 24483 4187 24517
rect 4242 24483 4281 24517
rect 4315 24483 4318 24517
rect 4388 24483 4427 24517
rect 4534 24483 4573 24517
rect 4632 24483 4646 24517
rect 4680 24483 4711 24517
rect 4763 24483 4792 24517
rect 4826 24483 4842 24517
rect 4899 24483 4938 24517
rect 4972 24483 4973 24517
rect 5045 24483 5084 24517
rect 5156 24483 5157 24517
rect 5191 24483 5230 24517
rect 5287 24483 5303 24517
rect 5337 24483 5365 24517
rect 5417 24483 5449 24517
rect 5483 24483 5495 24517
rect 5556 24483 5595 24517
rect 5701 24483 5739 24517
rect 5807 24483 5811 24517
rect 5845 24483 5883 24517
rect 5937 24483 5955 24517
rect 5989 24483 6015 24517
rect 4108 24470 4187 24483
rect 4239 24470 4318 24483
rect 4370 24470 4449 24483
rect 4501 24470 4580 24483
rect 4632 24470 4711 24483
rect 4763 24470 4842 24483
rect 4894 24470 4973 24483
rect 5025 24470 5104 24483
rect 5156 24470 5235 24483
rect 5287 24470 5365 24483
rect 5417 24470 5495 24483
rect 5547 24470 5625 24483
rect 5677 24470 5755 24483
rect 5807 24470 5885 24483
rect 5937 24470 6015 24483
rect 6067 24470 6218 24522
rect 4050 24458 6218 24470
rect 4050 24406 4056 24458
rect 4108 24406 4187 24458
rect 4239 24406 4318 24458
rect 4370 24406 4449 24458
rect 4501 24406 4580 24458
rect 4632 24406 4711 24458
rect 4763 24406 4842 24458
rect 4894 24406 4973 24458
rect 5025 24406 5104 24458
rect 5156 24406 5235 24458
rect 5287 24406 5365 24458
rect 5417 24406 5495 24458
rect 5547 24406 5625 24458
rect 5677 24406 5755 24458
rect 5807 24406 5885 24458
rect 5937 24406 6015 24458
rect 6067 24406 6218 24458
rect 4050 24394 6218 24406
rect 4050 24342 4056 24394
rect 4108 24381 4187 24394
rect 4239 24381 4318 24394
rect 4370 24381 4449 24394
rect 4501 24381 4580 24394
rect 4632 24381 4711 24394
rect 4763 24381 4842 24394
rect 4894 24381 4973 24394
rect 5025 24381 5104 24394
rect 5156 24381 5235 24394
rect 5287 24381 5365 24394
rect 5417 24381 5495 24394
rect 5547 24381 5625 24394
rect 5677 24381 5755 24394
rect 5807 24381 5885 24394
rect 5937 24381 6015 24394
rect 4108 24347 4135 24381
rect 4169 24347 4187 24381
rect 4242 24347 4281 24381
rect 4315 24347 4318 24381
rect 4388 24347 4427 24381
rect 4534 24347 4573 24381
rect 4632 24347 4646 24381
rect 4680 24347 4711 24381
rect 4763 24347 4792 24381
rect 4826 24347 4842 24381
rect 4899 24347 4938 24381
rect 4972 24347 4973 24381
rect 5045 24347 5084 24381
rect 5156 24347 5157 24381
rect 5191 24347 5230 24381
rect 5287 24347 5303 24381
rect 5337 24347 5365 24381
rect 5417 24347 5449 24381
rect 5483 24347 5495 24381
rect 5556 24347 5595 24381
rect 5701 24347 5739 24381
rect 5807 24347 5811 24381
rect 5845 24347 5883 24381
rect 5937 24347 5955 24381
rect 5989 24347 6015 24381
rect 4108 24342 4187 24347
rect 4239 24342 4318 24347
rect 4370 24342 4449 24347
rect 4501 24342 4580 24347
rect 4632 24342 4711 24347
rect 4763 24342 4842 24347
rect 4894 24342 4973 24347
rect 5025 24342 5104 24347
rect 5156 24342 5235 24347
rect 5287 24342 5365 24347
rect 5417 24342 5495 24347
rect 5547 24342 5625 24347
rect 5677 24342 5755 24347
rect 5807 24342 5885 24347
rect 5937 24342 6015 24347
rect 6067 24342 6218 24394
rect 4050 24341 6218 24342
rect 7074 24513 7192 24552
tri 9792 24537 9812 24557 sw
tri 9732 24523 9746 24537 se
rect 9792 24523 9812 24537
tri 9812 24523 9826 24537 sw
rect 7074 24479 7080 24513
rect 7114 24479 7152 24513
rect 7186 24479 7192 24513
rect 7074 24440 7192 24479
rect 7074 24406 7080 24440
rect 7114 24406 7152 24440
rect 7186 24406 7192 24440
rect 7074 24367 7192 24406
rect 7074 24333 7080 24367
rect 7114 24333 7152 24367
rect 7186 24333 7192 24367
rect 7988 24517 8040 24523
rect 7988 24399 8040 24465
rect 7988 24341 8040 24347
rect 9732 24517 9862 24523
rect 9784 24465 9810 24517
rect 9732 24399 9862 24465
rect 9784 24347 9810 24399
rect 9732 24341 9862 24347
rect 10710 24517 10828 24523
rect 10762 24465 10776 24517
rect 10710 24399 10828 24465
rect 10762 24347 10776 24399
rect 10710 24341 10828 24347
rect 7074 24294 7192 24333
tri 9732 24327 9746 24341 ne
rect 9792 24327 9812 24341
tri 9812 24327 9826 24341 nw
tri 9792 24307 9812 24327 nw
rect 7074 24260 7080 24294
rect 7114 24260 7152 24294
rect 7186 24260 7192 24294
rect 7074 24221 7192 24260
rect 4451 24144 4503 24190
rect 7074 24187 7080 24221
rect 7114 24187 7152 24221
rect 7186 24187 7192 24221
rect 7074 24148 7192 24187
rect 4451 24114 4507 24144
tri 4507 24114 4537 24144 nw
rect 7074 24114 7080 24148
rect 7114 24114 7152 24148
rect 7186 24114 7192 24148
rect 282 22749 334 22755
rect 282 22685 334 22697
rect 282 122 334 22633
rect 4451 19429 4503 24114
tri 4503 24110 4507 24114 nw
rect 7074 24075 7192 24114
rect 7074 24041 7080 24075
rect 7114 24041 7152 24075
rect 7186 24041 7192 24075
rect 7074 24002 7192 24041
rect 7074 23968 7080 24002
rect 7114 23968 7152 24002
rect 7186 23968 7192 24002
rect 7074 23929 7192 23968
rect 7074 23895 7080 23929
rect 7114 23895 7152 23929
rect 7186 23895 7192 23929
rect 7074 23856 7192 23895
rect 7074 23822 7080 23856
rect 7114 23822 7152 23856
rect 7186 23822 7192 23856
rect 7074 23782 7192 23822
rect 7074 23748 7080 23782
rect 7114 23748 7152 23782
rect 7186 23748 7192 23782
rect 7074 23708 7192 23748
rect 7074 23674 7080 23708
rect 7114 23674 7152 23708
rect 7186 23674 7192 23708
rect 7074 23634 7192 23674
rect 7074 23600 7080 23634
rect 7114 23600 7152 23634
rect 7186 23600 7192 23634
rect 7074 23560 7192 23600
rect 7074 23526 7080 23560
rect 7114 23526 7152 23560
rect 7186 23526 7192 23560
rect 7074 23486 7192 23526
rect 7074 23452 7080 23486
rect 7114 23452 7152 23486
rect 7186 23452 7192 23486
rect 7074 23412 7192 23452
rect 7074 23378 7080 23412
rect 7114 23378 7152 23412
rect 7186 23378 7192 23412
rect 7074 23268 7192 23378
rect 6050 23265 7774 23268
rect 6050 23213 6056 23265
rect 6108 23256 6123 23265
rect 6175 23256 6190 23265
rect 6242 23256 6257 23265
rect 6309 23256 6324 23265
rect 6376 23256 6391 23265
rect 6443 23256 6458 23265
rect 6510 23256 6525 23265
rect 6577 23256 6592 23265
rect 6644 23256 6659 23265
rect 6711 23256 6726 23265
rect 6778 23256 6792 23265
rect 6844 23256 6858 23265
rect 6910 23256 6924 23265
rect 6976 23256 6990 23265
rect 7042 23256 7056 23265
rect 7108 23256 7122 23265
rect 7174 23256 7188 23265
rect 7240 23256 7254 23265
rect 7306 23256 7320 23265
rect 7372 23256 7386 23265
rect 7438 23256 7452 23265
rect 7504 23256 7518 23265
rect 7570 23256 7584 23265
rect 7636 23256 7650 23265
rect 7702 23256 7716 23265
rect 7768 23213 7774 23265
rect 6050 23195 6067 23213
rect 7757 23195 7774 23213
rect 6050 23143 6056 23195
rect 7768 23143 7774 23195
rect 6050 23125 6067 23143
rect 7757 23125 7774 23143
rect 6050 23073 6056 23125
rect 7768 23073 7774 23125
rect 6050 23055 6067 23073
rect 7757 23055 7774 23073
rect 6050 23003 6056 23055
rect 7768 23003 7774 23055
rect 6050 22985 6067 23003
rect 7757 22985 7774 23003
rect 6050 22933 6056 22985
rect 7768 22933 7774 22985
rect 6050 22915 6067 22933
rect 7757 22915 7774 22933
rect 6050 22863 6056 22915
rect 7768 22863 7774 22915
rect 6050 22790 6067 22863
rect 7757 22790 7774 22863
rect 6050 22751 7774 22790
rect 6050 22717 6067 22751
rect 6101 22717 6139 22751
rect 6173 22717 6211 22751
rect 6245 22717 6283 22751
rect 6317 22717 6355 22751
rect 6389 22717 6427 22751
rect 6461 22717 6499 22751
rect 6533 22717 6571 22751
rect 6605 22717 6643 22751
rect 6677 22717 6715 22751
rect 6749 22717 6787 22751
rect 6821 22717 6859 22751
rect 6893 22717 6931 22751
rect 6965 22717 7003 22751
rect 7037 22717 7075 22751
rect 7109 22717 7147 22751
rect 7181 22717 7219 22751
rect 7253 22717 7291 22751
rect 7325 22717 7363 22751
rect 7397 22717 7435 22751
rect 7469 22717 7507 22751
rect 7541 22717 7579 22751
rect 7613 22717 7651 22751
rect 7685 22717 7723 22751
rect 7757 22717 7774 22751
rect 6050 22678 7774 22717
rect 8223 22703 8229 22755
rect 8281 22703 8293 22755
rect 8345 22703 8351 22755
rect 6050 22644 6067 22678
rect 6101 22644 6139 22678
rect 6173 22644 6211 22678
rect 6245 22644 6283 22678
rect 6317 22644 6355 22678
rect 6389 22644 6427 22678
rect 6461 22644 6499 22678
rect 6533 22644 6571 22678
rect 6605 22644 6643 22678
rect 6677 22644 6715 22678
rect 6749 22644 6787 22678
rect 6821 22644 6859 22678
rect 6893 22644 6931 22678
rect 6965 22644 7003 22678
rect 7037 22644 7075 22678
rect 7109 22644 7147 22678
rect 7181 22644 7219 22678
rect 7253 22644 7291 22678
rect 7325 22644 7363 22678
rect 7397 22644 7435 22678
rect 7469 22644 7507 22678
rect 7541 22644 7579 22678
rect 7613 22644 7651 22678
rect 7685 22644 7723 22678
rect 7757 22644 7774 22678
rect 6050 22605 7774 22644
rect 6050 22571 6067 22605
rect 6101 22571 6139 22605
rect 6173 22571 6211 22605
rect 6245 22571 6283 22605
rect 6317 22571 6355 22605
rect 6389 22571 6427 22605
rect 6461 22571 6499 22605
rect 6533 22571 6571 22605
rect 6605 22571 6643 22605
rect 6677 22571 6715 22605
rect 6749 22571 6787 22605
rect 6821 22571 6859 22605
rect 6893 22571 6931 22605
rect 6965 22571 7003 22605
rect 7037 22571 7075 22605
rect 7109 22571 7147 22605
rect 7181 22571 7219 22605
rect 7253 22571 7291 22605
rect 7325 22571 7363 22605
rect 7397 22571 7435 22605
rect 7469 22571 7507 22605
rect 7541 22571 7579 22605
rect 7613 22571 7651 22605
rect 7685 22571 7723 22605
rect 7757 22571 7774 22605
rect 6050 22532 7774 22571
rect 6050 22498 6067 22532
rect 6101 22498 6139 22532
rect 6173 22498 6211 22532
rect 6245 22498 6283 22532
rect 6317 22498 6355 22532
rect 6389 22498 6427 22532
rect 6461 22498 6499 22532
rect 6533 22498 6571 22532
rect 6605 22498 6643 22532
rect 6677 22498 6715 22532
rect 6749 22498 6787 22532
rect 6821 22498 6859 22532
rect 6893 22498 6931 22532
rect 6965 22498 7003 22532
rect 7037 22498 7075 22532
rect 7109 22498 7147 22532
rect 7181 22498 7219 22532
rect 7253 22498 7291 22532
rect 7325 22498 7363 22532
rect 7397 22498 7435 22532
rect 7469 22498 7507 22532
rect 7541 22498 7579 22532
rect 7613 22498 7651 22532
rect 7685 22498 7723 22532
rect 7757 22498 7774 22532
rect 6050 22486 7774 22498
rect 6846 21152 7104 21158
rect 6846 21100 6847 21152
rect 6899 21100 6949 21152
rect 7001 21100 7051 21152
rect 7103 21100 7104 21152
rect 6846 21068 7104 21100
rect 6846 21016 6847 21068
rect 6899 21016 6949 21068
rect 7001 21016 7051 21068
rect 7103 21016 7104 21068
rect 6846 20984 7104 21016
rect 6846 20932 6847 20984
rect 6899 20932 6949 20984
rect 7001 20932 7051 20984
rect 7103 20932 7104 20984
rect 6846 20900 7104 20932
rect 6846 20848 6847 20900
rect 6899 20848 6949 20900
rect 7001 20848 7051 20900
rect 7103 20848 7104 20900
rect 6846 20816 7104 20848
rect 6846 20764 6847 20816
rect 6899 20764 6949 20816
rect 7001 20764 7051 20816
rect 7103 20764 7104 20816
tri 4503 20099 4537 20133 sw
rect 4594 20048 4623 20053
tri 4623 20048 4628 20053 nw
tri 4594 20019 4623 20048 nw
tri 4693 19943 4727 19977 se
rect 4727 19924 4803 19980
tri 4769 19863 4803 19897 ne
tri 4594 19787 4628 19821 sw
tri 4594 19707 4628 19741 nw
tri 4798 19660 4803 19665 se
tri 4797 19659 4798 19660 se
rect 4798 19659 4803 19660
tri 4769 19631 4797 19659 se
rect 4797 19631 4803 19659
tri 4594 19508 4595 19509 sw
rect 4594 19503 4595 19508
tri 4595 19503 4600 19508 sw
rect 4594 19480 4600 19503
tri 4600 19480 4623 19503 sw
rect 4893 19480 4945 20048
rect 6009 19887 6015 19939
rect 6067 19887 6079 19939
rect 6131 19887 6283 19939
tri 6131 19780 6165 19814 se
rect 6165 19808 6217 19814
tri 6217 19780 6251 19814 sw
rect 6165 19744 6217 19756
tri 6131 19706 6159 19734 ne
rect 6159 19706 6165 19734
tri 6159 19700 6165 19706 ne
rect 6217 19706 6223 19734
tri 6223 19706 6251 19734 nw
tri 6217 19700 6223 19706 nw
rect 6165 19686 6217 19692
rect 6364 19694 6416 19706
rect 6364 19660 6373 19694
rect 6407 19660 6416 19694
rect 6009 19575 6015 19627
rect 6067 19575 6079 19627
rect 6131 19575 6283 19627
rect 6364 19622 6416 19660
rect 6364 19588 6373 19622
rect 6407 19588 6416 19622
rect 6364 19557 6416 19588
rect 6165 19507 6217 19513
tri 6143 19480 6165 19502 se
rect 4594 19478 4623 19480
tri 4623 19478 4625 19480 sw
tri 6141 19478 6143 19480 se
rect 6143 19478 6165 19480
rect 4594 19475 4625 19478
tri 4625 19475 4628 19478 sw
tri 6138 19475 6141 19478 se
rect 6141 19475 6165 19478
tri 6131 19468 6138 19475 se
rect 6138 19468 6165 19475
tri 6217 19478 6241 19502 sw
rect 6364 19493 6416 19505
rect 6217 19468 6241 19478
tri 6241 19468 6251 19478 sw
rect 6165 19443 6217 19455
rect 4451 19422 4530 19429
tri 4530 19422 4537 19429 nw
rect 4451 19416 4524 19422
tri 4524 19416 4530 19422 nw
tri 6131 19416 6137 19422 ne
rect 6137 19416 6165 19422
rect 4451 19414 4522 19416
tri 4522 19414 4524 19416 nw
tri 6137 19414 6139 19416 ne
rect 6139 19414 6165 19416
rect 4451 19405 4513 19414
tri 4513 19405 4522 19414 nw
tri 6139 19405 6148 19414 ne
rect 6148 19405 6165 19414
rect 4451 18542 4503 19405
tri 4503 19395 4513 19405 nw
tri 6148 19395 6158 19405 ne
rect 6158 19395 6165 19405
tri 6158 19388 6165 19395 ne
rect 6217 19416 6245 19422
tri 6245 19416 6251 19422 nw
rect 6217 19414 6243 19416
tri 6243 19414 6245 19416 nw
rect 6217 19405 6234 19414
tri 6234 19405 6243 19414 nw
rect 6364 19405 6416 19441
rect 6165 19385 6217 19391
tri 6217 19388 6234 19405 nw
rect 6364 19371 6373 19405
rect 6407 19371 6416 19405
rect 6364 19359 6416 19371
rect 6846 19666 7104 20764
rect 7710 21152 7762 21158
rect 7710 21085 7762 21100
rect 7710 21018 7762 21033
rect 7710 20951 7762 20966
rect 7710 20884 7762 20899
rect 7710 20816 7762 20832
tri 7104 19666 7137 19699 sw
rect 7710 19672 7762 20764
rect 6846 19665 7137 19666
tri 7137 19665 7138 19666 sw
rect 6846 19659 7576 19665
rect 6846 19625 6972 19659
rect 7006 19625 7052 19659
rect 7086 19625 7132 19659
rect 7166 19625 7212 19659
rect 7246 19625 7292 19659
rect 7326 19625 7372 19659
rect 7406 19625 7451 19659
rect 7485 19625 7530 19659
rect 7564 19625 7576 19659
rect 6846 19619 7576 19625
rect 6846 19602 7121 19619
tri 7121 19602 7138 19619 nw
rect 7618 19602 7664 19614
rect 6846 19522 7104 19602
tri 7104 19585 7121 19602 nw
rect 7618 19568 7624 19602
rect 7658 19568 7664 19602
tri 7104 19522 7125 19543 sw
tri 7597 19522 7618 19543 se
rect 7618 19522 7664 19568
rect 6846 19515 7125 19522
tri 7125 19515 7132 19522 sw
tri 7590 19515 7597 19522 se
rect 7597 19515 7664 19522
rect 6846 19509 7132 19515
tri 7132 19509 7138 19515 sw
tri 7584 19509 7590 19515 se
rect 7590 19509 7664 19515
rect 6846 19508 7664 19509
rect 6846 19503 7624 19508
rect 6846 19469 7116 19503
rect 7150 19469 7199 19503
rect 7233 19469 7282 19503
rect 7316 19469 7365 19503
rect 7399 19469 7448 19503
rect 7482 19469 7530 19503
rect 7564 19474 7624 19503
rect 7658 19474 7664 19508
rect 7564 19469 7664 19474
rect 6846 19463 7664 19469
rect 6846 19450 7125 19463
tri 7125 19450 7138 19463 nw
tri 7584 19450 7597 19463 ne
rect 7597 19450 7664 19463
rect 6846 19380 7104 19450
tri 7104 19429 7125 19450 nw
tri 7597 19429 7618 19450 ne
rect 7618 19414 7664 19450
tri 7104 19380 7111 19387 sw
rect 7618 19380 7624 19414
rect 7658 19380 7664 19414
rect 6846 19378 7111 19380
tri 7111 19378 7113 19380 sw
rect 6846 19353 7113 19378
tri 7113 19353 7138 19378 sw
rect 7618 19368 7664 19380
rect 7710 19594 7762 19620
rect 7710 19573 7716 19594
rect 7750 19573 7762 19594
rect 7710 19488 7716 19521
rect 7750 19515 7762 19521
rect 7750 19488 7756 19515
tri 7756 19509 7762 19515 nw
rect 8711 19808 8763 19814
rect 8711 19744 8763 19756
rect 7710 19450 7756 19488
rect 7710 19416 7716 19450
rect 7750 19416 7756 19450
rect 7710 19378 7756 19416
rect 6846 19347 7448 19353
rect 6009 19263 6015 19315
rect 6067 19263 6079 19315
rect 6131 19263 6283 19315
rect 6846 19313 6972 19347
rect 7006 19313 7058 19347
rect 7092 19313 7144 19347
rect 7178 19313 7230 19347
rect 7264 19313 7316 19347
rect 7350 19313 7402 19347
rect 7436 19313 7448 19347
rect 6846 19307 7448 19313
rect 7710 19344 7716 19378
rect 7750 19344 7756 19378
rect 6846 19306 7137 19307
tri 7137 19306 7138 19307 nw
rect 7710 19306 7756 19344
rect 6846 19292 7123 19306
tri 7123 19292 7137 19306 nw
rect 6846 19280 7111 19292
tri 7111 19280 7123 19292 nw
rect 7618 19280 7664 19292
rect 6364 19231 6416 19243
rect 6364 19197 6373 19231
rect 6407 19197 6416 19231
tri 6134 19157 6165 19188 se
rect 6165 19182 6217 19188
tri 6133 19156 6134 19157 se
rect 6134 19156 6165 19157
tri 6217 19157 6248 19188 sw
rect 6217 19156 6248 19157
tri 6248 19156 6249 19157 sw
rect 6364 19156 6416 19197
rect 6165 19118 6217 19130
tri 6131 19098 6143 19110 ne
rect 6143 19098 6165 19110
tri 6143 19090 6151 19098 ne
rect 6151 19090 6165 19098
tri 6151 19081 6160 19090 ne
rect 6160 19081 6165 19090
tri 6160 19076 6165 19081 ne
rect 6364 19122 6373 19156
rect 6407 19122 6416 19156
rect 6217 19098 6239 19110
tri 6239 19098 6251 19110 nw
rect 6217 19090 6231 19098
tri 6231 19090 6239 19098 nw
rect 6217 19081 6222 19090
tri 6222 19081 6231 19090 nw
rect 6364 19089 6416 19122
tri 6217 19076 6222 19081 nw
rect 6165 19060 6217 19066
rect 6364 19025 6416 19037
rect 6009 18951 6015 19003
rect 6067 18951 6079 19003
rect 6131 18951 6283 19003
rect 6364 18972 6373 18973
rect 6407 18972 6416 18973
rect 6364 18931 6416 18972
rect 6364 18897 6373 18931
rect 6407 18897 6416 18931
rect 6165 18886 6217 18892
tri 6143 18856 6165 18878 se
tri 6131 18844 6143 18856 se
rect 6143 18844 6165 18856
tri 6217 18856 6239 18878 sw
rect 6364 18856 6416 18897
rect 6217 18844 6239 18856
tri 6239 18844 6251 18856 sw
rect 6165 18822 6217 18834
tri 6131 18781 6148 18798 ne
rect 6148 18781 6165 18798
tri 6148 18764 6165 18781 ne
rect 6364 18822 6373 18856
rect 6407 18822 6416 18856
rect 6217 18781 6234 18798
tri 6234 18781 6251 18798 nw
rect 6364 18781 6416 18822
rect 6165 18764 6217 18770
tri 6217 18764 6234 18781 nw
rect 6364 18747 6373 18781
rect 6407 18747 6416 18781
rect 6364 18735 6416 18747
rect 6846 19058 7104 19280
tri 7104 19273 7111 19280 nw
rect 7618 19246 7624 19280
rect 7658 19246 7664 19280
rect 7618 19206 7664 19246
rect 7132 19191 7576 19197
rect 7132 19157 7144 19191
rect 7178 19157 7222 19191
rect 7256 19157 7299 19191
rect 7333 19157 7376 19191
rect 7410 19157 7453 19191
rect 7487 19157 7530 19191
rect 7564 19157 7576 19191
rect 7132 19151 7576 19157
tri 7442 19132 7461 19151 ne
rect 7461 19132 7576 19151
tri 7461 19117 7476 19132 ne
tri 7104 19058 7121 19075 sw
rect 6846 19041 7121 19058
tri 7121 19041 7138 19058 sw
rect 6846 19035 7448 19041
rect 6846 19001 6972 19035
rect 7006 19001 7058 19035
rect 7092 19001 7144 19035
rect 7178 19001 7230 19035
rect 7264 19001 7316 19035
rect 7350 19001 7402 19035
rect 7436 19001 7448 19035
rect 6846 18995 7448 19001
rect 6846 18984 7127 18995
tri 7127 18984 7138 18995 nw
rect 6846 18762 7104 18984
tri 7104 18961 7127 18984 nw
tri 7469 18912 7476 18919 se
rect 7476 18912 7576 19132
tri 7467 18910 7469 18912 se
rect 7469 18910 7576 18912
tri 7445 18888 7467 18910 se
rect 7467 18888 7576 18910
tri 7442 18885 7445 18888 se
rect 7445 18885 7576 18888
rect 7132 18879 7576 18885
rect 7132 18845 7144 18879
rect 7178 18845 7222 18879
rect 7256 18845 7299 18879
rect 7333 18845 7376 18879
rect 7410 18845 7453 18879
rect 7487 18856 7530 18879
rect 7564 18856 7576 18879
rect 7487 18845 7524 18856
rect 7132 18839 7524 18845
tri 7442 18836 7445 18839 ne
rect 7445 18836 7524 18839
tri 7445 18805 7476 18836 ne
rect 7476 18804 7524 18836
rect 7476 18792 7576 18804
tri 7104 18762 7105 18763 sw
rect 6846 18729 7105 18762
tri 7105 18729 7138 18762 sw
rect 7476 18740 7524 18792
rect 6846 18723 7448 18729
rect 6009 18639 6015 18691
rect 6067 18639 6079 18691
rect 6131 18639 6283 18691
rect 6846 18689 6972 18723
rect 7006 18689 7058 18723
rect 7092 18689 7144 18723
rect 7178 18689 7230 18723
rect 7264 18689 7316 18723
rect 7350 18689 7402 18723
rect 7436 18689 7448 18723
rect 6846 18683 7448 18689
rect 6846 18654 7109 18683
tri 7109 18654 7138 18683 nw
rect 6364 18625 6416 18631
tri 6235 18556 6245 18566 se
rect 6245 18562 6297 18568
tri 4503 18542 4517 18556 sw
tri 6221 18542 6235 18556 se
rect 6235 18542 6245 18556
rect 4451 18532 4517 18542
tri 4517 18532 4527 18542 sw
tri 6211 18532 6221 18542 se
rect 6221 18532 6245 18542
rect 4451 18522 4527 18532
tri 4527 18522 4537 18532 sw
rect 3833 18436 3839 18488
rect 3891 18436 3924 18488
rect 3976 18436 4009 18488
rect 4061 18436 4093 18488
rect 4145 18436 4177 18488
rect 4229 18436 4235 18488
rect 4451 18476 4503 18522
rect 6245 18498 6297 18510
tri 6211 18480 6217 18486 ne
rect 6217 18480 6245 18486
tri 6217 18476 6221 18480 ne
rect 6221 18476 6245 18480
tri 6221 18466 6231 18476 ne
rect 6231 18466 6245 18476
tri 6231 18452 6245 18466 ne
rect 6364 18561 6416 18573
rect 6364 18508 6373 18509
rect 6407 18508 6416 18509
rect 6364 18496 6416 18508
rect 6245 18440 6297 18446
rect 3833 18408 4235 18436
rect 3833 18356 3839 18408
rect 3891 18356 3924 18408
rect 3976 18356 4009 18408
rect 4061 18356 4093 18408
rect 4145 18356 4177 18408
rect 4229 18356 4235 18408
rect 6846 18432 7104 18654
tri 7104 18649 7109 18654 nw
tri 7449 18580 7476 18607 se
rect 7476 18580 7576 18740
tri 7442 18573 7449 18580 se
rect 7449 18573 7576 18580
rect 7132 18567 7576 18573
rect 7132 18533 7144 18567
rect 7178 18533 7222 18567
rect 7256 18533 7299 18567
rect 7333 18533 7376 18567
rect 7410 18533 7453 18567
rect 7487 18533 7530 18567
rect 7564 18533 7576 18567
rect 7132 18527 7576 18533
tri 7442 18506 7463 18527 ne
rect 7463 18506 7576 18527
tri 7463 18493 7476 18506 ne
tri 7104 18432 7123 18451 sw
rect 6846 18417 7123 18432
tri 7123 18417 7138 18432 sw
rect 6846 18411 7448 18417
rect 6846 18377 6972 18411
rect 7006 18377 7058 18411
rect 7092 18377 7144 18411
rect 7178 18377 7230 18411
rect 7264 18377 7316 18411
rect 7350 18377 7402 18411
rect 7436 18377 7448 18411
rect 6846 18371 7448 18377
rect 6846 18358 7125 18371
tri 7125 18358 7138 18371 nw
rect 6846 18136 7104 18358
tri 7104 18337 7125 18358 nw
tri 7465 18284 7476 18295 se
rect 7476 18284 7576 18506
tri 7442 18261 7465 18284 se
rect 7465 18261 7576 18284
rect 7132 18255 7576 18261
rect 7132 18221 7144 18255
rect 7178 18221 7222 18255
rect 7256 18221 7299 18255
rect 7333 18221 7376 18255
rect 7410 18221 7453 18255
rect 7487 18221 7530 18255
rect 7564 18221 7576 18255
rect 7132 18215 7576 18221
rect 7618 19172 7624 19206
rect 7658 19172 7664 19206
rect 7618 19132 7664 19172
rect 7618 19098 7624 19132
rect 7658 19098 7664 19132
rect 7618 19058 7664 19098
rect 7618 19024 7624 19058
rect 7658 19024 7664 19058
rect 7618 18984 7664 19024
rect 7618 18950 7624 18984
rect 7658 18950 7664 18984
rect 7618 18910 7664 18950
rect 7618 18876 7624 18910
rect 7658 18876 7664 18910
rect 7618 18836 7664 18876
rect 7618 18802 7624 18836
rect 7658 18802 7664 18836
rect 7618 18762 7664 18802
rect 7618 18728 7624 18762
rect 7658 18728 7664 18762
rect 7618 18688 7664 18728
rect 7618 18654 7624 18688
rect 7658 18654 7664 18688
rect 7618 18614 7664 18654
rect 7618 18580 7624 18614
rect 7658 18580 7664 18614
rect 7618 18540 7664 18580
rect 7618 18506 7624 18540
rect 7658 18506 7664 18540
rect 7618 18466 7664 18506
rect 7618 18432 7624 18466
rect 7658 18432 7664 18466
rect 7618 18392 7664 18432
rect 7618 18358 7624 18392
rect 7658 18358 7664 18392
rect 7618 18323 7664 18358
rect 7710 19272 7716 19306
rect 7750 19272 7756 19306
rect 7710 19234 7756 19272
rect 7710 19200 7716 19234
rect 7750 19200 7756 19234
rect 8631 19481 8683 19487
rect 8631 19417 8683 19429
rect 7710 19162 7756 19200
rect 7710 19128 7716 19162
rect 7750 19128 7756 19162
rect 7710 19090 7756 19128
rect 8551 19219 8603 19225
rect 8551 19155 8603 19167
rect 7710 19056 7716 19090
rect 7750 19056 7756 19090
rect 7710 19018 7756 19056
rect 7710 18984 7716 19018
rect 7750 18984 7756 19018
rect 7710 18946 7756 18984
rect 7710 18912 7716 18946
rect 7750 18912 7756 18946
rect 7710 18874 7756 18912
rect 7710 18840 7716 18874
rect 7750 18840 7756 18874
rect 7710 18802 7756 18840
rect 7710 18768 7716 18802
rect 7750 18768 7756 18802
rect 7710 18730 7756 18768
rect 7710 18696 7716 18730
rect 7750 18696 7756 18730
rect 7710 18658 7756 18696
rect 7710 18624 7716 18658
rect 7750 18624 7756 18658
rect 8471 19089 8523 19095
rect 8471 19025 8523 19037
rect 7710 18586 7756 18624
rect 7710 18552 7716 18586
rect 7750 18552 7756 18586
rect 7710 18514 7756 18552
rect 7710 18480 7716 18514
rect 7750 18480 7756 18514
rect 7710 18441 7756 18480
rect 7710 18407 7716 18441
rect 7750 18407 7756 18441
rect 7710 18368 7756 18407
rect 7710 18334 7716 18368
rect 7750 18334 7756 18368
tri 7664 18323 7670 18329 sw
rect 7618 18318 7670 18323
rect 7618 18317 7624 18318
rect 7658 18317 7670 18318
rect 7618 18253 7670 18265
tri 7602 18188 7618 18204 se
rect 7618 18195 7670 18201
rect 7618 18188 7664 18195
tri 7664 18189 7670 18195 nw
rect 7710 18295 7756 18334
rect 7710 18261 7716 18295
rect 7750 18261 7756 18295
rect 7710 18222 7756 18261
rect 8391 18625 8443 18631
rect 8391 18561 8443 18573
tri 7584 18170 7602 18188 se
rect 7602 18170 7664 18188
tri 7552 18139 7583 18170 se
rect 7583 18139 7624 18170
tri 7104 18136 7107 18139 sw
tri 7549 18136 7552 18139 se
rect 7552 18136 7624 18139
rect 7658 18136 7664 18170
rect 6846 18115 7107 18136
tri 7107 18115 7128 18136 sw
tri 7531 18118 7549 18136 se
rect 7549 18118 7664 18136
rect 7710 18188 7716 18222
rect 7750 18188 7756 18222
rect 7710 18149 7756 18188
tri 7528 18115 7531 18118 se
rect 7531 18115 7602 18118
tri 7602 18115 7605 18118 nw
rect 7710 18115 7716 18149
rect 7750 18115 7756 18149
rect 6846 18105 7128 18115
tri 7128 18105 7138 18115 sw
tri 7524 18111 7528 18115 se
rect 7528 18111 7592 18115
rect 7524 18105 7592 18111
tri 7592 18105 7602 18115 nw
rect 6846 18099 7448 18105
rect 6846 18065 6972 18099
rect 7006 18065 7058 18099
rect 7092 18065 7144 18099
rect 7178 18065 7230 18099
rect 7264 18065 7316 18099
rect 7350 18065 7402 18099
rect 7436 18065 7448 18099
rect 6846 18059 7448 18065
rect 6846 18052 7131 18059
tri 7131 18052 7138 18059 nw
rect 6846 18042 7121 18052
tri 7121 18042 7131 18052 nw
rect 6846 18040 7119 18042
tri 7119 18040 7121 18042 nw
rect 6846 17857 7104 18040
tri 7104 18025 7119 18040 nw
tri 7510 17969 7524 17983 se
rect 7524 17969 7576 18105
tri 7576 18089 7592 18105 nw
rect 7710 18076 7756 18115
tri 7509 17968 7510 17969 se
rect 7510 17968 7576 17969
tri 7490 17949 7509 17968 se
rect 7509 17949 7576 17968
rect 7132 17943 7576 17949
rect 7132 17909 7144 17943
rect 7178 17909 7222 17943
rect 7256 17909 7299 17943
rect 7333 17909 7376 17943
rect 7410 17909 7453 17943
rect 7487 17909 7530 17943
rect 7564 17909 7576 17943
rect 7616 18045 7668 18052
rect 7616 17981 7668 17993
rect 7616 17922 7668 17929
rect 7710 18042 7716 18076
rect 7750 18042 7756 18076
rect 8231 18241 8283 18247
rect 8231 18177 8283 18189
rect 7710 18003 7756 18042
rect 7710 17969 7716 18003
rect 7750 17969 7756 18003
rect 7710 17930 7756 17969
rect 7132 17903 7576 17909
rect 7710 17896 7716 17930
rect 7750 17896 7756 17930
tri 7104 17857 7120 17873 sw
rect 7710 17857 7756 17896
rect 6846 17839 7120 17857
tri 7120 17839 7138 17857 sw
rect 6846 17833 7576 17839
rect 6846 17799 6972 17833
rect 7006 17799 7052 17833
rect 7086 17799 7132 17833
rect 7166 17799 7212 17833
rect 7246 17799 7292 17833
rect 7326 17799 7372 17833
rect 7406 17799 7451 17833
rect 7485 17799 7530 17833
rect 7564 17799 7576 17833
rect 6846 17793 7576 17799
rect 7710 17823 7716 17857
rect 7750 17823 7756 17857
rect 6846 17784 7129 17793
tri 7129 17784 7138 17793 nw
rect 6846 17776 7121 17784
tri 7121 17776 7129 17784 nw
rect 7618 17776 7664 17788
rect 6846 17711 7104 17776
tri 7104 17759 7121 17776 nw
rect 7618 17742 7624 17776
rect 7658 17742 7664 17776
tri 7104 17711 7110 17717 sw
tri 7612 17711 7618 17717 se
rect 7618 17711 7664 17742
rect 6846 17683 7110 17711
tri 7110 17683 7138 17711 sw
tri 7584 17683 7612 17711 se
rect 7612 17683 7664 17711
rect 6846 17680 7664 17683
rect 6846 17677 7624 17680
rect 6846 17643 7116 17677
rect 7150 17643 7194 17677
rect 7228 17643 7271 17677
rect 7305 17643 7348 17677
rect 7382 17643 7425 17677
rect 7459 17643 7502 17677
rect 7536 17646 7624 17677
rect 7658 17646 7664 17680
rect 7536 17643 7664 17646
rect 6846 17637 7664 17643
rect 6846 17604 7105 17637
tri 7105 17604 7138 17637 nw
tri 7584 17604 7617 17637 ne
rect 7617 17604 7664 17637
rect 6846 17549 7104 17604
tri 7104 17603 7105 17604 nw
tri 7617 17603 7618 17604 ne
rect 7618 17583 7664 17604
tri 7104 17549 7116 17561 sw
rect 7618 17549 7624 17583
rect 7658 17549 7664 17583
rect 6846 17531 7116 17549
tri 7116 17531 7134 17549 sw
rect 7618 17537 7664 17549
rect 7710 17784 7756 17823
rect 7710 17750 7716 17784
rect 7750 17750 7756 17784
rect 7710 17711 7756 17750
rect 7710 17677 7716 17711
rect 7750 17677 7756 17711
rect 7710 17638 7756 17677
rect 7710 17604 7716 17638
rect 7750 17604 7756 17638
rect 7710 17565 7756 17604
rect 7710 17531 7716 17565
rect 7750 17531 7756 17565
rect 6846 17527 7134 17531
tri 7134 17527 7138 17531 sw
rect 6846 17521 7448 17527
rect 6846 17487 6972 17521
rect 7006 17487 7058 17521
rect 7092 17487 7144 17521
rect 7178 17487 7230 17521
rect 7264 17487 7316 17521
rect 7350 17487 7402 17521
rect 7436 17487 7448 17521
rect 6846 17481 7448 17487
rect 7710 17492 7756 17531
rect 6846 17468 7125 17481
tri 7125 17468 7138 17481 nw
rect 7618 17468 7664 17480
rect 6846 17330 7104 17468
tri 7104 17447 7125 17468 nw
rect 7618 17434 7624 17468
rect 7658 17434 7664 17468
rect 7618 17394 7664 17434
rect 6846 17278 6847 17330
rect 6899 17278 6915 17330
rect 6967 17278 6983 17330
rect 7035 17278 7051 17330
rect 7103 17278 7104 17330
rect 7132 17365 7576 17371
rect 7132 17331 7144 17365
rect 7178 17331 7222 17365
rect 7256 17331 7299 17365
rect 7333 17331 7376 17365
rect 7410 17331 7453 17365
rect 7487 17331 7530 17365
rect 7564 17331 7576 17365
rect 7132 17325 7576 17331
tri 7442 17319 7448 17325 ne
rect 7448 17319 7576 17325
tri 7448 17291 7476 17319 ne
rect 6846 17263 7104 17278
rect 6846 17211 6847 17263
rect 6899 17211 6915 17263
rect 6967 17211 6983 17263
rect 7035 17211 7051 17263
rect 7103 17244 7104 17263
tri 7104 17244 7109 17249 sw
rect 7103 17215 7109 17244
tri 7109 17215 7138 17244 sw
rect 7103 17211 7448 17215
rect 6846 17209 7448 17211
rect 6846 17196 6972 17209
rect 7006 17196 7058 17209
rect 7092 17196 7144 17209
rect 6846 17144 6847 17196
rect 6899 17144 6915 17196
rect 6967 17175 6972 17196
rect 6967 17144 6983 17175
rect 7035 17144 7051 17196
rect 7103 17175 7144 17196
rect 7178 17175 7230 17209
rect 7264 17175 7316 17209
rect 7350 17175 7402 17209
rect 7436 17175 7448 17209
rect 7103 17169 7448 17175
rect 7103 17144 7104 17169
rect 6846 17129 7104 17144
tri 7104 17135 7138 17169 nw
rect 6846 17077 6847 17129
rect 6899 17077 6915 17129
rect 6967 17077 6983 17129
rect 7035 17077 7051 17129
rect 7103 17077 7104 17129
rect 6846 17062 7104 17077
rect 6846 17010 6847 17062
rect 6899 17010 6915 17062
rect 6967 17010 6983 17062
rect 7035 17010 7051 17062
rect 7103 17010 7104 17062
tri 7443 17060 7476 17093 se
rect 7476 17076 7576 17319
rect 7476 17060 7524 17076
tri 7442 17059 7443 17060 se
rect 7443 17059 7524 17060
rect 7132 17053 7524 17059
rect 7132 17019 7144 17053
rect 7178 17019 7222 17053
rect 7256 17019 7299 17053
rect 7333 17019 7376 17053
rect 7410 17019 7453 17053
rect 7487 17024 7524 17053
rect 7487 17019 7530 17024
rect 7564 17019 7576 17024
rect 7132 17013 7576 17019
rect 6846 16994 7104 17010
rect 6846 16942 6847 16994
rect 6899 16942 6915 16994
rect 6967 16942 6983 16994
rect 7035 16942 7051 16994
rect 7103 16942 7104 16994
tri 7442 16985 7470 17013 ne
rect 7470 17012 7576 17013
rect 7470 16985 7524 17012
tri 7470 16981 7474 16985 ne
rect 7474 16981 7524 16985
tri 7474 16979 7476 16981 ne
rect 6846 16936 7104 16942
rect 7476 16960 7524 16981
tri 7104 16936 7105 16937 sw
rect 6846 16910 7105 16936
tri 7105 16910 7131 16936 sw
rect 6846 16908 7131 16910
tri 7131 16908 7133 16910 sw
rect 6846 16903 7133 16908
tri 7133 16903 7138 16908 sw
rect 6846 16897 7448 16903
rect 6846 16863 6972 16897
rect 7006 16863 7058 16897
rect 7092 16863 7144 16897
rect 7178 16863 7230 16897
rect 7264 16863 7316 16897
rect 7350 16863 7402 16897
rect 7436 16863 7448 16897
rect 6846 16857 7448 16863
rect 6846 16835 7116 16857
tri 7116 16835 7138 16857 nw
rect 6846 16610 7104 16835
tri 7104 16823 7116 16835 nw
tri 7455 16760 7476 16781 se
rect 7476 16760 7576 16960
tri 7442 16747 7455 16760 se
rect 7455 16747 7576 16760
rect 7132 16741 7576 16747
rect 7132 16707 7144 16741
rect 7178 16707 7222 16741
rect 7256 16707 7299 16741
rect 7333 16707 7376 16741
rect 7410 16707 7453 16741
rect 7487 16707 7530 16741
rect 7564 16707 7576 16741
rect 7132 16701 7576 16707
tri 7442 16685 7458 16701 ne
rect 7458 16685 7576 16701
tri 7458 16667 7476 16685 ne
tri 7104 16610 7119 16625 sw
rect 6846 16593 7119 16610
tri 7119 16593 7136 16610 sw
rect 6846 16591 7136 16593
tri 7136 16591 7138 16593 sw
rect 6846 16585 7448 16591
rect 6846 16551 6972 16585
rect 7006 16551 7058 16585
rect 7092 16551 7144 16585
rect 7178 16551 7230 16585
rect 7264 16551 7316 16585
rect 7350 16551 7402 16585
rect 7436 16551 7448 16585
rect 6846 16545 7448 16551
rect 6846 16535 7128 16545
tri 7128 16535 7138 16545 nw
rect 6846 16317 7104 16535
tri 7104 16511 7128 16535 nw
tri 7467 16460 7476 16469 se
rect 7476 16460 7576 16685
tri 7443 16436 7467 16460 se
rect 7467 16436 7576 16460
tri 7442 16435 7443 16436 se
rect 7443 16435 7576 16436
rect 7132 16429 7576 16435
rect 7132 16395 7144 16429
rect 7178 16395 7222 16429
rect 7256 16395 7299 16429
rect 7333 16395 7376 16429
rect 7410 16395 7453 16429
rect 7487 16395 7530 16429
rect 7564 16395 7576 16429
rect 7132 16389 7576 16395
rect 7618 17360 7624 17394
rect 7658 17360 7664 17394
rect 7618 17319 7664 17360
rect 7618 17285 7624 17319
rect 7658 17285 7664 17319
rect 7618 17244 7664 17285
rect 7618 17210 7624 17244
rect 7658 17210 7664 17244
rect 7618 17169 7664 17210
rect 7618 17135 7624 17169
rect 7658 17135 7664 17169
rect 7618 17094 7664 17135
rect 7618 17060 7624 17094
rect 7658 17060 7664 17094
rect 7618 17019 7664 17060
rect 7618 16985 7624 17019
rect 7658 16985 7664 17019
rect 7618 16944 7664 16985
rect 7618 16910 7624 16944
rect 7658 16910 7664 16944
rect 7618 16869 7664 16910
rect 7618 16835 7624 16869
rect 7658 16835 7664 16869
rect 7618 16794 7664 16835
rect 7618 16760 7624 16794
rect 7658 16760 7664 16794
rect 7618 16721 7664 16760
rect 7710 17458 7716 17492
rect 7750 17458 7756 17492
rect 7710 17419 7756 17458
rect 7710 17385 7716 17419
rect 7750 17385 7756 17419
rect 7710 17346 7756 17385
rect 7710 17312 7716 17346
rect 7750 17312 7756 17346
rect 7710 17273 7756 17312
rect 7710 17239 7716 17273
rect 7750 17239 7756 17273
rect 7710 17200 7756 17239
rect 7710 17166 7716 17200
rect 7750 17166 7756 17200
rect 7710 17127 7756 17166
rect 7710 17093 7716 17127
rect 7750 17093 7756 17127
rect 7710 17054 7756 17093
rect 7710 17020 7716 17054
rect 7750 17020 7756 17054
rect 7710 16981 7756 17020
rect 7710 16947 7716 16981
rect 7750 16947 7756 16981
rect 7710 16908 7756 16947
rect 7710 16874 7716 16908
rect 7750 16874 7756 16908
rect 7710 16835 7756 16874
rect 7710 16801 7716 16835
rect 7750 16801 7756 16835
rect 7710 16762 7756 16801
rect 7710 16728 7716 16762
rect 7750 16728 7756 16762
tri 7664 16721 7670 16727 sw
rect 7618 16719 7670 16721
rect 7618 16715 7624 16719
rect 7658 16715 7670 16719
rect 7618 16651 7670 16663
rect 7618 16593 7670 16599
rect 7618 16569 7664 16593
tri 7664 16587 7670 16593 nw
rect 7710 16689 7756 16728
rect 7710 16655 7716 16689
rect 7750 16655 7756 16689
rect 7710 16616 7756 16655
rect 7618 16535 7624 16569
rect 7658 16535 7664 16569
rect 7618 16494 7664 16535
rect 7618 16460 7624 16494
rect 7658 16460 7664 16494
rect 7618 16419 7664 16460
rect 7618 16385 7624 16419
rect 7658 16385 7664 16419
tri 7603 16363 7618 16378 se
rect 7618 16363 7664 16385
tri 7584 16344 7603 16363 se
rect 7603 16344 7664 16363
tri 7556 16317 7583 16344 se
rect 7583 16317 7624 16344
tri 6846 16310 6853 16317 ne
rect 6853 16310 7104 16317
tri 7552 16313 7556 16317 se
rect 7556 16313 7624 16317
tri 7104 16310 7107 16313 sw
tri 7549 16310 7552 16313 se
rect 7552 16310 7624 16313
rect 7658 16310 7664 16344
tri 6853 16290 6873 16310 ne
rect 6873 16290 7107 16310
tri 7107 16290 7127 16310 sw
tri 7531 16292 7549 16310 se
rect 7549 16292 7664 16310
rect 7710 16582 7716 16616
rect 7750 16582 7756 16616
rect 7710 16543 7756 16582
rect 7710 16509 7716 16543
rect 7750 16509 7756 16543
rect 7710 16470 7756 16509
rect 7710 16436 7716 16470
rect 7750 16436 7756 16470
rect 7710 16397 7756 16436
rect 7710 16363 7716 16397
rect 7750 16363 7756 16397
rect 7710 16324 7756 16363
tri 7529 16290 7531 16292 se
rect 7531 16290 7603 16292
tri 7603 16290 7605 16292 nw
rect 7710 16290 7716 16324
rect 7750 16290 7756 16324
tri 6873 16273 6890 16290 ne
rect 6890 16279 7127 16290
tri 7127 16279 7138 16290 sw
tri 7524 16285 7529 16290 se
rect 7529 16285 7592 16290
rect 7524 16279 7592 16285
tri 7592 16279 7603 16290 nw
rect 6890 16273 7448 16279
tri 6890 16239 6924 16273 ne
rect 6924 16239 6972 16273
rect 7006 16239 7058 16273
rect 7092 16239 7144 16273
rect 7178 16239 7230 16273
rect 7264 16239 7316 16273
rect 7350 16239 7402 16273
rect 7436 16239 7448 16273
tri 6924 16228 6935 16239 ne
rect 6935 16233 7448 16239
rect 6935 16228 7133 16233
tri 7133 16228 7138 16233 nw
rect 2654 16222 2706 16228
rect 2654 16158 2706 16170
rect 1648 15716 1700 15722
rect 1648 15652 1700 15664
rect 736 14139 742 14191
rect 794 14139 806 14191
rect 858 14139 864 14191
tri 731 3475 736 3480 se
rect 736 3475 764 14139
tri 764 14105 798 14139 nw
rect 1011 14059 1017 14111
rect 1069 14059 1081 14111
rect 1133 14059 1139 14111
tri 1077 14042 1094 14059 ne
rect 1094 14042 1139 14059
tri 1094 14037 1099 14042 ne
rect 1099 14037 1139 14042
tri 1099 14025 1111 14037 ne
tri 710 3454 731 3475 se
rect 731 3454 764 3475
tri 702 3446 710 3454 se
rect 710 3446 764 3454
rect 564 3418 764 3446
rect 792 13701 844 13707
rect 792 13637 844 13649
rect 792 13579 844 13585
rect 792 13561 826 13579
tri 826 13561 844 13579 nw
rect 564 3399 607 3418
tri 607 3399 626 3418 nw
tri 789 3399 792 3402 se
rect 792 3399 820 13561
tri 820 13555 826 13561 nw
rect 931 13497 983 13503
rect 931 13433 983 13445
tri 898 13376 931 13409 se
rect 931 13376 983 13381
tri 897 13375 898 13376 se
rect 898 13375 983 13376
tri 555 444 564 453 se
rect 564 444 592 3399
tri 592 3384 607 3399 nw
tri 774 3384 789 3399 se
rect 789 3384 820 3399
tri 758 3368 774 3384 se
rect 774 3368 820 3384
tri 540 429 555 444 se
rect 555 429 592 444
rect 540 423 592 429
rect 627 3340 820 3368
rect 848 13314 983 13375
rect 848 13304 900 13314
tri 900 13304 910 13314 nw
rect 848 13299 895 13304
tri 895 13299 900 13304 nw
rect 627 3323 672 3340
tri 672 3323 689 3340 nw
rect 627 3308 657 3323
tri 657 3308 672 3323 nw
rect 627 476 655 3308
tri 655 3306 657 3308 nw
tri 846 3306 848 3308 se
rect 848 3306 876 13299
tri 876 13280 895 13299 nw
tri 1105 13257 1111 13263 se
rect 1111 13257 1139 14037
rect 1648 14042 1700 15600
rect 2204 14139 2210 14191
rect 2262 14139 2274 14191
rect 2326 14139 2332 14191
tri 2246 14105 2280 14139 ne
tri 1700 14042 1723 14065 sw
rect 1648 14037 1723 14042
tri 1723 14037 1728 14042 sw
rect 1648 14031 1728 14037
tri 1728 14031 1734 14037 sw
tri 1081 13233 1105 13257 se
rect 1105 13233 1139 13257
tri 1080 13232 1081 13233 se
rect 1081 13232 1139 13233
tri 1077 13229 1080 13232 se
rect 1080 13229 1139 13232
tri 838 3298 846 3306 se
rect 846 3298 876 3306
tri 814 3274 838 3298 se
rect 838 3274 876 3298
rect 697 3246 876 3274
rect 904 13201 1139 13229
rect 1184 14025 1236 14031
rect 1648 13979 1654 14031
rect 1706 13979 1718 14031
rect 1770 13979 1776 14031
rect 1184 13961 1236 13973
rect 1184 13903 1236 13909
rect 1184 13898 1231 13903
tri 1231 13898 1236 13903 nw
rect 1184 13891 1224 13898
tri 1224 13891 1231 13898 nw
rect 904 13191 956 13201
tri 956 13191 966 13201 nw
rect 904 13186 951 13191
tri 951 13186 956 13191 nw
rect 697 3228 741 3246
tri 741 3228 759 3246 nw
rect 697 3213 726 3228
tri 726 3213 741 3228 nw
tri 889 3213 904 3228 se
rect 904 3213 932 13186
tri 932 13167 951 13186 nw
tri 1175 13061 1184 13070 se
rect 1184 13061 1212 13891
tri 1212 13879 1224 13891 nw
rect 1579 13795 1585 13847
rect 1637 13795 1649 13847
rect 1701 13795 1707 13847
rect 1299 13196 1351 13202
rect 1299 13132 1351 13144
rect 1299 13074 1351 13080
tri 1299 13070 1303 13074 ne
rect 1303 13070 1351 13074
tri 1303 13061 1312 13070 ne
rect 1312 13061 1351 13070
tri 1164 13050 1175 13061 se
rect 1175 13050 1212 13061
tri 1312 13050 1323 13061 ne
tri 1157 13043 1164 13050 se
rect 1164 13043 1212 13050
tri 1150 13036 1157 13043 se
rect 1157 13036 1212 13043
rect 697 558 725 3213
tri 725 3212 726 3213 nw
tri 888 3212 889 3213 se
rect 889 3212 932 3213
tri 884 3208 888 3212 se
rect 888 3208 932 3212
tri 870 3194 884 3208 se
rect 884 3194 932 3208
rect 771 3166 932 3194
rect 960 13008 1212 13036
rect 960 13003 1017 13008
tri 1017 13003 1022 13008 nw
rect 960 12988 1002 13003
tri 1002 12988 1017 13003 nw
rect 771 3143 810 3166
tri 810 3143 833 3166 nw
rect 771 3142 809 3143
tri 809 3142 810 3143 nw
tri 959 3142 960 3143 se
rect 960 3142 988 12988
tri 988 12974 1002 12988 nw
tri 1310 12337 1323 12350 se
rect 1323 12337 1351 13061
tri 1298 12325 1310 12337 se
rect 1310 12325 1351 12337
tri 1289 12316 1298 12325 se
rect 1298 12316 1351 12325
rect 771 632 799 3142
tri 799 3132 809 3142 nw
tri 949 3132 959 3142 se
rect 959 3132 988 3142
tri 926 3109 949 3132 se
rect 949 3109 988 3132
rect 827 3081 988 3109
rect 1072 12288 1351 12316
rect 1379 13131 1429 13183
rect 1481 13131 1493 13183
rect 1545 13131 1551 13183
rect 1379 13117 1427 13131
tri 1427 13117 1441 13131 nw
rect 1379 13105 1415 13117
tri 1415 13105 1427 13117 nw
rect 1072 12269 1115 12288
tri 1115 12269 1134 12288 nw
rect 1072 12265 1111 12269
tri 1111 12265 1115 12269 nw
tri 1375 12265 1379 12269 se
rect 1379 12265 1407 13105
tri 1407 13097 1415 13105 nw
rect 1491 12825 1543 12831
rect 1491 12761 1543 12773
rect 1491 12703 1543 12709
tri 1491 12679 1515 12703 ne
rect 1072 12263 1109 12265
tri 1109 12263 1111 12265 nw
tri 1373 12263 1375 12265 se
rect 1375 12263 1407 12265
rect 827 3061 869 3081
tri 869 3061 889 3081 nw
rect 827 740 855 3061
tri 855 3047 869 3061 nw
tri 1048 2952 1072 2976 se
rect 1072 2952 1100 12263
tri 1100 12254 1109 12263 nw
tri 1364 12254 1373 12263 se
rect 1373 12254 1407 12263
tri 1345 12235 1364 12254 se
rect 1364 12235 1407 12254
tri 1046 2950 1048 2952 se
rect 1048 2950 1100 2952
tri 1039 2943 1046 2950 se
rect 1046 2943 1100 2950
tri 1038 2942 1039 2943 se
rect 1039 2942 1100 2943
rect 957 2914 1100 2942
rect 1128 12207 1407 12235
rect 1435 12565 1487 12571
rect 1435 12501 1487 12513
rect 1435 12443 1487 12449
rect 1128 12203 1186 12207
tri 1186 12203 1190 12207 nw
rect 1128 12176 1159 12203
tri 1159 12176 1186 12203 nw
rect 957 2909 1014 2914
tri 1014 2909 1019 2914 nw
rect 957 2896 1001 2909
tri 1001 2896 1014 2909 nw
rect 957 927 985 2896
tri 985 2880 1001 2896 nw
tri 1112 2880 1128 2896 se
rect 1128 2880 1156 12176
tri 1156 12173 1159 12176 nw
tri 1432 12173 1435 12176 se
rect 1435 12173 1463 12443
tri 1463 12419 1487 12443 nw
tri 1428 12169 1432 12173 se
rect 1432 12169 1463 12173
tri 1426 12167 1428 12169 se
rect 1428 12167 1463 12169
tri 1401 12142 1426 12167 se
rect 1426 12142 1463 12167
tri 1109 2877 1112 2880 se
rect 1112 2877 1156 2880
tri 1099 2867 1109 2877 se
rect 1109 2867 1156 2877
tri 1094 2862 1099 2867 se
rect 1099 2862 1156 2867
rect 1032 2834 1156 2862
rect 1184 12114 1463 12142
rect 1184 12095 1227 12114
tri 1227 12095 1246 12114 nw
rect 1184 12085 1217 12095
tri 1217 12085 1227 12095 nw
rect 1032 2833 1093 2834
tri 1093 2833 1094 2834 nw
rect 1032 2830 1090 2833
tri 1090 2830 1093 2833 nw
rect 1032 2822 1082 2830
tri 1082 2822 1090 2830 nw
rect 1032 1000 1060 2822
tri 1060 2800 1082 2822 nw
tri 1162 2800 1184 2822 se
rect 1184 2800 1212 12085
tri 1212 12080 1217 12085 nw
tri 1509 12073 1515 12079 se
rect 1515 12073 1543 12703
tri 1487 12051 1509 12073 se
rect 1509 12051 1543 12073
tri 1481 12045 1487 12051 se
rect 1487 12045 1543 12051
tri 1158 2796 1162 2800 se
rect 1162 2796 1212 2800
tri 1153 2791 1158 2796 se
rect 1158 2791 1212 2796
tri 1150 2788 1153 2791 se
rect 1153 2788 1212 2791
rect 1104 2760 1212 2788
rect 1240 12017 1543 12045
rect 1104 2757 1163 2760
tri 1163 2757 1166 2760 nw
rect 1104 2750 1156 2757
tri 1156 2750 1163 2757 nw
rect 1104 1073 1132 2750
tri 1132 2726 1156 2750 nw
rect 1240 1180 1268 12017
tri 1268 11983 1302 12017 nw
tri 1545 11920 1579 11954 se
rect 1579 11920 1607 13795
tri 1607 13761 1641 13795 nw
rect 1296 11892 1607 11920
rect 1635 13666 1641 13718
rect 1693 13666 1705 13718
rect 1757 13666 1763 13718
rect 1635 13635 1666 13666
tri 1666 13635 1697 13666 nw
rect 1296 1252 1324 11892
tri 1324 11858 1358 11892 nw
tri 1621 11858 1635 11872 se
rect 1635 11858 1663 13635
tri 1663 13632 1666 13635 nw
tri 1601 11838 1621 11858 se
rect 1621 11838 1663 11858
rect 1352 11810 1663 11838
rect 1691 13371 1697 13423
rect 1749 13371 1761 13423
rect 1813 13371 1819 13423
rect 1691 13339 1721 13371
tri 1721 13339 1753 13371 nw
rect 1352 11786 1390 11810
tri 1390 11786 1414 11810 nw
tri 1685 11786 1691 11792 se
rect 1691 11786 1719 13339
tri 1719 13337 1721 13339 nw
rect 1775 13291 1781 13343
rect 1833 13291 1845 13343
rect 1897 13291 1903 13343
rect 1775 13280 1826 13291
tri 1826 13280 1837 13291 nw
rect 1775 13265 1811 13280
tri 1811 13265 1826 13280 nw
rect 1352 11782 1386 11786
tri 1386 11782 1390 11786 nw
tri 1681 11782 1685 11786 se
rect 1685 11782 1719 11786
rect 1352 1438 1380 11782
tri 1380 11776 1386 11782 nw
tri 1675 11776 1681 11782 se
rect 1681 11776 1719 11782
tri 1657 11758 1675 11776 se
rect 1675 11758 1719 11776
rect 1408 11730 1719 11758
tri 1747 13117 1775 13145 se
rect 1775 13117 1803 13265
tri 1803 13257 1811 13265 nw
rect 1747 13089 1803 13117
rect 1747 13077 1791 13089
tri 1791 13077 1803 13089 nw
rect 1903 13211 1937 13263
rect 1989 13211 2001 13263
rect 2053 13211 2059 13263
rect 1903 13201 1955 13211
tri 1955 13201 1965 13211 nw
rect 1903 13191 1945 13201
tri 1945 13191 1955 13201 nw
rect 1903 13186 1940 13191
tri 1940 13186 1945 13191 nw
rect 1408 11704 1444 11730
tri 1444 11704 1470 11730 nw
rect 1408 11697 1437 11704
tri 1437 11697 1444 11704 nw
tri 1740 11697 1747 11704 se
rect 1747 11697 1775 13077
tri 1775 13061 1791 13077 nw
tri 1896 13043 1903 13050 se
rect 1903 13043 1931 13186
tri 1931 13177 1940 13186 nw
tri 2273 13043 2280 13050 se
rect 2280 13043 2332 14139
tri 1877 13024 1896 13043 se
rect 1896 13024 1931 13043
tri 2254 13024 2273 13043 se
rect 2273 13024 2332 13043
tri 1869 13016 1877 13024 se
rect 1877 13016 1931 13024
tri 2246 13016 2254 13024 se
rect 2254 13016 2332 13024
rect 1408 1545 1436 11697
tri 1436 11696 1437 11697 nw
tri 1739 11696 1740 11697 se
rect 1740 11696 1775 11697
tri 1713 11670 1739 11696 se
rect 1739 11670 1775 11696
rect 1464 11642 1775 11670
rect 1803 12988 1931 13016
rect 1803 12969 1846 12988
tri 1846 12969 1865 12988 nw
rect 1803 12964 1841 12969
tri 1841 12964 1846 12969 nw
rect 2180 12964 2186 13016
rect 2238 12964 2274 13016
rect 2326 12964 2332 13016
rect 1464 11618 1502 11642
tri 1502 11618 1526 11642 nw
rect 1464 1807 1492 11618
tri 1492 11608 1502 11618 nw
tri 1793 11608 1803 11618 se
rect 1803 11608 1831 12964
tri 1831 12954 1841 12964 nw
tri 1792 11607 1793 11608 se
rect 1793 11607 1831 11608
tri 1769 11584 1792 11607 se
rect 1792 11584 1831 11607
rect 1520 11556 1831 11584
rect 1859 12835 1865 12887
rect 1917 12835 1929 12887
rect 1981 12835 1987 12887
rect 1520 2008 1548 11556
tri 1548 11522 1582 11556 nw
tri 1825 11468 1859 11502 se
rect 1859 11468 1887 12835
tri 1887 12801 1921 12835 nw
rect 2654 12773 2706 16106
rect 6818 16222 6870 16228
tri 6935 16219 6944 16228 ne
rect 6944 16219 7124 16228
tri 7124 16219 7133 16228 nw
rect 6818 16158 6870 16170
rect 5837 14865 5889 15229
tri 6742 15227 6744 15229 se
tri 6738 15223 6742 15227 se
rect 6742 15223 6744 15227
rect 6738 15217 6790 15223
rect 6738 15139 6790 15165
rect 6738 15060 6790 15087
rect 6738 14981 6790 15008
rect 6738 14923 6790 14929
tri 6738 14917 6744 14923 ne
rect 5977 14195 5983 14247
rect 6035 14195 6065 14247
rect 6117 14195 6147 14247
rect 6199 14195 6228 14247
rect 6280 14195 6309 14247
rect 6361 14195 6367 14247
rect 2955 14139 2961 14191
rect 3013 14139 3027 14191
rect 3079 14139 3085 14191
rect 5977 14151 6367 14195
rect 5977 14099 5983 14151
rect 6035 14099 6065 14151
rect 6117 14099 6147 14151
rect 6199 14099 6228 14151
rect 6280 14099 6309 14151
rect 6361 14099 6367 14151
tri 6796 14137 6818 14159 se
rect 6818 14137 6870 16106
rect 6944 16217 7122 16219
tri 7122 16217 7124 16219 nw
rect 6944 16216 7121 16217
tri 7121 16216 7122 16217 nw
rect 6944 16032 7104 16216
tri 7104 16199 7121 16216 nw
tri 7511 16144 7524 16157 se
rect 7524 16144 7576 16279
tri 7576 16263 7592 16279 nw
rect 7710 16251 7756 16290
tri 7490 16123 7511 16144 se
rect 7511 16123 7576 16144
rect 7132 16117 7576 16123
rect 7132 16083 7144 16117
rect 7178 16083 7222 16117
rect 7256 16083 7299 16117
rect 7333 16083 7376 16117
rect 7410 16083 7453 16117
rect 7487 16083 7530 16117
rect 7564 16083 7576 16117
rect 7615 16222 7667 16228
rect 7615 16158 7667 16170
rect 7615 16098 7667 16106
rect 7710 16217 7716 16251
rect 7750 16217 7756 16251
rect 7710 16178 7756 16217
rect 7710 16144 7716 16178
rect 7750 16144 7756 16178
rect 7710 16105 7756 16144
rect 7132 16077 7576 16083
rect 7710 16071 7716 16105
rect 7750 16071 7756 16105
tri 7104 16032 7119 16047 sw
rect 7710 16032 7756 16071
rect 6944 16013 7119 16032
tri 7119 16013 7138 16032 sw
rect 6944 16007 7576 16013
rect 6944 15973 6972 16007
rect 7006 15973 7052 16007
rect 7086 15973 7132 16007
rect 7166 15973 7212 16007
rect 7246 15973 7292 16007
rect 7326 15973 7372 16007
rect 7406 15973 7451 16007
rect 7485 15973 7530 16007
rect 7564 15973 7576 16007
rect 6944 15967 7576 15973
rect 7710 15998 7716 16032
rect 7750 15998 7756 16032
rect 6944 15962 7133 15967
tri 7133 15962 7138 15967 nw
rect 6944 15959 7130 15962
tri 7130 15959 7133 15962 nw
rect 6944 15950 7121 15959
tri 7121 15950 7130 15959 nw
rect 7618 15950 7664 15962
rect 6944 15886 7104 15950
tri 7104 15933 7121 15950 nw
rect 7618 15916 7624 15950
rect 7658 15916 7664 15950
tri 7104 15886 7109 15891 sw
tri 7613 15886 7618 15891 se
rect 7618 15886 7664 15916
rect 6944 15861 7109 15886
tri 7109 15861 7134 15886 sw
tri 7588 15861 7613 15886 se
rect 7613 15861 7664 15886
rect 6944 15857 7134 15861
tri 7134 15857 7138 15861 sw
tri 7584 15857 7588 15861 se
rect 7588 15857 7624 15861
rect 6944 15851 7624 15857
rect 6944 15817 7116 15851
rect 7150 15817 7194 15851
rect 7228 15817 7271 15851
rect 7305 15817 7348 15851
rect 7382 15817 7425 15851
rect 7459 15817 7502 15851
rect 7536 15827 7624 15851
rect 7658 15827 7664 15861
rect 7536 15817 7664 15827
rect 6944 15811 7664 15817
rect 6944 15779 7106 15811
tri 7106 15779 7138 15811 nw
tri 7584 15779 7616 15811 ne
rect 7616 15779 7664 15811
rect 6944 15726 7104 15779
tri 7104 15777 7106 15779 nw
tri 7616 15777 7618 15779 ne
rect 7618 15772 7664 15779
rect 7618 15738 7624 15772
rect 7658 15738 7664 15772
tri 7104 15726 7113 15735 sw
rect 7618 15726 7664 15738
rect 7710 15959 7756 15998
rect 7710 15925 7716 15959
rect 7750 15925 7756 15959
rect 7710 15886 7756 15925
rect 7710 15852 7716 15886
rect 7750 15852 7756 15886
rect 7710 15813 7756 15852
rect 7710 15779 7716 15813
rect 7750 15779 7756 15813
rect 7710 15740 7756 15779
rect 6944 15706 7113 15726
tri 7113 15706 7133 15726 sw
rect 7710 15706 7716 15740
rect 7750 15706 7756 15740
rect 6944 15701 7133 15706
tri 7133 15701 7138 15706 sw
rect 6944 15695 7448 15701
rect 6944 15661 6972 15695
rect 7006 15661 7058 15695
rect 7092 15661 7144 15695
rect 7178 15661 7230 15695
rect 7264 15661 7316 15695
rect 7350 15661 7402 15695
rect 7436 15661 7448 15695
rect 6944 15655 7448 15661
rect 7710 15667 7756 15706
rect 6944 15633 7116 15655
tri 7116 15633 7138 15655 nw
rect 6944 15630 7113 15633
tri 7113 15630 7116 15633 nw
rect 7618 15630 7664 15642
rect 6944 15414 7104 15630
tri 7104 15621 7113 15630 nw
rect 7476 15581 7576 15598
tri 7457 15560 7476 15579 se
rect 7476 15560 7508 15581
tri 7453 15556 7457 15560 se
rect 7457 15556 7508 15560
tri 7442 15545 7453 15556 se
rect 7453 15545 7508 15556
rect 7132 15539 7508 15545
rect 7560 15539 7576 15581
rect 7132 15505 7144 15539
rect 7178 15505 7222 15539
rect 7256 15505 7299 15539
rect 7333 15505 7376 15539
rect 7410 15505 7453 15539
rect 7487 15529 7508 15539
rect 7487 15517 7530 15529
rect 7487 15505 7508 15517
rect 7564 15505 7576 15539
rect 7132 15499 7508 15505
tri 7442 15487 7454 15499 ne
rect 7454 15487 7508 15499
tri 7454 15482 7459 15487 ne
rect 7459 15482 7508 15487
tri 7459 15465 7476 15482 ne
rect 7476 15465 7508 15482
rect 7560 15465 7576 15505
tri 7104 15414 7113 15423 sw
rect 6944 15408 7113 15414
tri 7113 15408 7119 15414 sw
rect 6944 15389 7119 15408
tri 7119 15389 7138 15408 sw
rect 6944 15383 7448 15389
rect 6944 15349 6972 15383
rect 7006 15349 7058 15383
rect 7092 15349 7144 15383
rect 7178 15349 7230 15383
rect 7264 15349 7316 15383
rect 7350 15349 7402 15383
rect 7436 15349 7448 15383
rect 6944 15343 7448 15349
rect 6944 15341 7136 15343
tri 7136 15341 7138 15343 nw
rect 6944 15334 7129 15341
tri 7129 15334 7136 15341 nw
rect 6944 15217 7104 15334
tri 7104 15309 7129 15334 nw
tri 7469 15260 7476 15267 se
rect 7476 15260 7576 15465
tri 7442 15233 7469 15260 se
rect 7469 15233 7576 15260
rect 6996 15165 7052 15217
rect 7132 15227 7576 15233
rect 7132 15193 7144 15227
rect 7178 15193 7222 15227
rect 7256 15193 7299 15227
rect 7333 15193 7376 15227
rect 7410 15193 7453 15227
rect 7487 15193 7530 15227
rect 7564 15193 7576 15227
rect 7132 15187 7576 15193
tri 7442 15186 7443 15187 ne
rect 7443 15186 7576 15187
rect 6944 15139 7104 15165
tri 7443 15153 7476 15186 ne
rect 6996 15087 7052 15139
rect 6944 15078 7104 15087
tri 7104 15078 7137 15111 sw
rect 6944 15077 7137 15078
tri 7137 15077 7138 15078 sw
rect 6944 15071 7448 15077
rect 6944 15060 6972 15071
rect 7006 15060 7058 15071
rect 7092 15060 7144 15071
rect 7006 15037 7052 15060
rect 7104 15037 7144 15060
rect 7178 15037 7230 15071
rect 7264 15037 7316 15071
rect 7350 15037 7402 15071
rect 7436 15037 7448 15071
rect 6996 15008 7052 15037
rect 7104 15031 7448 15037
rect 7104 15008 7111 15031
rect 6944 15004 7111 15008
tri 7111 15004 7138 15031 nw
rect 6944 14981 7104 15004
tri 7104 14997 7111 15004 nw
rect 6996 14929 7052 14981
tri 7451 14930 7476 14955 se
rect 7476 14930 7576 15186
rect 6944 14782 7104 14929
tri 7444 14923 7451 14930 se
rect 7451 14923 7576 14930
tri 7442 14921 7444 14923 se
rect 7444 14921 7576 14923
rect 7132 14915 7576 14921
rect 7132 14881 7144 14915
rect 7178 14881 7222 14915
rect 7256 14881 7299 14915
rect 7333 14881 7376 14915
rect 7410 14881 7453 14915
rect 7487 14881 7530 14915
rect 7564 14881 7576 14915
rect 7132 14875 7576 14881
tri 7442 14865 7452 14875 ne
rect 7452 14865 7576 14875
tri 7452 14856 7461 14865 ne
rect 7461 14856 7576 14865
tri 7461 14841 7476 14856 ne
tri 7104 14782 7121 14799 sw
rect 6944 14765 7121 14782
tri 7121 14765 7138 14782 sw
rect 6944 14759 7448 14765
rect 6944 14725 6972 14759
rect 7006 14725 7058 14759
rect 7092 14725 7144 14759
rect 7178 14725 7230 14759
rect 7264 14725 7316 14759
rect 7350 14725 7402 14759
rect 7436 14725 7448 14759
rect 6944 14719 7448 14725
rect 6944 14708 7127 14719
tri 7127 14708 7138 14719 nw
rect 6944 14484 7104 14708
tri 7104 14685 7127 14708 nw
tri 7467 14634 7476 14643 se
rect 7476 14634 7576 14856
tri 7444 14611 7467 14634 se
rect 7467 14611 7576 14634
tri 7442 14609 7444 14611 se
rect 7444 14609 7576 14611
rect 7132 14603 7576 14609
rect 7132 14569 7144 14603
rect 7178 14569 7222 14603
rect 7256 14569 7299 14603
rect 7333 14569 7376 14603
rect 7410 14569 7453 14603
rect 7487 14569 7530 14603
rect 7564 14569 7576 14603
rect 7132 14563 7576 14569
rect 7618 15596 7624 15630
rect 7658 15596 7664 15630
rect 7618 15556 7664 15596
rect 7618 15522 7624 15556
rect 7658 15522 7664 15556
rect 7618 15482 7664 15522
rect 7618 15448 7624 15482
rect 7658 15448 7664 15482
rect 7618 15408 7664 15448
rect 7618 15374 7624 15408
rect 7658 15374 7664 15408
rect 7618 15334 7664 15374
rect 7618 15300 7624 15334
rect 7658 15300 7664 15334
rect 7618 15260 7664 15300
rect 7618 15226 7624 15260
rect 7658 15226 7664 15260
rect 7618 15186 7664 15226
rect 7618 15152 7624 15186
rect 7658 15152 7664 15186
rect 7618 15112 7664 15152
rect 7618 15078 7624 15112
rect 7658 15078 7664 15112
rect 7618 15038 7664 15078
rect 7618 15004 7624 15038
rect 7658 15004 7664 15038
rect 7618 14964 7664 15004
rect 7618 14930 7624 14964
rect 7658 14930 7664 14964
rect 7618 14890 7664 14930
rect 7618 14876 7624 14890
rect 7658 14882 7664 14890
rect 7710 15633 7716 15667
rect 7750 15633 7756 15667
rect 7710 15594 7756 15633
rect 7710 15560 7716 15594
rect 7750 15560 7756 15594
rect 7710 15521 7756 15560
rect 7710 15487 7716 15521
rect 7750 15487 7756 15521
rect 7710 15448 7756 15487
rect 7710 15414 7716 15448
rect 7750 15414 7756 15448
rect 7710 15375 7756 15414
rect 7710 15341 7716 15375
rect 7750 15341 7756 15375
rect 7710 15302 7756 15341
rect 7710 15268 7716 15302
rect 7750 15268 7756 15302
rect 7710 15229 7756 15268
rect 7710 15195 7716 15229
rect 7750 15195 7756 15229
rect 7710 15156 7756 15195
rect 7710 15122 7716 15156
rect 7750 15122 7756 15156
rect 7710 15083 7756 15122
rect 7710 15049 7716 15083
rect 7750 15049 7756 15083
rect 7710 15010 7756 15049
rect 7710 14976 7716 15010
rect 7750 14976 7756 15010
rect 7710 14937 7756 14976
rect 7710 14903 7716 14937
rect 7750 14903 7756 14937
tri 7664 14882 7670 14888 sw
rect 7658 14876 7670 14882
rect 7618 14816 7670 14824
rect 7618 14812 7624 14816
rect 7658 14812 7670 14816
rect 7618 14754 7670 14760
rect 7618 14742 7664 14754
tri 7664 14748 7670 14754 nw
rect 7710 14864 7756 14903
rect 7710 14830 7716 14864
rect 7750 14830 7756 14864
rect 7710 14791 7756 14830
rect 7710 14757 7716 14791
rect 7750 14757 7756 14791
rect 7618 14708 7624 14742
rect 7658 14708 7664 14742
rect 7618 14668 7664 14708
rect 7618 14634 7624 14668
rect 7658 14634 7664 14668
rect 7618 14593 7664 14634
rect 7618 14559 7624 14593
rect 7658 14559 7664 14593
tri 7604 14538 7618 14552 se
rect 7618 14538 7664 14559
tri 7584 14518 7604 14538 se
rect 7604 14518 7664 14538
tri 7552 14487 7583 14518 se
rect 7583 14487 7624 14518
tri 7104 14484 7107 14487 sw
tri 7549 14484 7552 14487 se
rect 7552 14484 7624 14487
rect 7658 14484 7664 14518
rect 6944 14465 7107 14484
tri 7107 14465 7126 14484 sw
tri 7531 14466 7549 14484 se
rect 7549 14466 7664 14484
rect 7710 14718 7756 14757
rect 7710 14684 7716 14718
rect 7750 14684 7756 14718
rect 7710 14645 7756 14684
rect 7710 14611 7716 14645
rect 7750 14611 7756 14645
rect 7710 14572 7756 14611
rect 7710 14538 7716 14572
rect 7750 14538 7756 14572
rect 7710 14499 7756 14538
tri 7530 14465 7531 14466 se
rect 7531 14465 7604 14466
tri 7604 14465 7605 14466 nw
rect 7710 14465 7716 14499
rect 7750 14465 7756 14499
rect 6944 14453 7126 14465
tri 7126 14453 7138 14465 sw
tri 7524 14459 7530 14465 se
rect 7530 14459 7592 14465
rect 7524 14453 7592 14459
tri 7592 14453 7604 14465 nw
rect 6944 14447 7448 14453
rect 6944 14413 6972 14447
rect 7006 14413 7058 14447
rect 7092 14413 7144 14447
rect 7178 14413 7230 14447
rect 7264 14413 7316 14447
rect 7350 14413 7402 14447
rect 7436 14413 7448 14447
rect 6944 14407 7448 14413
rect 6944 14403 7134 14407
tri 7134 14403 7138 14407 nw
rect 6944 14392 7123 14403
tri 7123 14392 7134 14403 nw
rect 6944 14390 7121 14392
tri 7121 14390 7123 14392 nw
rect 6944 14248 7104 14390
tri 7104 14373 7121 14390 nw
tri 7512 14319 7524 14331 se
rect 7524 14319 7576 14453
tri 7576 14437 7592 14453 nw
rect 7710 14426 7756 14465
tri 7511 14318 7512 14319 se
rect 7512 14318 7576 14319
tri 7490 14297 7511 14318 se
rect 7511 14297 7576 14318
rect 7132 14291 7576 14297
rect 7132 14257 7144 14291
rect 7178 14257 7222 14291
rect 7256 14257 7299 14291
rect 7333 14257 7376 14291
rect 7410 14257 7453 14291
rect 7487 14257 7530 14291
rect 7564 14257 7576 14291
rect 7615 14411 7667 14417
rect 7615 14356 7624 14359
rect 7658 14356 7667 14359
rect 7615 14347 7667 14356
rect 7615 14284 7624 14295
rect 7658 14284 7667 14295
rect 7615 14272 7667 14284
rect 7710 14392 7716 14426
rect 7750 14392 7756 14426
rect 7710 14353 7756 14392
rect 7710 14319 7716 14353
rect 7750 14319 7756 14353
rect 7710 14280 7756 14319
rect 7132 14251 7576 14257
rect 7710 14246 7716 14280
rect 7750 14246 7756 14280
rect 7710 14234 7756 14246
rect 7910 18045 7962 18051
rect 7910 17981 7962 17993
rect 7910 15792 7962 17929
rect 7910 15728 7962 15740
tri 6793 14134 6796 14137 se
rect 6796 14134 6867 14137
tri 6867 14134 6870 14137 nw
rect 7191 14143 7197 14195
rect 7249 14143 7263 14195
rect 7315 14143 7329 14195
rect 7381 14143 7394 14195
rect 7446 14143 7452 14195
rect 5977 14076 6367 14099
tri 6742 14083 6793 14134 se
rect 6793 14116 6849 14134
tri 6849 14116 6867 14134 nw
rect 7191 14125 7452 14143
rect 6793 14083 6815 14116
tri 6367 14076 6374 14083 sw
tri 6741 14082 6742 14083 se
rect 6742 14082 6815 14083
tri 6815 14082 6849 14116 nw
tri 7157 14082 7191 14116 se
rect 7191 14082 7197 14125
rect 6741 14076 6809 14082
tri 6809 14076 6815 14082 nw
rect 7015 14076 7197 14082
rect 5977 14055 6374 14076
rect 5977 14003 5983 14055
rect 6035 14003 6065 14055
rect 6117 14003 6147 14055
rect 6199 14003 6228 14055
rect 6280 14003 6309 14055
rect 6361 14049 6374 14055
tri 6374 14049 6401 14076 sw
rect 6361 14037 6461 14049
rect 6361 14003 6364 14037
rect 6398 14003 6461 14037
rect 5977 13991 6426 14003
tri 6426 13991 6438 14003 nw
rect 5977 13985 6420 13991
tri 6420 13985 6426 13991 nw
rect 5977 13979 6414 13985
tri 6414 13979 6420 13985 nw
rect 6661 13979 6713 13991
rect 5977 13964 6404 13979
tri 6404 13969 6414 13979 nw
rect 5977 13930 6364 13964
rect 6398 13930 6404 13964
rect 6661 13945 6670 13979
rect 6704 13945 6713 13979
rect 5977 13891 6404 13930
rect 6501 13930 6553 13936
tri 6500 13926 6501 13927 se
tri 6494 13920 6500 13926 se
rect 6500 13920 6501 13926
tri 6472 13898 6494 13920 se
rect 6494 13898 6501 13920
tri 6467 13893 6472 13898 se
rect 6472 13893 6501 13898
rect 5977 13857 6364 13891
rect 6398 13857 6404 13891
rect 3336 13795 3342 13847
rect 3394 13795 3406 13847
rect 3458 13795 3920 13847
tri 3834 13783 3846 13795 ne
rect 3846 13783 3920 13795
tri 3846 13773 3856 13783 ne
rect 3856 13773 3920 13783
tri 3856 13761 3868 13773 ne
rect 3868 13743 3920 13773
rect 5977 13817 6404 13857
tri 6553 13920 6559 13926 sw
rect 6553 13898 6559 13920
tri 6559 13898 6581 13920 sw
rect 6661 13898 6713 13945
rect 6553 13893 6581 13898
tri 6581 13893 6586 13898 sw
rect 6501 13866 6553 13878
tri 6467 13846 6468 13847 ne
rect 6468 13846 6501 13847
tri 6468 13839 6475 13846 ne
rect 6475 13839 6501 13846
tri 6475 13817 6497 13839 ne
rect 6497 13817 6501 13839
rect 5977 13783 6364 13817
rect 6398 13783 6404 13817
tri 6497 13813 6501 13817 ne
rect 6661 13864 6670 13898
rect 6704 13864 6713 13898
rect 6553 13846 6585 13847
tri 6585 13846 6586 13847 nw
rect 6553 13839 6578 13846
tri 6578 13839 6585 13846 nw
rect 6553 13817 6556 13839
tri 6556 13817 6578 13839 nw
rect 6661 13817 6713 13864
tri 6553 13814 6556 13817 nw
rect 6501 13808 6553 13814
rect 5977 13761 6404 13783
rect 6661 13783 6670 13817
rect 6704 13783 6713 13817
tri 6404 13761 6414 13771 sw
rect 5977 13749 6414 13761
tri 6414 13749 6426 13761 sw
tri 3920 13743 3926 13749 sw
rect 5977 13743 6426 13749
rect 3329 13666 3335 13718
rect 3387 13666 3399 13718
rect 3451 13666 3750 13718
rect 3868 13715 3926 13743
tri 3926 13715 3954 13743 sw
rect 3868 13669 3920 13715
rect 5977 13709 6364 13743
rect 6398 13739 6426 13743
tri 6426 13739 6436 13749 sw
rect 6398 13737 6436 13739
tri 6436 13737 6438 13739 sw
rect 6398 13709 6461 13737
rect 5977 13691 6461 13709
rect 6661 13735 6713 13783
rect 6661 13701 6670 13735
rect 6704 13701 6713 13735
rect 5977 13669 6412 13691
rect 5977 13635 6364 13669
rect 6398 13665 6412 13669
tri 6412 13665 6438 13691 nw
rect 6398 13635 6404 13665
tri 6404 13657 6412 13665 nw
rect 6661 13657 6713 13701
rect 5977 13595 6404 13635
rect 6501 13621 6553 13627
tri 6500 13614 6501 13615 se
tri 6494 13608 6500 13614 se
rect 6500 13608 6501 13614
rect 5977 13561 6364 13595
rect 6398 13561 6404 13595
tri 6467 13581 6494 13608 se
rect 6494 13581 6501 13608
tri 3199 13522 3214 13537 sw
tri 3152 13521 3153 13522 se
tri 3134 13503 3152 13521 se
rect 3152 13503 3153 13521
rect 3199 13521 3214 13522
tri 3214 13521 3215 13522 sw
rect 5977 13521 6404 13561
tri 6553 13608 6559 13614 sw
rect 6553 13581 6559 13608
tri 6559 13581 6586 13608 sw
rect 6661 13593 6713 13605
rect 6501 13557 6553 13569
tri 6467 13522 6480 13535 ne
rect 6480 13522 6501 13535
rect 3199 13503 3215 13521
tri 3215 13503 3233 13521 sw
rect 3134 13451 3140 13503
rect 3192 13451 3204 13503
rect 3256 13451 3262 13503
rect 5977 13487 6364 13521
rect 6398 13487 6404 13521
tri 6480 13520 6482 13522 ne
rect 6482 13520 6501 13522
tri 6482 13513 6489 13520 ne
rect 6489 13513 6501 13520
tri 6489 13503 6499 13513 ne
rect 6499 13505 6501 13513
rect 6661 13537 6670 13541
rect 6704 13537 6713 13541
rect 6553 13520 6571 13535
tri 6571 13520 6586 13535 nw
rect 6553 13513 6564 13520
tri 6564 13513 6571 13520 nw
rect 6499 13503 6553 13505
tri 6499 13501 6501 13503 ne
rect 6501 13499 6553 13503
tri 6553 13502 6564 13513 nw
rect 5977 13455 6404 13487
rect 6661 13489 6713 13537
tri 6404 13455 6408 13459 sw
rect 6661 13455 6670 13489
rect 6704 13455 6713 13489
rect 5977 13448 6408 13455
tri 6408 13448 6415 13455 sw
rect 5977 13447 6415 13448
tri 5949 13413 5977 13441 se
rect 5977 13413 6364 13447
rect 6398 13441 6415 13447
tri 6415 13441 6422 13448 sw
rect 6661 13443 6713 13455
rect 6398 13425 6422 13441
tri 6422 13425 6438 13441 sw
rect 6398 13413 6461 13425
tri 5946 13410 5949 13413 se
rect 5949 13410 6461 13413
tri 5943 13407 5946 13410 se
rect 5946 13407 6461 13410
rect 5977 13379 6461 13407
rect 5977 13376 6435 13379
tri 6435 13376 6438 13379 nw
rect 5977 13373 6428 13376
rect 5977 13354 6364 13373
rect 2817 13339 6364 13354
rect 6398 13369 6428 13373
tri 6428 13369 6435 13376 nw
rect 6398 13348 6407 13369
tri 6407 13348 6428 13369 nw
rect 6661 13348 6713 13360
rect 6398 13339 6404 13348
tri 6404 13345 6407 13348 nw
rect 2817 13325 6404 13339
rect 5977 13299 6404 13325
rect 6661 13314 6670 13348
rect 6704 13314 6713 13348
rect 5977 13275 6364 13299
tri 5943 13265 5953 13275 ne
rect 5953 13265 6364 13275
rect 6398 13265 6404 13299
tri 6497 13297 6501 13301 se
rect 6501 13297 6553 13301
tri 6553 13297 6557 13301 sw
tri 6496 13296 6497 13297 se
rect 6497 13296 6557 13297
tri 6557 13296 6558 13297 sw
tri 6475 13275 6496 13296 se
rect 6496 13295 6558 13296
rect 6496 13275 6501 13295
tri 6469 13269 6475 13275 se
rect 6475 13269 6501 13275
tri 5953 13241 5977 13265 ne
rect 5977 13225 6404 13265
rect 3134 13183 3262 13217
rect 3134 13131 3140 13183
rect 3192 13131 3204 13183
rect 3256 13131 3262 13183
rect 3329 13141 3335 13193
rect 3387 13141 3399 13193
rect 3451 13141 3457 13193
rect 3134 13086 3262 13131
tri 3371 13117 3395 13141 ne
rect 3395 13117 3457 13141
tri 3395 13107 3405 13117 ne
rect 3405 13043 3457 13117
rect 5977 13191 6364 13225
rect 6398 13191 6404 13225
rect 6553 13275 6558 13295
tri 6558 13275 6579 13296 sw
rect 6553 13269 6579 13275
tri 6579 13269 6585 13275 sw
rect 6501 13231 6553 13243
tri 6467 13217 6473 13223 ne
rect 6473 13217 6501 13223
tri 6473 13194 6496 13217 ne
rect 6496 13194 6501 13217
rect 5977 13151 6404 13191
tri 6496 13189 6501 13194 ne
rect 6661 13267 6713 13314
rect 6661 13233 6670 13267
rect 6704 13233 6713 13267
rect 6553 13194 6557 13223
tri 6557 13194 6586 13223 nw
rect 6661 13198 6713 13233
tri 6553 13190 6557 13194 nw
rect 6501 13173 6553 13179
rect 5977 13117 6364 13151
rect 6398 13141 6404 13151
tri 6404 13141 6410 13147 sw
rect 6398 13140 6410 13141
tri 6410 13140 6411 13141 sw
rect 6398 13121 6411 13140
tri 6411 13121 6430 13140 sw
rect 6661 13134 6713 13146
rect 6398 13117 6430 13121
rect 5977 13113 6430 13117
tri 6430 13113 6438 13121 sw
rect 5977 13077 6461 13113
tri 3457 13043 3464 13050 sw
rect 5977 13043 6364 13077
rect 6398 13067 6461 13077
rect 6661 13071 6670 13082
rect 6704 13071 6713 13082
rect 6398 13050 6421 13067
tri 6421 13050 6438 13067 nw
rect 6398 13048 6419 13050
tri 6419 13048 6421 13050 nw
rect 6398 13043 6404 13048
rect 3405 13024 3464 13043
tri 3464 13024 3483 13043 sw
rect 3405 13016 3483 13024
tri 3483 13016 3491 13024 sw
rect 2862 12964 2868 13016
rect 2920 12964 2934 13016
rect 2986 12964 2992 13016
rect 3405 12962 3806 13016
rect 3868 12967 3920 13013
rect 5977 13003 6404 13043
tri 6404 13033 6419 13048 nw
rect 6661 13024 6713 13071
rect 5977 12969 6364 13003
rect 6398 12969 6404 13003
rect 6501 13004 6553 13010
tri 6496 12984 6501 12989 se
rect 3868 12950 3937 12967
tri 3937 12950 3954 12967 nw
rect 3868 12943 3930 12950
tri 3930 12943 3937 12950 nw
tri 3842 12895 3868 12921 se
rect 3868 12895 3920 12943
tri 3920 12933 3930 12943 nw
tri 3834 12887 3842 12895 se
rect 3842 12887 3920 12895
rect 3336 12835 3342 12887
rect 3394 12835 3406 12887
rect 3458 12835 3920 12887
rect 5977 12929 6404 12969
tri 6479 12967 6496 12984 se
rect 6496 12967 6501 12984
tri 6469 12957 6479 12967 se
rect 6479 12957 6501 12967
rect 5977 12895 6364 12929
rect 6398 12895 6404 12929
rect 6661 12990 6670 13024
rect 6704 12990 6713 13024
tri 6553 12984 6558 12989 sw
rect 6553 12967 6558 12984
tri 6558 12967 6575 12984 sw
rect 6553 12957 6575 12967
tri 6575 12957 6585 12967 sw
rect 6501 12940 6553 12952
tri 6472 12909 6474 12911 ne
rect 6474 12909 6501 12911
tri 6474 12899 6484 12909 ne
rect 6484 12899 6501 12909
rect 5977 12855 6404 12895
tri 6484 12887 6496 12899 ne
rect 6496 12888 6501 12899
rect 6661 12943 6713 12990
rect 6553 12909 6580 12911
tri 6580 12909 6582 12911 nw
rect 6661 12909 6670 12943
rect 6704 12909 6713 12943
rect 6553 12899 6570 12909
tri 6570 12899 6580 12909 nw
rect 6496 12887 6553 12888
tri 6496 12882 6501 12887 ne
rect 6501 12882 6553 12887
tri 6553 12882 6570 12899 nw
rect 2654 12709 2706 12721
rect 2654 12651 2706 12657
rect 5977 12821 6364 12855
rect 6398 12827 6404 12855
rect 6661 12861 6713 12909
tri 6404 12827 6412 12835 sw
rect 6661 12827 6670 12861
rect 6704 12827 6713 12861
rect 6398 12826 6412 12827
tri 6412 12826 6413 12827 sw
rect 6398 12821 6413 12826
rect 5977 12801 6413 12821
tri 6413 12801 6438 12826 sw
rect 6661 12815 6713 12827
rect 5977 12781 6461 12801
rect 5977 12747 6364 12781
rect 6398 12755 6461 12781
rect 6741 12787 6793 14076
tri 6793 14060 6809 14076 nw
rect 7015 14042 7027 14076
rect 7061 14042 7106 14076
rect 7140 14042 7185 14076
rect 7249 14073 7263 14125
rect 7315 14073 7329 14125
rect 7381 14073 7394 14125
rect 7446 14082 7452 14125
tri 7452 14082 7486 14116 sw
rect 7446 14076 7855 14082
rect 7446 14073 7530 14076
rect 7219 14055 7530 14073
rect 7015 14036 7197 14042
tri 7157 14025 7168 14036 ne
rect 7168 14025 7197 14036
tri 7168 14019 7174 14025 ne
rect 7174 14019 7197 14025
tri 7174 14002 7191 14019 ne
rect 7191 14003 7197 14019
rect 7249 14003 7263 14055
rect 7315 14003 7329 14055
rect 7381 14003 7394 14055
rect 7446 14042 7530 14055
rect 7564 14042 7629 14076
rect 7663 14042 7855 14076
rect 7446 14036 7855 14042
rect 7446 14019 7469 14036
tri 7469 14019 7486 14036 nw
tri 7775 14019 7792 14036 ne
rect 7792 14019 7855 14036
rect 7446 14003 7452 14019
tri 7188 13957 7191 13960 se
rect 7191 13957 7452 14003
tri 7452 14002 7469 14019 nw
tri 7792 14002 7809 14019 ne
rect 7809 13985 7815 14019
rect 7849 13985 7855 14019
tri 7176 13945 7188 13957 se
rect 7188 13945 7452 13957
tri 7157 13926 7176 13945 se
rect 7176 13926 7304 13945
rect 7015 13920 7304 13926
rect 6827 13880 6873 13892
rect 7015 13886 7027 13920
rect 7061 13886 7169 13920
rect 7203 13911 7304 13920
rect 7338 13931 7452 13945
tri 7452 13931 7481 13960 sw
rect 7809 13931 7855 13985
rect 7338 13926 7481 13931
tri 7481 13926 7486 13931 sw
rect 7338 13920 7675 13926
rect 7338 13911 7423 13920
rect 7203 13886 7423 13911
rect 7457 13886 7526 13920
rect 7560 13886 7629 13920
rect 7663 13886 7675 13920
rect 7015 13880 7675 13886
rect 7809 13897 7815 13931
rect 7849 13897 7855 13931
rect 6827 13846 6833 13880
rect 6867 13846 6873 13880
tri 7157 13873 7164 13880 ne
rect 7164 13873 7451 13880
tri 7164 13846 7191 13873 ne
rect 6827 13801 6873 13846
rect 7191 13839 7304 13873
rect 7338 13839 7451 13873
tri 7451 13846 7485 13880 nw
rect 7707 13850 7767 13856
tri 6873 13801 6876 13804 sw
tri 7188 13801 7191 13804 se
rect 7191 13801 7451 13839
rect 6827 13773 6876 13801
rect 6827 13739 6833 13773
rect 6867 13770 6876 13773
tri 6876 13770 6907 13801 sw
tri 7157 13770 7188 13801 se
rect 7188 13770 7304 13801
rect 6867 13767 7304 13770
rect 7338 13770 7451 13801
tri 7451 13770 7485 13804 sw
rect 7707 13798 7715 13850
rect 7707 13786 7767 13798
rect 7338 13767 7675 13770
rect 6867 13764 7675 13767
rect 6867 13739 6959 13764
rect 6827 13730 6959 13739
rect 6993 13730 7035 13764
rect 7069 13730 7110 13764
rect 7144 13730 7185 13764
rect 7219 13730 7521 13764
rect 7555 13730 7629 13764
rect 7663 13730 7675 13764
rect 6827 13729 7675 13730
rect 6827 13724 7304 13729
rect 6827 13695 6878 13724
tri 6878 13695 6907 13724 nw
tri 7157 13695 7186 13724 ne
rect 7186 13695 7304 13724
rect 7338 13724 7675 13729
rect 7707 13734 7715 13786
rect 7338 13720 7481 13724
tri 7481 13720 7485 13724 nw
rect 7338 13695 7451 13720
rect 6827 13665 6873 13695
tri 6873 13690 6878 13695 nw
tri 7186 13690 7191 13695 ne
rect 6827 13631 6833 13665
rect 6867 13631 6873 13665
rect 7191 13657 7451 13695
tri 7451 13690 7481 13720 nw
rect 6827 13619 6873 13631
tri 7166 13623 7191 13648 se
rect 7191 13623 7304 13657
rect 7338 13631 7451 13657
tri 7451 13631 7468 13648 sw
rect 7338 13623 7468 13631
tri 7162 13619 7166 13623 se
rect 7166 13619 7468 13623
tri 7157 13614 7162 13619 se
rect 7162 13614 7468 13619
tri 7468 13614 7485 13631 sw
rect 7015 13608 7675 13614
rect 6925 13571 6985 13577
rect 6827 13554 6873 13566
rect 6827 13520 6833 13554
rect 6867 13520 6873 13554
rect 6827 13482 6873 13520
rect 6827 13448 6833 13482
rect 6867 13448 6873 13482
rect 6827 13410 6873 13448
rect 6827 13376 6833 13410
rect 6867 13376 6873 13410
rect 6827 13338 6873 13376
tri 6821 13304 6827 13310 se
rect 6827 13304 6833 13338
rect 6867 13304 6873 13338
rect 6821 13298 6873 13304
rect 6821 13234 6833 13246
rect 6867 13234 6873 13246
rect 6821 13176 6833 13182
tri 6821 13170 6827 13176 ne
rect 6827 13160 6833 13176
rect 6867 13160 6873 13182
rect 6827 13121 6873 13160
rect 6827 13087 6833 13121
rect 6867 13087 6873 13121
rect 6925 13519 6933 13571
rect 7015 13574 7027 13608
rect 7061 13574 7169 13608
rect 7203 13585 7423 13608
rect 7203 13574 7304 13585
rect 7015 13568 7304 13574
tri 7157 13551 7174 13568 ne
rect 7174 13551 7304 13568
rect 7338 13574 7423 13585
rect 7457 13574 7526 13608
rect 7560 13574 7629 13608
rect 7663 13574 7675 13608
rect 7338 13568 7675 13574
rect 7338 13563 7480 13568
tri 7480 13563 7485 13568 nw
rect 7338 13551 7451 13563
tri 7174 13534 7191 13551 ne
rect 6925 13507 6985 13519
rect 6925 13455 6933 13507
rect 7191 13513 7451 13551
tri 7451 13534 7480 13563 nw
tri 6985 13479 6998 13492 sw
rect 7191 13479 7304 13513
rect 7338 13479 7451 13513
tri 7705 13490 7707 13492 se
rect 7707 13490 7767 13734
rect 7809 13843 7855 13897
rect 7809 13809 7815 13843
rect 7849 13809 7855 13843
rect 7809 13754 7855 13809
rect 7809 13720 7815 13754
rect 7849 13720 7855 13754
rect 7809 13665 7855 13720
rect 7809 13631 7815 13665
rect 7849 13631 7855 13665
rect 7809 13619 7855 13631
rect 6985 13458 6998 13479
tri 6998 13458 7019 13479 sw
rect 6985 13455 7141 13458
rect 6925 13452 7141 13455
rect 6925 13418 6937 13452
rect 6971 13418 7016 13452
rect 7050 13418 7095 13452
rect 7129 13418 7141 13452
rect 6925 13412 7141 13418
rect 7191 13441 7451 13479
tri 7673 13458 7705 13490 se
rect 7705 13458 7767 13490
rect 6925 13407 7014 13412
tri 7014 13407 7019 13412 nw
rect 7191 13407 7304 13441
rect 7338 13407 7451 13441
rect 7495 13452 7767 13458
rect 7495 13418 7507 13452
rect 7541 13418 7608 13452
rect 7642 13418 7709 13452
rect 7743 13418 7767 13452
rect 7495 13412 7767 13418
rect 6925 13383 6990 13407
tri 6990 13383 7014 13407 nw
rect 6925 13162 6985 13383
tri 6985 13378 6990 13383 nw
rect 7191 13369 7451 13407
tri 7673 13383 7702 13412 ne
rect 7702 13383 7767 13412
tri 7702 13378 7707 13383 ne
tri 7190 13335 7191 13336 se
rect 7191 13335 7304 13369
rect 7338 13335 7451 13369
tri 7165 13310 7190 13335 se
rect 7190 13310 7451 13335
tri 7451 13310 7477 13336 sw
tri 7157 13302 7165 13310 se
rect 7165 13302 7477 13310
tri 7477 13302 7485 13310 sw
rect 7015 13297 7675 13302
rect 7015 13296 7304 13297
rect 7015 13262 7027 13296
rect 7061 13262 7100 13296
rect 7134 13262 7173 13296
rect 7207 13263 7304 13296
rect 7338 13296 7675 13297
rect 7338 13263 7423 13296
rect 7207 13262 7423 13263
rect 7457 13262 7526 13296
rect 7560 13262 7629 13296
rect 7663 13262 7675 13296
rect 7015 13256 7675 13262
tri 7157 13236 7177 13256 ne
rect 7177 13236 7465 13256
tri 7465 13236 7485 13256 nw
tri 7177 13225 7188 13236 ne
rect 7188 13225 7451 13236
tri 7188 13222 7191 13225 ne
rect 7191 13191 7304 13225
rect 7338 13191 7451 13225
tri 7451 13222 7465 13236 nw
tri 6985 13162 7003 13180 sw
rect 6925 13152 7003 13162
tri 7003 13152 7013 13162 sw
rect 7191 13152 7451 13191
tri 7689 13162 7707 13180 se
rect 7707 13162 7767 13383
rect 6925 13146 7013 13152
tri 7013 13146 7019 13152 sw
rect 6925 13140 7141 13146
rect 6925 13106 6937 13140
rect 6971 13106 7016 13140
rect 7050 13106 7095 13140
rect 7129 13106 7141 13140
rect 6925 13100 7141 13106
rect 7191 13118 7304 13152
rect 7338 13118 7451 13152
tri 7673 13146 7689 13162 se
rect 7689 13146 7767 13162
rect 6827 13048 6873 13087
rect 6827 13014 6833 13048
rect 6867 13014 6873 13048
rect 7191 13079 7451 13118
rect 7493 13140 7767 13146
rect 7493 13106 7505 13140
rect 7539 13106 7607 13140
rect 7641 13106 7709 13140
rect 7743 13106 7767 13140
rect 7493 13100 7767 13106
rect 7809 13563 7855 13575
rect 7809 13529 7815 13563
rect 7849 13529 7855 13563
rect 7809 13490 7855 13529
rect 7809 13456 7815 13490
rect 7849 13456 7855 13490
rect 7809 13417 7855 13456
rect 7809 13383 7815 13417
rect 7849 13383 7855 13417
rect 7809 13344 7855 13383
rect 7809 13310 7815 13344
rect 7849 13310 7855 13344
rect 7809 13270 7855 13310
rect 7809 13236 7815 13270
rect 7849 13236 7855 13270
rect 7809 13196 7855 13236
rect 7809 13162 7815 13196
rect 7849 13162 7855 13196
rect 7809 13122 7855 13162
rect 7191 13045 7304 13079
rect 7338 13045 7451 13079
tri 7181 13014 7191 13024 se
rect 7191 13014 7451 13045
rect 7809 13088 7815 13122
rect 7849 13088 7855 13122
rect 7809 13048 7855 13088
tri 7855 13048 7861 13054 sw
rect 7809 13042 7815 13048
rect 7849 13042 7861 13048
tri 7451 13014 7461 13024 sw
rect 6827 12910 6873 13014
tri 7173 13006 7181 13014 se
rect 7181 13006 7461 13014
tri 7157 12990 7173 13006 se
rect 7173 12990 7304 13006
rect 7015 12984 7304 12990
rect 7015 12950 7027 12984
rect 7061 12950 7100 12984
rect 7134 12950 7173 12984
rect 7207 12972 7304 12984
rect 7338 12990 7461 13006
tri 7461 12990 7485 13014 sw
rect 7338 12984 7733 12990
rect 7338 12972 7439 12984
rect 7207 12950 7439 12972
rect 7473 12950 7522 12984
rect 7556 12950 7605 12984
rect 7639 12950 7687 12984
rect 7721 12950 7733 12984
rect 7015 12944 7733 12950
rect 7809 12978 7861 12990
tri 7067 12933 7078 12944 ne
rect 7078 12933 7555 12944
tri 7078 12924 7087 12933 ne
rect 7087 12924 7304 12933
tri 7087 12917 7094 12924 ne
rect 7094 12917 7304 12924
tri 6873 12910 6880 12917 sw
tri 7094 12910 7101 12917 ne
rect 6827 12899 6880 12910
tri 6880 12899 6891 12910 sw
rect 7101 12899 7304 12917
rect 7338 12924 7555 12933
tri 7555 12924 7575 12944 nw
rect 7338 12899 7541 12924
tri 7541 12910 7555 12924 nw
tri 7795 12910 7809 12924 se
rect 7809 12910 7861 12926
rect 6827 12897 6891 12899
tri 6827 12886 6838 12897 ne
rect 6838 12886 6891 12897
tri 6891 12886 6904 12899 sw
tri 6838 12874 6850 12886 ne
rect 6850 12874 7001 12886
tri 7001 12874 7013 12886 sw
rect 7101 12874 7541 12899
tri 7775 12890 7795 12910 se
rect 7795 12890 7861 12910
tri 6850 12851 6873 12874 ne
rect 6873 12869 7013 12874
tri 7013 12869 7018 12874 sw
rect 6873 12865 7018 12869
tri 7018 12865 7022 12869 sw
rect 6873 12851 7022 12865
tri 6873 12840 6884 12851 ne
rect 6884 12840 7022 12851
tri 7022 12840 7047 12865 sw
rect 7101 12840 7113 12874
rect 7147 12840 7185 12874
rect 7219 12860 7423 12874
rect 7219 12840 7304 12860
tri 6981 12830 6991 12840 ne
rect 6991 12838 7047 12840
tri 7047 12838 7049 12840 sw
rect 6991 12834 7049 12838
tri 7049 12834 7053 12838 sw
rect 7101 12834 7304 12840
rect 6991 12830 7053 12834
tri 7053 12830 7057 12834 sw
tri 6991 12826 6995 12830 ne
rect 6995 12826 7057 12830
tri 7157 12826 7165 12834 ne
rect 7165 12826 7304 12834
rect 7338 12840 7423 12860
rect 7457 12840 7495 12874
rect 7529 12840 7541 12874
tri 7603 12865 7628 12890 se
rect 7628 12865 7861 12890
rect 7338 12834 7541 12840
tri 7576 12838 7603 12865 se
rect 7603 12844 7861 12865
rect 7603 12838 7637 12844
tri 7572 12834 7576 12838 se
rect 7576 12834 7637 12838
rect 7338 12826 7451 12834
tri 6995 12820 7001 12826 ne
rect 7001 12820 7057 12826
tri 7001 12810 7011 12820 ne
tri 6793 12787 6806 12800 sw
rect 6741 12766 6806 12787
tri 6806 12766 6827 12787 sw
rect 6398 12754 6437 12755
tri 6437 12754 6438 12755 nw
rect 6741 12754 6983 12766
rect 6398 12747 6415 12754
rect 5977 12732 6415 12747
tri 6415 12732 6437 12754 nw
rect 6661 12743 6713 12749
rect 5977 12707 6404 12732
tri 6404 12721 6415 12732 nw
rect 6581 12721 6633 12727
rect 5977 12673 6364 12707
rect 6398 12673 6404 12707
rect 5977 12633 6404 12673
tri 6565 12663 6581 12679 se
rect 6581 12663 6633 12669
tri 6562 12660 6565 12663 se
rect 6565 12660 6633 12663
tri 6553 12651 6562 12660 se
rect 6562 12657 6633 12660
rect 6562 12651 6581 12657
tri 6547 12645 6553 12651 se
rect 6553 12645 6581 12651
rect 5977 12599 6364 12633
rect 6398 12599 6404 12633
rect 6741 12720 6943 12754
rect 6977 12720 6983 12754
rect 6741 12697 6983 12720
rect 6661 12679 6713 12691
tri 6903 12690 6910 12697 ne
rect 6910 12690 6983 12697
tri 6910 12682 6918 12690 ne
rect 6918 12682 6983 12690
rect 7011 12753 7057 12820
tri 7165 12800 7191 12826 ne
rect 7191 12787 7451 12826
tri 7451 12800 7485 12834 nw
tri 7571 12833 7572 12834 se
rect 7572 12833 7637 12834
tri 7637 12833 7648 12844 nw
tri 7057 12753 7068 12764 sw
rect 7191 12753 7304 12787
rect 7338 12753 7451 12787
tri 7567 12760 7571 12764 se
rect 7571 12760 7617 12833
tri 7617 12813 7637 12833 nw
tri 7871 12772 7910 12811 se
rect 7910 12772 7962 15676
rect 7011 12730 7068 12753
tri 7068 12730 7091 12753 sw
rect 7011 12724 7141 12730
rect 7011 12690 7023 12724
rect 7057 12690 7095 12724
rect 7129 12690 7141 12724
rect 7011 12684 7141 12690
rect 7191 12714 7451 12753
tri 7537 12730 7567 12760 se
rect 7567 12730 7617 12760
tri 6918 12663 6937 12682 ne
rect 6937 12648 6943 12682
rect 6977 12648 6983 12682
rect 7191 12680 7304 12714
rect 7338 12680 7451 12714
rect 7487 12724 7617 12730
rect 7487 12690 7499 12724
rect 7533 12690 7571 12724
rect 7605 12690 7617 12724
rect 7487 12684 7617 12690
rect 7659 12760 7962 12772
rect 7659 12726 7665 12760
rect 7699 12726 7962 12760
rect 7659 12698 7962 12726
rect 8148 14902 8203 14908
rect 8148 14850 8149 14902
rect 8201 14850 8203 14902
rect 8148 14812 8203 14850
rect 8148 14760 8149 14812
rect 8201 14760 8203 14812
rect 7659 12688 7705 12698
rect 7191 12653 7451 12680
rect 7659 12654 7665 12688
rect 7699 12654 7705 12688
tri 7705 12664 7739 12698 nw
rect 6937 12636 6983 12648
rect 7659 12642 7705 12654
rect 6661 12626 6670 12627
rect 6704 12626 6713 12627
rect 6661 12614 6713 12626
rect 6581 12599 6633 12605
rect 5977 12587 6404 12599
tri 7960 12539 7994 12573 se
rect 6536 12512 7995 12539
rect 6536 12460 6542 12512
rect 6594 12460 6608 12512
rect 6660 12460 6674 12512
rect 6726 12490 6740 12512
rect 6792 12490 6806 12512
rect 6858 12490 6872 12512
rect 6924 12490 6938 12512
rect 6735 12460 6740 12490
rect 6924 12460 6929 12490
rect 6990 12460 7004 12512
rect 7056 12460 7070 12512
rect 7122 12460 7136 12512
rect 7188 12490 7202 12512
rect 7254 12490 7268 12512
rect 7320 12490 7334 12512
rect 7386 12490 7400 12512
rect 7452 12490 7466 12512
rect 7191 12460 7202 12490
rect 7267 12460 7268 12490
rect 7452 12460 7461 12490
rect 7518 12460 7532 12512
rect 7584 12460 7598 12512
rect 7650 12460 7664 12512
rect 7716 12460 7729 12512
rect 7781 12460 7794 12512
rect 7846 12460 7859 12512
rect 7911 12460 7995 12512
rect 6536 12456 6548 12460
rect 6582 12456 6625 12460
rect 6659 12456 6701 12460
rect 6735 12456 6777 12460
rect 6811 12456 6853 12460
rect 6887 12456 6929 12460
rect 6963 12456 7005 12460
rect 7039 12456 7081 12460
rect 7115 12456 7157 12460
rect 7191 12456 7233 12460
rect 7267 12456 7309 12460
rect 7343 12456 7385 12460
rect 7419 12456 7461 12460
rect 7495 12456 7537 12460
rect 7571 12456 7613 12460
rect 7647 12456 7995 12460
rect 6386 12371 6432 12383
rect 6386 12337 6392 12371
rect 6426 12337 6432 12371
rect 6386 12299 6432 12337
rect 6386 12265 6392 12299
rect 6426 12265 6432 12299
rect 5187 12085 5649 12137
rect 5701 12085 5713 12137
rect 5765 12085 5771 12137
rect 5187 12073 5261 12085
tri 5261 12073 5273 12085 nw
tri 5165 12017 5187 12039 se
rect 5187 12017 5239 12073
tri 5239 12051 5261 12073 nw
tri 5153 12005 5165 12017 se
rect 5165 12005 5239 12017
rect 5187 11959 5239 12005
rect 5412 11956 5757 12008
rect 6115 11959 6121 12011
rect 6173 11959 6187 12011
rect 6239 11959 6245 12011
tri 5671 11954 5673 11956 ne
rect 5673 11954 5757 11956
tri 5673 11945 5682 11954 ne
rect 5682 11945 5757 11954
tri 5682 11922 5705 11945 ne
tri 5689 11838 5705 11854 se
rect 5705 11838 5757 11945
tri 5670 11819 5689 11838 se
rect 5689 11819 5757 11838
tri 5757 11819 5791 11853 sw
rect 5871 11837 5999 11885
rect 5670 11767 5676 11819
rect 5728 11767 5740 11819
rect 5792 11767 5798 11819
rect 5871 11785 5877 11837
rect 5929 11785 5941 11837
rect 5993 11785 5999 11837
rect 6386 11832 6432 12265
rect 6536 12371 7995 12456
rect 6536 12337 6542 12371
rect 6576 12359 7995 12371
rect 6576 12337 6798 12359
rect 6536 12325 6798 12337
rect 6832 12343 7120 12359
rect 6832 12325 6854 12343
tri 6854 12325 6872 12343 nw
tri 6924 12325 6942 12343 ne
rect 6942 12325 7020 12343
tri 7020 12325 7038 12343 nw
tri 7080 12325 7098 12343 ne
rect 7098 12325 7120 12343
rect 7154 12343 7432 12359
rect 7154 12325 7176 12343
tri 7176 12325 7194 12343 nw
tri 7392 12325 7410 12343 ne
rect 7410 12325 7432 12343
rect 7466 12343 7995 12359
rect 7466 12325 7472 12343
rect 6536 12299 6838 12325
tri 6838 12309 6854 12325 nw
tri 6942 12309 6958 12325 ne
rect 6536 12265 6542 12299
rect 6576 12265 6672 12299
rect 6706 12265 6838 12299
rect 6536 12263 6838 12265
rect 6536 12253 6798 12263
tri 6632 12229 6656 12253 ne
rect 6656 12229 6798 12253
rect 6832 12229 6838 12263
tri 6656 12219 6666 12229 ne
rect 6460 12165 6466 12217
rect 6518 12165 6530 12217
rect 6582 12165 6590 12217
rect 6460 12129 6590 12165
rect 6460 12095 6472 12129
rect 6506 12095 6544 12129
rect 6578 12095 6590 12129
rect 6460 12089 6590 12095
rect 6666 12167 6838 12229
rect 6666 12133 6672 12167
rect 6706 12133 6798 12167
rect 6832 12133 6838 12167
rect 6666 12121 6838 12133
rect 6958 12299 7004 12325
tri 7004 12309 7020 12325 nw
tri 7098 12309 7114 12325 ne
rect 6958 12265 6964 12299
rect 6998 12265 7004 12299
rect 6958 12167 7004 12265
rect 6958 12133 6964 12167
rect 6998 12133 7004 12167
rect 6958 12121 7004 12133
rect 7114 12263 7160 12325
tri 7160 12309 7176 12325 nw
tri 7410 12311 7424 12325 ne
rect 7424 12311 7472 12325
rect 7114 12229 7120 12263
rect 7154 12229 7160 12263
rect 7114 12167 7160 12229
rect 7114 12133 7120 12167
rect 7154 12133 7160 12167
rect 7114 12121 7160 12133
rect 7270 12299 7316 12311
tri 7424 12309 7426 12311 ne
rect 7270 12265 7276 12299
rect 7310 12265 7316 12299
rect 7270 12203 7316 12265
rect 7270 12169 7276 12203
rect 7310 12169 7316 12203
tri 7264 12121 7270 12127 se
rect 7270 12121 7316 12169
rect 7426 12263 7472 12311
tri 7472 12309 7506 12343 nw
tri 7704 12311 7736 12343 ne
rect 7736 12311 7995 12343
rect 7426 12229 7432 12263
rect 7466 12229 7472 12263
rect 7426 12167 7472 12229
rect 7426 12133 7432 12167
rect 7466 12133 7472 12167
tri 7316 12121 7322 12127 sw
rect 7426 12121 7472 12133
rect 7582 12299 7628 12311
tri 7736 12309 7738 12311 ne
rect 7582 12265 7588 12299
rect 7622 12265 7628 12299
rect 7582 12203 7628 12265
rect 7582 12169 7588 12203
rect 7622 12169 7628 12203
tri 7576 12121 7582 12127 se
rect 7582 12121 7628 12169
rect 6666 12120 6745 12121
tri 6745 12120 6746 12121 nw
tri 7263 12120 7264 12121 se
rect 7264 12120 7322 12121
tri 7322 12120 7323 12121 sw
tri 7575 12120 7576 12121 se
rect 7576 12120 7628 12121
rect 6666 12107 6732 12120
tri 6732 12107 6745 12120 nw
tri 7250 12107 7263 12120 se
rect 7263 12107 7323 12120
tri 7323 12107 7336 12120 sw
tri 7562 12107 7575 12120 se
rect 7575 12107 7628 12120
rect 6666 12100 6725 12107
tri 6725 12100 6732 12107 nw
tri 7243 12100 7250 12107 se
rect 7250 12100 7276 12107
rect 6666 12013 6712 12100
tri 6712 12087 6725 12100 nw
tri 7236 12093 7243 12100 se
rect 7243 12093 7276 12100
rect 6770 12041 6776 12093
rect 6828 12041 6840 12093
rect 6892 12073 7276 12093
rect 7310 12100 7336 12107
tri 7336 12100 7343 12107 sw
tri 7555 12100 7562 12107 se
rect 7562 12100 7588 12107
rect 7310 12093 7343 12100
tri 7343 12093 7350 12100 sw
tri 7548 12093 7555 12100 se
rect 7555 12093 7588 12100
rect 7310 12073 7588 12093
rect 7622 12073 7628 12107
rect 6892 12041 7628 12073
rect 7738 12299 7995 12311
rect 7738 12265 7744 12299
rect 7778 12265 7995 12299
rect 7738 12203 7995 12265
rect 7738 12169 7744 12203
rect 7778 12169 7995 12203
rect 7738 12107 7995 12169
rect 7738 12073 7744 12107
rect 7778 12073 7995 12107
rect 7738 12061 7995 12073
tri 6712 12013 6718 12019 sw
rect 6770 12013 7628 12041
tri 7960 12027 7994 12061 ne
rect 6666 11985 6718 12013
tri 6718 11985 6746 12013 sw
rect 6666 11979 7104 11985
rect 6666 11945 6724 11979
rect 6758 11945 6808 11979
rect 6842 11945 6892 11979
rect 6926 11945 6975 11979
rect 7009 11945 7058 11979
rect 7092 11945 7104 11979
rect 6666 11939 7104 11945
rect 7192 11979 7587 11985
rect 7192 11945 7204 11979
rect 7238 11945 7289 11979
rect 7323 11945 7373 11979
rect 7407 11945 7457 11979
rect 7491 11945 7541 11979
rect 7575 11945 7587 11979
tri 6432 11832 6466 11866 sw
tri 7158 11832 7192 11866 se
rect 7192 11838 7587 11945
rect 7192 11832 7465 11838
rect 6386 11786 7465 11832
rect 7517 11786 7529 11838
rect 7581 11786 7587 11838
rect 8148 11866 8203 14760
rect 8231 12972 8283 18125
rect 8311 16741 8363 16747
rect 8311 16651 8363 16689
rect 8311 13278 8363 16599
rect 8311 13214 8363 13226
rect 8311 13156 8363 13162
rect 8391 13733 8443 18509
rect 8391 13669 8443 13681
tri 8283 12972 8317 13006 sw
rect 8231 12920 8237 12972
rect 8289 12920 8301 12972
rect 8353 12920 8359 12972
rect 8391 12819 8443 13617
rect 8471 13122 8523 18973
rect 8551 13378 8603 19103
rect 8631 13733 8683 19365
rect 8711 14798 8763 19692
rect 8793 19435 8799 19487
rect 8851 19435 8863 19487
rect 8915 19435 8921 19487
rect 9005 18882 9145 18888
rect 9057 18830 9093 18882
rect 9005 18792 9145 18830
rect 9057 18740 9093 18792
rect 9005 15034 9145 18740
rect 9057 14982 9093 15034
rect 9005 14945 9145 14982
rect 9057 14893 9093 14945
rect 9385 17056 9391 17108
rect 9443 17056 9486 17108
rect 9538 17056 9544 17108
rect 9385 17006 9544 17056
rect 9385 16954 9391 17006
rect 9443 16954 9486 17006
rect 9538 16954 9544 17006
rect 9385 15059 9544 16954
rect 9385 15007 9391 15059
rect 9443 15007 9486 15059
rect 9538 15007 9544 15059
rect 9385 14991 9544 15007
rect 9385 14939 9391 14991
rect 9443 14939 9486 14991
rect 9538 14939 9544 14991
rect 9385 14938 9544 14939
rect 9005 14887 9145 14893
tri 8763 14798 8788 14823 sw
rect 8711 14746 9219 14798
rect 9271 14746 9283 14798
rect 9335 14792 9624 14798
rect 9335 14746 9572 14792
rect 8711 14740 9572 14746
rect 8711 14730 9624 14740
rect 8711 13969 8763 14730
tri 8763 14705 8788 14730 nw
tri 9165 14705 9190 14730 ne
rect 9190 14705 9353 14730
tri 9190 14696 9199 14705 ne
rect 9005 14558 9011 14610
rect 9063 14558 9087 14610
rect 9139 14558 9145 14610
rect 9199 14567 9353 14705
tri 9353 14696 9387 14730 nw
tri 9538 14696 9572 14730 ne
rect 9572 14724 9624 14730
rect 9572 14656 9624 14672
rect 9005 14528 9145 14558
rect 9005 14476 9011 14528
rect 9063 14476 9087 14528
rect 9139 14476 9145 14528
rect 9385 14541 9544 14571
tri 8763 13969 8764 13970 sw
rect 8711 13936 8764 13969
tri 8764 13936 8797 13969 sw
rect 8711 13884 8717 13936
rect 8769 13884 8781 13936
rect 8833 13884 8839 13936
rect 8631 13669 8683 13681
rect 8631 13611 8683 13617
rect 9005 13856 9145 14476
rect 9199 14241 9353 14507
rect 9251 14189 9301 14241
rect 9199 14151 9353 14189
rect 9251 14099 9301 14151
rect 9199 14061 9353 14099
rect 9251 14009 9301 14061
rect 9199 14003 9353 14009
rect 9385 14489 9391 14541
rect 9443 14489 9486 14541
rect 9538 14489 9544 14541
tri 9145 13856 9179 13890 sw
rect 9005 13804 9011 13856
rect 9063 13804 9087 13856
rect 9139 13804 9163 13856
rect 9215 13804 9221 13856
rect 8551 13314 8603 13326
rect 8551 13256 8603 13262
rect 8758 13378 8824 13384
rect 8758 13326 8763 13378
rect 8815 13326 8824 13378
rect 8758 13314 8824 13326
rect 8758 13262 8763 13314
rect 8815 13262 8824 13314
rect 8471 13058 8523 13070
rect 8471 13000 8523 13006
rect 8570 13038 8698 13044
rect 8391 12755 8443 12767
rect 8391 12697 8443 12703
rect 8622 12986 8646 13038
rect 8570 12953 8698 12986
rect 8622 12901 8646 12953
tri 8203 11866 8205 11868 sw
rect 8148 11835 8205 11866
tri 8205 11835 8236 11866 sw
rect 8148 11834 8236 11835
tri 8236 11834 8237 11835 sw
rect 5871 11755 5999 11785
rect 8148 11782 8154 11834
rect 8206 11782 8218 11834
rect 8270 11782 8276 11834
tri 6357 11730 6358 11731 sw
tri 7993 11730 7994 11731 se
rect 6357 11704 6358 11730
tri 6358 11704 6384 11730 sw
tri 7967 11704 7993 11730 se
rect 7993 11704 7994 11730
rect 6357 11697 6384 11704
tri 6384 11697 6391 11704 sw
tri 7960 11697 7967 11704 se
rect 7967 11697 7994 11704
rect 2661 11645 2667 11697
rect 2719 11645 2736 11697
rect 2788 11645 2805 11697
rect 2857 11645 2873 11697
rect 2925 11645 2941 11697
rect 2993 11645 3009 11697
rect 3061 11645 3077 11697
rect 3129 11645 3145 11697
rect 3197 11645 3213 11697
rect 3265 11645 3281 11697
rect 3333 11645 3349 11697
rect 3401 11645 3417 11697
rect 3469 11645 3485 11697
rect 3537 11645 7995 11697
rect 2661 11611 7995 11645
rect 1576 11440 1887 11468
rect 2213 11601 2265 11607
rect 2213 11537 2265 11549
rect 1576 2137 1604 11440
tri 1604 11406 1638 11440 nw
rect 2133 11433 2185 11439
tri 2099 11371 2133 11405 se
rect 2133 11371 2185 11381
rect 1639 11369 2185 11371
rect 1639 11317 2133 11369
rect 1639 11310 2185 11317
rect 1639 3994 1691 11310
tri 1691 11276 1725 11310 nw
tri 2099 11276 2133 11310 ne
rect 1802 11079 1808 11131
rect 1860 11079 1872 11131
rect 1924 11079 2073 11131
rect 1802 11075 2073 11079
rect 1639 3930 1691 3942
rect 1639 3872 1691 3878
rect 1733 11037 1785 11043
rect 1733 10973 1785 10985
rect 1733 3471 1785 10921
rect 1733 3407 1785 3419
rect 1632 2744 1684 2750
rect 1632 2680 1684 2692
rect 1632 2367 1684 2628
rect 1632 2303 1684 2315
rect 1632 2245 1684 2251
tri 1604 2137 1638 2171 sw
rect 1576 2085 1582 2137
rect 1634 2085 1646 2137
rect 1698 2085 1704 2137
tri 1618 2051 1652 2085 ne
tri 1548 2008 1572 2032 sw
rect 1520 2002 1572 2008
rect 1520 1938 1572 1950
rect 1520 1880 1572 1886
tri 1492 1807 1509 1824 sw
rect 1464 1800 1509 1807
tri 1509 1800 1516 1807 sw
rect 1464 1794 1516 1800
rect 1464 1730 1516 1742
rect 1464 1672 1516 1678
tri 1436 1545 1445 1554 sw
rect 1408 1520 1445 1545
tri 1445 1520 1470 1545 sw
rect 1408 1468 1414 1520
rect 1466 1468 1478 1520
rect 1530 1468 1536 1520
tri 1380 1438 1386 1444 sw
rect 1352 1410 1386 1438
tri 1386 1410 1414 1438 sw
rect 1352 1358 1358 1410
rect 1410 1358 1422 1410
rect 1474 1358 1480 1410
tri 1324 1252 1358 1286 sw
rect 1296 1200 1302 1252
rect 1354 1200 1366 1252
rect 1418 1200 1467 1252
tri 1268 1180 1272 1184 sw
rect 1240 1150 1272 1180
tri 1272 1150 1302 1180 sw
tri 1381 1166 1415 1200 ne
rect 1240 1098 1246 1150
rect 1298 1098 1310 1150
rect 1362 1098 1368 1150
tri 1132 1073 1152 1093 sw
rect 1104 1059 1152 1073
tri 1152 1059 1166 1073 sw
tri 1060 1000 1069 1009 sw
rect 1104 1007 1110 1059
rect 1162 1007 1174 1059
rect 1226 1007 1232 1059
rect 1032 975 1069 1000
tri 1069 975 1094 1000 sw
tri 985 927 987 929 sw
rect 957 895 987 927
tri 987 895 1019 927 sw
rect 1032 923 1038 975
rect 1090 923 1102 975
rect 1154 923 1160 975
rect 957 843 963 895
rect 1015 843 1027 895
rect 1079 843 1085 895
tri 855 740 860 745 sw
rect 827 711 860 740
tri 860 711 889 740 sw
rect 827 659 833 711
rect 885 659 897 711
rect 949 659 955 711
tri 799 632 809 642 sw
rect 771 608 809 632
tri 809 608 833 632 sw
tri 725 558 729 562 sw
rect 697 556 729 558
tri 729 556 731 558 sw
rect 771 556 910 608
rect 962 556 974 608
rect 1026 556 1032 608
rect 697 528 731 556
tri 731 528 759 556 sw
tri 655 476 657 478 sw
rect 697 476 703 528
rect 755 476 767 528
rect 819 476 1027 528
rect 627 444 657 476
tri 657 444 689 476 sw
tri 941 444 973 476 ne
rect 973 444 1027 476
rect 627 392 633 444
rect 685 392 697 444
rect 749 392 755 444
tri 973 442 975 444 ne
rect 540 359 592 371
rect 540 301 592 307
rect 282 58 334 70
rect 282 0 334 6
rect 975 0 1027 444
rect 1415 122 1467 1200
rect 1415 58 1467 70
rect 1415 0 1467 6
rect 1652 122 1704 2085
rect 1733 1866 1785 3355
rect 1813 10352 1865 10358
rect 1813 10288 1865 10300
rect 1813 2048 1865 10236
rect 2133 10247 2185 11310
rect 2213 10557 2265 11485
rect 2661 11559 2667 11611
rect 2719 11559 2736 11611
rect 2788 11559 2805 11611
rect 2857 11559 2873 11611
rect 2925 11559 2941 11611
rect 2993 11559 3009 11611
rect 3061 11559 3077 11611
rect 3129 11559 3145 11611
rect 3197 11559 3213 11611
rect 3265 11559 3281 11611
rect 3333 11559 3349 11611
rect 3401 11559 3417 11611
rect 3469 11559 3485 11611
rect 3537 11559 7995 11611
rect 2661 11465 7995 11559
tri 7960 11439 7986 11465 ne
rect 7986 11439 7994 11465
rect 2350 11433 2402 11439
tri 7986 11431 7994 11439 ne
rect 2350 11369 2402 11381
rect 2350 11311 2402 11317
tri 4968 11311 4987 11330 se
rect 4987 11314 5750 11330
tri 5750 11314 5766 11330 sw
rect 4987 11311 5766 11314
tri 4941 11284 4968 11311 se
rect 4968 11284 5766 11311
tri 5766 11284 5796 11314 sw
tri 4940 11283 4941 11284 se
rect 4941 11283 4997 11284
rect 2707 11277 2759 11283
rect 2707 11185 2759 11225
rect 2627 11117 2679 11123
rect 2627 11053 2679 11065
rect 2213 10493 2265 10505
rect 2213 10435 2265 10441
rect 2293 10515 2320 10567
rect 2372 10515 2384 10567
rect 2436 10515 2442 10567
rect 2293 10504 2368 10515
tri 2368 10504 2379 10515 nw
rect 2133 10183 2185 10195
rect 1977 10035 1983 10087
rect 2035 10035 2047 10087
rect 2099 10035 2105 10087
tri 2019 10011 2043 10035 ne
rect 2043 10011 2105 10035
tri 2043 10002 2052 10011 ne
rect 2052 10002 2105 10011
tri 2052 10001 2053 10002 ne
rect 1893 9677 1945 9683
rect 1893 9613 1945 9625
rect 1893 2744 1945 9561
rect 1893 2680 1945 2692
rect 1893 2622 1945 2628
rect 1973 9546 2025 9552
rect 1973 9482 2025 9494
rect 1973 2447 2025 9430
rect 2053 2661 2105 10002
rect 2053 2597 2105 2609
rect 2053 2539 2105 2545
tri 2130 2518 2133 2521 se
rect 2133 2518 2185 10131
rect 2213 10001 2265 10007
rect 2213 9937 2265 9949
rect 2213 2745 2265 9885
rect 2293 2877 2345 10504
tri 2345 10481 2368 10504 nw
rect 2293 2813 2345 2825
rect 2373 10453 2425 10459
rect 2373 10389 2425 10401
rect 2373 6312 2425 10337
rect 2373 6248 2425 6260
rect 2373 2928 2425 6196
rect 2627 3551 2679 11001
rect 2707 3837 2759 11133
tri 4931 11274 4940 11283 se
rect 4940 11274 4997 11283
tri 4997 11274 5007 11284 nw
tri 5730 11274 5740 11284 ne
rect 5740 11274 5796 11284
rect 3142 11118 3155 11127
rect 3142 11084 3154 11118
rect 3142 11075 3155 11084
rect 3207 11075 3219 11127
rect 3271 11075 3277 11127
rect 3343 11118 3610 11127
rect 3343 11084 3355 11118
rect 3389 11084 3437 11118
rect 3471 11084 3518 11118
rect 3552 11084 3599 11118
rect 3343 11075 3610 11084
rect 3662 11075 3674 11127
rect 3726 11118 3888 11127
rect 3726 11084 3761 11118
rect 3795 11084 3842 11118
rect 3876 11084 3888 11118
rect 3726 11075 3888 11084
rect 3971 11118 4069 11127
rect 3971 11084 3983 11118
rect 4017 11084 4065 11118
rect 3971 11075 4069 11084
rect 4121 11075 4133 11127
rect 4185 11118 4519 11127
rect 4185 11084 4229 11118
rect 4263 11084 4311 11118
rect 4345 11084 4392 11118
rect 4426 11084 4473 11118
rect 4507 11084 4519 11118
rect 4185 11075 4519 11084
rect 3081 10995 3087 11047
rect 3139 10995 3151 11047
rect 3203 10995 3209 11047
rect 4931 11016 4977 11274
tri 4977 11254 4997 11274 nw
tri 5740 11254 5760 11274 ne
rect 5760 11268 5796 11274
tri 5796 11268 5812 11284 sw
rect 5760 11254 5812 11268
tri 5760 11248 5766 11254 ne
rect 5006 11129 5012 11181
rect 5064 11129 5076 11181
rect 5128 11129 5136 11181
rect 5766 11178 5812 11254
tri 5812 11178 5846 11212 sw
tri 7009 11184 7025 11200 se
rect 7025 11184 7375 11200
tri 5984 11178 5990 11184 se
rect 5990 11178 5996 11184
rect 5315 11172 5680 11178
rect 5315 11138 5327 11172
rect 5361 11138 5404 11172
rect 5438 11138 5481 11172
rect 5515 11138 5558 11172
rect 5592 11138 5634 11172
rect 5668 11138 5680 11172
rect 5315 11132 5680 11138
rect 5766 11172 5996 11178
rect 6048 11172 6070 11184
rect 5766 11138 5803 11172
rect 5837 11138 5891 11172
rect 5925 11138 5979 11172
rect 6048 11138 6067 11172
rect 5766 11132 5996 11138
rect 6048 11132 6070 11138
rect 6122 11132 6143 11184
rect 6195 11132 6201 11184
tri 7003 11178 7009 11184 se
rect 7009 11178 7375 11184
tri 6979 11154 7003 11178 se
rect 7003 11154 7375 11178
tri 6959 11134 6979 11154 se
rect 6979 11134 7025 11154
tri 7025 11134 7045 11154 nw
tri 7289 11134 7309 11154 ne
rect 7309 11134 7375 11154
tri 6958 11133 6959 11134 se
rect 6959 11133 7024 11134
tri 7024 11133 7025 11134 nw
tri 7309 11133 7310 11134 ne
rect 7310 11133 7375 11134
rect 6958 11132 7023 11133
tri 7023 11132 7024 11133 nw
tri 7310 11132 7311 11133 ne
rect 7311 11132 7375 11133
tri 5375 11129 5378 11132 ne
rect 5378 11129 5455 11132
tri 5378 11098 5409 11129 ne
rect 5409 11078 5455 11129
tri 5455 11098 5489 11132 nw
rect 6958 11120 7011 11132
tri 7011 11120 7023 11132 nw
tri 7311 11120 7323 11132 ne
rect 6958 11116 7007 11120
tri 7007 11116 7011 11120 nw
tri 6944 11102 6958 11116 se
rect 6958 11102 7004 11116
tri 7004 11113 7007 11116 nw
rect 5714 11096 6281 11102
tri 6940 11098 6944 11102 se
rect 6944 11098 7004 11102
rect 5266 11050 5312 11062
tri 4977 11016 5009 11048 sw
tri 5234 11016 5266 11048 se
rect 5266 11016 5272 11050
rect 5306 11016 5312 11050
rect 4931 11014 5009 11016
tri 5009 11014 5011 11016 sw
tri 5232 11014 5234 11016 se
rect 5234 11014 5312 11016
rect 4931 11002 5039 11014
tri 3434 10995 3439 11000 se
tri 3093 10968 3120 10995 ne
rect 3120 10968 3127 10995
tri 3120 10961 3127 10968 ne
rect 3173 10968 3180 10995
tri 3180 10968 3207 10995 nw
tri 3407 10968 3434 10995 se
rect 3434 10968 3439 10995
tri 3173 10961 3180 10968 nw
tri 3406 10967 3407 10968 se
rect 3407 10967 3439 10968
tri 3485 10968 3517 11000 sw
tri 3719 10968 3751 11000 se
rect 3485 10967 3517 10968
tri 3517 10967 3518 10968 sw
tri 3718 10967 3719 10968 se
rect 3719 10967 3751 10968
tri 3797 10968 3829 11000 sw
tri 4031 10968 4063 11000 se
rect 3797 10967 3829 10968
tri 3829 10967 3830 10968 sw
tri 4030 10967 4031 10968 se
rect 4031 10967 4063 10968
tri 4109 10968 4141 11000 sw
tri 4343 10968 4375 11000 se
rect 4109 10967 4141 10968
tri 4141 10967 4142 10968 sw
tri 4342 10967 4343 10968 se
rect 4343 10967 4375 10968
tri 4421 10968 4453 11000 sw
rect 4931 10968 4999 11002
rect 5033 10968 5039 11002
rect 4421 10967 4453 10968
tri 4453 10967 4454 10968 sw
rect 3405 10915 3411 10967
rect 3463 10915 3480 10967
rect 3532 10915 3538 10967
rect 3701 10915 3707 10967
rect 3759 10915 3772 10967
rect 3824 10915 3830 10967
rect 4027 10915 4033 10967
rect 4085 10915 4097 10967
rect 4149 10915 4155 10967
rect 4336 10915 4342 10967
rect 4394 10915 4406 10967
rect 4458 10915 4464 10967
rect 4931 10930 5039 10968
tri 3405 10896 3424 10915 ne
rect 3424 10896 3439 10915
tri 3424 10882 3438 10896 ne
rect 3438 10882 3439 10896
rect 3485 10896 3499 10915
tri 3499 10896 3518 10915 nw
tri 3717 10896 3736 10915 ne
rect 3736 10896 3751 10915
rect 3485 10884 3487 10896
tri 3487 10884 3499 10896 nw
tri 3736 10884 3748 10896 ne
rect 3748 10884 3751 10896
tri 3485 10882 3487 10884 nw
tri 3748 10882 3750 10884 ne
rect 3750 10882 3751 10884
rect 3797 10896 3811 10915
tri 3811 10896 3830 10915 nw
tri 4029 10896 4048 10915 ne
rect 4048 10896 4063 10915
rect 3797 10884 3799 10896
tri 3799 10884 3811 10896 nw
tri 4048 10884 4060 10896 ne
rect 4060 10884 4063 10896
tri 3797 10882 3799 10884 nw
tri 4060 10882 4062 10884 ne
rect 4062 10882 4063 10884
tri 3438 10881 3439 10882 ne
tri 3750 10881 3751 10882 ne
tri 4062 10881 4063 10882 ne
rect 4109 10896 4124 10915
tri 4124 10896 4143 10915 nw
tri 4341 10896 4360 10915 ne
rect 4360 10896 4375 10915
rect 4109 10884 4112 10896
tri 4112 10884 4124 10896 nw
tri 4360 10884 4372 10896 ne
rect 4372 10884 4375 10896
tri 4109 10881 4112 10884 nw
tri 4372 10881 4375 10884 ne
rect 4421 10896 4436 10915
tri 4436 10896 4455 10915 nw
rect 4931 10896 4999 10930
rect 5033 10896 5039 10930
rect 4421 10884 4424 10896
tri 4424 10884 4436 10896 nw
rect 4931 10884 5039 10896
rect 5143 11002 5312 11014
rect 5143 10968 5149 11002
rect 5183 10970 5312 11002
rect 5183 10968 5272 10970
rect 5143 10936 5272 10968
rect 5306 10936 5312 10970
rect 5409 11044 5415 11078
rect 5449 11044 5455 11078
rect 5409 10993 5455 11044
rect 5409 10959 5415 10993
rect 5449 10959 5455 10993
tri 5312 10936 5334 10958 sw
tri 5387 10936 5409 10958 se
rect 5409 10936 5455 10959
rect 5565 11078 5611 11090
rect 5565 11044 5571 11078
rect 5605 11044 5611 11078
rect 5565 10970 5611 11044
rect 5714 11044 5721 11096
rect 5773 11044 5842 11096
rect 5894 11078 5963 11096
rect 5917 11044 5963 11078
rect 6015 11044 6083 11096
rect 6135 11078 6203 11096
rect 6135 11044 6195 11078
rect 6255 11044 6281 11096
tri 6924 11082 6940 11098 se
rect 6940 11082 7004 11098
rect 6824 11076 7004 11082
rect 5714 11042 6281 11044
rect 6683 11060 6757 11072
tri 5843 11026 5859 11042 ne
rect 5859 11026 5941 11042
tri 5941 11026 5957 11042 nw
tri 6155 11026 6171 11042 ne
rect 6171 11026 6253 11042
tri 6253 11026 6269 11042 nw
rect 6683 11026 6717 11060
rect 6751 11026 6757 11060
rect 6824 11042 6836 11076
rect 6870 11042 6908 11076
rect 6942 11042 7004 11076
rect 6824 11036 7004 11042
rect 7069 11057 7121 11069
tri 5859 11023 5862 11026 ne
rect 5862 11023 5938 11026
tri 5938 11023 5941 11026 nw
tri 6171 11023 6174 11026 ne
rect 6174 11023 6250 11026
tri 6250 11023 6253 11026 nw
tri 5862 11014 5871 11023 ne
rect 5871 11014 5923 11023
tri 5455 10936 5477 10958 sw
tri 5543 10936 5565 10958 se
rect 5565 10936 5571 10970
rect 5605 10953 5611 10970
rect 5721 11002 5767 11014
tri 5871 11008 5877 11014 ne
rect 5721 10968 5727 11002
rect 5761 10968 5767 11002
tri 5611 10953 5616 10958 sw
tri 5716 10953 5721 10958 se
rect 5721 10953 5767 10968
rect 5877 10998 5923 11014
tri 5923 11008 5938 11023 nw
tri 6174 11014 6183 11023 ne
rect 6183 11014 6235 11023
rect 5877 10964 5883 10998
rect 5917 10964 5923 10998
tri 5767 10953 5772 10958 sw
rect 5605 10951 5616 10953
tri 5616 10951 5618 10953 sw
tri 5714 10951 5716 10953 se
rect 5716 10951 5772 10953
tri 5772 10951 5774 10953 sw
rect 5877 10952 5923 10964
rect 6033 11002 6079 11014
tri 6183 11008 6189 11014 ne
rect 6033 10968 6039 11002
rect 6073 10968 6079 11002
tri 6028 10953 6033 10958 se
rect 6033 10953 6079 10968
rect 6189 10998 6235 11014
tri 6235 11008 6250 11023 nw
rect 6189 10964 6195 10998
rect 6229 10964 6235 10998
tri 6079 10953 6084 10958 sw
tri 6027 10952 6028 10953 se
rect 6028 10952 6084 10953
tri 6026 10951 6027 10952 se
rect 6027 10951 6084 10952
tri 6084 10951 6086 10953 sw
rect 6189 10952 6235 10964
rect 6345 11002 6391 11014
rect 6345 10968 6351 11002
rect 6385 10968 6391 11002
tri 6340 10953 6345 10958 se
rect 6345 10953 6391 10968
tri 6339 10952 6340 10953 se
rect 6340 10952 6391 10953
tri 6338 10951 6339 10952 se
rect 6339 10951 6391 10952
rect 5605 10936 5618 10951
rect 5143 10930 5334 10936
rect 5143 10896 5149 10930
rect 5183 10926 5334 10930
tri 5334 10926 5344 10936 sw
tri 5377 10926 5387 10936 se
rect 5387 10926 5477 10936
tri 5477 10926 5487 10936 sw
tri 5533 10926 5543 10936 se
rect 5543 10926 5618 10936
tri 5618 10926 5643 10951 sw
tri 5689 10926 5714 10951 se
rect 5714 10926 5774 10951
tri 5774 10926 5799 10951 sw
tri 6001 10926 6026 10951 se
rect 6026 10926 6086 10951
tri 6086 10926 6111 10951 sw
tri 6313 10926 6338 10951 se
rect 6338 10926 6391 10951
rect 5183 10924 5344 10926
tri 5344 10924 5346 10926 sw
tri 5375 10924 5377 10926 se
rect 5377 10924 5487 10926
tri 5487 10924 5489 10926 sw
tri 5531 10924 5533 10926 se
rect 5533 10924 5643 10926
tri 5643 10924 5645 10926 sw
tri 5687 10924 5689 10926 se
rect 5689 10924 5799 10926
tri 5799 10924 5801 10926 sw
tri 5999 10924 6001 10926 se
rect 6001 10924 6111 10926
tri 6111 10924 6113 10926 sw
tri 6311 10924 6313 10926 se
rect 6313 10924 6351 10926
rect 5183 10917 6351 10924
rect 5183 10908 5727 10917
rect 5183 10896 5415 10908
tri 4421 10881 4424 10884 nw
tri 3282 10875 3283 10876 se
tri 3329 10875 3330 10876 sw
tri 3594 10875 3595 10876 se
tri 3641 10875 3642 10876 sw
tri 3906 10875 3907 10876 se
tri 3953 10875 3954 10876 sw
tri 4218 10875 4219 10876 se
tri 4265 10875 4266 10876 sw
tri 4530 10875 4531 10876 se
tri 4577 10875 4578 10876 sw
tri 3281 10874 3282 10875 se
rect 3282 10874 3330 10875
tri 3330 10874 3331 10875 sw
tri 3593 10874 3594 10875 se
rect 3594 10874 3642 10875
tri 3642 10874 3643 10875 sw
tri 3905 10874 3906 10875 se
rect 3906 10874 3954 10875
tri 3954 10874 3955 10875 sw
tri 4217 10874 4218 10875 se
rect 4218 10874 4266 10875
tri 4266 10874 4267 10875 sw
tri 4529 10874 4530 10875 se
rect 4530 10874 4578 10875
tri 4578 10874 4579 10875 sw
tri 5142 10874 5143 10875 se
rect 5143 10874 5415 10896
rect 5449 10883 5727 10908
rect 5761 10916 6351 10917
rect 5761 10883 6039 10916
rect 5449 10882 6039 10883
rect 6073 10892 6351 10916
rect 6385 10892 6391 10926
rect 6073 10882 6391 10892
rect 5449 10874 6391 10882
tri 3257 10850 3281 10874 se
rect 3281 10850 3331 10874
tri 3331 10850 3355 10874 sw
tri 3569 10850 3593 10874 se
rect 3593 10850 3643 10874
tri 3643 10850 3667 10874 sw
tri 3881 10850 3905 10874 se
rect 3905 10850 3955 10874
tri 3955 10850 3979 10874 sw
tri 4193 10850 4217 10874 se
rect 4217 10850 4267 10874
tri 4267 10850 4291 10874 sw
tri 4505 10850 4529 10874 se
rect 4529 10850 4579 10874
tri 4579 10850 4603 10874 sw
tri 5118 10850 5142 10874 se
rect 5142 10850 6391 10874
tri 3249 10842 3257 10850 se
rect 3257 10842 3355 10850
tri 3355 10842 3363 10850 sw
tri 3561 10842 3569 10850 se
rect 3569 10842 3667 10850
tri 3667 10842 3675 10850 sw
tri 3873 10842 3881 10850 se
rect 3881 10842 3979 10850
tri 3979 10842 3987 10850 sw
tri 4185 10842 4193 10850 se
rect 4193 10842 4291 10850
tri 4291 10842 4299 10850 sw
tri 4497 10842 4505 10850 se
rect 4505 10842 4603 10850
tri 4603 10842 4611 10850 sw
tri 5110 10842 5118 10850 se
rect 5118 10842 6351 10850
rect 3115 10841 4618 10842
tri 4618 10841 4619 10842 sw
tri 5109 10841 5110 10842 se
rect 5110 10841 6351 10842
rect 3115 10789 3121 10841
rect 3173 10789 3186 10841
rect 3238 10789 3251 10841
rect 3303 10812 3316 10841
rect 3368 10812 3381 10841
rect 3433 10812 3446 10841
rect 3498 10812 3511 10841
rect 3563 10812 3576 10841
rect 3310 10789 3316 10812
rect 3563 10789 3572 10812
rect 3628 10789 3641 10841
rect 3693 10789 3706 10841
rect 3758 10789 3771 10841
rect 3823 10812 3836 10841
rect 3888 10812 3901 10841
rect 3953 10812 3966 10841
rect 4018 10812 4031 10841
rect 4083 10812 4096 10841
rect 3828 10789 3836 10812
rect 4083 10789 4090 10812
rect 4148 10789 4160 10841
rect 4212 10789 4224 10841
rect 4276 10789 4288 10841
rect 4340 10812 4352 10841
rect 4404 10812 4416 10841
rect 4468 10812 4480 10841
rect 4532 10812 4544 10841
rect 4346 10789 4352 10812
rect 4532 10789 4534 10812
rect 4596 10789 4608 10841
rect 4660 10789 4672 10841
rect 4724 10789 4736 10841
rect 4788 10789 4800 10841
rect 4852 10789 4864 10841
rect 4916 10789 4928 10841
rect 4980 10789 4992 10841
rect 5044 10789 5056 10841
rect 5108 10789 5120 10841
rect 5172 10789 5184 10841
rect 5236 10789 5248 10841
rect 5300 10789 5312 10841
rect 5364 10789 5376 10841
rect 5428 10789 5440 10841
rect 5492 10789 5504 10841
rect 5556 10789 5568 10841
rect 5620 10789 5632 10841
rect 5684 10789 5696 10841
rect 5748 10832 5760 10841
rect 5748 10789 5760 10798
rect 5812 10789 5824 10841
rect 5876 10789 5888 10841
rect 5940 10789 5952 10841
rect 6004 10789 6016 10841
rect 6068 10831 6080 10841
rect 6073 10797 6080 10831
rect 6068 10789 6080 10797
rect 6132 10789 6144 10841
rect 6196 10789 6208 10841
rect 6260 10816 6351 10841
rect 6385 10816 6391 10850
rect 6260 10804 6391 10816
rect 6683 10987 6757 11026
rect 6683 10953 6717 10987
rect 6751 10953 6757 10987
rect 7069 10993 7121 11005
rect 6683 10951 6757 10953
tri 6757 10951 6772 10966 sw
rect 6683 10932 6772 10951
tri 6772 10932 6791 10951 sw
rect 7069 10935 7121 10941
rect 6683 10926 6954 10932
rect 6683 10914 6836 10926
rect 6683 10880 6717 10914
rect 6751 10892 6836 10914
rect 6870 10892 6908 10926
rect 6942 10892 6954 10926
rect 6751 10880 6954 10892
rect 6683 10841 6954 10880
rect 6683 10835 6717 10841
rect 6751 10835 6954 10841
rect 6260 10789 6280 10804
rect 3115 10778 3127 10789
rect 3161 10778 3202 10789
rect 3236 10778 3276 10789
rect 3310 10778 3350 10789
rect 3384 10778 3424 10789
rect 3458 10778 3498 10789
rect 3532 10778 3572 10789
rect 3606 10778 3646 10789
rect 3680 10778 3720 10789
rect 3754 10778 3794 10789
rect 3828 10778 3868 10789
rect 3902 10778 3942 10789
rect 3976 10778 4016 10789
rect 4050 10778 4090 10789
rect 4124 10778 4164 10789
rect 4198 10778 4238 10789
rect 4272 10778 4312 10789
rect 4346 10778 4386 10789
rect 4420 10778 4460 10789
rect 4494 10778 4534 10789
rect 4568 10784 6280 10789
tri 6280 10784 6300 10804 nw
rect 4568 10778 6266 10784
rect 3115 10771 6266 10778
rect 3115 10719 3121 10771
rect 3173 10719 3186 10771
rect 3238 10719 3251 10771
rect 3303 10719 3316 10771
rect 3368 10719 3381 10771
rect 3433 10719 3446 10771
rect 3498 10719 3511 10771
rect 3563 10719 3576 10771
rect 3628 10719 3641 10771
rect 3693 10719 3706 10771
rect 3758 10719 3771 10771
rect 3823 10719 3836 10771
rect 3888 10719 3901 10771
rect 3953 10719 3966 10771
rect 4018 10719 4031 10771
rect 4083 10719 4096 10771
rect 4148 10719 4160 10771
rect 4212 10719 4224 10771
rect 4276 10719 4288 10771
rect 4340 10719 4352 10771
rect 4404 10719 4416 10771
rect 4468 10719 4480 10771
rect 4532 10719 4544 10771
rect 4596 10719 4608 10771
rect 4660 10719 4672 10771
rect 4724 10719 4736 10771
rect 4788 10719 4800 10771
rect 4852 10719 4864 10771
rect 4916 10719 4928 10771
rect 4980 10719 4992 10771
rect 5044 10719 5056 10771
rect 5108 10719 5120 10771
rect 5172 10719 5184 10771
rect 5236 10719 5248 10771
rect 5300 10719 5312 10771
rect 5364 10719 5376 10771
rect 5428 10719 5440 10771
rect 5492 10719 5504 10771
rect 5556 10719 5568 10771
rect 5620 10719 5632 10771
rect 5684 10719 5696 10771
rect 5748 10719 5760 10771
rect 5812 10719 5824 10771
rect 5876 10719 5888 10771
rect 5940 10719 5952 10771
rect 6004 10719 6016 10771
rect 6068 10719 6080 10771
rect 6132 10719 6144 10771
rect 6196 10719 6208 10771
rect 6260 10719 6266 10771
tri 6266 10770 6280 10784 nw
rect 6683 10783 6711 10835
rect 6763 10783 6811 10835
rect 6863 10824 6954 10835
tri 6954 10824 6988 10858 sw
rect 6863 10818 7268 10824
rect 6863 10784 6923 10818
rect 6957 10784 7022 10818
rect 7056 10784 7122 10818
rect 7156 10784 7268 10818
rect 6863 10783 7268 10784
rect 6683 10778 7268 10783
rect 6683 10771 6864 10778
rect 3115 10714 6266 10719
rect 3115 10701 4989 10714
rect 5023 10701 5062 10714
rect 5096 10701 5135 10714
rect 5169 10701 5208 10714
rect 5242 10701 5281 10714
rect 5315 10701 5354 10714
rect 5388 10701 5427 10714
rect 5461 10701 5500 10714
rect 5534 10701 5572 10714
rect 5606 10701 5644 10714
rect 5678 10701 5716 10714
rect 5750 10701 5788 10714
rect 5822 10701 5860 10714
rect 5894 10701 5932 10714
rect 5966 10701 6004 10714
rect 6038 10701 6076 10714
rect 6110 10701 6148 10714
rect 6182 10701 6220 10714
rect 6254 10701 6266 10714
rect 3115 10649 3121 10701
rect 3173 10649 3186 10701
rect 3238 10649 3251 10701
rect 3303 10649 3316 10701
rect 3368 10649 3381 10701
rect 3433 10649 3446 10701
rect 3498 10649 3511 10701
rect 3563 10649 3576 10701
rect 3628 10649 3641 10701
rect 3693 10649 3706 10701
rect 3758 10649 3771 10701
rect 3823 10649 3836 10701
rect 3888 10649 3901 10701
rect 3953 10649 3966 10701
rect 4018 10649 4031 10701
rect 4083 10649 4096 10701
rect 4148 10649 4160 10701
rect 4212 10649 4224 10701
rect 4276 10649 4288 10701
rect 4340 10649 4352 10701
rect 4404 10649 4416 10701
rect 4468 10649 4480 10701
rect 4532 10649 4544 10701
rect 4596 10649 4608 10701
rect 4660 10649 4672 10701
rect 4724 10649 4736 10701
rect 4788 10649 4800 10701
rect 4852 10649 4864 10701
rect 4916 10649 4928 10701
rect 4980 10680 4989 10701
rect 4980 10649 4992 10680
rect 5044 10649 5056 10701
rect 5108 10649 5120 10701
rect 5172 10649 5184 10701
rect 5242 10680 5248 10701
rect 5492 10680 5500 10701
rect 5236 10649 5248 10680
rect 5300 10649 5312 10680
rect 5364 10649 5376 10680
rect 5428 10649 5440 10680
rect 5492 10649 5504 10680
rect 5556 10649 5568 10701
rect 5620 10649 5632 10701
rect 5684 10649 5696 10701
rect 5750 10680 5760 10701
rect 5822 10680 5824 10701
rect 6068 10680 6076 10701
rect 5748 10649 5760 10680
rect 5812 10649 5824 10680
rect 5876 10649 5888 10680
rect 5940 10649 5952 10680
rect 6004 10649 6016 10680
rect 6068 10649 6080 10680
rect 6132 10649 6144 10701
rect 6196 10649 6208 10701
rect 6260 10649 6266 10701
rect 6683 10719 6711 10771
rect 6763 10719 6811 10771
rect 6863 10719 6864 10771
tri 6864 10744 6898 10778 nw
tri 7188 10744 7222 10778 ne
rect 6683 10707 6864 10719
rect 6683 10655 6711 10707
rect 6763 10655 6811 10707
rect 6863 10692 6864 10707
rect 7222 10726 7268 10778
tri 6864 10692 6872 10700 sw
rect 7222 10692 7228 10726
rect 7262 10692 7268 10726
rect 6863 10666 6872 10692
tri 6872 10666 6898 10692 sw
rect 6863 10660 7086 10666
rect 6683 10626 6836 10655
rect 6870 10626 6938 10660
rect 6972 10626 7040 10660
rect 7074 10626 7086 10660
rect 6683 10622 7086 10626
rect 6683 10588 6717 10622
rect 6751 10620 7086 10622
rect 7222 10651 7268 10692
rect 6751 10617 6895 10620
tri 6895 10617 6898 10620 nw
rect 7222 10617 7228 10651
rect 7262 10617 7268 10651
rect 6751 10588 6864 10617
rect 6683 10549 6864 10588
tri 6864 10586 6895 10617 nw
rect 7222 10576 7268 10617
rect 6314 10521 6519 10527
rect 6366 10469 6390 10521
rect 6442 10469 6466 10521
rect 6518 10469 6519 10521
rect 6314 10449 6519 10469
rect 6366 10397 6390 10449
rect 6442 10397 6466 10449
rect 6518 10397 6519 10449
rect 6314 10377 6519 10397
rect 6366 10325 6390 10377
rect 6442 10325 6466 10377
rect 6518 10325 6519 10377
rect 6314 10305 6519 10325
rect 3729 10251 3735 10303
rect 3787 10251 3799 10303
rect 3851 10251 4313 10303
tri 4227 10227 4251 10251 ne
rect 4251 10227 4313 10251
tri 4251 10217 4261 10227 ne
rect 4261 10203 4313 10227
rect 6366 10253 6390 10305
rect 6442 10253 6466 10305
rect 6518 10253 6519 10305
rect 6314 10233 6519 10253
tri 4313 10203 4315 10205 sw
rect 4261 10192 4315 10203
tri 4315 10192 4326 10203 sw
rect 4261 10189 4326 10192
tri 4326 10189 4329 10192 sw
rect 3255 10125 3261 10177
rect 3313 10125 3327 10177
rect 3379 10125 3385 10177
rect 3743 10122 4088 10174
rect 4261 10171 4329 10189
tri 4329 10171 4347 10189 sw
rect 6366 10181 6390 10233
rect 6442 10181 6466 10233
rect 6518 10181 6519 10233
rect 4261 10125 4313 10171
rect 6314 10161 6519 10181
rect 3743 10117 3824 10122
tri 3824 10117 3829 10122 nw
rect 3505 10007 3633 10051
tri 3735 10011 3743 10019 se
rect 3743 10011 3795 10117
tri 3795 10088 3824 10117 nw
rect 6366 10109 6390 10161
rect 6442 10109 6466 10161
rect 6518 10109 6519 10161
tri 3795 10011 3803 10019 sw
rect 3505 9955 3511 10007
rect 3563 9955 3575 10007
rect 3627 9955 3633 10007
tri 3726 10002 3735 10011 se
rect 3735 10002 3803 10011
tri 3803 10002 3812 10011 sw
tri 3725 10001 3726 10002 se
rect 3726 10001 3812 10002
tri 3709 9985 3725 10001 se
rect 3725 9985 3812 10001
tri 3812 9985 3829 10002 sw
rect 3505 9921 3633 9955
rect 3702 9933 3708 9985
rect 3760 9933 3772 9985
rect 3824 9933 3830 9985
tri 3113 9867 3143 9897 se
tri 6284 9867 6314 9897 se
rect 6314 9867 6519 10109
tri 3109 9863 3113 9867 se
rect 3113 9863 3143 9867
tri 6280 9863 6284 9867 se
rect 6284 9863 6519 9867
rect 3093 9851 3690 9863
rect 3093 9799 3099 9851
rect 3151 9799 3166 9851
rect 3218 9799 3233 9851
rect 3285 9799 3300 9851
rect 3352 9799 3367 9851
rect 3419 9799 3434 9851
rect 3486 9799 3500 9851
rect 3552 9799 3566 9851
rect 3618 9799 3632 9851
rect 3684 9812 3690 9851
rect 6314 9814 6519 9863
rect 6683 10515 6717 10549
rect 6751 10542 6864 10549
rect 7120 10545 7180 10551
tri 6864 10542 6866 10544 sw
rect 6751 10521 6866 10542
rect 6683 10477 6744 10515
rect 6683 10443 6717 10477
rect 6796 10469 6812 10521
rect 6864 10510 6866 10521
tri 6866 10510 6898 10542 sw
rect 6864 10504 7086 10510
rect 6864 10470 6922 10504
rect 6956 10470 7040 10504
rect 7074 10470 7086 10504
rect 6864 10469 7086 10470
rect 6751 10464 7086 10469
rect 7120 10493 7128 10545
rect 7120 10481 7180 10493
rect 6751 10449 6869 10464
rect 6683 10405 6744 10443
rect 6683 10371 6717 10405
rect 6796 10397 6812 10449
rect 6864 10435 6869 10449
tri 6869 10435 6898 10464 nw
tri 6864 10430 6869 10435 nw
rect 6751 10377 6864 10397
rect 7120 10429 7128 10481
rect 6683 10333 6744 10371
rect 6683 10299 6717 10333
rect 6796 10325 6812 10377
tri 6864 10354 6898 10388 sw
rect 6864 10348 7086 10354
rect 6751 10314 6836 10325
rect 6870 10314 6938 10348
rect 6972 10314 7040 10348
rect 7074 10314 7086 10348
rect 6751 10308 7086 10314
rect 6751 10305 6871 10308
rect 6683 10261 6744 10299
rect 6683 10227 6717 10261
rect 6796 10253 6812 10305
rect 6864 10281 6871 10305
tri 6871 10281 6898 10308 nw
tri 6864 10274 6871 10281 nw
rect 6751 10233 6864 10253
rect 6683 10189 6744 10227
rect 6683 10155 6717 10189
rect 6796 10181 6812 10233
tri 7091 10203 7120 10232 se
rect 7120 10203 7180 10429
rect 7222 10542 7228 10576
rect 7262 10542 7268 10576
rect 7222 10501 7268 10542
rect 7222 10467 7228 10501
rect 7262 10467 7268 10501
rect 7222 10426 7268 10467
rect 7222 10392 7228 10426
rect 7262 10392 7268 10426
rect 7222 10380 7268 10392
rect 7323 10315 7375 11132
tri 7086 10198 7091 10203 se
rect 7091 10198 7180 10203
rect 6751 10161 6864 10181
rect 6683 10117 6744 10155
rect 6683 10083 6717 10117
rect 6796 10109 6812 10161
rect 6909 10192 7180 10198
rect 6909 10158 6921 10192
rect 6955 10158 7021 10192
rect 7055 10158 7122 10192
rect 7156 10158 7180 10192
rect 6909 10152 7180 10158
tri 7086 10125 7113 10152 ne
rect 7113 10125 7180 10152
tri 7113 10118 7120 10125 ne
rect 6751 10083 6864 10109
rect 6683 10048 6864 10083
tri 6864 10048 6892 10076 sw
rect 6683 10045 6892 10048
rect 6683 10011 6717 10045
rect 6751 10042 6892 10045
tri 6892 10042 6898 10048 sw
rect 6751 10036 7086 10042
rect 6751 10011 6836 10036
rect 6683 10002 6836 10011
rect 6870 10002 6938 10036
rect 6972 10002 7040 10036
rect 7074 10002 7086 10036
rect 6683 9996 7086 10002
rect 6683 9973 6873 9996
rect 6683 9939 6717 9973
rect 6751 9971 6873 9973
tri 6873 9971 6898 9996 nw
rect 6751 9939 6864 9971
tri 6864 9962 6873 9971 nw
rect 6683 9901 6864 9939
rect 6683 9867 6717 9901
rect 6751 9867 6864 9901
tri 7094 9894 7120 9920 se
rect 7120 9894 7180 10125
tri 7086 9886 7094 9894 se
rect 7094 9886 7180 9894
rect 6683 9829 6864 9867
rect 6912 9880 7180 9886
rect 6912 9846 6924 9880
rect 6958 9846 7023 9880
rect 7057 9846 7122 9880
rect 7156 9846 7180 9880
rect 7222 10281 7268 10293
rect 7222 10247 7228 10281
rect 7262 10247 7268 10281
rect 7323 10251 7375 10263
rect 7222 10245 7268 10247
tri 7268 10245 7274 10251 sw
rect 7222 10239 7274 10245
rect 7323 10193 7375 10199
rect 8465 10994 8517 11000
rect 8465 10930 8517 10942
rect 7222 10175 7228 10187
rect 7262 10175 7274 10187
rect 7222 10091 7228 10123
rect 7262 10117 7274 10123
rect 7262 10091 7268 10117
tri 7268 10111 7274 10117 nw
rect 7715 10159 7843 10165
rect 7222 10048 7268 10091
rect 7222 10014 7228 10048
rect 7262 10014 7268 10048
rect 7222 9971 7268 10014
rect 7222 9937 7228 9971
rect 7262 9937 7268 9971
rect 7222 9894 7268 9937
rect 7222 9860 7228 9894
rect 7262 9860 7268 9894
rect 7222 9848 7268 9860
rect 7767 10107 7791 10159
rect 7715 10069 7843 10107
rect 7767 10017 7791 10069
rect 6912 9840 7180 9846
rect 3684 9799 6451 9812
rect 3093 9778 6451 9799
rect 3093 9771 3690 9778
rect 3093 9719 3099 9771
rect 3151 9719 3166 9771
rect 3218 9719 3233 9771
rect 3285 9719 3300 9771
rect 3352 9719 3367 9771
rect 3419 9719 3434 9771
rect 3486 9719 3500 9771
rect 3552 9719 3566 9771
rect 3618 9719 3632 9771
rect 3684 9731 3690 9771
rect 3684 9724 3695 9731
tri 3695 9724 3702 9731 nw
rect 3684 9719 3690 9724
tri 3690 9719 3695 9724 nw
rect 5831 9609 5837 9661
rect 5889 9609 5901 9661
rect 5953 9609 5959 9661
rect 6028 9643 6156 9673
tri 5832 9595 5846 9609 ne
rect 5846 9595 5938 9609
tri 5938 9595 5952 9609 nw
tri 5846 9575 5866 9595 ne
tri 5853 9493 5866 9506 se
rect 5866 9493 5918 9595
tri 5918 9575 5938 9595 nw
rect 6028 9591 6034 9643
rect 6086 9591 6098 9643
rect 6150 9591 6156 9643
rect 6028 9543 6156 9591
tri 5843 9483 5853 9493 se
rect 5853 9483 5918 9493
tri 5832 9472 5843 9483 se
rect 5843 9472 5918 9483
rect 5348 9423 5400 9469
tri 5314 9415 5322 9423 ne
rect 5322 9415 5400 9423
rect 5573 9420 5918 9472
rect 6276 9417 6282 9469
rect 6334 9417 6348 9469
rect 6400 9417 6406 9469
tri 5322 9412 5325 9415 ne
rect 5325 9412 5400 9415
tri 5325 9410 5327 9412 ne
rect 5327 9410 5400 9412
tri 5327 9389 5348 9410 ne
rect 5348 9376 5400 9410
tri 5400 9376 5401 9377 sw
rect 5348 9343 5401 9376
tri 5401 9343 5434 9376 sw
rect 5348 9291 5810 9343
rect 5862 9291 5874 9343
rect 5926 9291 5932 9343
rect 6491 9195 6519 9805
rect 6683 9795 6717 9829
rect 6751 9795 6864 9829
rect 6683 9733 6864 9795
tri 6864 9733 6895 9764 sw
rect 6683 9730 6895 9733
tri 6895 9730 6898 9733 sw
rect 6571 9720 6623 9726
rect 6571 9656 6623 9668
rect 5348 8541 5810 8593
rect 5862 8541 5874 8593
rect 5926 8541 5932 8593
rect 5348 8509 5402 8541
tri 5402 8509 5434 8541 nw
tri 5341 8488 5348 8495 se
rect 5348 8488 5400 8509
tri 5400 8507 5402 8509 nw
tri 5324 8471 5341 8488 se
rect 5341 8471 5400 8488
tri 5314 8461 5324 8471 se
rect 5324 8461 5400 8471
rect 5348 8415 5400 8461
rect 5573 8412 5918 8464
rect 6276 8415 6282 8467
rect 6334 8415 6348 8467
rect 6400 8415 6406 8467
tri 5832 8400 5844 8412 ne
rect 5844 8400 5918 8412
tri 5844 8378 5866 8400 ne
tri 5850 8293 5866 8309 se
rect 5866 8293 5918 8400
tri 5918 8293 5934 8309 sw
rect 6028 8293 6156 8341
tri 5832 8275 5850 8293 se
rect 5850 8275 5934 8293
tri 5934 8275 5952 8293 sw
rect 5831 8223 5837 8275
rect 5889 8223 5901 8275
rect 5953 8223 5959 8275
rect 6028 8241 6034 8293
rect 6086 8241 6098 8293
rect 6150 8241 6156 8293
rect 6028 8211 6156 8241
rect 6571 8254 6623 9604
rect 6683 9724 7086 9730
rect 6683 9702 6836 9724
rect 6683 9668 6717 9702
rect 6751 9690 6836 9702
rect 6870 9690 6938 9724
rect 6972 9690 7040 9724
rect 7074 9690 7086 9724
rect 6751 9684 7086 9690
rect 6751 9668 6873 9684
rect 6683 9659 6873 9668
tri 6873 9659 6898 9684 nw
rect 6683 9629 6864 9659
tri 6864 9650 6873 9659 nw
rect 6683 9595 6717 9629
rect 6751 9595 6864 9629
rect 6683 9556 6864 9595
rect 7222 9608 7228 9660
rect 7280 9608 7292 9660
rect 7344 9608 7350 9660
rect 6683 9522 6717 9556
rect 6751 9522 6864 9556
rect 6912 9568 7170 9574
rect 6912 9534 6924 9568
rect 6958 9534 7023 9568
rect 7057 9534 7122 9568
rect 7156 9534 7170 9568
rect 6912 9528 7170 9534
rect 6683 9483 6864 9522
tri 7084 9494 7118 9528 ne
rect 6683 9449 6717 9483
rect 6751 9449 6864 9483
rect 6683 9418 6864 9449
tri 6864 9418 6898 9452 sw
rect 6683 9412 7086 9418
rect 6683 9410 6836 9412
rect 6683 9376 6717 9410
rect 6751 9378 6836 9410
rect 6870 9378 6938 9412
rect 6972 9378 7040 9412
rect 7074 9378 7086 9412
rect 6751 9376 7086 9378
rect 6683 9372 7086 9376
rect 6683 9337 6864 9372
tri 6864 9338 6898 9372 nw
rect 6683 9303 6717 9337
rect 6751 9303 6864 9337
rect 6683 9264 6864 9303
rect 6683 9230 6717 9264
rect 6751 9230 6864 9264
tri 7084 9262 7118 9296 se
rect 7118 9262 7170 9528
rect 6683 9191 6864 9230
rect 6912 9256 7040 9262
rect 6912 9222 6924 9256
rect 6958 9222 7023 9256
rect 6912 9210 7040 9222
rect 7092 9210 7112 9262
rect 7164 9210 7170 9262
rect 7222 9571 7268 9608
tri 7268 9574 7302 9608 nw
rect 7222 9537 7228 9571
rect 7262 9537 7268 9571
rect 7222 9493 7268 9537
rect 7222 9459 7228 9493
rect 7262 9459 7268 9493
rect 7222 9415 7268 9459
rect 7222 9381 7228 9415
rect 7262 9381 7268 9415
rect 7222 9337 7268 9381
rect 7222 9303 7228 9337
rect 7262 9303 7268 9337
rect 7222 9259 7268 9303
rect 7222 9225 7228 9259
rect 7262 9225 7268 9259
rect 6683 9157 6717 9191
rect 6751 9157 6864 9191
rect 6683 9119 6864 9157
rect 7222 9181 7268 9225
rect 7715 9262 7843 10017
rect 8465 9955 8517 10878
rect 8570 10633 8698 12901
rect 8570 10581 8576 10633
rect 8628 10581 8640 10633
rect 8692 10581 8698 10633
rect 8758 10635 8824 13262
tri 8824 10635 8858 10669 sw
rect 8758 10583 8764 10635
rect 8816 10583 8846 10635
rect 8898 10583 8904 10635
rect 9005 10391 9145 13804
tri 9145 13770 9179 13804 nw
rect 9385 13577 9544 14489
rect 9385 13525 9391 13577
rect 9443 13525 9486 13577
rect 9538 13525 9544 13577
rect 9385 13501 9544 13525
rect 9385 13449 9391 13501
rect 9443 13449 9486 13501
rect 9538 13449 9544 13501
rect 9385 13044 9544 13449
rect 9385 12992 9391 13044
rect 9443 12992 9486 13044
rect 9538 12992 9544 13044
rect 9385 12948 9544 12992
rect 9385 12896 9391 12948
rect 9443 12896 9486 12948
rect 9538 12896 9544 12948
rect 9385 12895 9544 12896
rect 9336 12349 9342 12401
rect 9394 12349 9406 12401
rect 9458 12349 9464 12401
tri 9378 12321 9406 12349 ne
rect 9406 12321 9464 12349
rect 9226 12269 9232 12321
rect 9284 12269 9296 12321
rect 9348 12269 9354 12321
tri 9406 12315 9412 12321 ne
rect 9226 12244 9287 12269
tri 9287 12244 9312 12269 nw
rect 9226 12100 9278 12244
tri 9278 12235 9287 12244 nw
tri 9278 12100 9289 12111 sw
rect 9226 12087 9289 12100
tri 9289 12087 9302 12100 sw
rect 9226 12077 9302 12087
tri 9302 12077 9312 12087 sw
rect 9226 12025 9384 12077
tri 9298 11991 9332 12025 ne
rect 9176 11869 9182 11921
rect 9234 11869 9246 11921
rect 9298 11869 9304 11921
tri 9218 11866 9221 11869 ne
rect 9221 11866 9304 11869
tri 9221 11835 9252 11866 ne
rect 9005 10339 9011 10391
rect 9063 10339 9087 10391
rect 9139 10339 9145 10391
rect 9005 10325 9145 10339
rect 9005 10273 9011 10325
rect 9063 10273 9087 10325
rect 9139 10273 9145 10325
rect 8856 10193 8862 10245
rect 8914 10193 8926 10245
rect 8978 10193 8984 10245
tri 8898 10159 8932 10193 ne
tri 8517 9955 8528 9966 sw
rect 8465 9944 8528 9955
tri 8465 9881 8528 9944 ne
tri 8528 9881 8602 9955 sw
tri 8528 9807 8602 9881 ne
tri 8602 9807 8676 9881 sw
tri 8602 9733 8676 9807 ne
tri 8676 9733 8750 9807 sw
tri 8676 9659 8750 9733 ne
tri 8750 9659 8824 9733 sw
tri 8750 9637 8772 9659 ne
rect 8292 9417 8298 9469
rect 8350 9417 8362 9469
rect 8414 9417 8420 9469
tri 8334 9383 8368 9417 ne
rect 7715 9210 7721 9262
rect 7773 9210 7785 9262
rect 7837 9210 7843 9262
rect 7222 9147 7228 9181
rect 7262 9151 7268 9181
tri 7268 9151 7302 9185 sw
rect 7262 9147 7331 9151
rect 6683 9085 6717 9119
rect 6751 9106 6864 9119
tri 6864 9106 6898 9140 sw
rect 7222 9121 7331 9147
tri 7331 9121 7361 9151 sw
rect 6751 9100 7086 9106
rect 7222 9105 7361 9121
rect 6751 9085 6836 9100
rect 6683 9066 6836 9085
rect 6870 9066 6938 9100
rect 6972 9066 7040 9100
rect 7074 9066 7086 9100
tri 7281 9071 7315 9105 ne
rect 6683 9060 7086 9066
rect 6683 9047 6871 9060
rect 6683 9013 6717 9047
rect 6751 9033 6871 9047
tri 6871 9033 6898 9060 nw
rect 7222 9033 7268 9045
rect 6751 9013 6864 9033
tri 6864 9026 6871 9033 nw
rect 6683 8975 6864 9013
rect 7222 8999 7228 9033
rect 7262 8999 7268 9033
rect 6683 8941 6717 8975
rect 6751 8950 6864 8975
tri 6864 8950 6898 8984 sw
tri 7188 8950 7222 8984 se
rect 7222 8950 7268 8999
rect 6751 8946 7268 8950
rect 6751 8944 7228 8946
rect 6751 8941 6924 8944
rect 6683 8910 6924 8941
rect 6958 8910 7023 8944
rect 7057 8910 7122 8944
rect 7156 8912 7228 8944
rect 7262 8912 7268 8946
rect 7156 8910 7268 8912
rect 6683 8904 7268 8910
rect 6683 8903 6864 8904
rect 6683 8869 6717 8903
rect 6751 8869 6864 8903
tri 6864 8870 6898 8904 nw
tri 7188 8870 7222 8904 ne
rect 6683 8831 6864 8869
rect 6683 8797 6717 8831
rect 6751 8825 6864 8831
rect 7222 8859 7268 8904
tri 6864 8825 6867 8828 sw
rect 7222 8825 7228 8859
rect 7262 8825 7268 8859
rect 6751 8797 6867 8825
rect 6683 8794 6867 8797
tri 6867 8794 6898 8825 sw
rect 6683 8788 7086 8794
rect 6683 8759 6836 8788
rect 6683 8725 6717 8759
rect 6751 8754 6836 8759
rect 6870 8754 6938 8788
rect 6972 8754 7040 8788
rect 7074 8754 7086 8788
rect 6751 8748 7086 8754
rect 7222 8772 7268 8825
rect 6751 8738 6888 8748
tri 6888 8738 6898 8748 nw
rect 7222 8738 7228 8772
rect 7262 8738 7268 8772
rect 6751 8725 6864 8738
rect 6683 8687 6864 8725
tri 6864 8714 6888 8738 nw
tri 7206 8714 7222 8730 se
rect 7222 8714 7268 8738
tri 7188 8696 7206 8714 se
rect 7206 8696 7268 8714
rect 6683 8653 6717 8687
rect 6751 8653 6864 8687
rect 6683 8615 6864 8653
rect 6683 8581 6717 8615
rect 6751 8581 6864 8615
rect 6912 8685 7268 8696
rect 6912 8651 7228 8685
rect 7262 8651 7268 8685
rect 6912 8632 7268 8651
rect 6912 8598 6924 8632
rect 6958 8598 7023 8632
rect 7057 8598 7122 8632
rect 7156 8598 7268 8632
rect 6912 8592 7268 8598
rect 6683 8543 6864 8581
rect 6683 8509 6717 8543
rect 6751 8509 6864 8543
tri 7281 8528 7315 8562 se
rect 7315 8528 7361 9105
rect 8208 8927 8260 8933
rect 8208 8863 8260 8875
rect 6683 8471 6864 8509
rect 6899 8522 7361 8528
rect 6899 8488 6911 8522
rect 6945 8488 6983 8522
rect 7017 8488 7361 8522
rect 6899 8482 7361 8488
rect 7903 8771 7955 8777
rect 7903 8707 7955 8719
rect 6683 8437 6717 8471
rect 6751 8437 6864 8471
rect 6683 8425 6864 8437
tri 6683 8400 6708 8425 ne
rect 6708 8400 6864 8425
rect 7072 8434 7118 8446
tri 6864 8400 6870 8406 sw
rect 7072 8400 7078 8434
rect 7112 8400 7118 8434
tri 6708 8366 6742 8400 ne
rect 6742 8372 6870 8400
tri 6870 8372 6898 8400 sw
rect 6742 8366 6954 8372
tri 6742 8364 6744 8366 ne
rect 6744 8332 6836 8366
rect 6870 8332 6908 8366
rect 6942 8332 6954 8366
rect 6744 8326 6954 8332
rect 7072 8327 7118 8400
tri 6623 8254 6657 8288 sw
rect 6571 8202 6902 8254
rect 7072 8242 7078 8327
rect 7112 8294 7118 8327
tri 7118 8294 7152 8328 sw
tri 7869 8294 7903 8328 se
rect 7903 8294 7955 8655
rect 7130 8242 7143 8294
rect 7195 8242 7201 8294
rect 7827 8242 7833 8294
rect 7885 8242 7897 8294
rect 7949 8242 7955 8294
tri 7869 8208 7903 8242 ne
tri 6816 8168 6850 8202 ne
rect 3142 8152 6518 8153
rect 3142 8100 3148 8152
rect 3200 8100 3213 8152
rect 3265 8100 3278 8152
rect 3330 8100 3343 8152
rect 3395 8100 3408 8152
rect 3460 8100 3473 8152
rect 3525 8100 3538 8152
rect 3590 8100 3603 8152
rect 3655 8100 3668 8152
rect 3720 8100 3733 8152
rect 3785 8100 3798 8152
rect 3850 8100 3863 8152
rect 3915 8100 3928 8152
rect 3980 8100 3993 8152
rect 4045 8100 4058 8152
rect 4110 8100 4123 8152
rect 4175 8100 4188 8152
rect 4240 8100 4253 8152
rect 4305 8100 4318 8152
rect 4370 8100 4383 8152
rect 3142 8088 4383 8100
rect 3142 8036 3148 8088
rect 3200 8036 3213 8088
rect 3265 8036 3278 8088
rect 3330 8036 3343 8088
rect 3395 8036 3408 8088
rect 3460 8036 3473 8088
rect 3525 8036 3538 8088
rect 3590 8036 3603 8088
rect 3655 8036 3668 8088
rect 3720 8036 3733 8088
rect 3785 8036 3798 8088
rect 3850 8036 3863 8088
rect 3915 8036 3928 8088
rect 3980 8036 3993 8088
rect 4045 8036 4058 8088
rect 4110 8036 4123 8088
rect 4175 8036 4188 8088
rect 4240 8036 4253 8088
rect 4305 8036 4318 8088
rect 4370 8036 4383 8088
rect 3142 8024 4383 8036
rect 3142 7972 3148 8024
rect 3200 7972 3213 8024
rect 3265 7972 3278 8024
rect 3330 7972 3343 8024
rect 3395 7972 3408 8024
rect 3460 7972 3473 8024
rect 3525 7972 3538 8024
rect 3590 7972 3603 8024
rect 3655 7972 3668 8024
rect 3720 7972 3733 8024
rect 3785 7972 3798 8024
rect 3850 7972 3863 8024
rect 3915 7972 3928 8024
rect 3980 7972 3993 8024
rect 4045 7972 4058 8024
rect 4110 7972 4123 8024
rect 4175 7972 4188 8024
rect 4240 7972 4253 8024
rect 4305 7972 4318 8024
rect 4370 7972 4383 8024
rect 5459 7972 6518 8152
rect 3142 7970 6518 7972
tri 2842 7926 2876 7960 sw
tri 6710 7926 6744 7960 se
rect 2842 7920 6744 7926
rect 2842 7886 2874 7920
rect 2908 7886 2948 7920
rect 2982 7886 3022 7920
rect 3056 7886 3096 7920
rect 3130 7886 3170 7920
rect 3204 7886 3244 7920
rect 3278 7886 3318 7920
rect 3352 7886 3392 7920
rect 3426 7886 3466 7920
rect 3500 7886 3539 7920
rect 3573 7886 3612 7920
rect 3646 7886 3685 7920
rect 3719 7886 3758 7920
rect 3792 7886 3831 7920
rect 3865 7886 3904 7920
rect 3938 7886 3977 7920
rect 4011 7886 4050 7920
rect 4084 7886 4123 7920
rect 4157 7886 4196 7920
rect 4230 7886 4269 7920
rect 4303 7886 4342 7920
rect 4376 7886 4415 7920
rect 4449 7886 4488 7920
rect 4522 7886 4561 7920
rect 4595 7886 4634 7920
rect 4668 7886 4707 7920
rect 4741 7886 4780 7920
rect 4814 7886 4853 7920
rect 4887 7886 4926 7920
rect 4960 7886 4999 7920
rect 5033 7886 5072 7920
rect 5106 7886 5145 7920
rect 5179 7886 5218 7920
rect 5252 7886 5291 7920
rect 5325 7886 5364 7920
rect 5398 7886 5437 7920
rect 5471 7886 5510 7920
rect 5544 7886 5583 7920
rect 5617 7886 5656 7920
rect 5690 7886 5729 7920
rect 5763 7886 5802 7920
rect 5836 7886 5875 7920
rect 5909 7886 5948 7920
rect 5982 7886 6021 7920
rect 6055 7886 6094 7920
rect 6128 7886 6167 7920
rect 6201 7886 6240 7920
rect 6274 7886 6313 7920
rect 6347 7886 6386 7920
rect 6420 7886 6459 7920
rect 6493 7886 6532 7920
rect 6566 7886 6605 7920
rect 6639 7886 6678 7920
rect 6712 7886 6744 7920
rect 2842 7880 6744 7886
rect 2842 7852 2848 7880
tri 2848 7852 2876 7880 nw
tri 6710 7852 6738 7880 ne
rect 6738 7852 6744 7880
rect 2842 7847 2843 7852
tri 2843 7847 2848 7852 nw
tri 6738 7847 6743 7852 ne
rect 6743 7847 6744 7852
tri 2842 7846 2843 7847 nw
tri 6743 7846 6744 7847 ne
tri 5648 7285 5649 7286 ne
rect 5649 7285 5653 7286
tri 5649 7281 5653 7285 ne
rect 5699 7285 5732 7286
tri 5732 7285 5733 7286 nw
rect 5699 7281 5728 7285
tri 5728 7281 5732 7285 nw
rect 5699 7262 5709 7281
tri 5709 7262 5728 7281 nw
tri 5699 7252 5709 7262 nw
tri 5855 6595 5861 6601 sw
tri 5855 6461 5861 6467 nw
tri 5595 5759 5618 5782 sw
rect 5595 5748 5618 5759
tri 5618 5748 5629 5759 sw
tri 5806 5490 5809 5493 se
tri 5787 5471 5806 5490 se
rect 5806 5471 5809 5490
tri 5775 5459 5787 5471 se
rect 5787 5459 5809 5471
tri 5855 5490 5858 5493 sw
rect 5855 5471 5858 5490
tri 5858 5471 5877 5490 sw
rect 5855 5459 5877 5471
tri 5877 5459 5889 5471 sw
rect 6418 4219 6634 4257
rect 5894 4159 5917 4170
rect 5894 4009 5918 4159
tri 5641 4003 5647 4009 ne
tri 5775 4003 5781 4009 nw
rect 5546 3872 5552 3924
rect 5604 3872 5616 3924
rect 5668 3872 5674 3924
tri 5560 3865 5567 3872 ne
rect 5567 3865 5674 3872
tri 5567 3850 5582 3865 ne
rect 5582 3850 5674 3865
tri 5582 3843 5589 3850 ne
rect 5589 3843 5674 3850
rect 2707 3760 2759 3785
rect 2707 3683 2759 3708
rect 5421 3791 5427 3843
rect 5479 3791 5491 3843
rect 5543 3791 5549 3843
tri 5589 3838 5594 3843 ne
rect 2707 3606 2759 3631
tri 5415 3625 5421 3631 se
rect 5421 3625 5549 3791
tri 5400 3610 5415 3625 se
rect 5415 3610 5549 3625
tri 5390 3600 5400 3610 se
rect 5400 3600 5549 3610
rect 2707 3548 2759 3554
rect 4356 3591 4369 3600
rect 4356 3557 4368 3591
rect 4356 3548 4369 3557
rect 4421 3548 4433 3600
rect 4485 3548 4491 3600
rect 4595 3591 4833 3600
rect 4595 3557 4607 3591
rect 4641 3557 4682 3591
rect 4716 3557 4757 3591
rect 4791 3557 4832 3591
rect 4595 3548 4833 3557
rect 4885 3548 4897 3600
rect 4949 3591 5103 3600
tri 5387 3597 5390 3600 se
rect 5390 3597 5407 3600
rect 4949 3557 4982 3591
rect 5016 3557 5057 3591
rect 5091 3557 5103 3591
rect 4949 3548 5103 3557
rect 5216 3591 5407 3597
rect 5216 3557 5228 3591
rect 5262 3557 5320 3591
rect 5354 3557 5407 3591
rect 5216 3548 5407 3557
rect 5459 3548 5491 3600
rect 5543 3548 5549 3600
rect 2627 3487 2679 3499
rect 2627 3429 2679 3435
rect 4300 3429 4306 3481
rect 4358 3429 4370 3481
rect 4422 3429 4428 3481
tri 4312 3420 4321 3429 ne
rect 4321 3420 4346 3429
tri 4321 3399 4342 3420 ne
rect 4342 3399 4346 3420
tri 4342 3395 4346 3399 ne
rect 4392 3420 4417 3429
tri 4417 3420 4426 3429 nw
rect 4392 3399 4396 3420
tri 4396 3399 4417 3420 nw
tri 4392 3395 4396 3399 nw
tri 3853 3365 3856 3368 se
tri 3842 3354 3853 3365 se
rect 3853 3354 3856 3365
tri 3811 3323 3842 3354 se
rect 3842 3323 3856 3354
tri 3786 3298 3811 3323 se
rect 3811 3298 3856 3323
tri 3752 3264 3786 3298 se
rect 3786 3264 3856 3298
tri 3735 3247 3752 3264 se
rect 3752 3247 3856 3264
tri 3701 3213 3735 3247 se
rect 3735 3213 3856 3247
tri 3696 3208 3701 3213 se
rect 3701 3208 3856 3213
tri 3659 3171 3696 3208 se
rect 3696 3171 3856 3208
tri 3652 3164 3659 3171 se
rect 3659 3164 3856 3171
tri 4056 3323 4086 3353 sw
rect 4056 3298 4086 3323
tri 4086 3298 4111 3323 sw
rect 4499 3315 4551 3467
tri 4643 3420 4658 3435 se
tri 4624 3401 4643 3420 se
rect 4643 3401 4658 3420
tri 4704 3420 4719 3435 sw
rect 4704 3401 4719 3420
tri 4719 3401 4738 3420 sw
rect 4624 3349 4630 3401
rect 4682 3349 4694 3401
rect 4746 3349 4752 3401
tri 4624 3323 4650 3349 ne
rect 4650 3323 4658 3349
tri 4650 3315 4658 3323 ne
rect 4704 3323 4712 3349
tri 4712 3323 4738 3349 nw
tri 4704 3315 4712 3323 nw
rect 4811 3315 4863 3467
tri 4955 3420 4970 3435 se
tri 4936 3401 4955 3420 se
rect 4955 3401 4970 3420
tri 5016 3420 5029 3433 sw
rect 5016 3401 5029 3420
tri 5029 3401 5048 3420 sw
rect 4920 3349 4926 3401
rect 4978 3349 4990 3401
rect 5042 3349 5048 3401
tri 4936 3323 4962 3349 ne
rect 4962 3323 4970 3349
tri 4962 3317 4968 3323 ne
rect 4968 3317 4970 3323
rect 5016 3323 5022 3349
tri 5022 3323 5048 3349 nw
tri 5016 3317 5022 3323 nw
tri 4968 3315 4970 3317 ne
rect 5123 3315 5175 3467
tri 5267 3420 5282 3435 se
tri 5248 3401 5267 3420 se
rect 5267 3401 5282 3420
tri 5328 3420 5343 3435 sw
rect 5328 3401 5343 3420
tri 5343 3401 5362 3420 sw
rect 5245 3349 5251 3401
rect 5303 3349 5315 3401
rect 5367 3349 5373 3401
tri 5248 3323 5274 3349 ne
rect 5274 3323 5282 3349
tri 5274 3315 5282 3323 ne
rect 5328 3323 5336 3349
tri 5336 3323 5362 3349 nw
tri 5328 3315 5336 3323 nw
rect 5435 3315 5487 3467
tri 5579 3420 5594 3435 se
rect 5594 3420 5674 3843
tri 5560 3401 5579 3420 se
rect 5579 3401 5674 3420
rect 5546 3349 5552 3401
rect 5604 3349 5616 3401
rect 5668 3349 5674 3401
tri 5560 3323 5586 3349 ne
rect 5586 3323 5594 3349
tri 5586 3315 5594 3323 ne
rect 5640 3323 5648 3349
tri 5648 3323 5674 3349 nw
tri 5640 3315 5648 3323 nw
rect 5747 3315 5799 3467
rect 4056 3264 4111 3298
tri 4111 3264 4145 3298 sw
rect 4056 3247 4145 3264
tri 4145 3247 4162 3264 sw
rect 4499 3251 4551 3263
rect 4056 3213 4162 3247
tri 4162 3213 4196 3247 sw
rect 4056 3208 4196 3213
tri 4196 3208 4201 3213 sw
rect 4056 3171 4201 3208
tri 4201 3171 4238 3208 sw
rect 4499 3193 4551 3199
rect 4811 3251 4863 3263
rect 4811 3193 4863 3199
rect 5123 3251 5175 3263
rect 5123 3193 5175 3199
rect 5435 3251 5487 3263
rect 5435 3193 5487 3199
rect 5747 3251 5799 3263
rect 5747 3193 5799 3199
rect 4056 3164 4238 3171
tri 4238 3164 4245 3171 sw
rect 4056 3142 4245 3164
tri 4245 3142 4267 3164 sw
rect 4056 3137 4267 3142
tri 4267 3137 4272 3142 sw
rect 2889 3136 6623 3137
rect 2889 3118 5629 3136
tri 2855 3108 2865 3118 ne
rect 2865 3108 5629 3118
tri 2865 3096 2877 3108 ne
rect 2877 3096 5629 3108
tri 2877 3095 2878 3096 ne
rect 2878 3095 5629 3096
tri 2878 3091 2882 3095 ne
rect 2882 3091 5629 3095
tri 2882 3084 2889 3091 ne
rect 2889 3084 5629 3091
rect 5681 3084 5696 3136
rect 5748 3084 5763 3136
rect 5815 3084 5830 3136
rect 5882 3084 5897 3136
rect 5949 3084 5964 3136
rect 6016 3084 6031 3136
rect 6083 3084 6098 3136
rect 6150 3084 6165 3136
rect 6217 3084 6232 3136
rect 6284 3084 6299 3136
rect 6351 3084 6366 3136
rect 6418 3084 6433 3136
rect 6485 3084 6499 3136
rect 6551 3084 6565 3136
rect 6617 3084 6623 3136
rect 2889 3061 6623 3084
tri 6623 3061 6653 3091 sw
rect 2889 3057 6653 3061
tri 6653 3057 6657 3061 sw
rect 2889 3048 6623 3057
rect 2889 2996 5629 3048
rect 5681 2996 5696 3048
rect 5748 2996 5763 3048
rect 5815 2996 5830 3048
rect 5882 2996 5897 3048
rect 5949 2996 5964 3048
rect 6016 2996 6031 3048
rect 6083 2996 6098 3048
rect 6150 2996 6165 3048
rect 6217 2996 6232 3048
rect 6284 2996 6299 3048
rect 6351 2996 6366 3048
rect 6418 2996 6433 3048
rect 6485 2996 6499 3048
rect 6551 2996 6565 3048
rect 6617 2996 6623 3048
rect 2373 2864 2425 2876
rect 2373 2806 2425 2812
rect 3604 2806 3610 2858
rect 3662 2806 3674 2858
rect 3726 2806 3910 2858
rect 2293 2703 2345 2761
tri 3263 2703 3269 2709 se
rect 2213 2681 2265 2693
tri 3235 2675 3263 2703 se
rect 3263 2675 3269 2703
tri 3315 2675 3349 2709 sw
rect 3706 2703 3712 2755
rect 3764 2703 3776 2755
rect 3828 2703 3834 2755
rect 2213 2623 2265 2629
tri 2955 2623 2957 2625 se
tri 2954 2622 2955 2623 se
rect 2955 2622 2957 2623
tri 2949 2617 2954 2622 se
rect 2954 2617 2957 2622
tri 2923 2591 2949 2617 se
rect 2949 2591 2957 2617
tri 3003 2623 3005 2625 sw
rect 3226 2623 3232 2675
rect 3284 2623 3296 2675
rect 3348 2623 3354 2675
rect 4264 2672 4316 2854
rect 3003 2622 3005 2623
tri 3005 2622 3006 2623 sw
tri 3235 2622 3236 2623 ne
rect 3236 2622 3269 2623
rect 3003 2617 3006 2622
tri 3006 2617 3011 2622 sw
tri 3236 2617 3241 2622 ne
rect 3241 2617 3269 2622
rect 3003 2591 3011 2617
tri 3011 2591 3037 2617 sw
tri 3241 2591 3267 2617 ne
rect 3267 2591 3269 2617
rect 2917 2539 2923 2591
rect 2975 2539 2987 2591
rect 3039 2539 3045 2591
tri 3267 2589 3269 2591 ne
rect 3315 2617 3343 2623
tri 3343 2617 3349 2623 nw
tri 3315 2589 3343 2617 nw
rect 4264 2608 4316 2620
rect 4264 2542 4316 2556
rect 4577 2737 4629 2854
rect 4914 2809 4920 2861
rect 4972 2809 4984 2861
rect 5036 2809 5042 2861
tri 5042 2855 5048 2861 sw
tri 5970 2855 5976 2861 se
rect 5976 2809 5982 2861
rect 6034 2809 6046 2861
rect 6098 2809 6104 2861
rect 5874 2706 5880 2758
rect 5932 2706 5944 2758
rect 5996 2706 6002 2758
tri 6387 2706 6393 2712 se
rect 4577 2673 4629 2685
tri 6359 2678 6387 2706 se
rect 6387 2678 6393 2706
tri 6439 2678 6473 2712 sw
rect 6354 2626 6360 2678
rect 6412 2626 6424 2678
rect 6476 2626 6482 2678
tri 6703 2626 6705 2628 se
tri 6359 2622 6363 2626 ne
rect 6363 2622 6393 2626
rect 4577 2542 4629 2621
tri 6363 2617 6368 2622 ne
rect 6368 2617 6393 2622
tri 6368 2594 6391 2617 ne
rect 6391 2594 6393 2617
tri 6391 2592 6393 2594 ne
rect 6439 2617 6464 2626
tri 6464 2617 6473 2626 nw
tri 6694 2617 6703 2626 se
rect 6703 2617 6705 2626
rect 6439 2594 6441 2617
tri 6441 2594 6464 2617 nw
tri 6671 2594 6694 2617 se
rect 6694 2594 6705 2617
tri 6751 2622 6757 2628 sw
rect 6751 2617 6757 2622
tri 6757 2617 6762 2622 sw
rect 6751 2594 6762 2617
tri 6762 2594 6785 2617 sw
tri 6439 2592 6441 2594 nw
rect 6663 2542 6669 2594
rect 6721 2542 6733 2594
rect 6785 2542 6791 2594
tri 2099 2487 2130 2518 se
rect 2130 2487 2185 2518
rect 2057 2435 2063 2487
rect 2115 2435 2127 2487
rect 2179 2435 2185 2487
rect 2981 2448 2987 2500
rect 3039 2448 3053 2500
rect 3105 2448 3111 2500
rect 4291 2451 4297 2503
rect 4349 2451 4363 2503
rect 4415 2451 4421 2503
rect 4969 2493 5021 2499
tri 4935 2435 4942 2442 ne
rect 4942 2441 4969 2442
rect 6597 2451 6603 2503
rect 6655 2451 6669 2503
rect 6721 2451 6727 2503
rect 4942 2435 5021 2441
tri 4942 2408 4969 2435 ne
rect 4969 2429 5021 2435
rect 1973 2383 2025 2395
tri 5021 2425 5038 2442 nw
rect 1973 2325 2025 2331
rect 4116 2325 4122 2377
rect 4174 2325 4186 2377
rect 4238 2373 4244 2377
tri 4244 2373 4248 2377 sw
rect 4238 2350 4248 2373
tri 4248 2350 4271 2373 sw
rect 4969 2371 5021 2377
tri 6844 2371 6850 2377 se
rect 6850 2371 6902 8202
tri 7397 8118 7431 8152 se
rect 6944 7937 7576 7938
rect 6944 7885 6950 7937
rect 7002 7886 7046 7937
rect 7098 7886 7576 7937
rect 7006 7885 7046 7886
rect 7098 7885 7132 7886
rect 6944 7852 6972 7885
rect 7006 7852 7052 7885
rect 7086 7852 7132 7885
rect 7166 7852 7212 7886
rect 7246 7852 7292 7886
rect 7326 7852 7372 7886
rect 7406 7852 7451 7886
rect 7485 7852 7530 7886
rect 7564 7852 7576 7886
rect 6944 7846 7576 7852
rect 7710 7881 7756 7893
rect 7710 7847 7716 7881
rect 7750 7847 7756 7881
rect 6944 7841 7121 7846
rect 6944 7789 6950 7841
rect 7002 7789 7046 7841
rect 7098 7829 7121 7841
tri 7121 7829 7138 7846 nw
rect 7618 7829 7664 7841
rect 7098 7789 7104 7829
tri 7104 7812 7121 7829 nw
rect 6944 7738 7104 7789
rect 7618 7795 7624 7829
rect 7658 7795 7664 7829
tri 7104 7738 7136 7770 sw
tri 7586 7738 7618 7770 se
rect 7618 7738 7664 7795
rect 6944 7736 7136 7738
tri 7136 7736 7138 7738 sw
tri 7584 7736 7586 7738 se
rect 7586 7736 7624 7738
rect 6944 7730 7624 7736
rect 6944 7696 7144 7730
rect 7178 7696 7222 7730
rect 7256 7696 7299 7730
rect 7333 7696 7376 7730
rect 7410 7696 7453 7730
rect 7487 7696 7530 7730
rect 7564 7704 7624 7730
rect 7658 7704 7664 7738
rect 7564 7696 7664 7704
rect 6944 7690 7664 7696
rect 6944 7665 7113 7690
tri 7113 7665 7138 7690 nw
tri 7584 7665 7609 7690 ne
rect 7609 7665 7664 7690
rect 6944 7612 7104 7665
tri 7104 7656 7113 7665 nw
tri 7609 7656 7618 7665 ne
rect 7618 7646 7664 7665
tri 7104 7612 7106 7614 sw
rect 7618 7612 7624 7646
rect 7658 7612 7664 7646
rect 6944 7593 7106 7612
tri 7106 7593 7125 7612 sw
rect 7618 7600 7664 7612
rect 7710 7809 7756 7847
rect 7710 7775 7716 7809
rect 7750 7775 7756 7809
rect 7710 7737 7756 7775
rect 7710 7703 7716 7737
rect 7750 7703 7756 7737
rect 7710 7665 7756 7703
rect 7710 7631 7716 7665
rect 7750 7631 7756 7665
rect 7710 7593 7756 7631
rect 6944 7580 7125 7593
tri 7125 7580 7138 7593 sw
rect 6944 7574 7448 7580
rect 6944 7540 6972 7574
rect 7006 7540 7058 7574
rect 7092 7540 7144 7574
rect 7178 7540 7230 7574
rect 7264 7540 7316 7574
rect 7350 7540 7402 7574
rect 7436 7540 7448 7574
rect 6944 7534 7448 7540
rect 7710 7559 7716 7593
rect 7750 7559 7756 7593
rect 6944 7521 7125 7534
tri 7125 7521 7138 7534 nw
rect 7710 7521 7756 7559
rect 6944 7504 7108 7521
tri 7108 7504 7125 7521 nw
rect 7618 7504 7664 7516
rect 6944 7286 7104 7504
tri 7104 7500 7108 7504 nw
rect 7618 7470 7624 7504
rect 7658 7470 7664 7504
rect 7618 7431 7664 7470
rect 7132 7418 7576 7424
rect 7132 7384 7144 7418
rect 7178 7384 7222 7418
rect 7256 7384 7299 7418
rect 7333 7384 7376 7418
rect 7410 7384 7453 7418
rect 7487 7384 7530 7418
rect 7564 7384 7576 7418
rect 7132 7378 7576 7384
tri 7442 7377 7443 7378 ne
rect 7443 7377 7576 7378
tri 7443 7358 7462 7377 ne
rect 7462 7358 7576 7377
tri 7462 7344 7476 7358 ne
rect 7476 7339 7576 7358
tri 7104 7286 7120 7302 sw
rect 7476 7287 7500 7339
rect 7552 7287 7576 7339
rect 6944 7285 7120 7286
tri 7120 7285 7121 7286 sw
rect 6944 7268 7121 7285
tri 7121 7268 7138 7285 sw
rect 6944 7262 7448 7268
rect 6944 7228 6972 7262
rect 7006 7228 7058 7262
rect 7092 7228 7144 7262
rect 7178 7228 7230 7262
rect 7264 7228 7316 7262
rect 7350 7228 7402 7262
rect 7436 7228 7448 7262
rect 6944 7222 7448 7228
rect 7476 7249 7576 7287
rect 6944 7211 7127 7222
tri 7127 7211 7138 7222 nw
rect 6944 6989 7104 7211
tri 7104 7188 7127 7211 nw
rect 7476 7197 7500 7249
rect 7552 7197 7576 7249
tri 7467 7137 7476 7146 se
rect 7476 7137 7576 7197
tri 7442 7112 7467 7137 se
rect 7467 7112 7576 7137
rect 7132 7106 7576 7112
rect 7132 7072 7144 7106
rect 7178 7072 7222 7106
rect 7256 7072 7299 7106
rect 7333 7072 7376 7106
rect 7410 7072 7453 7106
rect 7487 7072 7530 7106
rect 7564 7072 7576 7106
rect 7132 7066 7576 7072
tri 7442 7063 7445 7066 ne
rect 7445 7063 7576 7066
tri 7445 7051 7457 7063 ne
rect 7457 7051 7576 7063
tri 7457 7045 7463 7051 ne
rect 7463 7045 7576 7051
tri 7463 7032 7476 7045 ne
tri 7104 6989 7105 6990 sw
rect 6944 6956 7105 6989
tri 7105 6956 7138 6989 sw
rect 6944 6950 7448 6956
rect 6944 6916 6972 6950
rect 7006 6916 7058 6950
rect 7092 6916 7144 6950
rect 7178 6916 7230 6950
rect 7264 6916 7316 6950
rect 7350 6916 7402 6950
rect 7436 6916 7448 6950
rect 6944 6910 7448 6916
rect 6944 6881 7109 6910
tri 7109 6881 7138 6910 nw
rect 6944 6659 7104 6881
tri 7104 6876 7109 6881 nw
tri 7449 6807 7476 6834 se
rect 7476 6807 7576 7045
tri 7443 6801 7449 6807 se
rect 7449 6801 7576 6807
tri 7442 6800 7443 6801 se
rect 7443 6800 7576 6801
rect 7132 6794 7576 6800
rect 7132 6760 7144 6794
rect 7178 6760 7222 6794
rect 7256 6760 7299 6794
rect 7333 6760 7376 6794
rect 7410 6760 7453 6794
rect 7487 6760 7530 6794
rect 7564 6760 7576 6794
rect 7132 6754 7576 6760
tri 7442 6733 7463 6754 ne
rect 7463 6733 7576 6754
tri 7463 6729 7467 6733 ne
rect 7467 6729 7576 6733
tri 7467 6720 7476 6729 ne
tri 7104 6659 7123 6678 sw
rect 6944 6657 7123 6659
tri 7123 6657 7125 6659 sw
rect 6944 6644 7125 6657
tri 7125 6644 7138 6657 sw
rect 6944 6638 7448 6644
rect 6944 6604 6972 6638
rect 7006 6604 7058 6638
rect 7092 6604 7144 6638
rect 7178 6604 7230 6638
rect 7264 6604 7316 6638
rect 7350 6604 7402 6638
rect 7436 6604 7448 6638
rect 6944 6598 7448 6604
rect 6944 6595 7135 6598
tri 7135 6595 7138 6598 nw
rect 6944 6585 7125 6595
tri 7125 6585 7135 6595 nw
rect 6944 6363 7104 6585
tri 7104 6564 7125 6585 nw
tri 7465 6511 7476 6522 se
rect 7476 6511 7576 6729
tri 7442 6488 7465 6511 se
rect 7465 6488 7576 6511
rect 7132 6482 7576 6488
rect 7132 6448 7144 6482
rect 7178 6448 7222 6482
rect 7256 6448 7299 6482
rect 7333 6448 7376 6482
rect 7410 6448 7453 6482
rect 7487 6448 7530 6482
rect 7564 6448 7576 6482
rect 7132 6442 7576 6448
rect 7618 7397 7624 7431
rect 7658 7397 7664 7431
rect 7618 7358 7664 7397
rect 7618 7324 7624 7358
rect 7658 7324 7664 7358
rect 7618 7285 7664 7324
rect 7618 7251 7624 7285
rect 7658 7251 7664 7285
rect 7618 7211 7664 7251
rect 7618 7177 7624 7211
rect 7658 7177 7664 7211
rect 7618 7137 7664 7177
rect 7618 7103 7624 7137
rect 7658 7103 7664 7137
rect 7618 7063 7664 7103
rect 7618 7039 7624 7063
rect 7658 7045 7664 7063
rect 7710 7487 7716 7521
rect 7750 7487 7756 7521
rect 7710 7449 7756 7487
rect 7710 7415 7716 7449
rect 7750 7415 7756 7449
rect 7710 7377 7756 7415
rect 7710 7343 7716 7377
rect 7750 7343 7756 7377
rect 7710 7305 7756 7343
rect 7710 7271 7716 7305
rect 7750 7271 7756 7305
rect 7710 7233 7756 7271
rect 7710 7199 7716 7233
rect 7750 7199 7756 7233
rect 7710 7161 7756 7199
rect 7710 7127 7716 7161
rect 7750 7127 7756 7161
rect 7710 7089 7756 7127
rect 7710 7055 7716 7089
rect 7750 7055 7756 7089
tri 7664 7045 7670 7051 sw
rect 7658 7039 7670 7045
rect 7618 6975 7624 6987
rect 7658 6975 7670 6987
rect 7618 6917 7670 6923
rect 7618 6915 7664 6917
rect 7618 6881 7624 6915
rect 7658 6881 7664 6915
tri 7664 6911 7670 6917 nw
rect 7710 7017 7756 7055
rect 7710 6983 7716 7017
rect 7750 6983 7756 7017
rect 7710 6945 7756 6983
rect 7710 6911 7716 6945
rect 7750 6911 7756 6945
rect 7618 6841 7664 6881
rect 7618 6807 7624 6841
rect 7658 6807 7664 6841
rect 7618 6767 7664 6807
rect 7618 6733 7624 6767
rect 7658 6733 7664 6767
rect 7618 6693 7664 6733
rect 7618 6659 7624 6693
rect 7658 6659 7664 6693
rect 7618 6619 7664 6659
rect 7618 6585 7624 6619
rect 7658 6585 7664 6619
rect 7618 6545 7664 6585
rect 7618 6511 7624 6545
rect 7658 6511 7664 6545
rect 7618 6471 7664 6511
rect 7618 6437 7624 6471
rect 7658 6437 7664 6471
tri 7594 6407 7618 6431 se
rect 7618 6407 7664 6437
tri 7584 6397 7594 6407 se
rect 7594 6397 7664 6407
tri 7552 6366 7583 6397 se
rect 7583 6366 7624 6397
tri 7104 6363 7107 6366 sw
tri 7549 6363 7552 6366 se
rect 7552 6363 7624 6366
rect 7658 6363 7664 6397
rect 6944 6335 7107 6363
tri 7107 6335 7135 6363 sw
tri 7537 6351 7549 6363 se
rect 7549 6351 7664 6363
tri 7531 6345 7537 6351 se
rect 7537 6345 7664 6351
rect 7710 6873 7756 6911
rect 7710 6839 7716 6873
rect 7750 6839 7756 6873
rect 7710 6801 7756 6839
rect 7710 6767 7716 6801
rect 7750 6767 7756 6801
rect 7710 6729 7756 6767
rect 7710 6695 7716 6729
rect 7750 6695 7756 6729
rect 7710 6657 7756 6695
rect 7710 6623 7716 6657
rect 7750 6623 7756 6657
rect 7710 6585 7756 6623
rect 7710 6551 7716 6585
rect 7750 6551 7756 6585
rect 7710 6513 7756 6551
rect 7710 6479 7716 6513
rect 7750 6479 7756 6513
rect 7710 6441 7756 6479
rect 7710 6407 7716 6441
rect 7750 6407 7756 6441
rect 7710 6369 7756 6407
tri 7524 6338 7531 6345 se
rect 7531 6338 7595 6345
rect 7524 6335 7595 6338
tri 7595 6335 7605 6345 nw
rect 7710 6335 7716 6369
rect 7750 6335 7756 6369
rect 6944 6332 7135 6335
tri 7135 6332 7138 6335 sw
rect 7524 6332 7592 6335
tri 7592 6332 7595 6335 nw
rect 6944 6326 7448 6332
rect 6944 6292 6972 6326
rect 7006 6292 7058 6326
rect 7092 6292 7144 6326
rect 7178 6292 7230 6326
rect 7264 6292 7316 6326
rect 7350 6292 7402 6326
rect 7436 6292 7448 6326
rect 6944 6286 7448 6292
rect 6944 6279 7131 6286
tri 7131 6279 7138 6286 nw
rect 6944 6267 7119 6279
tri 7119 6267 7131 6279 nw
rect 6944 6127 7104 6267
tri 7104 6252 7119 6267 nw
tri 7509 6195 7524 6210 se
rect 7524 6195 7576 6332
tri 7576 6316 7592 6332 nw
rect 7710 6297 7756 6335
tri 7490 6176 7509 6195 se
rect 7509 6176 7576 6195
rect 7132 6170 7576 6176
rect 7132 6136 7144 6170
rect 7178 6136 7222 6170
rect 7256 6136 7299 6170
rect 7333 6136 7376 6170
rect 7410 6136 7453 6170
rect 7487 6136 7530 6170
rect 7564 6136 7576 6170
rect 7615 6267 7667 6279
rect 7615 6262 7624 6267
rect 7658 6262 7667 6267
rect 7615 6198 7667 6210
rect 7615 6140 7667 6146
rect 7710 6263 7716 6297
rect 7750 6263 7756 6297
rect 7710 6225 7756 6263
rect 7710 6191 7716 6225
rect 7750 6191 7756 6225
rect 7710 6153 7756 6191
rect 7132 6130 7576 6136
rect 6996 6075 7052 6127
rect 7710 6119 7716 6153
rect 7750 6119 7756 6153
tri 7104 6081 7123 6100 sw
rect 7710 6081 7756 6119
rect 7104 6075 7123 6081
rect 6944 6066 7123 6075
tri 7123 6066 7138 6081 sw
rect 6944 6060 7576 6066
rect 6944 6057 6972 6060
rect 7006 6026 7052 6060
rect 7086 6057 7132 6060
rect 7104 6026 7132 6057
rect 7166 6026 7212 6060
rect 7246 6026 7292 6060
rect 7326 6026 7372 6060
rect 7406 6026 7451 6060
rect 7485 6026 7530 6060
rect 7564 6026 7576 6060
rect 6996 6005 7052 6026
rect 7104 6020 7576 6026
rect 7710 6047 7716 6081
rect 7750 6047 7756 6081
rect 7104 6009 7127 6020
tri 7127 6009 7138 6020 nw
rect 7104 6005 7121 6009
rect 6944 6003 7121 6005
tri 7121 6003 7127 6009 nw
rect 7618 6003 7664 6015
rect 6944 5987 7104 6003
rect 6996 5935 7052 5987
tri 7104 5986 7121 6003 nw
rect 7618 5969 7624 6003
rect 7658 5969 7664 6003
tri 7104 5937 7111 5944 sw
tri 7611 5937 7618 5944 se
rect 7618 5937 7664 5969
rect 7104 5935 7111 5937
rect 6944 5917 7111 5935
rect 6996 5865 7052 5917
rect 7104 5916 7111 5917
tri 7111 5916 7132 5937 sw
tri 7590 5916 7611 5937 se
rect 7611 5916 7664 5937
rect 7104 5910 7132 5916
tri 7132 5910 7138 5916 sw
tri 7584 5910 7590 5916 se
rect 7590 5910 7624 5916
rect 7104 5904 7624 5910
rect 7104 5870 7144 5904
rect 7178 5870 7222 5904
rect 7256 5870 7299 5904
rect 7333 5870 7376 5904
rect 7410 5870 7453 5904
rect 7487 5870 7530 5904
rect 7564 5882 7624 5904
rect 7658 5882 7664 5916
rect 7710 6009 7756 6047
rect 7710 5975 7716 6009
rect 7750 5975 7756 6009
rect 7710 5937 7756 5975
tri 7706 5910 7710 5914 se
rect 7710 5910 7716 5937
rect 7564 5870 7664 5882
rect 7104 5865 7664 5870
rect 6944 5864 7664 5865
rect 6944 5847 7105 5864
rect 6996 5795 7052 5847
rect 7104 5831 7105 5847
tri 7105 5831 7138 5864 nw
tri 7584 5831 7617 5864 ne
rect 7617 5831 7664 5864
tri 7104 5830 7105 5831 nw
tri 7617 5830 7618 5831 ne
rect 6944 5782 7104 5795
rect 7618 5828 7664 5831
rect 7618 5794 7624 5828
rect 7658 5794 7664 5828
tri 7104 5782 7110 5788 sw
rect 7618 5782 7664 5794
tri 7704 5908 7706 5910 se
rect 7706 5908 7716 5910
rect 7704 5903 7716 5908
rect 7750 5903 7756 5937
rect 7704 5902 7756 5903
rect 7704 5835 7716 5850
rect 7750 5835 7756 5850
rect 6944 5777 7110 5782
rect 6996 5748 7052 5777
rect 7104 5759 7110 5777
tri 7110 5759 7133 5782 sw
rect 7704 5768 7716 5783
rect 7750 5768 7756 5783
rect 7104 5754 7133 5759
tri 7133 5754 7138 5759 sw
rect 7104 5748 7448 5754
rect 7006 5725 7052 5748
rect 7104 5725 7144 5748
rect 6944 5714 6972 5725
rect 7006 5714 7058 5725
rect 7092 5714 7144 5725
rect 7178 5714 7230 5748
rect 7264 5714 7316 5748
rect 7350 5714 7402 5748
rect 7436 5714 7448 5748
rect 6944 5708 7448 5714
rect 6944 5706 7117 5708
rect 6996 5654 7052 5706
rect 7104 5687 7117 5706
tri 7117 5687 7138 5708 nw
rect 7704 5700 7716 5716
rect 7750 5700 7756 5716
tri 7104 5674 7117 5687 nw
rect 6944 5635 7104 5654
rect 6996 5583 7052 5635
rect 7618 5670 7664 5682
rect 7618 5636 7624 5670
rect 7658 5636 7664 5670
rect 6944 5564 7104 5583
rect 6996 5512 7052 5564
rect 7132 5592 7576 5598
rect 7132 5558 7144 5592
rect 7178 5558 7222 5592
rect 7256 5558 7299 5592
rect 7333 5558 7376 5592
rect 7410 5558 7453 5592
rect 7487 5558 7530 5592
rect 7564 5558 7576 5592
rect 7132 5552 7576 5558
tri 7442 5543 7451 5552 ne
rect 7451 5543 7576 5552
tri 7451 5524 7470 5543 ne
rect 7470 5524 7576 5543
tri 7470 5518 7476 5524 ne
rect 6944 5471 7104 5512
tri 7104 5471 7109 5476 sw
rect 6944 5459 7109 5471
tri 7109 5459 7121 5471 sw
rect 6944 5451 7121 5459
tri 7121 5451 7129 5459 sw
rect 6944 5442 7129 5451
tri 7129 5442 7138 5451 sw
rect 6944 5436 7448 5442
rect 6944 5402 6972 5436
rect 7006 5402 7058 5436
rect 7092 5402 7144 5436
rect 7178 5402 7230 5436
rect 7264 5402 7316 5436
rect 7350 5402 7402 5436
rect 7436 5402 7448 5436
rect 6944 5396 7448 5402
rect 6944 5378 7120 5396
tri 7120 5378 7138 5396 nw
rect 6944 5159 7104 5378
tri 7104 5362 7120 5378 nw
tri 7461 5305 7476 5320 se
rect 7476 5305 7576 5524
tri 7442 5286 7461 5305 se
rect 7461 5286 7576 5305
rect 7132 5280 7576 5286
rect 7132 5246 7144 5280
rect 7178 5246 7222 5280
rect 7256 5246 7299 5280
rect 7333 5246 7376 5280
rect 7410 5246 7453 5280
rect 7487 5246 7530 5280
rect 7564 5246 7576 5280
rect 7132 5240 7576 5246
tri 7442 5232 7450 5240 ne
rect 7450 5232 7524 5240
tri 7450 5206 7476 5232 ne
rect 7476 5188 7524 5232
tri 7104 5159 7109 5164 sw
rect 6944 5130 7109 5159
tri 7109 5130 7138 5159 sw
rect 7476 5150 7576 5188
rect 6944 5124 7448 5130
rect 6944 5090 6972 5124
rect 7006 5090 7058 5124
rect 7092 5090 7144 5124
rect 7178 5090 7230 5124
rect 7264 5090 7316 5124
rect 7350 5090 7402 5124
rect 7436 5090 7448 5124
rect 6944 5084 7448 5090
rect 7476 5098 7524 5150
rect 6944 5052 7106 5084
tri 7106 5052 7138 5084 nw
rect 6944 4833 7104 5052
tri 7104 5050 7106 5052 nw
tri 7470 5002 7476 5008 se
rect 7476 5002 7576 5098
tri 7464 4996 7470 5002 se
rect 7470 4996 7576 5002
tri 7447 4979 7464 4996 se
rect 7464 4979 7576 4996
tri 7442 4974 7447 4979 se
rect 7447 4974 7576 4979
rect 7132 4968 7576 4974
rect 7132 4934 7144 4968
rect 7178 4934 7222 4968
rect 7256 4934 7299 4968
rect 7333 4934 7376 4968
rect 7410 4934 7453 4968
rect 7487 4934 7530 4968
rect 7564 4934 7576 4968
rect 7132 4928 7576 4934
tri 7442 4906 7464 4928 ne
rect 7464 4906 7576 4928
tri 7464 4894 7476 4906 ne
tri 7104 4833 7123 4852 sw
rect 6944 4818 7123 4833
tri 7123 4818 7138 4833 sw
rect 6944 4812 7448 4818
rect 6944 4778 6972 4812
rect 7006 4778 7058 4812
rect 7092 4778 7144 4812
rect 7178 4778 7230 4812
rect 7264 4778 7316 4812
rect 7350 4778 7402 4812
rect 7436 4778 7448 4812
rect 6944 4772 7448 4778
rect 6944 4759 7125 4772
tri 7125 4759 7138 4772 nw
rect 6944 4741 7107 4759
tri 7107 4741 7125 4759 nw
rect 6944 4537 7104 4741
tri 7104 4738 7107 4741 nw
tri 7465 4685 7476 4696 se
rect 7476 4685 7576 4906
tri 7448 4668 7465 4685 se
rect 7465 4668 7576 4685
tri 7442 4662 7448 4668 se
rect 7448 4662 7576 4668
rect 7132 4656 7576 4662
rect 7132 4622 7144 4656
rect 7178 4622 7222 4656
rect 7256 4622 7299 4656
rect 7333 4622 7376 4656
rect 7410 4622 7453 4656
rect 7487 4622 7530 4656
rect 7564 4622 7576 4656
rect 7132 4616 7576 4622
rect 7618 5597 7664 5636
rect 7618 5563 7624 5597
rect 7658 5563 7664 5597
rect 7618 5524 7664 5563
rect 7618 5490 7624 5524
rect 7658 5490 7664 5524
rect 7704 5632 7716 5648
rect 7750 5632 7756 5648
rect 7704 5577 7756 5580
rect 7704 5564 7716 5577
rect 7750 5564 7756 5577
rect 7704 5506 7756 5512
tri 7704 5505 7705 5506 ne
rect 7705 5505 7756 5506
tri 7705 5500 7710 5505 ne
rect 7618 5451 7664 5490
rect 7618 5417 7624 5451
rect 7658 5417 7664 5451
rect 7618 5378 7664 5417
rect 7618 5344 7624 5378
rect 7658 5344 7664 5378
rect 7618 5305 7664 5344
rect 7618 5271 7624 5305
rect 7658 5271 7664 5305
rect 7618 5232 7664 5271
rect 7618 5198 7624 5232
rect 7658 5198 7664 5232
rect 7618 5159 7664 5198
rect 7618 5125 7624 5159
rect 7658 5125 7664 5159
rect 7618 5086 7664 5125
rect 7618 5052 7624 5086
rect 7658 5052 7664 5086
rect 7618 5013 7664 5052
rect 7618 4990 7624 5013
rect 7658 4996 7664 5013
rect 7710 5471 7716 5505
rect 7750 5471 7756 5505
rect 7710 5432 7756 5471
rect 7710 5398 7716 5432
rect 7750 5398 7756 5432
rect 7710 5359 7756 5398
rect 7710 5325 7716 5359
rect 7750 5325 7756 5359
rect 7710 5286 7756 5325
rect 7710 5252 7716 5286
rect 7750 5252 7756 5286
rect 7710 5213 7756 5252
rect 7710 5179 7716 5213
rect 7750 5179 7756 5213
rect 7710 5140 7756 5179
rect 7710 5106 7716 5140
rect 7750 5106 7756 5140
rect 7710 5067 7756 5106
rect 7710 5033 7716 5067
rect 7750 5033 7756 5067
tri 7664 4996 7670 5002 sw
rect 7658 4990 7670 4996
rect 7618 4926 7624 4938
rect 7658 4926 7670 4938
rect 7618 4868 7670 4874
rect 7618 4867 7664 4868
rect 7618 4833 7624 4867
rect 7658 4833 7664 4867
tri 7664 4862 7670 4868 nw
rect 7710 4994 7756 5033
rect 7710 4960 7716 4994
rect 7750 4960 7756 4994
rect 7710 4921 7756 4960
rect 7710 4887 7716 4921
rect 7750 4887 7756 4921
rect 7618 4793 7664 4833
rect 7618 4759 7624 4793
rect 7658 4759 7664 4793
rect 7618 4719 7664 4759
rect 7618 4685 7624 4719
rect 7658 4685 7664 4719
rect 7618 4645 7664 4685
rect 7618 4611 7624 4645
rect 7658 4611 7664 4645
tri 7608 4595 7618 4605 se
rect 7618 4595 7664 4611
tri 7584 4571 7608 4595 se
rect 7608 4571 7664 4595
tri 7552 4540 7583 4571 se
rect 7583 4540 7624 4571
tri 7104 4537 7107 4540 sw
tri 7549 4537 7552 4540 se
rect 7552 4537 7624 4540
rect 7658 4537 7664 4571
rect 6944 4522 7107 4537
tri 7107 4522 7122 4537 sw
tri 7537 4525 7549 4537 se
rect 7549 4525 7664 4537
tri 7534 4522 7537 4525 se
rect 7537 4522 7664 4525
rect 6944 4506 7122 4522
tri 7122 4506 7138 4522 sw
tri 7531 4519 7534 4522 se
rect 7534 4519 7664 4522
rect 7710 4848 7756 4887
rect 7710 4814 7716 4848
rect 7750 4814 7756 4848
rect 7710 4775 7756 4814
rect 7710 4741 7716 4775
rect 7750 4741 7756 4775
rect 7710 4702 7756 4741
rect 7710 4668 7716 4702
rect 7750 4668 7756 4702
rect 7710 4629 7756 4668
rect 7710 4595 7716 4629
rect 7750 4595 7756 4629
rect 7710 4556 7756 4595
rect 7710 4522 7716 4556
rect 7750 4522 7756 4556
tri 7524 4512 7531 4519 se
rect 7531 4512 7592 4519
rect 7524 4506 7592 4512
tri 7592 4506 7605 4519 nw
rect 6944 4500 7448 4506
rect 6944 4466 6972 4500
rect 7006 4466 7058 4500
rect 7092 4466 7144 4500
rect 7178 4466 7230 4500
rect 7264 4466 7316 4500
rect 7350 4466 7402 4500
rect 7436 4466 7448 4500
rect 6944 4460 7448 4466
rect 6944 4449 7127 4460
tri 7127 4449 7138 4460 nw
rect 6944 4439 7117 4449
tri 7117 4439 7127 4449 nw
rect 6944 4264 7104 4439
tri 7104 4426 7117 4439 nw
tri 7516 4376 7524 4384 se
rect 7524 4376 7576 4506
tri 7576 4490 7592 4506 nw
rect 7710 4483 7756 4522
tri 7507 4367 7516 4376 se
rect 7516 4367 7576 4376
tri 7490 4350 7507 4367 se
rect 7507 4350 7576 4367
rect 7132 4344 7576 4350
rect 7132 4310 7144 4344
rect 7178 4310 7222 4344
rect 7256 4310 7299 4344
rect 7333 4310 7376 4344
rect 7410 4310 7453 4344
rect 7487 4310 7530 4344
rect 7564 4310 7576 4344
rect 7615 4448 7667 4454
rect 7615 4384 7667 4396
rect 7615 4321 7667 4332
rect 7710 4449 7716 4483
rect 7750 4449 7756 4483
rect 7710 4410 7756 4449
rect 7710 4376 7716 4410
rect 7750 4376 7756 4410
rect 7710 4337 7756 4376
rect 7132 4304 7576 4310
rect 7710 4303 7716 4337
rect 7750 4303 7756 4337
tri 7104 4264 7114 4274 sw
rect 7710 4264 7756 4303
rect 6944 4257 7114 4264
tri 7114 4257 7121 4264 sw
rect 6944 4240 7121 4257
tri 7121 4240 7138 4257 sw
rect 6944 4234 7576 4240
rect 6944 4200 6972 4234
rect 7006 4200 7052 4234
rect 7086 4200 7132 4234
rect 7166 4200 7212 4234
rect 7246 4200 7292 4234
rect 7326 4200 7372 4234
rect 7406 4200 7451 4234
rect 7485 4200 7530 4234
rect 7564 4200 7576 4234
rect 6944 4194 7576 4200
rect 7710 4230 7716 4264
rect 7750 4230 7756 4264
rect 6944 4191 7135 4194
tri 7135 4191 7138 4194 nw
rect 7710 4191 7756 4230
rect 6944 4177 7121 4191
tri 7121 4177 7135 4191 nw
rect 7618 4177 7664 4189
rect 6944 4170 7114 4177
tri 7114 4170 7121 4177 nw
rect 6944 4099 7104 4170
tri 7104 4160 7114 4170 nw
rect 7618 4143 7624 4177
rect 7658 4143 7664 4177
tri 7104 4099 7123 4118 sw
tri 7599 4099 7618 4118 se
rect 7618 4099 7664 4143
rect 6944 4084 7123 4099
tri 7123 4084 7138 4099 sw
tri 7584 4084 7599 4099 se
rect 7599 4084 7624 4099
rect 6944 4078 7624 4084
rect 6944 4054 7144 4078
rect 6996 4002 7052 4054
rect 7104 4044 7144 4054
rect 7178 4044 7222 4078
rect 7256 4044 7299 4078
rect 7333 4044 7376 4078
rect 7410 4044 7453 4078
rect 7487 4044 7530 4078
rect 7564 4065 7624 4078
rect 7658 4065 7664 4099
rect 7564 4044 7664 4065
rect 7104 4038 7664 4044
rect 7104 4020 7120 4038
tri 7120 4020 7138 4038 nw
tri 7584 4020 7602 4038 ne
rect 7602 4020 7664 4038
rect 7104 4009 7109 4020
tri 7109 4009 7120 4020 nw
tri 7602 4009 7613 4020 ne
rect 7613 4009 7624 4020
tri 7104 4004 7109 4009 nw
tri 7613 4004 7618 4009 ne
rect 6944 3987 7104 4002
rect 6996 3935 7052 3987
rect 7618 3986 7624 4009
rect 7658 3986 7664 4020
rect 7618 3974 7664 3986
rect 7710 4157 7716 4191
rect 7750 4157 7756 4191
rect 7710 4118 7756 4157
rect 7710 4084 7716 4118
rect 7750 4084 7756 4118
rect 7710 4045 7756 4084
rect 7710 4011 7716 4045
rect 7750 4011 7756 4045
rect 7710 3972 7756 4011
tri 7104 3938 7128 3962 sw
rect 7710 3938 7716 3972
rect 7750 3938 7756 3972
rect 7104 3935 7128 3938
rect 6944 3928 7128 3935
tri 7128 3928 7138 3938 sw
rect 6944 3922 7448 3928
rect 6944 3920 6972 3922
rect 7006 3920 7058 3922
rect 7092 3920 7144 3922
rect 7006 3888 7052 3920
rect 7104 3888 7144 3920
rect 7178 3888 7230 3922
rect 7264 3888 7316 3922
rect 7350 3888 7402 3922
rect 7436 3888 7448 3922
rect 6996 3868 7052 3888
rect 7104 3882 7448 3888
rect 7710 3899 7756 3938
rect 7104 3868 7121 3882
rect 6944 3865 7121 3868
tri 7121 3865 7138 3882 nw
rect 7615 3871 7667 3877
rect 6944 3853 7106 3865
rect 6996 3801 7052 3853
rect 7104 3850 7106 3853
tri 7106 3850 7121 3865 nw
tri 7104 3848 7106 3850 nw
rect 6944 3786 7104 3801
rect 6996 3734 7052 3786
rect 7615 3816 7624 3819
rect 7658 3816 7667 3819
rect 7615 3807 7667 3816
rect 6944 3718 7104 3734
rect 7132 3766 7576 3772
rect 7132 3732 7144 3766
rect 7178 3732 7222 3766
rect 7256 3732 7299 3766
rect 7333 3732 7376 3766
rect 7410 3732 7453 3766
rect 7487 3732 7530 3766
rect 7564 3732 7576 3766
rect 7615 3749 7624 3755
tri 7615 3746 7618 3749 ne
rect 7132 3726 7576 3732
tri 7442 3719 7449 3726 ne
rect 7449 3719 7576 3726
rect 6996 3666 7052 3718
tri 7449 3700 7468 3719 ne
rect 7468 3700 7576 3719
tri 7468 3692 7476 3700 ne
rect 6944 3646 7104 3666
tri 7104 3646 7108 3650 sw
rect 6944 3625 7108 3646
tri 7108 3625 7129 3646 sw
rect 6944 3616 7129 3625
tri 7129 3616 7138 3625 sw
rect 6944 3610 7448 3616
rect 6944 3576 6972 3610
rect 7006 3576 7058 3610
rect 7092 3576 7144 3610
rect 7178 3576 7230 3610
rect 7264 3576 7316 3610
rect 7350 3576 7402 3610
rect 7436 3576 7448 3610
rect 6944 3570 7448 3576
rect 6944 3550 7118 3570
tri 7118 3550 7138 3570 nw
rect 6944 3323 7104 3550
tri 7104 3536 7118 3550 nw
tri 7457 3475 7476 3494 se
rect 7476 3475 7576 3700
tri 7442 3460 7457 3475 se
rect 7457 3460 7576 3475
rect 7132 3454 7576 3460
rect 7132 3420 7144 3454
rect 7178 3420 7222 3454
rect 7256 3420 7299 3454
rect 7333 3420 7376 3454
rect 7410 3420 7453 3454
rect 7487 3420 7530 3454
rect 7564 3420 7576 3454
rect 7132 3414 7576 3420
tri 7442 3399 7457 3414 ne
rect 7457 3399 7576 3414
tri 7457 3380 7476 3399 ne
tri 7104 3323 7119 3338 sw
rect 6944 3315 7119 3323
rect 6996 3298 7052 3315
rect 7104 3304 7119 3315
tri 7119 3304 7138 3323 sw
rect 7104 3298 7448 3304
rect 7006 3264 7052 3298
rect 7104 3264 7144 3298
rect 7178 3264 7230 3298
rect 7264 3264 7316 3298
rect 7350 3264 7402 3298
rect 7436 3264 7448 3298
rect 6996 3263 7052 3264
rect 7104 3263 7448 3264
rect 6944 3258 7448 3263
rect 7476 3272 7576 3399
rect 6944 3247 7127 3258
tri 7127 3247 7138 3258 nw
rect 6944 3244 7104 3247
rect 6996 3192 7052 3244
tri 7104 3224 7127 3247 nw
rect 6944 3172 7104 3192
rect 7476 3220 7524 3272
rect 7476 3208 7576 3220
rect 6996 3120 7052 3172
tri 7465 3171 7476 3182 se
rect 7476 3171 7524 3208
tri 7442 3148 7465 3171 se
rect 7465 3156 7524 3171
rect 7465 3148 7576 3156
rect 6944 3100 7104 3120
rect 7132 3142 7576 3148
rect 7132 3108 7144 3142
rect 7178 3108 7222 3142
rect 7256 3108 7299 3142
rect 7333 3108 7376 3142
rect 7410 3108 7453 3142
rect 7487 3108 7530 3142
rect 7564 3108 7576 3142
rect 7132 3102 7576 3108
rect 6996 3048 7052 3100
tri 7442 3096 7448 3102 ne
rect 7448 3096 7576 3102
tri 7448 3095 7449 3096 ne
rect 7449 3095 7576 3096
tri 7449 3068 7476 3095 ne
rect 6944 3028 7104 3048
rect 6996 2986 7052 3028
tri 7104 3023 7107 3026 sw
rect 7104 3019 7107 3023
tri 7107 3019 7111 3023 sw
rect 7104 2992 7111 3019
tri 7111 2992 7138 3019 sw
rect 7104 2986 7448 2992
rect 7006 2976 7052 2986
rect 7104 2976 7144 2986
rect 6944 2952 6972 2976
rect 7006 2952 7058 2976
rect 7092 2952 7144 2976
rect 7178 2952 7230 2986
rect 7264 2952 7316 2986
rect 7350 2952 7402 2986
rect 7436 2952 7448 2986
rect 6944 2946 7448 2952
rect 6944 2943 7135 2946
tri 7135 2943 7138 2946 nw
rect 6944 2680 7104 2943
tri 7104 2912 7135 2943 nw
tri 7473 2867 7476 2870 se
rect 7476 2867 7576 3095
tri 7442 2836 7473 2867 se
rect 7473 2836 7576 2867
rect 7132 2830 7576 2836
rect 7132 2796 7144 2830
rect 7178 2796 7227 2830
rect 7261 2796 7310 2830
rect 7344 2796 7392 2830
rect 7426 2796 7474 2830
rect 7508 2805 7576 2830
rect 7618 3741 7624 3749
rect 7658 3741 7667 3755
rect 7618 3700 7667 3741
rect 7618 3666 7624 3700
rect 7658 3666 7667 3700
rect 7618 3625 7667 3666
rect 7618 3591 7624 3625
rect 7658 3591 7667 3625
rect 7618 3550 7667 3591
rect 7618 3516 7624 3550
rect 7658 3516 7667 3550
rect 7618 3475 7667 3516
rect 7618 3441 7624 3475
rect 7658 3441 7667 3475
rect 7618 3399 7667 3441
rect 7618 3365 7624 3399
rect 7658 3365 7667 3399
rect 7618 3323 7667 3365
rect 7618 3289 7624 3323
rect 7658 3289 7667 3323
rect 7618 3247 7667 3289
rect 7618 3213 7624 3247
rect 7658 3213 7667 3247
rect 7618 3171 7667 3213
rect 7618 3137 7624 3171
rect 7658 3137 7667 3171
rect 7618 3095 7667 3137
rect 7618 3061 7624 3095
rect 7658 3061 7667 3095
rect 7618 3019 7667 3061
rect 7618 2985 7624 3019
rect 7658 2985 7667 3019
rect 7618 2943 7667 2985
rect 7618 2909 7624 2943
rect 7658 2909 7667 2943
rect 7618 2867 7667 2909
rect 7618 2833 7624 2867
rect 7658 2833 7667 2867
rect 7508 2804 7534 2805
tri 7534 2804 7535 2805 nw
rect 7508 2796 7525 2804
rect 7132 2795 7525 2796
tri 7525 2795 7534 2804 nw
rect 7132 2791 7521 2795
tri 7521 2791 7525 2795 nw
tri 7614 2791 7618 2795 se
rect 7618 2791 7667 2833
rect 7132 2790 7520 2791
tri 7520 2790 7521 2791 nw
tri 7613 2790 7614 2791 se
rect 7614 2790 7624 2791
tri 7585 2762 7613 2790 se
rect 7613 2762 7624 2790
tri 7578 2758 7582 2762 se
rect 7582 2758 7624 2762
tri 7577 2757 7578 2758 se
rect 7578 2757 7624 2758
rect 7658 2757 7667 2791
rect 7710 3865 7716 3899
rect 7750 3865 7756 3899
rect 7710 3826 7756 3865
rect 7710 3792 7716 3826
rect 7750 3792 7756 3826
rect 7710 3753 7756 3792
rect 7710 3719 7716 3753
rect 7750 3719 7756 3753
rect 7710 3680 7756 3719
rect 7710 3646 7716 3680
rect 7750 3646 7756 3680
rect 7710 3607 7756 3646
rect 7710 3573 7716 3607
rect 7750 3573 7756 3607
rect 7710 3534 7756 3573
rect 7784 3687 7875 4039
rect 7784 3635 7823 3687
rect 7784 3606 7875 3635
rect 7784 3554 7823 3606
rect 7784 3548 7875 3554
rect 7710 3500 7716 3534
rect 7750 3500 7756 3534
rect 7710 3461 7756 3500
rect 7710 3427 7716 3461
rect 7750 3427 7756 3461
rect 7710 3388 7756 3427
rect 7710 3354 7716 3388
rect 7750 3354 7756 3388
rect 7710 3315 7756 3354
rect 7710 3281 7716 3315
rect 7750 3281 7756 3315
rect 7710 3242 7756 3281
rect 7710 3208 7716 3242
rect 7750 3208 7756 3242
rect 7710 3169 7756 3208
rect 7710 3135 7716 3169
rect 7750 3135 7756 3169
rect 7710 3096 7756 3135
rect 7710 3062 7716 3096
rect 7750 3062 7756 3096
rect 7710 3023 7756 3062
rect 7710 2989 7716 3023
rect 7750 2989 7756 3023
rect 7710 2950 7756 2989
rect 7710 2916 7716 2950
rect 7750 2916 7756 2950
rect 7710 2877 7756 2916
rect 7710 2843 7716 2877
rect 7750 2843 7756 2877
rect 7710 2804 7756 2843
rect 7710 2770 7716 2804
rect 7750 2770 7756 2804
rect 7710 2758 7756 2770
rect 7903 2931 7955 8242
rect 7903 2867 7955 2879
tri 7534 2714 7577 2757 se
rect 7577 2714 7667 2757
tri 7104 2680 7138 2714 sw
tri 7531 2711 7534 2714 se
rect 7534 2711 7667 2714
tri 7524 2704 7531 2711 se
rect 7531 2704 7576 2711
rect 6944 2674 7448 2680
rect 6944 2640 6972 2674
rect 7006 2640 7058 2674
rect 7092 2640 7144 2674
rect 7178 2640 7230 2674
rect 7264 2640 7316 2674
rect 7350 2640 7402 2674
rect 7436 2640 7448 2674
rect 6944 2634 7448 2640
rect 6944 2626 7130 2634
tri 7130 2626 7138 2634 nw
rect 6944 2617 7121 2626
tri 7121 2617 7130 2626 nw
rect 6944 2484 7104 2617
tri 7104 2600 7121 2617 nw
tri 7509 2543 7524 2558 se
rect 7524 2543 7576 2704
tri 7576 2682 7605 2711 nw
tri 7874 2634 7903 2663 se
rect 7903 2634 7955 2815
rect 8208 2880 8260 8811
rect 8368 8562 8420 9417
tri 8738 9219 8772 9253 se
rect 8772 9219 8824 9659
rect 8696 9167 8702 9219
rect 8754 9167 8766 9219
rect 8818 9167 8824 9219
tri 8738 9151 8754 9167 ne
rect 8754 9151 8824 9167
tri 8754 9133 8772 9151 ne
rect 8368 8498 8420 8510
rect 8208 2816 8260 2828
rect 8208 2758 8260 2764
rect 8288 8280 8340 8286
rect 8288 8216 8340 8228
tri 7869 2629 7874 2634 se
rect 7874 2629 7955 2634
tri 7490 2524 7509 2543 se
rect 7509 2524 7576 2543
rect 7132 2518 7576 2524
rect 7132 2484 7144 2518
rect 7178 2484 7222 2518
rect 7256 2484 7299 2518
rect 7333 2484 7376 2518
rect 7410 2484 7453 2518
rect 7487 2484 7530 2518
rect 7564 2484 7576 2518
rect 7132 2478 7576 2484
rect 7619 2617 7955 2629
rect 8288 2748 8340 8164
rect 8288 2684 8340 2696
rect 8288 2626 8340 2632
rect 7619 2583 7625 2617
rect 7659 2583 7955 2617
rect 7619 2577 7955 2583
rect 7619 2523 7665 2577
tri 7665 2543 7699 2577 nw
rect 7619 2489 7625 2523
rect 7659 2489 7665 2523
rect 7619 2477 7665 2489
rect 8368 2503 8420 8446
rect 8528 8642 8580 8648
rect 8528 8578 8580 8590
rect 8448 8406 8500 8412
rect 8448 8342 8500 8354
rect 8448 2716 8500 8290
rect 8448 2652 8500 2664
rect 8448 2594 8500 2600
tri 8420 2503 8454 2537 sw
tri 6823 2350 6844 2371 se
rect 6844 2350 6902 2371
rect 8368 2451 8374 2503
rect 8426 2451 8438 2503
rect 8490 2451 8496 2503
rect 4238 2343 4271 2350
tri 4271 2343 4278 2350 sw
tri 6816 2343 6823 2350 se
rect 6823 2343 6902 2350
rect 4238 2325 5462 2343
rect 3799 2245 3805 2297
rect 3857 2245 3869 2297
rect 3921 2291 4069 2297
tri 4069 2291 4075 2297 sw
rect 4116 2291 5462 2325
rect 6774 2291 6780 2343
rect 6832 2291 6844 2343
rect 6896 2291 6902 2343
tri 7960 2316 7994 2350 se
rect 7044 2309 7996 2316
rect 3921 2275 4075 2291
tri 4075 2275 4091 2291 sw
tri 5376 2275 5392 2291 ne
rect 5392 2275 5462 2291
rect 3921 2257 4091 2275
tri 4091 2257 4109 2275 sw
tri 5392 2257 5410 2275 ne
rect 3921 2245 4109 2257
tri 4047 2241 4051 2245 ne
rect 4051 2241 4109 2245
tri 4109 2241 4125 2257 sw
tri 4051 2231 4061 2241 ne
rect 4061 2231 5264 2241
tri 5264 2231 5274 2241 sw
tri 4061 2223 4069 2231 ne
rect 4069 2223 5274 2231
tri 4069 2217 4075 2223 ne
rect 4075 2217 5274 2223
rect 2087 2165 2093 2217
rect 2145 2165 2157 2217
rect 2209 2165 2215 2217
rect 3771 2165 3777 2217
rect 3829 2165 3841 2217
rect 3893 2171 3899 2217
tri 4075 2197 4095 2217 ne
rect 4095 2197 5274 2217
tri 5274 2197 5308 2231 sw
tri 4095 2189 4103 2197 ne
rect 4103 2189 5308 2197
tri 5308 2189 5316 2197 sw
tri 5242 2184 5247 2189 ne
rect 5247 2184 5316 2189
tri 5316 2184 5321 2189 sw
tri 3899 2171 3912 2184 sw
tri 5247 2171 5260 2184 ne
rect 5260 2171 5321 2184
tri 5321 2171 5334 2184 sw
rect 3893 2165 3912 2171
tri 3912 2165 3918 2171 sw
tri 5260 2165 5266 2171 ne
rect 5266 2165 5334 2171
tri 5334 2165 5340 2171 sw
tri 2129 2131 2163 2165 ne
tri 1865 2048 1899 2082 sw
tri 2129 2048 2163 2082 se
rect 2163 2048 2215 2165
tri 3813 2153 3825 2165 ne
rect 3825 2153 3918 2165
tri 3918 2153 3930 2165 sw
tri 5266 2157 5274 2165 ne
rect 5274 2157 5340 2165
tri 5340 2157 5348 2165 sw
tri 5274 2153 5278 2157 ne
rect 5278 2153 5348 2157
tri 3825 2131 3847 2153 ne
rect 3847 2150 3930 2153
tri 3930 2150 3933 2153 sw
tri 5278 2150 5281 2153 ne
rect 5281 2150 5348 2153
rect 3847 2098 5241 2150
tri 5281 2135 5296 2150 ne
tri 5077 2085 5090 2098 ne
rect 5090 2085 5241 2098
tri 5090 2082 5093 2085 ne
rect 5093 2082 5241 2085
tri 5093 2075 5100 2082 ne
rect 5100 2075 5241 2082
tri 5100 2064 5111 2075 ne
rect 1813 1996 2215 2048
tri 2129 1962 2163 1996 ne
tri 1785 1866 1819 1900 sw
rect 1733 1814 1961 1866
tri 1875 1780 1909 1814 ne
rect 1652 58 1704 70
rect 1652 0 1704 6
rect 1909 122 1961 1814
rect 1909 58 1961 70
rect 1909 0 1961 6
rect 2163 122 2215 1996
rect 3195 1984 3201 2036
rect 3253 1984 3267 2036
rect 3319 1984 3325 2036
rect 3911 1984 3917 2036
rect 3969 1984 3994 2036
rect 4046 1984 4052 2036
rect 5111 1986 5241 2075
tri 5293 1963 5296 1966 se
rect 5296 1963 5348 2150
tri 5292 1962 5293 1963 se
rect 5293 1962 5348 1963
tri 5278 1948 5292 1962 se
rect 5292 1948 5348 1962
rect 3708 1942 3760 1948
tri 2994 1885 2995 1886 se
tri 2975 1866 2994 1885 se
rect 2994 1866 2995 1885
tri 2961 1852 2975 1866 se
rect 2975 1852 2995 1866
tri 3041 1885 3042 1886 sw
rect 3041 1852 3042 1885
tri 3042 1852 3075 1885 sw
rect 3708 1858 3760 1890
rect 2955 1800 2961 1852
rect 3013 1800 3025 1852
rect 3077 1800 3083 1852
rect 3708 1800 3760 1806
rect 4908 1942 4960 1948
tri 5262 1932 5278 1948 se
rect 5278 1932 5348 1948
rect 4908 1858 4960 1890
rect 5296 1880 5348 1932
rect 5410 1918 5462 2275
rect 7044 2275 7076 2309
rect 7110 2275 7155 2309
rect 7189 2275 7234 2309
rect 7268 2275 7313 2309
rect 7347 2275 7392 2309
rect 7426 2275 7470 2309
rect 7504 2275 7548 2309
rect 7582 2275 7626 2309
rect 7660 2275 7704 2309
rect 7738 2275 7782 2309
rect 7816 2275 7860 2309
rect 7894 2275 7996 2309
rect 7044 2231 7996 2275
rect 7044 2197 7076 2231
rect 7110 2197 7155 2231
rect 7189 2197 7234 2231
rect 7268 2197 7313 2231
rect 7347 2197 7392 2231
rect 7426 2197 7470 2231
rect 7504 2197 7548 2231
rect 7582 2197 7626 2231
rect 7660 2197 7704 2231
rect 7738 2197 7782 2231
rect 7816 2197 7860 2231
rect 7894 2197 7996 2231
rect 7044 2153 7996 2197
rect 7044 2119 7076 2153
rect 7110 2119 7155 2153
rect 7189 2119 7234 2153
rect 7268 2119 7313 2153
rect 7347 2119 7392 2153
rect 7426 2119 7470 2153
rect 7504 2119 7548 2153
rect 7582 2119 7626 2153
rect 7660 2119 7704 2153
rect 7738 2119 7782 2153
rect 7816 2119 7860 2153
rect 7894 2119 7996 2153
rect 8368 2183 8420 2451
tri 8420 2417 8454 2451 nw
tri 8420 2183 8454 2217 sw
rect 8368 2131 8374 2183
rect 8426 2131 8438 2183
rect 8490 2131 8496 2183
rect 7044 2075 7996 2119
rect 7044 2041 7076 2075
rect 7110 2041 7155 2075
rect 7189 2041 7234 2075
rect 7268 2041 7313 2075
rect 7347 2041 7392 2075
rect 7426 2041 7470 2075
rect 7504 2041 7548 2075
rect 7582 2041 7626 2075
rect 7660 2041 7704 2075
rect 7738 2041 7782 2075
rect 7816 2041 7860 2075
rect 7894 2041 7996 2075
rect 5827 1980 5833 2032
rect 5885 1980 5910 2032
rect 5962 1980 5968 2032
rect 6543 1984 6549 2036
rect 6601 1984 6626 2036
rect 6678 1984 6684 2036
rect 7044 1997 7996 2041
tri 8494 2036 8528 2070 se
rect 8528 2036 8580 8526
rect 7044 1963 7076 1997
rect 7110 1963 7155 1997
rect 7189 1963 7234 1997
rect 7268 1963 7313 1997
rect 7347 1963 7392 1997
rect 7426 1963 7470 1997
rect 7504 1963 7548 1997
rect 7582 1963 7626 1997
rect 7660 1963 7704 1997
rect 7738 1963 7782 1997
rect 7816 1963 7860 1997
rect 7894 1963 7996 1997
rect 8452 1984 8458 2036
rect 8510 1984 8522 2036
rect 8574 1984 8580 2036
rect 8608 8221 8660 8227
rect 8608 8157 8660 8169
rect 4908 1800 4960 1806
rect 5410 1854 5462 1866
rect 5410 1796 5462 1802
rect 5621 1942 5673 1948
rect 5621 1858 5673 1890
rect 5621 1800 5673 1806
rect 6340 1942 6392 1948
rect 6340 1858 6392 1890
rect 6340 1800 6392 1806
rect 7044 1919 7996 1963
tri 8592 1950 8608 1966 se
rect 8608 1950 8660 8105
tri 8574 1932 8592 1950 se
rect 8592 1932 8660 1950
rect 7044 1885 7076 1919
rect 7110 1885 7155 1919
rect 7189 1885 7234 1919
rect 7268 1885 7313 1919
rect 7347 1885 7392 1919
rect 7426 1885 7470 1919
rect 7504 1885 7548 1919
rect 7582 1885 7626 1919
rect 7660 1885 7704 1919
rect 7738 1885 7782 1919
rect 7816 1885 7860 1919
rect 7894 1885 7996 1919
rect 7044 1841 7996 1885
rect 8532 1880 8538 1932
rect 8590 1880 8602 1932
rect 8654 1880 8660 1932
rect 8688 8120 8740 8126
rect 8688 8056 8740 8068
rect 7044 1807 7076 1841
rect 7110 1807 7155 1841
rect 7189 1807 7234 1841
rect 7268 1807 7313 1841
rect 7347 1807 7392 1841
rect 7426 1807 7470 1841
rect 7504 1807 7548 1841
rect 7582 1807 7626 1841
rect 7660 1807 7704 1841
rect 7738 1807 7782 1841
rect 7816 1807 7860 1841
rect 7894 1807 7996 1841
rect 7044 1800 7996 1807
rect 8688 1846 8740 8004
rect 8772 4524 8824 9151
rect 8772 4460 8824 4472
rect 8772 3101 8824 4408
rect 8772 3037 8824 3049
rect 8772 2979 8824 2985
rect 8852 9149 8904 9155
rect 8852 9085 8904 9097
tri 8818 2932 8852 2966 se
rect 8852 2932 8904 9033
rect 8932 5010 8984 10193
rect 8932 4946 8984 4958
rect 8932 4888 8984 4894
rect 9012 9956 9064 9962
rect 9012 9892 9064 9904
rect 8805 2880 8904 2932
rect 8805 2493 8857 2880
tri 8857 2846 8891 2880 nw
rect 8805 2429 8857 2441
rect 8805 2371 8857 2377
tri 9001 2634 9012 2645 se
rect 9012 2634 9064 9840
rect 9001 2582 9064 2634
tri 7960 1796 7964 1800 ne
rect 7964 1796 7994 1800
tri 7964 1766 7994 1796 ne
rect 8688 1782 8740 1794
rect 3469 1619 4397 1746
tri 4397 1619 4524 1746 sw
rect 4747 1694 6479 1746
rect 6531 1694 6580 1746
rect 6632 1694 6681 1746
rect 6733 1694 6782 1746
rect 6834 1694 6882 1746
rect 6934 1694 6982 1746
rect 7034 1694 7082 1746
rect 7134 1694 7182 1746
rect 7234 1694 7282 1746
rect 7334 1694 7382 1746
rect 7434 1694 7482 1746
rect 7534 1694 7582 1746
rect 7634 1694 7682 1746
rect 7734 1694 7782 1746
rect 7834 1694 7840 1746
rect 8688 1724 8740 1730
rect 8788 1984 8794 2036
rect 8846 1984 8858 2036
rect 8910 1984 8916 2036
rect 4747 1672 7840 1694
rect 4747 1620 6479 1672
rect 6531 1620 6580 1672
rect 6632 1620 6681 1672
rect 6733 1620 6782 1672
rect 6834 1620 6882 1672
rect 6934 1620 6982 1672
rect 7034 1620 7082 1672
rect 7134 1620 7182 1672
rect 7234 1620 7282 1672
rect 7334 1620 7382 1672
rect 7434 1620 7482 1672
rect 7534 1620 7582 1672
rect 7634 1620 7682 1672
rect 7734 1620 7782 1672
rect 7834 1620 7840 1672
rect 4747 1619 7840 1620
rect 3469 1591 4524 1619
tri 4524 1591 4552 1619 sw
rect 3469 1574 4552 1591
tri 4552 1574 4569 1591 sw
tri 7977 1574 7994 1591 se
tri 4327 1557 4344 1574 ne
rect 4344 1557 4569 1574
tri 4569 1557 4586 1574 sw
tri 7960 1557 7977 1574 se
rect 7977 1557 7994 1574
tri 4344 1545 4356 1557 ne
rect 4356 1545 4586 1557
tri 4586 1545 4598 1557 sw
rect 7038 1545 7994 1557
tri 4356 1520 4381 1545 ne
rect 4381 1520 4598 1545
rect 2955 1468 2961 1520
rect 3013 1468 3025 1520
rect 3077 1468 3083 1520
tri 4381 1518 4383 1520 ne
rect 4383 1518 4598 1520
rect 3521 1516 4126 1518
tri 2961 1444 2985 1468 ne
rect 2985 1444 2995 1468
tri 2985 1438 2991 1444 ne
rect 2991 1438 2995 1444
tri 2991 1434 2995 1438 ne
rect 3041 1438 3045 1468
tri 3045 1438 3075 1468 nw
rect 3521 1464 3527 1516
rect 3579 1464 3595 1516
rect 3647 1464 3663 1516
rect 3715 1464 3731 1516
rect 3783 1464 3799 1516
rect 3851 1464 3867 1516
rect 3919 1464 3934 1516
rect 3986 1464 4001 1516
rect 4053 1464 4068 1516
rect 4120 1464 4126 1516
tri 4383 1511 4390 1518 ne
rect 4390 1511 4598 1518
tri 4598 1511 4632 1545 sw
rect 7038 1511 7049 1545
rect 7083 1511 7121 1545
rect 7155 1511 7193 1545
rect 7227 1511 7265 1545
rect 7299 1511 7337 1545
rect 7371 1511 7409 1545
rect 7443 1511 7481 1545
rect 7515 1511 7553 1545
rect 7587 1511 7625 1545
rect 7659 1511 7697 1545
rect 7731 1511 7769 1545
rect 7803 1511 7841 1545
rect 7875 1511 7994 1545
tri 4390 1472 4429 1511 ne
rect 4429 1472 4632 1511
tri 4632 1472 4671 1511 sw
rect 7038 1472 7994 1511
tri 4429 1468 4433 1472 ne
rect 4433 1468 4671 1472
rect 3521 1452 4126 1464
tri 3041 1434 3045 1438 nw
rect 3521 1400 3527 1452
rect 3579 1400 3595 1452
rect 3647 1400 3663 1452
rect 3715 1400 3731 1452
rect 3783 1400 3799 1452
rect 3851 1400 3867 1452
rect 3919 1400 3934 1452
rect 3986 1400 4001 1452
rect 4053 1400 4068 1452
rect 4120 1400 4126 1452
tri 4433 1438 4463 1468 ne
rect 4463 1438 4671 1468
tri 4671 1438 4705 1472 sw
rect 7038 1438 7049 1472
rect 7083 1438 7121 1472
rect 7155 1438 7193 1472
rect 7227 1438 7265 1472
rect 7299 1438 7337 1472
rect 7371 1438 7409 1472
rect 7443 1438 7481 1472
rect 7515 1438 7553 1472
rect 7587 1438 7625 1472
rect 7659 1438 7697 1472
rect 7731 1438 7769 1472
rect 7803 1438 7841 1472
rect 7875 1438 7994 1472
tri 4463 1434 4467 1438 ne
rect 4467 1434 4705 1438
rect 3521 1388 4126 1400
tri 4467 1399 4502 1434 ne
rect 4502 1399 4705 1434
tri 4705 1399 4744 1438 sw
rect 7038 1399 7994 1438
rect 3195 1285 3201 1337
rect 3253 1285 3267 1337
rect 3319 1285 3325 1337
rect 3521 1336 3527 1388
rect 3579 1336 3595 1388
rect 3647 1336 3663 1388
rect 3715 1336 3731 1388
rect 3783 1336 3799 1388
rect 3851 1336 3867 1388
rect 3919 1336 3934 1388
rect 3986 1336 4001 1388
rect 4053 1336 4068 1388
rect 4120 1336 4126 1388
tri 4502 1365 4536 1399 ne
rect 4536 1365 4744 1399
tri 4744 1365 4778 1399 sw
rect 7038 1365 7049 1399
rect 7083 1365 7121 1399
rect 7155 1365 7193 1399
rect 7227 1365 7265 1399
rect 7299 1365 7337 1399
rect 7371 1365 7409 1399
rect 7443 1365 7481 1399
rect 7515 1365 7553 1399
rect 7587 1365 7625 1399
rect 7659 1365 7697 1399
rect 7731 1365 7769 1399
rect 7803 1365 7841 1399
rect 7875 1365 7994 1399
tri 4536 1337 4564 1365 ne
rect 4564 1337 4778 1365
rect 3521 1324 4126 1336
tri 4564 1332 4569 1337 ne
rect 4569 1332 4778 1337
tri 4778 1332 4811 1365 sw
tri 4569 1326 4575 1332 ne
rect 4575 1326 4811 1332
tri 4811 1326 4817 1332 sw
rect 7038 1326 7994 1365
rect 3521 1272 3527 1324
rect 3579 1272 3595 1324
rect 3647 1272 3663 1324
rect 3715 1272 3731 1324
rect 3783 1272 3799 1324
rect 3851 1272 3867 1324
rect 3919 1272 3934 1324
rect 3986 1272 4001 1324
rect 4053 1272 4068 1324
rect 4120 1272 4126 1324
tri 4575 1292 4609 1326 ne
rect 4609 1292 4817 1326
tri 4817 1292 4851 1326 sw
rect 7038 1292 7049 1326
rect 7083 1292 7121 1326
rect 7155 1292 7193 1326
rect 7227 1292 7265 1326
rect 7299 1292 7337 1326
rect 7371 1292 7409 1326
rect 7443 1292 7481 1326
rect 7515 1292 7553 1326
rect 7587 1292 7625 1326
rect 7659 1292 7697 1326
rect 7731 1292 7769 1326
rect 7803 1292 7841 1326
rect 7875 1292 7994 1326
tri 4609 1285 4616 1292 ne
rect 4616 1285 4851 1292
rect 3521 1260 4126 1272
rect 3521 1208 3527 1260
rect 3579 1208 3595 1260
rect 3647 1208 3663 1260
rect 3715 1208 3731 1260
rect 3783 1208 3799 1260
rect 3851 1208 3867 1260
rect 3919 1208 3934 1260
rect 3986 1208 4001 1260
rect 4053 1208 4068 1260
rect 4120 1208 4126 1260
tri 4616 1253 4648 1285 ne
rect 4648 1253 4851 1285
tri 4851 1253 4890 1292 sw
rect 7038 1253 7994 1292
tri 4648 1219 4682 1253 ne
rect 4682 1219 4890 1253
tri 4890 1219 4924 1253 sw
rect 7038 1219 7049 1253
rect 7083 1219 7121 1253
rect 7155 1219 7193 1253
rect 7227 1219 7265 1253
rect 7299 1219 7337 1253
rect 7371 1219 7409 1253
rect 7443 1219 7481 1253
rect 7515 1219 7553 1253
rect 7587 1219 7625 1253
rect 7659 1219 7697 1253
rect 7731 1219 7769 1253
rect 7803 1219 7841 1253
rect 7875 1219 7994 1253
tri 3506 929 3521 944 se
rect 3521 929 4126 1208
tri 4682 1180 4721 1219 ne
rect 4721 1208 4924 1219
tri 4924 1208 4935 1219 sw
rect 4721 1180 4935 1208
tri 4935 1180 4963 1208 sw
rect 7038 1180 7994 1219
tri 4721 1146 4755 1180 ne
rect 4755 1146 4963 1180
tri 4963 1146 4997 1180 sw
rect 7038 1146 7049 1180
rect 7083 1146 7121 1180
rect 7155 1146 7193 1180
rect 7227 1146 7265 1180
rect 7299 1146 7337 1180
rect 7371 1146 7409 1180
rect 7443 1146 7481 1180
rect 7515 1146 7553 1180
rect 7587 1146 7625 1180
rect 7659 1146 7697 1180
rect 7731 1146 7769 1180
rect 7803 1146 7841 1180
rect 7875 1146 7994 1180
tri 4755 1107 4794 1146 ne
rect 4794 1107 4997 1146
tri 4997 1107 5036 1146 sw
rect 7038 1107 7994 1146
tri 4794 1090 4811 1107 ne
rect 4811 1090 5036 1107
tri 5036 1090 5053 1107 sw
tri 4811 1078 4823 1090 ne
rect 4823 1078 5053 1090
tri 5053 1078 5065 1090 sw
tri 4823 1073 4828 1078 ne
rect 4828 1073 6623 1078
tri 4828 1034 4867 1073 ne
rect 4867 1048 6623 1073
rect 4867 1034 5829 1048
tri 4867 1000 4901 1034 ne
rect 4901 1000 5829 1034
tri 4901 966 4935 1000 ne
rect 4935 996 5829 1000
rect 5881 996 5896 1048
rect 5948 996 5963 1048
rect 6015 996 6030 1048
rect 6082 996 6097 1048
rect 6149 996 6164 1048
rect 6216 996 6231 1048
rect 6283 996 6298 1048
rect 6350 996 6365 1048
rect 6417 996 6432 1048
rect 6484 996 6499 1048
rect 6551 996 6565 1048
rect 6617 996 6623 1048
rect 4935 966 6623 996
rect 7038 1073 7049 1107
rect 7083 1073 7121 1107
rect 7155 1073 7193 1107
rect 7227 1073 7265 1107
rect 7299 1073 7337 1107
rect 7371 1073 7409 1107
rect 7443 1073 7481 1107
rect 7515 1073 7553 1107
rect 7587 1073 7625 1107
rect 7659 1073 7697 1107
rect 7731 1073 7769 1107
rect 7803 1073 7841 1107
rect 7875 1073 7994 1107
rect 7038 1034 7994 1073
rect 7038 1000 7049 1034
rect 7083 1000 7121 1034
rect 7155 1000 7193 1034
rect 7227 1000 7265 1034
rect 7299 1000 7337 1034
rect 7371 1000 7409 1034
rect 7443 1000 7481 1034
rect 7515 1000 7553 1034
rect 7587 1000 7625 1034
rect 7659 1000 7697 1034
rect 7731 1000 7769 1034
rect 7803 1000 7841 1034
rect 7875 1000 7994 1034
rect 7038 961 7994 1000
tri 4126 929 4141 944 sw
tri 3504 927 3506 929 se
rect 3506 927 4141 929
tri 4141 927 4143 929 sw
rect 7038 927 7049 961
rect 7083 927 7121 961
rect 7155 927 7193 961
rect 7227 927 7265 961
rect 7299 927 7337 961
rect 7371 927 7409 961
rect 7443 927 7481 961
rect 7515 927 7553 961
rect 7587 927 7625 961
rect 7659 927 7697 961
rect 7731 927 7769 961
rect 7803 927 7841 961
rect 7875 927 7994 961
tri 3487 910 3504 927 se
rect 3504 910 4143 927
tri 4143 910 4160 927 sw
rect 7038 888 7994 927
rect 7038 854 7049 888
rect 7083 854 7121 888
rect 7155 854 7193 888
rect 7227 854 7265 888
rect 7299 854 7337 888
rect 7371 854 7409 888
rect 7443 854 7481 888
rect 7515 854 7553 888
rect 7587 854 7625 888
rect 7659 854 7697 888
rect 7731 854 7769 888
rect 7803 854 7841 888
rect 7875 854 7994 888
rect 8388 1064 8440 1095
rect 8388 1000 8440 1012
rect 7038 814 7994 854
tri 8354 844 8388 878 se
rect 8388 844 8440 948
rect 7038 780 7049 814
rect 7083 780 7121 814
rect 7155 780 7193 814
rect 7227 780 7265 814
rect 7299 780 7337 814
rect 7371 780 7409 814
rect 7443 780 7481 814
rect 7515 780 7553 814
rect 7587 780 7625 814
rect 7659 780 7697 814
rect 7731 780 7769 814
rect 7803 780 7841 814
rect 7875 780 7994 814
rect 7038 740 7994 780
tri 5009 711 5012 714 se
rect 5012 711 5018 714
tri 5006 708 5009 711 se
rect 5009 708 5018 711
rect 3604 656 3610 708
rect 3662 656 3674 708
rect 3726 656 3732 708
rect 4264 701 4316 707
tri 3732 656 3738 662 nw
rect 4264 637 4316 649
tri 3265 558 3269 562 se
tri 3263 556 3265 558 se
rect 3265 556 3269 558
tri 3235 528 3263 556 se
rect 3263 528 3269 556
tri 3315 558 3319 562 sw
rect 3315 528 3319 558
tri 3319 528 3349 558 sw
rect 3706 556 3712 608
rect 3764 556 3776 608
rect 3828 556 3834 608
tri 2955 476 2957 478 se
tri 2923 444 2955 476 se
rect 2955 444 2957 476
tri 3003 444 3037 478 sw
rect 3226 476 3232 528
rect 3284 476 3296 528
rect 3348 476 3354 528
tri 3235 444 3267 476 ne
rect 3267 444 3269 476
rect 2917 392 2923 444
rect 2975 392 2987 444
rect 3039 392 3045 444
tri 3267 442 3269 444 ne
rect 3315 444 3317 476
tri 3317 444 3349 476 nw
tri 3315 442 3317 444 nw
rect 4264 395 4316 585
rect 4576 701 4628 707
rect 5012 662 5018 708
rect 5070 662 5082 714
rect 5134 662 5140 714
tri 5140 708 5146 714 sw
tri 5973 708 5976 711 se
tri 5973 659 5976 662 ne
rect 5976 659 5982 711
rect 6034 659 6046 711
rect 6098 659 6104 711
rect 7038 706 7049 740
rect 7083 706 7121 740
rect 7155 706 7193 740
rect 7227 706 7265 740
rect 7299 706 7337 740
rect 7371 706 7409 740
rect 7443 706 7481 740
rect 7515 706 7553 740
rect 7587 706 7625 740
rect 7659 706 7697 740
rect 7731 706 7769 740
rect 7803 706 7841 740
rect 7875 706 7994 740
rect 7038 666 7994 706
rect 4576 626 4628 649
rect 7038 632 7049 666
rect 7083 632 7121 666
rect 7155 632 7193 666
rect 7227 632 7265 666
rect 7299 632 7337 666
rect 7371 632 7409 666
rect 7443 632 7481 666
rect 7515 632 7553 666
rect 7587 632 7625 666
rect 7659 632 7697 666
rect 7731 632 7769 666
rect 7803 632 7841 666
rect 7875 632 7994 666
rect 4576 395 4628 574
rect 5016 559 5022 611
rect 5074 559 5086 611
rect 5138 559 5144 611
rect 5874 556 5880 608
rect 5932 556 5944 608
rect 5996 556 6002 608
rect 7038 592 7994 632
tri 6389 558 6393 562 se
tri 6387 556 6389 558 se
rect 6389 556 6393 558
tri 6359 528 6387 556 se
rect 6387 528 6393 556
tri 6439 558 6443 562 sw
rect 7038 558 7049 592
rect 7083 558 7121 592
rect 7155 558 7193 592
rect 7227 558 7265 592
rect 7299 558 7337 592
rect 7371 558 7409 592
rect 7443 558 7481 592
rect 7515 558 7553 592
rect 7587 558 7625 592
rect 7659 558 7697 592
rect 7731 558 7769 592
rect 7803 558 7841 592
rect 7875 558 7994 592
rect 6439 528 6443 558
tri 6443 528 6473 558 sw
rect 6354 476 6360 528
rect 6412 476 6424 528
rect 6476 476 6482 528
rect 7038 518 7994 558
rect 7038 484 7049 518
rect 7083 484 7121 518
rect 7155 484 7193 518
rect 7227 484 7265 518
rect 7299 484 7337 518
rect 7371 484 7409 518
rect 7443 484 7481 518
rect 7515 484 7553 518
rect 7587 484 7625 518
rect 7659 484 7697 518
rect 7731 484 7769 518
rect 7803 484 7841 518
rect 7875 484 7994 518
tri 6703 476 6705 478 se
tri 6359 444 6391 476 ne
rect 6391 444 6393 476
tri 6391 442 6393 444 ne
rect 6439 444 6441 476
tri 6441 444 6473 476 nw
tri 6671 444 6703 476 se
rect 6703 444 6705 476
tri 6751 444 6785 478 sw
rect 7038 444 7994 484
tri 6439 442 6441 444 nw
rect 6663 392 6669 444
rect 6721 392 6733 444
rect 6785 392 6791 444
rect 7038 410 7049 444
rect 7083 410 7121 444
rect 7155 410 7193 444
rect 7227 410 7265 444
rect 7299 410 7337 444
rect 7371 410 7409 444
rect 7443 410 7481 444
rect 7515 410 7553 444
rect 7587 410 7625 444
rect 7659 410 7697 444
rect 7731 410 7769 444
rect 7803 410 7841 444
rect 7875 410 7994 444
rect 7038 370 7994 410
rect 2981 301 2987 353
rect 3039 301 3053 353
rect 3105 301 3111 353
rect 4291 304 4297 356
rect 4349 304 4363 356
rect 4415 304 4421 356
rect 6597 301 6603 353
rect 6655 301 6669 353
rect 6721 301 6727 353
rect 7038 336 7049 370
rect 7083 336 7121 370
rect 7155 336 7193 370
rect 7227 336 7265 370
rect 7299 336 7337 370
rect 7371 336 7409 370
rect 7443 336 7481 370
rect 7515 336 7553 370
rect 7587 336 7625 370
rect 7659 336 7697 370
rect 7731 336 7769 370
rect 7803 336 7841 370
rect 7875 336 7994 370
rect 7038 296 7994 336
rect 7038 262 7049 296
rect 7083 262 7121 296
rect 7155 262 7193 296
rect 7227 262 7265 296
rect 7299 262 7337 296
rect 7371 262 7409 296
rect 7443 262 7481 296
rect 7515 262 7553 296
rect 7587 262 7625 296
rect 7659 262 7697 296
rect 7731 262 7769 296
rect 7803 262 7841 296
rect 7875 262 7994 296
rect 7038 222 7994 262
rect 7038 188 7049 222
rect 7083 188 7121 222
rect 7155 188 7193 222
rect 7227 188 7265 222
rect 7299 188 7337 222
rect 7371 188 7409 222
rect 7443 188 7481 222
rect 7515 188 7553 222
rect 7587 188 7625 222
rect 7659 188 7697 222
rect 7731 188 7769 222
rect 7803 188 7841 222
rect 7875 188 7994 222
rect 2163 58 2215 70
rect 2163 0 2215 6
rect 2483 158 2561 164
rect 2483 106 2496 158
rect 2548 106 2561 158
rect 7038 148 7994 188
rect 2483 58 2561 106
rect 2483 6 2496 58
rect 2548 6 2561 58
rect 2483 0 2561 6
rect 6843 122 6895 128
rect 6843 58 6895 70
rect 7038 114 7049 148
rect 7083 114 7121 148
rect 7155 114 7193 148
rect 7227 114 7265 148
rect 7299 114 7337 148
rect 7371 114 7409 148
rect 7443 114 7481 148
rect 7515 114 7553 148
rect 7587 114 7625 148
rect 7659 114 7697 148
rect 7731 114 7769 148
rect 7803 114 7841 148
rect 7875 114 7994 148
rect 7038 74 7994 114
rect 7038 40 7049 74
rect 7083 40 7121 74
rect 7155 40 7193 74
rect 7227 40 7265 74
rect 7299 40 7337 74
rect 7371 40 7409 74
rect 7443 40 7481 74
rect 7515 40 7553 74
rect 7587 40 7625 74
rect 7659 40 7697 74
rect 7731 40 7769 74
rect 7803 40 7841 74
rect 7875 50 7994 74
rect 8176 792 8440 844
rect 8788 876 8840 1984
tri 8840 1950 8874 1984 nw
tri 8936 1788 9001 1853 se
rect 9001 1831 9053 2582
tri 9053 2571 9064 2582 nw
rect 9092 9632 9144 9642
rect 9092 9568 9144 9580
rect 9092 2333 9144 9516
rect 9092 2269 9144 2281
rect 9092 2211 9144 2217
rect 9172 9358 9224 9364
rect 9172 9294 9224 9306
rect 9001 1788 9010 1831
tri 9010 1788 9053 1831 nw
tri 8902 1426 8936 1460 se
rect 8936 1426 8996 1788
tri 8996 1774 9010 1788 nw
tri 9171 1619 9172 1620 se
rect 9172 1619 9224 9242
tri 9143 1591 9171 1619 se
rect 9171 1591 9224 1619
tri 9138 1586 9143 1591 se
rect 9143 1586 9224 1591
rect 9044 1534 9050 1586
rect 9102 1534 9114 1586
rect 9166 1534 9224 1586
tri 9138 1500 9172 1534 ne
rect 8868 1374 8874 1426
rect 8926 1374 8938 1426
rect 8990 1374 8996 1426
rect 9172 1080 9224 1534
rect 9172 1016 9224 1028
rect 9172 958 9224 964
tri 8840 876 8874 910 sw
rect 8788 824 8794 876
rect 8846 824 8858 876
rect 8910 824 8916 876
rect 8176 122 8228 792
tri 8228 758 8262 792 nw
rect 9252 444 9304 11866
rect 9332 781 9384 12025
rect 9332 717 9384 729
rect 9332 659 9384 665
rect 9412 678 9464 12321
rect 9572 12081 9624 14604
rect 9890 14466 9942 14472
rect 9890 14402 9942 14414
tri 9792 14261 9812 14281 sw
tri 9732 14247 9746 14261 se
rect 9792 14247 9812 14261
tri 9812 14247 9826 14261 sw
rect 9732 14241 9862 14247
rect 9784 14189 9808 14241
rect 9860 14189 9862 14241
rect 9732 14151 9862 14189
rect 9784 14099 9808 14151
rect 9860 14099 9862 14151
rect 9732 14061 9862 14099
rect 9784 14009 9808 14061
rect 9860 14009 9862 14061
rect 9732 14003 9862 14009
tri 9732 13989 9746 14003 ne
rect 9792 13989 9812 14003
tri 9812 13989 9826 14003 nw
tri 9792 13969 9812 13989 nw
tri 9792 12553 9812 12573 sw
tri 9732 12539 9746 12553 se
rect 9792 12539 9812 12553
tri 9812 12539 9826 12553 sw
rect 9732 12512 9862 12539
rect 9732 12460 9738 12512
rect 9790 12460 9804 12512
rect 9856 12460 9862 12512
rect 9732 12433 9862 12460
tri 9732 12419 9746 12433 ne
rect 9792 12419 9812 12433
tri 9812 12419 9826 12433 nw
tri 9792 12399 9812 12419 nw
rect 9890 12366 9942 14350
rect 10710 14255 10828 14261
rect 10762 14203 10776 14255
rect 10710 14158 10828 14203
rect 10762 14106 10776 14158
rect 10710 14061 10828 14106
rect 10762 14009 10776 14061
rect 10710 14003 10828 14009
rect 9890 12302 9942 12314
rect 9572 12017 9624 12029
rect 9572 11959 9624 11965
rect 9652 12262 9704 12268
rect 9890 12244 9942 12250
rect 9652 12198 9704 12210
rect 9572 11588 9624 11594
rect 9572 11524 9624 11536
rect 9492 9876 9544 9882
rect 9492 9812 9544 9824
rect 9492 1576 9544 9760
rect 9492 1512 9544 1524
rect 9492 1454 9544 1460
tri 9538 1186 9572 1220 se
rect 9572 1186 9624 11472
rect 9496 1134 9502 1186
rect 9554 1134 9566 1186
rect 9618 1134 9624 1186
rect 9652 1416 9704 12146
rect 9652 1352 9704 1364
rect 9572 1080 9624 1086
rect 9572 1016 9624 1028
rect 9412 614 9464 626
rect 9412 556 9464 562
rect 9492 946 9544 952
rect 9492 882 9544 894
tri 9304 444 9338 478 sw
rect 9252 392 9258 444
rect 9310 392 9322 444
rect 9374 392 9380 444
tri 9458 352 9492 386 se
rect 9492 352 9544 830
rect 9232 300 9544 352
rect 8176 58 8228 70
rect 7875 40 8040 50
rect 7038 28 8040 40
rect 6843 0 6895 6
rect 8176 0 8228 6
rect 8469 122 8521 128
rect 8469 58 8521 70
rect 8469 0 8521 6
rect 8701 122 8753 128
rect 8701 58 8753 70
rect 8701 0 8753 6
rect 8918 122 8970 128
rect 8918 58 8970 70
rect 8918 0 8970 6
rect 9232 122 9284 300
tri 9284 266 9318 300 nw
rect 9232 58 9284 70
rect 9232 0 9284 6
rect 9572 122 9624 964
rect 9652 343 9704 1300
rect 9890 11894 9942 11900
rect 9890 11812 9942 11842
rect 9890 598 9942 11760
rect 9970 11744 10022 11750
rect 9970 11680 10022 11692
rect 9970 1336 10022 11628
rect 9970 1272 10022 1284
rect 9970 1214 10022 1220
rect 9890 534 9942 546
rect 9890 476 9942 482
tri 9704 343 9738 377 sw
rect 9652 291 9836 343
tri 9750 257 9784 291 ne
rect 9572 58 9624 70
rect 9572 0 9624 6
rect 9784 122 9836 291
rect 9784 58 9836 70
rect 9784 0 9836 6
rect 10031 122 10083 128
rect 10031 58 10083 70
rect 10031 0 10083 6
rect 10263 122 10315 128
rect 10263 58 10315 70
rect 10263 0 10315 6
<< via1 >>
rect 8488 30284 8540 30336
rect 8552 30284 8604 30336
rect 8487 30082 8539 30134
rect 8551 30082 8603 30134
rect 8487 30002 8539 30054
rect 8551 30002 8603 30054
rect 8487 29922 8539 29974
rect 8551 29922 8603 29974
rect 8487 29842 8539 29894
rect 8551 29842 8603 29894
rect 8487 29762 8539 29814
rect 8551 29762 8603 29814
rect 8487 29647 8539 29699
rect 8551 29647 8603 29699
rect 8488 29408 8540 29460
rect 8552 29408 8604 29460
rect 366 27936 418 27988
rect 432 27936 484 27988
rect 366 27869 418 27921
rect 432 27869 484 27921
rect 366 27802 418 27854
rect 432 27802 484 27854
rect 366 27735 418 27787
rect 432 27735 484 27787
rect 366 27668 418 27720
rect 432 27668 484 27720
rect 366 27601 418 27653
rect 432 27601 484 27653
rect 366 27534 418 27586
rect 432 27534 484 27586
rect 366 27467 418 27519
rect 432 27467 484 27519
rect 366 27400 418 27452
rect 432 27400 484 27452
rect 2481 27936 2533 27988
rect 2547 27936 2599 27988
rect 2481 27869 2533 27921
rect 2547 27869 2599 27921
rect 2481 27802 2533 27854
rect 2547 27802 2599 27854
rect 2481 27735 2533 27787
rect 2547 27735 2599 27787
rect 2481 27668 2533 27720
rect 2547 27668 2599 27720
rect 2481 27601 2533 27653
rect 2547 27601 2599 27653
rect 2481 27534 2533 27586
rect 2547 27534 2599 27586
rect 2481 27467 2533 27519
rect 2547 27467 2599 27519
rect 2878 27903 2930 27912
rect 3008 27903 3060 27912
rect 3138 27903 3190 27912
rect 3268 27903 3320 27912
rect 3398 27903 3450 27912
rect 3528 27903 3580 27912
rect 3658 27903 3710 27912
rect 3788 27903 3840 27912
rect 3918 27903 3970 27912
rect 4048 27903 4100 27912
rect 4178 27903 4230 27912
rect 4308 27903 4360 27912
rect 4438 27903 4490 27912
rect 4568 27903 4620 27912
rect 4698 27903 4750 27912
rect 4828 27903 4880 27912
rect 4958 27903 5010 27912
rect 5088 27903 5140 27912
rect 5218 27903 5270 27912
rect 5348 27903 5400 27912
rect 5478 27903 5530 27912
rect 5608 27903 5660 27912
rect 5738 27903 5790 27912
rect 5868 27903 5920 27912
rect 5998 27903 6050 27912
rect 2878 27869 2884 27903
rect 2884 27869 2918 27903
rect 2918 27869 2930 27903
rect 3008 27869 3030 27903
rect 3030 27869 3060 27903
rect 3138 27869 3176 27903
rect 3176 27869 3190 27903
rect 3268 27869 3283 27903
rect 3283 27869 3320 27903
rect 3398 27869 3429 27903
rect 3429 27869 3450 27903
rect 3528 27869 3541 27903
rect 3541 27869 3575 27903
rect 3575 27869 3580 27903
rect 3658 27869 3687 27903
rect 3687 27869 3710 27903
rect 3788 27869 3794 27903
rect 3794 27869 3833 27903
rect 3833 27869 3840 27903
rect 3918 27869 3940 27903
rect 3940 27869 3970 27903
rect 4048 27869 4052 27903
rect 4052 27869 4086 27903
rect 4086 27869 4100 27903
rect 4178 27869 4198 27903
rect 4198 27869 4230 27903
rect 4308 27869 4344 27903
rect 4344 27869 4360 27903
rect 4438 27869 4451 27903
rect 4451 27869 4490 27903
rect 4568 27869 4597 27903
rect 4597 27869 4620 27903
rect 4698 27869 4709 27903
rect 4709 27869 4743 27903
rect 4743 27869 4750 27903
rect 4828 27869 4855 27903
rect 4855 27869 4880 27903
rect 4958 27869 4962 27903
rect 4962 27869 5001 27903
rect 5001 27869 5010 27903
rect 5088 27869 5108 27903
rect 5108 27869 5140 27903
rect 5218 27869 5220 27903
rect 5220 27869 5254 27903
rect 5254 27869 5270 27903
rect 5348 27869 5366 27903
rect 5366 27869 5400 27903
rect 5478 27869 5512 27903
rect 5512 27869 5530 27903
rect 5608 27869 5619 27903
rect 5619 27869 5658 27903
rect 5658 27869 5660 27903
rect 5738 27869 5765 27903
rect 5765 27869 5790 27903
rect 5868 27869 5877 27903
rect 5877 27869 5911 27903
rect 5911 27869 5920 27903
rect 5998 27869 6023 27903
rect 6023 27869 6050 27903
rect 2878 27860 2930 27869
rect 3008 27860 3060 27869
rect 3138 27860 3190 27869
rect 3268 27860 3320 27869
rect 3398 27860 3450 27869
rect 3528 27860 3580 27869
rect 3658 27860 3710 27869
rect 3788 27860 3840 27869
rect 3918 27860 3970 27869
rect 4048 27860 4100 27869
rect 4178 27860 4230 27869
rect 4308 27860 4360 27869
rect 4438 27860 4490 27869
rect 4568 27860 4620 27869
rect 4698 27860 4750 27869
rect 4828 27860 4880 27869
rect 4958 27860 5010 27869
rect 5088 27860 5140 27869
rect 5218 27860 5270 27869
rect 5348 27860 5400 27869
rect 5478 27860 5530 27869
rect 5608 27860 5660 27869
rect 5738 27860 5790 27869
rect 5868 27860 5920 27869
rect 5998 27860 6050 27869
rect 6128 27860 6180 27912
rect 6258 27860 6310 27912
rect 6388 27860 6440 27912
rect 6517 27860 6569 27912
rect 6646 27860 6698 27912
rect 6775 27860 6827 27912
rect 6904 27860 6956 27912
rect 7033 27860 7085 27912
rect 7162 27860 7214 27912
rect 7291 27860 7343 27912
rect 7420 27860 7472 27912
rect 7549 27860 7601 27912
rect 7678 27860 7730 27912
rect 7807 27860 7859 27912
rect 7936 27860 7988 27912
rect 2878 27823 2930 27832
rect 3008 27823 3060 27832
rect 3138 27823 3190 27832
rect 3268 27823 3320 27832
rect 3398 27823 3450 27832
rect 3528 27823 3580 27832
rect 3658 27823 3710 27832
rect 3788 27823 3840 27832
rect 3918 27823 3970 27832
rect 4048 27823 4100 27832
rect 4178 27823 4230 27832
rect 4308 27823 4360 27832
rect 4438 27823 4490 27832
rect 4568 27823 4620 27832
rect 4698 27823 4750 27832
rect 4828 27823 4880 27832
rect 4958 27823 5010 27832
rect 5088 27823 5140 27832
rect 5218 27823 5270 27832
rect 5348 27823 5400 27832
rect 5478 27823 5530 27832
rect 5608 27823 5660 27832
rect 5738 27823 5790 27832
rect 5868 27823 5920 27832
rect 5998 27823 6050 27832
rect 2878 27789 2884 27823
rect 2884 27789 2918 27823
rect 2918 27789 2930 27823
rect 3008 27789 3030 27823
rect 3030 27789 3060 27823
rect 3138 27789 3176 27823
rect 3176 27789 3190 27823
rect 3268 27789 3283 27823
rect 3283 27789 3320 27823
rect 3398 27789 3429 27823
rect 3429 27789 3450 27823
rect 3528 27789 3541 27823
rect 3541 27789 3575 27823
rect 3575 27789 3580 27823
rect 3658 27789 3687 27823
rect 3687 27789 3710 27823
rect 3788 27789 3794 27823
rect 3794 27789 3833 27823
rect 3833 27789 3840 27823
rect 3918 27789 3940 27823
rect 3940 27789 3970 27823
rect 4048 27789 4052 27823
rect 4052 27789 4086 27823
rect 4086 27789 4100 27823
rect 4178 27789 4198 27823
rect 4198 27789 4230 27823
rect 4308 27789 4344 27823
rect 4344 27789 4360 27823
rect 4438 27789 4451 27823
rect 4451 27789 4490 27823
rect 4568 27789 4597 27823
rect 4597 27789 4620 27823
rect 4698 27789 4709 27823
rect 4709 27789 4743 27823
rect 4743 27789 4750 27823
rect 4828 27789 4855 27823
rect 4855 27789 4880 27823
rect 4958 27789 4962 27823
rect 4962 27789 5001 27823
rect 5001 27789 5010 27823
rect 5088 27789 5108 27823
rect 5108 27789 5140 27823
rect 5218 27789 5220 27823
rect 5220 27789 5254 27823
rect 5254 27789 5270 27823
rect 5348 27789 5366 27823
rect 5366 27789 5400 27823
rect 5478 27789 5512 27823
rect 5512 27789 5530 27823
rect 5608 27789 5619 27823
rect 5619 27789 5658 27823
rect 5658 27789 5660 27823
rect 5738 27789 5765 27823
rect 5765 27789 5790 27823
rect 5868 27789 5877 27823
rect 5877 27789 5911 27823
rect 5911 27789 5920 27823
rect 5998 27789 6023 27823
rect 6023 27789 6050 27823
rect 2878 27780 2930 27789
rect 3008 27780 3060 27789
rect 3138 27780 3190 27789
rect 3268 27780 3320 27789
rect 3398 27780 3450 27789
rect 3528 27780 3580 27789
rect 3658 27780 3710 27789
rect 3788 27780 3840 27789
rect 3918 27780 3970 27789
rect 4048 27780 4100 27789
rect 4178 27780 4230 27789
rect 4308 27780 4360 27789
rect 4438 27780 4490 27789
rect 4568 27780 4620 27789
rect 4698 27780 4750 27789
rect 4828 27780 4880 27789
rect 4958 27780 5010 27789
rect 5088 27780 5140 27789
rect 5218 27780 5270 27789
rect 5348 27780 5400 27789
rect 5478 27780 5530 27789
rect 5608 27780 5660 27789
rect 5738 27780 5790 27789
rect 5868 27780 5920 27789
rect 5998 27780 6050 27789
rect 6128 27780 6180 27832
rect 6258 27780 6310 27832
rect 6388 27780 6440 27832
rect 6517 27780 6569 27832
rect 6646 27780 6698 27832
rect 6775 27780 6827 27832
rect 6904 27780 6956 27832
rect 7033 27780 7085 27832
rect 7162 27780 7214 27832
rect 7291 27780 7343 27832
rect 7420 27780 7472 27832
rect 7549 27780 7601 27832
rect 7678 27780 7730 27832
rect 7807 27780 7859 27832
rect 7936 27780 7988 27832
rect 2878 27743 2930 27752
rect 3008 27743 3060 27752
rect 3138 27743 3190 27752
rect 3268 27743 3320 27752
rect 3398 27743 3450 27752
rect 3528 27743 3580 27752
rect 3658 27743 3710 27752
rect 3788 27743 3840 27752
rect 3918 27743 3970 27752
rect 4048 27743 4100 27752
rect 4178 27743 4230 27752
rect 4308 27743 4360 27752
rect 4438 27743 4490 27752
rect 4568 27743 4620 27752
rect 4698 27743 4750 27752
rect 4828 27743 4880 27752
rect 4958 27743 5010 27752
rect 5088 27743 5140 27752
rect 5218 27743 5270 27752
rect 5348 27743 5400 27752
rect 5478 27743 5530 27752
rect 5608 27743 5660 27752
rect 5738 27743 5790 27752
rect 5868 27743 5920 27752
rect 5998 27743 6050 27752
rect 2878 27709 2884 27743
rect 2884 27709 2918 27743
rect 2918 27709 2930 27743
rect 3008 27709 3030 27743
rect 3030 27709 3060 27743
rect 3138 27709 3176 27743
rect 3176 27709 3190 27743
rect 3268 27709 3283 27743
rect 3283 27709 3320 27743
rect 3398 27709 3429 27743
rect 3429 27709 3450 27743
rect 3528 27709 3541 27743
rect 3541 27709 3575 27743
rect 3575 27709 3580 27743
rect 3658 27709 3687 27743
rect 3687 27709 3710 27743
rect 3788 27709 3794 27743
rect 3794 27709 3833 27743
rect 3833 27709 3840 27743
rect 3918 27709 3940 27743
rect 3940 27709 3970 27743
rect 4048 27709 4052 27743
rect 4052 27709 4086 27743
rect 4086 27709 4100 27743
rect 4178 27709 4198 27743
rect 4198 27709 4230 27743
rect 4308 27709 4344 27743
rect 4344 27709 4360 27743
rect 4438 27709 4451 27743
rect 4451 27709 4490 27743
rect 4568 27709 4597 27743
rect 4597 27709 4620 27743
rect 4698 27709 4709 27743
rect 4709 27709 4743 27743
rect 4743 27709 4750 27743
rect 4828 27709 4855 27743
rect 4855 27709 4880 27743
rect 4958 27709 4962 27743
rect 4962 27709 5001 27743
rect 5001 27709 5010 27743
rect 5088 27709 5108 27743
rect 5108 27709 5140 27743
rect 5218 27709 5220 27743
rect 5220 27709 5254 27743
rect 5254 27709 5270 27743
rect 5348 27709 5366 27743
rect 5366 27709 5400 27743
rect 5478 27709 5512 27743
rect 5512 27709 5530 27743
rect 5608 27709 5619 27743
rect 5619 27709 5658 27743
rect 5658 27709 5660 27743
rect 5738 27709 5765 27743
rect 5765 27709 5790 27743
rect 5868 27709 5877 27743
rect 5877 27709 5911 27743
rect 5911 27709 5920 27743
rect 5998 27709 6023 27743
rect 6023 27709 6050 27743
rect 2878 27700 2930 27709
rect 3008 27700 3060 27709
rect 3138 27700 3190 27709
rect 3268 27700 3320 27709
rect 3398 27700 3450 27709
rect 3528 27700 3580 27709
rect 3658 27700 3710 27709
rect 3788 27700 3840 27709
rect 3918 27700 3970 27709
rect 4048 27700 4100 27709
rect 4178 27700 4230 27709
rect 4308 27700 4360 27709
rect 4438 27700 4490 27709
rect 4568 27700 4620 27709
rect 4698 27700 4750 27709
rect 4828 27700 4880 27709
rect 4958 27700 5010 27709
rect 5088 27700 5140 27709
rect 5218 27700 5270 27709
rect 5348 27700 5400 27709
rect 5478 27700 5530 27709
rect 5608 27700 5660 27709
rect 5738 27700 5790 27709
rect 5868 27700 5920 27709
rect 5998 27700 6050 27709
rect 6128 27700 6180 27752
rect 6258 27700 6310 27752
rect 6388 27700 6440 27752
rect 6517 27700 6569 27752
rect 6646 27700 6698 27752
rect 6775 27700 6827 27752
rect 6904 27700 6956 27752
rect 7033 27700 7085 27752
rect 7162 27700 7214 27752
rect 7291 27700 7343 27752
rect 7420 27700 7472 27752
rect 7549 27700 7601 27752
rect 7678 27700 7730 27752
rect 7807 27700 7859 27752
rect 7936 27700 7988 27752
rect 2878 27663 2930 27672
rect 3008 27663 3060 27672
rect 3138 27663 3190 27672
rect 3268 27663 3320 27672
rect 3398 27663 3450 27672
rect 3528 27663 3580 27672
rect 3658 27663 3710 27672
rect 3788 27663 3840 27672
rect 3918 27663 3970 27672
rect 4048 27663 4100 27672
rect 4178 27663 4230 27672
rect 4308 27663 4360 27672
rect 4438 27663 4490 27672
rect 4568 27663 4620 27672
rect 4698 27663 4750 27672
rect 4828 27663 4880 27672
rect 4958 27663 5010 27672
rect 5088 27663 5140 27672
rect 5218 27663 5270 27672
rect 5348 27663 5400 27672
rect 5478 27663 5530 27672
rect 5608 27663 5660 27672
rect 5738 27663 5790 27672
rect 5868 27663 5920 27672
rect 5998 27663 6050 27672
rect 2878 27629 2884 27663
rect 2884 27629 2918 27663
rect 2918 27629 2930 27663
rect 3008 27629 3030 27663
rect 3030 27629 3060 27663
rect 3138 27629 3176 27663
rect 3176 27629 3190 27663
rect 3268 27629 3283 27663
rect 3283 27629 3320 27663
rect 3398 27629 3429 27663
rect 3429 27629 3450 27663
rect 3528 27629 3541 27663
rect 3541 27629 3575 27663
rect 3575 27629 3580 27663
rect 3658 27629 3687 27663
rect 3687 27629 3710 27663
rect 3788 27629 3794 27663
rect 3794 27629 3833 27663
rect 3833 27629 3840 27663
rect 3918 27629 3940 27663
rect 3940 27629 3970 27663
rect 4048 27629 4052 27663
rect 4052 27629 4086 27663
rect 4086 27629 4100 27663
rect 4178 27629 4198 27663
rect 4198 27629 4230 27663
rect 4308 27629 4344 27663
rect 4344 27629 4360 27663
rect 4438 27629 4451 27663
rect 4451 27629 4490 27663
rect 4568 27629 4597 27663
rect 4597 27629 4620 27663
rect 4698 27629 4709 27663
rect 4709 27629 4743 27663
rect 4743 27629 4750 27663
rect 4828 27629 4855 27663
rect 4855 27629 4880 27663
rect 4958 27629 4962 27663
rect 4962 27629 5001 27663
rect 5001 27629 5010 27663
rect 5088 27629 5108 27663
rect 5108 27629 5140 27663
rect 5218 27629 5220 27663
rect 5220 27629 5254 27663
rect 5254 27629 5270 27663
rect 5348 27629 5366 27663
rect 5366 27629 5400 27663
rect 5478 27629 5512 27663
rect 5512 27629 5530 27663
rect 5608 27629 5619 27663
rect 5619 27629 5658 27663
rect 5658 27629 5660 27663
rect 5738 27629 5765 27663
rect 5765 27629 5790 27663
rect 5868 27629 5877 27663
rect 5877 27629 5911 27663
rect 5911 27629 5920 27663
rect 5998 27629 6023 27663
rect 6023 27629 6050 27663
rect 2878 27620 2930 27629
rect 3008 27620 3060 27629
rect 3138 27620 3190 27629
rect 3268 27620 3320 27629
rect 3398 27620 3450 27629
rect 3528 27620 3580 27629
rect 3658 27620 3710 27629
rect 3788 27620 3840 27629
rect 3918 27620 3970 27629
rect 4048 27620 4100 27629
rect 4178 27620 4230 27629
rect 4308 27620 4360 27629
rect 4438 27620 4490 27629
rect 4568 27620 4620 27629
rect 4698 27620 4750 27629
rect 4828 27620 4880 27629
rect 4958 27620 5010 27629
rect 5088 27620 5140 27629
rect 5218 27620 5270 27629
rect 5348 27620 5400 27629
rect 5478 27620 5530 27629
rect 5608 27620 5660 27629
rect 5738 27620 5790 27629
rect 5868 27620 5920 27629
rect 5998 27620 6050 27629
rect 6128 27620 6180 27672
rect 6258 27620 6310 27672
rect 6388 27620 6440 27672
rect 6517 27620 6569 27672
rect 6646 27620 6698 27672
rect 6775 27620 6827 27672
rect 6904 27620 6956 27672
rect 7033 27620 7085 27672
rect 7162 27620 7214 27672
rect 7291 27620 7343 27672
rect 7420 27620 7472 27672
rect 7549 27620 7601 27672
rect 7678 27620 7730 27672
rect 7807 27620 7859 27672
rect 7936 27620 7988 27672
rect 2878 27583 2930 27592
rect 3008 27583 3060 27592
rect 3138 27583 3190 27592
rect 3268 27583 3320 27592
rect 3398 27583 3450 27592
rect 3528 27583 3580 27592
rect 3658 27583 3710 27592
rect 3788 27583 3840 27592
rect 3918 27583 3970 27592
rect 4048 27583 4100 27592
rect 4178 27583 4230 27592
rect 4308 27583 4360 27592
rect 4438 27583 4490 27592
rect 4568 27583 4620 27592
rect 4698 27583 4750 27592
rect 4828 27583 4880 27592
rect 4958 27583 5010 27592
rect 5088 27583 5140 27592
rect 5218 27583 5270 27592
rect 5348 27583 5400 27592
rect 5478 27583 5530 27592
rect 5608 27583 5660 27592
rect 5738 27583 5790 27592
rect 5868 27583 5920 27592
rect 5998 27583 6050 27592
rect 2878 27549 2884 27583
rect 2884 27549 2918 27583
rect 2918 27549 2930 27583
rect 3008 27549 3030 27583
rect 3030 27549 3060 27583
rect 3138 27549 3176 27583
rect 3176 27549 3190 27583
rect 3268 27549 3283 27583
rect 3283 27549 3320 27583
rect 3398 27549 3429 27583
rect 3429 27549 3450 27583
rect 3528 27549 3541 27583
rect 3541 27549 3575 27583
rect 3575 27549 3580 27583
rect 3658 27549 3687 27583
rect 3687 27549 3710 27583
rect 3788 27549 3794 27583
rect 3794 27549 3833 27583
rect 3833 27549 3840 27583
rect 3918 27549 3940 27583
rect 3940 27549 3970 27583
rect 4048 27549 4052 27583
rect 4052 27549 4086 27583
rect 4086 27549 4100 27583
rect 4178 27549 4198 27583
rect 4198 27549 4230 27583
rect 4308 27549 4344 27583
rect 4344 27549 4360 27583
rect 4438 27549 4451 27583
rect 4451 27549 4490 27583
rect 4568 27549 4597 27583
rect 4597 27549 4620 27583
rect 4698 27549 4709 27583
rect 4709 27549 4743 27583
rect 4743 27549 4750 27583
rect 4828 27549 4855 27583
rect 4855 27549 4880 27583
rect 4958 27549 4962 27583
rect 4962 27549 5001 27583
rect 5001 27549 5010 27583
rect 5088 27549 5108 27583
rect 5108 27549 5140 27583
rect 5218 27549 5220 27583
rect 5220 27549 5254 27583
rect 5254 27549 5270 27583
rect 5348 27549 5366 27583
rect 5366 27549 5400 27583
rect 5478 27549 5512 27583
rect 5512 27549 5530 27583
rect 5608 27549 5619 27583
rect 5619 27549 5658 27583
rect 5658 27549 5660 27583
rect 5738 27549 5765 27583
rect 5765 27549 5790 27583
rect 5868 27549 5877 27583
rect 5877 27549 5911 27583
rect 5911 27549 5920 27583
rect 5998 27549 6023 27583
rect 6023 27549 6050 27583
rect 2878 27540 2930 27549
rect 3008 27540 3060 27549
rect 3138 27540 3190 27549
rect 3268 27540 3320 27549
rect 3398 27540 3450 27549
rect 3528 27540 3580 27549
rect 3658 27540 3710 27549
rect 3788 27540 3840 27549
rect 3918 27540 3970 27549
rect 4048 27540 4100 27549
rect 4178 27540 4230 27549
rect 4308 27540 4360 27549
rect 4438 27540 4490 27549
rect 4568 27540 4620 27549
rect 4698 27540 4750 27549
rect 4828 27540 4880 27549
rect 4958 27540 5010 27549
rect 5088 27540 5140 27549
rect 5218 27540 5270 27549
rect 5348 27540 5400 27549
rect 5478 27540 5530 27549
rect 5608 27540 5660 27549
rect 5738 27540 5790 27549
rect 5868 27540 5920 27549
rect 5998 27540 6050 27549
rect 6128 27540 6180 27592
rect 6258 27540 6310 27592
rect 6388 27540 6440 27592
rect 6517 27540 6569 27592
rect 6646 27540 6698 27592
rect 6775 27540 6827 27592
rect 6904 27540 6956 27592
rect 7033 27540 7085 27592
rect 7162 27540 7214 27592
rect 7291 27540 7343 27592
rect 7420 27540 7472 27592
rect 7549 27540 7601 27592
rect 7678 27540 7730 27592
rect 7807 27540 7859 27592
rect 7936 27540 7988 27592
rect 2878 27503 2930 27512
rect 3008 27503 3060 27512
rect 3138 27503 3190 27512
rect 3268 27503 3320 27512
rect 3398 27503 3450 27512
rect 3528 27503 3580 27512
rect 3658 27503 3710 27512
rect 3788 27503 3840 27512
rect 3918 27503 3970 27512
rect 4048 27503 4100 27512
rect 4178 27503 4230 27512
rect 4308 27503 4360 27512
rect 4438 27503 4490 27512
rect 4568 27503 4620 27512
rect 4698 27503 4750 27512
rect 4828 27503 4880 27512
rect 4958 27503 5010 27512
rect 5088 27503 5140 27512
rect 5218 27503 5270 27512
rect 5348 27503 5400 27512
rect 5478 27503 5530 27512
rect 5608 27503 5660 27512
rect 5738 27503 5790 27512
rect 5868 27503 5920 27512
rect 5998 27503 6050 27512
rect 2878 27469 2884 27503
rect 2884 27469 2918 27503
rect 2918 27469 2930 27503
rect 3008 27469 3030 27503
rect 3030 27469 3060 27503
rect 3138 27469 3176 27503
rect 3176 27469 3190 27503
rect 3268 27469 3283 27503
rect 3283 27469 3320 27503
rect 3398 27469 3429 27503
rect 3429 27469 3450 27503
rect 3528 27469 3541 27503
rect 3541 27469 3575 27503
rect 3575 27469 3580 27503
rect 3658 27469 3687 27503
rect 3687 27469 3710 27503
rect 3788 27469 3794 27503
rect 3794 27469 3833 27503
rect 3833 27469 3840 27503
rect 3918 27469 3940 27503
rect 3940 27469 3970 27503
rect 4048 27469 4052 27503
rect 4052 27469 4086 27503
rect 4086 27469 4100 27503
rect 4178 27469 4198 27503
rect 4198 27469 4230 27503
rect 4308 27469 4344 27503
rect 4344 27469 4360 27503
rect 4438 27469 4451 27503
rect 4451 27469 4490 27503
rect 4568 27469 4597 27503
rect 4597 27469 4620 27503
rect 4698 27469 4709 27503
rect 4709 27469 4743 27503
rect 4743 27469 4750 27503
rect 4828 27469 4855 27503
rect 4855 27469 4880 27503
rect 4958 27469 4962 27503
rect 4962 27469 5001 27503
rect 5001 27469 5010 27503
rect 5088 27469 5108 27503
rect 5108 27469 5140 27503
rect 5218 27469 5220 27503
rect 5220 27469 5254 27503
rect 5254 27469 5270 27503
rect 5348 27469 5366 27503
rect 5366 27469 5400 27503
rect 5478 27469 5512 27503
rect 5512 27469 5530 27503
rect 5608 27469 5619 27503
rect 5619 27469 5658 27503
rect 5658 27469 5660 27503
rect 5738 27469 5765 27503
rect 5765 27469 5790 27503
rect 5868 27469 5877 27503
rect 5877 27469 5911 27503
rect 5911 27469 5920 27503
rect 5998 27469 6023 27503
rect 6023 27469 6050 27503
rect 2878 27460 2930 27469
rect 3008 27460 3060 27469
rect 3138 27460 3190 27469
rect 3268 27460 3320 27469
rect 3398 27460 3450 27469
rect 3528 27460 3580 27469
rect 3658 27460 3710 27469
rect 3788 27460 3840 27469
rect 3918 27460 3970 27469
rect 4048 27460 4100 27469
rect 4178 27460 4230 27469
rect 4308 27460 4360 27469
rect 4438 27460 4490 27469
rect 4568 27460 4620 27469
rect 4698 27460 4750 27469
rect 4828 27460 4880 27469
rect 4958 27460 5010 27469
rect 5088 27460 5140 27469
rect 5218 27460 5270 27469
rect 5348 27460 5400 27469
rect 5478 27460 5530 27469
rect 5608 27460 5660 27469
rect 5738 27460 5790 27469
rect 5868 27460 5920 27469
rect 5998 27460 6050 27469
rect 6128 27460 6180 27512
rect 6258 27460 6310 27512
rect 6388 27460 6440 27512
rect 6517 27460 6569 27512
rect 6646 27460 6698 27512
rect 6775 27460 6827 27512
rect 6904 27460 6956 27512
rect 7033 27460 7085 27512
rect 7162 27460 7214 27512
rect 7291 27460 7343 27512
rect 7420 27460 7472 27512
rect 7549 27460 7601 27512
rect 7678 27460 7730 27512
rect 7807 27460 7859 27512
rect 7936 27460 7988 27512
rect 2481 27400 2533 27452
rect 2547 27400 2599 27452
rect 9732 27936 9784 27988
rect 9810 27936 9862 27988
rect 9732 27869 9784 27921
rect 9810 27869 9862 27921
rect 9732 27802 9784 27854
rect 9810 27802 9862 27854
rect 9732 27735 9784 27787
rect 9810 27735 9862 27787
rect 9732 27668 9784 27720
rect 9810 27668 9862 27720
rect 9732 27601 9784 27653
rect 9810 27601 9862 27653
rect 9732 27534 9784 27586
rect 9810 27534 9862 27586
rect 9732 27467 9784 27519
rect 9810 27467 9862 27519
rect 9732 27400 9784 27452
rect 9810 27400 9862 27452
rect 3310 27330 3362 27336
rect 3376 27330 3428 27336
rect 3310 27284 3316 27330
rect 3316 27284 3362 27330
rect 3376 27284 3422 27330
rect 3422 27284 3428 27330
rect 3310 27224 3316 27270
rect 3316 27224 3362 27270
rect 3376 27224 3422 27270
rect 3422 27224 3428 27270
rect 3310 27218 3362 27224
rect 3376 27218 3428 27224
rect 5389 27329 5505 27334
rect 5389 27223 5395 27329
rect 5395 27223 5501 27329
rect 5501 27223 5505 27329
rect 5389 27218 5505 27223
rect 3269 26795 3321 26847
rect 3337 26795 3389 26847
rect 3405 26795 3457 26847
rect 3269 26711 3321 26763
rect 3337 26711 3389 26763
rect 3405 26711 3457 26763
rect 3269 26627 3321 26679
rect 3337 26627 3389 26679
rect 3405 26627 3457 26679
rect 3269 26542 3321 26594
rect 3337 26542 3389 26594
rect 3405 26542 3457 26594
rect 3269 26457 3321 26509
rect 3337 26457 3389 26509
rect 3405 26457 3457 26509
rect 4056 24517 4108 24522
rect 4187 24517 4239 24522
rect 4318 24517 4370 24522
rect 4449 24517 4501 24522
rect 4580 24517 4632 24522
rect 4711 24517 4763 24522
rect 4842 24517 4894 24522
rect 4973 24517 5025 24522
rect 5104 24517 5156 24522
rect 5235 24517 5287 24522
rect 5365 24517 5417 24522
rect 5495 24517 5547 24522
rect 5625 24517 5677 24522
rect 5755 24517 5807 24522
rect 5885 24517 5937 24522
rect 6015 24517 6067 24522
rect 4056 24483 4062 24517
rect 4062 24483 4096 24517
rect 4096 24483 4108 24517
rect 4187 24483 4208 24517
rect 4208 24483 4239 24517
rect 4318 24483 4354 24517
rect 4354 24483 4370 24517
rect 4449 24483 4461 24517
rect 4461 24483 4500 24517
rect 4500 24483 4501 24517
rect 4580 24483 4607 24517
rect 4607 24483 4632 24517
rect 4711 24483 4719 24517
rect 4719 24483 4753 24517
rect 4753 24483 4763 24517
rect 4842 24483 4865 24517
rect 4865 24483 4894 24517
rect 4973 24483 5011 24517
rect 5011 24483 5025 24517
rect 5104 24483 5118 24517
rect 5118 24483 5156 24517
rect 5235 24483 5264 24517
rect 5264 24483 5287 24517
rect 5365 24483 5376 24517
rect 5376 24483 5410 24517
rect 5410 24483 5417 24517
rect 5495 24483 5522 24517
rect 5522 24483 5547 24517
rect 5625 24483 5629 24517
rect 5629 24483 5667 24517
rect 5667 24483 5677 24517
rect 5755 24483 5773 24517
rect 5773 24483 5807 24517
rect 5885 24483 5917 24517
rect 5917 24483 5937 24517
rect 6015 24483 6027 24517
rect 6027 24483 6061 24517
rect 6061 24483 6067 24517
rect 4056 24470 4108 24483
rect 4187 24470 4239 24483
rect 4318 24470 4370 24483
rect 4449 24470 4501 24483
rect 4580 24470 4632 24483
rect 4711 24470 4763 24483
rect 4842 24470 4894 24483
rect 4973 24470 5025 24483
rect 5104 24470 5156 24483
rect 5235 24470 5287 24483
rect 5365 24470 5417 24483
rect 5495 24470 5547 24483
rect 5625 24470 5677 24483
rect 5755 24470 5807 24483
rect 5885 24470 5937 24483
rect 6015 24470 6067 24483
rect 4056 24406 4108 24458
rect 4187 24406 4239 24458
rect 4318 24406 4370 24458
rect 4449 24406 4501 24458
rect 4580 24406 4632 24458
rect 4711 24406 4763 24458
rect 4842 24406 4894 24458
rect 4973 24406 5025 24458
rect 5104 24406 5156 24458
rect 5235 24406 5287 24458
rect 5365 24406 5417 24458
rect 5495 24406 5547 24458
rect 5625 24406 5677 24458
rect 5755 24406 5807 24458
rect 5885 24406 5937 24458
rect 6015 24406 6067 24458
rect 4056 24381 4108 24394
rect 4187 24381 4239 24394
rect 4318 24381 4370 24394
rect 4449 24381 4501 24394
rect 4580 24381 4632 24394
rect 4711 24381 4763 24394
rect 4842 24381 4894 24394
rect 4973 24381 5025 24394
rect 5104 24381 5156 24394
rect 5235 24381 5287 24394
rect 5365 24381 5417 24394
rect 5495 24381 5547 24394
rect 5625 24381 5677 24394
rect 5755 24381 5807 24394
rect 5885 24381 5937 24394
rect 6015 24381 6067 24394
rect 4056 24347 4062 24381
rect 4062 24347 4096 24381
rect 4096 24347 4108 24381
rect 4187 24347 4208 24381
rect 4208 24347 4239 24381
rect 4318 24347 4354 24381
rect 4354 24347 4370 24381
rect 4449 24347 4461 24381
rect 4461 24347 4500 24381
rect 4500 24347 4501 24381
rect 4580 24347 4607 24381
rect 4607 24347 4632 24381
rect 4711 24347 4719 24381
rect 4719 24347 4753 24381
rect 4753 24347 4763 24381
rect 4842 24347 4865 24381
rect 4865 24347 4894 24381
rect 4973 24347 5011 24381
rect 5011 24347 5025 24381
rect 5104 24347 5118 24381
rect 5118 24347 5156 24381
rect 5235 24347 5264 24381
rect 5264 24347 5287 24381
rect 5365 24347 5376 24381
rect 5376 24347 5410 24381
rect 5410 24347 5417 24381
rect 5495 24347 5522 24381
rect 5522 24347 5547 24381
rect 5625 24347 5629 24381
rect 5629 24347 5667 24381
rect 5667 24347 5677 24381
rect 5755 24347 5773 24381
rect 5773 24347 5807 24381
rect 5885 24347 5917 24381
rect 5917 24347 5937 24381
rect 6015 24347 6027 24381
rect 6027 24347 6061 24381
rect 6061 24347 6067 24381
rect 4056 24342 4108 24347
rect 4187 24342 4239 24347
rect 4318 24342 4370 24347
rect 4449 24342 4501 24347
rect 4580 24342 4632 24347
rect 4711 24342 4763 24347
rect 4842 24342 4894 24347
rect 4973 24342 5025 24347
rect 5104 24342 5156 24347
rect 5235 24342 5287 24347
rect 5365 24342 5417 24347
rect 5495 24342 5547 24347
rect 5625 24342 5677 24347
rect 5755 24342 5807 24347
rect 5885 24342 5937 24347
rect 6015 24342 6067 24347
rect 7988 24465 8040 24517
rect 7988 24347 8040 24399
rect 9732 24465 9784 24517
rect 9810 24465 9862 24517
rect 9732 24347 9784 24399
rect 9810 24347 9862 24399
rect 10710 24465 10762 24517
rect 10776 24465 10828 24517
rect 10710 24347 10762 24399
rect 10776 24347 10828 24399
rect 282 22697 334 22749
rect 282 22633 334 22685
rect 6056 23256 6108 23265
rect 6123 23256 6175 23265
rect 6190 23256 6242 23265
rect 6257 23256 6309 23265
rect 6324 23256 6376 23265
rect 6391 23256 6443 23265
rect 6458 23256 6510 23265
rect 6525 23256 6577 23265
rect 6592 23256 6644 23265
rect 6659 23256 6711 23265
rect 6726 23256 6778 23265
rect 6792 23256 6844 23265
rect 6858 23256 6910 23265
rect 6924 23256 6976 23265
rect 6990 23256 7042 23265
rect 7056 23256 7108 23265
rect 7122 23256 7174 23265
rect 7188 23256 7240 23265
rect 7254 23256 7306 23265
rect 7320 23256 7372 23265
rect 7386 23256 7438 23265
rect 7452 23256 7504 23265
rect 7518 23256 7570 23265
rect 7584 23256 7636 23265
rect 7650 23256 7702 23265
rect 7716 23256 7768 23265
rect 6056 23213 6067 23256
rect 6067 23213 6108 23256
rect 6123 23213 6175 23256
rect 6190 23213 6242 23256
rect 6257 23213 6309 23256
rect 6324 23213 6376 23256
rect 6391 23213 6443 23256
rect 6458 23213 6510 23256
rect 6525 23213 6577 23256
rect 6592 23213 6644 23256
rect 6659 23213 6711 23256
rect 6726 23213 6778 23256
rect 6792 23213 6844 23256
rect 6858 23213 6910 23256
rect 6924 23213 6976 23256
rect 6990 23213 7042 23256
rect 7056 23213 7108 23256
rect 7122 23213 7174 23256
rect 7188 23213 7240 23256
rect 7254 23213 7306 23256
rect 7320 23213 7372 23256
rect 7386 23213 7438 23256
rect 7452 23213 7504 23256
rect 7518 23213 7570 23256
rect 7584 23213 7636 23256
rect 7650 23213 7702 23256
rect 7716 23213 7757 23256
rect 7757 23213 7768 23256
rect 6056 23143 6067 23195
rect 6067 23143 6108 23195
rect 6123 23143 6175 23195
rect 6190 23143 6242 23195
rect 6257 23143 6309 23195
rect 6324 23143 6376 23195
rect 6391 23143 6443 23195
rect 6458 23143 6510 23195
rect 6525 23143 6577 23195
rect 6592 23143 6644 23195
rect 6659 23143 6711 23195
rect 6726 23143 6778 23195
rect 6792 23143 6844 23195
rect 6858 23143 6910 23195
rect 6924 23143 6976 23195
rect 6990 23143 7042 23195
rect 7056 23143 7108 23195
rect 7122 23143 7174 23195
rect 7188 23143 7240 23195
rect 7254 23143 7306 23195
rect 7320 23143 7372 23195
rect 7386 23143 7438 23195
rect 7452 23143 7504 23195
rect 7518 23143 7570 23195
rect 7584 23143 7636 23195
rect 7650 23143 7702 23195
rect 7716 23143 7757 23195
rect 7757 23143 7768 23195
rect 6056 23073 6067 23125
rect 6067 23073 6108 23125
rect 6123 23073 6175 23125
rect 6190 23073 6242 23125
rect 6257 23073 6309 23125
rect 6324 23073 6376 23125
rect 6391 23073 6443 23125
rect 6458 23073 6510 23125
rect 6525 23073 6577 23125
rect 6592 23073 6644 23125
rect 6659 23073 6711 23125
rect 6726 23073 6778 23125
rect 6792 23073 6844 23125
rect 6858 23073 6910 23125
rect 6924 23073 6976 23125
rect 6990 23073 7042 23125
rect 7056 23073 7108 23125
rect 7122 23073 7174 23125
rect 7188 23073 7240 23125
rect 7254 23073 7306 23125
rect 7320 23073 7372 23125
rect 7386 23073 7438 23125
rect 7452 23073 7504 23125
rect 7518 23073 7570 23125
rect 7584 23073 7636 23125
rect 7650 23073 7702 23125
rect 7716 23073 7757 23125
rect 7757 23073 7768 23125
rect 6056 23003 6067 23055
rect 6067 23003 6108 23055
rect 6123 23003 6175 23055
rect 6190 23003 6242 23055
rect 6257 23003 6309 23055
rect 6324 23003 6376 23055
rect 6391 23003 6443 23055
rect 6458 23003 6510 23055
rect 6525 23003 6577 23055
rect 6592 23003 6644 23055
rect 6659 23003 6711 23055
rect 6726 23003 6778 23055
rect 6792 23003 6844 23055
rect 6858 23003 6910 23055
rect 6924 23003 6976 23055
rect 6990 23003 7042 23055
rect 7056 23003 7108 23055
rect 7122 23003 7174 23055
rect 7188 23003 7240 23055
rect 7254 23003 7306 23055
rect 7320 23003 7372 23055
rect 7386 23003 7438 23055
rect 7452 23003 7504 23055
rect 7518 23003 7570 23055
rect 7584 23003 7636 23055
rect 7650 23003 7702 23055
rect 7716 23003 7757 23055
rect 7757 23003 7768 23055
rect 6056 22933 6067 22985
rect 6067 22933 6108 22985
rect 6123 22933 6175 22985
rect 6190 22933 6242 22985
rect 6257 22933 6309 22985
rect 6324 22933 6376 22985
rect 6391 22933 6443 22985
rect 6458 22933 6510 22985
rect 6525 22933 6577 22985
rect 6592 22933 6644 22985
rect 6659 22933 6711 22985
rect 6726 22933 6778 22985
rect 6792 22933 6844 22985
rect 6858 22933 6910 22985
rect 6924 22933 6976 22985
rect 6990 22933 7042 22985
rect 7056 22933 7108 22985
rect 7122 22933 7174 22985
rect 7188 22933 7240 22985
rect 7254 22933 7306 22985
rect 7320 22933 7372 22985
rect 7386 22933 7438 22985
rect 7452 22933 7504 22985
rect 7518 22933 7570 22985
rect 7584 22933 7636 22985
rect 7650 22933 7702 22985
rect 7716 22933 7757 22985
rect 7757 22933 7768 22985
rect 6056 22863 6067 22915
rect 6067 22863 6108 22915
rect 6123 22863 6175 22915
rect 6190 22863 6242 22915
rect 6257 22863 6309 22915
rect 6324 22863 6376 22915
rect 6391 22863 6443 22915
rect 6458 22863 6510 22915
rect 6525 22863 6577 22915
rect 6592 22863 6644 22915
rect 6659 22863 6711 22915
rect 6726 22863 6778 22915
rect 6792 22863 6844 22915
rect 6858 22863 6910 22915
rect 6924 22863 6976 22915
rect 6990 22863 7042 22915
rect 7056 22863 7108 22915
rect 7122 22863 7174 22915
rect 7188 22863 7240 22915
rect 7254 22863 7306 22915
rect 7320 22863 7372 22915
rect 7386 22863 7438 22915
rect 7452 22863 7504 22915
rect 7518 22863 7570 22915
rect 7584 22863 7636 22915
rect 7650 22863 7702 22915
rect 7716 22863 7757 22915
rect 7757 22863 7768 22915
rect 8229 22703 8281 22755
rect 8293 22703 8345 22755
rect 6847 21100 6899 21152
rect 6949 21100 7001 21152
rect 7051 21100 7103 21152
rect 6847 21016 6899 21068
rect 6949 21016 7001 21068
rect 7051 21016 7103 21068
rect 6847 20932 6899 20984
rect 6949 20932 7001 20984
rect 7051 20932 7103 20984
rect 6847 20848 6899 20900
rect 6949 20848 7001 20900
rect 7051 20848 7103 20900
rect 6847 20764 6899 20816
rect 6949 20764 7001 20816
rect 7051 20764 7103 20816
rect 6015 19887 6067 19939
rect 6079 19887 6131 19939
rect 6165 19756 6217 19808
rect 6165 19692 6217 19744
rect 6015 19575 6067 19627
rect 6079 19575 6131 19627
rect 6364 19550 6416 19557
rect 6364 19516 6373 19550
rect 6373 19516 6407 19550
rect 6407 19516 6416 19550
rect 6165 19455 6217 19507
rect 6364 19505 6416 19516
rect 6364 19478 6416 19493
rect 6165 19391 6217 19443
rect 6364 19444 6373 19478
rect 6373 19444 6407 19478
rect 6407 19444 6416 19478
rect 6364 19441 6416 19444
rect 7710 21100 7762 21152
rect 7710 21033 7762 21085
rect 7710 20966 7762 21018
rect 7710 20899 7762 20951
rect 7710 20832 7762 20884
rect 7710 20764 7762 20816
rect 7710 19666 7762 19672
rect 7710 19632 7716 19666
rect 7716 19632 7750 19666
rect 7750 19632 7762 19666
rect 7710 19620 7762 19632
rect 7710 19560 7716 19573
rect 7716 19560 7750 19573
rect 7750 19560 7762 19573
rect 7710 19522 7762 19560
rect 7710 19521 7716 19522
rect 7716 19521 7750 19522
rect 7750 19521 7762 19522
rect 8711 19756 8763 19808
rect 8711 19692 8763 19744
rect 6015 19263 6067 19315
rect 6079 19263 6131 19315
rect 6165 19130 6217 19182
rect 6165 19066 6217 19118
rect 6364 19081 6416 19089
rect 6364 19047 6373 19081
rect 6373 19047 6407 19081
rect 6407 19047 6416 19081
rect 6364 19037 6416 19047
rect 6364 19006 6416 19025
rect 6015 18951 6067 19003
rect 6079 18951 6131 19003
rect 6364 18973 6373 19006
rect 6373 18973 6407 19006
rect 6407 18973 6416 19006
rect 6165 18834 6217 18886
rect 6165 18770 6217 18822
rect 7524 18845 7530 18856
rect 7530 18845 7564 18856
rect 7564 18845 7576 18856
rect 7524 18804 7576 18845
rect 7524 18740 7576 18792
rect 6015 18639 6067 18691
rect 6079 18639 6131 18691
rect 6364 18614 6416 18625
rect 6364 18580 6373 18614
rect 6373 18580 6407 18614
rect 6407 18580 6416 18614
rect 6364 18573 6416 18580
rect 3839 18436 3891 18488
rect 3924 18436 3976 18488
rect 4009 18436 4061 18488
rect 4093 18436 4145 18488
rect 4177 18436 4229 18488
rect 6245 18510 6297 18562
rect 6245 18446 6297 18498
rect 6364 18542 6416 18561
rect 6364 18509 6373 18542
rect 6373 18509 6407 18542
rect 6407 18509 6416 18542
rect 3839 18356 3891 18408
rect 3924 18356 3976 18408
rect 4009 18356 4061 18408
rect 4093 18356 4145 18408
rect 4177 18356 4229 18408
rect 8631 19429 8683 19481
rect 8631 19365 8683 19417
rect 8551 19167 8603 19219
rect 8551 19103 8603 19155
rect 8471 19037 8523 19089
rect 8471 18973 8523 19025
rect 7618 18284 7624 18317
rect 7624 18284 7658 18317
rect 7658 18284 7670 18317
rect 7618 18265 7670 18284
rect 7618 18244 7670 18253
rect 7618 18210 7624 18244
rect 7624 18210 7658 18244
rect 7658 18210 7670 18244
rect 7618 18201 7670 18210
rect 8391 18573 8443 18625
rect 8391 18509 8443 18561
rect 7616 18040 7668 18045
rect 7616 18006 7624 18040
rect 7624 18006 7658 18040
rect 7658 18006 7668 18040
rect 7616 17993 7668 18006
rect 7616 17968 7668 17981
rect 7616 17934 7624 17968
rect 7624 17934 7658 17968
rect 7658 17934 7668 17968
rect 7616 17929 7668 17934
rect 8231 18189 8283 18241
rect 8231 18125 8283 18177
rect 6847 17278 6899 17330
rect 6915 17278 6967 17330
rect 6983 17278 7035 17330
rect 7051 17278 7103 17330
rect 6847 17211 6899 17263
rect 6915 17211 6967 17263
rect 6983 17211 7035 17263
rect 7051 17211 7103 17263
rect 6847 17144 6899 17196
rect 6915 17144 6967 17196
rect 6983 17175 7006 17196
rect 7006 17175 7035 17196
rect 6983 17144 7035 17175
rect 7051 17175 7058 17196
rect 7058 17175 7092 17196
rect 7092 17175 7103 17196
rect 7051 17144 7103 17175
rect 6847 17077 6899 17129
rect 6915 17077 6967 17129
rect 6983 17077 7035 17129
rect 7051 17077 7103 17129
rect 6847 17010 6899 17062
rect 6915 17010 6967 17062
rect 6983 17010 7035 17062
rect 7051 17010 7103 17062
rect 7524 17053 7576 17076
rect 7524 17024 7530 17053
rect 7530 17024 7564 17053
rect 7564 17024 7576 17053
rect 6847 16942 6899 16994
rect 6915 16942 6967 16994
rect 6983 16942 7035 16994
rect 7051 16942 7103 16994
rect 7524 16960 7576 17012
rect 7618 16685 7624 16715
rect 7624 16685 7658 16715
rect 7658 16685 7670 16715
rect 7618 16663 7670 16685
rect 7618 16644 7670 16651
rect 7618 16610 7624 16644
rect 7624 16610 7658 16644
rect 7658 16610 7670 16644
rect 7618 16599 7670 16610
rect 2654 16170 2706 16222
rect 2654 16106 2706 16158
rect 1648 15664 1700 15716
rect 1648 15600 1700 15652
rect 742 14139 794 14191
rect 806 14139 858 14191
rect 1017 14059 1069 14111
rect 1081 14059 1133 14111
rect 792 13649 844 13701
rect 792 13585 844 13637
rect 931 13445 983 13497
rect 931 13381 983 13433
rect 540 371 592 423
rect 2210 14139 2262 14191
rect 2274 14139 2326 14191
rect 1184 13973 1236 14025
rect 1654 13979 1706 14031
rect 1718 13979 1770 14031
rect 1184 13909 1236 13961
rect 1585 13795 1637 13847
rect 1649 13795 1701 13847
rect 1299 13144 1351 13196
rect 1299 13080 1351 13132
rect 1429 13131 1481 13183
rect 1493 13131 1545 13183
rect 1491 12773 1543 12825
rect 1491 12709 1543 12761
rect 1435 12513 1487 12565
rect 1435 12449 1487 12501
rect 1641 13666 1693 13718
rect 1705 13666 1757 13718
rect 1697 13371 1749 13423
rect 1761 13371 1813 13423
rect 1781 13291 1833 13343
rect 1845 13291 1897 13343
rect 1937 13211 1989 13263
rect 2001 13211 2053 13263
rect 2186 12964 2238 13016
rect 2274 12964 2326 13016
rect 1865 12835 1917 12887
rect 1929 12835 1981 12887
rect 6818 16170 6870 16222
rect 6818 16106 6870 16158
rect 6738 15165 6790 15217
rect 6738 15087 6790 15139
rect 6738 15008 6790 15060
rect 6738 14929 6790 14981
rect 5983 14195 6035 14247
rect 6065 14195 6117 14247
rect 6147 14195 6199 14247
rect 6228 14195 6280 14247
rect 6309 14195 6361 14247
rect 2961 14139 3013 14191
rect 3027 14139 3079 14191
rect 5983 14099 6035 14151
rect 6065 14099 6117 14151
rect 6147 14099 6199 14151
rect 6228 14099 6280 14151
rect 6309 14099 6361 14151
rect 7615 16216 7667 16222
rect 7615 16182 7624 16216
rect 7624 16182 7658 16216
rect 7658 16182 7667 16216
rect 7615 16170 7667 16182
rect 7615 16144 7667 16158
rect 7615 16110 7624 16144
rect 7624 16110 7658 16144
rect 7658 16110 7667 16144
rect 7615 16106 7667 16110
rect 7508 15539 7560 15581
rect 7508 15529 7530 15539
rect 7530 15529 7560 15539
rect 7508 15505 7530 15517
rect 7530 15505 7560 15517
rect 7508 15465 7560 15505
rect 6944 15165 6996 15217
rect 7052 15165 7104 15217
rect 6944 15087 6996 15139
rect 7052 15087 7104 15139
rect 6944 15037 6972 15060
rect 6972 15037 6996 15060
rect 7052 15037 7058 15060
rect 7058 15037 7092 15060
rect 7092 15037 7104 15060
rect 6944 15008 6996 15037
rect 7052 15008 7104 15037
rect 6944 14929 6996 14981
rect 7052 14929 7104 14981
rect 7618 14856 7624 14876
rect 7624 14856 7658 14876
rect 7658 14856 7670 14876
rect 7618 14824 7670 14856
rect 7618 14782 7624 14812
rect 7624 14782 7658 14812
rect 7658 14782 7670 14812
rect 7618 14760 7670 14782
rect 7615 14390 7667 14411
rect 7615 14359 7624 14390
rect 7624 14359 7658 14390
rect 7658 14359 7667 14390
rect 7615 14318 7667 14347
rect 7615 14295 7624 14318
rect 7624 14295 7658 14318
rect 7658 14295 7667 14318
rect 7910 17993 7962 18045
rect 7910 17929 7962 17981
rect 7910 15740 7962 15792
rect 7910 15676 7962 15728
rect 7197 14143 7249 14195
rect 7263 14143 7315 14195
rect 7329 14143 7381 14195
rect 7394 14143 7446 14195
rect 7197 14076 7249 14125
rect 5983 14003 6035 14055
rect 6065 14003 6117 14055
rect 6147 14003 6199 14055
rect 6228 14003 6280 14055
rect 6309 14003 6361 14055
rect 3342 13795 3394 13847
rect 3406 13795 3458 13847
rect 6501 13878 6553 13930
rect 6501 13814 6553 13866
rect 3335 13666 3387 13718
rect 3399 13666 3451 13718
rect 6661 13653 6713 13657
rect 6501 13569 6553 13621
rect 6661 13619 6670 13653
rect 6670 13619 6704 13653
rect 6704 13619 6713 13653
rect 6661 13605 6713 13619
rect 3140 13451 3192 13503
rect 3204 13451 3256 13503
rect 6501 13505 6553 13557
rect 6661 13571 6713 13593
rect 6661 13541 6670 13571
rect 6670 13541 6704 13571
rect 6704 13541 6713 13571
rect 3140 13131 3192 13183
rect 3204 13131 3256 13183
rect 3335 13141 3387 13193
rect 3399 13141 3451 13193
rect 6501 13243 6553 13295
rect 6501 13179 6553 13231
rect 6661 13186 6713 13198
rect 6661 13152 6670 13186
rect 6670 13152 6704 13186
rect 6704 13152 6713 13186
rect 6661 13146 6713 13152
rect 6661 13105 6713 13134
rect 6661 13082 6670 13105
rect 6670 13082 6704 13105
rect 6704 13082 6713 13105
rect 2868 12964 2920 13016
rect 2934 12964 2986 13016
rect 3342 12835 3394 12887
rect 3406 12835 3458 12887
rect 6501 12952 6553 13004
rect 6501 12888 6553 12940
rect 2654 12721 2706 12773
rect 2654 12657 2706 12709
rect 7197 14073 7219 14076
rect 7219 14073 7249 14076
rect 7263 14073 7315 14125
rect 7329 14073 7381 14125
rect 7394 14073 7446 14125
rect 7197 14042 7219 14055
rect 7219 14042 7249 14055
rect 7197 14003 7249 14042
rect 7263 14003 7315 14055
rect 7329 14003 7381 14055
rect 7394 14003 7446 14055
rect 7715 13798 7767 13850
rect 7715 13734 7767 13786
rect 6821 13266 6873 13298
rect 6821 13246 6833 13266
rect 6833 13246 6867 13266
rect 6867 13246 6873 13266
rect 6821 13232 6833 13234
rect 6833 13232 6867 13234
rect 6867 13232 6873 13234
rect 6821 13194 6873 13232
rect 6821 13182 6833 13194
rect 6833 13182 6867 13194
rect 6867 13182 6873 13194
rect 6933 13519 6985 13571
rect 6933 13455 6985 13507
rect 7809 13014 7815 13042
rect 7815 13014 7849 13042
rect 7849 13014 7861 13042
rect 7809 12990 7861 13014
rect 7809 12926 7861 12978
rect 6661 12732 6713 12743
rect 6581 12669 6633 12721
rect 6581 12605 6633 12657
rect 6661 12698 6670 12732
rect 6670 12698 6704 12732
rect 6704 12698 6713 12732
rect 6661 12691 6713 12698
rect 6661 12660 6713 12679
rect 6661 12627 6670 12660
rect 6670 12627 6704 12660
rect 6704 12627 6713 12660
rect 8149 14850 8201 14902
rect 8149 14760 8201 14812
rect 6542 12490 6594 12512
rect 6542 12460 6548 12490
rect 6548 12460 6582 12490
rect 6582 12460 6594 12490
rect 6608 12490 6660 12512
rect 6608 12460 6625 12490
rect 6625 12460 6659 12490
rect 6659 12460 6660 12490
rect 6674 12490 6726 12512
rect 6740 12490 6792 12512
rect 6806 12490 6858 12512
rect 6872 12490 6924 12512
rect 6938 12490 6990 12512
rect 6674 12460 6701 12490
rect 6701 12460 6726 12490
rect 6740 12460 6777 12490
rect 6777 12460 6792 12490
rect 6806 12460 6811 12490
rect 6811 12460 6853 12490
rect 6853 12460 6858 12490
rect 6872 12460 6887 12490
rect 6887 12460 6924 12490
rect 6938 12460 6963 12490
rect 6963 12460 6990 12490
rect 7004 12490 7056 12512
rect 7004 12460 7005 12490
rect 7005 12460 7039 12490
rect 7039 12460 7056 12490
rect 7070 12490 7122 12512
rect 7070 12460 7081 12490
rect 7081 12460 7115 12490
rect 7115 12460 7122 12490
rect 7136 12490 7188 12512
rect 7202 12490 7254 12512
rect 7268 12490 7320 12512
rect 7334 12490 7386 12512
rect 7400 12490 7452 12512
rect 7466 12490 7518 12512
rect 7136 12460 7157 12490
rect 7157 12460 7188 12490
rect 7202 12460 7233 12490
rect 7233 12460 7254 12490
rect 7268 12460 7309 12490
rect 7309 12460 7320 12490
rect 7334 12460 7343 12490
rect 7343 12460 7385 12490
rect 7385 12460 7386 12490
rect 7400 12460 7419 12490
rect 7419 12460 7452 12490
rect 7466 12460 7495 12490
rect 7495 12460 7518 12490
rect 7532 12490 7584 12512
rect 7532 12460 7537 12490
rect 7537 12460 7571 12490
rect 7571 12460 7584 12490
rect 7598 12490 7650 12512
rect 7598 12460 7613 12490
rect 7613 12460 7647 12490
rect 7647 12460 7650 12490
rect 7664 12460 7716 12512
rect 7729 12460 7781 12512
rect 7794 12460 7846 12512
rect 7859 12460 7911 12512
rect 5649 12085 5701 12137
rect 5713 12085 5765 12137
rect 6121 11959 6173 12011
rect 6187 11959 6239 12011
rect 5676 11767 5728 11819
rect 5740 11767 5792 11819
rect 5877 11785 5929 11837
rect 5941 11785 5993 11837
rect 6466 12165 6518 12217
rect 6530 12165 6582 12217
rect 6776 12041 6828 12093
rect 6840 12041 6892 12093
rect 7465 11786 7517 11838
rect 7529 11786 7581 11838
rect 8311 16689 8363 16741
rect 8311 16599 8363 16651
rect 8311 13226 8363 13278
rect 8311 13162 8363 13214
rect 8391 13681 8443 13733
rect 8391 13617 8443 13669
rect 8237 12920 8289 12972
rect 8301 12920 8353 12972
rect 8799 19435 8851 19487
rect 8863 19435 8915 19487
rect 9005 18830 9057 18882
rect 9093 18830 9145 18882
rect 9005 18740 9057 18792
rect 9093 18740 9145 18792
rect 9005 14982 9057 15034
rect 9093 14982 9145 15034
rect 9005 14893 9057 14945
rect 9093 14893 9145 14945
rect 9391 17056 9443 17108
rect 9486 17056 9538 17108
rect 9391 16954 9443 17006
rect 9486 16954 9538 17006
rect 9391 15007 9443 15059
rect 9486 15007 9538 15059
rect 9391 14939 9443 14991
rect 9486 14939 9538 14991
rect 9219 14746 9271 14798
rect 9283 14746 9335 14798
rect 9572 14740 9624 14792
rect 9011 14558 9063 14610
rect 9087 14558 9139 14610
rect 9572 14672 9624 14724
rect 9572 14604 9624 14656
rect 9011 14476 9063 14528
rect 9087 14476 9139 14528
rect 8717 13884 8769 13936
rect 8781 13884 8833 13936
rect 8631 13681 8683 13733
rect 8631 13617 8683 13669
rect 9199 14189 9251 14241
rect 9301 14189 9353 14241
rect 9199 14099 9251 14151
rect 9301 14099 9353 14151
rect 9199 14009 9251 14061
rect 9301 14009 9353 14061
rect 9391 14489 9443 14541
rect 9486 14489 9538 14541
rect 9011 13804 9063 13856
rect 9087 13804 9139 13856
rect 9163 13804 9215 13856
rect 8551 13326 8603 13378
rect 8551 13262 8603 13314
rect 8763 13326 8815 13378
rect 8763 13262 8815 13314
rect 8471 13070 8523 13122
rect 8471 13006 8523 13058
rect 8391 12767 8443 12819
rect 8391 12703 8443 12755
rect 8570 12986 8622 13038
rect 8646 12986 8698 13038
rect 8570 12901 8622 12953
rect 8646 12901 8698 12953
rect 8154 11782 8206 11834
rect 8218 11782 8270 11834
rect 2667 11645 2719 11697
rect 2736 11645 2788 11697
rect 2805 11645 2857 11697
rect 2873 11645 2925 11697
rect 2941 11645 2993 11697
rect 3009 11645 3061 11697
rect 3077 11645 3129 11697
rect 3145 11645 3197 11697
rect 3213 11645 3265 11697
rect 3281 11645 3333 11697
rect 3349 11645 3401 11697
rect 3417 11645 3469 11697
rect 3485 11645 3537 11697
rect 2213 11549 2265 11601
rect 2213 11485 2265 11537
rect 2133 11381 2185 11433
rect 2133 11317 2185 11369
rect 1808 11079 1860 11131
rect 1872 11079 1924 11131
rect 1639 3942 1691 3994
rect 1639 3878 1691 3930
rect 1733 10985 1785 11037
rect 1733 10921 1785 10973
rect 1733 3419 1785 3471
rect 1733 3355 1785 3407
rect 1632 2692 1684 2744
rect 1632 2628 1684 2680
rect 1632 2315 1684 2367
rect 1632 2251 1684 2303
rect 1582 2085 1634 2137
rect 1646 2085 1698 2137
rect 1520 1950 1572 2002
rect 1520 1886 1572 1938
rect 1464 1742 1516 1794
rect 1464 1678 1516 1730
rect 1414 1468 1466 1520
rect 1478 1468 1530 1520
rect 1358 1358 1410 1410
rect 1422 1358 1474 1410
rect 1302 1200 1354 1252
rect 1366 1200 1418 1252
rect 1246 1098 1298 1150
rect 1310 1098 1362 1150
rect 1110 1007 1162 1059
rect 1174 1007 1226 1059
rect 1038 923 1090 975
rect 1102 923 1154 975
rect 963 843 1015 895
rect 1027 843 1079 895
rect 833 659 885 711
rect 897 659 949 711
rect 910 556 962 608
rect 974 556 1026 608
rect 703 476 755 528
rect 767 476 819 528
rect 633 392 685 444
rect 697 392 749 444
rect 540 307 592 359
rect 282 70 334 122
rect 282 6 334 58
rect 1415 70 1467 122
rect 1415 6 1467 58
rect 1813 10300 1865 10352
rect 1813 10236 1865 10288
rect 2667 11559 2719 11611
rect 2736 11559 2788 11611
rect 2805 11559 2857 11611
rect 2873 11559 2925 11611
rect 2941 11559 2993 11611
rect 3009 11559 3061 11611
rect 3077 11559 3129 11611
rect 3145 11559 3197 11611
rect 3213 11559 3265 11611
rect 3281 11559 3333 11611
rect 3349 11559 3401 11611
rect 3417 11559 3469 11611
rect 3485 11559 3537 11611
rect 2350 11381 2402 11433
rect 2350 11317 2402 11369
rect 2707 11225 2759 11277
rect 2707 11133 2759 11185
rect 2627 11065 2679 11117
rect 2627 11001 2679 11053
rect 2213 10505 2265 10557
rect 2213 10441 2265 10493
rect 2320 10515 2372 10567
rect 2384 10515 2436 10567
rect 2133 10195 2185 10247
rect 2133 10131 2185 10183
rect 1983 10035 2035 10087
rect 2047 10035 2099 10087
rect 1893 9625 1945 9677
rect 1893 9561 1945 9613
rect 1893 2692 1945 2744
rect 1893 2628 1945 2680
rect 1973 9494 2025 9546
rect 1973 9430 2025 9482
rect 2053 2609 2105 2661
rect 2053 2545 2105 2597
rect 2213 9949 2265 10001
rect 2213 9885 2265 9937
rect 2213 2693 2265 2745
rect 2293 2825 2345 2877
rect 2293 2761 2345 2813
rect 2373 10401 2425 10453
rect 2373 10337 2425 10389
rect 2373 6260 2425 6312
rect 2373 6196 2425 6248
rect 2627 3499 2679 3551
rect 3155 11118 3207 11127
rect 3155 11084 3188 11118
rect 3188 11084 3207 11118
rect 3155 11075 3207 11084
rect 3219 11118 3271 11127
rect 3219 11084 3226 11118
rect 3226 11084 3260 11118
rect 3260 11084 3271 11118
rect 3219 11075 3271 11084
rect 3610 11118 3662 11127
rect 3610 11084 3633 11118
rect 3633 11084 3662 11118
rect 3610 11075 3662 11084
rect 3674 11118 3726 11127
rect 3674 11084 3680 11118
rect 3680 11084 3714 11118
rect 3714 11084 3726 11118
rect 3674 11075 3726 11084
rect 4069 11118 4121 11127
rect 4069 11084 4099 11118
rect 4099 11084 4121 11118
rect 4069 11075 4121 11084
rect 4133 11118 4185 11127
rect 4133 11084 4147 11118
rect 4147 11084 4181 11118
rect 4181 11084 4185 11118
rect 4133 11075 4185 11084
rect 3087 10995 3139 11047
rect 3151 10995 3203 11047
rect 5012 11172 5064 11181
rect 5012 11138 5018 11172
rect 5018 11138 5052 11172
rect 5052 11138 5064 11172
rect 5012 11129 5064 11138
rect 5076 11172 5128 11181
rect 5076 11138 5090 11172
rect 5090 11138 5124 11172
rect 5124 11138 5128 11172
rect 5076 11129 5128 11138
rect 5996 11172 6048 11184
rect 6070 11172 6122 11184
rect 5996 11138 6013 11172
rect 6013 11138 6048 11172
rect 6070 11138 6101 11172
rect 6101 11138 6122 11172
rect 5996 11132 6048 11138
rect 6070 11132 6122 11138
rect 6143 11172 6195 11184
rect 6143 11138 6155 11172
rect 6155 11138 6189 11172
rect 6189 11138 6195 11172
rect 6143 11132 6195 11138
rect 3411 10915 3463 10967
rect 3480 10915 3532 10967
rect 3707 10915 3759 10967
rect 3772 10915 3824 10967
rect 4033 10915 4085 10967
rect 4097 10915 4149 10967
rect 4342 10915 4394 10967
rect 4406 10915 4458 10967
rect 5721 11044 5773 11096
rect 5842 11078 5894 11096
rect 5842 11044 5883 11078
rect 5883 11044 5894 11078
rect 5963 11044 6015 11096
rect 6083 11044 6135 11096
rect 6203 11078 6255 11096
rect 6203 11044 6229 11078
rect 6229 11044 6255 11078
rect 3121 10812 3173 10841
rect 3121 10789 3127 10812
rect 3127 10789 3161 10812
rect 3161 10789 3173 10812
rect 3186 10812 3238 10841
rect 3186 10789 3202 10812
rect 3202 10789 3236 10812
rect 3236 10789 3238 10812
rect 3251 10812 3303 10841
rect 3316 10812 3368 10841
rect 3381 10812 3433 10841
rect 3446 10812 3498 10841
rect 3511 10812 3563 10841
rect 3576 10812 3628 10841
rect 3251 10789 3276 10812
rect 3276 10789 3303 10812
rect 3316 10789 3350 10812
rect 3350 10789 3368 10812
rect 3381 10789 3384 10812
rect 3384 10789 3424 10812
rect 3424 10789 3433 10812
rect 3446 10789 3458 10812
rect 3458 10789 3498 10812
rect 3511 10789 3532 10812
rect 3532 10789 3563 10812
rect 3576 10789 3606 10812
rect 3606 10789 3628 10812
rect 3641 10812 3693 10841
rect 3641 10789 3646 10812
rect 3646 10789 3680 10812
rect 3680 10789 3693 10812
rect 3706 10812 3758 10841
rect 3706 10789 3720 10812
rect 3720 10789 3754 10812
rect 3754 10789 3758 10812
rect 3771 10812 3823 10841
rect 3836 10812 3888 10841
rect 3901 10812 3953 10841
rect 3966 10812 4018 10841
rect 4031 10812 4083 10841
rect 4096 10812 4148 10841
rect 3771 10789 3794 10812
rect 3794 10789 3823 10812
rect 3836 10789 3868 10812
rect 3868 10789 3888 10812
rect 3901 10789 3902 10812
rect 3902 10789 3942 10812
rect 3942 10789 3953 10812
rect 3966 10789 3976 10812
rect 3976 10789 4016 10812
rect 4016 10789 4018 10812
rect 4031 10789 4050 10812
rect 4050 10789 4083 10812
rect 4096 10789 4124 10812
rect 4124 10789 4148 10812
rect 4160 10812 4212 10841
rect 4160 10789 4164 10812
rect 4164 10789 4198 10812
rect 4198 10789 4212 10812
rect 4224 10812 4276 10841
rect 4224 10789 4238 10812
rect 4238 10789 4272 10812
rect 4272 10789 4276 10812
rect 4288 10812 4340 10841
rect 4352 10812 4404 10841
rect 4416 10812 4468 10841
rect 4480 10812 4532 10841
rect 4544 10812 4596 10841
rect 4288 10789 4312 10812
rect 4312 10789 4340 10812
rect 4352 10789 4386 10812
rect 4386 10789 4404 10812
rect 4416 10789 4420 10812
rect 4420 10789 4460 10812
rect 4460 10789 4468 10812
rect 4480 10789 4494 10812
rect 4494 10789 4532 10812
rect 4544 10789 4568 10812
rect 4568 10789 4596 10812
rect 4608 10789 4660 10841
rect 4672 10789 4724 10841
rect 4736 10789 4788 10841
rect 4800 10789 4852 10841
rect 4864 10789 4916 10841
rect 4928 10789 4980 10841
rect 4992 10789 5044 10841
rect 5056 10789 5108 10841
rect 5120 10789 5172 10841
rect 5184 10789 5236 10841
rect 5248 10789 5300 10841
rect 5312 10789 5364 10841
rect 5376 10789 5428 10841
rect 5440 10789 5492 10841
rect 5504 10789 5556 10841
rect 5568 10789 5620 10841
rect 5632 10789 5684 10841
rect 5696 10832 5748 10841
rect 5760 10832 5812 10841
rect 5696 10798 5727 10832
rect 5727 10798 5748 10832
rect 5760 10798 5761 10832
rect 5761 10798 5812 10832
rect 5696 10789 5748 10798
rect 5760 10789 5812 10798
rect 5824 10789 5876 10841
rect 5888 10789 5940 10841
rect 5952 10789 6004 10841
rect 6016 10831 6068 10841
rect 6016 10797 6039 10831
rect 6039 10797 6068 10831
rect 6016 10789 6068 10797
rect 6080 10789 6132 10841
rect 6144 10789 6196 10841
rect 6208 10789 6260 10841
rect 7069 11023 7078 11057
rect 7078 11023 7112 11057
rect 7112 11023 7121 11057
rect 7069 11005 7121 11023
rect 7069 10985 7121 10993
rect 7069 10951 7078 10985
rect 7078 10951 7112 10985
rect 7112 10951 7121 10985
rect 7069 10941 7121 10951
rect 3121 10719 3173 10771
rect 3186 10719 3238 10771
rect 3251 10719 3303 10771
rect 3316 10719 3368 10771
rect 3381 10719 3433 10771
rect 3446 10719 3498 10771
rect 3511 10719 3563 10771
rect 3576 10719 3628 10771
rect 3641 10719 3693 10771
rect 3706 10719 3758 10771
rect 3771 10719 3823 10771
rect 3836 10719 3888 10771
rect 3901 10719 3953 10771
rect 3966 10719 4018 10771
rect 4031 10719 4083 10771
rect 4096 10719 4148 10771
rect 4160 10719 4212 10771
rect 4224 10719 4276 10771
rect 4288 10719 4340 10771
rect 4352 10719 4404 10771
rect 4416 10719 4468 10771
rect 4480 10719 4532 10771
rect 4544 10719 4596 10771
rect 4608 10719 4660 10771
rect 4672 10719 4724 10771
rect 4736 10719 4788 10771
rect 4800 10719 4852 10771
rect 4864 10719 4916 10771
rect 4928 10719 4980 10771
rect 4992 10719 5044 10771
rect 5056 10719 5108 10771
rect 5120 10719 5172 10771
rect 5184 10719 5236 10771
rect 5248 10719 5300 10771
rect 5312 10719 5364 10771
rect 5376 10719 5428 10771
rect 5440 10719 5492 10771
rect 5504 10719 5556 10771
rect 5568 10719 5620 10771
rect 5632 10719 5684 10771
rect 5696 10719 5748 10771
rect 5760 10719 5812 10771
rect 5824 10719 5876 10771
rect 5888 10719 5940 10771
rect 5952 10719 6004 10771
rect 6016 10719 6068 10771
rect 6080 10719 6132 10771
rect 6144 10719 6196 10771
rect 6208 10719 6260 10771
rect 6711 10807 6717 10835
rect 6717 10807 6751 10835
rect 6751 10807 6763 10835
rect 6711 10783 6763 10807
rect 6811 10783 6863 10835
rect 3121 10649 3173 10701
rect 3186 10649 3238 10701
rect 3251 10649 3303 10701
rect 3316 10649 3368 10701
rect 3381 10649 3433 10701
rect 3446 10649 3498 10701
rect 3511 10649 3563 10701
rect 3576 10649 3628 10701
rect 3641 10649 3693 10701
rect 3706 10649 3758 10701
rect 3771 10649 3823 10701
rect 3836 10649 3888 10701
rect 3901 10649 3953 10701
rect 3966 10649 4018 10701
rect 4031 10649 4083 10701
rect 4096 10649 4148 10701
rect 4160 10649 4212 10701
rect 4224 10649 4276 10701
rect 4288 10649 4340 10701
rect 4352 10649 4404 10701
rect 4416 10649 4468 10701
rect 4480 10649 4532 10701
rect 4544 10649 4596 10701
rect 4608 10649 4660 10701
rect 4672 10649 4724 10701
rect 4736 10649 4788 10701
rect 4800 10649 4852 10701
rect 4864 10649 4916 10701
rect 4928 10649 4980 10701
rect 4992 10680 5023 10701
rect 5023 10680 5044 10701
rect 4992 10649 5044 10680
rect 5056 10680 5062 10701
rect 5062 10680 5096 10701
rect 5096 10680 5108 10701
rect 5056 10649 5108 10680
rect 5120 10680 5135 10701
rect 5135 10680 5169 10701
rect 5169 10680 5172 10701
rect 5120 10649 5172 10680
rect 5184 10680 5208 10701
rect 5208 10680 5236 10701
rect 5248 10680 5281 10701
rect 5281 10680 5300 10701
rect 5312 10680 5315 10701
rect 5315 10680 5354 10701
rect 5354 10680 5364 10701
rect 5376 10680 5388 10701
rect 5388 10680 5427 10701
rect 5427 10680 5428 10701
rect 5440 10680 5461 10701
rect 5461 10680 5492 10701
rect 5504 10680 5534 10701
rect 5534 10680 5556 10701
rect 5184 10649 5236 10680
rect 5248 10649 5300 10680
rect 5312 10649 5364 10680
rect 5376 10649 5428 10680
rect 5440 10649 5492 10680
rect 5504 10649 5556 10680
rect 5568 10680 5572 10701
rect 5572 10680 5606 10701
rect 5606 10680 5620 10701
rect 5568 10649 5620 10680
rect 5632 10680 5644 10701
rect 5644 10680 5678 10701
rect 5678 10680 5684 10701
rect 5632 10649 5684 10680
rect 5696 10680 5716 10701
rect 5716 10680 5748 10701
rect 5760 10680 5788 10701
rect 5788 10680 5812 10701
rect 5824 10680 5860 10701
rect 5860 10680 5876 10701
rect 5888 10680 5894 10701
rect 5894 10680 5932 10701
rect 5932 10680 5940 10701
rect 5952 10680 5966 10701
rect 5966 10680 6004 10701
rect 6016 10680 6038 10701
rect 6038 10680 6068 10701
rect 6080 10680 6110 10701
rect 6110 10680 6132 10701
rect 5696 10649 5748 10680
rect 5760 10649 5812 10680
rect 5824 10649 5876 10680
rect 5888 10649 5940 10680
rect 5952 10649 6004 10680
rect 6016 10649 6068 10680
rect 6080 10649 6132 10680
rect 6144 10680 6148 10701
rect 6148 10680 6182 10701
rect 6182 10680 6196 10701
rect 6144 10649 6196 10680
rect 6208 10680 6220 10701
rect 6220 10680 6254 10701
rect 6254 10680 6260 10701
rect 6208 10649 6260 10680
rect 6711 10768 6763 10771
rect 6711 10734 6717 10768
rect 6717 10734 6751 10768
rect 6751 10734 6763 10768
rect 6711 10719 6763 10734
rect 6811 10719 6863 10771
rect 6711 10695 6763 10707
rect 6711 10661 6717 10695
rect 6717 10661 6751 10695
rect 6751 10661 6763 10695
rect 6711 10655 6763 10661
rect 6811 10660 6863 10707
rect 6811 10655 6836 10660
rect 6836 10655 6863 10660
rect 6314 10469 6366 10521
rect 6390 10469 6442 10521
rect 6466 10469 6518 10521
rect 6314 10397 6366 10449
rect 6390 10397 6442 10449
rect 6466 10397 6518 10449
rect 6314 10325 6366 10377
rect 6390 10325 6442 10377
rect 6466 10325 6518 10377
rect 3735 10251 3787 10303
rect 3799 10251 3851 10303
rect 6314 10253 6366 10305
rect 6390 10253 6442 10305
rect 6466 10253 6518 10305
rect 3261 10125 3313 10177
rect 3327 10125 3379 10177
rect 6314 10181 6366 10233
rect 6390 10181 6442 10233
rect 6466 10181 6518 10233
rect 6314 10109 6366 10161
rect 6390 10109 6442 10161
rect 6466 10109 6518 10161
rect 3511 9955 3563 10007
rect 3575 9955 3627 10007
rect 3708 9933 3760 9985
rect 3772 9933 3824 9985
rect 3099 9799 3151 9851
rect 3166 9799 3218 9851
rect 3233 9799 3285 9851
rect 3300 9799 3352 9851
rect 3367 9799 3419 9851
rect 3434 9799 3486 9851
rect 3500 9799 3552 9851
rect 3566 9799 3618 9851
rect 3632 9799 3684 9851
rect 6744 10515 6751 10521
rect 6751 10515 6796 10521
rect 6744 10477 6796 10515
rect 6744 10469 6751 10477
rect 6751 10469 6796 10477
rect 6812 10469 6864 10521
rect 7128 10493 7180 10545
rect 6744 10443 6751 10449
rect 6751 10443 6796 10449
rect 6744 10405 6796 10443
rect 6744 10397 6751 10405
rect 6751 10397 6796 10405
rect 6812 10397 6864 10449
rect 7128 10429 7180 10481
rect 6744 10371 6751 10377
rect 6751 10371 6796 10377
rect 6744 10333 6796 10371
rect 6744 10325 6751 10333
rect 6751 10325 6796 10333
rect 6812 10348 6864 10377
rect 6812 10325 6836 10348
rect 6836 10325 6864 10348
rect 6744 10299 6751 10305
rect 6751 10299 6796 10305
rect 6744 10261 6796 10299
rect 6744 10253 6751 10261
rect 6751 10253 6796 10261
rect 6812 10253 6864 10305
rect 6744 10227 6751 10233
rect 6751 10227 6796 10233
rect 6744 10189 6796 10227
rect 6744 10181 6751 10189
rect 6751 10181 6796 10189
rect 6812 10181 6864 10233
rect 6744 10155 6751 10161
rect 6751 10155 6796 10161
rect 6744 10117 6796 10155
rect 6744 10109 6751 10117
rect 6751 10109 6796 10117
rect 6812 10109 6864 10161
rect 7323 10263 7375 10315
rect 7222 10203 7274 10239
rect 7222 10187 7228 10203
rect 7228 10187 7262 10203
rect 7262 10187 7274 10203
rect 7323 10199 7375 10251
rect 8465 10942 8517 10994
rect 8465 10878 8517 10930
rect 7222 10169 7228 10175
rect 7228 10169 7262 10175
rect 7262 10169 7274 10175
rect 7222 10125 7274 10169
rect 7222 10123 7228 10125
rect 7228 10123 7262 10125
rect 7262 10123 7274 10125
rect 7715 10107 7767 10159
rect 7791 10107 7843 10159
rect 7715 10017 7767 10069
rect 7791 10017 7843 10069
rect 3099 9719 3151 9771
rect 3166 9719 3218 9771
rect 3233 9719 3285 9771
rect 3300 9719 3352 9771
rect 3367 9719 3419 9771
rect 3434 9719 3486 9771
rect 3500 9719 3552 9771
rect 3566 9719 3618 9771
rect 3632 9719 3684 9771
rect 5837 9609 5889 9661
rect 5901 9609 5953 9661
rect 6034 9591 6086 9643
rect 6098 9591 6150 9643
rect 6282 9417 6334 9469
rect 6348 9417 6400 9469
rect 5810 9291 5862 9343
rect 5874 9291 5926 9343
rect 6571 9668 6623 9720
rect 6571 9604 6623 9656
rect 5810 8541 5862 8593
rect 5874 8541 5926 8593
rect 6282 8415 6334 8467
rect 6348 8415 6400 8467
rect 5837 8223 5889 8275
rect 5901 8223 5953 8275
rect 6034 8241 6086 8293
rect 6098 8241 6150 8293
rect 7228 9648 7280 9660
rect 7228 9614 7262 9648
rect 7262 9614 7280 9648
rect 7228 9608 7280 9614
rect 7292 9608 7344 9660
rect 7040 9256 7092 9262
rect 7040 9222 7057 9256
rect 7057 9222 7092 9256
rect 7040 9210 7092 9222
rect 7112 9256 7164 9262
rect 7112 9222 7122 9256
rect 7122 9222 7156 9256
rect 7156 9222 7164 9256
rect 7112 9210 7164 9222
rect 8576 10581 8628 10633
rect 8640 10581 8692 10633
rect 8764 10583 8816 10635
rect 8846 10583 8898 10635
rect 9391 13525 9443 13577
rect 9486 13525 9538 13577
rect 9391 13449 9443 13501
rect 9486 13449 9538 13501
rect 9391 12992 9443 13044
rect 9486 12992 9538 13044
rect 9391 12896 9443 12948
rect 9486 12896 9538 12948
rect 9342 12349 9394 12401
rect 9406 12349 9458 12401
rect 9232 12269 9284 12321
rect 9296 12269 9348 12321
rect 9182 11869 9234 11921
rect 9246 11869 9298 11921
rect 9011 10339 9063 10391
rect 9087 10339 9139 10391
rect 9011 10273 9063 10325
rect 9087 10273 9139 10325
rect 8862 10193 8914 10245
rect 8926 10193 8978 10245
rect 8298 9417 8350 9469
rect 8362 9417 8414 9469
rect 7721 9210 7773 9262
rect 7785 9210 7837 9262
rect 8208 8875 8260 8927
rect 8208 8811 8260 8863
rect 7903 8719 7955 8771
rect 7903 8655 7955 8707
rect 7078 8293 7112 8294
rect 7112 8293 7130 8294
rect 7078 8242 7130 8293
rect 7143 8242 7195 8294
rect 7833 8242 7885 8294
rect 7897 8242 7949 8294
rect 3148 8100 3200 8152
rect 3213 8100 3265 8152
rect 3278 8100 3330 8152
rect 3343 8100 3395 8152
rect 3408 8100 3460 8152
rect 3473 8100 3525 8152
rect 3538 8100 3590 8152
rect 3603 8100 3655 8152
rect 3668 8100 3720 8152
rect 3733 8100 3785 8152
rect 3798 8100 3850 8152
rect 3863 8100 3915 8152
rect 3928 8100 3980 8152
rect 3993 8100 4045 8152
rect 4058 8100 4110 8152
rect 4123 8100 4175 8152
rect 4188 8100 4240 8152
rect 4253 8100 4305 8152
rect 4318 8100 4370 8152
rect 3148 8036 3200 8088
rect 3213 8036 3265 8088
rect 3278 8036 3330 8088
rect 3343 8036 3395 8088
rect 3408 8036 3460 8088
rect 3473 8036 3525 8088
rect 3538 8036 3590 8088
rect 3603 8036 3655 8088
rect 3668 8036 3720 8088
rect 3733 8036 3785 8088
rect 3798 8036 3850 8088
rect 3863 8036 3915 8088
rect 3928 8036 3980 8088
rect 3993 8036 4045 8088
rect 4058 8036 4110 8088
rect 4123 8036 4175 8088
rect 4188 8036 4240 8088
rect 4253 8036 4305 8088
rect 4318 8036 4370 8088
rect 3148 7972 3200 8024
rect 3213 7972 3265 8024
rect 3278 7972 3330 8024
rect 3343 7972 3395 8024
rect 3408 7972 3460 8024
rect 3473 7972 3525 8024
rect 3538 7972 3590 8024
rect 3603 7972 3655 8024
rect 3668 7972 3720 8024
rect 3733 7972 3785 8024
rect 3798 7972 3850 8024
rect 3863 7972 3915 8024
rect 3928 7972 3980 8024
rect 3993 7972 4045 8024
rect 4058 7972 4110 8024
rect 4123 7972 4175 8024
rect 4188 7972 4240 8024
rect 4253 7972 4305 8024
rect 4318 7972 4370 8024
rect 4383 7972 5459 8152
rect 5552 3872 5604 3924
rect 5616 3872 5668 3924
rect 2707 3785 2759 3837
rect 2707 3708 2759 3760
rect 2707 3631 2759 3683
rect 5427 3791 5479 3843
rect 5491 3791 5543 3843
rect 2707 3554 2759 3606
rect 4369 3591 4421 3600
rect 4369 3557 4402 3591
rect 4402 3557 4421 3591
rect 4369 3548 4421 3557
rect 4433 3591 4485 3600
rect 4433 3557 4440 3591
rect 4440 3557 4474 3591
rect 4474 3557 4485 3591
rect 4433 3548 4485 3557
rect 4833 3591 4885 3600
rect 4833 3557 4866 3591
rect 4866 3557 4885 3591
rect 4833 3548 4885 3557
rect 4897 3591 4949 3600
rect 4897 3557 4907 3591
rect 4907 3557 4941 3591
rect 4941 3557 4949 3591
rect 4897 3548 4949 3557
rect 5407 3591 5459 3600
rect 5407 3557 5412 3591
rect 5412 3557 5446 3591
rect 5446 3557 5459 3591
rect 5407 3548 5459 3557
rect 5491 3591 5543 3600
rect 5491 3557 5503 3591
rect 5503 3557 5537 3591
rect 5537 3557 5543 3591
rect 5491 3548 5543 3557
rect 2627 3435 2679 3487
rect 4306 3429 4358 3481
rect 4370 3429 4422 3481
rect 4630 3349 4682 3401
rect 4694 3349 4746 3401
rect 4926 3349 4978 3401
rect 4990 3349 5042 3401
rect 5251 3349 5303 3401
rect 5315 3349 5367 3401
rect 5552 3349 5604 3401
rect 5616 3349 5668 3401
rect 4499 3263 4551 3315
rect 4499 3199 4551 3251
rect 4811 3263 4863 3315
rect 4811 3199 4863 3251
rect 5123 3263 5175 3315
rect 5123 3199 5175 3251
rect 5435 3263 5487 3315
rect 5435 3199 5487 3251
rect 5747 3263 5799 3315
rect 5747 3199 5799 3251
rect 5629 3084 5681 3136
rect 5696 3084 5748 3136
rect 5763 3084 5815 3136
rect 5830 3084 5882 3136
rect 5897 3084 5949 3136
rect 5964 3084 6016 3136
rect 6031 3084 6083 3136
rect 6098 3084 6150 3136
rect 6165 3084 6217 3136
rect 6232 3084 6284 3136
rect 6299 3084 6351 3136
rect 6366 3084 6418 3136
rect 6433 3084 6485 3136
rect 6499 3084 6551 3136
rect 6565 3084 6617 3136
rect 5629 2996 5681 3048
rect 5696 2996 5748 3048
rect 5763 2996 5815 3048
rect 5830 2996 5882 3048
rect 5897 2996 5949 3048
rect 5964 2996 6016 3048
rect 6031 2996 6083 3048
rect 6098 2996 6150 3048
rect 6165 2996 6217 3048
rect 6232 2996 6284 3048
rect 6299 2996 6351 3048
rect 6366 2996 6418 3048
rect 6433 2996 6485 3048
rect 6499 2996 6551 3048
rect 6565 2996 6617 3048
rect 2373 2876 2425 2928
rect 2373 2812 2425 2864
rect 3610 2806 3662 2858
rect 3674 2806 3726 2858
rect 2213 2629 2265 2681
rect 3712 2703 3764 2755
rect 3776 2703 3828 2755
rect 3232 2623 3284 2675
rect 3296 2623 3348 2675
rect 2923 2539 2975 2591
rect 2987 2539 3039 2591
rect 4264 2620 4316 2672
rect 4264 2556 4316 2608
rect 4920 2809 4972 2861
rect 4984 2809 5036 2861
rect 5982 2809 6034 2861
rect 6046 2809 6098 2861
rect 4577 2685 4629 2737
rect 5880 2706 5932 2758
rect 5944 2706 5996 2758
rect 4577 2621 4629 2673
rect 6360 2626 6412 2678
rect 6424 2626 6476 2678
rect 6669 2542 6721 2594
rect 6733 2542 6785 2594
rect 1973 2395 2025 2447
rect 2063 2435 2115 2487
rect 2127 2435 2179 2487
rect 2987 2448 3039 2500
rect 3053 2448 3105 2500
rect 4297 2451 4349 2503
rect 4363 2451 4415 2503
rect 4969 2441 5021 2493
rect 6603 2451 6655 2503
rect 6669 2451 6721 2503
rect 1973 2331 2025 2383
rect 4969 2377 5021 2429
rect 4122 2325 4174 2377
rect 4186 2325 4238 2377
rect 6950 7886 7002 7937
rect 7046 7886 7098 7937
rect 6950 7885 6972 7886
rect 6972 7885 7002 7886
rect 7046 7885 7052 7886
rect 7052 7885 7086 7886
rect 7086 7885 7098 7886
rect 6950 7789 7002 7841
rect 7046 7789 7098 7841
rect 7500 7287 7552 7339
rect 7500 7197 7552 7249
rect 7618 7029 7624 7039
rect 7624 7029 7658 7039
rect 7658 7029 7670 7039
rect 7618 6989 7670 7029
rect 7618 6987 7624 6989
rect 7624 6987 7658 6989
rect 7658 6987 7670 6989
rect 7618 6955 7624 6975
rect 7624 6955 7658 6975
rect 7658 6955 7670 6975
rect 7618 6923 7670 6955
rect 7615 6233 7624 6262
rect 7624 6233 7658 6262
rect 7658 6233 7667 6262
rect 7615 6210 7667 6233
rect 7615 6195 7667 6198
rect 7615 6161 7624 6195
rect 7624 6161 7658 6195
rect 7658 6161 7667 6195
rect 7615 6146 7667 6161
rect 6944 6075 6996 6127
rect 7052 6075 7104 6127
rect 6944 6026 6972 6057
rect 6972 6026 6996 6057
rect 7052 6026 7086 6057
rect 7086 6026 7104 6057
rect 6944 6005 6996 6026
rect 7052 6005 7104 6026
rect 6944 5935 6996 5987
rect 7052 5935 7104 5987
rect 6944 5865 6996 5917
rect 7052 5865 7104 5917
rect 6944 5795 6996 5847
rect 7052 5795 7104 5847
rect 7704 5865 7756 5902
rect 7704 5850 7716 5865
rect 7716 5850 7750 5865
rect 7750 5850 7756 5865
rect 7704 5831 7716 5835
rect 7716 5831 7750 5835
rect 7750 5831 7756 5835
rect 7704 5793 7756 5831
rect 7704 5783 7716 5793
rect 7716 5783 7750 5793
rect 7750 5783 7756 5793
rect 6944 5748 6996 5777
rect 7052 5748 7104 5777
rect 7704 5759 7716 5768
rect 7716 5759 7750 5768
rect 7750 5759 7756 5768
rect 6944 5725 6972 5748
rect 6972 5725 6996 5748
rect 7052 5725 7058 5748
rect 7058 5725 7092 5748
rect 7092 5725 7104 5748
rect 7704 5721 7756 5759
rect 7704 5716 7716 5721
rect 7716 5716 7750 5721
rect 7750 5716 7756 5721
rect 6944 5654 6996 5706
rect 7052 5654 7104 5706
rect 7704 5687 7716 5700
rect 7716 5687 7750 5700
rect 7750 5687 7756 5700
rect 6944 5583 6996 5635
rect 7052 5583 7104 5635
rect 6944 5512 6996 5564
rect 7052 5512 7104 5564
rect 7524 5188 7576 5240
rect 7524 5098 7576 5150
rect 7704 5649 7756 5687
rect 7704 5648 7716 5649
rect 7716 5648 7750 5649
rect 7750 5648 7756 5649
rect 7704 5615 7716 5632
rect 7716 5615 7750 5632
rect 7750 5615 7756 5632
rect 7704 5580 7756 5615
rect 7704 5543 7716 5564
rect 7716 5543 7750 5564
rect 7750 5543 7756 5564
rect 7704 5512 7756 5543
rect 7618 4979 7624 4990
rect 7624 4979 7658 4990
rect 7658 4979 7670 4990
rect 7618 4940 7670 4979
rect 7618 4938 7624 4940
rect 7624 4938 7658 4940
rect 7658 4938 7670 4940
rect 7618 4906 7624 4926
rect 7624 4906 7658 4926
rect 7658 4906 7670 4926
rect 7618 4874 7670 4906
rect 7615 4439 7667 4448
rect 7615 4405 7624 4439
rect 7624 4405 7658 4439
rect 7658 4405 7667 4439
rect 7615 4396 7667 4405
rect 7615 4367 7667 4384
rect 7615 4333 7624 4367
rect 7624 4333 7658 4367
rect 7658 4333 7667 4367
rect 7615 4332 7667 4333
rect 6944 4002 6996 4054
rect 7052 4002 7104 4054
rect 6944 3935 6996 3987
rect 7052 3935 7104 3987
rect 6944 3888 6972 3920
rect 6972 3888 6996 3920
rect 7052 3888 7058 3920
rect 7058 3888 7092 3920
rect 7092 3888 7104 3920
rect 6944 3868 6996 3888
rect 7052 3868 7104 3888
rect 6944 3801 6996 3853
rect 7052 3801 7104 3853
rect 7615 3850 7667 3871
rect 6944 3734 6996 3786
rect 7052 3734 7104 3786
rect 7615 3819 7624 3850
rect 7624 3819 7658 3850
rect 7658 3819 7667 3850
rect 7615 3775 7667 3807
rect 7615 3755 7624 3775
rect 7624 3755 7658 3775
rect 7658 3755 7667 3775
rect 6944 3666 6996 3718
rect 7052 3666 7104 3718
rect 6944 3298 6996 3315
rect 7052 3298 7104 3315
rect 6944 3264 6972 3298
rect 6972 3264 6996 3298
rect 7052 3264 7058 3298
rect 7058 3264 7092 3298
rect 7092 3264 7104 3298
rect 6944 3263 6996 3264
rect 7052 3263 7104 3264
rect 6944 3192 6996 3244
rect 7052 3192 7104 3244
rect 7524 3220 7576 3272
rect 6944 3120 6996 3172
rect 7052 3120 7104 3172
rect 7524 3156 7576 3208
rect 6944 3048 6996 3100
rect 7052 3048 7104 3100
rect 6944 2986 6996 3028
rect 7052 2986 7104 3028
rect 6944 2976 6972 2986
rect 6972 2976 6996 2986
rect 7052 2976 7058 2986
rect 7058 2976 7092 2986
rect 7092 2976 7104 2986
rect 7823 3635 7875 3687
rect 7823 3554 7875 3606
rect 7903 2879 7955 2931
rect 7903 2815 7955 2867
rect 8702 9167 8754 9219
rect 8766 9167 8818 9219
rect 8368 8510 8420 8562
rect 8368 8446 8420 8498
rect 8208 2828 8260 2880
rect 8208 2764 8260 2816
rect 8288 8228 8340 8280
rect 8288 8164 8340 8216
rect 8288 2696 8340 2748
rect 8288 2632 8340 2684
rect 8528 8590 8580 8642
rect 8528 8526 8580 8578
rect 8448 8354 8500 8406
rect 8448 8290 8500 8342
rect 8448 2664 8500 2716
rect 8448 2600 8500 2652
rect 8374 2451 8426 2503
rect 8438 2451 8490 2503
rect 3805 2245 3857 2297
rect 3869 2245 3921 2297
rect 6780 2291 6832 2343
rect 6844 2291 6896 2343
rect 2093 2165 2145 2217
rect 2157 2165 2209 2217
rect 3777 2165 3829 2217
rect 3841 2165 3893 2217
rect 1652 70 1704 122
rect 1652 6 1704 58
rect 1909 70 1961 122
rect 1909 6 1961 58
rect 3201 1984 3253 2036
rect 3267 1984 3319 2036
rect 3917 1984 3969 2036
rect 3994 1984 4046 2036
rect 3708 1890 3760 1942
rect 2961 1800 3013 1852
rect 3025 1800 3077 1852
rect 3708 1806 3760 1858
rect 4908 1890 4960 1942
rect 8374 2131 8426 2183
rect 8438 2131 8490 2183
rect 5833 1980 5885 2032
rect 5910 1980 5962 2032
rect 6549 1984 6601 2036
rect 6626 1984 6678 2036
rect 8458 1984 8510 2036
rect 8522 1984 8574 2036
rect 8608 8169 8660 8221
rect 8608 8105 8660 8157
rect 4908 1806 4960 1858
rect 5410 1866 5462 1918
rect 5410 1802 5462 1854
rect 5621 1890 5673 1942
rect 5621 1806 5673 1858
rect 6340 1890 6392 1942
rect 6340 1806 6392 1858
rect 8538 1880 8590 1932
rect 8602 1880 8654 1932
rect 8688 8068 8740 8120
rect 8688 8004 8740 8056
rect 8772 4472 8824 4524
rect 8772 4408 8824 4460
rect 8772 3049 8824 3101
rect 8772 2985 8824 3037
rect 8852 9097 8904 9149
rect 8852 9033 8904 9085
rect 8932 4958 8984 5010
rect 8932 4894 8984 4946
rect 9012 9904 9064 9956
rect 9012 9840 9064 9892
rect 8805 2441 8857 2493
rect 8805 2377 8857 2429
rect 8688 1794 8740 1846
rect 6479 1694 6531 1746
rect 6580 1694 6632 1746
rect 6681 1694 6733 1746
rect 6782 1694 6834 1746
rect 6882 1694 6934 1746
rect 6982 1694 7034 1746
rect 7082 1694 7134 1746
rect 7182 1694 7234 1746
rect 7282 1694 7334 1746
rect 7382 1694 7434 1746
rect 7482 1694 7534 1746
rect 7582 1694 7634 1746
rect 7682 1694 7734 1746
rect 7782 1694 7834 1746
rect 8688 1730 8740 1782
rect 8794 1984 8846 2036
rect 8858 1984 8910 2036
rect 6479 1620 6531 1672
rect 6580 1620 6632 1672
rect 6681 1620 6733 1672
rect 6782 1620 6834 1672
rect 6882 1620 6934 1672
rect 6982 1620 7034 1672
rect 7082 1620 7134 1672
rect 7182 1620 7234 1672
rect 7282 1620 7334 1672
rect 7382 1620 7434 1672
rect 7482 1620 7534 1672
rect 7582 1620 7634 1672
rect 7682 1620 7734 1672
rect 7782 1620 7834 1672
rect 2961 1468 3013 1520
rect 3025 1468 3077 1520
rect 3527 1464 3579 1516
rect 3595 1464 3647 1516
rect 3663 1464 3715 1516
rect 3731 1464 3783 1516
rect 3799 1464 3851 1516
rect 3867 1464 3919 1516
rect 3934 1464 3986 1516
rect 4001 1464 4053 1516
rect 4068 1464 4120 1516
rect 3527 1400 3579 1452
rect 3595 1400 3647 1452
rect 3663 1400 3715 1452
rect 3731 1400 3783 1452
rect 3799 1400 3851 1452
rect 3867 1400 3919 1452
rect 3934 1400 3986 1452
rect 4001 1400 4053 1452
rect 4068 1400 4120 1452
rect 3201 1285 3253 1337
rect 3267 1285 3319 1337
rect 3527 1336 3579 1388
rect 3595 1336 3647 1388
rect 3663 1336 3715 1388
rect 3731 1336 3783 1388
rect 3799 1336 3851 1388
rect 3867 1336 3919 1388
rect 3934 1336 3986 1388
rect 4001 1336 4053 1388
rect 4068 1336 4120 1388
rect 3527 1272 3579 1324
rect 3595 1272 3647 1324
rect 3663 1272 3715 1324
rect 3731 1272 3783 1324
rect 3799 1272 3851 1324
rect 3867 1272 3919 1324
rect 3934 1272 3986 1324
rect 4001 1272 4053 1324
rect 4068 1272 4120 1324
rect 3527 1208 3579 1260
rect 3595 1208 3647 1260
rect 3663 1208 3715 1260
rect 3731 1208 3783 1260
rect 3799 1208 3851 1260
rect 3867 1208 3919 1260
rect 3934 1208 3986 1260
rect 4001 1208 4053 1260
rect 4068 1208 4120 1260
rect 5829 996 5881 1048
rect 5896 996 5948 1048
rect 5963 996 6015 1048
rect 6030 996 6082 1048
rect 6097 996 6149 1048
rect 6164 996 6216 1048
rect 6231 996 6283 1048
rect 6298 996 6350 1048
rect 6365 996 6417 1048
rect 6432 996 6484 1048
rect 6499 996 6551 1048
rect 6565 996 6617 1048
rect 8388 1012 8440 1064
rect 8388 948 8440 1000
rect 3610 656 3662 708
rect 3674 656 3726 708
rect 4264 649 4316 701
rect 3712 556 3764 608
rect 3776 556 3828 608
rect 4264 585 4316 637
rect 3232 476 3284 528
rect 3296 476 3348 528
rect 2923 392 2975 444
rect 2987 392 3039 444
rect 4576 649 4628 701
rect 5018 662 5070 714
rect 5082 662 5134 714
rect 5982 659 6034 711
rect 6046 659 6098 711
rect 4576 574 4628 626
rect 5022 559 5074 611
rect 5086 559 5138 611
rect 5880 556 5932 608
rect 5944 556 5996 608
rect 6360 476 6412 528
rect 6424 476 6476 528
rect 6669 392 6721 444
rect 6733 392 6785 444
rect 2987 301 3039 353
rect 3053 301 3105 353
rect 4297 304 4349 356
rect 4363 304 4415 356
rect 6603 301 6655 353
rect 6669 301 6721 353
rect 2163 70 2215 122
rect 2163 6 2215 58
rect 2496 106 2548 158
rect 2496 6 2548 58
rect 6843 70 6895 122
rect 6843 6 6895 58
rect 9092 9580 9144 9632
rect 9092 9516 9144 9568
rect 9092 2281 9144 2333
rect 9092 2217 9144 2269
rect 9172 9306 9224 9358
rect 9172 9242 9224 9294
rect 9050 1534 9102 1586
rect 9114 1534 9166 1586
rect 8874 1374 8926 1426
rect 8938 1374 8990 1426
rect 9172 1028 9224 1080
rect 9172 964 9224 1016
rect 8794 824 8846 876
rect 8858 824 8910 876
rect 9332 729 9384 781
rect 9332 665 9384 717
rect 9890 14414 9942 14466
rect 9890 14350 9942 14402
rect 9732 14189 9784 14241
rect 9808 14189 9860 14241
rect 9732 14099 9784 14151
rect 9808 14099 9860 14151
rect 9732 14009 9784 14061
rect 9808 14009 9860 14061
rect 9738 12460 9790 12512
rect 9804 12460 9856 12512
rect 10710 14203 10762 14255
rect 10776 14203 10828 14255
rect 10710 14106 10762 14158
rect 10776 14106 10828 14158
rect 10710 14009 10762 14061
rect 10776 14009 10828 14061
rect 9890 12314 9942 12366
rect 9572 12029 9624 12081
rect 9572 11965 9624 12017
rect 9652 12210 9704 12262
rect 9890 12250 9942 12302
rect 9652 12146 9704 12198
rect 9572 11536 9624 11588
rect 9572 11472 9624 11524
rect 9492 9824 9544 9876
rect 9492 9760 9544 9812
rect 9492 1524 9544 1576
rect 9492 1460 9544 1512
rect 9502 1134 9554 1186
rect 9566 1134 9618 1186
rect 9652 1364 9704 1416
rect 9652 1300 9704 1352
rect 9572 1028 9624 1080
rect 9572 964 9624 1016
rect 9412 626 9464 678
rect 9412 562 9464 614
rect 9492 894 9544 946
rect 9492 830 9544 882
rect 9258 392 9310 444
rect 9322 392 9374 444
rect 8176 70 8228 122
rect 8176 6 8228 58
rect 8469 70 8521 122
rect 8469 6 8521 58
rect 8701 70 8753 122
rect 8701 6 8753 58
rect 8918 70 8970 122
rect 8918 6 8970 58
rect 9232 70 9284 122
rect 9232 6 9284 58
rect 9890 11842 9942 11894
rect 9890 11760 9942 11812
rect 9970 11692 10022 11744
rect 9970 11628 10022 11680
rect 9970 1284 10022 1336
rect 9970 1220 10022 1272
rect 9890 546 9942 598
rect 9890 482 9942 534
rect 9572 70 9624 122
rect 9572 6 9624 58
rect 9784 70 9836 122
rect 9784 6 9836 58
rect 10031 70 10083 122
rect 10031 6 10083 58
rect 10263 70 10315 122
rect 10263 6 10315 58
<< metal2 >>
rect 282 38979 3543 38988
rect 282 38946 2714 38979
rect 282 38890 291 38946
rect 347 38890 374 38946
rect 430 38890 456 38946
rect 512 38890 538 38946
rect 594 38890 620 38946
rect 676 38890 702 38946
rect 758 38890 784 38946
rect 840 38890 866 38946
rect 922 38890 948 38946
rect 1004 38890 1030 38946
rect 1086 38890 1112 38946
rect 1168 38890 1194 38946
rect 1250 38890 1276 38946
rect 1332 38890 1358 38946
rect 1414 38923 2714 38946
rect 2770 38923 2794 38979
rect 2850 38923 2874 38979
rect 2930 38923 2954 38979
rect 3010 38923 3034 38979
rect 3090 38923 3114 38979
rect 3170 38923 3194 38979
rect 3250 38923 3274 38979
rect 3330 38923 3354 38979
rect 3410 38923 3434 38979
rect 3490 38923 3543 38979
rect 1414 38895 3543 38923
rect 1414 38890 2714 38895
rect 282 38860 2714 38890
rect 282 38804 291 38860
rect 347 38804 374 38860
rect 430 38804 456 38860
rect 512 38804 538 38860
rect 594 38804 620 38860
rect 676 38804 702 38860
rect 758 38804 784 38860
rect 840 38804 866 38860
rect 922 38804 948 38860
rect 1004 38804 1030 38860
rect 1086 38804 1112 38860
rect 1168 38804 1194 38860
rect 1250 38804 1276 38860
rect 1332 38804 1358 38860
rect 1414 38839 2714 38860
rect 2770 38839 2794 38895
rect 2850 38839 2874 38895
rect 2930 38839 2954 38895
rect 3010 38839 3034 38895
rect 3090 38839 3114 38895
rect 3170 38839 3194 38895
rect 3250 38839 3274 38895
rect 3330 38839 3354 38895
rect 3410 38839 3434 38895
rect 3490 38839 3543 38895
rect 1414 38811 3543 38839
rect 1414 38804 2714 38811
rect 282 38774 2714 38804
rect 282 38718 291 38774
rect 347 38718 374 38774
rect 430 38718 456 38774
rect 512 38718 538 38774
rect 594 38718 620 38774
rect 676 38718 702 38774
rect 758 38718 784 38774
rect 840 38718 866 38774
rect 922 38718 948 38774
rect 1004 38718 1030 38774
rect 1086 38718 1112 38774
rect 1168 38718 1194 38774
rect 1250 38718 1276 38774
rect 1332 38718 1358 38774
rect 1414 38755 2714 38774
rect 2770 38755 2794 38811
rect 2850 38755 2874 38811
rect 2930 38755 2954 38811
rect 3010 38755 3034 38811
rect 3090 38755 3114 38811
rect 3170 38755 3194 38811
rect 3250 38755 3274 38811
rect 3330 38755 3354 38811
rect 3410 38755 3434 38811
rect 3490 38755 3543 38811
rect 1414 38727 3543 38755
rect 1414 38718 2714 38727
rect 282 38688 2714 38718
rect 282 38632 291 38688
rect 347 38632 374 38688
rect 430 38632 456 38688
rect 512 38632 538 38688
rect 594 38632 620 38688
rect 676 38632 702 38688
rect 758 38632 784 38688
rect 840 38632 866 38688
rect 922 38632 948 38688
rect 1004 38632 1030 38688
rect 1086 38632 1112 38688
rect 1168 38632 1194 38688
rect 1250 38632 1276 38688
rect 1332 38632 1358 38688
rect 1414 38671 2714 38688
rect 2770 38671 2794 38727
rect 2850 38671 2874 38727
rect 2930 38671 2954 38727
rect 3010 38671 3034 38727
rect 3090 38671 3114 38727
rect 3170 38671 3194 38727
rect 3250 38671 3274 38727
rect 3330 38671 3354 38727
rect 3410 38671 3434 38727
rect 3490 38671 3543 38727
rect 1414 38643 3543 38671
rect 1414 38632 2714 38643
rect 282 38602 2714 38632
rect 282 38546 291 38602
rect 347 38546 374 38602
rect 430 38546 456 38602
rect 512 38546 538 38602
rect 594 38546 620 38602
rect 676 38546 702 38602
rect 758 38546 784 38602
rect 840 38546 866 38602
rect 922 38546 948 38602
rect 1004 38546 1030 38602
rect 1086 38546 1112 38602
rect 1168 38546 1194 38602
rect 1250 38546 1276 38602
rect 1332 38546 1358 38602
rect 1414 38587 2714 38602
rect 2770 38587 2794 38643
rect 2850 38587 2874 38643
rect 2930 38587 2954 38643
rect 3010 38587 3034 38643
rect 3090 38587 3114 38643
rect 3170 38587 3194 38643
rect 3250 38587 3274 38643
rect 3330 38587 3354 38643
rect 3410 38587 3434 38643
rect 3490 38587 3543 38643
rect 1414 38559 3543 38587
rect 1414 38546 2714 38559
rect 282 38516 2714 38546
rect 282 38460 291 38516
rect 347 38460 374 38516
rect 430 38460 456 38516
rect 512 38460 538 38516
rect 594 38460 620 38516
rect 676 38460 702 38516
rect 758 38460 784 38516
rect 840 38460 866 38516
rect 922 38460 948 38516
rect 1004 38460 1030 38516
rect 1086 38460 1112 38516
rect 1168 38460 1194 38516
rect 1250 38460 1276 38516
rect 1332 38460 1358 38516
rect 1414 38503 2714 38516
rect 2770 38503 2794 38559
rect 2850 38503 2874 38559
rect 2930 38503 2954 38559
rect 3010 38503 3034 38559
rect 3090 38503 3114 38559
rect 3170 38503 3194 38559
rect 3250 38503 3274 38559
rect 3330 38503 3354 38559
rect 3410 38503 3434 38559
rect 3490 38503 3543 38559
rect 1414 38475 3543 38503
rect 1414 38460 2714 38475
rect 282 38430 2714 38460
rect 282 38374 291 38430
rect 347 38374 374 38430
rect 430 38374 456 38430
rect 512 38374 538 38430
rect 594 38374 620 38430
rect 676 38374 702 38430
rect 758 38374 784 38430
rect 840 38374 866 38430
rect 922 38374 948 38430
rect 1004 38374 1030 38430
rect 1086 38374 1112 38430
rect 1168 38374 1194 38430
rect 1250 38374 1276 38430
rect 1332 38374 1358 38430
rect 1414 38419 2714 38430
rect 2770 38419 2794 38475
rect 2850 38419 2874 38475
rect 2930 38419 2954 38475
rect 3010 38419 3034 38475
rect 3090 38419 3114 38475
rect 3170 38419 3194 38475
rect 3250 38419 3274 38475
rect 3330 38419 3354 38475
rect 3410 38419 3434 38475
rect 3490 38419 3543 38475
rect 1414 38391 3543 38419
rect 1414 38374 2714 38391
rect 282 38344 2714 38374
rect 282 38288 291 38344
rect 347 38288 374 38344
rect 430 38288 456 38344
rect 512 38288 538 38344
rect 594 38288 620 38344
rect 676 38288 702 38344
rect 758 38288 784 38344
rect 840 38288 866 38344
rect 922 38288 948 38344
rect 1004 38288 1030 38344
rect 1086 38288 1112 38344
rect 1168 38288 1194 38344
rect 1250 38288 1276 38344
rect 1332 38288 1358 38344
rect 1414 38335 2714 38344
rect 2770 38335 2794 38391
rect 2850 38335 2874 38391
rect 2930 38335 2954 38391
rect 3010 38335 3034 38391
rect 3090 38335 3114 38391
rect 3170 38335 3194 38391
rect 3250 38335 3274 38391
rect 3330 38335 3354 38391
rect 3410 38335 3434 38391
rect 3490 38335 3543 38391
rect 1414 38307 3543 38335
rect 1414 38288 2714 38307
rect 282 38258 2714 38288
rect 282 38202 291 38258
rect 347 38202 374 38258
rect 430 38202 456 38258
rect 512 38202 538 38258
rect 594 38202 620 38258
rect 676 38202 702 38258
rect 758 38202 784 38258
rect 840 38202 866 38258
rect 922 38202 948 38258
rect 1004 38202 1030 38258
rect 1086 38202 1112 38258
rect 1168 38202 1194 38258
rect 1250 38202 1276 38258
rect 1332 38202 1358 38258
rect 1414 38251 2714 38258
rect 2770 38251 2794 38307
rect 2850 38251 2874 38307
rect 2930 38251 2954 38307
rect 3010 38251 3034 38307
rect 3090 38251 3114 38307
rect 3170 38251 3194 38307
rect 3250 38251 3274 38307
rect 3330 38251 3354 38307
rect 3410 38251 3434 38307
rect 3490 38251 3543 38307
rect 1414 38223 3543 38251
rect 1414 38202 2714 38223
rect 282 38172 2714 38202
rect 282 38116 291 38172
rect 347 38116 374 38172
rect 430 38116 456 38172
rect 512 38116 538 38172
rect 594 38116 620 38172
rect 676 38116 702 38172
rect 758 38116 784 38172
rect 840 38116 866 38172
rect 922 38116 948 38172
rect 1004 38116 1030 38172
rect 1086 38116 1112 38172
rect 1168 38116 1194 38172
rect 1250 38116 1276 38172
rect 1332 38116 1358 38172
rect 1414 38167 2714 38172
rect 2770 38167 2794 38223
rect 2850 38167 2874 38223
rect 2930 38167 2954 38223
rect 3010 38167 3034 38223
rect 3090 38167 3114 38223
rect 3170 38167 3194 38223
rect 3250 38167 3274 38223
rect 3330 38167 3354 38223
rect 3410 38167 3434 38223
rect 3490 38167 3543 38223
rect 1414 38138 3543 38167
rect 1414 38116 2714 38138
rect 282 38086 2714 38116
rect 282 38030 291 38086
rect 347 38030 374 38086
rect 430 38030 456 38086
rect 512 38030 538 38086
rect 594 38030 620 38086
rect 676 38030 702 38086
rect 758 38030 784 38086
rect 840 38030 866 38086
rect 922 38030 948 38086
rect 1004 38030 1030 38086
rect 1086 38030 1112 38086
rect 1168 38030 1194 38086
rect 1250 38030 1276 38086
rect 1332 38030 1358 38086
rect 1414 38082 2714 38086
rect 2770 38082 2794 38138
rect 2850 38082 2874 38138
rect 2930 38082 2954 38138
rect 3010 38082 3034 38138
rect 3090 38082 3114 38138
rect 3170 38082 3194 38138
rect 3250 38082 3274 38138
rect 3330 38082 3354 38138
rect 3410 38082 3434 38138
rect 3490 38082 3543 38138
rect 1414 38053 3543 38082
rect 1414 38030 2714 38053
rect 282 37997 2714 38030
rect 2770 37997 2794 38053
rect 2850 37997 2874 38053
rect 2930 37997 2954 38053
rect 3010 37997 3034 38053
rect 3090 37997 3114 38053
rect 3170 37997 3194 38053
rect 3250 37997 3274 38053
rect 3330 37997 3354 38053
rect 3410 37997 3434 38053
rect 3490 37997 3543 38053
rect 282 37988 3543 37997
tri 5663 36372 6673 37382 sw
rect 4663 36330 10022 36372
rect 4663 36274 8035 36330
rect 8091 36274 8116 36330
rect 8172 36274 8197 36330
rect 8253 36274 8277 36330
rect 8333 36274 8357 36330
rect 8413 36274 8437 36330
rect 8493 36274 8517 36330
rect 8573 36274 8597 36330
rect 8653 36274 8677 36330
rect 8733 36274 8757 36330
rect 8813 36274 8837 36330
rect 8893 36274 8917 36330
rect 8973 36274 8997 36330
rect 9053 36274 9077 36330
rect 9133 36274 9157 36330
rect 9213 36274 9237 36330
rect 9293 36274 9317 36330
rect 9373 36274 9397 36330
rect 9453 36274 9477 36330
rect 9533 36274 9557 36330
rect 9613 36274 9637 36330
rect 9693 36274 9717 36330
rect 9773 36274 9797 36330
rect 9853 36274 9877 36330
rect 9933 36274 9957 36330
rect 10013 36274 10022 36330
rect 4663 36244 10022 36274
rect 4663 36188 8035 36244
rect 8091 36188 8116 36244
rect 8172 36188 8197 36244
rect 8253 36188 8277 36244
rect 8333 36188 8357 36244
rect 8413 36188 8437 36244
rect 8493 36188 8517 36244
rect 8573 36188 8597 36244
rect 8653 36188 8677 36244
rect 8733 36188 8757 36244
rect 8813 36188 8837 36244
rect 8893 36188 8917 36244
rect 8973 36188 8997 36244
rect 9053 36188 9077 36244
rect 9133 36188 9157 36244
rect 9213 36188 9237 36244
rect 9293 36188 9317 36244
rect 9373 36188 9397 36244
rect 9453 36188 9477 36244
rect 9533 36188 9557 36244
rect 9613 36188 9637 36244
rect 9693 36188 9717 36244
rect 9773 36188 9797 36244
rect 9853 36188 9877 36244
rect 9933 36188 9957 36244
rect 10013 36188 10022 36244
rect 4663 36158 10022 36188
rect 4663 36102 8035 36158
rect 8091 36102 8116 36158
rect 8172 36102 8197 36158
rect 8253 36102 8277 36158
rect 8333 36102 8357 36158
rect 8413 36102 8437 36158
rect 8493 36102 8517 36158
rect 8573 36102 8597 36158
rect 8653 36102 8677 36158
rect 8733 36102 8757 36158
rect 8813 36102 8837 36158
rect 8893 36102 8917 36158
rect 8973 36102 8997 36158
rect 9053 36102 9077 36158
rect 9133 36102 9157 36158
rect 9213 36102 9237 36158
rect 9293 36102 9317 36158
rect 9373 36102 9397 36158
rect 9453 36102 9477 36158
rect 9533 36102 9557 36158
rect 9613 36102 9637 36158
rect 9693 36102 9717 36158
rect 9773 36102 9797 36158
rect 9853 36102 9877 36158
rect 9933 36102 9957 36158
rect 10013 36102 10022 36158
rect 4663 36072 10022 36102
rect 4663 36016 8035 36072
rect 8091 36016 8116 36072
rect 8172 36016 8197 36072
rect 8253 36016 8277 36072
rect 8333 36016 8357 36072
rect 8413 36016 8437 36072
rect 8493 36016 8517 36072
rect 8573 36016 8597 36072
rect 8653 36016 8677 36072
rect 8733 36016 8757 36072
rect 8813 36016 8837 36072
rect 8893 36016 8917 36072
rect 8973 36016 8997 36072
rect 9053 36016 9077 36072
rect 9133 36016 9157 36072
rect 9213 36016 9237 36072
rect 9293 36016 9317 36072
rect 9373 36016 9397 36072
rect 9453 36016 9477 36072
rect 9533 36016 9557 36072
rect 9613 36016 9637 36072
rect 9693 36016 9717 36072
rect 9773 36016 9797 36072
rect 9853 36016 9877 36072
rect 9933 36016 9957 36072
rect 10013 36016 10022 36072
rect 4663 35986 10022 36016
rect 4663 35930 8035 35986
rect 8091 35930 8116 35986
rect 8172 35930 8197 35986
rect 8253 35930 8277 35986
rect 8333 35930 8357 35986
rect 8413 35930 8437 35986
rect 8493 35930 8517 35986
rect 8573 35930 8597 35986
rect 8653 35930 8677 35986
rect 8733 35930 8757 35986
rect 8813 35930 8837 35986
rect 8893 35930 8917 35986
rect 8973 35930 8997 35986
rect 9053 35930 9077 35986
rect 9133 35930 9157 35986
rect 9213 35930 9237 35986
rect 9293 35930 9317 35986
rect 9373 35930 9397 35986
rect 9453 35930 9477 35986
rect 9533 35930 9557 35986
rect 9613 35930 9637 35986
rect 9693 35930 9717 35986
rect 9773 35930 9797 35986
rect 9853 35930 9877 35986
rect 9933 35930 9957 35986
rect 10013 35930 10022 35986
rect 4663 35900 10022 35930
rect 4663 35844 8035 35900
rect 8091 35844 8116 35900
rect 8172 35844 8197 35900
rect 8253 35844 8277 35900
rect 8333 35844 8357 35900
rect 8413 35844 8437 35900
rect 8493 35844 8517 35900
rect 8573 35844 8597 35900
rect 8653 35844 8677 35900
rect 8733 35844 8757 35900
rect 8813 35844 8837 35900
rect 8893 35844 8917 35900
rect 8973 35844 8997 35900
rect 9053 35844 9077 35900
rect 9133 35844 9157 35900
rect 9213 35844 9237 35900
rect 9293 35844 9317 35900
rect 9373 35844 9397 35900
rect 9453 35844 9477 35900
rect 9533 35844 9557 35900
rect 9613 35844 9637 35900
rect 9693 35844 9717 35900
rect 9773 35844 9797 35900
rect 9853 35844 9877 35900
rect 9933 35844 9957 35900
rect 10013 35844 10022 35900
rect 4663 35814 10022 35844
rect 4663 35758 8035 35814
rect 8091 35758 8116 35814
rect 8172 35758 8197 35814
rect 8253 35758 8277 35814
rect 8333 35758 8357 35814
rect 8413 35758 8437 35814
rect 8493 35758 8517 35814
rect 8573 35758 8597 35814
rect 8653 35758 8677 35814
rect 8733 35758 8757 35814
rect 8813 35758 8837 35814
rect 8893 35758 8917 35814
rect 8973 35758 8997 35814
rect 9053 35758 9077 35814
rect 9133 35758 9157 35814
rect 9213 35758 9237 35814
rect 9293 35758 9317 35814
rect 9373 35758 9397 35814
rect 9453 35758 9477 35814
rect 9533 35758 9557 35814
rect 9613 35758 9637 35814
rect 9693 35758 9717 35814
rect 9773 35758 9797 35814
rect 9853 35758 9877 35814
rect 9933 35758 9957 35814
rect 10013 35758 10022 35814
rect 4663 35728 10022 35758
rect 4663 35672 8035 35728
rect 8091 35672 8116 35728
rect 8172 35672 8197 35728
rect 8253 35672 8277 35728
rect 8333 35672 8357 35728
rect 8413 35672 8437 35728
rect 8493 35672 8517 35728
rect 8573 35672 8597 35728
rect 8653 35672 8677 35728
rect 8733 35672 8757 35728
rect 8813 35672 8837 35728
rect 8893 35672 8917 35728
rect 8973 35672 8997 35728
rect 9053 35672 9077 35728
rect 9133 35672 9157 35728
rect 9213 35672 9237 35728
rect 9293 35672 9317 35728
rect 9373 35672 9397 35728
rect 9453 35672 9477 35728
rect 9533 35672 9557 35728
rect 9613 35672 9637 35728
rect 9693 35672 9717 35728
rect 9773 35672 9797 35728
rect 9853 35672 9877 35728
rect 9933 35672 9957 35728
rect 10013 35672 10022 35728
rect 4663 35642 10022 35672
rect 4663 35586 8035 35642
rect 8091 35586 8116 35642
rect 8172 35586 8197 35642
rect 8253 35586 8277 35642
rect 8333 35586 8357 35642
rect 8413 35586 8437 35642
rect 8493 35586 8517 35642
rect 8573 35586 8597 35642
rect 8653 35586 8677 35642
rect 8733 35586 8757 35642
rect 8813 35586 8837 35642
rect 8893 35586 8917 35642
rect 8973 35586 8997 35642
rect 9053 35586 9077 35642
rect 9133 35586 9157 35642
rect 9213 35586 9237 35642
rect 9293 35586 9317 35642
rect 9373 35586 9397 35642
rect 9453 35586 9477 35642
rect 9533 35586 9557 35642
rect 9613 35586 9637 35642
rect 9693 35586 9717 35642
rect 9773 35586 9797 35642
rect 9853 35586 9877 35642
rect 9933 35586 9957 35642
rect 10013 35586 10022 35642
rect 4663 35556 10022 35586
rect 4663 35500 8035 35556
rect 8091 35500 8116 35556
rect 8172 35500 8197 35556
rect 8253 35500 8277 35556
rect 8333 35500 8357 35556
rect 8413 35500 8437 35556
rect 8493 35500 8517 35556
rect 8573 35500 8597 35556
rect 8653 35500 8677 35556
rect 8733 35500 8757 35556
rect 8813 35500 8837 35556
rect 8893 35500 8917 35556
rect 8973 35500 8997 35556
rect 9053 35500 9077 35556
rect 9133 35500 9157 35556
rect 9213 35500 9237 35556
rect 9293 35500 9317 35556
rect 9373 35500 9397 35556
rect 9453 35500 9477 35556
rect 9533 35500 9557 35556
rect 9613 35500 9637 35556
rect 9693 35500 9717 35556
rect 9773 35500 9797 35556
rect 9853 35500 9877 35556
rect 9933 35500 9957 35556
rect 10013 35500 10022 35556
rect 4663 35470 10022 35500
rect 4663 35414 8035 35470
rect 8091 35414 8116 35470
rect 8172 35414 8197 35470
rect 8253 35414 8277 35470
rect 8333 35414 8357 35470
rect 8413 35414 8437 35470
rect 8493 35414 8517 35470
rect 8573 35414 8597 35470
rect 8653 35414 8677 35470
rect 8733 35414 8757 35470
rect 8813 35414 8837 35470
rect 8893 35414 8917 35470
rect 8973 35414 8997 35470
rect 9053 35414 9077 35470
rect 9133 35414 9157 35470
rect 9213 35414 9237 35470
rect 9293 35414 9317 35470
rect 9373 35414 9397 35470
rect 9453 35414 9477 35470
rect 9533 35414 9557 35470
rect 9613 35414 9637 35470
rect 9693 35414 9717 35470
rect 9773 35414 9797 35470
rect 9853 35414 9877 35470
rect 9933 35414 9957 35470
rect 10013 35414 10022 35470
rect 4663 35372 10022 35414
tri 5663 34362 6673 35372 nw
rect 8481 30336 8490 30338
rect 8546 30336 8570 30338
rect 8481 30284 8488 30336
rect 8546 30284 8552 30336
rect 8481 30282 8490 30284
rect 8546 30282 8570 30284
rect 8626 30282 8635 30338
rect 8481 30082 8487 30134
rect 8539 30082 8551 30134
rect 8603 30082 8609 30134
rect 8481 30002 8487 30054
rect 8539 30002 8551 30054
rect 8603 30002 8609 30054
rect 8481 29922 8487 29974
rect 8539 29922 8551 29974
rect 8603 29922 8609 29974
rect 8481 29842 8487 29894
rect 8539 29842 8551 29894
rect 8603 29842 8609 29894
rect 8481 29762 8487 29814
rect 8539 29762 8551 29814
rect 8603 29762 8609 29814
rect 8481 29647 8487 29699
rect 8539 29647 8551 29699
rect 8603 29647 8609 29699
rect 8481 29460 8490 29462
rect 8546 29460 8570 29462
rect 8481 29408 8488 29460
rect 8546 29408 8552 29460
rect 8481 29406 8490 29408
rect 8546 29406 8570 29408
rect 8626 29406 8635 29462
rect 3550 28871 8035 28927
rect 8091 28871 8116 28927
rect 8172 28871 8197 28927
rect 8253 28871 8277 28927
rect 8333 28871 8357 28927
rect 8413 28871 8437 28927
rect 8493 28871 8517 28927
rect 8573 28871 8597 28927
rect 8653 28871 8677 28927
rect 8733 28871 8757 28927
rect 8813 28871 8837 28927
rect 8893 28871 8917 28927
rect 8973 28871 8997 28927
rect 9053 28871 9077 28927
rect 9133 28871 9157 28927
rect 9213 28871 9237 28927
rect 9293 28871 9317 28927
rect 9373 28871 9397 28927
rect 9453 28871 9477 28927
rect 9533 28871 9557 28927
rect 9613 28871 9637 28927
rect 9693 28871 9717 28927
rect 9773 28871 9797 28927
rect 9853 28871 9877 28927
rect 9933 28871 9957 28927
rect 10013 28871 10022 28927
rect 3550 28815 10022 28871
rect 3550 28759 8035 28815
rect 8091 28759 8116 28815
rect 8172 28759 8197 28815
rect 8253 28759 8277 28815
rect 8333 28759 8357 28815
rect 8413 28759 8437 28815
rect 8493 28759 8517 28815
rect 8573 28759 8597 28815
rect 8653 28759 8677 28815
rect 8733 28759 8757 28815
rect 8813 28759 8837 28815
rect 8893 28759 8917 28815
rect 8973 28759 8997 28815
rect 9053 28759 9077 28815
rect 9133 28759 9157 28815
rect 9213 28759 9237 28815
rect 9293 28759 9317 28815
rect 9373 28759 9397 28815
rect 9453 28759 9477 28815
rect 9533 28759 9557 28815
rect 9613 28759 9637 28815
rect 9693 28759 9717 28815
rect 9773 28759 9797 28815
rect 9853 28759 9877 28815
rect 9933 28759 9957 28815
rect 10013 28759 10022 28815
rect 3550 28703 10022 28759
rect 3550 28647 8035 28703
rect 8091 28647 8116 28703
rect 8172 28647 8197 28703
rect 8253 28647 8277 28703
rect 8333 28647 8357 28703
rect 8413 28647 8437 28703
rect 8493 28647 8517 28703
rect 8573 28647 8597 28703
rect 8653 28647 8677 28703
rect 8733 28647 8757 28703
rect 8813 28647 8837 28703
rect 8893 28647 8917 28703
rect 8973 28647 8997 28703
rect 9053 28647 9077 28703
rect 9133 28647 9157 28703
rect 9213 28647 9237 28703
rect 9293 28647 9317 28703
rect 9373 28647 9397 28703
rect 9453 28647 9477 28703
rect 9533 28647 9557 28703
rect 9613 28647 9637 28703
rect 9693 28647 9717 28703
rect 9773 28647 9797 28703
rect 9853 28647 9877 28703
rect 9933 28647 9957 28703
rect 10013 28647 10022 28703
rect 354 27992 9862 27994
rect 354 27988 2670 27992
rect 354 27936 366 27988
rect 418 27936 432 27988
rect 484 27936 2481 27988
rect 2533 27936 2547 27988
rect 2599 27936 2670 27988
rect 2726 27936 2759 27992
rect 2815 27936 2848 27992
rect 2904 27936 2937 27992
rect 2993 27936 3025 27992
rect 3081 27936 3113 27992
rect 3169 27936 3201 27992
rect 3257 27936 3289 27992
rect 3345 27936 3377 27992
rect 3433 27988 9862 27992
rect 3433 27936 9732 27988
rect 9784 27936 9810 27988
rect 354 27921 9862 27936
rect 354 27869 366 27921
rect 418 27869 432 27921
rect 484 27869 2481 27921
rect 2533 27869 2547 27921
rect 2599 27912 9732 27921
rect 2599 27902 2878 27912
rect 2930 27902 3008 27912
rect 3060 27902 3138 27912
rect 3190 27902 3268 27912
rect 3320 27902 3398 27912
rect 2599 27869 2670 27902
rect 354 27854 2670 27869
rect 354 27802 366 27854
rect 418 27802 432 27854
rect 484 27802 2481 27854
rect 2533 27802 2547 27854
rect 2599 27846 2670 27854
rect 2726 27846 2759 27902
rect 2815 27846 2848 27902
rect 2930 27860 2937 27902
rect 2904 27846 2937 27860
rect 2993 27860 3008 27902
rect 2993 27846 3025 27860
rect 3081 27846 3113 27902
rect 3190 27860 3201 27902
rect 3169 27846 3201 27860
rect 3257 27860 3268 27902
rect 3257 27846 3289 27860
rect 3345 27846 3377 27902
rect 3450 27860 3528 27912
rect 3580 27860 3658 27912
rect 3710 27860 3788 27912
rect 3840 27860 3918 27912
rect 3970 27860 4048 27912
rect 4100 27860 4178 27912
rect 4230 27860 4308 27912
rect 4360 27860 4438 27912
rect 4490 27860 4568 27912
rect 4620 27860 4698 27912
rect 4750 27860 4828 27912
rect 4880 27860 4958 27912
rect 5010 27860 5088 27912
rect 5140 27860 5218 27912
rect 5270 27860 5348 27912
rect 5400 27860 5478 27912
rect 5530 27860 5608 27912
rect 5660 27860 5738 27912
rect 5790 27860 5868 27912
rect 5920 27860 5998 27912
rect 6050 27860 6128 27912
rect 6180 27860 6258 27912
rect 6310 27860 6388 27912
rect 6440 27860 6517 27912
rect 6569 27860 6646 27912
rect 6698 27860 6775 27912
rect 6827 27860 6904 27912
rect 6956 27860 7033 27912
rect 7085 27860 7162 27912
rect 7214 27860 7291 27912
rect 7343 27860 7420 27912
rect 7472 27860 7549 27912
rect 7601 27860 7678 27912
rect 7730 27860 7807 27912
rect 7859 27860 7936 27912
rect 7988 27869 9732 27912
rect 9784 27869 9810 27921
rect 7988 27860 9862 27869
rect 3433 27854 9862 27860
rect 3433 27846 9732 27854
rect 2599 27832 9732 27846
rect 2599 27812 2878 27832
rect 2930 27812 3008 27832
rect 3060 27812 3138 27832
rect 3190 27812 3268 27832
rect 3320 27812 3398 27832
rect 2599 27802 2670 27812
rect 354 27787 2670 27802
rect 354 27735 366 27787
rect 418 27735 432 27787
rect 484 27735 2481 27787
rect 2533 27735 2547 27787
rect 2599 27756 2670 27787
rect 2726 27756 2759 27812
rect 2815 27756 2848 27812
rect 2930 27780 2937 27812
rect 2904 27756 2937 27780
rect 2993 27780 3008 27812
rect 2993 27756 3025 27780
rect 3081 27756 3113 27812
rect 3190 27780 3201 27812
rect 3169 27756 3201 27780
rect 3257 27780 3268 27812
rect 3257 27756 3289 27780
rect 3345 27756 3377 27812
rect 3450 27780 3528 27832
rect 3580 27780 3658 27832
rect 3710 27780 3788 27832
rect 3840 27780 3918 27832
rect 3970 27780 4048 27832
rect 4100 27780 4178 27832
rect 4230 27780 4308 27832
rect 4360 27780 4438 27832
rect 4490 27780 4568 27832
rect 4620 27780 4698 27832
rect 4750 27780 4828 27832
rect 4880 27780 4958 27832
rect 5010 27780 5088 27832
rect 5140 27780 5218 27832
rect 5270 27780 5348 27832
rect 5400 27780 5478 27832
rect 5530 27780 5608 27832
rect 5660 27780 5738 27832
rect 5790 27780 5868 27832
rect 5920 27780 5998 27832
rect 6050 27780 6128 27832
rect 6180 27780 6258 27832
rect 6310 27780 6388 27832
rect 6440 27780 6517 27832
rect 6569 27780 6646 27832
rect 6698 27780 6775 27832
rect 6827 27780 6904 27832
rect 6956 27780 7033 27832
rect 7085 27780 7162 27832
rect 7214 27780 7291 27832
rect 7343 27780 7420 27832
rect 7472 27780 7549 27832
rect 7601 27780 7678 27832
rect 7730 27780 7807 27832
rect 7859 27780 7936 27832
rect 7988 27802 9732 27832
rect 9784 27802 9810 27854
rect 7988 27787 9862 27802
rect 7988 27780 9732 27787
rect 3433 27756 9732 27780
rect 2599 27752 9732 27756
rect 2599 27735 2878 27752
rect 354 27722 2878 27735
rect 2930 27722 3008 27752
rect 3060 27722 3138 27752
rect 3190 27722 3268 27752
rect 3320 27722 3398 27752
rect 354 27720 2670 27722
rect 354 27668 366 27720
rect 418 27668 432 27720
rect 484 27668 2481 27720
rect 2533 27668 2547 27720
rect 2599 27668 2670 27720
rect 354 27666 2670 27668
rect 2726 27666 2759 27722
rect 2815 27666 2848 27722
rect 2930 27700 2937 27722
rect 2904 27672 2937 27700
rect 2930 27666 2937 27672
rect 2993 27700 3008 27722
rect 2993 27672 3025 27700
rect 2993 27666 3008 27672
rect 3081 27666 3113 27722
rect 3190 27700 3201 27722
rect 3169 27672 3201 27700
rect 3190 27666 3201 27672
rect 3257 27700 3268 27722
rect 3257 27672 3289 27700
rect 3257 27666 3268 27672
rect 3345 27666 3377 27722
rect 3450 27700 3528 27752
rect 3580 27700 3658 27752
rect 3710 27700 3788 27752
rect 3840 27700 3918 27752
rect 3970 27700 4048 27752
rect 4100 27700 4178 27752
rect 4230 27700 4308 27752
rect 4360 27700 4438 27752
rect 4490 27700 4568 27752
rect 4620 27700 4698 27752
rect 4750 27700 4828 27752
rect 4880 27700 4958 27752
rect 5010 27700 5088 27752
rect 5140 27700 5218 27752
rect 5270 27700 5348 27752
rect 5400 27700 5478 27752
rect 5530 27700 5608 27752
rect 5660 27700 5738 27752
rect 5790 27700 5868 27752
rect 5920 27700 5998 27752
rect 6050 27700 6128 27752
rect 6180 27700 6258 27752
rect 6310 27700 6388 27752
rect 6440 27700 6517 27752
rect 6569 27700 6646 27752
rect 6698 27700 6775 27752
rect 6827 27700 6904 27752
rect 6956 27700 7033 27752
rect 7085 27700 7162 27752
rect 7214 27700 7291 27752
rect 7343 27700 7420 27752
rect 7472 27700 7549 27752
rect 7601 27700 7678 27752
rect 7730 27700 7807 27752
rect 7859 27700 7936 27752
rect 7988 27735 9732 27752
rect 9784 27735 9810 27787
rect 7988 27720 9862 27735
rect 7988 27700 9732 27720
rect 3433 27672 9732 27700
rect 354 27653 2878 27666
rect 354 27601 366 27653
rect 418 27601 432 27653
rect 484 27601 2481 27653
rect 2533 27601 2547 27653
rect 2599 27632 2878 27653
rect 2930 27632 3008 27666
rect 3060 27632 3138 27666
rect 3190 27632 3268 27666
rect 3320 27632 3398 27666
rect 2599 27601 2670 27632
rect 354 27586 2670 27601
rect 354 27534 366 27586
rect 418 27534 432 27586
rect 484 27534 2481 27586
rect 2533 27534 2547 27586
rect 2599 27576 2670 27586
rect 2726 27576 2759 27632
rect 2815 27576 2848 27632
rect 2930 27620 2937 27632
rect 2904 27592 2937 27620
rect 2930 27576 2937 27592
rect 2993 27620 3008 27632
rect 2993 27592 3025 27620
rect 2993 27576 3008 27592
rect 3081 27576 3113 27632
rect 3190 27620 3201 27632
rect 3169 27592 3201 27620
rect 3190 27576 3201 27592
rect 3257 27620 3268 27632
rect 3257 27592 3289 27620
rect 3257 27576 3268 27592
rect 3345 27576 3377 27632
rect 3450 27620 3528 27672
rect 3580 27620 3658 27672
rect 3710 27620 3788 27672
rect 3840 27620 3918 27672
rect 3970 27620 4048 27672
rect 4100 27620 4178 27672
rect 4230 27620 4308 27672
rect 4360 27620 4438 27672
rect 4490 27620 4568 27672
rect 4620 27620 4698 27672
rect 4750 27620 4828 27672
rect 4880 27620 4958 27672
rect 5010 27620 5088 27672
rect 5140 27620 5218 27672
rect 5270 27620 5348 27672
rect 5400 27620 5478 27672
rect 5530 27620 5608 27672
rect 5660 27620 5738 27672
rect 5790 27620 5868 27672
rect 5920 27620 5998 27672
rect 6050 27620 6128 27672
rect 6180 27620 6258 27672
rect 6310 27620 6388 27672
rect 6440 27620 6517 27672
rect 6569 27620 6646 27672
rect 6698 27620 6775 27672
rect 6827 27620 6904 27672
rect 6956 27620 7033 27672
rect 7085 27620 7162 27672
rect 7214 27620 7291 27672
rect 7343 27620 7420 27672
rect 7472 27620 7549 27672
rect 7601 27620 7678 27672
rect 7730 27620 7807 27672
rect 7859 27620 7936 27672
rect 7988 27668 9732 27672
rect 9784 27668 9810 27720
rect 7988 27653 9862 27668
rect 7988 27620 9732 27653
rect 3433 27601 9732 27620
rect 9784 27601 9810 27653
rect 3433 27592 9862 27601
rect 2599 27542 2878 27576
rect 2930 27542 3008 27576
rect 3060 27542 3138 27576
rect 3190 27542 3268 27576
rect 3320 27542 3398 27576
rect 2599 27534 2670 27542
rect 354 27519 2670 27534
rect 354 27467 366 27519
rect 418 27467 432 27519
rect 484 27467 2481 27519
rect 2533 27467 2547 27519
rect 2599 27486 2670 27519
rect 2726 27486 2759 27542
rect 2815 27486 2848 27542
rect 2930 27540 2937 27542
rect 2904 27512 2937 27540
rect 2930 27486 2937 27512
rect 2993 27540 3008 27542
rect 2993 27512 3025 27540
rect 2993 27486 3008 27512
rect 3081 27486 3113 27542
rect 3190 27540 3201 27542
rect 3169 27512 3201 27540
rect 3190 27486 3201 27512
rect 3257 27540 3268 27542
rect 3257 27512 3289 27540
rect 3257 27486 3268 27512
rect 3345 27486 3377 27542
rect 3450 27540 3528 27592
rect 3580 27540 3658 27592
rect 3710 27540 3788 27592
rect 3840 27540 3918 27592
rect 3970 27540 4048 27592
rect 4100 27540 4178 27592
rect 4230 27540 4308 27592
rect 4360 27540 4438 27592
rect 4490 27540 4568 27592
rect 4620 27540 4698 27592
rect 4750 27540 4828 27592
rect 4880 27540 4958 27592
rect 5010 27540 5088 27592
rect 5140 27540 5218 27592
rect 5270 27540 5348 27592
rect 5400 27540 5478 27592
rect 5530 27540 5608 27592
rect 5660 27540 5738 27592
rect 5790 27540 5868 27592
rect 5920 27540 5998 27592
rect 6050 27540 6128 27592
rect 6180 27540 6258 27592
rect 6310 27540 6388 27592
rect 6440 27540 6517 27592
rect 6569 27540 6646 27592
rect 6698 27540 6775 27592
rect 6827 27540 6904 27592
rect 6956 27540 7033 27592
rect 7085 27540 7162 27592
rect 7214 27540 7291 27592
rect 7343 27540 7420 27592
rect 7472 27540 7549 27592
rect 7601 27540 7678 27592
rect 7730 27540 7807 27592
rect 7859 27540 7936 27592
rect 7988 27586 9862 27592
rect 7988 27540 9732 27586
rect 3433 27534 9732 27540
rect 9784 27534 9810 27586
rect 3433 27519 9862 27534
rect 3433 27512 9732 27519
rect 2599 27467 2878 27486
rect 354 27460 2878 27467
rect 2930 27460 3008 27486
rect 3060 27460 3138 27486
rect 3190 27460 3268 27486
rect 3320 27460 3398 27486
rect 3450 27460 3528 27512
rect 3580 27460 3658 27512
rect 3710 27460 3788 27512
rect 3840 27460 3918 27512
rect 3970 27460 4048 27512
rect 4100 27460 4178 27512
rect 4230 27460 4308 27512
rect 4360 27460 4438 27512
rect 4490 27460 4568 27512
rect 4620 27460 4698 27512
rect 4750 27460 4828 27512
rect 4880 27460 4958 27512
rect 5010 27460 5088 27512
rect 5140 27460 5218 27512
rect 5270 27460 5348 27512
rect 5400 27460 5478 27512
rect 5530 27460 5608 27512
rect 5660 27460 5738 27512
rect 5790 27460 5868 27512
rect 5920 27460 5998 27512
rect 6050 27460 6128 27512
rect 6180 27460 6258 27512
rect 6310 27460 6388 27512
rect 6440 27460 6517 27512
rect 6569 27460 6646 27512
rect 6698 27460 6775 27512
rect 6827 27460 6904 27512
rect 6956 27460 7033 27512
rect 7085 27460 7162 27512
rect 7214 27460 7291 27512
rect 7343 27460 7420 27512
rect 7472 27460 7549 27512
rect 7601 27460 7678 27512
rect 7730 27460 7807 27512
rect 7859 27460 7936 27512
rect 7988 27467 9732 27512
rect 9784 27467 9810 27519
rect 7988 27460 9862 27467
rect 354 27452 9862 27460
rect 354 27400 366 27452
rect 418 27400 432 27452
rect 484 27400 2481 27452
rect 2533 27400 2547 27452
rect 2599 27400 2670 27452
rect 354 27396 2670 27400
rect 2726 27396 2759 27452
rect 2815 27396 2848 27452
rect 2904 27396 2937 27452
rect 2993 27396 3025 27452
rect 3081 27396 3113 27452
rect 3169 27396 3201 27452
rect 3257 27396 3289 27452
rect 3345 27396 3377 27452
rect 3433 27400 9732 27452
rect 9784 27400 9810 27452
rect 3433 27396 9862 27400
rect 354 27394 9862 27396
tri 5349 27360 5383 27394 ne
rect 2494 27327 3310 27336
rect 2550 27284 3310 27327
rect 3362 27284 3376 27336
rect 3428 27284 3434 27336
rect 2550 27271 3434 27284
rect 2494 27270 3434 27271
rect 2494 27247 3310 27270
rect 2550 27218 3310 27247
rect 3362 27218 3376 27270
rect 3428 27218 3434 27270
rect 5383 27334 5511 27394
tri 5511 27360 5545 27394 nw
rect 5383 27218 5389 27334
rect 5505 27218 5511 27334
rect 2494 27182 2550 27191
tri 2550 27184 2584 27218 nw
rect 3268 26852 7908 26853
rect 3268 26847 6742 26852
rect 3268 26795 3269 26847
rect 3321 26795 3337 26847
rect 3389 26795 3405 26847
rect 3457 26796 6742 26847
rect 6798 26796 6827 26852
rect 6883 26796 6912 26852
rect 6968 26796 6997 26852
rect 7053 26796 7082 26852
rect 7138 26796 7167 26852
rect 7223 26796 7252 26852
rect 7308 26796 7337 26852
rect 7393 26796 7422 26852
rect 7478 26796 7507 26852
rect 7563 26796 7591 26852
rect 7647 26796 7675 26852
rect 7731 26796 7759 26852
rect 7815 26796 7843 26852
rect 7899 26796 7908 26852
rect 3457 26795 7908 26796
rect 3268 26766 7908 26795
rect 3268 26763 6742 26766
rect 3268 26711 3269 26763
rect 3321 26711 3337 26763
rect 3389 26711 3405 26763
rect 3457 26711 6742 26763
rect 3268 26710 6742 26711
rect 6798 26710 6827 26766
rect 6883 26710 6912 26766
rect 6968 26710 6997 26766
rect 7053 26710 7082 26766
rect 7138 26710 7167 26766
rect 7223 26710 7252 26766
rect 7308 26710 7337 26766
rect 7393 26710 7422 26766
rect 7478 26710 7507 26766
rect 7563 26710 7591 26766
rect 7647 26710 7675 26766
rect 7731 26710 7759 26766
rect 7815 26710 7843 26766
rect 7899 26710 7908 26766
rect 3268 26680 7908 26710
rect 3268 26679 6742 26680
rect 3268 26627 3269 26679
rect 3321 26627 3337 26679
rect 3389 26627 3405 26679
rect 3457 26627 6742 26679
rect 3268 26624 6742 26627
rect 6798 26624 6827 26680
rect 6883 26624 6912 26680
rect 6968 26624 6997 26680
rect 7053 26624 7082 26680
rect 7138 26624 7167 26680
rect 7223 26624 7252 26680
rect 7308 26624 7337 26680
rect 7393 26624 7422 26680
rect 7478 26624 7507 26680
rect 7563 26624 7591 26680
rect 7647 26624 7675 26680
rect 7731 26624 7759 26680
rect 7815 26624 7843 26680
rect 7899 26624 7908 26680
rect 3268 26594 7908 26624
rect 3268 26542 3269 26594
rect 3321 26542 3337 26594
rect 3389 26542 3405 26594
rect 3457 26542 6742 26594
rect 3268 26538 6742 26542
rect 6798 26538 6827 26594
rect 6883 26538 6912 26594
rect 6968 26538 6997 26594
rect 7053 26538 7082 26594
rect 7138 26538 7167 26594
rect 7223 26538 7252 26594
rect 7308 26538 7337 26594
rect 7393 26538 7422 26594
rect 7478 26538 7507 26594
rect 7563 26538 7591 26594
rect 7647 26538 7675 26594
rect 7731 26538 7759 26594
rect 7815 26538 7843 26594
rect 7899 26538 7908 26594
rect 3268 26509 7908 26538
rect 3268 26457 3269 26509
rect 3321 26457 3337 26509
rect 3389 26457 3405 26509
rect 3457 26508 7908 26509
rect 3457 26457 6742 26508
rect 3268 26452 6742 26457
rect 6798 26452 6827 26508
rect 6883 26452 6912 26508
rect 6968 26452 6997 26508
rect 7053 26452 7082 26508
rect 7138 26452 7167 26508
rect 7223 26452 7252 26508
rect 7308 26452 7337 26508
rect 7393 26452 7422 26508
rect 7478 26452 7507 26508
rect 7563 26452 7591 26508
rect 7647 26452 7675 26508
rect 7731 26452 7759 26508
rect 7815 26452 7843 26508
rect 7899 26452 7908 26508
rect 3268 26451 7908 26452
rect 2661 24467 2670 24523
rect 2726 24467 2751 24523
rect 2807 24467 2832 24523
rect 2888 24467 2913 24523
rect 2969 24467 2994 24523
rect 3050 24467 3075 24523
rect 3131 24467 3156 24523
rect 3212 24467 3237 24523
rect 3293 24467 3318 24523
rect 3374 24467 3398 24523
rect 3454 24467 3478 24523
rect 3534 24522 10828 24523
rect 3534 24470 4056 24522
rect 4108 24470 4187 24522
rect 4239 24470 4318 24522
rect 4370 24470 4449 24522
rect 4501 24470 4580 24522
rect 4632 24470 4711 24522
rect 4763 24470 4842 24522
rect 4894 24470 4973 24522
rect 5025 24470 5104 24522
rect 5156 24470 5235 24522
rect 5287 24470 5365 24522
rect 5417 24470 5495 24522
rect 5547 24470 5625 24522
rect 5677 24470 5755 24522
rect 5807 24470 5885 24522
rect 5937 24470 6015 24522
rect 6067 24517 10828 24522
rect 6067 24470 7988 24517
rect 3534 24467 7988 24470
rect 2661 24465 7988 24467
rect 8040 24465 9732 24517
rect 9784 24465 9810 24517
rect 9862 24465 10710 24517
rect 10762 24465 10776 24517
rect 2661 24458 10828 24465
rect 2661 24406 4056 24458
rect 4108 24406 4187 24458
rect 4239 24406 4318 24458
rect 4370 24406 4449 24458
rect 4501 24406 4580 24458
rect 4632 24406 4711 24458
rect 4763 24406 4842 24458
rect 4894 24406 4973 24458
rect 5025 24406 5104 24458
rect 5156 24406 5235 24458
rect 5287 24406 5365 24458
rect 5417 24406 5495 24458
rect 5547 24406 5625 24458
rect 5677 24406 5755 24458
rect 5807 24406 5885 24458
rect 5937 24406 6015 24458
rect 6067 24406 10828 24458
rect 2661 24399 10828 24406
rect 2661 24397 7988 24399
rect 2661 24341 2670 24397
rect 2726 24341 2751 24397
rect 2807 24341 2832 24397
rect 2888 24341 2913 24397
rect 2969 24341 2994 24397
rect 3050 24341 3075 24397
rect 3131 24341 3156 24397
rect 3212 24341 3237 24397
rect 3293 24341 3318 24397
rect 3374 24341 3398 24397
rect 3454 24341 3478 24397
rect 3534 24394 7988 24397
rect 3534 24342 4056 24394
rect 4108 24342 4187 24394
rect 4239 24342 4318 24394
rect 4370 24342 4449 24394
rect 4501 24342 4580 24394
rect 4632 24342 4711 24394
rect 4763 24342 4842 24394
rect 4894 24342 4973 24394
rect 5025 24342 5104 24394
rect 5156 24342 5235 24394
rect 5287 24342 5365 24394
rect 5417 24342 5495 24394
rect 5547 24342 5625 24394
rect 5677 24342 5755 24394
rect 5807 24342 5885 24394
rect 5937 24342 6015 24394
rect 6067 24347 7988 24394
rect 8040 24347 9732 24399
rect 9784 24347 9810 24399
rect 9862 24347 10710 24399
rect 10762 24347 10776 24399
rect 6067 24342 10828 24347
rect 3534 24341 10828 24342
rect 2661 23212 2670 23268
rect 2726 23212 2751 23268
rect 2807 23212 2832 23268
rect 2888 23212 2913 23268
rect 2969 23212 2994 23268
rect 3050 23212 3075 23268
rect 3131 23212 3156 23268
rect 3212 23212 3237 23268
rect 3293 23212 3318 23268
rect 3374 23212 3398 23268
rect 3454 23212 3478 23268
rect 3534 23265 7775 23268
rect 3534 23213 6056 23265
rect 6108 23213 6123 23265
rect 6175 23213 6190 23265
rect 6242 23213 6257 23265
rect 6309 23213 6324 23265
rect 6376 23213 6391 23265
rect 6443 23213 6458 23265
rect 6510 23213 6525 23265
rect 6577 23213 6592 23265
rect 6644 23213 6659 23265
rect 6711 23213 6726 23265
rect 6778 23213 6792 23265
rect 6844 23213 6858 23265
rect 6910 23213 6924 23265
rect 6976 23213 6990 23265
rect 7042 23213 7056 23265
rect 7108 23213 7122 23265
rect 7174 23213 7188 23265
rect 7240 23213 7254 23265
rect 7306 23213 7320 23265
rect 7372 23213 7386 23265
rect 7438 23213 7452 23265
rect 7504 23213 7518 23265
rect 7570 23213 7584 23265
rect 7636 23213 7650 23265
rect 7702 23213 7716 23265
rect 7768 23213 7775 23265
rect 3534 23212 7775 23213
rect 2661 23195 7775 23212
rect 2661 23180 6056 23195
rect 2661 23124 2670 23180
rect 2726 23124 2751 23180
rect 2807 23124 2832 23180
rect 2888 23124 2913 23180
rect 2969 23124 2994 23180
rect 3050 23124 3075 23180
rect 3131 23124 3156 23180
rect 3212 23124 3237 23180
rect 3293 23124 3318 23180
rect 3374 23124 3398 23180
rect 3454 23124 3478 23180
rect 3534 23143 6056 23180
rect 6108 23143 6123 23195
rect 6175 23143 6190 23195
rect 6242 23143 6257 23195
rect 6309 23143 6324 23195
rect 6376 23143 6391 23195
rect 6443 23143 6458 23195
rect 6510 23143 6525 23195
rect 6577 23143 6592 23195
rect 6644 23143 6659 23195
rect 6711 23143 6726 23195
rect 6778 23143 6792 23195
rect 6844 23143 6858 23195
rect 6910 23143 6924 23195
rect 6976 23143 6990 23195
rect 7042 23143 7056 23195
rect 7108 23143 7122 23195
rect 7174 23143 7188 23195
rect 7240 23143 7254 23195
rect 7306 23143 7320 23195
rect 7372 23143 7386 23195
rect 7438 23143 7452 23195
rect 7504 23143 7518 23195
rect 7570 23143 7584 23195
rect 7636 23143 7650 23195
rect 7702 23143 7716 23195
rect 7768 23143 7775 23195
rect 3534 23125 7775 23143
rect 3534 23124 6056 23125
rect 2661 23092 6056 23124
rect 2661 23036 2670 23092
rect 2726 23036 2751 23092
rect 2807 23036 2832 23092
rect 2888 23036 2913 23092
rect 2969 23036 2994 23092
rect 3050 23036 3075 23092
rect 3131 23036 3156 23092
rect 3212 23036 3237 23092
rect 3293 23036 3318 23092
rect 3374 23036 3398 23092
rect 3454 23036 3478 23092
rect 3534 23073 6056 23092
rect 6108 23073 6123 23125
rect 6175 23073 6190 23125
rect 6242 23073 6257 23125
rect 6309 23073 6324 23125
rect 6376 23073 6391 23125
rect 6443 23073 6458 23125
rect 6510 23073 6525 23125
rect 6577 23073 6592 23125
rect 6644 23073 6659 23125
rect 6711 23073 6726 23125
rect 6778 23073 6792 23125
rect 6844 23073 6858 23125
rect 6910 23073 6924 23125
rect 6976 23073 6990 23125
rect 7042 23073 7056 23125
rect 7108 23073 7122 23125
rect 7174 23073 7188 23125
rect 7240 23073 7254 23125
rect 7306 23073 7320 23125
rect 7372 23073 7386 23125
rect 7438 23073 7452 23125
rect 7504 23073 7518 23125
rect 7570 23073 7584 23125
rect 7636 23073 7650 23125
rect 7702 23073 7716 23125
rect 7768 23073 7775 23125
rect 3534 23055 7775 23073
rect 3534 23036 6056 23055
rect 2661 23004 6056 23036
rect 2661 22948 2670 23004
rect 2726 22948 2751 23004
rect 2807 22948 2832 23004
rect 2888 22948 2913 23004
rect 2969 22948 2994 23004
rect 3050 22948 3075 23004
rect 3131 22948 3156 23004
rect 3212 22948 3237 23004
rect 3293 22948 3318 23004
rect 3374 22948 3398 23004
rect 3454 22948 3478 23004
rect 3534 23003 6056 23004
rect 6108 23003 6123 23055
rect 6175 23003 6190 23055
rect 6242 23003 6257 23055
rect 6309 23003 6324 23055
rect 6376 23003 6391 23055
rect 6443 23003 6458 23055
rect 6510 23003 6525 23055
rect 6577 23003 6592 23055
rect 6644 23003 6659 23055
rect 6711 23003 6726 23055
rect 6778 23003 6792 23055
rect 6844 23003 6858 23055
rect 6910 23003 6924 23055
rect 6976 23003 6990 23055
rect 7042 23003 7056 23055
rect 7108 23003 7122 23055
rect 7174 23003 7188 23055
rect 7240 23003 7254 23055
rect 7306 23003 7320 23055
rect 7372 23003 7386 23055
rect 7438 23003 7452 23055
rect 7504 23003 7518 23055
rect 7570 23003 7584 23055
rect 7636 23003 7650 23055
rect 7702 23003 7716 23055
rect 7768 23003 7775 23055
rect 3534 22985 7775 23003
rect 3534 22948 6056 22985
rect 2661 22933 6056 22948
rect 6108 22933 6123 22985
rect 6175 22933 6190 22985
rect 6242 22933 6257 22985
rect 6309 22933 6324 22985
rect 6376 22933 6391 22985
rect 6443 22933 6458 22985
rect 6510 22933 6525 22985
rect 6577 22933 6592 22985
rect 6644 22933 6659 22985
rect 6711 22933 6726 22985
rect 6778 22933 6792 22985
rect 6844 22933 6858 22985
rect 6910 22933 6924 22985
rect 6976 22933 6990 22985
rect 7042 22933 7056 22985
rect 7108 22933 7122 22985
rect 7174 22933 7188 22985
rect 7240 22933 7254 22985
rect 7306 22933 7320 22985
rect 7372 22933 7386 22985
rect 7438 22933 7452 22985
rect 7504 22933 7518 22985
rect 7570 22933 7584 22985
rect 7636 22933 7650 22985
rect 7702 22933 7716 22985
rect 7768 22933 7775 22985
rect 2661 22916 7775 22933
rect 2661 22860 2670 22916
rect 2726 22860 2751 22916
rect 2807 22860 2832 22916
rect 2888 22860 2913 22916
rect 2969 22860 2994 22916
rect 3050 22860 3075 22916
rect 3131 22860 3156 22916
rect 3212 22860 3237 22916
rect 3293 22860 3318 22916
rect 3374 22860 3398 22916
rect 3454 22860 3478 22916
rect 3534 22915 7775 22916
rect 3534 22863 6056 22915
rect 6108 22863 6123 22915
rect 6175 22863 6190 22915
rect 6242 22863 6257 22915
rect 6309 22863 6324 22915
rect 6376 22863 6391 22915
rect 6443 22863 6458 22915
rect 6510 22863 6525 22915
rect 6577 22863 6592 22915
rect 6644 22863 6659 22915
rect 6711 22863 6726 22915
rect 6778 22863 6792 22915
rect 6844 22863 6858 22915
rect 6910 22863 6924 22915
rect 6976 22863 6990 22915
rect 7042 22863 7056 22915
rect 7108 22863 7122 22915
rect 7174 22863 7188 22915
rect 7240 22863 7254 22915
rect 7306 22863 7320 22915
rect 7372 22863 7386 22915
rect 7438 22863 7452 22915
rect 7504 22863 7518 22915
rect 7570 22863 7584 22915
rect 7636 22863 7650 22915
rect 7702 22863 7716 22915
rect 7768 22863 7775 22915
rect 3534 22860 7775 22863
rect 282 22749 8229 22755
rect 334 22703 8229 22749
rect 8281 22703 8293 22755
rect 8345 22703 8351 22755
rect 282 22685 334 22697
tri 334 22669 368 22703 nw
rect 282 22627 334 22633
rect 3703 21102 3712 21158
rect 3768 21102 3793 21158
rect 3849 21102 3874 21158
rect 3930 21102 3955 21158
rect 4011 21102 4036 21158
rect 4092 21102 4117 21158
rect 4173 21102 4198 21158
rect 4254 21102 4278 21158
rect 4334 21102 4358 21158
rect 4414 21102 4438 21158
rect 4494 21152 7762 21158
rect 4494 21102 6847 21152
rect 3703 21100 6847 21102
rect 6899 21100 6949 21152
rect 7001 21100 7051 21152
rect 7103 21100 7710 21152
rect 3703 21085 7762 21100
rect 3703 21072 7710 21085
rect 3703 21016 3712 21072
rect 3768 21016 3793 21072
rect 3849 21016 3874 21072
rect 3930 21016 3955 21072
rect 4011 21016 4036 21072
rect 4092 21016 4117 21072
rect 4173 21016 4198 21072
rect 4254 21016 4278 21072
rect 4334 21016 4358 21072
rect 4414 21016 4438 21072
rect 4494 21068 7710 21072
rect 4494 21016 6847 21068
rect 6899 21016 6949 21068
rect 7001 21016 7051 21068
rect 7103 21033 7710 21068
rect 7103 21018 7762 21033
rect 7103 21016 7710 21018
rect 3703 20986 7710 21016
rect 3703 20930 3712 20986
rect 3768 20930 3793 20986
rect 3849 20930 3874 20986
rect 3930 20930 3955 20986
rect 4011 20930 4036 20986
rect 4092 20930 4117 20986
rect 4173 20930 4198 20986
rect 4254 20930 4278 20986
rect 4334 20930 4358 20986
rect 4414 20930 4438 20986
rect 4494 20984 7710 20986
rect 4494 20932 6847 20984
rect 6899 20932 6949 20984
rect 7001 20932 7051 20984
rect 7103 20966 7710 20984
rect 7103 20951 7762 20966
rect 7103 20932 7710 20951
rect 4494 20930 7710 20932
rect 3703 20900 7710 20930
rect 3703 20844 3712 20900
rect 3768 20844 3793 20900
rect 3849 20844 3874 20900
rect 3930 20844 3955 20900
rect 4011 20844 4036 20900
rect 4092 20844 4117 20900
rect 4173 20844 4198 20900
rect 4254 20844 4278 20900
rect 4334 20844 4358 20900
rect 4414 20844 4438 20900
rect 4494 20848 6847 20900
rect 6899 20848 6949 20900
rect 7001 20848 7051 20900
rect 7103 20899 7710 20900
rect 7103 20884 7762 20899
rect 7103 20848 7710 20884
rect 4494 20844 7710 20848
rect 3703 20832 7710 20844
rect 3703 20816 7762 20832
rect 3703 20814 6847 20816
rect 3703 20758 3712 20814
rect 3768 20758 3793 20814
rect 3849 20758 3874 20814
rect 3930 20758 3955 20814
rect 4011 20758 4036 20814
rect 4092 20758 4117 20814
rect 4173 20758 4198 20814
rect 4254 20758 4278 20814
rect 4334 20758 4358 20814
rect 4414 20758 4438 20814
rect 4494 20764 6847 20814
rect 6899 20764 6949 20816
rect 7001 20764 7051 20816
rect 7103 20764 7710 20816
rect 4494 20758 7762 20764
rect 5937 19887 6015 19939
rect 6067 19887 6079 19939
rect 6131 19887 6137 19939
rect 5937 19627 6137 19887
rect 5937 19575 6015 19627
rect 6067 19575 6079 19627
rect 6131 19575 6137 19627
tri 5901 19315 5937 19351 se
rect 5937 19315 6137 19575
rect 6165 19808 8763 19814
rect 6217 19762 8711 19808
rect 6217 19756 6245 19762
tri 6245 19756 6251 19762 nw
tri 8677 19756 8683 19762 ne
rect 8683 19756 8711 19762
rect 6165 19744 6233 19756
tri 6233 19744 6245 19756 nw
tri 8683 19744 8695 19756 ne
rect 8695 19744 8763 19756
tri 6217 19728 6233 19744 nw
tri 8695 19728 8711 19744 ne
rect 6165 19507 6217 19692
rect 8711 19686 8763 19692
rect 7710 19672 7762 19678
rect 7710 19573 7762 19620
rect 6165 19443 6217 19455
rect 6364 19557 6416 19563
tri 6416 19515 6422 19521 sw
rect 7710 19515 7762 19521
rect 6416 19505 6422 19515
rect 6364 19493 6422 19505
rect 6416 19487 6422 19493
tri 6422 19487 6450 19515 sw
rect 6416 19481 8799 19487
rect 6416 19441 8631 19481
rect 6364 19435 8631 19441
tri 8597 19429 8603 19435 ne
rect 8603 19429 8631 19435
rect 8683 19435 8799 19481
rect 8851 19435 8863 19487
rect 8915 19435 8921 19487
tri 8603 19417 8615 19429 ne
rect 8615 19417 8683 19429
tri 8615 19401 8631 19417 ne
rect 6165 19385 6217 19391
tri 8683 19401 8717 19435 nw
rect 8631 19359 8683 19365
tri 5849 19263 5901 19315 se
rect 5901 19263 6015 19315
rect 6067 19263 6079 19315
rect 6131 19263 6137 19315
tri 5805 19219 5849 19263 se
rect 5849 19219 6137 19263
tri 5768 19182 5805 19219 se
rect 5805 19182 6137 19219
tri 5716 19130 5768 19182 se
rect 5768 19130 6137 19182
tri 5715 19129 5716 19130 se
rect 5716 19129 6137 19130
tri 5704 19118 5715 19129 se
rect 5715 19118 6137 19129
tri 5681 19095 5704 19118 se
rect 5704 19095 6137 19118
rect 3321 19039 3712 19095
rect 3768 19039 3793 19095
rect 3849 19039 3874 19095
rect 3930 19039 3955 19095
rect 4011 19039 4036 19095
rect 4092 19039 4117 19095
rect 4173 19039 4198 19095
rect 4254 19039 4278 19095
rect 4334 19039 4358 19095
rect 4414 19039 4438 19095
rect 4494 19039 6137 19095
rect 3321 19003 6137 19039
rect 3321 18951 6015 19003
rect 6067 18951 6079 19003
rect 6131 18951 6137 19003
rect 3321 18895 3712 18951
rect 3768 18895 3793 18951
rect 3849 18895 3874 18951
rect 3930 18895 3955 18951
rect 4011 18895 4036 18951
rect 4092 18895 4117 18951
rect 4173 18895 4198 18951
rect 4254 18895 4278 18951
rect 4334 18895 4358 18951
rect 4414 18895 4438 18951
rect 4494 18895 6137 18951
tri 4966 18886 4975 18895 ne
rect 4975 18886 4987 18895
tri 4975 18874 4987 18886 ne
rect 5039 18886 5051 18895
tri 5051 18886 5060 18895 nw
tri 5681 18888 5688 18895 ne
rect 5688 18888 6137 18895
tri 5688 18886 5690 18888 ne
rect 5690 18886 6137 18888
tri 5039 18874 5051 18886 nw
tri 5690 18874 5702 18886 ne
rect 5702 18874 6137 18886
tri 5702 18834 5742 18874 ne
rect 5742 18834 6137 18874
tri 5742 18822 5754 18834 ne
rect 5754 18822 6137 18834
tri 5754 18780 5796 18822 ne
rect 5796 18780 6137 18822
tri 5237 18770 5247 18780 se
tri 5796 18770 5806 18780 ne
rect 5806 18770 6137 18780
tri 5213 18746 5237 18770 se
rect 5237 18746 5247 18770
tri 5806 18746 5830 18770 ne
rect 5830 18746 6137 18770
rect 6165 19219 8603 19225
rect 6165 19182 8551 19219
rect 6217 19173 8551 19182
rect 6217 19167 6245 19173
tri 6245 19167 6251 19173 nw
tri 8517 19167 8523 19173 ne
rect 8523 19167 8551 19173
rect 6217 19155 6233 19167
tri 6233 19155 6245 19167 nw
tri 8523 19155 8535 19167 ne
rect 8535 19155 8603 19167
tri 6217 19139 6233 19155 nw
tri 8535 19139 8551 19155 ne
rect 6165 19118 6217 19130
rect 8551 19097 8603 19103
rect 6165 18886 6217 19066
rect 6364 19089 6416 19095
tri 6359 19037 6364 19042 se
rect 8471 19089 8523 19095
tri 6416 19042 6427 19053 sw
tri 8460 19042 8471 19053 se
rect 6416 19037 6427 19042
tri 6427 19037 6432 19042 sw
tri 8455 19037 8460 19042 se
rect 8460 19037 8471 19042
tri 6347 19025 6359 19037 se
rect 6359 19025 6432 19037
tri 6432 19025 6444 19037 sw
tri 8443 19025 8455 19037 se
rect 8455 19025 8523 19037
tri 6341 19019 6347 19025 se
rect 6347 19019 6364 19025
tri 6319 18997 6341 19019 se
rect 6341 18997 6364 19019
tri 6295 18973 6319 18997 se
rect 6319 18973 6364 18997
rect 6416 19019 6444 19025
tri 6444 19019 6450 19025 sw
tri 8437 19019 8443 19025 se
rect 8443 19019 8471 19025
rect 6416 18973 8471 19019
rect 6165 18822 6217 18834
rect 6165 18764 6217 18770
tri 6245 18923 6295 18973 se
rect 6295 18967 8523 18973
rect 6295 18923 6319 18967
tri 6319 18923 6363 18967 nw
tri 5830 18740 5836 18746 ne
rect 5836 18740 6137 18746
tri 5836 18734 5842 18740 ne
rect 5842 18734 6137 18740
tri 5842 18691 5885 18734 ne
rect 5885 18691 6137 18734
tri 5885 18639 5937 18691 ne
rect 5937 18639 6015 18691
rect 6067 18639 6079 18691
rect 6131 18639 6137 18691
rect 6245 18562 6297 18923
tri 6297 18901 6319 18923 nw
rect 7524 18882 9146 18888
rect 7524 18856 9005 18882
rect 7576 18830 9005 18856
rect 9057 18830 9093 18882
rect 9145 18830 9146 18882
rect 7576 18804 9146 18830
rect 7524 18792 9146 18804
rect 7576 18740 9005 18792
rect 9057 18740 9093 18792
rect 9145 18740 9146 18792
rect 7524 18734 9146 18740
rect 6245 18498 6297 18510
rect 6364 18625 8443 18631
rect 6416 18579 8391 18625
rect 6416 18573 6444 18579
tri 6444 18573 6450 18579 nw
tri 8357 18573 8363 18579 ne
rect 8363 18573 8391 18579
rect 6364 18561 6432 18573
tri 6432 18561 6444 18573 nw
tri 8363 18561 8375 18573 ne
rect 8375 18561 8443 18573
tri 6416 18545 6432 18561 nw
tri 8375 18545 8391 18561 ne
rect 6364 18503 6416 18509
rect 8391 18503 8443 18509
rect 3833 18436 3839 18488
rect 3891 18436 3924 18488
rect 3976 18436 4009 18488
rect 4061 18436 4093 18488
rect 4145 18436 4177 18488
rect 4229 18446 5185 18488
tri 5185 18446 5227 18488 sw
rect 4229 18436 5227 18446
rect 3833 18408 5227 18436
rect 3833 18356 3839 18408
rect 3891 18356 3924 18408
rect 3976 18356 4009 18408
rect 4061 18356 4093 18408
rect 4145 18356 4177 18408
rect 4229 18356 5227 18408
tri 5227 18356 5317 18446 sw
rect 6245 18440 6297 18446
tri 5131 18323 5164 18356 ne
rect 5164 18323 5317 18356
tri 5317 18323 5350 18356 sw
tri 5164 18317 5170 18323 ne
rect 5170 18317 5350 18323
tri 5350 18317 5356 18323 sw
rect 7618 18317 7670 18323
tri 5170 18265 5222 18317 ne
rect 5222 18265 5356 18317
tri 5356 18265 5408 18317 sw
tri 5222 18262 5225 18265 ne
rect 5225 18262 5408 18265
tri 5408 18262 5411 18265 sw
tri 5225 18253 5234 18262 ne
rect 5234 18253 5832 18262
tri 5234 18201 5286 18253 ne
rect 5286 18206 5832 18253
rect 5888 18206 5914 18262
rect 5970 18206 5995 18262
rect 6051 18206 6076 18262
rect 6132 18206 6157 18262
rect 6213 18206 6238 18262
rect 6294 18206 6319 18262
rect 6375 18206 6400 18262
rect 6456 18206 6481 18262
rect 6537 18206 6562 18262
rect 6618 18206 6627 18262
rect 5286 18201 6627 18206
tri 5286 18189 5298 18201 ne
rect 5298 18189 6627 18201
rect 7618 18253 7670 18265
tri 7670 18247 7704 18281 sw
rect 7670 18241 8283 18247
rect 7670 18201 8231 18241
rect 7618 18195 8231 18201
tri 8197 18189 8203 18195 ne
rect 8203 18189 8231 18195
tri 5298 18177 5310 18189 ne
rect 5310 18182 6627 18189
rect 5310 18177 5832 18182
tri 5310 18170 5317 18177 ne
rect 5317 18170 5832 18177
tri 5317 18126 5361 18170 ne
rect 5361 18126 5832 18170
rect 5888 18126 5914 18182
rect 5970 18126 5995 18182
rect 6051 18126 6076 18182
rect 6132 18126 6157 18182
rect 6213 18126 6238 18182
rect 6294 18126 6319 18182
rect 6375 18126 6400 18182
rect 6456 18126 6481 18182
rect 6537 18126 6562 18182
rect 6618 18126 6627 18182
tri 8203 18177 8215 18189 ne
rect 8215 18177 8283 18189
tri 8215 18161 8231 18177 ne
rect 8231 18119 8283 18125
rect 7616 18045 7962 18051
rect 7668 17993 7910 18045
rect 7616 17981 7962 17993
rect 7668 17929 7910 17981
rect 7616 17923 7962 17929
rect 8910 17403 8921 17463
rect 3703 17280 3712 17336
rect 3768 17280 3793 17336
rect 3849 17280 3874 17336
rect 3930 17280 3955 17336
rect 4011 17280 4036 17336
rect 4092 17280 4117 17336
rect 4173 17280 4198 17336
rect 4254 17280 4278 17336
rect 4334 17280 4358 17336
rect 4414 17280 4438 17336
rect 4494 17330 7104 17336
rect 4494 17280 6847 17330
rect 3703 17278 6847 17280
rect 6899 17278 6915 17330
rect 6967 17278 6983 17330
rect 7035 17278 7051 17330
rect 7103 17278 7104 17330
rect 3703 17263 7104 17278
rect 3703 17250 6847 17263
rect 3703 17194 3712 17250
rect 3768 17194 3793 17250
rect 3849 17194 3874 17250
rect 3930 17194 3955 17250
rect 4011 17194 4036 17250
rect 4092 17194 4117 17250
rect 4173 17194 4198 17250
rect 4254 17194 4278 17250
rect 4334 17194 4358 17250
rect 4414 17194 4438 17250
rect 4494 17211 6847 17250
rect 6899 17211 6915 17263
rect 6967 17211 6983 17263
rect 7035 17211 7051 17263
rect 7103 17211 7104 17263
rect 4494 17196 7104 17211
rect 4494 17194 6847 17196
rect 3703 17164 6847 17194
rect 3703 17108 3712 17164
rect 3768 17108 3793 17164
rect 3849 17108 3874 17164
rect 3930 17108 3955 17164
rect 4011 17108 4036 17164
rect 4092 17108 4117 17164
rect 4173 17108 4198 17164
rect 4254 17108 4278 17164
rect 4334 17108 4358 17164
rect 4414 17108 4438 17164
rect 4494 17144 6847 17164
rect 6899 17144 6915 17196
rect 6967 17144 6983 17196
rect 7035 17144 7051 17196
rect 7103 17144 7104 17196
rect 4494 17129 7104 17144
rect 4494 17108 6847 17129
rect 3703 17078 6847 17108
rect 3703 17022 3712 17078
rect 3768 17022 3793 17078
rect 3849 17022 3874 17078
rect 3930 17022 3955 17078
rect 4011 17022 4036 17078
rect 4092 17022 4117 17078
rect 4173 17022 4198 17078
rect 4254 17022 4278 17078
rect 4334 17022 4358 17078
rect 4414 17022 4438 17078
rect 4494 17077 6847 17078
rect 6899 17077 6915 17129
rect 6967 17077 6983 17129
rect 7035 17077 7051 17129
rect 7103 17077 7104 17129
rect 4494 17062 7104 17077
rect 4494 17022 6847 17062
rect 3703 17010 6847 17022
rect 6899 17010 6915 17062
rect 6967 17010 6983 17062
rect 7035 17010 7051 17062
rect 7103 17010 7104 17062
rect 3703 16994 7104 17010
rect 3703 16992 6847 16994
rect 3703 16936 3712 16992
rect 3768 16936 3793 16992
rect 3849 16936 3874 16992
rect 3930 16936 3955 16992
rect 4011 16936 4036 16992
rect 4092 16936 4117 16992
rect 4173 16936 4198 16992
rect 4254 16936 4278 16992
rect 4334 16936 4358 16992
rect 4414 16936 4438 16992
rect 4494 16942 6847 16992
rect 6899 16942 6915 16994
rect 6967 16942 6983 16994
rect 7035 16942 7051 16994
rect 7103 16942 7104 16994
rect 7524 17076 9391 17108
rect 7576 17056 9391 17076
rect 9443 17056 9486 17108
rect 9538 17056 9544 17108
rect 7576 17024 9544 17056
rect 7524 17012 9544 17024
rect 7576 17006 9544 17012
rect 7576 16960 9391 17006
rect 7524 16954 9391 16960
rect 9443 16954 9486 17006
rect 9538 16954 9544 17006
rect 4494 16936 7104 16942
rect 7618 16741 8363 16747
rect 7618 16715 8311 16741
rect 7670 16689 8311 16715
rect 7670 16663 8363 16689
rect 7618 16651 8363 16663
rect 7670 16599 8311 16651
rect 7618 16593 8363 16599
rect 2654 16222 7667 16228
rect 2706 16176 6818 16222
rect 2706 16170 2734 16176
tri 2734 16170 2740 16176 nw
tri 6784 16170 6790 16176 ne
rect 6790 16170 6818 16176
rect 6870 16176 7615 16222
rect 6870 16170 6898 16176
tri 6898 16170 6904 16176 nw
tri 7581 16170 7587 16176 ne
rect 7587 16170 7615 16176
rect 2654 16158 2722 16170
tri 2722 16158 2734 16170 nw
tri 6790 16158 6802 16170 ne
rect 6802 16158 6886 16170
tri 6886 16158 6898 16170 nw
tri 7587 16158 7599 16170 ne
rect 7599 16158 7667 16170
tri 2706 16142 2722 16158 nw
tri 6802 16142 6818 16158 ne
rect 2654 16100 2706 16106
tri 6870 16142 6886 16158 nw
tri 7599 16142 7615 16158 ne
rect 6818 16100 6870 16106
rect 7615 16100 7667 16106
rect 7910 15792 7962 15798
tri 7894 15740 7910 15756 se
tri 7882 15728 7894 15740 se
rect 7894 15728 7962 15740
tri 7876 15722 7882 15728 se
rect 7882 15722 7910 15728
rect 1648 15716 7910 15722
rect 1700 15676 7910 15716
rect 1700 15670 7962 15676
rect 1648 15652 1700 15664
tri 1700 15636 1734 15670 nw
rect 1648 15594 1700 15600
rect 7508 15589 10191 15598
rect 7508 15581 10135 15589
rect 7560 15533 10135 15581
rect 7560 15529 10191 15533
rect 7508 15517 10191 15529
rect 7560 15509 10191 15517
rect 7560 15465 10135 15509
rect 7508 15453 10135 15465
rect 7508 15444 10191 15453
rect 770 15319 9624 15371
tri 740 14195 770 14225 se
rect 770 14195 846 15319
tri 846 15285 880 15319 nw
tri 9538 15285 9572 15319 ne
rect 3703 15221 7104 15223
rect 3703 15165 3712 15221
rect 3768 15165 3793 15221
rect 3849 15165 3874 15221
rect 3930 15165 3955 15221
rect 4011 15165 4036 15221
rect 4092 15165 4117 15221
rect 4173 15165 4198 15221
rect 3703 15141 4198 15165
rect 3703 15085 3712 15141
rect 3768 15085 3793 15141
rect 3849 15085 3874 15141
rect 3930 15085 3955 15141
rect 4011 15085 4036 15141
rect 4092 15085 4117 15141
rect 4173 15085 4198 15141
rect 3703 15061 4198 15085
rect 3703 15005 3712 15061
rect 3768 15005 3793 15061
rect 3849 15005 3874 15061
rect 3930 15005 3955 15061
rect 4011 15005 4036 15061
rect 4092 15005 4117 15061
rect 4173 15005 4198 15061
rect 3703 14981 4198 15005
rect 3703 14925 3712 14981
rect 3768 14925 3793 14981
rect 3849 14925 3874 14981
rect 3930 14925 3955 14981
rect 4011 14925 4036 14981
rect 4092 14925 4117 14981
rect 4173 14925 4198 14981
rect 4494 15217 7104 15221
rect 4494 15165 6738 15217
rect 6790 15165 6944 15217
rect 6996 15165 7052 15217
rect 4494 15139 7104 15165
rect 4494 15087 6738 15139
rect 6790 15087 6944 15139
rect 6996 15087 7052 15139
rect 4494 15060 7104 15087
rect 4494 15008 6738 15060
rect 6790 15008 6944 15060
rect 6996 15008 7052 15060
rect 4494 14981 7104 15008
rect 4494 14929 6738 14981
rect 6790 14929 6944 14981
rect 6996 14929 7052 14981
rect 4494 14925 7104 14929
rect 3703 14923 7104 14925
rect 9005 15034 9145 15040
rect 9057 14982 9093 15034
rect 9005 14945 9145 14982
rect 7618 14902 8203 14908
rect 7618 14876 8149 14902
rect 7670 14850 8149 14876
rect 8201 14850 8203 14902
rect 7670 14824 8203 14850
rect 7618 14812 8203 14824
rect 7670 14760 8149 14812
rect 8201 14760 8203 14812
rect 7618 14754 8203 14760
rect 9057 14893 9093 14945
rect 2661 14611 5858 14625
rect 2661 14555 2670 14611
rect 2726 14555 2751 14611
rect 2807 14555 2832 14611
rect 2888 14555 2913 14611
rect 2969 14555 2994 14611
rect 3050 14555 3075 14611
rect 3131 14555 3156 14611
rect 3212 14555 3237 14611
rect 3293 14555 3318 14611
rect 3374 14555 3398 14611
rect 3454 14555 3478 14611
rect 3534 14610 5858 14611
tri 5858 14610 5873 14625 sw
rect 9005 14610 9145 14893
rect 9385 15007 9391 15059
rect 9443 15007 9486 15059
rect 9538 15007 9544 15059
rect 9385 14991 9544 15007
rect 9385 14939 9391 14991
rect 9443 14939 9486 14991
rect 9538 14939 9544 14991
rect 3534 14558 5873 14610
tri 5873 14558 5925 14610 sw
rect 9005 14558 9011 14610
rect 9063 14558 9087 14610
rect 9139 14558 9145 14610
rect 9199 14746 9219 14798
rect 9271 14746 9283 14798
rect 9335 14746 9353 14798
rect 9199 14567 9353 14746
rect 3534 14555 5925 14558
rect 2661 14541 5925 14555
tri 5925 14541 5942 14558 sw
rect 2661 14528 5942 14541
tri 5942 14528 5955 14541 sw
rect 9005 14528 9145 14558
rect 2661 14527 5955 14528
rect 2661 14471 2670 14527
rect 2726 14471 2751 14527
rect 2807 14471 2832 14527
rect 2888 14471 2913 14527
rect 2969 14471 2994 14527
rect 3050 14471 3075 14527
rect 3131 14471 3156 14527
rect 3212 14471 3237 14527
rect 3293 14471 3318 14527
rect 3374 14471 3398 14527
rect 3454 14471 3478 14527
rect 3534 14476 5955 14527
tri 5955 14476 6007 14528 sw
rect 9005 14476 9011 14528
rect 9063 14476 9087 14528
rect 9139 14476 9145 14528
rect 3534 14471 6007 14476
rect 2661 14466 6007 14471
tri 6007 14466 6017 14476 sw
rect 9005 14475 9145 14476
rect 9385 14541 9544 14939
rect 9572 14792 9624 15319
rect 9572 14724 9624 14740
rect 9572 14656 9624 14672
rect 9572 14598 9624 14604
rect 9385 14489 9391 14541
rect 9443 14489 9486 14541
rect 9538 14489 9544 14541
rect 2661 14459 6017 14466
tri 6017 14459 6024 14466 sw
rect 9385 14459 9544 14489
rect 9890 14466 9942 14472
rect 2661 14443 6024 14459
rect 2661 14387 2670 14443
rect 2726 14387 2751 14443
rect 2807 14387 2832 14443
rect 2888 14387 2913 14443
rect 2969 14387 2994 14443
rect 3050 14387 3075 14443
rect 3131 14387 3156 14443
rect 3212 14387 3237 14443
rect 3293 14387 3318 14443
rect 3374 14387 3398 14443
rect 3454 14387 3478 14443
rect 3534 14430 6024 14443
tri 6024 14430 6053 14459 sw
rect 3534 14417 6053 14430
tri 6053 14417 6066 14430 sw
tri 9877 14417 9890 14430 se
rect 3534 14414 6066 14417
tri 6066 14414 6069 14417 sw
rect 7615 14414 7667 14417
tri 7667 14414 7670 14417 sw
tri 9874 14414 9877 14417 se
rect 9877 14414 9890 14417
rect 3534 14411 6069 14414
tri 6069 14411 6072 14414 sw
rect 7615 14411 7670 14414
rect 3534 14387 6072 14411
rect 2661 14359 6072 14387
tri 6072 14359 6124 14411 sw
rect 7667 14402 7670 14411
tri 7670 14402 7682 14414 sw
tri 9862 14402 9874 14414 se
rect 9874 14402 9942 14414
rect 7667 14396 7682 14402
tri 7682 14396 7688 14402 sw
tri 9856 14396 9862 14402 se
rect 9862 14396 9890 14402
rect 7667 14359 9890 14396
rect 2661 14350 6124 14359
tri 6124 14350 6133 14359 sw
rect 7615 14350 9890 14359
rect 2661 14347 6133 14350
tri 6133 14347 6136 14350 sw
rect 7615 14347 9942 14350
rect 2661 14295 6136 14347
tri 6136 14295 6188 14347 sw
rect 7667 14344 9942 14347
tri 7667 14310 7701 14344 nw
rect 2661 14289 6188 14295
tri 6188 14289 6194 14295 sw
rect 7615 14289 7667 14295
rect 2661 14261 6194 14289
tri 6194 14261 6222 14289 sw
rect 2661 14255 10828 14261
rect 2661 14251 10710 14255
tri 5619 14247 5623 14251 ne
rect 5623 14247 10710 14251
tri 5623 14225 5645 14247 ne
rect 5645 14225 5983 14247
tri 846 14195 876 14225 sw
tri 5645 14195 5675 14225 ne
rect 5675 14195 5983 14225
rect 6035 14195 6065 14247
rect 6117 14195 6147 14247
rect 6199 14195 6228 14247
rect 6280 14195 6309 14247
rect 6361 14241 10710 14247
rect 6361 14195 9199 14241
tri 736 14191 740 14195 se
rect 740 14191 876 14195
tri 876 14191 880 14195 sw
tri 5675 14191 5679 14195 ne
rect 5679 14191 7197 14195
rect 736 14139 742 14191
rect 794 14139 806 14191
rect 858 14139 2210 14191
rect 2262 14139 2274 14191
rect 2326 14139 2961 14191
rect 3013 14139 3027 14191
rect 3079 14139 3085 14191
tri 5679 14151 5719 14191 ne
rect 5719 14151 7197 14191
tri 5719 14139 5731 14151 ne
rect 5731 14139 5983 14151
tri 5731 14111 5759 14139 ne
rect 5759 14111 5983 14139
rect 1011 14059 1017 14111
rect 1069 14059 1081 14111
rect 1133 14059 3201 14111
tri 5759 14099 5771 14111 ne
rect 5771 14099 5983 14111
rect 6035 14099 6065 14151
rect 6117 14099 6147 14151
rect 6199 14099 6228 14151
rect 6280 14099 6309 14151
rect 6361 14143 7197 14151
rect 7249 14143 7263 14195
rect 7315 14143 7329 14195
rect 7381 14143 7394 14195
rect 7446 14189 9199 14195
rect 9251 14189 9301 14241
rect 9353 14189 9732 14241
rect 9784 14189 9808 14241
rect 9860 14203 10710 14241
rect 10762 14203 10776 14255
rect 9860 14189 10828 14203
rect 7446 14158 10828 14189
rect 7446 14151 10710 14158
rect 7446 14143 9199 14151
rect 6361 14125 9199 14143
rect 6361 14099 7197 14125
tri 5771 14073 5797 14099 ne
rect 5797 14073 7197 14099
rect 7249 14073 7263 14125
rect 7315 14073 7329 14125
rect 7381 14073 7394 14125
rect 7446 14099 9199 14125
rect 9251 14099 9301 14151
rect 9353 14099 9732 14151
rect 9784 14099 9808 14151
rect 9860 14106 10710 14151
rect 10762 14106 10776 14158
rect 9860 14099 10828 14106
rect 7446 14073 10828 14099
tri 5797 14061 5809 14073 ne
rect 5809 14061 10828 14073
tri 5809 14059 5811 14061 ne
rect 5811 14059 9199 14061
tri 5811 14055 5815 14059 ne
rect 5815 14055 9199 14059
tri 5815 14031 5839 14055 ne
rect 5839 14031 5983 14055
rect 1184 14025 1654 14031
rect 1236 13979 1654 14025
rect 1706 13979 1718 14031
rect 1770 13979 3107 14031
tri 5839 14003 5867 14031 ne
rect 5867 14003 5983 14031
rect 6035 14003 6065 14055
rect 6117 14003 6147 14055
rect 6199 14003 6228 14055
rect 6280 14003 6309 14055
rect 6361 14003 7197 14055
rect 7249 14003 7263 14055
rect 7315 14003 7329 14055
rect 7381 14003 7394 14055
rect 7446 14009 9199 14055
rect 9251 14009 9301 14061
rect 9353 14009 9732 14061
rect 9784 14009 9808 14061
rect 9860 14009 10710 14061
rect 10762 14009 10776 14061
rect 7446 14003 10828 14009
rect 1184 13961 1236 13973
tri 1236 13945 1270 13979 nw
tri 3061 13945 3095 13979 ne
rect 1184 13903 1236 13909
rect 6501 13930 8717 13936
rect 6553 13884 8717 13930
rect 8769 13884 8781 13936
rect 8833 13884 8839 13936
rect 6553 13878 6559 13884
rect 6501 13866 6559 13878
rect 1579 13795 1585 13847
rect 1637 13795 1649 13847
rect 1701 13795 3342 13847
rect 3394 13795 3406 13847
rect 3458 13795 3464 13847
rect 6553 13856 6559 13866
tri 6559 13856 6587 13884 nw
tri 6553 13850 6559 13856 nw
rect 7715 13850 9011 13856
rect 792 13701 844 13707
rect 1635 13666 1641 13718
rect 1693 13666 1705 13718
rect 1757 13666 3335 13718
rect 3387 13666 3399 13718
rect 3451 13666 3457 13718
tri 844 13657 852 13665 sw
rect 844 13649 852 13657
rect 792 13637 852 13649
rect 844 13631 852 13637
tri 852 13631 878 13657 sw
rect 844 13585 2838 13631
rect 792 13579 2838 13585
rect 6501 13621 6553 13814
rect 7767 13804 9011 13850
rect 9063 13804 9087 13856
rect 9139 13804 9163 13856
rect 9215 13804 9221 13856
rect 7715 13786 7767 13798
tri 7767 13770 7801 13804 nw
rect 7715 13728 7767 13734
rect 8391 13733 8443 13739
tri 8375 13681 8391 13697 se
rect 8631 13733 8683 13739
tri 8443 13681 8459 13697 sw
tri 8615 13681 8631 13697 se
tri 8363 13669 8375 13681 se
rect 8375 13669 8459 13681
tri 8459 13669 8471 13681 sw
tri 8603 13669 8615 13681 se
rect 8615 13669 8683 13681
tri 8359 13665 8363 13669 se
rect 8363 13665 8391 13669
tri 8357 13663 8359 13665 se
rect 8359 13663 8391 13665
rect 6501 13557 6553 13569
rect 931 13497 3140 13503
rect 983 13451 3140 13497
rect 3192 13451 3204 13503
rect 3256 13451 3262 13503
tri 3571 13455 3573 13457 se
rect 3573 13455 3625 13530
rect 6661 13657 8391 13663
rect 6713 13617 8391 13657
rect 8443 13663 8471 13669
tri 8471 13663 8477 13669 sw
tri 8597 13663 8603 13669 se
rect 8603 13663 8631 13669
rect 8443 13617 8631 13663
rect 6713 13611 8683 13617
rect 6661 13593 6713 13605
tri 6713 13577 6747 13611 nw
rect 6661 13535 6713 13541
rect 6933 13571 9391 13577
rect 6501 13499 6553 13505
rect 6985 13525 9391 13571
rect 9443 13525 9486 13577
rect 9538 13525 9544 13577
rect 6985 13519 9544 13525
rect 6933 13507 9544 13519
tri 3625 13461 3659 13495 nw
tri 3567 13451 3571 13455 se
rect 3571 13451 3625 13455
rect 983 13449 1015 13451
tri 1015 13449 1017 13451 nw
tri 3565 13449 3567 13451 se
rect 3567 13449 3625 13451
rect 6985 13501 9544 13507
rect 6985 13455 9391 13501
rect 6933 13449 9391 13455
rect 9443 13449 9486 13501
rect 9538 13449 9544 13501
rect 983 13445 989 13449
rect 931 13433 989 13445
rect 983 13423 989 13433
tri 989 13423 1015 13449 nw
tri 3539 13423 3565 13449 se
rect 3565 13423 3625 13449
tri 983 13417 989 13423 nw
rect 931 13375 983 13381
rect 1691 13371 1697 13423
rect 1749 13371 1761 13423
rect 1813 13371 3625 13423
tri 9351 13415 9385 13449 ne
rect 6501 13378 8815 13384
rect 1775 13291 1781 13343
rect 1833 13291 1845 13343
rect 1897 13291 3625 13343
tri 3539 13290 3540 13291 ne
rect 3540 13290 3625 13291
tri 3540 13263 3567 13290 ne
rect 3567 13263 3625 13290
rect 1903 13211 1937 13263
rect 1989 13211 2001 13263
rect 2053 13211 3457 13263
tri 3567 13257 3573 13263 ne
tri 3295 13202 3304 13211 ne
rect 3304 13202 3457 13211
rect 1299 13196 1351 13202
tri 3304 13193 3313 13202 ne
rect 3313 13193 3457 13202
tri 3313 13187 3319 13193 ne
rect 3319 13187 3335 13193
tri 3319 13183 3323 13187 ne
rect 3323 13183 3335 13187
rect 1299 13132 1351 13144
tri 1351 13131 1357 13137 sw
rect 1423 13131 1429 13183
rect 1481 13131 1493 13183
rect 1545 13131 3140 13183
rect 3192 13131 3204 13183
rect 3256 13131 3262 13183
tri 3323 13177 3329 13183 ne
rect 3329 13141 3335 13183
rect 3387 13141 3399 13193
rect 3451 13141 3457 13193
rect 3573 13200 3625 13263
rect 6501 13332 8551 13378
rect 6501 13326 6581 13332
tri 6581 13326 6587 13332 nw
tri 8517 13326 8523 13332 ne
rect 8523 13326 8551 13332
rect 8603 13332 8763 13378
rect 8603 13326 8631 13332
tri 8631 13326 8637 13332 nw
tri 8729 13326 8735 13332 ne
rect 8735 13326 8763 13332
rect 6501 13314 6569 13326
tri 6569 13314 6581 13326 nw
tri 8523 13314 8535 13326 ne
rect 8535 13314 8619 13326
tri 8619 13314 8631 13326 nw
tri 8735 13314 8747 13326 ne
rect 8747 13314 8815 13326
rect 6501 13295 6553 13314
tri 6553 13298 6569 13314 nw
tri 8535 13304 8545 13314 ne
rect 8545 13304 8551 13314
rect 6821 13298 6873 13304
tri 8545 13298 8551 13304 ne
rect 6501 13231 6553 13243
tri 3625 13200 3646 13221 sw
rect 3573 13187 3646 13200
tri 3646 13187 3659 13200 sw
rect 3573 13184 3625 13187
tri 6873 13284 6879 13290 sw
rect 6873 13278 6879 13284
tri 6879 13278 6885 13284 sw
tri 8305 13278 8311 13284 se
rect 8311 13278 8363 13284
rect 6873 13256 6885 13278
tri 6885 13256 6907 13278 sw
tri 8283 13256 8305 13278 se
rect 8305 13256 8311 13278
rect 6873 13246 8311 13256
rect 6821 13234 8311 13246
rect 1351 13103 1357 13131
tri 1357 13103 1385 13131 sw
rect 1351 13080 2838 13103
rect 1299 13051 2838 13080
rect 2180 12964 2186 13016
rect 2238 12964 2274 13016
rect 2326 12964 2868 13016
rect 2920 12964 2934 13016
rect 2986 12964 2992 13016
rect 6501 13004 6553 13179
rect 6661 13198 6713 13204
rect 6873 13226 8311 13234
tri 8603 13298 8619 13314 nw
tri 8747 13298 8763 13314 ne
rect 8551 13256 8603 13262
rect 8763 13256 8815 13262
rect 6873 13214 8363 13226
rect 6873 13200 8311 13214
rect 6821 13176 6873 13182
tri 6873 13176 6897 13200 nw
tri 8277 13176 8301 13200 ne
rect 8301 13176 8311 13200
tri 8301 13166 8311 13176 ne
tri 6713 13156 6719 13162 sw
rect 8311 13156 8363 13162
rect 6713 13146 6719 13156
rect 6661 13141 6719 13146
tri 6719 13141 6734 13156 sw
tri 6657 13137 6661 13141 se
rect 6661 13137 6734 13141
tri 6654 13134 6657 13137 se
rect 6657 13134 6734 13137
tri 6648 13128 6654 13134 se
rect 6654 13128 6661 13134
tri 6623 13103 6648 13128 se
rect 6648 13103 6661 13128
tri 6602 13082 6623 13103 se
rect 6623 13082 6661 13103
rect 6713 13128 6734 13134
tri 6734 13128 6747 13141 sw
rect 6713 13122 8523 13128
rect 6713 13082 8471 13122
tri 6596 13076 6602 13082 se
rect 6602 13076 8471 13082
tri 6590 13070 6596 13076 se
rect 6596 13070 6664 13076
tri 6664 13070 6670 13076 nw
tri 8437 13070 8443 13076 ne
rect 8443 13070 8471 13076
rect 6501 12940 6553 12952
rect 1859 12835 1865 12887
rect 1917 12835 1929 12887
rect 1981 12835 3342 12887
rect 3394 12835 3406 12887
rect 3458 12835 3464 12887
rect 6501 12882 6553 12888
tri 6581 13061 6590 13070 se
rect 6590 13061 6655 13070
tri 6655 13061 6664 13070 nw
tri 8443 13061 8452 13070 ne
rect 8452 13061 8523 13070
rect 6581 13058 6652 13061
tri 6652 13058 6655 13061 nw
tri 8452 13058 8455 13061 ne
rect 8455 13058 8523 13061
rect 6581 13054 6648 13058
tri 6648 13054 6652 13058 nw
tri 8455 13054 8459 13058 ne
rect 8459 13054 8471 13058
rect 6581 13051 6645 13054
tri 6645 13051 6648 13054 nw
tri 8459 13051 8462 13054 ne
rect 8462 13051 8471 13054
rect 6581 13048 6642 13051
tri 6642 13048 6645 13051 nw
tri 8462 13048 8465 13051 ne
rect 8465 13048 8471 13051
rect 6581 13042 6636 13048
tri 6636 13042 6642 13048 nw
rect 7809 13042 7861 13048
tri 8465 13044 8469 13048 ne
rect 8469 13044 8471 13048
tri 8469 13042 8471 13044 ne
rect 1491 12825 1543 12831
rect 1491 12761 1543 12773
rect 2654 12773 2706 12779
tri 1543 12721 1559 12737 sw
tri 2638 12721 2654 12737 se
tri 2706 12721 2722 12737 sw
tri 3079 12721 3095 12737 se
rect 1543 12709 1559 12721
tri 1559 12709 1571 12721 sw
tri 2626 12709 2638 12721 se
rect 2638 12709 2722 12721
rect 1491 12703 1571 12709
tri 1571 12703 1577 12709 sw
tri 2620 12703 2626 12709 se
rect 2626 12703 2654 12709
tri 1491 12677 1517 12703 ne
rect 1517 12657 2654 12703
rect 2706 12703 2722 12709
tri 2722 12703 2740 12721 sw
tri 3061 12703 3079 12721 se
rect 3079 12703 3095 12721
rect 6581 12721 6633 13042
tri 6633 13039 6636 13042 nw
tri 9351 13044 9385 13078 se
rect 9385 13044 9544 13449
rect 7809 12986 7861 12990
tri 7861 12986 7881 13006 sw
rect 8471 13000 8523 13006
rect 8570 13038 9391 13044
rect 8622 12986 8646 13038
rect 8698 12992 9391 13038
rect 9443 12992 9486 13044
rect 9538 12992 9544 13044
rect 8698 12986 9544 12992
rect 7809 12978 7881 12986
rect 7861 12972 7881 12978
tri 7881 12972 7895 12986 sw
rect 7861 12926 8237 12972
rect 7809 12920 8237 12926
rect 8289 12920 8301 12972
rect 8353 12920 8359 12972
rect 8570 12953 9544 12986
rect 8622 12901 8646 12953
rect 8698 12948 9544 12953
rect 8698 12901 9391 12948
rect 8570 12896 9391 12901
rect 9443 12896 9486 12948
rect 9538 12896 9544 12948
rect 8570 12895 9544 12896
rect 8391 12819 8443 12825
tri 8387 12779 8391 12783 se
tri 8375 12767 8387 12779 se
rect 8387 12767 8391 12779
tri 8363 12755 8375 12767 se
rect 8375 12755 8443 12767
tri 8357 12749 8363 12755 se
rect 8363 12749 8391 12755
rect 2706 12657 3107 12703
rect 1517 12651 3107 12657
rect 6581 12657 6633 12669
rect 1435 12571 3201 12623
rect 6661 12743 8391 12749
rect 6713 12703 8391 12743
rect 6713 12697 8443 12703
rect 6713 12691 6719 12697
rect 6661 12679 6719 12691
rect 6713 12669 6719 12679
tri 6719 12669 6747 12697 nw
tri 6713 12663 6719 12669 nw
rect 6661 12621 6713 12627
rect 6770 12660 10191 12669
rect 6770 12625 10135 12660
rect 6581 12599 6633 12605
rect 1435 12569 1519 12571
tri 1519 12569 1521 12571 nw
rect 6770 12569 6779 12625
rect 6835 12569 6859 12625
rect 6915 12604 10135 12625
rect 6915 12569 10191 12604
rect 1435 12565 1489 12569
rect 1487 12539 1489 12565
tri 1489 12539 1519 12569 nw
tri 10101 12539 10131 12569 ne
rect 10131 12539 10191 12569
tri 1487 12537 1489 12539 nw
rect 1435 12501 1487 12513
rect 1435 12443 1487 12449
rect 6536 12512 9862 12539
tri 10131 12535 10135 12539 ne
rect 10135 12536 10191 12539
rect 6536 12460 6542 12512
rect 6594 12460 6608 12512
rect 6660 12460 6674 12512
rect 6726 12460 6740 12512
rect 6792 12460 6806 12512
rect 6858 12460 6872 12512
rect 6924 12460 6938 12512
rect 6990 12460 7004 12512
rect 7056 12460 7070 12512
rect 7122 12460 7136 12512
rect 7188 12460 7202 12512
rect 7254 12460 7268 12512
rect 7320 12460 7334 12512
rect 7386 12460 7400 12512
rect 7452 12460 7466 12512
rect 7518 12460 7532 12512
rect 7584 12460 7598 12512
rect 7650 12460 7664 12512
rect 7716 12460 7729 12512
rect 7781 12460 7794 12512
rect 7846 12460 7859 12512
rect 7911 12460 9738 12512
rect 9790 12460 9804 12512
rect 9856 12460 9862 12512
rect 10135 12471 10191 12480
rect 6536 12433 9862 12460
rect 5906 12349 9342 12401
rect 9394 12349 9406 12401
rect 9458 12349 9464 12401
tri 9573 12366 9579 12372 se
rect 9579 12366 9942 12372
tri 9556 12349 9573 12366 se
rect 9573 12349 9890 12366
tri 9528 12321 9556 12349 se
rect 9556 12321 9890 12349
rect 6008 12269 9232 12321
rect 9284 12269 9296 12321
rect 9348 12320 9890 12321
rect 9348 12314 9595 12320
tri 9595 12314 9601 12320 nw
tri 9856 12314 9862 12320 ne
rect 9862 12314 9890 12320
rect 9348 12302 9583 12314
tri 9583 12302 9595 12314 nw
tri 9862 12302 9874 12314 ne
rect 9874 12302 9942 12314
rect 9348 12269 9550 12302
tri 9550 12269 9583 12302 nw
tri 9874 12286 9890 12302 ne
rect 6012 12262 6039 12269
tri 6039 12262 6046 12269 nw
tri 6426 12262 6433 12269 ne
rect 6433 12262 6615 12269
tri 6615 12262 6622 12269 nw
rect 9652 12262 9704 12268
tri 6012 12235 6039 12262 nw
tri 6433 12235 6460 12262 ne
rect 6460 12244 6597 12262
tri 6597 12244 6615 12262 nw
rect 6460 12217 6588 12244
tri 6588 12235 6597 12244 nw
rect 6460 12165 6466 12217
rect 6518 12165 6530 12217
rect 6582 12165 6588 12217
tri 9618 12192 9652 12226 se
rect 9890 12244 9942 12250
rect 9652 12198 9704 12210
rect 6659 12146 9652 12192
rect 6659 12140 9704 12146
rect 5643 12085 5649 12137
rect 5701 12085 5713 12137
rect 5765 12093 5771 12137
tri 5771 12093 5803 12125 sw
tri 6627 12093 6659 12125 se
rect 6659 12093 6711 12140
tri 6711 12106 6745 12140 nw
rect 5765 12091 5803 12093
tri 5803 12091 5805 12093 sw
tri 6625 12091 6627 12093 se
rect 6627 12091 6711 12093
rect 5765 12085 6711 12091
rect 5643 12039 6711 12085
rect 6770 12093 6779 12095
rect 6835 12093 6859 12095
rect 6770 12041 6776 12093
rect 6835 12041 6840 12093
rect 6770 12039 6779 12041
rect 6835 12039 6859 12041
rect 6915 12039 6924 12095
rect 9572 12081 9624 12087
tri 9566 12039 9572 12045 se
tri 9556 12029 9566 12039 se
rect 9566 12029 9572 12039
tri 9544 12017 9556 12029 se
rect 9556 12017 9624 12029
tri 9538 12011 9544 12017 se
rect 9544 12011 9572 12017
rect 6115 11959 6121 12011
rect 6173 11959 6187 12011
rect 6239 11965 9572 12011
rect 6239 11959 9624 11965
rect 6257 11869 9182 11921
rect 9234 11869 9246 11921
rect 9298 11869 9304 11921
rect 9890 11894 9942 11900
rect 5482 11785 5534 11837
tri 5448 11767 5466 11785 ne
rect 5466 11767 5534 11785
rect 5670 11767 5676 11819
rect 5728 11767 5740 11819
rect 5792 11767 5798 11819
rect 5871 11785 5877 11837
rect 5929 11785 5941 11837
rect 5993 11804 6081 11837
tri 6081 11804 6114 11837 sw
rect 5993 11788 6114 11804
tri 6114 11788 6130 11804 sw
rect 5993 11786 6130 11788
tri 6130 11786 6132 11788 sw
rect 7459 11786 7465 11838
rect 7517 11786 7529 11838
rect 7581 11834 8276 11838
rect 7581 11786 8154 11834
rect 5993 11785 6132 11786
tri 6132 11785 6133 11786 sw
tri 6059 11782 6062 11785 ne
rect 6062 11782 6133 11785
tri 6133 11782 6136 11785 sw
rect 7459 11782 8154 11786
rect 8206 11782 8218 11834
rect 8270 11782 8276 11834
tri 9864 11812 9890 11838 se
rect 9890 11812 9942 11842
tri 9856 11804 9864 11812 se
rect 9864 11804 9890 11812
tri 8999 11782 9005 11788 se
rect 9005 11782 9890 11804
tri 5466 11760 5473 11767 ne
rect 5473 11760 5534 11767
tri 5671 11760 5678 11767 ne
rect 5678 11760 5798 11767
tri 6062 11760 6084 11782 ne
rect 6084 11760 6136 11782
tri 6136 11760 6158 11782 sw
tri 8977 11760 8999 11782 se
rect 8999 11760 9890 11782
tri 5473 11754 5479 11760 ne
rect 5479 11754 5534 11760
tri 5678 11754 5684 11760 ne
rect 5684 11754 5798 11760
tri 6084 11754 6090 11760 ne
rect 6090 11754 6158 11760
tri 6158 11754 6164 11760 sw
tri 8971 11754 8977 11760 se
rect 8977 11754 9942 11760
tri 5479 11751 5482 11754 ne
rect 2661 11645 2667 11697
rect 2726 11645 2736 11697
rect 2993 11645 2994 11697
rect 3061 11645 3075 11697
rect 3131 11645 3145 11697
rect 3212 11645 3213 11697
rect 3469 11645 3478 11697
rect 3537 11645 3543 11697
rect 2661 11641 2670 11645
rect 2726 11641 2751 11645
rect 2807 11641 2832 11645
rect 2888 11641 2913 11645
rect 2969 11641 2994 11645
rect 3050 11641 3075 11645
rect 3131 11641 3156 11645
rect 3212 11641 3237 11645
rect 3293 11641 3318 11645
rect 3374 11641 3398 11645
rect 3454 11641 3478 11645
rect 3534 11641 3543 11645
rect 2661 11615 3543 11641
rect 2661 11611 2670 11615
rect 2726 11611 2751 11615
rect 2807 11611 2832 11615
rect 2888 11611 2913 11615
rect 2969 11611 2994 11615
rect 3050 11611 3075 11615
rect 3131 11611 3156 11615
rect 3212 11611 3237 11615
rect 3293 11611 3318 11615
rect 3374 11611 3398 11615
rect 3454 11611 3478 11615
rect 3534 11611 3543 11615
rect 2213 11601 2265 11607
tri 2265 11559 2271 11565 sw
rect 2661 11559 2667 11611
rect 2726 11559 2736 11611
rect 2993 11559 2994 11611
rect 3061 11559 3075 11611
rect 3131 11559 3145 11611
rect 3212 11559 3213 11611
rect 3469 11559 3478 11611
rect 3537 11559 3543 11611
rect 5482 11628 5534 11754
tri 5684 11751 5687 11754 ne
rect 5687 11751 5798 11754
tri 5687 11744 5694 11751 ne
rect 5694 11744 5798 11751
tri 6090 11744 6100 11754 ne
rect 6100 11744 9081 11754
tri 9081 11744 9091 11754 nw
rect 9970 11744 10022 11750
tri 5694 11733 5705 11744 ne
rect 5705 11697 5798 11744
tri 6100 11720 6124 11744 ne
rect 6124 11720 9057 11744
tri 9057 11720 9081 11744 nw
tri 6124 11711 6133 11720 ne
rect 6133 11711 9057 11720
tri 6133 11708 6136 11711 ne
rect 6136 11708 9057 11711
tri 5798 11697 5809 11708 sw
tri 6136 11702 6142 11708 ne
rect 6142 11702 9057 11708
tri 9964 11702 9970 11708 se
tri 9959 11697 9964 11702 se
rect 9964 11697 9970 11702
rect 5705 11692 5809 11697
tri 5809 11692 5814 11697 sw
tri 9954 11692 9959 11697 se
rect 9959 11692 9970 11697
rect 5705 11680 5814 11692
tri 5814 11680 5826 11692 sw
tri 9942 11680 9954 11692 se
rect 9954 11680 10022 11692
rect 5705 11674 5826 11680
tri 5826 11674 5832 11680 sw
tri 9936 11674 9942 11680 se
rect 9942 11674 9970 11680
tri 5534 11628 5536 11630 sw
rect 5705 11628 9970 11674
rect 5482 11622 5536 11628
tri 5536 11622 5542 11628 sw
rect 5705 11622 10022 11628
rect 5482 11608 5542 11622
tri 5482 11594 5496 11608 ne
rect 5496 11594 5542 11608
tri 5542 11594 5570 11622 sw
tri 5496 11588 5502 11594 ne
rect 5502 11588 9624 11594
tri 5502 11559 5531 11588 ne
rect 5531 11559 9572 11588
rect 2265 11549 2271 11559
rect 2213 11537 2271 11549
rect 2265 11536 2271 11537
tri 2271 11536 2294 11559 sw
tri 5531 11556 5534 11559 ne
rect 5534 11556 9572 11559
tri 5534 11542 5548 11556 ne
rect 5548 11542 9572 11556
tri 9538 11536 9544 11542 ne
rect 9544 11536 9572 11542
rect 2265 11531 2294 11536
tri 2294 11531 2299 11536 sw
tri 9544 11531 9549 11536 ne
rect 9549 11531 9624 11536
rect 2265 11524 4460 11531
tri 4460 11524 4467 11531 sw
tri 9549 11524 9556 11531 ne
rect 9556 11524 9624 11531
rect 2265 11485 4467 11524
rect 2213 11479 4467 11485
tri 4467 11479 4512 11524 sw
tri 9556 11508 9572 11524 ne
tri 4438 11477 4440 11479 ne
rect 4440 11477 4512 11479
tri 4512 11477 4514 11479 sw
tri 4440 11472 4445 11477 ne
rect 4445 11472 4514 11477
tri 4514 11472 4519 11477 sw
tri 4445 11457 4460 11472 ne
rect 4460 11457 4519 11472
tri 4460 11439 4478 11457 ne
rect 4478 11439 4519 11457
tri 4519 11439 4552 11472 sw
rect 9572 11466 9624 11472
rect 2133 11433 2402 11439
rect 2185 11381 2350 11433
tri 4478 11403 4514 11439 ne
rect 4514 11403 4552 11439
tri 4552 11403 4588 11439 sw
tri 4514 11397 4520 11403 ne
rect 4520 11397 4588 11403
rect 2133 11369 2402 11381
rect 2185 11317 2350 11369
tri 2402 11363 2436 11397 sw
tri 4520 11363 4554 11397 ne
rect 4554 11363 4588 11397
rect 2402 11355 4009 11363
tri 4009 11355 4017 11363 sw
tri 4554 11355 4562 11363 ne
rect 4562 11355 4588 11363
rect 2402 11329 4017 11355
tri 4017 11329 4043 11355 sw
tri 4562 11329 4588 11355 ne
tri 4588 11329 4662 11403 sw
rect 2402 11317 4043 11329
rect 2133 11311 4043 11317
tri 4043 11311 4061 11329 sw
tri 4588 11311 4606 11329 ne
rect 4606 11311 4662 11329
tri 4662 11311 4680 11329 sw
tri 3987 11283 4015 11311 ne
rect 4015 11283 4061 11311
rect 2707 11281 3868 11283
tri 3868 11281 3870 11283 sw
tri 4015 11281 4017 11283 ne
rect 4017 11281 4061 11283
tri 4061 11281 4091 11311 sw
tri 4606 11281 4636 11311 ne
rect 4636 11283 4680 11311
tri 4680 11283 4708 11311 sw
rect 4636 11281 4708 11283
rect 2707 11277 3870 11281
rect 2759 11275 3870 11277
tri 3870 11275 3876 11281 sw
tri 4017 11275 4023 11281 ne
rect 4023 11275 4091 11281
rect 2759 11238 3876 11275
tri 3876 11238 3913 11275 sw
tri 4023 11238 4060 11275 ne
rect 4060 11255 4091 11275
tri 4091 11255 4117 11281 sw
tri 4636 11255 4662 11281 ne
rect 4662 11255 4708 11281
tri 4708 11255 4736 11283 sw
rect 6714 11274 6770 11283
rect 4060 11238 4117 11255
tri 4117 11238 4134 11255 sw
tri 4662 11238 4679 11255 ne
rect 4679 11238 4736 11255
rect 2759 11231 3913 11238
tri 3913 11231 3920 11238 sw
tri 4060 11231 4067 11238 ne
rect 4067 11231 4134 11238
tri 4134 11231 4141 11238 sw
tri 4679 11231 4686 11238 ne
rect 4686 11231 4736 11238
rect 2707 11185 2759 11225
tri 2759 11197 2793 11231 nw
tri 3115 11197 3149 11231 ne
rect 623 11075 632 11131
rect 688 11075 713 11131
rect 769 11075 794 11131
rect 850 11075 875 11131
rect 931 11075 956 11131
rect 1012 11075 1037 11131
rect 1093 11075 1118 11131
rect 1174 11075 1198 11131
rect 1254 11075 1278 11131
rect 1334 11075 1358 11131
rect 1414 11079 1808 11131
rect 1860 11079 1872 11131
rect 1924 11079 1993 11131
rect 2707 11127 2759 11133
rect 3149 11127 3277 11231
tri 3277 11197 3311 11231 nw
tri 3846 11201 3876 11231 ne
rect 3876 11207 3920 11231
tri 3920 11207 3944 11231 sw
tri 4067 11207 4091 11231 ne
rect 4091 11207 4141 11231
tri 4141 11207 4165 11231 sw
tri 4686 11207 4710 11231 ne
rect 4710 11218 4736 11231
tri 4736 11218 4773 11255 sw
rect 4710 11207 4773 11218
rect 3876 11201 3944 11207
tri 3944 11201 3950 11207 sw
tri 4091 11201 4097 11207 ne
rect 4097 11201 4464 11207
tri 3876 11197 3880 11201 ne
rect 3880 11197 3950 11201
tri 3950 11197 3954 11201 sw
tri 4097 11197 4101 11201 ne
rect 4101 11197 4464 11201
tri 3880 11184 3893 11197 ne
rect 3893 11184 3954 11197
tri 3954 11184 3967 11197 sw
tri 4101 11184 4114 11197 ne
rect 4114 11184 4464 11197
tri 4710 11184 4733 11207 ne
rect 4733 11184 4773 11207
tri 4773 11184 4807 11218 sw
tri 6680 11184 6714 11218 se
rect 6714 11194 6770 11218
tri 3893 11181 3896 11184 ne
rect 3896 11181 3967 11184
tri 3967 11181 3970 11184 sw
tri 4114 11181 4117 11184 ne
rect 4117 11181 4464 11184
tri 4733 11181 4736 11184 ne
rect 4736 11181 4807 11184
tri 4807 11181 4810 11184 sw
tri 3896 11129 3948 11181 ne
rect 3948 11155 3970 11181
tri 3970 11155 3996 11181 sw
tri 4117 11155 4143 11181 ne
rect 4143 11155 4464 11181
rect 3948 11129 3996 11155
tri 3996 11129 4022 11155 sw
tri 4352 11129 4378 11155 ne
rect 4378 11129 4464 11155
tri 4736 11129 4788 11181 ne
rect 4788 11129 5012 11181
rect 5064 11129 5076 11181
rect 5128 11129 5134 11181
rect 5990 11132 5996 11184
rect 6048 11132 6070 11184
rect 6122 11132 6143 11184
rect 6195 11138 6714 11184
rect 6195 11132 6770 11138
rect 5990 11129 6770 11132
rect 6840 11189 6896 11198
tri 6839 11129 6840 11130 se
rect 6840 11129 6896 11133
tri 3948 11127 3950 11129 ne
rect 3950 11127 4022 11129
tri 4022 11127 4024 11129 sw
tri 4378 11127 4380 11129 ne
rect 4380 11127 4464 11129
rect 1414 11075 1993 11079
rect 2627 11117 2679 11123
tri 2679 11075 2685 11081 sw
rect 3149 11075 3155 11127
rect 3207 11075 3219 11127
rect 3271 11075 3277 11127
tri 3598 11075 3604 11081 se
rect 3604 11075 3610 11127
rect 3662 11075 3674 11127
rect 3726 11075 3732 11127
tri 3950 11121 3956 11127 ne
rect 3956 11121 4069 11127
tri 3956 11115 3962 11121 ne
rect 3962 11115 4069 11121
tri 3962 11081 3996 11115 ne
rect 3996 11081 4069 11115
tri 3996 11075 4002 11081 ne
rect 4002 11075 4069 11081
rect 4121 11075 4133 11127
rect 4185 11075 4191 11127
tri 4380 11121 4386 11127 ne
rect 2679 11065 2685 11075
rect 2627 11053 2685 11065
rect 1733 11037 1785 11043
rect 2679 11047 2685 11053
tri 2685 11047 2713 11075 sw
tri 3570 11047 3598 11075 se
rect 3598 11047 3662 11075
tri 3662 11047 3690 11075 nw
rect 2679 11001 3087 11047
rect 1733 10973 1785 10985
tri 1785 10967 1819 11001 sw
rect 2627 10995 3087 11001
rect 3139 10995 3151 11047
rect 3203 11044 3659 11047
tri 3659 11044 3662 11047 nw
rect 3203 10995 3656 11044
tri 3656 11041 3659 11044 nw
tri 4380 10995 4386 11001 se
rect 4386 10995 4464 11127
tri 6806 11096 6839 11129 se
rect 6839 11109 6896 11129
rect 6839 11096 6840 11109
rect 5715 11044 5721 11096
rect 5773 11044 5842 11096
rect 5894 11044 5963 11096
rect 6015 11044 6083 11096
rect 6135 11044 6203 11096
rect 6255 11053 6840 11096
rect 6255 11044 6896 11053
rect 7069 11057 7121 11063
tri 4379 10994 4380 10995 se
rect 4380 10994 4464 10995
tri 4378 10993 4379 10994 se
rect 4379 10993 4464 10994
tri 4352 10967 4378 10993 se
rect 4378 10967 4464 10993
rect 1785 10921 3411 10967
rect 1733 10915 3411 10921
rect 3463 10915 3480 10967
rect 3532 10915 3707 10967
rect 3759 10915 3772 10967
rect 3824 10915 3830 10967
rect 4027 10915 4033 10967
rect 4085 10915 4097 10967
rect 4149 10915 4342 10967
rect 4394 10915 4406 10967
rect 4458 10915 4464 10967
rect 7069 11000 7121 11005
tri 7121 11000 7155 11034 sw
rect 7069 10994 8517 11000
rect 7069 10993 8465 10994
rect 7121 10948 8465 10993
rect 7121 10942 7128 10948
tri 7128 10942 7134 10948 nw
tri 8431 10942 8437 10948 ne
rect 8437 10942 8465 10948
rect 7069 10935 7121 10941
tri 7121 10935 7128 10942 nw
tri 8437 10935 8444 10942 ne
rect 8444 10935 8517 10942
tri 8444 10930 8449 10935 ne
rect 8449 10930 8517 10935
tri 8449 10915 8464 10930 ne
rect 8464 10915 8465 10930
tri 8464 10914 8465 10915 ne
rect 8465 10872 8517 10878
rect 623 10841 6864 10842
rect 623 10785 632 10841
rect 688 10785 713 10841
rect 769 10785 794 10841
rect 850 10785 875 10841
rect 931 10785 956 10841
rect 1012 10785 1037 10841
rect 1093 10785 1118 10841
rect 1174 10785 1198 10841
rect 1254 10785 1278 10841
rect 1334 10785 1358 10841
rect 1414 10789 3121 10841
rect 3173 10789 3186 10841
rect 3238 10789 3251 10841
rect 3303 10789 3316 10841
rect 3368 10789 3381 10841
rect 3433 10789 3446 10841
rect 3498 10789 3511 10841
rect 3563 10789 3576 10841
rect 3628 10789 3641 10841
rect 3693 10789 3706 10841
rect 3758 10789 3771 10841
rect 3823 10789 3836 10841
rect 3888 10789 3901 10841
rect 3953 10789 3966 10841
rect 4018 10789 4031 10841
rect 4083 10789 4096 10841
rect 4148 10789 4160 10841
rect 4212 10789 4224 10841
rect 4276 10789 4288 10841
rect 4340 10789 4352 10841
rect 4404 10789 4416 10841
rect 4468 10789 4480 10841
rect 4532 10789 4544 10841
rect 4596 10789 4608 10841
rect 4660 10789 4672 10841
rect 4724 10789 4736 10841
rect 4788 10789 4800 10841
rect 4852 10789 4864 10841
rect 4916 10789 4928 10841
rect 4980 10789 4992 10841
rect 5044 10789 5056 10841
rect 5108 10789 5120 10841
rect 5172 10789 5184 10841
rect 5236 10789 5248 10841
rect 5300 10789 5312 10841
rect 5364 10789 5376 10841
rect 5428 10789 5440 10841
rect 5492 10789 5504 10841
rect 5556 10789 5568 10841
rect 5620 10789 5632 10841
rect 5684 10789 5696 10841
rect 5748 10789 5760 10841
rect 5812 10789 5824 10841
rect 5876 10789 5888 10841
rect 5940 10789 5952 10841
rect 6004 10789 6016 10841
rect 6068 10789 6080 10841
rect 6132 10789 6144 10841
rect 6196 10789 6208 10841
rect 6260 10835 6864 10841
rect 6260 10789 6711 10835
rect 1414 10785 6711 10789
rect 623 10783 6711 10785
rect 6763 10783 6811 10835
rect 6863 10783 6864 10835
rect 623 10771 6864 10783
rect 623 10719 3121 10771
rect 3173 10719 3186 10771
rect 3238 10719 3251 10771
rect 3303 10719 3316 10771
rect 3368 10719 3381 10771
rect 3433 10719 3446 10771
rect 3498 10719 3511 10771
rect 3563 10719 3576 10771
rect 3628 10719 3641 10771
rect 3693 10719 3706 10771
rect 3758 10719 3771 10771
rect 3823 10719 3836 10771
rect 3888 10719 3901 10771
rect 3953 10719 3966 10771
rect 4018 10719 4031 10771
rect 4083 10719 4096 10771
rect 4148 10719 4160 10771
rect 4212 10719 4224 10771
rect 4276 10719 4288 10771
rect 4340 10719 4352 10771
rect 4404 10719 4416 10771
rect 4468 10719 4480 10771
rect 4532 10719 4544 10771
rect 4596 10719 4608 10771
rect 4660 10719 4672 10771
rect 4724 10719 4736 10771
rect 4788 10719 4800 10771
rect 4852 10719 4864 10771
rect 4916 10719 4928 10771
rect 4980 10719 4992 10771
rect 5044 10719 5056 10771
rect 5108 10719 5120 10771
rect 5172 10719 5184 10771
rect 5236 10719 5248 10771
rect 5300 10719 5312 10771
rect 5364 10719 5376 10771
rect 5428 10719 5440 10771
rect 5492 10719 5504 10771
rect 5556 10719 5568 10771
rect 5620 10719 5632 10771
rect 5684 10719 5696 10771
rect 5748 10719 5760 10771
rect 5812 10719 5824 10771
rect 5876 10719 5888 10771
rect 5940 10719 5952 10771
rect 6004 10719 6016 10771
rect 6068 10719 6080 10771
rect 6132 10719 6144 10771
rect 6196 10719 6208 10771
rect 6260 10719 6711 10771
rect 6763 10719 6811 10771
rect 6863 10719 6864 10771
rect 623 10707 6864 10719
rect 623 10705 6711 10707
rect 623 10649 632 10705
rect 688 10649 713 10705
rect 769 10649 794 10705
rect 850 10649 875 10705
rect 931 10649 956 10705
rect 1012 10649 1037 10705
rect 1093 10649 1118 10705
rect 1174 10649 1198 10705
rect 1254 10649 1278 10705
rect 1334 10649 1358 10705
rect 1414 10701 6711 10705
rect 1414 10649 3121 10701
rect 3173 10649 3186 10701
rect 3238 10649 3251 10701
rect 3303 10649 3316 10701
rect 3368 10649 3381 10701
rect 3433 10649 3446 10701
rect 3498 10649 3511 10701
rect 3563 10649 3576 10701
rect 3628 10649 3641 10701
rect 3693 10649 3706 10701
rect 3758 10649 3771 10701
rect 3823 10649 3836 10701
rect 3888 10649 3901 10701
rect 3953 10649 3966 10701
rect 4018 10649 4031 10701
rect 4083 10649 4096 10701
rect 4148 10649 4160 10701
rect 4212 10649 4224 10701
rect 4276 10649 4288 10701
rect 4340 10649 4352 10701
rect 4404 10649 4416 10701
rect 4468 10649 4480 10701
rect 4532 10649 4544 10701
rect 4596 10649 4608 10701
rect 4660 10649 4672 10701
rect 4724 10649 4736 10701
rect 4788 10649 4800 10701
rect 4852 10649 4864 10701
rect 4916 10649 4928 10701
rect 4980 10649 4992 10701
rect 5044 10649 5056 10701
rect 5108 10649 5120 10701
rect 5172 10649 5184 10701
rect 5236 10649 5248 10701
rect 5300 10649 5312 10701
rect 5364 10649 5376 10701
rect 5428 10649 5440 10701
rect 5492 10649 5504 10701
rect 5556 10649 5568 10701
rect 5620 10649 5632 10701
rect 5684 10649 5696 10701
rect 5748 10649 5760 10701
rect 5812 10649 5824 10701
rect 5876 10649 5888 10701
rect 5940 10649 5952 10701
rect 6004 10649 6016 10701
rect 6068 10649 6080 10701
rect 6132 10649 6144 10701
rect 6196 10649 6208 10701
rect 6260 10655 6711 10701
rect 6763 10655 6811 10707
rect 6863 10655 6864 10707
rect 6260 10649 6864 10655
rect 8758 10635 8767 10639
rect 8823 10635 8847 10639
rect 8544 10579 8553 10635
rect 8609 10633 8633 10635
rect 8689 10633 8698 10635
rect 8628 10581 8633 10633
rect 8692 10581 8698 10633
rect 8758 10583 8764 10635
rect 8823 10583 8846 10635
rect 8903 10583 8912 10639
rect 8609 10579 8633 10581
rect 8689 10579 8698 10581
tri 10251 10567 10261 10577 se
rect 10261 10568 10317 10577
rect 2213 10557 2265 10563
tri 2265 10515 2271 10521 sw
rect 2314 10515 2320 10567
rect 2372 10515 2384 10567
rect 2436 10515 3595 10567
tri 10247 10563 10251 10567 se
rect 10251 10563 10261 10567
tri 10235 10551 10247 10563 se
rect 10247 10551 10261 10563
rect 7120 10545 10261 10551
rect 6314 10521 6864 10527
rect 2265 10505 2271 10515
rect 2213 10493 2271 10505
rect 2265 10487 2271 10493
tri 2271 10487 2299 10515 sw
rect 2265 10453 3493 10487
rect 2265 10441 2373 10453
rect 2213 10435 2373 10441
tri 2339 10401 2373 10435 ne
rect 2425 10435 3493 10453
rect 6366 10469 6390 10521
rect 6442 10469 6466 10521
rect 6518 10469 6744 10521
rect 6796 10469 6812 10521
rect 6314 10449 6864 10469
tri 2425 10401 2459 10435 nw
tri 3454 10401 3488 10435 ne
rect 2373 10389 2425 10401
rect 1813 10352 2286 10358
rect 1865 10325 2286 10352
tri 2286 10325 2298 10337 sw
rect 2373 10331 2425 10337
rect 6366 10397 6390 10449
rect 6442 10397 6466 10449
rect 6518 10397 6744 10449
rect 6796 10397 6812 10449
rect 7120 10493 7128 10545
rect 7180 10512 10261 10545
rect 7180 10493 10317 10512
rect 7120 10488 10317 10493
rect 7120 10481 10261 10488
rect 7120 10429 7128 10481
rect 7180 10432 10261 10481
rect 7180 10429 10317 10432
rect 7120 10423 10317 10429
rect 6314 10377 6864 10397
rect 6366 10325 6390 10377
rect 6442 10325 6466 10377
rect 6518 10325 6744 10377
rect 6796 10325 6812 10377
rect 1865 10315 2298 10325
tri 2298 10315 2308 10325 sw
rect 1865 10306 2308 10315
tri 2308 10306 2317 10315 sw
rect 1865 10305 1898 10306
tri 1898 10305 1899 10306 nw
tri 2200 10305 2201 10306 ne
rect 2201 10305 2317 10306
tri 2317 10305 2318 10306 sw
rect 6314 10305 6864 10325
rect 8374 10360 9011 10391
rect 1865 10303 1896 10305
tri 1896 10303 1898 10305 nw
tri 2201 10303 2203 10305 ne
rect 2203 10303 2318 10305
tri 2318 10303 2320 10305 sw
rect 1813 10288 1865 10300
tri 1865 10272 1896 10303 nw
tri 2203 10272 2234 10303 ne
rect 1813 10230 1865 10236
rect 2133 10247 2185 10253
rect 2234 10251 3735 10303
rect 3787 10251 3799 10303
rect 3851 10251 3857 10303
rect 6366 10253 6390 10305
rect 6442 10253 6466 10305
rect 6518 10253 6744 10305
rect 6796 10253 6812 10305
rect 7323 10315 7375 10321
tri 7307 10263 7323 10279 se
rect 8374 10304 8383 10360
rect 8439 10304 8463 10360
rect 8519 10339 9011 10360
rect 9063 10339 9087 10391
rect 9139 10339 9145 10391
rect 8519 10325 9145 10339
rect 8519 10304 9011 10325
tri 7375 10273 7381 10279 sw
rect 8374 10273 9011 10304
rect 9063 10273 9087 10325
rect 9139 10273 9145 10325
rect 7375 10263 7381 10273
rect 6314 10233 6864 10253
tri 7295 10251 7307 10263 se
rect 7307 10251 7381 10263
tri 7289 10245 7295 10251 se
rect 7295 10245 7323 10251
rect 2133 10183 2185 10195
tri 2185 10181 2215 10211 sw
rect 6366 10181 6390 10233
rect 6442 10181 6466 10233
rect 6518 10181 6744 10233
rect 6796 10181 6812 10233
rect 2185 10177 2215 10181
tri 2215 10177 2219 10181 sw
rect 2185 10131 3261 10177
rect 2133 10125 3261 10131
rect 3313 10125 3327 10177
rect 3379 10125 3385 10177
rect 6314 10161 6864 10181
rect 6366 10109 6390 10161
rect 6442 10109 6466 10161
rect 6518 10109 6744 10161
rect 6796 10109 6812 10161
rect 7222 10239 7323 10245
rect 7274 10199 7323 10239
rect 7375 10245 7381 10251
tri 7381 10245 7409 10273 sw
rect 7375 10199 8862 10245
rect 7274 10193 8862 10199
rect 8914 10193 8926 10245
rect 8978 10193 8984 10245
rect 7274 10187 7280 10193
rect 7222 10175 7280 10187
rect 7274 10165 7280 10175
tri 7280 10165 7308 10193 nw
tri 7274 10159 7280 10165 nw
rect 7715 10159 8977 10165
rect 7222 10117 7274 10123
rect 6314 10103 6864 10109
rect 7767 10107 7791 10159
rect 7843 10156 8977 10159
rect 7843 10107 8916 10156
rect 7715 10100 8916 10107
rect 8972 10100 8977 10156
rect 1977 10035 1983 10087
rect 2035 10035 2047 10087
rect 2099 10035 3244 10087
rect 7715 10076 8977 10100
rect 7715 10069 8916 10076
rect 7767 10017 7791 10069
rect 7843 10020 8916 10069
rect 8972 10020 8977 10076
rect 7843 10017 8977 10020
rect 7715 10011 8977 10017
rect 2213 10001 3511 10007
rect 2265 9955 3511 10001
rect 3563 9955 3575 10007
rect 3627 9955 3633 10007
rect 2265 9949 2277 9955
rect 2213 9937 2277 9949
rect 2265 9933 2277 9937
tri 2277 9933 2299 9955 nw
rect 3702 9933 3708 9985
rect 3760 9933 3772 9985
rect 3824 9933 3830 9985
rect 3966 9951 4018 10003
rect 8011 9956 9064 9962
rect 3966 9933 4034 9951
tri 4034 9933 4052 9951 nw
tri 2265 9921 2277 9933 nw
tri 3709 9921 3721 9933 ne
rect 3721 9921 3816 9933
tri 3721 9920 3722 9921 ne
rect 3722 9920 3816 9921
tri 3816 9920 3829 9933 nw
rect 3966 9920 4021 9933
tri 4021 9920 4034 9933 nw
tri 3722 9909 3733 9920 ne
rect 3733 9909 3805 9920
tri 3805 9909 3816 9920 nw
tri 3733 9904 3738 9909 ne
rect 3738 9904 3800 9909
tri 3800 9904 3805 9909 nw
tri 3738 9899 3743 9904 ne
rect 2213 9879 2265 9885
rect 623 9813 3099 9851
rect 623 9757 632 9813
rect 688 9757 713 9813
rect 769 9757 794 9813
rect 850 9757 875 9813
rect 931 9757 956 9813
rect 1012 9757 1037 9813
rect 1093 9757 1118 9813
rect 1174 9757 1198 9813
rect 1254 9757 1278 9813
rect 1334 9757 1358 9813
rect 1414 9799 3099 9813
rect 3151 9799 3166 9851
rect 3218 9799 3233 9851
rect 3285 9799 3300 9851
rect 3352 9799 3367 9851
rect 3419 9799 3434 9851
rect 3486 9799 3500 9851
rect 3552 9799 3566 9851
rect 3618 9799 3632 9851
rect 3684 9799 3690 9851
rect 1414 9771 3690 9799
rect 1414 9757 3099 9771
rect 623 9719 3099 9757
rect 3151 9719 3166 9771
rect 3218 9719 3233 9771
rect 3285 9719 3300 9771
rect 3352 9719 3367 9771
rect 3419 9719 3434 9771
rect 3486 9719 3500 9771
rect 3552 9719 3566 9771
rect 3618 9719 3632 9771
rect 3684 9719 3690 9771
rect 1893 9677 3318 9683
rect 1945 9661 3318 9677
tri 3741 9666 3743 9668 se
rect 3743 9666 3795 9904
tri 3795 9899 3800 9904 nw
tri 3318 9661 3323 9666 sw
tri 3736 9661 3741 9666 se
rect 3741 9661 3795 9666
rect 1945 9643 3323 9661
tri 3323 9643 3341 9661 sw
tri 3718 9643 3736 9661 se
rect 3736 9646 3795 9661
rect 3736 9643 3792 9646
tri 3792 9643 3795 9646 nw
rect 1945 9632 3341 9643
tri 3341 9632 3352 9643 sw
tri 3707 9632 3718 9643 se
rect 3718 9632 3781 9643
tri 3781 9632 3792 9643 nw
rect 1945 9625 1956 9632
rect 1893 9613 1956 9625
rect 1945 9609 1956 9613
tri 1956 9609 1979 9632 nw
tri 3232 9609 3255 9632 ne
rect 3255 9609 3758 9632
tri 3758 9609 3781 9632 nw
tri 1945 9598 1956 9609 nw
tri 3255 9598 3266 9609 ne
rect 3266 9598 3747 9609
tri 3747 9598 3758 9609 nw
rect 3266 9594 3743 9598
tri 3743 9594 3747 9598 nw
rect 3266 9591 3740 9594
tri 3740 9591 3743 9594 nw
rect 3266 9580 3729 9591
tri 3729 9580 3740 9591 nw
tri 3958 9580 3966 9588 se
rect 3966 9580 4018 9920
tri 4018 9917 4021 9920 nw
tri 8008 9917 8011 9920 se
rect 8011 9917 9012 9956
tri 8000 9909 8008 9917 se
rect 8008 9909 9012 9917
tri 7995 9904 8000 9909 se
rect 8000 9904 8092 9909
tri 8092 9904 8097 9909 nw
tri 8978 9904 8983 9909 ne
rect 8983 9904 9012 9909
tri 7983 9892 7995 9904 se
rect 7995 9892 8080 9904
tri 8080 9892 8092 9904 nw
tri 8983 9892 8995 9904 ne
rect 8995 9892 9064 9904
tri 7977 9886 7983 9892 se
rect 7983 9886 8074 9892
tri 8074 9886 8080 9892 nw
tri 8995 9886 9001 9892 ne
rect 9001 9886 9012 9892
tri 5698 9875 5709 9886 se
rect 5709 9875 8063 9886
tri 8063 9875 8074 9886 nw
tri 9001 9875 9012 9886 ne
tri 5663 9840 5698 9875 se
rect 5698 9840 8063 9875
tri 5647 9824 5663 9840 se
rect 5663 9834 8063 9840
rect 9492 9876 9544 9882
rect 9012 9834 9064 9840
tri 9486 9834 9492 9840 se
rect 5663 9824 5721 9834
tri 5721 9824 5731 9834 nw
tri 9476 9824 9486 9834 se
rect 9486 9824 9492 9834
tri 5643 9820 5647 9824 se
rect 5647 9820 5717 9824
tri 5717 9820 5721 9824 nw
tri 9472 9820 9476 9824 se
rect 9476 9820 9544 9824
rect 5643 9812 5709 9820
tri 5709 9812 5717 9820 nw
tri 9464 9812 9472 9820 se
rect 9472 9812 9544 9820
rect 5643 9806 5703 9812
tri 5703 9806 5709 9812 nw
tri 9458 9806 9464 9812 se
rect 9464 9806 9492 9812
tri 5634 9668 5643 9677 se
rect 5643 9668 5695 9806
tri 5695 9798 5703 9806 nw
rect 5866 9760 9492 9806
rect 5866 9754 9544 9760
rect 5866 9726 5965 9754
tri 5965 9726 5993 9754 nw
tri 5845 9674 5866 9695 se
rect 5866 9674 5959 9726
tri 5959 9720 5965 9726 nw
tri 6297 9720 6303 9726 se
rect 6303 9720 6623 9726
tri 6251 9674 6297 9720 se
rect 6297 9674 6571 9720
tri 5839 9668 5845 9674 se
rect 5845 9668 5959 9674
tri 6245 9668 6251 9674 se
rect 6251 9668 6319 9674
tri 6319 9668 6325 9674 nw
tri 6537 9668 6543 9674 ne
rect 6543 9668 6571 9674
tri 5627 9661 5634 9668 se
rect 5634 9661 5695 9668
tri 5832 9661 5839 9668 se
rect 5839 9661 5959 9668
tri 5609 9643 5627 9661 se
rect 5627 9643 5695 9661
rect 5643 9591 5695 9643
rect 5831 9609 5837 9661
rect 5889 9609 5901 9661
rect 5953 9609 5959 9661
tri 6237 9660 6245 9668 se
rect 6245 9660 6311 9668
tri 6311 9660 6319 9668 nw
tri 6543 9660 6551 9668 ne
rect 6551 9660 6623 9668
tri 6233 9656 6237 9660 se
rect 6237 9656 6307 9660
tri 6307 9656 6311 9660 nw
tri 6551 9656 6555 9660 ne
rect 6555 9656 6623 9660
tri 6229 9652 6233 9656 se
rect 6233 9652 6303 9656
tri 6303 9652 6307 9656 nw
tri 6555 9652 6559 9656 ne
rect 6559 9652 6571 9656
tri 6220 9643 6229 9652 se
rect 6229 9643 6294 9652
tri 6294 9643 6303 9652 nw
tri 6559 9643 6568 9652 ne
rect 6568 9643 6571 9652
rect 6028 9591 6034 9643
rect 6086 9591 6098 9643
rect 6150 9640 6291 9643
tri 6291 9640 6294 9643 nw
tri 6568 9640 6571 9643 ne
rect 6150 9608 6259 9640
tri 6259 9608 6291 9640 nw
rect 6150 9604 6255 9608
tri 6255 9604 6259 9608 nw
rect 7222 9608 7228 9660
rect 7280 9608 7292 9660
rect 7344 9608 7943 9660
rect 7222 9604 7943 9608
rect 7999 9604 8023 9660
rect 8079 9604 8089 9660
rect 9092 9632 9144 9638
rect 6150 9591 6242 9604
tri 6242 9591 6255 9604 nw
rect 6571 9598 6623 9604
tri 9090 9591 9092 9593 se
tri 9079 9580 9090 9591 se
rect 9090 9580 9092 9591
tri 3946 9568 3958 9580 se
rect 3958 9568 4018 9580
tri 9067 9568 9079 9580 se
rect 9079 9568 9144 9580
rect 1893 9555 1945 9561
tri 3937 9559 3946 9568 se
rect 3946 9566 4018 9568
rect 3946 9559 4011 9566
tri 4011 9559 4018 9566 nw
tri 9058 9559 9067 9568 se
rect 9067 9559 9092 9568
tri 3933 9555 3937 9559 se
rect 3937 9555 4004 9559
tri 3930 9552 3933 9555 se
rect 3933 9552 4004 9555
tri 4004 9552 4011 9559 nw
rect 1973 9546 3968 9552
rect 2025 9516 3968 9546
tri 3968 9516 4004 9552 nw
rect 6418 9516 9092 9559
rect 2025 9500 3952 9516
tri 3952 9500 3968 9516 nw
rect 6418 9507 9144 9516
rect 2025 9494 2028 9500
rect 1973 9482 2028 9494
rect 2025 9469 2028 9482
tri 2028 9469 2059 9500 nw
tri 2025 9466 2028 9469 nw
rect 1973 9424 2025 9430
rect 6276 9417 6282 9469
rect 6334 9417 6348 9469
rect 6400 9417 8298 9469
rect 8350 9417 8362 9469
rect 8414 9417 8420 9469
rect 9172 9358 9224 9364
rect 5804 9291 5810 9343
rect 5862 9291 5874 9343
rect 5926 9306 8925 9343
tri 8925 9306 8941 9322 sw
tri 9156 9306 9172 9322 se
rect 5926 9294 8941 9306
tri 8941 9294 8953 9306 sw
tri 9144 9294 9156 9306 se
rect 9156 9294 9224 9306
rect 5926 9291 8953 9294
tri 8839 9288 8842 9291 ne
rect 8842 9288 8953 9291
tri 8953 9288 8959 9294 sw
tri 9138 9288 9144 9294 se
rect 9144 9288 9172 9294
tri 8842 9262 8868 9288 ne
rect 8868 9262 9172 9288
rect 7034 9210 7040 9262
rect 7092 9210 7112 9262
rect 7164 9210 7721 9262
rect 7773 9210 7785 9262
rect 7837 9210 7843 9262
tri 8868 9257 8873 9262 ne
rect 8873 9242 9172 9262
rect 8873 9236 9224 9242
tri 8394 9210 8403 9219 se
rect 8403 9210 8702 9219
tri 8377 9193 8394 9210 se
rect 8394 9193 8702 9210
tri 6173 9167 6199 9193 sw
tri 8351 9167 8377 9193 se
rect 8377 9167 8702 9193
rect 8754 9167 8766 9219
rect 8818 9167 8824 9219
rect 6173 9159 6199 9167
tri 6199 9159 6207 9167 sw
tri 8343 9159 8351 9167 se
rect 8351 9159 8407 9167
rect 6169 9149 8407 9159
tri 8407 9149 8425 9167 nw
rect 8852 9149 8904 9155
rect 6169 9107 8365 9149
tri 8365 9107 8407 9149 nw
tri 8846 9107 8852 9113 se
tri 8836 9097 8846 9107 se
rect 8846 9097 8852 9107
tri 8824 9085 8836 9097 se
rect 8836 9085 8904 9097
tri 8818 9079 8824 9085 se
rect 8824 9079 8852 9085
rect 6067 9033 8852 9079
rect 6067 9027 8904 9033
rect 8208 8927 8260 8933
tri 8192 8875 8208 8891 se
tri 8180 8863 8192 8875 se
rect 8192 8863 8260 8875
tri 8174 8857 8180 8863 se
rect 8180 8857 8208 8863
rect 6067 8811 8208 8857
rect 6067 8805 8260 8811
rect 6169 8771 7955 8777
rect 6169 8725 7903 8771
rect 6173 8719 6201 8725
tri 6201 8719 6207 8725 nw
tri 7869 8719 7875 8725 ne
rect 7875 8719 7903 8725
rect 6173 8707 6189 8719
tri 6189 8707 6201 8719 nw
tri 7875 8707 7887 8719 ne
rect 7887 8707 7955 8719
tri 6173 8691 6189 8707 nw
tri 7887 8691 7903 8707 ne
rect 7903 8649 7955 8655
rect 8004 8642 8580 8648
tri 7973 8596 8004 8627 se
rect 8004 8596 8528 8642
tri 7970 8593 7973 8596 se
rect 7973 8593 8087 8596
tri 8087 8593 8090 8596 nw
tri 8494 8593 8497 8596 ne
rect 8497 8593 8528 8596
rect 5804 8541 5810 8593
rect 5862 8541 5874 8593
rect 5926 8590 8084 8593
tri 8084 8590 8087 8593 nw
tri 8497 8590 8500 8593 ne
rect 8500 8590 8528 8593
rect 5926 8578 8072 8590
tri 8072 8578 8084 8590 nw
tri 8500 8578 8512 8590 ne
rect 8512 8578 8580 8590
rect 5926 8541 8056 8578
tri 8056 8562 8072 8578 nw
tri 8512 8568 8522 8578 ne
rect 8522 8568 8528 8578
rect 8368 8562 8420 8568
tri 8522 8562 8528 8568 ne
rect 8528 8520 8580 8526
tri 8365 8498 8368 8501 se
rect 8368 8498 8420 8510
tri 8334 8467 8365 8498 se
rect 8365 8467 8368 8498
rect 6276 8415 6282 8467
rect 6334 8415 6348 8467
rect 6400 8446 8368 8467
rect 6400 8440 8420 8446
rect 6400 8415 8368 8440
tri 8368 8415 8393 8440 nw
tri 8447 8406 8448 8407 se
rect 8448 8406 8500 8412
tri 8418 8377 8447 8406 se
rect 8447 8377 8448 8406
rect 6418 8354 8448 8377
rect 6418 8342 8500 8354
rect 6418 8325 8448 8342
tri 8414 8294 8445 8325 ne
rect 8445 8294 8448 8325
rect 5643 8241 5695 8293
tri 5609 8223 5627 8241 ne
rect 5627 8223 5695 8241
rect 5831 8223 5837 8275
rect 5889 8223 5901 8275
rect 5953 8223 5959 8275
rect 6028 8241 6034 8293
rect 6086 8241 6098 8293
rect 6150 8242 6242 8293
tri 6242 8242 6293 8293 sw
rect 7072 8242 7078 8294
rect 7130 8242 7143 8294
rect 7195 8242 7833 8294
rect 7885 8242 7897 8294
rect 7949 8242 7955 8294
tri 8445 8291 8448 8294 ne
rect 8288 8280 8340 8286
rect 8448 8284 8500 8290
tri 8286 8242 8288 8244 se
rect 6150 8241 6293 8242
tri 6293 8241 6294 8242 sw
tri 8285 8241 8286 8242 se
rect 8286 8241 8288 8242
tri 6220 8228 6233 8241 ne
rect 6233 8228 6294 8241
tri 6294 8228 6307 8241 sw
tri 8272 8228 8285 8241 se
rect 8285 8228 8288 8241
tri 6233 8223 6238 8228 ne
rect 6238 8223 6307 8228
tri 6307 8223 6312 8228 sw
tri 8267 8223 8272 8228 se
rect 8272 8223 8340 8228
tri 5627 8221 5629 8223 ne
rect 5629 8221 5695 8223
tri 5832 8221 5834 8223 ne
rect 5834 8221 5959 8223
tri 6238 8221 6240 8223 ne
rect 6240 8221 6312 8223
tri 6312 8221 6314 8223 sw
tri 8265 8221 8267 8223 se
rect 8267 8221 8340 8223
tri 5629 8216 5634 8221 ne
rect 5634 8216 5695 8221
tri 5834 8216 5839 8221 ne
rect 5839 8216 5959 8221
tri 6240 8216 6245 8221 ne
rect 6245 8216 6314 8221
tri 6314 8216 6319 8221 sw
tri 8260 8216 8265 8221 se
rect 8265 8216 8340 8221
tri 5634 8207 5643 8216 ne
rect 628 8097 637 8153
rect 693 8097 718 8153
rect 774 8097 798 8153
rect 854 8097 878 8153
rect 934 8097 958 8153
rect 1014 8097 1038 8153
rect 1094 8097 1118 8153
rect 1174 8097 1198 8153
rect 1254 8097 1278 8153
rect 1334 8097 1358 8153
rect 1414 8152 5465 8153
rect 1414 8100 3148 8152
rect 3200 8100 3213 8152
rect 3265 8100 3278 8152
rect 3330 8100 3343 8152
rect 3395 8100 3408 8152
rect 3460 8100 3473 8152
rect 3525 8100 3538 8152
rect 3590 8100 3603 8152
rect 3655 8100 3668 8152
rect 3720 8100 3733 8152
rect 3785 8100 3798 8152
rect 3850 8100 3863 8152
rect 3915 8100 3928 8152
rect 3980 8100 3993 8152
rect 4045 8100 4058 8152
rect 4110 8100 4123 8152
rect 4175 8100 4188 8152
rect 4240 8100 4253 8152
rect 4305 8100 4318 8152
rect 4370 8100 4383 8152
rect 1414 8097 4383 8100
rect 628 8088 4383 8097
rect 628 8036 3148 8088
rect 3200 8036 3213 8088
rect 3265 8036 3278 8088
rect 3330 8036 3343 8088
rect 3395 8036 3408 8088
rect 3460 8036 3473 8088
rect 3525 8036 3538 8088
rect 3590 8036 3603 8088
rect 3655 8036 3668 8088
rect 3720 8036 3733 8088
rect 3785 8036 3798 8088
rect 3850 8036 3863 8088
rect 3915 8036 3928 8088
rect 3980 8036 3993 8088
rect 4045 8036 4058 8088
rect 4110 8036 4123 8088
rect 4175 8036 4188 8088
rect 4240 8036 4253 8088
rect 4305 8036 4318 8088
rect 4370 8036 4383 8088
rect 628 8027 4383 8036
rect 628 7971 637 8027
rect 693 7971 718 8027
rect 774 7971 798 8027
rect 854 7971 878 8027
rect 934 7971 958 8027
rect 1014 7971 1038 8027
rect 1094 7971 1118 8027
rect 1174 7971 1198 8027
rect 1254 7971 1278 8027
rect 1334 7971 1358 8027
rect 1414 8024 4383 8027
rect 1414 7972 3148 8024
rect 3200 7972 3213 8024
rect 3265 7972 3278 8024
rect 3330 7972 3343 8024
rect 3395 7972 3408 8024
rect 3460 7972 3473 8024
rect 3525 7972 3538 8024
rect 3590 7972 3603 8024
rect 3655 7972 3668 8024
rect 3720 7972 3733 8024
rect 3785 7972 3798 8024
rect 3850 7972 3863 8024
rect 3915 7972 3928 8024
rect 3980 7972 3993 8024
rect 4045 7972 4058 8024
rect 4110 7972 4123 8024
rect 4175 7972 4188 8024
rect 4240 7972 4253 8024
rect 4305 7972 4318 8024
rect 4370 7972 4383 8024
rect 5459 7972 5465 8152
rect 5643 8078 5695 8216
tri 5839 8207 5848 8216 ne
rect 5848 8207 5959 8216
tri 6245 8210 6251 8216 ne
rect 6251 8210 6319 8216
tri 6319 8210 6325 8216 sw
tri 8254 8210 8260 8216 se
rect 8260 8210 8288 8216
tri 5848 8189 5866 8207 ne
rect 5866 8157 5959 8207
tri 6251 8167 6294 8210 ne
rect 6294 8167 8288 8210
tri 6294 8164 6297 8167 ne
rect 6297 8164 8288 8167
rect 8608 8221 8660 8227
tri 5959 8157 5966 8164 sw
tri 6297 8158 6303 8164 ne
rect 6303 8158 8340 8164
tri 8602 8158 8608 8164 se
rect 8608 8158 8660 8169
tri 8601 8157 8602 8158 se
rect 8602 8157 8660 8158
rect 5866 8153 5966 8157
tri 5966 8153 5970 8157 sw
tri 8597 8153 8601 8157 se
rect 8601 8153 8608 8157
rect 5866 8130 5970 8153
tri 5970 8130 5993 8153 sw
tri 8574 8130 8597 8153 se
rect 8597 8130 8608 8153
rect 5866 8105 8608 8130
rect 5866 8099 8660 8105
rect 8688 8120 8740 8126
tri 5695 8078 5703 8086 sw
rect 5866 8084 8642 8099
tri 8642 8084 8657 8099 nw
rect 5866 8078 8636 8084
tri 8636 8078 8642 8084 nw
tri 8682 8078 8688 8084 se
rect 5643 8068 5703 8078
tri 5703 8068 5713 8078 sw
tri 8672 8068 8682 8078 se
rect 8682 8068 8688 8078
rect 5643 8064 5713 8068
tri 5643 8056 5651 8064 ne
rect 5651 8056 5713 8064
tri 5713 8056 5725 8068 sw
tri 8660 8056 8672 8068 se
rect 8672 8056 8740 8068
tri 5651 8050 5657 8056 ne
rect 5657 8050 5725 8056
tri 5725 8050 5731 8056 sw
tri 8654 8050 8660 8056 se
rect 8660 8050 8688 8056
tri 5657 8012 5695 8050 ne
rect 5695 8012 8688 8050
tri 5695 8004 5703 8012 ne
rect 5703 8004 8688 8012
tri 5703 7998 5709 8004 ne
rect 5709 7998 8740 8004
rect 1414 7971 5465 7972
rect 628 7970 5465 7971
rect 5823 7937 7104 7938
rect 5823 7881 5832 7937
rect 5888 7881 5913 7937
rect 5969 7881 5994 7937
rect 6050 7881 6075 7937
rect 6131 7881 6156 7937
rect 6212 7881 6237 7937
rect 6293 7881 6318 7937
rect 6374 7881 6398 7937
rect 6454 7881 6478 7937
rect 6534 7881 6558 7937
rect 6614 7885 6950 7937
rect 7002 7885 7046 7937
rect 7098 7885 7104 7937
rect 6614 7881 7104 7885
rect 5823 7845 7104 7881
rect 5823 7789 5832 7845
rect 5888 7789 5913 7845
rect 5969 7789 5994 7845
rect 6050 7789 6075 7845
rect 6131 7789 6156 7845
rect 6212 7789 6237 7845
rect 6293 7789 6318 7845
rect 6374 7789 6398 7845
rect 6454 7789 6478 7845
rect 6534 7789 6558 7845
rect 6614 7841 7104 7845
rect 6614 7789 6950 7841
rect 7002 7789 7046 7841
rect 7098 7789 7104 7841
rect 282 7756 3543 7765
rect 282 7723 2714 7756
rect 282 7667 291 7723
rect 347 7667 374 7723
rect 430 7667 456 7723
rect 512 7667 538 7723
rect 594 7667 620 7723
rect 676 7667 702 7723
rect 758 7667 784 7723
rect 840 7667 866 7723
rect 922 7667 948 7723
rect 1004 7667 1030 7723
rect 1086 7667 1112 7723
rect 1168 7667 1194 7723
rect 1250 7667 1276 7723
rect 1332 7667 1358 7723
rect 1414 7700 2714 7723
rect 2770 7700 2794 7756
rect 2850 7700 2874 7756
rect 2930 7700 2954 7756
rect 3010 7700 3034 7756
rect 3090 7700 3114 7756
rect 3170 7700 3194 7756
rect 3250 7700 3274 7756
rect 3330 7700 3354 7756
rect 3410 7700 3434 7756
rect 3490 7700 3543 7756
rect 1414 7672 3543 7700
rect 1414 7667 2714 7672
rect 282 7637 2714 7667
rect 282 7581 291 7637
rect 347 7581 374 7637
rect 430 7581 456 7637
rect 512 7581 538 7637
rect 594 7581 620 7637
rect 676 7581 702 7637
rect 758 7581 784 7637
rect 840 7581 866 7637
rect 922 7581 948 7637
rect 1004 7581 1030 7637
rect 1086 7581 1112 7637
rect 1168 7581 1194 7637
rect 1250 7581 1276 7637
rect 1332 7581 1358 7637
rect 1414 7616 2714 7637
rect 2770 7616 2794 7672
rect 2850 7616 2874 7672
rect 2930 7616 2954 7672
rect 3010 7616 3034 7672
rect 3090 7616 3114 7672
rect 3170 7616 3194 7672
rect 3250 7616 3274 7672
rect 3330 7616 3354 7672
rect 3410 7616 3434 7672
rect 3490 7616 3543 7672
rect 1414 7588 3543 7616
rect 1414 7581 2714 7588
rect 282 7551 2714 7581
rect 282 7495 291 7551
rect 347 7495 374 7551
rect 430 7495 456 7551
rect 512 7495 538 7551
rect 594 7495 620 7551
rect 676 7495 702 7551
rect 758 7495 784 7551
rect 840 7495 866 7551
rect 922 7495 948 7551
rect 1004 7495 1030 7551
rect 1086 7495 1112 7551
rect 1168 7495 1194 7551
rect 1250 7495 1276 7551
rect 1332 7495 1358 7551
rect 1414 7532 2714 7551
rect 2770 7532 2794 7588
rect 2850 7532 2874 7588
rect 2930 7532 2954 7588
rect 3010 7532 3034 7588
rect 3090 7532 3114 7588
rect 3170 7532 3194 7588
rect 3250 7532 3274 7588
rect 3330 7532 3354 7588
rect 3410 7532 3434 7588
rect 3490 7532 3543 7588
rect 1414 7504 3543 7532
rect 1414 7495 2714 7504
rect 282 7465 2714 7495
rect 282 7409 291 7465
rect 347 7409 374 7465
rect 430 7409 456 7465
rect 512 7409 538 7465
rect 594 7409 620 7465
rect 676 7409 702 7465
rect 758 7409 784 7465
rect 840 7409 866 7465
rect 922 7409 948 7465
rect 1004 7409 1030 7465
rect 1086 7409 1112 7465
rect 1168 7409 1194 7465
rect 1250 7409 1276 7465
rect 1332 7409 1358 7465
rect 1414 7448 2714 7465
rect 2770 7448 2794 7504
rect 2850 7448 2874 7504
rect 2930 7448 2954 7504
rect 3010 7448 3034 7504
rect 3090 7448 3114 7504
rect 3170 7448 3194 7504
rect 3250 7448 3274 7504
rect 3330 7448 3354 7504
rect 3410 7448 3434 7504
rect 3490 7448 3543 7504
rect 1414 7420 3543 7448
rect 1414 7409 2714 7420
rect 282 7379 2714 7409
rect 282 7323 291 7379
rect 347 7323 374 7379
rect 430 7323 456 7379
rect 512 7323 538 7379
rect 594 7323 620 7379
rect 676 7323 702 7379
rect 758 7323 784 7379
rect 840 7323 866 7379
rect 922 7323 948 7379
rect 1004 7323 1030 7379
rect 1086 7323 1112 7379
rect 1168 7323 1194 7379
rect 1250 7323 1276 7379
rect 1332 7323 1358 7379
rect 1414 7364 2714 7379
rect 2770 7364 2794 7420
rect 2850 7364 2874 7420
rect 2930 7364 2954 7420
rect 3010 7364 3034 7420
rect 3090 7364 3114 7420
rect 3170 7364 3194 7420
rect 3250 7364 3274 7420
rect 3330 7364 3354 7420
rect 3410 7364 3434 7420
rect 3490 7364 3543 7420
rect 1414 7336 3543 7364
rect 1414 7323 2714 7336
rect 282 7293 2714 7323
rect 282 7237 291 7293
rect 347 7237 374 7293
rect 430 7237 456 7293
rect 512 7237 538 7293
rect 594 7237 620 7293
rect 676 7237 702 7293
rect 758 7237 784 7293
rect 840 7237 866 7293
rect 922 7237 948 7293
rect 1004 7237 1030 7293
rect 1086 7237 1112 7293
rect 1168 7237 1194 7293
rect 1250 7237 1276 7293
rect 1332 7237 1358 7293
rect 1414 7280 2714 7293
rect 2770 7280 2794 7336
rect 2850 7280 2874 7336
rect 2930 7280 2954 7336
rect 3010 7280 3034 7336
rect 3090 7280 3114 7336
rect 3170 7280 3194 7336
rect 3250 7280 3274 7336
rect 3330 7280 3354 7336
rect 3410 7280 3434 7336
rect 3490 7280 3543 7336
rect 1414 7252 3543 7280
rect 1414 7237 2714 7252
rect 282 7207 2714 7237
rect 282 7151 291 7207
rect 347 7151 374 7207
rect 430 7151 456 7207
rect 512 7151 538 7207
rect 594 7151 620 7207
rect 676 7151 702 7207
rect 758 7151 784 7207
rect 840 7151 866 7207
rect 922 7151 948 7207
rect 1004 7151 1030 7207
rect 1086 7151 1112 7207
rect 1168 7151 1194 7207
rect 1250 7151 1276 7207
rect 1332 7151 1358 7207
rect 1414 7196 2714 7207
rect 2770 7196 2794 7252
rect 2850 7196 2874 7252
rect 2930 7196 2954 7252
rect 3010 7196 3034 7252
rect 3090 7196 3114 7252
rect 3170 7196 3194 7252
rect 3250 7196 3274 7252
rect 3330 7196 3354 7252
rect 3410 7196 3434 7252
rect 3490 7196 3543 7252
rect 1414 7168 3543 7196
rect 6840 7339 7576 7345
rect 6840 7336 7500 7339
rect 6896 7287 7500 7336
rect 7552 7287 7576 7339
rect 6896 7280 7576 7287
rect 6840 7256 7576 7280
rect 6896 7249 7576 7256
rect 6896 7200 7500 7249
rect 6840 7197 7500 7200
rect 7552 7197 7576 7249
rect 6840 7191 7576 7197
rect 1414 7151 2714 7168
rect 282 7121 2714 7151
rect 282 7065 291 7121
rect 347 7065 374 7121
rect 430 7065 456 7121
rect 512 7065 538 7121
rect 594 7065 620 7121
rect 676 7065 702 7121
rect 758 7065 784 7121
rect 840 7065 866 7121
rect 922 7065 948 7121
rect 1004 7065 1030 7121
rect 1086 7065 1112 7121
rect 1168 7065 1194 7121
rect 1250 7065 1276 7121
rect 1332 7065 1358 7121
rect 1414 7112 2714 7121
rect 2770 7112 2794 7168
rect 2850 7112 2874 7168
rect 2930 7112 2954 7168
rect 3010 7112 3034 7168
rect 3090 7112 3114 7168
rect 3170 7112 3194 7168
rect 3250 7112 3274 7168
rect 3330 7112 3354 7168
rect 3410 7112 3434 7168
rect 3490 7112 3543 7168
rect 1414 7084 3543 7112
rect 1414 7065 2714 7084
rect 282 7035 2714 7065
rect 282 6979 291 7035
rect 347 6979 374 7035
rect 430 6979 456 7035
rect 512 6979 538 7035
rect 594 6979 620 7035
rect 676 6979 702 7035
rect 758 6979 784 7035
rect 840 6979 866 7035
rect 922 6979 948 7035
rect 1004 6979 1030 7035
rect 1086 6979 1112 7035
rect 1168 6979 1194 7035
rect 1250 6979 1276 7035
rect 1332 6979 1358 7035
rect 1414 7028 2714 7035
rect 2770 7028 2794 7084
rect 2850 7028 2874 7084
rect 2930 7028 2954 7084
rect 3010 7028 3034 7084
rect 3090 7028 3114 7084
rect 3170 7028 3194 7084
rect 3250 7028 3274 7084
rect 3330 7028 3354 7084
rect 3410 7028 3434 7084
rect 3490 7028 3543 7084
rect 1414 7000 3543 7028
rect 1414 6979 2714 7000
rect 282 6949 2714 6979
rect 282 6893 291 6949
rect 347 6893 374 6949
rect 430 6893 456 6949
rect 512 6893 538 6949
rect 594 6893 620 6949
rect 676 6893 702 6949
rect 758 6893 784 6949
rect 840 6893 866 6949
rect 922 6893 948 6949
rect 1004 6893 1030 6949
rect 1086 6893 1112 6949
rect 1168 6893 1194 6949
rect 1250 6893 1276 6949
rect 1332 6893 1358 6949
rect 1414 6944 2714 6949
rect 2770 6944 2794 7000
rect 2850 6944 2874 7000
rect 2930 6944 2954 7000
rect 3010 6944 3034 7000
rect 3090 6944 3114 7000
rect 3170 6944 3194 7000
rect 3250 6944 3274 7000
rect 3330 6944 3354 7000
rect 3410 6944 3434 7000
rect 3490 6944 3543 7000
rect 1414 6915 3543 6944
rect 6714 7062 6770 7071
rect 6714 6987 6770 7006
rect 7618 7039 7670 7045
tri 6770 6987 6786 7003 sw
tri 7602 6987 7618 7003 se
rect 6714 6982 6786 6987
rect 6770 6975 6786 6982
tri 6786 6975 6798 6987 sw
tri 7590 6975 7602 6987 se
rect 7602 6975 7670 6987
rect 6770 6969 6798 6975
tri 6798 6969 6804 6975 sw
tri 7584 6969 7590 6975 se
rect 7590 6969 7618 6975
rect 6770 6926 7618 6969
rect 6714 6923 7618 6926
rect 6714 6917 7670 6923
rect 1414 6893 2714 6915
rect 282 6863 2714 6893
rect 282 6807 291 6863
rect 347 6807 374 6863
rect 430 6807 456 6863
rect 512 6807 538 6863
rect 594 6807 620 6863
rect 676 6807 702 6863
rect 758 6807 784 6863
rect 840 6807 866 6863
rect 922 6807 948 6863
rect 1004 6807 1030 6863
rect 1086 6807 1112 6863
rect 1168 6807 1194 6863
rect 1250 6807 1276 6863
rect 1332 6807 1358 6863
rect 1414 6859 2714 6863
rect 2770 6859 2794 6915
rect 2850 6859 2874 6915
rect 2930 6859 2954 6915
rect 3010 6859 3034 6915
rect 3090 6859 3114 6915
rect 3170 6859 3194 6915
rect 3250 6859 3274 6915
rect 3330 6859 3354 6915
rect 3410 6859 3434 6915
rect 3490 6859 3543 6915
rect 1414 6830 3543 6859
rect 1414 6807 2714 6830
rect 282 6774 2714 6807
rect 2770 6774 2794 6830
rect 2850 6774 2874 6830
rect 2930 6774 2954 6830
rect 3010 6774 3034 6830
rect 3090 6774 3114 6830
rect 3170 6774 3194 6830
rect 3250 6774 3274 6830
rect 3330 6774 3354 6830
rect 3410 6774 3434 6830
rect 3490 6774 3543 6830
rect 282 6765 3543 6774
tri 5861 6519 5895 6553 sw
tri 8094 6519 8128 6553 se
tri 5666 6342 5727 6403 se
rect 5727 6351 7318 6403
rect 5727 6342 5740 6351
tri 5740 6342 5749 6351 nw
tri 7296 6342 7305 6351 ne
rect 7305 6342 7318 6351
tri 7318 6342 7379 6403 sw
tri 5653 6329 5666 6342 se
rect 5666 6329 5727 6342
tri 5727 6329 5740 6342 nw
tri 7305 6329 7318 6342 ne
rect 7318 6329 7379 6342
tri 5642 6318 5653 6329 se
rect 5653 6318 5716 6329
tri 5716 6318 5727 6329 nw
tri 7318 6318 7329 6329 ne
rect 7329 6318 7379 6329
rect 2373 6312 5666 6318
rect 2425 6268 5666 6312
tri 5666 6268 5716 6318 nw
tri 7329 6268 7379 6318 ne
tri 7379 6268 7453 6342 sw
rect 2425 6266 5664 6268
tri 5664 6266 5666 6268 nw
tri 7379 6266 7381 6268 ne
rect 7381 6266 7667 6268
rect 2425 6262 2455 6266
tri 2455 6262 2459 6266 nw
tri 7381 6262 7385 6266 ne
rect 7385 6262 7667 6266
rect 2373 6248 2425 6260
tri 2425 6232 2455 6262 nw
tri 7385 6232 7415 6262 ne
rect 7415 6232 7615 6262
tri 7415 6216 7431 6232 ne
rect 7431 6216 7615 6232
tri 7581 6210 7587 6216 ne
rect 7587 6210 7615 6216
tri 7587 6198 7599 6210 ne
rect 7599 6198 7667 6210
rect 2373 6190 2425 6196
tri 7599 6190 7607 6198 ne
rect 7607 6190 7615 6198
tri 7607 6182 7615 6190 ne
rect 7615 6140 7667 6146
rect 6507 6127 7104 6133
rect 6507 6124 6944 6127
rect 6563 6068 6587 6124
rect 6643 6075 6944 6124
rect 6996 6075 7052 6127
rect 6643 6068 7104 6075
rect 6507 6057 7104 6068
rect 6507 6032 6944 6057
rect 6563 5976 6587 6032
rect 6643 6005 6944 6032
rect 6996 6005 7052 6057
rect 6643 5987 7104 6005
rect 6643 5976 6944 5987
rect 6507 5940 6944 5976
rect 6563 5884 6587 5940
rect 6643 5935 6944 5940
rect 6996 5935 7052 5987
rect 6643 5917 7104 5935
rect 6643 5884 6944 5917
rect 6507 5865 6944 5884
rect 6996 5865 7052 5917
tri 7104 5908 7329 6133 sw
rect 7104 5902 7756 5908
rect 7104 5865 7704 5902
rect 6507 5850 7704 5865
rect 6507 5848 7756 5850
rect 6563 5792 6587 5848
rect 6643 5847 7756 5848
rect 6643 5795 6944 5847
rect 6996 5795 7052 5847
rect 7104 5835 7756 5847
rect 7104 5795 7704 5835
rect 6643 5792 7704 5795
rect 6507 5783 7704 5792
rect 6507 5777 7756 5783
rect 6507 5756 6944 5777
rect 6563 5700 6587 5756
rect 6643 5725 6944 5756
rect 6996 5725 7052 5777
rect 7104 5768 7756 5777
rect 7104 5725 7704 5768
rect 6643 5716 7704 5725
rect 6643 5706 7756 5716
rect 6643 5700 6944 5706
rect 6507 5664 6944 5700
rect 6563 5608 6587 5664
rect 6643 5654 6944 5664
rect 6996 5654 7052 5706
rect 7104 5700 7756 5706
rect 7104 5654 7704 5700
rect 6643 5648 7704 5654
rect 6643 5635 7756 5648
rect 6643 5608 6944 5635
rect 6507 5583 6944 5608
rect 6996 5583 7052 5635
rect 7104 5632 7756 5635
rect 7104 5583 7704 5632
rect 6507 5580 7704 5583
rect 6507 5571 7756 5580
rect 6563 5515 6587 5571
rect 6643 5564 7756 5571
rect 6643 5515 6944 5564
rect 6507 5512 6944 5515
rect 6996 5512 7052 5564
rect 7104 5512 7704 5564
rect 6507 5506 7756 5512
rect 7524 5240 10317 5246
rect 7576 5237 10317 5240
rect 7576 5188 10261 5237
rect 7524 5181 10261 5188
rect 7524 5157 10317 5181
rect 7524 5150 10261 5157
rect 7576 5101 10261 5150
rect 7576 5098 10317 5101
rect 7524 5092 10317 5098
rect 8932 5010 8984 5016
rect 7618 4990 7670 4996
tri 7670 4958 7686 4974 sw
tri 8916 4958 8932 4974 se
rect 7670 4946 7686 4958
tri 7686 4946 7698 4958 sw
tri 8904 4946 8916 4958 se
rect 8916 4946 8984 4958
rect 7670 4940 7698 4946
tri 7698 4940 7704 4946 sw
tri 8898 4940 8904 4946 se
rect 8904 4940 8932 4946
rect 7670 4938 8932 4940
rect 7618 4926 8932 4938
rect 7670 4894 8932 4926
rect 7670 4888 8984 4894
rect 7618 4868 7670 4874
tri 7670 4868 7690 4888 nw
rect 8772 4524 8824 4530
tri 8756 4472 8772 4488 se
tri 8744 4460 8756 4472 se
rect 8756 4460 8824 4472
tri 8738 4454 8744 4460 se
rect 8744 4454 8772 4460
rect 7615 4448 8772 4454
rect 7667 4408 8772 4448
rect 7667 4402 8824 4408
rect 7615 4384 7667 4396
tri 7667 4368 7701 4402 nw
rect 7615 4326 7667 4332
tri 6471 4219 6477 4225 ne
tri 6605 4219 6611 4225 nw
rect 6458 4054 7104 4060
rect 6458 4051 6944 4054
rect 1639 3994 1691 4000
rect 6458 3995 6459 4051
rect 6515 3995 6561 4051
rect 6617 3995 6663 4051
rect 6719 4002 6944 4051
rect 6996 4002 7052 4054
rect 6719 3995 7104 4002
rect 6458 3987 7104 3995
rect 6458 3970 6944 3987
rect 1639 3935 1691 3942
tri 1691 3935 1714 3958 sw
rect 1639 3930 1714 3935
rect 1691 3924 1714 3930
tri 1714 3924 1725 3935 sw
rect 1691 3878 5552 3924
rect 1639 3872 5552 3878
rect 5604 3872 5616 3924
rect 5668 3872 5674 3924
rect 6458 3914 6459 3970
rect 6515 3914 6561 3970
rect 6617 3914 6663 3970
rect 6719 3935 6944 3970
rect 6996 3935 7052 3987
rect 6719 3920 7104 3935
rect 6719 3914 6944 3920
rect 6458 3889 6944 3914
rect 2707 3837 5427 3843
rect 2759 3791 5427 3837
rect 5479 3791 5491 3843
rect 5543 3791 5549 3843
rect 6458 3833 6459 3889
rect 6515 3833 6561 3889
rect 6617 3833 6663 3889
rect 6719 3868 6944 3889
rect 6996 3868 7052 3920
rect 6719 3853 7104 3868
rect 6719 3833 6944 3853
rect 6458 3807 6944 3833
rect 2759 3786 2788 3791
tri 2788 3786 2793 3791 nw
rect 2707 3760 2759 3785
tri 2759 3757 2788 3786 nw
rect 2707 3683 2759 3708
rect 6458 3751 6459 3807
rect 6515 3751 6561 3807
rect 6617 3751 6663 3807
rect 6719 3801 6944 3807
rect 6996 3801 7052 3853
rect 6719 3786 7104 3801
rect 6719 3751 6944 3786
rect 6458 3734 6944 3751
rect 6996 3734 7052 3786
rect 6458 3725 7104 3734
rect 6458 3669 6459 3725
rect 6515 3669 6561 3725
rect 6617 3669 6663 3725
rect 6719 3718 7104 3725
rect 7615 3871 8084 3878
rect 7667 3869 8084 3871
rect 7667 3819 8023 3869
rect 7615 3813 8023 3819
rect 8079 3813 8084 3869
rect 7615 3807 8084 3813
rect 7667 3789 8084 3807
rect 7667 3755 8023 3789
rect 7615 3733 8023 3755
rect 8079 3733 8084 3789
rect 7615 3724 8084 3733
rect 6719 3669 6944 3718
rect 6458 3666 6944 3669
rect 6996 3666 7052 3718
rect 6458 3660 7104 3666
rect 7823 3687 7875 3693
rect 2707 3606 2759 3631
tri 2759 3606 2787 3634 sw
tri 7795 3606 7823 3634 se
rect 7823 3606 7875 3635
rect 2627 3551 2679 3557
rect 2759 3600 2787 3606
tri 2787 3600 2793 3606 sw
tri 7789 3600 7795 3606 se
rect 7795 3600 7823 3606
rect 2759 3554 4369 3600
rect 2707 3548 4369 3554
rect 4421 3548 4433 3600
rect 4485 3548 4491 3600
rect 4827 3548 4833 3600
rect 4885 3548 4897 3600
rect 4949 3548 4955 3600
rect 5401 3548 5407 3600
rect 5459 3548 5491 3600
rect 5543 3554 7823 3600
rect 5543 3548 7875 3554
tri 4805 3525 4827 3547 se
rect 4827 3525 4879 3548
tri 4879 3525 4902 3548 nw
tri 4795 3515 4805 3525 se
rect 4805 3515 4869 3525
tri 4869 3515 4879 3525 nw
rect 2627 3487 2679 3499
rect 1733 3471 1785 3477
tri 2679 3481 2713 3515 sw
tri 4783 3503 4795 3515 se
rect 4795 3503 4857 3515
tri 4857 3503 4869 3515 nw
tri 4761 3481 4783 3503 se
rect 4783 3481 4835 3503
tri 4835 3481 4857 3503 nw
rect 2679 3435 4306 3481
rect 1733 3407 1785 3419
tri 1785 3401 1819 3435 sw
rect 2627 3429 4306 3435
rect 4358 3429 4370 3481
rect 4422 3435 4789 3481
tri 4789 3435 4835 3481 nw
rect 4422 3429 4783 3435
tri 4783 3429 4789 3435 nw
rect 1785 3355 4630 3401
rect 1733 3349 4630 3355
rect 4682 3349 4694 3401
rect 4746 3349 4926 3401
rect 4978 3349 4990 3401
rect 5042 3349 5048 3401
rect 5245 3349 5251 3401
rect 5303 3349 5315 3401
rect 5367 3349 5552 3401
rect 5604 3349 5616 3401
rect 5668 3349 5674 3401
rect 4195 3315 5832 3321
rect 4195 3263 4499 3315
rect 4551 3263 4811 3315
rect 4863 3263 5123 3315
rect 5175 3263 5435 3315
rect 5487 3263 5747 3315
rect 5799 3265 5832 3315
rect 5888 3265 5914 3321
rect 5970 3265 5995 3321
rect 6051 3265 6076 3321
rect 6132 3265 6157 3321
rect 6213 3265 6238 3321
rect 6294 3265 6319 3321
rect 6375 3265 6400 3321
rect 6456 3265 6481 3321
rect 6537 3265 6562 3321
rect 6618 3315 7106 3321
rect 6618 3265 6944 3315
rect 5799 3263 6944 3265
rect 6996 3263 7052 3315
rect 7104 3263 7106 3315
rect 4195 3251 7106 3263
rect 4195 3199 4499 3251
rect 4551 3199 4811 3251
rect 4863 3199 5123 3251
rect 5175 3199 5435 3251
rect 5487 3199 5747 3251
rect 5799 3244 7106 3251
rect 5799 3241 6944 3244
rect 5799 3199 5832 3241
rect 4195 3193 5832 3199
tri 5589 3192 5590 3193 ne
rect 5590 3192 5832 3193
tri 5590 3172 5610 3192 ne
rect 5610 3185 5832 3192
rect 5888 3185 5914 3241
rect 5970 3185 5995 3241
rect 6051 3185 6076 3241
rect 6132 3185 6157 3241
rect 6213 3185 6238 3241
rect 6294 3185 6319 3241
rect 6375 3185 6400 3241
rect 6456 3185 6481 3241
rect 6537 3185 6562 3241
rect 6618 3192 6944 3241
rect 6996 3192 7052 3244
rect 7104 3192 7106 3244
rect 6618 3185 7106 3192
rect 5610 3172 7106 3185
tri 5610 3159 5623 3172 ne
rect 5623 3137 6944 3172
rect 5623 3136 5832 3137
rect 5888 3136 5914 3137
rect 5970 3136 5995 3137
rect 6051 3136 6076 3137
rect 6132 3136 6157 3137
rect 6213 3136 6238 3137
rect 6294 3136 6319 3137
rect 6375 3136 6400 3137
rect 6456 3136 6481 3137
rect 6537 3136 6562 3137
rect 5623 3084 5629 3136
rect 5681 3084 5696 3136
rect 5748 3084 5763 3136
rect 5815 3084 5830 3136
rect 5888 3084 5897 3136
rect 6150 3084 6157 3136
rect 6217 3084 6232 3136
rect 6294 3084 6299 3136
rect 6551 3084 6562 3136
rect 6618 3120 6944 3137
rect 6996 3120 7052 3172
rect 7104 3120 7106 3172
rect 7524 3295 8977 3304
rect 7524 3272 8916 3295
rect 7576 3239 8916 3272
rect 8972 3239 8977 3295
rect 7576 3220 8977 3239
rect 7524 3215 8977 3220
rect 7524 3208 8916 3215
rect 7576 3159 8916 3208
rect 8972 3159 8977 3215
rect 7576 3156 8977 3159
rect 7524 3150 8977 3156
rect 6618 3100 7106 3120
rect 5623 3081 5832 3084
rect 5888 3081 5914 3084
rect 5970 3081 5995 3084
rect 6051 3081 6076 3084
rect 6132 3081 6157 3084
rect 6213 3081 6238 3084
rect 6294 3081 6319 3084
rect 6375 3081 6400 3084
rect 6456 3081 6481 3084
rect 6537 3081 6562 3084
rect 6618 3081 6944 3100
rect 5623 3057 6944 3081
rect 5623 3048 5832 3057
rect 5888 3048 5914 3057
rect 5970 3048 5995 3057
rect 6051 3048 6076 3057
rect 6132 3048 6157 3057
rect 6213 3048 6238 3057
rect 6294 3048 6319 3057
rect 6375 3048 6400 3057
rect 6456 3048 6481 3057
rect 6537 3048 6562 3057
rect 6618 3048 6944 3057
rect 6996 3048 7052 3100
rect 7104 3048 7106 3100
rect 8772 3101 8824 3107
tri 8756 3049 8772 3065 se
rect 5623 2996 5629 3048
rect 5681 2996 5696 3048
rect 5748 2996 5763 3048
rect 5815 2996 5830 3048
rect 5888 3001 5897 3048
rect 6150 3001 6157 3048
rect 5882 2996 5897 3001
rect 5949 2996 5964 3001
rect 6016 2996 6031 3001
rect 6083 2996 6098 3001
rect 6150 2996 6165 3001
rect 6217 2996 6232 3048
rect 6294 3001 6299 3048
rect 6551 3001 6562 3048
rect 6618 3028 7106 3048
tri 8744 3037 8756 3049 se
rect 8756 3037 8824 3049
tri 8738 3031 8744 3037 se
rect 8744 3031 8772 3037
rect 6618 3001 6944 3028
rect 6284 2996 6299 3001
rect 6351 2996 6366 3001
rect 6418 2996 6433 3001
rect 6485 2996 6499 3001
rect 6551 2996 6565 3001
rect 6617 2996 6944 3001
rect 5623 2976 6944 2996
rect 6996 2976 7052 3028
rect 7104 2976 7106 3028
rect 5623 2970 7106 2976
rect 7639 2985 8772 3031
rect 7639 2979 8824 2985
rect 7639 2975 7721 2979
tri 7721 2975 7725 2979 nw
tri 7634 2970 7639 2975 se
rect 7639 2970 7691 2975
tri 7605 2941 7634 2970 se
rect 7634 2941 7691 2970
tri 7691 2945 7721 2975 nw
rect 2373 2928 2425 2934
rect 2293 2877 2345 2883
rect 2293 2813 2345 2825
tri 2425 2889 2428 2892 sw
rect 4914 2889 7691 2941
rect 7903 2931 7955 2937
tri 7900 2892 7903 2895 se
tri 7897 2889 7900 2892 se
rect 7900 2889 7903 2892
rect 2425 2879 2428 2889
tri 2428 2879 2438 2889 sw
rect 4914 2879 5066 2889
tri 5066 2879 5076 2889 nw
tri 7887 2879 7897 2889 se
rect 7897 2879 7903 2889
rect 2425 2876 2438 2879
rect 2373 2867 2438 2876
tri 2438 2867 2450 2879 sw
rect 4914 2867 5054 2879
tri 5054 2867 5066 2879 nw
tri 7875 2867 7887 2879 se
rect 7887 2867 7955 2879
rect 2373 2864 2450 2867
rect 2425 2861 2450 2864
tri 2450 2861 2456 2867 sw
rect 4914 2861 5048 2867
tri 5048 2861 5054 2867 nw
tri 7869 2861 7875 2867 se
rect 7875 2861 7903 2867
rect 2425 2858 2456 2861
tri 2456 2858 2459 2861 sw
rect 2425 2812 3610 2858
rect 2373 2806 3610 2812
rect 3662 2806 3674 2858
rect 3726 2806 3732 2858
rect 4914 2809 4920 2861
rect 4972 2809 4984 2861
rect 5036 2809 5042 2861
tri 5042 2855 5048 2861 nw
rect 5976 2809 5982 2861
rect 6034 2809 6046 2861
rect 6098 2815 7903 2861
rect 6098 2809 7955 2815
rect 8208 2880 8260 2886
rect 8208 2816 8260 2828
tri 8205 2789 8208 2792 se
tri 2345 2764 2370 2789 sw
tri 8180 2764 8205 2789 se
rect 8205 2764 8208 2789
rect 2345 2761 2370 2764
rect 2293 2758 2370 2761
tri 2370 2758 2376 2764 sw
tri 8174 2758 8180 2764 se
rect 8180 2758 8260 2764
rect 2293 2755 2376 2758
tri 2376 2755 2379 2758 sw
tri 2293 2751 2297 2755 ne
rect 2297 2751 3712 2755
rect 1632 2744 1945 2750
rect 1684 2692 1893 2744
rect 1632 2680 1945 2692
rect 1684 2628 1893 2680
rect 2213 2745 2265 2751
tri 2297 2750 2298 2751 ne
rect 2298 2750 3712 2751
tri 2298 2743 2305 2750 ne
rect 2305 2743 3712 2750
tri 2305 2731 2317 2743 ne
tri 2265 2703 2271 2709 sw
rect 2317 2703 3712 2743
rect 3764 2703 3776 2755
rect 3828 2703 3834 2755
rect 4577 2737 4629 2743
rect 2265 2693 2271 2703
rect 2213 2685 2271 2693
tri 2271 2685 2289 2703 sw
rect 5874 2706 5880 2758
rect 5932 2706 5944 2758
rect 5996 2755 8257 2758
tri 8257 2755 8260 2758 nw
rect 5996 2750 8252 2755
tri 8252 2750 8257 2755 nw
rect 5996 2748 8250 2750
tri 8250 2748 8252 2750 nw
rect 8288 2748 8340 2754
rect 5996 2743 8245 2748
tri 8245 2743 8250 2748 nw
rect 5996 2706 8236 2743
tri 8236 2734 8245 2743 nw
tri 8282 2706 8288 2712 se
tri 8272 2696 8282 2706 se
rect 8282 2696 8288 2706
rect 2213 2684 2289 2685
tri 2289 2684 2290 2685 sw
rect 2213 2681 2290 2684
rect 1632 2622 1945 2628
rect 2053 2661 2105 2667
rect 2265 2678 2290 2681
tri 2290 2678 2296 2684 sw
rect 2265 2675 2296 2678
tri 2296 2675 2299 2678 sw
rect 2265 2629 3232 2675
tri 2105 2623 2107 2625 sw
rect 2213 2623 3232 2629
rect 3284 2623 3296 2675
rect 3348 2623 3354 2675
rect 4264 2672 4316 2678
rect 2105 2622 2107 2623
tri 2107 2622 2108 2623 sw
rect 2105 2620 2108 2622
tri 2108 2620 2110 2622 sw
rect 4577 2673 4629 2685
tri 8260 2684 8272 2696 se
rect 8272 2684 8340 2696
tri 8254 2678 8260 2684 se
rect 8260 2678 8288 2684
tri 4316 2622 4330 2636 sw
rect 4316 2621 4330 2622
tri 4330 2621 4331 2622 sw
rect 6354 2626 6360 2678
rect 6412 2626 6424 2678
rect 6476 2632 8288 2678
rect 6476 2626 8340 2632
rect 8448 2716 8500 2722
rect 8448 2652 8500 2664
tri 8446 2626 8448 2628 se
rect 4316 2620 4331 2621
rect 2105 2609 2110 2620
rect 2053 2608 2110 2609
tri 2110 2608 2122 2620 sw
rect 4264 2608 4331 2620
rect 2053 2602 2122 2608
tri 2122 2602 2128 2608 sw
rect 2053 2597 2128 2602
rect 2105 2591 2128 2597
tri 2128 2591 2139 2602 sw
rect 2105 2545 2923 2591
rect 2053 2539 2923 2545
rect 2975 2539 2987 2591
rect 3039 2539 3045 2591
rect 4316 2602 4331 2608
tri 4331 2602 4350 2621 sw
rect 4316 2600 4477 2602
tri 4477 2600 4479 2602 sw
rect 4316 2594 4479 2600
tri 4479 2594 4485 2600 sw
rect 4316 2591 4485 2594
tri 4485 2591 4488 2594 sw
rect 4316 2556 4488 2591
rect 4264 2550 4488 2556
tri 4455 2546 4459 2550 ne
rect 4459 2546 4488 2550
tri 4488 2546 4533 2591 sw
tri 4459 2542 4463 2546 ne
rect 4463 2542 4533 2546
tri 4463 2539 4466 2542 ne
rect 4466 2539 4533 2542
tri 4466 2528 4477 2539 ne
rect 4477 2528 4533 2539
tri 4477 2524 4481 2528 ne
tri 4288 2500 4291 2503 se
rect 4291 2500 4297 2503
tri 2120 2487 2133 2500 se
rect 2133 2487 2987 2500
rect 1973 2447 2025 2453
rect 2057 2435 2063 2487
rect 2115 2435 2127 2487
rect 2179 2448 2987 2487
rect 3039 2448 3053 2500
rect 3105 2451 4297 2500
rect 4349 2451 4363 2503
rect 4415 2451 4421 2503
rect 3105 2448 4387 2451
tri 4387 2448 4390 2451 nw
rect 2179 2447 2197 2448
tri 2197 2447 2198 2448 nw
tri 4270 2447 4271 2448 ne
rect 4271 2447 4386 2448
tri 4386 2447 4387 2448 nw
rect 2179 2441 2191 2447
tri 2191 2441 2197 2447 nw
tri 4271 2441 4277 2447 ne
rect 4277 2441 4380 2447
tri 4380 2441 4386 2447 nw
rect 2179 2435 2185 2441
tri 2185 2435 2191 2441 nw
tri 4277 2435 4283 2441 ne
rect 4283 2435 4374 2441
tri 4374 2435 4380 2441 nw
tri 4283 2429 4289 2435 ne
rect 4289 2429 4368 2435
tri 4368 2429 4374 2435 nw
tri 4289 2417 4301 2429 ne
rect 4301 2417 4356 2429
tri 4356 2417 4368 2429 nw
tri 4301 2414 4304 2417 ne
rect 1973 2383 2025 2395
rect 1632 2367 1684 2373
tri 2025 2377 2059 2411 sw
rect 2025 2331 4122 2377
tri 1684 2327 1688 2331 sw
rect 1684 2325 1688 2327
tri 1688 2325 1690 2327 sw
rect 1973 2325 4122 2331
rect 4174 2325 4186 2377
rect 4238 2325 4244 2377
rect 1684 2315 1690 2325
rect 1632 2303 1690 2315
rect 1684 2297 1690 2303
tri 1690 2297 1718 2325 sw
rect 1684 2251 3805 2297
rect 1632 2245 3805 2251
rect 3857 2245 3869 2297
rect 3921 2245 3927 2297
rect 4304 2217 4356 2417
rect 4481 2327 4533 2528
rect 4577 2379 4629 2621
tri 8420 2600 8446 2626 se
rect 8446 2600 8448 2626
tri 8414 2594 8420 2600 se
rect 8420 2594 8500 2600
rect 6663 2542 6669 2594
rect 6721 2542 6733 2594
rect 6785 2542 8500 2594
rect 4969 2493 5021 2499
tri 5021 2451 5027 2457 sw
rect 6597 2451 6603 2503
rect 6655 2451 6669 2503
rect 6721 2451 8374 2503
rect 8426 2451 8438 2503
rect 8490 2451 8496 2503
rect 8805 2493 8857 2499
tri 8799 2451 8805 2457 se
rect 5021 2441 5027 2451
tri 5027 2441 5037 2451 sw
tri 8789 2441 8799 2451 se
rect 8799 2441 8805 2451
rect 4969 2429 5037 2441
tri 5037 2429 5049 2441 sw
tri 8777 2429 8789 2441 se
rect 8789 2429 8857 2441
tri 4577 2377 4579 2379 ne
rect 4579 2377 4629 2379
tri 4629 2377 4653 2401 sw
rect 5021 2423 5049 2429
tri 5049 2423 5055 2429 sw
tri 8771 2423 8777 2429 se
rect 8777 2423 8805 2429
rect 5021 2377 8805 2423
tri 4579 2343 4613 2377 ne
rect 4613 2343 4653 2377
tri 4653 2343 4687 2377 sw
rect 4969 2371 8857 2377
tri 4613 2328 4628 2343 ne
rect 4628 2328 6780 2343
tri 4533 2327 4534 2328 sw
tri 4628 2327 4629 2328 ne
rect 4629 2327 6780 2328
rect 4481 2325 4534 2327
tri 4534 2325 4536 2327 sw
tri 4629 2325 4631 2327 ne
rect 4631 2325 6780 2327
rect 4481 2306 4536 2325
tri 4481 2297 4490 2306 ne
rect 4490 2297 4536 2306
tri 4536 2297 4564 2325 sw
tri 4631 2297 4659 2325 ne
rect 4659 2297 6780 2325
tri 4490 2291 4496 2297 ne
rect 4496 2291 4564 2297
tri 4564 2291 4570 2297 sw
tri 4659 2291 4665 2297 ne
rect 4665 2291 6780 2297
rect 6832 2291 6844 2343
rect 6896 2291 6902 2343
rect 9092 2333 9144 2339
tri 9086 2291 9092 2297 se
tri 4496 2281 4506 2291 ne
rect 4506 2281 4570 2291
tri 4570 2281 4580 2291 sw
tri 9076 2281 9086 2291 se
rect 9086 2281 9092 2291
tri 4506 2269 4518 2281 ne
rect 4518 2269 4580 2281
tri 4580 2269 4592 2281 sw
tri 9064 2269 9076 2281 se
rect 9076 2269 9144 2281
tri 4518 2263 4524 2269 ne
rect 4524 2263 4592 2269
tri 4592 2263 4598 2269 sw
tri 9058 2263 9064 2269 se
rect 9064 2263 9092 2269
tri 4524 2254 4533 2263 ne
rect 4533 2254 9092 2263
tri 4533 2245 4542 2254 ne
rect 4542 2245 9092 2254
tri 4542 2235 4552 2245 ne
rect 4552 2235 9092 2245
tri 4356 2217 4374 2235 sw
tri 4552 2217 4570 2235 ne
rect 4570 2217 9092 2235
rect 2087 2165 2093 2217
rect 2145 2165 2157 2217
rect 2209 2165 3777 2217
rect 3829 2165 3841 2217
rect 3893 2165 3899 2217
rect 4304 2213 4374 2217
tri 4304 2183 4334 2213 ne
rect 4334 2211 4374 2213
tri 4374 2211 4380 2217 sw
tri 4570 2211 4576 2217 ne
rect 4576 2211 9144 2217
rect 4334 2183 4380 2211
tri 4380 2183 4408 2211 sw
tri 4334 2165 4352 2183 ne
rect 4352 2165 8374 2183
tri 4352 2161 4356 2165 ne
rect 4356 2161 8374 2165
tri 4356 2137 4380 2161 ne
rect 4380 2137 8374 2161
rect 1576 2085 1582 2137
rect 1634 2085 1646 2137
rect 1698 2085 3325 2137
tri 4380 2131 4386 2137 ne
rect 4386 2131 8374 2137
rect 8426 2131 8438 2183
rect 8490 2131 8496 2183
tri 3161 2051 3195 2085 ne
rect 3195 2036 3325 2085
rect 1520 2002 1572 2008
rect 1520 1949 1572 1950
tri 1572 1949 1589 1966 sw
tri 3001 1949 3018 1966 se
rect 3018 1949 3146 1996
rect 3195 1984 3201 2036
rect 3253 1984 3267 2036
rect 3319 1984 3325 2036
rect 3911 1984 3917 2036
rect 3969 1984 3994 2036
rect 4046 1984 4841 2036
tri 4755 1983 4756 1984 ne
rect 4756 1983 4841 1984
tri 3776 1980 3779 1983 ne
rect 3779 1980 3810 1983
tri 4756 1980 4759 1983 ne
rect 4759 1980 4841 1983
tri 4976 1980 4979 1983 ne
rect 4979 1980 5010 1983
tri 5692 1980 5695 1983 ne
rect 5695 1980 5726 1983
rect 5827 1980 5833 2032
rect 5885 1980 5910 2032
rect 5962 1980 6278 2032
rect 6543 1984 6549 2036
rect 6601 1984 6626 2036
rect 6678 1984 8458 2036
rect 8510 1984 8522 2036
rect 8574 1984 8794 2036
rect 8846 1984 8858 2036
rect 8910 1984 8916 2036
tri 6408 1980 6411 1983 ne
rect 6411 1980 6442 1983
tri 3779 1949 3810 1980 ne
tri 4759 1950 4789 1980 ne
rect 1520 1946 1589 1949
tri 1589 1946 1592 1949 sw
tri 2998 1946 3001 1949 se
rect 3001 1946 3146 1949
rect 1520 1942 1592 1946
tri 1592 1942 1596 1946 sw
tri 2994 1942 2998 1946 se
rect 2998 1942 3146 1946
rect 1520 1938 1596 1942
rect 1572 1932 1596 1938
tri 1596 1932 1606 1942 sw
tri 2984 1932 2994 1942 se
rect 2994 1932 3146 1942
rect 3708 1942 3760 1948
rect 1572 1886 3184 1932
rect 1520 1880 3184 1886
rect 3708 1866 3760 1890
tri 3760 1866 3780 1886 sw
rect 4046 1880 4745 1932
tri 4659 1866 4673 1880 ne
rect 4673 1866 4745 1880
rect 3708 1858 3780 1866
tri 3780 1858 3788 1866 sw
tri 4673 1858 4681 1866 ne
rect 4681 1858 4745 1866
rect 1464 1800 2961 1852
rect 3013 1800 3025 1852
rect 3077 1800 3083 1852
rect 3760 1852 3788 1858
tri 3788 1852 3794 1858 sw
tri 4681 1852 4687 1858 ne
rect 4687 1852 4745 1858
rect 3760 1806 4579 1852
tri 4687 1846 4693 1852 ne
rect 3708 1800 4579 1806
rect 1464 1794 1544 1800
tri 1544 1794 1550 1800 nw
tri 4493 1794 4499 1800 ne
rect 4499 1794 4579 1800
rect 1516 1782 1532 1794
tri 1532 1782 1544 1794 nw
tri 4499 1782 4511 1794 ne
rect 4511 1782 4579 1794
tri 1516 1766 1532 1782 nw
tri 4511 1766 4527 1782 ne
rect 1464 1730 1516 1742
rect 1464 1672 1516 1678
rect 1408 1468 1414 1520
rect 1466 1468 1478 1520
rect 1530 1468 2961 1520
rect 3013 1468 3025 1520
rect 3077 1468 3083 1520
rect 3521 1516 4464 1518
rect 3521 1464 3527 1516
rect 3579 1464 3595 1516
rect 3647 1464 3663 1516
rect 3783 1464 3798 1516
rect 3854 1464 3867 1516
rect 4053 1464 4056 1516
rect 4120 1464 4142 1516
rect 3521 1460 3712 1464
rect 3768 1460 3798 1464
rect 3854 1460 3884 1464
rect 3940 1460 3970 1464
rect 4026 1460 4056 1464
rect 4112 1460 4142 1464
rect 4198 1460 4228 1516
rect 4284 1460 4314 1516
rect 4370 1460 4399 1516
rect 4455 1460 4464 1516
rect 3521 1452 4464 1460
rect 1352 1415 3100 1440
rect 1352 1410 3146 1415
rect 1352 1358 1358 1410
rect 1410 1358 1422 1410
rect 1474 1388 3146 1410
rect 1474 1374 1496 1388
tri 1496 1374 1510 1388 nw
tri 2984 1374 2998 1388 ne
rect 2998 1374 3146 1388
rect 1474 1358 1480 1374
tri 1480 1358 1496 1374 nw
tri 2998 1358 3014 1374 ne
rect 3014 1358 3146 1374
tri 3014 1354 3018 1358 ne
rect 3018 1334 3146 1358
rect 3521 1400 3527 1452
rect 3579 1400 3595 1452
rect 3647 1400 3663 1452
rect 3715 1432 3731 1452
rect 3783 1432 3799 1452
rect 3851 1432 3867 1452
rect 3919 1432 3934 1452
rect 3986 1432 4001 1452
rect 4053 1432 4068 1452
rect 4120 1432 4464 1452
rect 3783 1400 3798 1432
rect 3854 1400 3867 1432
rect 4053 1400 4056 1432
rect 4120 1400 4142 1432
rect 3521 1388 3712 1400
rect 3768 1388 3798 1400
rect 3854 1388 3884 1400
rect 3940 1388 3970 1400
rect 4026 1388 4056 1400
rect 4112 1388 4142 1400
tri 3194 1285 3195 1286 se
rect 3195 1285 3201 1337
rect 3253 1285 3267 1337
rect 3319 1285 3325 1337
tri 3181 1272 3194 1285 se
rect 3194 1272 3325 1285
tri 3175 1266 3181 1272 se
rect 3181 1266 3325 1272
tri 3169 1260 3175 1266 se
rect 3175 1260 3325 1266
tri 3161 1252 3169 1260 se
rect 3169 1252 3325 1260
rect 1296 1200 1302 1252
rect 1354 1200 1366 1252
rect 1418 1200 3325 1252
rect 3521 1336 3527 1388
rect 3579 1336 3595 1388
rect 3647 1336 3663 1388
rect 3783 1376 3798 1388
rect 3854 1376 3867 1388
rect 4053 1376 4056 1388
rect 4120 1376 4142 1388
rect 4198 1376 4228 1432
rect 4284 1376 4314 1432
rect 4370 1376 4399 1432
rect 4455 1376 4464 1432
rect 3715 1348 3731 1376
rect 3783 1348 3799 1376
rect 3851 1348 3867 1376
rect 3919 1348 3934 1376
rect 3986 1348 4001 1376
rect 4053 1348 4068 1376
rect 4120 1348 4464 1376
rect 3783 1336 3798 1348
rect 3854 1336 3867 1348
rect 4053 1336 4056 1348
rect 4120 1336 4142 1348
rect 3521 1324 3712 1336
rect 3768 1324 3798 1336
rect 3854 1324 3884 1336
rect 3940 1324 3970 1336
rect 4026 1324 4056 1336
rect 4112 1324 4142 1336
rect 3521 1272 3527 1324
rect 3579 1272 3595 1324
rect 3647 1272 3663 1324
rect 3783 1292 3798 1324
rect 3854 1292 3867 1324
rect 4053 1292 4056 1324
rect 4120 1292 4142 1324
rect 4198 1292 4228 1348
rect 4284 1292 4314 1348
rect 4370 1292 4399 1348
rect 4455 1292 4464 1348
rect 3715 1272 3731 1292
rect 3783 1272 3799 1292
rect 3851 1272 3867 1292
rect 3919 1272 3934 1292
rect 3986 1272 4001 1292
rect 4053 1272 4068 1292
rect 4120 1272 4464 1292
rect 4527 1300 4579 1782
tri 4579 1300 4601 1322 sw
rect 4693 1301 4745 1852
rect 4789 1381 4841 1980
tri 4979 1949 5010 1980 ne
tri 5695 1949 5726 1980 ne
tri 6192 1949 6223 1980 ne
rect 6223 1949 6278 1980
tri 6411 1949 6442 1980 ne
tri 6223 1948 6224 1949 ne
rect 6224 1948 6278 1949
rect 4908 1942 4960 1948
rect 5621 1942 5673 1948
tri 6224 1946 6226 1948 ne
rect 4908 1880 4960 1890
rect 5410 1918 5462 1924
tri 4960 1880 4962 1882 sw
tri 5408 1880 5410 1882 se
rect 4908 1866 4962 1880
tri 4962 1866 4976 1880 sw
tri 5394 1866 5408 1880 se
rect 5408 1866 5410 1880
rect 4908 1858 4976 1866
tri 4976 1858 4984 1866 sw
tri 5386 1858 5394 1866 se
rect 5394 1858 5462 1866
rect 4960 1854 4984 1858
tri 4984 1854 4988 1858 sw
tri 5382 1854 5386 1858 se
rect 5386 1854 5462 1858
rect 4960 1848 4988 1854
tri 4988 1848 4994 1854 sw
tri 5376 1848 5382 1854 se
rect 5382 1848 5410 1854
rect 4960 1806 5410 1848
rect 4908 1802 5410 1806
rect 4908 1796 5462 1802
rect 5621 1858 5673 1890
rect 5794 1880 6140 1932
tri 6054 1858 6076 1880 ne
rect 6076 1858 6140 1880
tri 6076 1846 6088 1858 ne
rect 5621 1512 5673 1806
rect 6088 1586 6140 1858
rect 6226 1694 6278 1948
rect 6340 1942 6392 1948
rect 6340 1880 6392 1890
tri 6392 1880 6398 1886 sw
rect 6678 1880 8538 1932
rect 8590 1880 8602 1932
rect 8654 1880 8660 1932
rect 6340 1858 6398 1880
rect 6392 1852 6398 1858
tri 6398 1852 6426 1880 sw
rect 6392 1846 8740 1852
rect 6392 1806 8688 1846
rect 6340 1800 8688 1806
tri 8654 1794 8660 1800 ne
rect 8660 1794 8688 1800
tri 8660 1782 8672 1794 ne
rect 8672 1782 8740 1794
tri 8672 1766 8688 1782 ne
tri 6278 1694 6283 1699 sw
rect 6473 1694 6479 1746
rect 6531 1694 6580 1746
rect 6632 1694 6681 1746
rect 6733 1694 6782 1746
rect 6834 1694 6882 1746
rect 6934 1694 6982 1746
rect 7034 1711 7082 1746
rect 7065 1694 7082 1711
rect 7134 1711 7182 1746
rect 7234 1711 7282 1746
rect 7134 1694 7137 1711
rect 7234 1694 7265 1711
rect 7334 1694 7382 1746
rect 7434 1711 7482 1746
rect 7534 1711 7582 1746
rect 7449 1694 7482 1711
rect 7577 1694 7582 1711
rect 7634 1711 7682 1746
rect 7734 1711 7782 1746
rect 7634 1694 7649 1711
rect 7734 1694 7776 1711
rect 7834 1694 7841 1746
rect 8688 1724 8740 1730
rect 6226 1677 6283 1694
tri 6226 1672 6231 1677 ne
rect 6231 1672 6283 1677
tri 6283 1672 6305 1694 sw
rect 6473 1672 7009 1694
rect 7065 1672 7137 1694
rect 7193 1672 7265 1694
rect 7321 1672 7393 1694
rect 7449 1672 7521 1694
rect 7577 1672 7649 1694
rect 7705 1672 7776 1694
rect 7832 1672 7841 1694
tri 6231 1660 6243 1672 ne
rect 6243 1660 6305 1672
tri 6305 1660 6317 1672 sw
tri 6243 1625 6278 1660 ne
rect 6278 1625 6317 1660
tri 6278 1620 6283 1625 ne
rect 6283 1620 6317 1625
tri 6317 1620 6357 1660 sw
rect 6473 1620 6479 1672
rect 6531 1620 6580 1672
rect 6632 1620 6681 1672
rect 6733 1620 6782 1672
rect 6834 1620 6882 1672
rect 6934 1620 6982 1672
rect 7065 1655 7082 1672
rect 7034 1620 7082 1655
rect 7134 1655 7137 1672
rect 7234 1655 7265 1672
rect 7134 1620 7182 1655
rect 7234 1620 7282 1655
rect 7334 1620 7382 1672
rect 7449 1655 7482 1672
rect 7577 1655 7582 1672
rect 7434 1620 7482 1655
rect 7534 1620 7582 1655
rect 7634 1655 7649 1672
rect 7734 1655 7776 1672
rect 7634 1620 7682 1655
rect 7734 1620 7782 1655
rect 7834 1620 7841 1672
tri 6283 1599 6304 1620 ne
rect 6304 1599 6357 1620
tri 6140 1586 6153 1599 sw
tri 6304 1586 6317 1599 ne
rect 6317 1586 6357 1599
tri 6357 1586 6391 1620 sw
rect 6473 1619 7841 1620
rect 6088 1580 6153 1586
tri 6153 1580 6159 1586 sw
tri 6317 1580 6323 1586 ne
rect 6323 1580 9050 1586
rect 6088 1577 6159 1580
tri 6088 1534 6131 1577 ne
rect 6131 1534 6159 1577
tri 6159 1534 6205 1580 sw
tri 6323 1534 6369 1580 ne
rect 6369 1534 9050 1580
rect 9102 1534 9114 1586
rect 9166 1534 9172 1586
rect 9492 1576 9544 1582
tri 9486 1534 9492 1540 se
tri 6131 1524 6141 1534 ne
rect 6141 1524 6205 1534
tri 6205 1524 6215 1534 sw
tri 9476 1524 9486 1534 se
rect 9486 1524 9492 1534
tri 6141 1522 6143 1524 ne
rect 6143 1522 6215 1524
tri 6215 1522 6217 1524 sw
tri 9474 1522 9476 1524 se
rect 9476 1522 9544 1524
tri 5673 1512 5683 1522 sw
tri 6143 1512 6153 1522 ne
rect 6153 1512 6217 1522
tri 6217 1512 6227 1522 sw
tri 9464 1512 9474 1522 se
rect 9474 1512 9544 1522
rect 5621 1500 5683 1512
tri 5683 1500 5695 1512 sw
tri 6153 1506 6159 1512 ne
rect 6159 1506 6227 1512
tri 6227 1506 6233 1512 sw
tri 9458 1506 9464 1512 se
rect 9464 1506 9492 1512
tri 6159 1500 6165 1506 ne
rect 6165 1500 9492 1506
tri 5621 1460 5661 1500 ne
rect 5661 1460 5695 1500
tri 5695 1460 5735 1500 sw
tri 6165 1460 6205 1500 ne
rect 6205 1460 9492 1500
tri 5661 1426 5695 1460 ne
rect 5695 1454 5735 1460
tri 5735 1454 5741 1460 sw
tri 6205 1454 6211 1460 ne
rect 6211 1454 9544 1460
rect 5695 1426 5741 1454
tri 5741 1426 5769 1454 sw
tri 5695 1403 5718 1426 ne
rect 5718 1403 8874 1426
tri 4789 1374 4796 1381 ne
rect 4796 1374 4841 1381
tri 4841 1374 4870 1403 sw
tri 5718 1374 5747 1403 ne
rect 5747 1374 8874 1403
rect 8926 1374 8938 1426
rect 8990 1374 8996 1426
rect 9652 1416 9704 1422
tri 4796 1364 4806 1374 ne
rect 4806 1364 4870 1374
tri 4870 1364 4880 1374 sw
tri 4806 1352 4818 1364 ne
rect 4818 1352 4880 1364
tri 4880 1352 4892 1364 sw
tri 4818 1346 4824 1352 ne
rect 4824 1346 4892 1352
tri 4892 1346 4898 1352 sw
tri 9618 1346 9652 1380 se
rect 9652 1352 9704 1364
tri 4824 1329 4841 1346 ne
rect 4841 1329 9652 1346
tri 4841 1323 4847 1329 ne
rect 4847 1323 9652 1329
tri 4693 1300 4694 1301 ne
rect 4694 1300 4745 1301
tri 4745 1300 4768 1323 sw
tri 4847 1300 4870 1323 ne
rect 4870 1300 9652 1323
rect 9970 1336 10022 1342
tri 4527 1284 4543 1300 ne
rect 4543 1284 4601 1300
tri 4601 1284 4617 1300 sw
tri 4694 1284 4710 1300 ne
rect 4710 1294 4768 1300
tri 4768 1294 4774 1300 sw
tri 4870 1294 4876 1300 ne
rect 4876 1294 9704 1300
tri 9964 1294 9970 1300 se
rect 4710 1284 4774 1294
tri 4774 1284 4784 1294 sw
tri 9954 1284 9964 1294 se
rect 9964 1284 9970 1294
tri 4543 1272 4555 1284 ne
rect 4555 1272 4617 1284
tri 4617 1272 4629 1284 sw
tri 4710 1272 4722 1284 ne
rect 4722 1272 4784 1284
tri 4784 1272 4796 1284 sw
tri 9942 1272 9954 1284 se
rect 9954 1272 10022 1284
rect 3521 1264 4464 1272
rect 3521 1260 3712 1264
rect 3768 1260 3798 1264
rect 3854 1260 3884 1264
rect 3940 1260 3970 1264
rect 4026 1260 4056 1264
rect 4112 1260 4142 1264
rect 3521 1208 3527 1260
rect 3579 1208 3595 1260
rect 3647 1208 3663 1260
rect 3783 1208 3798 1260
rect 3854 1208 3867 1260
rect 4053 1208 4056 1260
rect 4120 1208 4142 1260
rect 4198 1208 4228 1264
rect 4284 1208 4314 1264
rect 4370 1208 4399 1264
rect 4455 1208 4464 1264
tri 4555 1260 4567 1272 ne
rect 4567 1266 4629 1272
tri 4629 1266 4635 1272 sw
tri 4722 1266 4728 1272 ne
rect 4728 1266 4796 1272
tri 4796 1266 4802 1272 sw
tri 9936 1266 9942 1272 se
rect 9942 1266 9970 1272
rect 4567 1260 4635 1266
tri 4635 1260 4641 1266 sw
tri 4728 1260 4734 1266 ne
rect 4734 1260 9970 1266
tri 4567 1248 4579 1260 ne
rect 4579 1249 4641 1260
tri 4641 1249 4652 1260 sw
tri 4734 1249 4745 1260 ne
rect 4745 1249 9970 1260
rect 4579 1248 4652 1249
tri 4579 1220 4607 1248 ne
rect 4607 1220 4652 1248
tri 4652 1220 4681 1249 sw
tri 4745 1220 4774 1249 ne
rect 4774 1220 9970 1249
rect 3521 1206 4464 1208
tri 4607 1206 4621 1220 ne
rect 4621 1214 4681 1220
tri 4681 1214 4687 1220 sw
tri 4774 1214 4780 1220 ne
rect 4780 1214 10022 1220
rect 4621 1206 4687 1214
tri 4687 1206 4695 1214 sw
tri 4621 1200 4627 1206 ne
rect 4627 1200 4695 1206
tri 4695 1200 4701 1206 sw
tri 4627 1186 4641 1200 ne
rect 4641 1186 4701 1200
tri 4701 1186 4715 1200 sw
tri 4641 1150 4677 1186 ne
rect 4677 1150 9502 1186
rect 1240 1098 1246 1150
rect 1298 1098 1310 1150
rect 1362 1134 4530 1150
tri 4530 1134 4546 1150 sw
tri 4677 1134 4693 1150 ne
rect 4693 1134 9502 1150
rect 9554 1134 9566 1186
rect 9618 1134 9624 1186
rect 1362 1098 4546 1134
tri 4508 1084 4522 1098 ne
rect 4522 1095 4546 1098
tri 4546 1095 4585 1134 sw
rect 4522 1084 4585 1095
tri 4585 1084 4596 1095 sw
rect 8388 1086 8819 1095
tri 4522 1080 4526 1084 ne
rect 4526 1080 4596 1084
tri 4596 1080 4600 1084 sw
tri 4526 1076 4530 1080 ne
rect 4530 1078 4600 1080
tri 4600 1078 4602 1080 sw
rect 4530 1076 4602 1078
tri 4530 1064 4542 1076 ne
rect 4542 1064 4602 1076
tri 4602 1064 4616 1078 sw
tri 4542 1059 4547 1064 ne
rect 4547 1059 4616 1064
rect 1104 1007 1110 1059
rect 1162 1007 1174 1059
rect 1226 1055 4453 1059
tri 4453 1055 4457 1059 sw
tri 4547 1055 4551 1059 ne
rect 4551 1055 4616 1059
rect 1226 1048 4457 1055
tri 4457 1048 4464 1055 sw
tri 4551 1048 4558 1055 ne
rect 4558 1048 4616 1055
tri 4616 1048 4632 1064 sw
rect 5823 1050 6623 1078
rect 5823 1048 5832 1050
rect 5888 1048 5913 1050
rect 5969 1048 5994 1050
rect 6050 1048 6075 1050
rect 6131 1048 6156 1050
rect 6212 1048 6237 1050
rect 6293 1048 6318 1050
rect 6374 1048 6398 1050
rect 6454 1048 6478 1050
rect 6534 1048 6558 1050
rect 6614 1048 6623 1050
rect 1226 1010 4464 1048
tri 4464 1010 4502 1048 sw
tri 4558 1010 4596 1048 ne
rect 4596 1010 4632 1048
tri 4632 1010 4670 1048 sw
rect 1226 1007 4502 1010
tri 4431 996 4442 1007 ne
rect 4442 996 4502 1007
tri 4502 996 4516 1010 sw
tri 4596 996 4610 1010 ne
rect 4610 996 4670 1010
tri 4670 996 4684 1010 sw
rect 5823 996 5829 1048
rect 5888 996 5896 1048
rect 6149 996 6156 1048
rect 6216 996 6231 1048
rect 6293 996 6298 1048
rect 6551 996 6558 1048
rect 6617 996 6623 1048
tri 4442 981 4457 996 ne
rect 4457 981 4516 996
tri 4516 981 4531 996 sw
tri 4610 981 4625 996 ne
rect 4625 981 4684 996
tri 4457 975 4463 981 ne
rect 4463 975 4531 981
tri 4531 975 4537 981 sw
tri 4625 975 4631 981 ne
rect 4631 975 4684 981
rect 1032 923 1038 975
rect 1090 923 1102 975
rect 1154 970 4401 975
tri 4401 970 4406 975 sw
tri 4463 970 4468 975 ne
rect 4468 970 4537 975
tri 4537 970 4542 975 sw
tri 4631 970 4636 975 ne
rect 4636 970 4684 975
rect 1154 948 4406 970
tri 4406 948 4428 970 sw
tri 4468 948 4490 970 ne
rect 4490 948 4542 970
tri 4542 948 4564 970 sw
tri 4636 948 4658 970 ne
rect 4658 966 4684 970
tri 4684 966 4714 996 sw
rect 5823 994 5832 996
rect 5888 994 5913 996
rect 5969 994 5994 996
rect 6050 994 6075 996
rect 6131 994 6156 996
rect 6212 994 6237 996
rect 6293 994 6318 996
rect 6374 994 6398 996
rect 6454 994 6478 996
rect 6534 994 6558 996
rect 6614 994 6623 996
rect 5823 966 6623 994
rect 8388 1064 8763 1086
rect 8440 1030 8763 1064
rect 8440 1012 8819 1030
rect 8388 1006 8819 1012
rect 8388 1000 8763 1006
rect 4658 948 4714 966
tri 4714 948 4732 966 sw
rect 8440 950 8763 1000
rect 9172 1080 9624 1086
rect 9224 1033 9572 1080
rect 9224 1028 9253 1033
tri 9253 1028 9258 1033 nw
tri 9538 1028 9543 1033 ne
rect 9543 1028 9572 1033
rect 9172 1016 9241 1028
tri 9241 1016 9253 1028 nw
tri 9543 1016 9555 1028 ne
rect 9555 1016 9624 1028
tri 9224 999 9241 1016 nw
tri 9555 999 9572 1016 ne
rect 9172 958 9224 964
rect 9572 958 9624 964
rect 8440 948 8819 950
rect 1154 946 4428 948
tri 4428 946 4430 948 sw
tri 4490 946 4492 948 ne
rect 4492 946 4564 948
tri 4564 946 4566 948 sw
tri 4658 946 4660 948 ne
rect 4660 946 4732 948
tri 4732 946 4734 948 sw
rect 1154 936 4430 946
tri 4430 936 4440 946 sw
tri 4492 936 4502 946 ne
rect 4502 936 4566 946
tri 4566 936 4576 946 sw
tri 4660 936 4670 946 ne
rect 4670 941 4734 946
tri 4734 941 4739 946 sw
rect 8388 941 8819 948
rect 9492 946 9544 952
rect 4670 936 4739 941
tri 4739 936 4744 941 sw
rect 1154 923 4440 936
tri 4379 896 4406 923 ne
rect 4406 919 4440 923
tri 4440 919 4457 936 sw
tri 4502 919 4519 936 ne
rect 4519 919 4576 936
rect 4406 907 4457 919
tri 4457 907 4469 919 sw
tri 4519 907 4531 919 ne
rect 4531 907 4576 919
tri 4576 907 4605 936 sw
tri 4670 907 4699 936 ne
rect 4699 910 4744 936
tri 4744 910 4770 936 sw
rect 4699 907 4770 910
rect 4406 896 4469 907
tri 4469 896 4480 907 sw
tri 4531 896 4542 907 ne
rect 4542 896 4605 907
tri 4605 896 4616 907 sw
tri 4699 896 4710 907 ne
rect 4710 896 4770 907
tri 4406 895 4407 896 ne
rect 4407 895 4480 896
rect 957 843 963 895
rect 1015 843 1027 895
rect 1079 894 4211 895
tri 4211 894 4212 895 sw
tri 4407 894 4408 895 ne
rect 4408 894 4480 895
tri 4480 894 4482 896 sw
tri 4542 894 4544 896 ne
rect 4544 894 4616 896
tri 4616 894 4618 896 sw
tri 4710 894 4712 896 ne
rect 4712 894 4770 896
tri 4770 894 4786 910 sw
rect 1079 882 4212 894
tri 4212 882 4224 894 sw
tri 4408 882 4420 894 ne
rect 4420 882 4482 894
tri 4482 882 4494 894 sw
tri 4544 882 4556 894 ne
rect 4556 882 4618 894
tri 4618 882 4630 894 sw
tri 4712 882 4724 894 ne
rect 4724 882 4786 894
tri 4786 882 4798 894 sw
rect 1079 876 4224 882
tri 4224 876 4230 882 sw
tri 4420 876 4426 882 ne
rect 4426 876 4494 882
tri 4494 876 4500 882 sw
tri 4556 876 4562 882 ne
rect 4562 876 4630 882
tri 4630 876 4636 882 sw
tri 4724 876 4730 882 ne
rect 4730 876 4798 882
tri 4798 876 4804 882 sw
tri 9458 876 9492 910 se
rect 9492 882 9544 894
rect 1079 843 4230 876
tri 4230 843 4263 876 sw
tri 4426 843 4459 876 ne
rect 4459 862 4500 876
tri 4500 862 4514 876 sw
tri 4562 862 4576 876 ne
rect 4576 862 4636 876
tri 4636 862 4650 876 sw
tri 4730 862 4744 876 ne
rect 4744 862 4804 876
tri 4804 862 4818 876 sw
rect 4459 845 4514 862
tri 4514 845 4531 862 sw
tri 4576 845 4593 862 ne
rect 4593 845 4650 862
rect 4459 843 4531 845
tri 4189 824 4208 843 ne
rect 4208 824 4263 843
tri 4263 824 4282 843 sw
tri 4459 824 4478 843 ne
rect 4478 833 4531 843
tri 4531 833 4543 845 sw
tri 4593 833 4605 845 ne
rect 4605 833 4650 845
tri 4650 833 4679 862 sw
tri 4744 833 4773 862 ne
rect 4773 833 4818 862
rect 4478 824 4543 833
tri 4543 824 4552 833 sw
tri 4605 824 4614 833 ne
rect 4614 824 4679 833
tri 4679 824 4688 833 sw
tri 4773 824 4782 833 ne
rect 4782 824 4818 833
tri 4818 824 4856 862 sw
rect 8788 824 8794 876
rect 8846 824 8858 876
rect 8910 830 9492 876
rect 8910 824 9544 830
tri 4208 822 4210 824 ne
rect 4210 822 4282 824
tri 4282 822 4284 824 sw
tri 4478 822 4480 824 ne
rect 4480 822 4552 824
tri 4552 822 4554 824 sw
tri 4614 822 4616 824 ne
rect 4616 822 4688 824
tri 4688 822 4690 824 sw
tri 4782 822 4784 824 ne
rect 4784 822 4856 824
tri 4210 781 4251 822 ne
rect 4251 790 4284 822
tri 4284 790 4316 822 sw
rect 4251 781 4316 790
tri 4480 781 4521 822 ne
rect 4521 788 4554 822
tri 4554 788 4588 822 sw
tri 4616 788 4650 822 ne
rect 4650 788 4690 822
tri 4690 788 4724 822 sw
tri 4784 788 4818 822 ne
rect 4818 788 4856 822
tri 4856 788 4892 824 sw
rect 4521 781 4588 788
tri 4588 781 4595 788 sw
tri 4650 781 4657 788 ne
rect 4657 781 4724 788
tri 4724 781 4731 788 sw
tri 4818 781 4825 788 ne
rect 4825 787 4892 788
tri 4892 787 4893 788 sw
rect 4825 781 4893 787
tri 4893 781 4899 787 sw
rect 9332 781 9384 787
tri 4251 769 4263 781 ne
rect 4263 769 4316 781
tri 4263 768 4264 769 ne
rect 827 659 833 711
rect 885 659 897 711
rect 949 708 3732 711
rect 949 659 3610 708
tri 3601 656 3604 659 ne
rect 3604 656 3610 659
rect 3662 656 3674 708
rect 3726 656 3732 708
rect 4264 701 4316 769
tri 4521 748 4554 781 ne
rect 4554 771 4595 781
tri 4595 771 4605 781 sw
tri 4657 771 4667 781 ne
rect 4667 771 4731 781
rect 4554 759 4605 771
tri 4605 759 4617 771 sw
tri 4667 759 4679 771 ne
rect 4679 759 4731 771
tri 4731 759 4753 781 sw
tri 4825 759 4847 781 ne
rect 4847 759 4899 781
rect 4554 748 4617 759
tri 4617 748 4628 759 sw
tri 4554 729 4573 748 ne
rect 4573 729 4628 748
tri 4679 729 4709 759 ne
rect 4709 729 4753 759
tri 4753 729 4783 759 sw
tri 4847 729 4877 759 ne
rect 4877 745 4899 759
tri 4899 745 4935 781 sw
rect 4877 729 4935 745
tri 4935 729 4951 745 sw
tri 9316 729 9332 745 se
tri 4573 726 4576 729 ne
rect 4264 637 4316 649
rect 904 556 910 608
rect 962 556 974 608
rect 1026 556 3712 608
rect 3764 556 3776 608
rect 3828 556 3834 608
rect 4264 579 4316 585
rect 4576 701 4628 729
tri 4709 717 4721 729 ne
rect 4721 717 4783 729
tri 4783 717 4795 729 sw
tri 4877 717 4889 729 ne
rect 4889 717 4951 729
tri 4951 717 4963 729 sw
tri 9304 717 9316 729 se
rect 9316 717 9384 729
tri 4721 714 4724 717 ne
rect 4724 714 4795 717
tri 4795 714 4798 717 sw
tri 4889 714 4892 717 ne
rect 4892 714 4963 717
tri 4963 714 4966 717 sw
tri 9301 714 9304 717 se
rect 9304 714 9332 717
tri 4724 685 4753 714 ne
rect 4753 711 4798 714
tri 4798 711 4801 714 sw
tri 4892 711 4895 714 ne
rect 4895 711 5018 714
rect 4753 685 4801 711
tri 4801 685 4827 711 sw
tri 4895 685 4921 711 ne
rect 4921 685 5018 711
tri 4753 662 4776 685 ne
rect 4776 662 4827 685
tri 4827 662 4850 685 sw
tri 4921 662 4944 685 ne
rect 4944 662 5018 685
rect 5070 662 5082 714
rect 5134 662 5140 714
tri 9298 711 9301 714 se
rect 9301 711 9332 714
tri 4776 659 4779 662 ne
rect 4779 659 4850 662
tri 4850 659 4853 662 sw
rect 5976 659 5982 711
rect 6034 659 6046 711
rect 6098 665 9332 711
rect 6098 659 9384 665
rect 9412 678 9464 684
rect 4576 626 4628 649
tri 4779 626 4812 659 ne
rect 4812 642 4853 659
tri 4853 642 4870 659 sw
rect 4812 626 4870 642
tri 4870 626 4886 642 sw
tri 9396 626 9412 642 se
tri 4812 614 4824 626 ne
rect 4824 614 4886 626
tri 4886 614 4898 626 sw
tri 9384 614 9396 626 se
rect 9396 614 9464 626
tri 4824 611 4827 614 ne
rect 4827 611 4898 614
tri 4898 611 4901 614 sw
tri 9381 611 9384 614 se
rect 9384 611 9412 614
tri 4827 608 4830 611 ne
rect 4830 608 5022 611
rect 4576 568 4628 574
tri 4830 568 4870 608 ne
rect 4870 568 5022 608
tri 4870 559 4879 568 ne
rect 4879 559 5022 568
rect 5074 559 5086 611
rect 5138 559 5144 611
tri 9378 608 9381 611 se
rect 9381 608 9412 611
rect 5874 556 5880 608
rect 5932 556 5944 608
rect 5996 562 9412 608
rect 9890 598 9942 604
rect 5996 556 9464 562
tri 9884 556 9890 562 se
tri 9874 546 9884 556 se
rect 9884 546 9890 556
tri 9862 534 9874 546 se
rect 9874 534 9942 546
tri 9856 528 9862 534 se
rect 9862 528 9890 534
rect 697 476 703 528
rect 755 476 767 528
rect 819 476 3232 528
rect 3284 476 3296 528
rect 3348 476 3354 528
rect 6354 476 6360 528
rect 6412 476 6424 528
rect 6476 482 9890 528
rect 6476 476 9942 482
rect 540 423 592 429
rect 627 392 633 444
rect 685 392 697 444
rect 749 392 2923 444
rect 2975 392 2987 444
rect 3039 392 3045 444
rect 6663 392 6669 444
rect 6721 392 6733 444
rect 6785 392 9258 444
rect 9310 392 9322 444
rect 9374 392 9380 444
rect 540 359 592 371
tri 592 356 623 387 sw
rect 592 353 623 356
tri 623 353 626 356 sw
tri 3108 353 3111 356 se
rect 3111 353 4297 356
rect 592 307 2987 353
rect 540 301 2987 307
rect 3039 301 3053 353
rect 3105 304 4297 353
rect 4349 304 4363 356
rect 4415 353 6727 356
rect 4415 304 6603 353
rect 3105 301 3111 304
tri 3111 301 3114 304 nw
tri 6594 301 6597 304 ne
rect 6597 301 6603 304
rect 6655 301 6669 353
rect 6721 301 6727 353
rect 2483 158 2561 164
rect 2483 145 2496 158
rect 2548 145 2561 158
rect 282 122 334 128
rect 282 58 334 70
rect 282 0 334 6
rect 1415 122 1467 128
rect 1415 58 1467 70
rect 1415 0 1467 6
rect 1652 122 1704 128
rect 1652 58 1704 70
rect 1652 0 1704 6
rect 1909 122 1961 128
rect 1909 58 1961 70
rect 1909 0 1961 6
rect 2163 122 2215 128
rect 2163 58 2215 70
rect 2163 0 2215 6
rect 2483 89 2494 145
rect 2550 89 2561 145
rect 2483 65 2561 89
rect 2483 9 2494 65
rect 2550 9 2561 65
rect 2483 6 2496 9
rect 2548 6 2561 9
rect 2483 0 2561 6
rect 6840 145 6896 154
rect 8467 145 8523 154
rect 6840 70 6843 89
rect 6895 70 6896 89
rect 6840 65 6896 70
rect 6840 6 6843 9
rect 6895 6 6896 9
rect 6840 0 6896 6
rect 8176 122 8228 128
rect 8176 58 8228 70
rect 8176 0 8228 6
rect 8467 70 8469 89
rect 8521 70 8523 89
rect 8467 65 8523 70
rect 8467 6 8469 9
rect 8521 6 8523 9
rect 8467 0 8523 6
rect 8700 145 8756 154
rect 8700 70 8701 89
rect 8753 70 8756 89
rect 8700 65 8756 70
rect 8700 6 8701 9
rect 8753 6 8756 9
rect 8700 0 8756 6
rect 8916 145 8972 154
rect 10029 145 10085 154
rect 8916 70 8918 89
rect 8970 70 8972 89
rect 8916 65 8972 70
rect 8916 6 8918 9
rect 8970 6 8972 9
rect 8916 0 8972 6
rect 9232 122 9284 128
rect 9232 58 9284 70
rect 9232 0 9284 6
rect 9572 122 9624 128
rect 9572 58 9624 70
rect 9572 0 9624 6
rect 9784 122 9836 128
rect 9784 58 9836 70
rect 9784 0 9836 6
rect 10029 70 10031 89
rect 10083 70 10085 89
rect 10029 65 10085 70
rect 10029 6 10031 9
rect 10083 6 10085 9
rect 10029 0 10085 6
rect 10261 145 10317 154
rect 10261 70 10263 89
rect 10315 70 10317 89
rect 10261 65 10317 70
rect 10261 6 10263 9
rect 10315 6 10317 9
rect 10261 0 10317 6
<< via2 >>
rect 291 38890 347 38946
rect 374 38890 430 38946
rect 456 38890 512 38946
rect 538 38890 594 38946
rect 620 38890 676 38946
rect 702 38890 758 38946
rect 784 38890 840 38946
rect 866 38890 922 38946
rect 948 38890 1004 38946
rect 1030 38890 1086 38946
rect 1112 38890 1168 38946
rect 1194 38890 1250 38946
rect 1276 38890 1332 38946
rect 1358 38890 1414 38946
rect 2714 38923 2770 38979
rect 2794 38923 2850 38979
rect 2874 38923 2930 38979
rect 2954 38923 3010 38979
rect 3034 38923 3090 38979
rect 3114 38923 3170 38979
rect 3194 38923 3250 38979
rect 3274 38923 3330 38979
rect 3354 38923 3410 38979
rect 3434 38923 3490 38979
rect 291 38804 347 38860
rect 374 38804 430 38860
rect 456 38804 512 38860
rect 538 38804 594 38860
rect 620 38804 676 38860
rect 702 38804 758 38860
rect 784 38804 840 38860
rect 866 38804 922 38860
rect 948 38804 1004 38860
rect 1030 38804 1086 38860
rect 1112 38804 1168 38860
rect 1194 38804 1250 38860
rect 1276 38804 1332 38860
rect 1358 38804 1414 38860
rect 2714 38839 2770 38895
rect 2794 38839 2850 38895
rect 2874 38839 2930 38895
rect 2954 38839 3010 38895
rect 3034 38839 3090 38895
rect 3114 38839 3170 38895
rect 3194 38839 3250 38895
rect 3274 38839 3330 38895
rect 3354 38839 3410 38895
rect 3434 38839 3490 38895
rect 291 38718 347 38774
rect 374 38718 430 38774
rect 456 38718 512 38774
rect 538 38718 594 38774
rect 620 38718 676 38774
rect 702 38718 758 38774
rect 784 38718 840 38774
rect 866 38718 922 38774
rect 948 38718 1004 38774
rect 1030 38718 1086 38774
rect 1112 38718 1168 38774
rect 1194 38718 1250 38774
rect 1276 38718 1332 38774
rect 1358 38718 1414 38774
rect 2714 38755 2770 38811
rect 2794 38755 2850 38811
rect 2874 38755 2930 38811
rect 2954 38755 3010 38811
rect 3034 38755 3090 38811
rect 3114 38755 3170 38811
rect 3194 38755 3250 38811
rect 3274 38755 3330 38811
rect 3354 38755 3410 38811
rect 3434 38755 3490 38811
rect 291 38632 347 38688
rect 374 38632 430 38688
rect 456 38632 512 38688
rect 538 38632 594 38688
rect 620 38632 676 38688
rect 702 38632 758 38688
rect 784 38632 840 38688
rect 866 38632 922 38688
rect 948 38632 1004 38688
rect 1030 38632 1086 38688
rect 1112 38632 1168 38688
rect 1194 38632 1250 38688
rect 1276 38632 1332 38688
rect 1358 38632 1414 38688
rect 2714 38671 2770 38727
rect 2794 38671 2850 38727
rect 2874 38671 2930 38727
rect 2954 38671 3010 38727
rect 3034 38671 3090 38727
rect 3114 38671 3170 38727
rect 3194 38671 3250 38727
rect 3274 38671 3330 38727
rect 3354 38671 3410 38727
rect 3434 38671 3490 38727
rect 291 38546 347 38602
rect 374 38546 430 38602
rect 456 38546 512 38602
rect 538 38546 594 38602
rect 620 38546 676 38602
rect 702 38546 758 38602
rect 784 38546 840 38602
rect 866 38546 922 38602
rect 948 38546 1004 38602
rect 1030 38546 1086 38602
rect 1112 38546 1168 38602
rect 1194 38546 1250 38602
rect 1276 38546 1332 38602
rect 1358 38546 1414 38602
rect 2714 38587 2770 38643
rect 2794 38587 2850 38643
rect 2874 38587 2930 38643
rect 2954 38587 3010 38643
rect 3034 38587 3090 38643
rect 3114 38587 3170 38643
rect 3194 38587 3250 38643
rect 3274 38587 3330 38643
rect 3354 38587 3410 38643
rect 3434 38587 3490 38643
rect 291 38460 347 38516
rect 374 38460 430 38516
rect 456 38460 512 38516
rect 538 38460 594 38516
rect 620 38460 676 38516
rect 702 38460 758 38516
rect 784 38460 840 38516
rect 866 38460 922 38516
rect 948 38460 1004 38516
rect 1030 38460 1086 38516
rect 1112 38460 1168 38516
rect 1194 38460 1250 38516
rect 1276 38460 1332 38516
rect 1358 38460 1414 38516
rect 2714 38503 2770 38559
rect 2794 38503 2850 38559
rect 2874 38503 2930 38559
rect 2954 38503 3010 38559
rect 3034 38503 3090 38559
rect 3114 38503 3170 38559
rect 3194 38503 3250 38559
rect 3274 38503 3330 38559
rect 3354 38503 3410 38559
rect 3434 38503 3490 38559
rect 291 38374 347 38430
rect 374 38374 430 38430
rect 456 38374 512 38430
rect 538 38374 594 38430
rect 620 38374 676 38430
rect 702 38374 758 38430
rect 784 38374 840 38430
rect 866 38374 922 38430
rect 948 38374 1004 38430
rect 1030 38374 1086 38430
rect 1112 38374 1168 38430
rect 1194 38374 1250 38430
rect 1276 38374 1332 38430
rect 1358 38374 1414 38430
rect 2714 38419 2770 38475
rect 2794 38419 2850 38475
rect 2874 38419 2930 38475
rect 2954 38419 3010 38475
rect 3034 38419 3090 38475
rect 3114 38419 3170 38475
rect 3194 38419 3250 38475
rect 3274 38419 3330 38475
rect 3354 38419 3410 38475
rect 3434 38419 3490 38475
rect 291 38288 347 38344
rect 374 38288 430 38344
rect 456 38288 512 38344
rect 538 38288 594 38344
rect 620 38288 676 38344
rect 702 38288 758 38344
rect 784 38288 840 38344
rect 866 38288 922 38344
rect 948 38288 1004 38344
rect 1030 38288 1086 38344
rect 1112 38288 1168 38344
rect 1194 38288 1250 38344
rect 1276 38288 1332 38344
rect 1358 38288 1414 38344
rect 2714 38335 2770 38391
rect 2794 38335 2850 38391
rect 2874 38335 2930 38391
rect 2954 38335 3010 38391
rect 3034 38335 3090 38391
rect 3114 38335 3170 38391
rect 3194 38335 3250 38391
rect 3274 38335 3330 38391
rect 3354 38335 3410 38391
rect 3434 38335 3490 38391
rect 291 38202 347 38258
rect 374 38202 430 38258
rect 456 38202 512 38258
rect 538 38202 594 38258
rect 620 38202 676 38258
rect 702 38202 758 38258
rect 784 38202 840 38258
rect 866 38202 922 38258
rect 948 38202 1004 38258
rect 1030 38202 1086 38258
rect 1112 38202 1168 38258
rect 1194 38202 1250 38258
rect 1276 38202 1332 38258
rect 1358 38202 1414 38258
rect 2714 38251 2770 38307
rect 2794 38251 2850 38307
rect 2874 38251 2930 38307
rect 2954 38251 3010 38307
rect 3034 38251 3090 38307
rect 3114 38251 3170 38307
rect 3194 38251 3250 38307
rect 3274 38251 3330 38307
rect 3354 38251 3410 38307
rect 3434 38251 3490 38307
rect 291 38116 347 38172
rect 374 38116 430 38172
rect 456 38116 512 38172
rect 538 38116 594 38172
rect 620 38116 676 38172
rect 702 38116 758 38172
rect 784 38116 840 38172
rect 866 38116 922 38172
rect 948 38116 1004 38172
rect 1030 38116 1086 38172
rect 1112 38116 1168 38172
rect 1194 38116 1250 38172
rect 1276 38116 1332 38172
rect 1358 38116 1414 38172
rect 2714 38167 2770 38223
rect 2794 38167 2850 38223
rect 2874 38167 2930 38223
rect 2954 38167 3010 38223
rect 3034 38167 3090 38223
rect 3114 38167 3170 38223
rect 3194 38167 3250 38223
rect 3274 38167 3330 38223
rect 3354 38167 3410 38223
rect 3434 38167 3490 38223
rect 291 38030 347 38086
rect 374 38030 430 38086
rect 456 38030 512 38086
rect 538 38030 594 38086
rect 620 38030 676 38086
rect 702 38030 758 38086
rect 784 38030 840 38086
rect 866 38030 922 38086
rect 948 38030 1004 38086
rect 1030 38030 1086 38086
rect 1112 38030 1168 38086
rect 1194 38030 1250 38086
rect 1276 38030 1332 38086
rect 1358 38030 1414 38086
rect 2714 38082 2770 38138
rect 2794 38082 2850 38138
rect 2874 38082 2930 38138
rect 2954 38082 3010 38138
rect 3034 38082 3090 38138
rect 3114 38082 3170 38138
rect 3194 38082 3250 38138
rect 3274 38082 3330 38138
rect 3354 38082 3410 38138
rect 3434 38082 3490 38138
rect 2714 37997 2770 38053
rect 2794 37997 2850 38053
rect 2874 37997 2930 38053
rect 2954 37997 3010 38053
rect 3034 37997 3090 38053
rect 3114 37997 3170 38053
rect 3194 37997 3250 38053
rect 3274 37997 3330 38053
rect 3354 37997 3410 38053
rect 3434 37997 3490 38053
rect 8035 36274 8091 36330
rect 8116 36274 8172 36330
rect 8197 36274 8253 36330
rect 8277 36274 8333 36330
rect 8357 36274 8413 36330
rect 8437 36274 8493 36330
rect 8517 36274 8573 36330
rect 8597 36274 8653 36330
rect 8677 36274 8733 36330
rect 8757 36274 8813 36330
rect 8837 36274 8893 36330
rect 8917 36274 8973 36330
rect 8997 36274 9053 36330
rect 9077 36274 9133 36330
rect 9157 36274 9213 36330
rect 9237 36274 9293 36330
rect 9317 36274 9373 36330
rect 9397 36274 9453 36330
rect 9477 36274 9533 36330
rect 9557 36274 9613 36330
rect 9637 36274 9693 36330
rect 9717 36274 9773 36330
rect 9797 36274 9853 36330
rect 9877 36274 9933 36330
rect 9957 36274 10013 36330
rect 8035 36188 8091 36244
rect 8116 36188 8172 36244
rect 8197 36188 8253 36244
rect 8277 36188 8333 36244
rect 8357 36188 8413 36244
rect 8437 36188 8493 36244
rect 8517 36188 8573 36244
rect 8597 36188 8653 36244
rect 8677 36188 8733 36244
rect 8757 36188 8813 36244
rect 8837 36188 8893 36244
rect 8917 36188 8973 36244
rect 8997 36188 9053 36244
rect 9077 36188 9133 36244
rect 9157 36188 9213 36244
rect 9237 36188 9293 36244
rect 9317 36188 9373 36244
rect 9397 36188 9453 36244
rect 9477 36188 9533 36244
rect 9557 36188 9613 36244
rect 9637 36188 9693 36244
rect 9717 36188 9773 36244
rect 9797 36188 9853 36244
rect 9877 36188 9933 36244
rect 9957 36188 10013 36244
rect 8035 36102 8091 36158
rect 8116 36102 8172 36158
rect 8197 36102 8253 36158
rect 8277 36102 8333 36158
rect 8357 36102 8413 36158
rect 8437 36102 8493 36158
rect 8517 36102 8573 36158
rect 8597 36102 8653 36158
rect 8677 36102 8733 36158
rect 8757 36102 8813 36158
rect 8837 36102 8893 36158
rect 8917 36102 8973 36158
rect 8997 36102 9053 36158
rect 9077 36102 9133 36158
rect 9157 36102 9213 36158
rect 9237 36102 9293 36158
rect 9317 36102 9373 36158
rect 9397 36102 9453 36158
rect 9477 36102 9533 36158
rect 9557 36102 9613 36158
rect 9637 36102 9693 36158
rect 9717 36102 9773 36158
rect 9797 36102 9853 36158
rect 9877 36102 9933 36158
rect 9957 36102 10013 36158
rect 8035 36016 8091 36072
rect 8116 36016 8172 36072
rect 8197 36016 8253 36072
rect 8277 36016 8333 36072
rect 8357 36016 8413 36072
rect 8437 36016 8493 36072
rect 8517 36016 8573 36072
rect 8597 36016 8653 36072
rect 8677 36016 8733 36072
rect 8757 36016 8813 36072
rect 8837 36016 8893 36072
rect 8917 36016 8973 36072
rect 8997 36016 9053 36072
rect 9077 36016 9133 36072
rect 9157 36016 9213 36072
rect 9237 36016 9293 36072
rect 9317 36016 9373 36072
rect 9397 36016 9453 36072
rect 9477 36016 9533 36072
rect 9557 36016 9613 36072
rect 9637 36016 9693 36072
rect 9717 36016 9773 36072
rect 9797 36016 9853 36072
rect 9877 36016 9933 36072
rect 9957 36016 10013 36072
rect 8035 35930 8091 35986
rect 8116 35930 8172 35986
rect 8197 35930 8253 35986
rect 8277 35930 8333 35986
rect 8357 35930 8413 35986
rect 8437 35930 8493 35986
rect 8517 35930 8573 35986
rect 8597 35930 8653 35986
rect 8677 35930 8733 35986
rect 8757 35930 8813 35986
rect 8837 35930 8893 35986
rect 8917 35930 8973 35986
rect 8997 35930 9053 35986
rect 9077 35930 9133 35986
rect 9157 35930 9213 35986
rect 9237 35930 9293 35986
rect 9317 35930 9373 35986
rect 9397 35930 9453 35986
rect 9477 35930 9533 35986
rect 9557 35930 9613 35986
rect 9637 35930 9693 35986
rect 9717 35930 9773 35986
rect 9797 35930 9853 35986
rect 9877 35930 9933 35986
rect 9957 35930 10013 35986
rect 8035 35844 8091 35900
rect 8116 35844 8172 35900
rect 8197 35844 8253 35900
rect 8277 35844 8333 35900
rect 8357 35844 8413 35900
rect 8437 35844 8493 35900
rect 8517 35844 8573 35900
rect 8597 35844 8653 35900
rect 8677 35844 8733 35900
rect 8757 35844 8813 35900
rect 8837 35844 8893 35900
rect 8917 35844 8973 35900
rect 8997 35844 9053 35900
rect 9077 35844 9133 35900
rect 9157 35844 9213 35900
rect 9237 35844 9293 35900
rect 9317 35844 9373 35900
rect 9397 35844 9453 35900
rect 9477 35844 9533 35900
rect 9557 35844 9613 35900
rect 9637 35844 9693 35900
rect 9717 35844 9773 35900
rect 9797 35844 9853 35900
rect 9877 35844 9933 35900
rect 9957 35844 10013 35900
rect 8035 35758 8091 35814
rect 8116 35758 8172 35814
rect 8197 35758 8253 35814
rect 8277 35758 8333 35814
rect 8357 35758 8413 35814
rect 8437 35758 8493 35814
rect 8517 35758 8573 35814
rect 8597 35758 8653 35814
rect 8677 35758 8733 35814
rect 8757 35758 8813 35814
rect 8837 35758 8893 35814
rect 8917 35758 8973 35814
rect 8997 35758 9053 35814
rect 9077 35758 9133 35814
rect 9157 35758 9213 35814
rect 9237 35758 9293 35814
rect 9317 35758 9373 35814
rect 9397 35758 9453 35814
rect 9477 35758 9533 35814
rect 9557 35758 9613 35814
rect 9637 35758 9693 35814
rect 9717 35758 9773 35814
rect 9797 35758 9853 35814
rect 9877 35758 9933 35814
rect 9957 35758 10013 35814
rect 8035 35672 8091 35728
rect 8116 35672 8172 35728
rect 8197 35672 8253 35728
rect 8277 35672 8333 35728
rect 8357 35672 8413 35728
rect 8437 35672 8493 35728
rect 8517 35672 8573 35728
rect 8597 35672 8653 35728
rect 8677 35672 8733 35728
rect 8757 35672 8813 35728
rect 8837 35672 8893 35728
rect 8917 35672 8973 35728
rect 8997 35672 9053 35728
rect 9077 35672 9133 35728
rect 9157 35672 9213 35728
rect 9237 35672 9293 35728
rect 9317 35672 9373 35728
rect 9397 35672 9453 35728
rect 9477 35672 9533 35728
rect 9557 35672 9613 35728
rect 9637 35672 9693 35728
rect 9717 35672 9773 35728
rect 9797 35672 9853 35728
rect 9877 35672 9933 35728
rect 9957 35672 10013 35728
rect 8035 35586 8091 35642
rect 8116 35586 8172 35642
rect 8197 35586 8253 35642
rect 8277 35586 8333 35642
rect 8357 35586 8413 35642
rect 8437 35586 8493 35642
rect 8517 35586 8573 35642
rect 8597 35586 8653 35642
rect 8677 35586 8733 35642
rect 8757 35586 8813 35642
rect 8837 35586 8893 35642
rect 8917 35586 8973 35642
rect 8997 35586 9053 35642
rect 9077 35586 9133 35642
rect 9157 35586 9213 35642
rect 9237 35586 9293 35642
rect 9317 35586 9373 35642
rect 9397 35586 9453 35642
rect 9477 35586 9533 35642
rect 9557 35586 9613 35642
rect 9637 35586 9693 35642
rect 9717 35586 9773 35642
rect 9797 35586 9853 35642
rect 9877 35586 9933 35642
rect 9957 35586 10013 35642
rect 8035 35500 8091 35556
rect 8116 35500 8172 35556
rect 8197 35500 8253 35556
rect 8277 35500 8333 35556
rect 8357 35500 8413 35556
rect 8437 35500 8493 35556
rect 8517 35500 8573 35556
rect 8597 35500 8653 35556
rect 8677 35500 8733 35556
rect 8757 35500 8813 35556
rect 8837 35500 8893 35556
rect 8917 35500 8973 35556
rect 8997 35500 9053 35556
rect 9077 35500 9133 35556
rect 9157 35500 9213 35556
rect 9237 35500 9293 35556
rect 9317 35500 9373 35556
rect 9397 35500 9453 35556
rect 9477 35500 9533 35556
rect 9557 35500 9613 35556
rect 9637 35500 9693 35556
rect 9717 35500 9773 35556
rect 9797 35500 9853 35556
rect 9877 35500 9933 35556
rect 9957 35500 10013 35556
rect 8035 35414 8091 35470
rect 8116 35414 8172 35470
rect 8197 35414 8253 35470
rect 8277 35414 8333 35470
rect 8357 35414 8413 35470
rect 8437 35414 8493 35470
rect 8517 35414 8573 35470
rect 8597 35414 8653 35470
rect 8677 35414 8733 35470
rect 8757 35414 8813 35470
rect 8837 35414 8893 35470
rect 8917 35414 8973 35470
rect 8997 35414 9053 35470
rect 9077 35414 9133 35470
rect 9157 35414 9213 35470
rect 9237 35414 9293 35470
rect 9317 35414 9373 35470
rect 9397 35414 9453 35470
rect 9477 35414 9533 35470
rect 9557 35414 9613 35470
rect 9637 35414 9693 35470
rect 9717 35414 9773 35470
rect 9797 35414 9853 35470
rect 9877 35414 9933 35470
rect 9957 35414 10013 35470
rect 8490 30336 8546 30338
rect 8570 30336 8626 30338
rect 8490 30284 8540 30336
rect 8540 30284 8546 30336
rect 8570 30284 8604 30336
rect 8604 30284 8626 30336
rect 8490 30282 8546 30284
rect 8570 30282 8626 30284
rect 8490 29460 8546 29462
rect 8570 29460 8626 29462
rect 8490 29408 8540 29460
rect 8540 29408 8546 29460
rect 8570 29408 8604 29460
rect 8604 29408 8626 29460
rect 8490 29406 8546 29408
rect 8570 29406 8626 29408
rect 8035 28871 8091 28927
rect 8116 28871 8172 28927
rect 8197 28871 8253 28927
rect 8277 28871 8333 28927
rect 8357 28871 8413 28927
rect 8437 28871 8493 28927
rect 8517 28871 8573 28927
rect 8597 28871 8653 28927
rect 8677 28871 8733 28927
rect 8757 28871 8813 28927
rect 8837 28871 8893 28927
rect 8917 28871 8973 28927
rect 8997 28871 9053 28927
rect 9077 28871 9133 28927
rect 9157 28871 9213 28927
rect 9237 28871 9293 28927
rect 9317 28871 9373 28927
rect 9397 28871 9453 28927
rect 9477 28871 9533 28927
rect 9557 28871 9613 28927
rect 9637 28871 9693 28927
rect 9717 28871 9773 28927
rect 9797 28871 9853 28927
rect 9877 28871 9933 28927
rect 9957 28871 10013 28927
rect 8035 28759 8091 28815
rect 8116 28759 8172 28815
rect 8197 28759 8253 28815
rect 8277 28759 8333 28815
rect 8357 28759 8413 28815
rect 8437 28759 8493 28815
rect 8517 28759 8573 28815
rect 8597 28759 8653 28815
rect 8677 28759 8733 28815
rect 8757 28759 8813 28815
rect 8837 28759 8893 28815
rect 8917 28759 8973 28815
rect 8997 28759 9053 28815
rect 9077 28759 9133 28815
rect 9157 28759 9213 28815
rect 9237 28759 9293 28815
rect 9317 28759 9373 28815
rect 9397 28759 9453 28815
rect 9477 28759 9533 28815
rect 9557 28759 9613 28815
rect 9637 28759 9693 28815
rect 9717 28759 9773 28815
rect 9797 28759 9853 28815
rect 9877 28759 9933 28815
rect 9957 28759 10013 28815
rect 8035 28647 8091 28703
rect 8116 28647 8172 28703
rect 8197 28647 8253 28703
rect 8277 28647 8333 28703
rect 8357 28647 8413 28703
rect 8437 28647 8493 28703
rect 8517 28647 8573 28703
rect 8597 28647 8653 28703
rect 8677 28647 8733 28703
rect 8757 28647 8813 28703
rect 8837 28647 8893 28703
rect 8917 28647 8973 28703
rect 8997 28647 9053 28703
rect 9077 28647 9133 28703
rect 9157 28647 9213 28703
rect 9237 28647 9293 28703
rect 9317 28647 9373 28703
rect 9397 28647 9453 28703
rect 9477 28647 9533 28703
rect 9557 28647 9613 28703
rect 9637 28647 9693 28703
rect 9717 28647 9773 28703
rect 9797 28647 9853 28703
rect 9877 28647 9933 28703
rect 9957 28647 10013 28703
rect 2670 27936 2726 27992
rect 2759 27936 2815 27992
rect 2848 27936 2904 27992
rect 2937 27936 2993 27992
rect 3025 27936 3081 27992
rect 3113 27936 3169 27992
rect 3201 27936 3257 27992
rect 3289 27936 3345 27992
rect 3377 27936 3433 27992
rect 2670 27846 2726 27902
rect 2759 27846 2815 27902
rect 2848 27860 2878 27902
rect 2878 27860 2904 27902
rect 2848 27846 2904 27860
rect 2937 27846 2993 27902
rect 3025 27860 3060 27902
rect 3060 27860 3081 27902
rect 3025 27846 3081 27860
rect 3113 27860 3138 27902
rect 3138 27860 3169 27902
rect 3113 27846 3169 27860
rect 3201 27846 3257 27902
rect 3289 27860 3320 27902
rect 3320 27860 3345 27902
rect 3289 27846 3345 27860
rect 3377 27860 3398 27902
rect 3398 27860 3433 27902
rect 3377 27846 3433 27860
rect 2670 27756 2726 27812
rect 2759 27756 2815 27812
rect 2848 27780 2878 27812
rect 2878 27780 2904 27812
rect 2848 27756 2904 27780
rect 2937 27756 2993 27812
rect 3025 27780 3060 27812
rect 3060 27780 3081 27812
rect 3025 27756 3081 27780
rect 3113 27780 3138 27812
rect 3138 27780 3169 27812
rect 3113 27756 3169 27780
rect 3201 27756 3257 27812
rect 3289 27780 3320 27812
rect 3320 27780 3345 27812
rect 3289 27756 3345 27780
rect 3377 27780 3398 27812
rect 3398 27780 3433 27812
rect 3377 27756 3433 27780
rect 2670 27666 2726 27722
rect 2759 27666 2815 27722
rect 2848 27700 2878 27722
rect 2878 27700 2904 27722
rect 2848 27672 2904 27700
rect 2848 27666 2878 27672
rect 2878 27666 2904 27672
rect 2937 27666 2993 27722
rect 3025 27700 3060 27722
rect 3060 27700 3081 27722
rect 3025 27672 3081 27700
rect 3025 27666 3060 27672
rect 3060 27666 3081 27672
rect 3113 27700 3138 27722
rect 3138 27700 3169 27722
rect 3113 27672 3169 27700
rect 3113 27666 3138 27672
rect 3138 27666 3169 27672
rect 3201 27666 3257 27722
rect 3289 27700 3320 27722
rect 3320 27700 3345 27722
rect 3289 27672 3345 27700
rect 3289 27666 3320 27672
rect 3320 27666 3345 27672
rect 3377 27700 3398 27722
rect 3398 27700 3433 27722
rect 3377 27672 3433 27700
rect 3377 27666 3398 27672
rect 3398 27666 3433 27672
rect 2670 27576 2726 27632
rect 2759 27576 2815 27632
rect 2848 27620 2878 27632
rect 2878 27620 2904 27632
rect 2848 27592 2904 27620
rect 2848 27576 2878 27592
rect 2878 27576 2904 27592
rect 2937 27576 2993 27632
rect 3025 27620 3060 27632
rect 3060 27620 3081 27632
rect 3025 27592 3081 27620
rect 3025 27576 3060 27592
rect 3060 27576 3081 27592
rect 3113 27620 3138 27632
rect 3138 27620 3169 27632
rect 3113 27592 3169 27620
rect 3113 27576 3138 27592
rect 3138 27576 3169 27592
rect 3201 27576 3257 27632
rect 3289 27620 3320 27632
rect 3320 27620 3345 27632
rect 3289 27592 3345 27620
rect 3289 27576 3320 27592
rect 3320 27576 3345 27592
rect 3377 27620 3398 27632
rect 3398 27620 3433 27632
rect 3377 27592 3433 27620
rect 3377 27576 3398 27592
rect 3398 27576 3433 27592
rect 2670 27486 2726 27542
rect 2759 27486 2815 27542
rect 2848 27540 2878 27542
rect 2878 27540 2904 27542
rect 2848 27512 2904 27540
rect 2848 27486 2878 27512
rect 2878 27486 2904 27512
rect 2937 27486 2993 27542
rect 3025 27540 3060 27542
rect 3060 27540 3081 27542
rect 3025 27512 3081 27540
rect 3025 27486 3060 27512
rect 3060 27486 3081 27512
rect 3113 27540 3138 27542
rect 3138 27540 3169 27542
rect 3113 27512 3169 27540
rect 3113 27486 3138 27512
rect 3138 27486 3169 27512
rect 3201 27486 3257 27542
rect 3289 27540 3320 27542
rect 3320 27540 3345 27542
rect 3289 27512 3345 27540
rect 3289 27486 3320 27512
rect 3320 27486 3345 27512
rect 3377 27540 3398 27542
rect 3398 27540 3433 27542
rect 3377 27512 3433 27540
rect 3377 27486 3398 27512
rect 3398 27486 3433 27512
rect 2670 27396 2726 27452
rect 2759 27396 2815 27452
rect 2848 27396 2904 27452
rect 2937 27396 2993 27452
rect 3025 27396 3081 27452
rect 3113 27396 3169 27452
rect 3201 27396 3257 27452
rect 3289 27396 3345 27452
rect 3377 27396 3433 27452
rect 2494 27271 2550 27327
rect 2494 27191 2550 27247
rect 6742 26796 6798 26852
rect 6827 26796 6883 26852
rect 6912 26796 6968 26852
rect 6997 26796 7053 26852
rect 7082 26796 7138 26852
rect 7167 26796 7223 26852
rect 7252 26796 7308 26852
rect 7337 26796 7393 26852
rect 7422 26796 7478 26852
rect 7507 26796 7563 26852
rect 7591 26796 7647 26852
rect 7675 26796 7731 26852
rect 7759 26796 7815 26852
rect 7843 26796 7899 26852
rect 6742 26710 6798 26766
rect 6827 26710 6883 26766
rect 6912 26710 6968 26766
rect 6997 26710 7053 26766
rect 7082 26710 7138 26766
rect 7167 26710 7223 26766
rect 7252 26710 7308 26766
rect 7337 26710 7393 26766
rect 7422 26710 7478 26766
rect 7507 26710 7563 26766
rect 7591 26710 7647 26766
rect 7675 26710 7731 26766
rect 7759 26710 7815 26766
rect 7843 26710 7899 26766
rect 6742 26624 6798 26680
rect 6827 26624 6883 26680
rect 6912 26624 6968 26680
rect 6997 26624 7053 26680
rect 7082 26624 7138 26680
rect 7167 26624 7223 26680
rect 7252 26624 7308 26680
rect 7337 26624 7393 26680
rect 7422 26624 7478 26680
rect 7507 26624 7563 26680
rect 7591 26624 7647 26680
rect 7675 26624 7731 26680
rect 7759 26624 7815 26680
rect 7843 26624 7899 26680
rect 6742 26538 6798 26594
rect 6827 26538 6883 26594
rect 6912 26538 6968 26594
rect 6997 26538 7053 26594
rect 7082 26538 7138 26594
rect 7167 26538 7223 26594
rect 7252 26538 7308 26594
rect 7337 26538 7393 26594
rect 7422 26538 7478 26594
rect 7507 26538 7563 26594
rect 7591 26538 7647 26594
rect 7675 26538 7731 26594
rect 7759 26538 7815 26594
rect 7843 26538 7899 26594
rect 6742 26452 6798 26508
rect 6827 26452 6883 26508
rect 6912 26452 6968 26508
rect 6997 26452 7053 26508
rect 7082 26452 7138 26508
rect 7167 26452 7223 26508
rect 7252 26452 7308 26508
rect 7337 26452 7393 26508
rect 7422 26452 7478 26508
rect 7507 26452 7563 26508
rect 7591 26452 7647 26508
rect 7675 26452 7731 26508
rect 7759 26452 7815 26508
rect 7843 26452 7899 26508
rect 2670 24467 2726 24523
rect 2751 24467 2807 24523
rect 2832 24467 2888 24523
rect 2913 24467 2969 24523
rect 2994 24467 3050 24523
rect 3075 24467 3131 24523
rect 3156 24467 3212 24523
rect 3237 24467 3293 24523
rect 3318 24467 3374 24523
rect 3398 24467 3454 24523
rect 3478 24467 3534 24523
rect 2670 24341 2726 24397
rect 2751 24341 2807 24397
rect 2832 24341 2888 24397
rect 2913 24341 2969 24397
rect 2994 24341 3050 24397
rect 3075 24341 3131 24397
rect 3156 24341 3212 24397
rect 3237 24341 3293 24397
rect 3318 24341 3374 24397
rect 3398 24341 3454 24397
rect 3478 24341 3534 24397
rect 2670 23212 2726 23268
rect 2751 23212 2807 23268
rect 2832 23212 2888 23268
rect 2913 23212 2969 23268
rect 2994 23212 3050 23268
rect 3075 23212 3131 23268
rect 3156 23212 3212 23268
rect 3237 23212 3293 23268
rect 3318 23212 3374 23268
rect 3398 23212 3454 23268
rect 3478 23212 3534 23268
rect 2670 23124 2726 23180
rect 2751 23124 2807 23180
rect 2832 23124 2888 23180
rect 2913 23124 2969 23180
rect 2994 23124 3050 23180
rect 3075 23124 3131 23180
rect 3156 23124 3212 23180
rect 3237 23124 3293 23180
rect 3318 23124 3374 23180
rect 3398 23124 3454 23180
rect 3478 23124 3534 23180
rect 2670 23036 2726 23092
rect 2751 23036 2807 23092
rect 2832 23036 2888 23092
rect 2913 23036 2969 23092
rect 2994 23036 3050 23092
rect 3075 23036 3131 23092
rect 3156 23036 3212 23092
rect 3237 23036 3293 23092
rect 3318 23036 3374 23092
rect 3398 23036 3454 23092
rect 3478 23036 3534 23092
rect 2670 22948 2726 23004
rect 2751 22948 2807 23004
rect 2832 22948 2888 23004
rect 2913 22948 2969 23004
rect 2994 22948 3050 23004
rect 3075 22948 3131 23004
rect 3156 22948 3212 23004
rect 3237 22948 3293 23004
rect 3318 22948 3374 23004
rect 3398 22948 3454 23004
rect 3478 22948 3534 23004
rect 2670 22860 2726 22916
rect 2751 22860 2807 22916
rect 2832 22860 2888 22916
rect 2913 22860 2969 22916
rect 2994 22860 3050 22916
rect 3075 22860 3131 22916
rect 3156 22860 3212 22916
rect 3237 22860 3293 22916
rect 3318 22860 3374 22916
rect 3398 22860 3454 22916
rect 3478 22860 3534 22916
rect 3712 21102 3768 21158
rect 3793 21102 3849 21158
rect 3874 21102 3930 21158
rect 3955 21102 4011 21158
rect 4036 21102 4092 21158
rect 4117 21102 4173 21158
rect 4198 21102 4254 21158
rect 4278 21102 4334 21158
rect 4358 21102 4414 21158
rect 4438 21102 4494 21158
rect 3712 21016 3768 21072
rect 3793 21016 3849 21072
rect 3874 21016 3930 21072
rect 3955 21016 4011 21072
rect 4036 21016 4092 21072
rect 4117 21016 4173 21072
rect 4198 21016 4254 21072
rect 4278 21016 4334 21072
rect 4358 21016 4414 21072
rect 4438 21016 4494 21072
rect 3712 20930 3768 20986
rect 3793 20930 3849 20986
rect 3874 20930 3930 20986
rect 3955 20930 4011 20986
rect 4036 20930 4092 20986
rect 4117 20930 4173 20986
rect 4198 20930 4254 20986
rect 4278 20930 4334 20986
rect 4358 20930 4414 20986
rect 4438 20930 4494 20986
rect 3712 20844 3768 20900
rect 3793 20844 3849 20900
rect 3874 20844 3930 20900
rect 3955 20844 4011 20900
rect 4036 20844 4092 20900
rect 4117 20844 4173 20900
rect 4198 20844 4254 20900
rect 4278 20844 4334 20900
rect 4358 20844 4414 20900
rect 4438 20844 4494 20900
rect 3712 20758 3768 20814
rect 3793 20758 3849 20814
rect 3874 20758 3930 20814
rect 3955 20758 4011 20814
rect 4036 20758 4092 20814
rect 4117 20758 4173 20814
rect 4198 20758 4254 20814
rect 4278 20758 4334 20814
rect 4358 20758 4414 20814
rect 4438 20758 4494 20814
rect 3712 19039 3768 19095
rect 3793 19039 3849 19095
rect 3874 19039 3930 19095
rect 3955 19039 4011 19095
rect 4036 19039 4092 19095
rect 4117 19039 4173 19095
rect 4198 19039 4254 19095
rect 4278 19039 4334 19095
rect 4358 19039 4414 19095
rect 4438 19039 4494 19095
rect 3712 18895 3768 18951
rect 3793 18895 3849 18951
rect 3874 18895 3930 18951
rect 3955 18895 4011 18951
rect 4036 18895 4092 18951
rect 4117 18895 4173 18951
rect 4198 18895 4254 18951
rect 4278 18895 4334 18951
rect 4358 18895 4414 18951
rect 4438 18895 4494 18951
rect 5832 18206 5888 18262
rect 5914 18206 5970 18262
rect 5995 18206 6051 18262
rect 6076 18206 6132 18262
rect 6157 18206 6213 18262
rect 6238 18206 6294 18262
rect 6319 18206 6375 18262
rect 6400 18206 6456 18262
rect 6481 18206 6537 18262
rect 6562 18206 6618 18262
rect 5832 18126 5888 18182
rect 5914 18126 5970 18182
rect 5995 18126 6051 18182
rect 6076 18126 6132 18182
rect 6157 18126 6213 18182
rect 6238 18126 6294 18182
rect 6319 18126 6375 18182
rect 6400 18126 6456 18182
rect 6481 18126 6537 18182
rect 6562 18126 6618 18182
rect 3712 17280 3768 17336
rect 3793 17280 3849 17336
rect 3874 17280 3930 17336
rect 3955 17280 4011 17336
rect 4036 17280 4092 17336
rect 4117 17280 4173 17336
rect 4198 17280 4254 17336
rect 4278 17280 4334 17336
rect 4358 17280 4414 17336
rect 4438 17280 4494 17336
rect 3712 17194 3768 17250
rect 3793 17194 3849 17250
rect 3874 17194 3930 17250
rect 3955 17194 4011 17250
rect 4036 17194 4092 17250
rect 4117 17194 4173 17250
rect 4198 17194 4254 17250
rect 4278 17194 4334 17250
rect 4358 17194 4414 17250
rect 4438 17194 4494 17250
rect 3712 17108 3768 17164
rect 3793 17108 3849 17164
rect 3874 17108 3930 17164
rect 3955 17108 4011 17164
rect 4036 17108 4092 17164
rect 4117 17108 4173 17164
rect 4198 17108 4254 17164
rect 4278 17108 4334 17164
rect 4358 17108 4414 17164
rect 4438 17108 4494 17164
rect 3712 17022 3768 17078
rect 3793 17022 3849 17078
rect 3874 17022 3930 17078
rect 3955 17022 4011 17078
rect 4036 17022 4092 17078
rect 4117 17022 4173 17078
rect 4198 17022 4254 17078
rect 4278 17022 4334 17078
rect 4358 17022 4414 17078
rect 4438 17022 4494 17078
rect 3712 16936 3768 16992
rect 3793 16936 3849 16992
rect 3874 16936 3930 16992
rect 3955 16936 4011 16992
rect 4036 16936 4092 16992
rect 4117 16936 4173 16992
rect 4198 16936 4254 16992
rect 4278 16936 4334 16992
rect 4358 16936 4414 16992
rect 4438 16936 4494 16992
rect 10135 15533 10191 15589
rect 10135 15453 10191 15509
rect 3712 15165 3768 15221
rect 3793 15165 3849 15221
rect 3874 15165 3930 15221
rect 3955 15165 4011 15221
rect 4036 15165 4092 15221
rect 4117 15165 4173 15221
rect 3712 15085 3768 15141
rect 3793 15085 3849 15141
rect 3874 15085 3930 15141
rect 3955 15085 4011 15141
rect 4036 15085 4092 15141
rect 4117 15085 4173 15141
rect 3712 15005 3768 15061
rect 3793 15005 3849 15061
rect 3874 15005 3930 15061
rect 3955 15005 4011 15061
rect 4036 15005 4092 15061
rect 4117 15005 4173 15061
rect 3712 14925 3768 14981
rect 3793 14925 3849 14981
rect 3874 14925 3930 14981
rect 3955 14925 4011 14981
rect 4036 14925 4092 14981
rect 4117 14925 4173 14981
rect 4198 14925 4494 15221
rect 2670 14555 2726 14611
rect 2751 14555 2807 14611
rect 2832 14555 2888 14611
rect 2913 14555 2969 14611
rect 2994 14555 3050 14611
rect 3075 14555 3131 14611
rect 3156 14555 3212 14611
rect 3237 14555 3293 14611
rect 3318 14555 3374 14611
rect 3398 14555 3454 14611
rect 3478 14555 3534 14611
rect 2670 14471 2726 14527
rect 2751 14471 2807 14527
rect 2832 14471 2888 14527
rect 2913 14471 2969 14527
rect 2994 14471 3050 14527
rect 3075 14471 3131 14527
rect 3156 14471 3212 14527
rect 3237 14471 3293 14527
rect 3318 14471 3374 14527
rect 3398 14471 3454 14527
rect 3478 14471 3534 14527
rect 2670 14387 2726 14443
rect 2751 14387 2807 14443
rect 2832 14387 2888 14443
rect 2913 14387 2969 14443
rect 2994 14387 3050 14443
rect 3075 14387 3131 14443
rect 3156 14387 3212 14443
rect 3237 14387 3293 14443
rect 3318 14387 3374 14443
rect 3398 14387 3454 14443
rect 3478 14387 3534 14443
rect 6779 12569 6835 12625
rect 6859 12569 6915 12625
rect 10135 12604 10191 12660
rect 10135 12480 10191 12536
rect 6779 12093 6835 12095
rect 6859 12093 6915 12095
rect 6779 12041 6828 12093
rect 6828 12041 6835 12093
rect 6859 12041 6892 12093
rect 6892 12041 6915 12093
rect 6779 12039 6835 12041
rect 6859 12039 6915 12041
rect 2670 11645 2719 11697
rect 2719 11645 2726 11697
rect 2751 11645 2788 11697
rect 2788 11645 2805 11697
rect 2805 11645 2807 11697
rect 2832 11645 2857 11697
rect 2857 11645 2873 11697
rect 2873 11645 2888 11697
rect 2913 11645 2925 11697
rect 2925 11645 2941 11697
rect 2941 11645 2969 11697
rect 2994 11645 3009 11697
rect 3009 11645 3050 11697
rect 3075 11645 3077 11697
rect 3077 11645 3129 11697
rect 3129 11645 3131 11697
rect 3156 11645 3197 11697
rect 3197 11645 3212 11697
rect 3237 11645 3265 11697
rect 3265 11645 3281 11697
rect 3281 11645 3293 11697
rect 3318 11645 3333 11697
rect 3333 11645 3349 11697
rect 3349 11645 3374 11697
rect 3398 11645 3401 11697
rect 3401 11645 3417 11697
rect 3417 11645 3454 11697
rect 3478 11645 3485 11697
rect 3485 11645 3534 11697
rect 2670 11641 2726 11645
rect 2751 11641 2807 11645
rect 2832 11641 2888 11645
rect 2913 11641 2969 11645
rect 2994 11641 3050 11645
rect 3075 11641 3131 11645
rect 3156 11641 3212 11645
rect 3237 11641 3293 11645
rect 3318 11641 3374 11645
rect 3398 11641 3454 11645
rect 3478 11641 3534 11645
rect 2670 11611 2726 11615
rect 2751 11611 2807 11615
rect 2832 11611 2888 11615
rect 2913 11611 2969 11615
rect 2994 11611 3050 11615
rect 3075 11611 3131 11615
rect 3156 11611 3212 11615
rect 3237 11611 3293 11615
rect 3318 11611 3374 11615
rect 3398 11611 3454 11615
rect 3478 11611 3534 11615
rect 2670 11559 2719 11611
rect 2719 11559 2726 11611
rect 2751 11559 2788 11611
rect 2788 11559 2805 11611
rect 2805 11559 2807 11611
rect 2832 11559 2857 11611
rect 2857 11559 2873 11611
rect 2873 11559 2888 11611
rect 2913 11559 2925 11611
rect 2925 11559 2941 11611
rect 2941 11559 2969 11611
rect 2994 11559 3009 11611
rect 3009 11559 3050 11611
rect 3075 11559 3077 11611
rect 3077 11559 3129 11611
rect 3129 11559 3131 11611
rect 3156 11559 3197 11611
rect 3197 11559 3212 11611
rect 3237 11559 3265 11611
rect 3265 11559 3281 11611
rect 3281 11559 3293 11611
rect 3318 11559 3333 11611
rect 3333 11559 3349 11611
rect 3349 11559 3374 11611
rect 3398 11559 3401 11611
rect 3401 11559 3417 11611
rect 3417 11559 3454 11611
rect 3478 11559 3485 11611
rect 3485 11559 3534 11611
rect 632 11075 688 11131
rect 713 11075 769 11131
rect 794 11075 850 11131
rect 875 11075 931 11131
rect 956 11075 1012 11131
rect 1037 11075 1093 11131
rect 1118 11075 1174 11131
rect 1198 11075 1254 11131
rect 1278 11075 1334 11131
rect 1358 11075 1414 11131
rect 6714 11218 6770 11274
rect 6714 11138 6770 11194
rect 6840 11133 6896 11189
rect 6840 11053 6896 11109
rect 632 10785 688 10841
rect 713 10785 769 10841
rect 794 10785 850 10841
rect 875 10785 931 10841
rect 956 10785 1012 10841
rect 1037 10785 1093 10841
rect 1118 10785 1174 10841
rect 1198 10785 1254 10841
rect 1278 10785 1334 10841
rect 1358 10785 1414 10841
rect 632 10649 688 10705
rect 713 10649 769 10705
rect 794 10649 850 10705
rect 875 10649 931 10705
rect 956 10649 1012 10705
rect 1037 10649 1093 10705
rect 1118 10649 1174 10705
rect 1198 10649 1254 10705
rect 1278 10649 1334 10705
rect 1358 10649 1414 10705
rect 8767 10635 8823 10639
rect 8847 10635 8903 10639
rect 8553 10633 8609 10635
rect 8633 10633 8689 10635
rect 8553 10581 8576 10633
rect 8576 10581 8609 10633
rect 8633 10581 8640 10633
rect 8640 10581 8689 10633
rect 8767 10583 8816 10635
rect 8816 10583 8823 10635
rect 8847 10583 8898 10635
rect 8898 10583 8903 10635
rect 8553 10579 8609 10581
rect 8633 10579 8689 10581
rect 10261 10512 10317 10568
rect 10261 10432 10317 10488
rect 8383 10304 8439 10360
rect 8463 10304 8519 10360
rect 8916 10100 8972 10156
rect 8916 10020 8972 10076
rect 632 9757 688 9813
rect 713 9757 769 9813
rect 794 9757 850 9813
rect 875 9757 931 9813
rect 956 9757 1012 9813
rect 1037 9757 1093 9813
rect 1118 9757 1174 9813
rect 1198 9757 1254 9813
rect 1278 9757 1334 9813
rect 1358 9757 1414 9813
rect 7943 9604 7999 9660
rect 8023 9604 8079 9660
rect 637 8097 693 8153
rect 718 8097 774 8153
rect 798 8097 854 8153
rect 878 8097 934 8153
rect 958 8097 1014 8153
rect 1038 8097 1094 8153
rect 1118 8097 1174 8153
rect 1198 8097 1254 8153
rect 1278 8097 1334 8153
rect 1358 8097 1414 8153
rect 637 7971 693 8027
rect 718 7971 774 8027
rect 798 7971 854 8027
rect 878 7971 934 8027
rect 958 7971 1014 8027
rect 1038 7971 1094 8027
rect 1118 7971 1174 8027
rect 1198 7971 1254 8027
rect 1278 7971 1334 8027
rect 1358 7971 1414 8027
rect 5832 7881 5888 7937
rect 5913 7881 5969 7937
rect 5994 7881 6050 7937
rect 6075 7881 6131 7937
rect 6156 7881 6212 7937
rect 6237 7881 6293 7937
rect 6318 7881 6374 7937
rect 6398 7881 6454 7937
rect 6478 7881 6534 7937
rect 6558 7881 6614 7937
rect 5832 7789 5888 7845
rect 5913 7789 5969 7845
rect 5994 7789 6050 7845
rect 6075 7789 6131 7845
rect 6156 7789 6212 7845
rect 6237 7789 6293 7845
rect 6318 7789 6374 7845
rect 6398 7789 6454 7845
rect 6478 7789 6534 7845
rect 6558 7789 6614 7845
rect 291 7667 347 7723
rect 374 7667 430 7723
rect 456 7667 512 7723
rect 538 7667 594 7723
rect 620 7667 676 7723
rect 702 7667 758 7723
rect 784 7667 840 7723
rect 866 7667 922 7723
rect 948 7667 1004 7723
rect 1030 7667 1086 7723
rect 1112 7667 1168 7723
rect 1194 7667 1250 7723
rect 1276 7667 1332 7723
rect 1358 7667 1414 7723
rect 2714 7700 2770 7756
rect 2794 7700 2850 7756
rect 2874 7700 2930 7756
rect 2954 7700 3010 7756
rect 3034 7700 3090 7756
rect 3114 7700 3170 7756
rect 3194 7700 3250 7756
rect 3274 7700 3330 7756
rect 3354 7700 3410 7756
rect 3434 7700 3490 7756
rect 291 7581 347 7637
rect 374 7581 430 7637
rect 456 7581 512 7637
rect 538 7581 594 7637
rect 620 7581 676 7637
rect 702 7581 758 7637
rect 784 7581 840 7637
rect 866 7581 922 7637
rect 948 7581 1004 7637
rect 1030 7581 1086 7637
rect 1112 7581 1168 7637
rect 1194 7581 1250 7637
rect 1276 7581 1332 7637
rect 1358 7581 1414 7637
rect 2714 7616 2770 7672
rect 2794 7616 2850 7672
rect 2874 7616 2930 7672
rect 2954 7616 3010 7672
rect 3034 7616 3090 7672
rect 3114 7616 3170 7672
rect 3194 7616 3250 7672
rect 3274 7616 3330 7672
rect 3354 7616 3410 7672
rect 3434 7616 3490 7672
rect 291 7495 347 7551
rect 374 7495 430 7551
rect 456 7495 512 7551
rect 538 7495 594 7551
rect 620 7495 676 7551
rect 702 7495 758 7551
rect 784 7495 840 7551
rect 866 7495 922 7551
rect 948 7495 1004 7551
rect 1030 7495 1086 7551
rect 1112 7495 1168 7551
rect 1194 7495 1250 7551
rect 1276 7495 1332 7551
rect 1358 7495 1414 7551
rect 2714 7532 2770 7588
rect 2794 7532 2850 7588
rect 2874 7532 2930 7588
rect 2954 7532 3010 7588
rect 3034 7532 3090 7588
rect 3114 7532 3170 7588
rect 3194 7532 3250 7588
rect 3274 7532 3330 7588
rect 3354 7532 3410 7588
rect 3434 7532 3490 7588
rect 291 7409 347 7465
rect 374 7409 430 7465
rect 456 7409 512 7465
rect 538 7409 594 7465
rect 620 7409 676 7465
rect 702 7409 758 7465
rect 784 7409 840 7465
rect 866 7409 922 7465
rect 948 7409 1004 7465
rect 1030 7409 1086 7465
rect 1112 7409 1168 7465
rect 1194 7409 1250 7465
rect 1276 7409 1332 7465
rect 1358 7409 1414 7465
rect 2714 7448 2770 7504
rect 2794 7448 2850 7504
rect 2874 7448 2930 7504
rect 2954 7448 3010 7504
rect 3034 7448 3090 7504
rect 3114 7448 3170 7504
rect 3194 7448 3250 7504
rect 3274 7448 3330 7504
rect 3354 7448 3410 7504
rect 3434 7448 3490 7504
rect 291 7323 347 7379
rect 374 7323 430 7379
rect 456 7323 512 7379
rect 538 7323 594 7379
rect 620 7323 676 7379
rect 702 7323 758 7379
rect 784 7323 840 7379
rect 866 7323 922 7379
rect 948 7323 1004 7379
rect 1030 7323 1086 7379
rect 1112 7323 1168 7379
rect 1194 7323 1250 7379
rect 1276 7323 1332 7379
rect 1358 7323 1414 7379
rect 2714 7364 2770 7420
rect 2794 7364 2850 7420
rect 2874 7364 2930 7420
rect 2954 7364 3010 7420
rect 3034 7364 3090 7420
rect 3114 7364 3170 7420
rect 3194 7364 3250 7420
rect 3274 7364 3330 7420
rect 3354 7364 3410 7420
rect 3434 7364 3490 7420
rect 291 7237 347 7293
rect 374 7237 430 7293
rect 456 7237 512 7293
rect 538 7237 594 7293
rect 620 7237 676 7293
rect 702 7237 758 7293
rect 784 7237 840 7293
rect 866 7237 922 7293
rect 948 7237 1004 7293
rect 1030 7237 1086 7293
rect 1112 7237 1168 7293
rect 1194 7237 1250 7293
rect 1276 7237 1332 7293
rect 1358 7237 1414 7293
rect 2714 7280 2770 7336
rect 2794 7280 2850 7336
rect 2874 7280 2930 7336
rect 2954 7280 3010 7336
rect 3034 7280 3090 7336
rect 3114 7280 3170 7336
rect 3194 7280 3250 7336
rect 3274 7280 3330 7336
rect 3354 7280 3410 7336
rect 3434 7280 3490 7336
rect 291 7151 347 7207
rect 374 7151 430 7207
rect 456 7151 512 7207
rect 538 7151 594 7207
rect 620 7151 676 7207
rect 702 7151 758 7207
rect 784 7151 840 7207
rect 866 7151 922 7207
rect 948 7151 1004 7207
rect 1030 7151 1086 7207
rect 1112 7151 1168 7207
rect 1194 7151 1250 7207
rect 1276 7151 1332 7207
rect 1358 7151 1414 7207
rect 2714 7196 2770 7252
rect 2794 7196 2850 7252
rect 2874 7196 2930 7252
rect 2954 7196 3010 7252
rect 3034 7196 3090 7252
rect 3114 7196 3170 7252
rect 3194 7196 3250 7252
rect 3274 7196 3330 7252
rect 3354 7196 3410 7252
rect 3434 7196 3490 7252
rect 6840 7280 6896 7336
rect 6840 7200 6896 7256
rect 291 7065 347 7121
rect 374 7065 430 7121
rect 456 7065 512 7121
rect 538 7065 594 7121
rect 620 7065 676 7121
rect 702 7065 758 7121
rect 784 7065 840 7121
rect 866 7065 922 7121
rect 948 7065 1004 7121
rect 1030 7065 1086 7121
rect 1112 7065 1168 7121
rect 1194 7065 1250 7121
rect 1276 7065 1332 7121
rect 1358 7065 1414 7121
rect 2714 7112 2770 7168
rect 2794 7112 2850 7168
rect 2874 7112 2930 7168
rect 2954 7112 3010 7168
rect 3034 7112 3090 7168
rect 3114 7112 3170 7168
rect 3194 7112 3250 7168
rect 3274 7112 3330 7168
rect 3354 7112 3410 7168
rect 3434 7112 3490 7168
rect 291 6979 347 7035
rect 374 6979 430 7035
rect 456 6979 512 7035
rect 538 6979 594 7035
rect 620 6979 676 7035
rect 702 6979 758 7035
rect 784 6979 840 7035
rect 866 6979 922 7035
rect 948 6979 1004 7035
rect 1030 6979 1086 7035
rect 1112 6979 1168 7035
rect 1194 6979 1250 7035
rect 1276 6979 1332 7035
rect 1358 6979 1414 7035
rect 2714 7028 2770 7084
rect 2794 7028 2850 7084
rect 2874 7028 2930 7084
rect 2954 7028 3010 7084
rect 3034 7028 3090 7084
rect 3114 7028 3170 7084
rect 3194 7028 3250 7084
rect 3274 7028 3330 7084
rect 3354 7028 3410 7084
rect 3434 7028 3490 7084
rect 291 6893 347 6949
rect 374 6893 430 6949
rect 456 6893 512 6949
rect 538 6893 594 6949
rect 620 6893 676 6949
rect 702 6893 758 6949
rect 784 6893 840 6949
rect 866 6893 922 6949
rect 948 6893 1004 6949
rect 1030 6893 1086 6949
rect 1112 6893 1168 6949
rect 1194 6893 1250 6949
rect 1276 6893 1332 6949
rect 1358 6893 1414 6949
rect 2714 6944 2770 7000
rect 2794 6944 2850 7000
rect 2874 6944 2930 7000
rect 2954 6944 3010 7000
rect 3034 6944 3090 7000
rect 3114 6944 3170 7000
rect 3194 6944 3250 7000
rect 3274 6944 3330 7000
rect 3354 6944 3410 7000
rect 3434 6944 3490 7000
rect 6714 7006 6770 7062
rect 6714 6926 6770 6982
rect 291 6807 347 6863
rect 374 6807 430 6863
rect 456 6807 512 6863
rect 538 6807 594 6863
rect 620 6807 676 6863
rect 702 6807 758 6863
rect 784 6807 840 6863
rect 866 6807 922 6863
rect 948 6807 1004 6863
rect 1030 6807 1086 6863
rect 1112 6807 1168 6863
rect 1194 6807 1250 6863
rect 1276 6807 1332 6863
rect 1358 6807 1414 6863
rect 2714 6859 2770 6915
rect 2794 6859 2850 6915
rect 2874 6859 2930 6915
rect 2954 6859 3010 6915
rect 3034 6859 3090 6915
rect 3114 6859 3170 6915
rect 3194 6859 3250 6915
rect 3274 6859 3330 6915
rect 3354 6859 3410 6915
rect 3434 6859 3490 6915
rect 2714 6774 2770 6830
rect 2794 6774 2850 6830
rect 2874 6774 2930 6830
rect 2954 6774 3010 6830
rect 3034 6774 3090 6830
rect 3114 6774 3170 6830
rect 3194 6774 3250 6830
rect 3274 6774 3330 6830
rect 3354 6774 3410 6830
rect 3434 6774 3490 6830
rect 6507 6068 6563 6124
rect 6587 6068 6643 6124
rect 6507 5976 6563 6032
rect 6587 5976 6643 6032
rect 6507 5884 6563 5940
rect 6587 5884 6643 5940
rect 6507 5792 6563 5848
rect 6587 5792 6643 5848
rect 6507 5700 6563 5756
rect 6587 5700 6643 5756
rect 6507 5608 6563 5664
rect 6587 5608 6643 5664
rect 6507 5515 6563 5571
rect 6587 5515 6643 5571
rect 10261 5181 10317 5237
rect 10261 5101 10317 5157
rect 6459 3995 6515 4051
rect 6561 3995 6617 4051
rect 6663 3995 6719 4051
rect 6459 3914 6515 3970
rect 6561 3914 6617 3970
rect 6663 3914 6719 3970
rect 6459 3833 6515 3889
rect 6561 3833 6617 3889
rect 6663 3833 6719 3889
rect 6459 3751 6515 3807
rect 6561 3751 6617 3807
rect 6663 3751 6719 3807
rect 6459 3669 6515 3725
rect 6561 3669 6617 3725
rect 6663 3669 6719 3725
rect 8023 3813 8079 3869
rect 8023 3733 8079 3789
rect 5832 3265 5888 3321
rect 5914 3265 5970 3321
rect 5995 3265 6051 3321
rect 6076 3265 6132 3321
rect 6157 3265 6213 3321
rect 6238 3265 6294 3321
rect 6319 3265 6375 3321
rect 6400 3265 6456 3321
rect 6481 3265 6537 3321
rect 6562 3265 6618 3321
rect 5832 3185 5888 3241
rect 5914 3185 5970 3241
rect 5995 3185 6051 3241
rect 6076 3185 6132 3241
rect 6157 3185 6213 3241
rect 6238 3185 6294 3241
rect 6319 3185 6375 3241
rect 6400 3185 6456 3241
rect 6481 3185 6537 3241
rect 6562 3185 6618 3241
rect 5832 3136 5888 3137
rect 5914 3136 5970 3137
rect 5995 3136 6051 3137
rect 6076 3136 6132 3137
rect 6157 3136 6213 3137
rect 6238 3136 6294 3137
rect 6319 3136 6375 3137
rect 6400 3136 6456 3137
rect 6481 3136 6537 3137
rect 6562 3136 6618 3137
rect 5832 3084 5882 3136
rect 5882 3084 5888 3136
rect 5914 3084 5949 3136
rect 5949 3084 5964 3136
rect 5964 3084 5970 3136
rect 5995 3084 6016 3136
rect 6016 3084 6031 3136
rect 6031 3084 6051 3136
rect 6076 3084 6083 3136
rect 6083 3084 6098 3136
rect 6098 3084 6132 3136
rect 6157 3084 6165 3136
rect 6165 3084 6213 3136
rect 6238 3084 6284 3136
rect 6284 3084 6294 3136
rect 6319 3084 6351 3136
rect 6351 3084 6366 3136
rect 6366 3084 6375 3136
rect 6400 3084 6418 3136
rect 6418 3084 6433 3136
rect 6433 3084 6456 3136
rect 6481 3084 6485 3136
rect 6485 3084 6499 3136
rect 6499 3084 6537 3136
rect 6562 3084 6565 3136
rect 6565 3084 6617 3136
rect 6617 3084 6618 3136
rect 8916 3239 8972 3295
rect 8916 3159 8972 3215
rect 5832 3081 5888 3084
rect 5914 3081 5970 3084
rect 5995 3081 6051 3084
rect 6076 3081 6132 3084
rect 6157 3081 6213 3084
rect 6238 3081 6294 3084
rect 6319 3081 6375 3084
rect 6400 3081 6456 3084
rect 6481 3081 6537 3084
rect 6562 3081 6618 3084
rect 5832 3048 5888 3057
rect 5914 3048 5970 3057
rect 5995 3048 6051 3057
rect 6076 3048 6132 3057
rect 6157 3048 6213 3057
rect 6238 3048 6294 3057
rect 6319 3048 6375 3057
rect 6400 3048 6456 3057
rect 6481 3048 6537 3057
rect 6562 3048 6618 3057
rect 5832 3001 5882 3048
rect 5882 3001 5888 3048
rect 5914 3001 5949 3048
rect 5949 3001 5964 3048
rect 5964 3001 5970 3048
rect 5995 3001 6016 3048
rect 6016 3001 6031 3048
rect 6031 3001 6051 3048
rect 6076 3001 6083 3048
rect 6083 3001 6098 3048
rect 6098 3001 6132 3048
rect 6157 3001 6165 3048
rect 6165 3001 6213 3048
rect 6238 3001 6284 3048
rect 6284 3001 6294 3048
rect 6319 3001 6351 3048
rect 6351 3001 6366 3048
rect 6366 3001 6375 3048
rect 6400 3001 6418 3048
rect 6418 3001 6433 3048
rect 6433 3001 6456 3048
rect 6481 3001 6485 3048
rect 6485 3001 6499 3048
rect 6499 3001 6537 3048
rect 6562 3001 6565 3048
rect 6565 3001 6617 3048
rect 6617 3001 6618 3048
rect 3712 1464 3715 1516
rect 3715 1464 3731 1516
rect 3731 1464 3768 1516
rect 3798 1464 3799 1516
rect 3799 1464 3851 1516
rect 3851 1464 3854 1516
rect 3884 1464 3919 1516
rect 3919 1464 3934 1516
rect 3934 1464 3940 1516
rect 3970 1464 3986 1516
rect 3986 1464 4001 1516
rect 4001 1464 4026 1516
rect 4056 1464 4068 1516
rect 4068 1464 4112 1516
rect 3712 1460 3768 1464
rect 3798 1460 3854 1464
rect 3884 1460 3940 1464
rect 3970 1460 4026 1464
rect 4056 1460 4112 1464
rect 4142 1460 4198 1516
rect 4228 1460 4284 1516
rect 4314 1460 4370 1516
rect 4399 1460 4455 1516
rect 3712 1400 3715 1432
rect 3715 1400 3731 1432
rect 3731 1400 3768 1432
rect 3798 1400 3799 1432
rect 3799 1400 3851 1432
rect 3851 1400 3854 1432
rect 3884 1400 3919 1432
rect 3919 1400 3934 1432
rect 3934 1400 3940 1432
rect 3970 1400 3986 1432
rect 3986 1400 4001 1432
rect 4001 1400 4026 1432
rect 4056 1400 4068 1432
rect 4068 1400 4112 1432
rect 3712 1388 3768 1400
rect 3798 1388 3854 1400
rect 3884 1388 3940 1400
rect 3970 1388 4026 1400
rect 4056 1388 4112 1400
rect 3712 1376 3715 1388
rect 3715 1376 3731 1388
rect 3731 1376 3768 1388
rect 3798 1376 3799 1388
rect 3799 1376 3851 1388
rect 3851 1376 3854 1388
rect 3884 1376 3919 1388
rect 3919 1376 3934 1388
rect 3934 1376 3940 1388
rect 3970 1376 3986 1388
rect 3986 1376 4001 1388
rect 4001 1376 4026 1388
rect 4056 1376 4068 1388
rect 4068 1376 4112 1388
rect 4142 1376 4198 1432
rect 4228 1376 4284 1432
rect 4314 1376 4370 1432
rect 4399 1376 4455 1432
rect 3712 1336 3715 1348
rect 3715 1336 3731 1348
rect 3731 1336 3768 1348
rect 3798 1336 3799 1348
rect 3799 1336 3851 1348
rect 3851 1336 3854 1348
rect 3884 1336 3919 1348
rect 3919 1336 3934 1348
rect 3934 1336 3940 1348
rect 3970 1336 3986 1348
rect 3986 1336 4001 1348
rect 4001 1336 4026 1348
rect 4056 1336 4068 1348
rect 4068 1336 4112 1348
rect 3712 1324 3768 1336
rect 3798 1324 3854 1336
rect 3884 1324 3940 1336
rect 3970 1324 4026 1336
rect 4056 1324 4112 1336
rect 3712 1292 3715 1324
rect 3715 1292 3731 1324
rect 3731 1292 3768 1324
rect 3798 1292 3799 1324
rect 3799 1292 3851 1324
rect 3851 1292 3854 1324
rect 3884 1292 3919 1324
rect 3919 1292 3934 1324
rect 3934 1292 3940 1324
rect 3970 1292 3986 1324
rect 3986 1292 4001 1324
rect 4001 1292 4026 1324
rect 4056 1292 4068 1324
rect 4068 1292 4112 1324
rect 4142 1292 4198 1348
rect 4228 1292 4284 1348
rect 4314 1292 4370 1348
rect 4399 1292 4455 1348
rect 7009 1694 7034 1711
rect 7034 1694 7065 1711
rect 7137 1694 7182 1711
rect 7182 1694 7193 1711
rect 7265 1694 7282 1711
rect 7282 1694 7321 1711
rect 7393 1694 7434 1711
rect 7434 1694 7449 1711
rect 7521 1694 7534 1711
rect 7534 1694 7577 1711
rect 7649 1694 7682 1711
rect 7682 1694 7705 1711
rect 7776 1694 7782 1711
rect 7782 1694 7832 1711
rect 7009 1672 7065 1694
rect 7137 1672 7193 1694
rect 7265 1672 7321 1694
rect 7393 1672 7449 1694
rect 7521 1672 7577 1694
rect 7649 1672 7705 1694
rect 7776 1672 7832 1694
rect 7009 1655 7034 1672
rect 7034 1655 7065 1672
rect 7137 1655 7182 1672
rect 7182 1655 7193 1672
rect 7265 1655 7282 1672
rect 7282 1655 7321 1672
rect 7393 1655 7434 1672
rect 7434 1655 7449 1672
rect 7521 1655 7534 1672
rect 7534 1655 7577 1672
rect 7649 1655 7682 1672
rect 7682 1655 7705 1672
rect 7776 1655 7782 1672
rect 7782 1655 7832 1672
rect 3712 1260 3768 1264
rect 3798 1260 3854 1264
rect 3884 1260 3940 1264
rect 3970 1260 4026 1264
rect 4056 1260 4112 1264
rect 3712 1208 3715 1260
rect 3715 1208 3731 1260
rect 3731 1208 3768 1260
rect 3798 1208 3799 1260
rect 3799 1208 3851 1260
rect 3851 1208 3854 1260
rect 3884 1208 3919 1260
rect 3919 1208 3934 1260
rect 3934 1208 3940 1260
rect 3970 1208 3986 1260
rect 3986 1208 4001 1260
rect 4001 1208 4026 1260
rect 4056 1208 4068 1260
rect 4068 1208 4112 1260
rect 4142 1208 4198 1264
rect 4228 1208 4284 1264
rect 4314 1208 4370 1264
rect 4399 1208 4455 1264
rect 5832 1048 5888 1050
rect 5913 1048 5969 1050
rect 5994 1048 6050 1050
rect 6075 1048 6131 1050
rect 6156 1048 6212 1050
rect 6237 1048 6293 1050
rect 6318 1048 6374 1050
rect 6398 1048 6454 1050
rect 6478 1048 6534 1050
rect 6558 1048 6614 1050
rect 5832 996 5881 1048
rect 5881 996 5888 1048
rect 5913 996 5948 1048
rect 5948 996 5963 1048
rect 5963 996 5969 1048
rect 5994 996 6015 1048
rect 6015 996 6030 1048
rect 6030 996 6050 1048
rect 6075 996 6082 1048
rect 6082 996 6097 1048
rect 6097 996 6131 1048
rect 6156 996 6164 1048
rect 6164 996 6212 1048
rect 6237 996 6283 1048
rect 6283 996 6293 1048
rect 6318 996 6350 1048
rect 6350 996 6365 1048
rect 6365 996 6374 1048
rect 6398 996 6417 1048
rect 6417 996 6432 1048
rect 6432 996 6454 1048
rect 6478 996 6484 1048
rect 6484 996 6499 1048
rect 6499 996 6534 1048
rect 6558 996 6565 1048
rect 6565 996 6614 1048
rect 5832 994 5888 996
rect 5913 994 5969 996
rect 5994 994 6050 996
rect 6075 994 6131 996
rect 6156 994 6212 996
rect 6237 994 6293 996
rect 6318 994 6374 996
rect 6398 994 6454 996
rect 6478 994 6534 996
rect 6558 994 6614 996
rect 8763 1030 8819 1086
rect 8763 950 8819 1006
rect 2494 106 2496 145
rect 2496 106 2548 145
rect 2548 106 2550 145
rect 2494 89 2550 106
rect 2494 58 2550 65
rect 2494 9 2496 58
rect 2496 9 2548 58
rect 2548 9 2550 58
rect 6840 122 6896 145
rect 6840 89 6843 122
rect 6843 89 6895 122
rect 6895 89 6896 122
rect 6840 58 6896 65
rect 6840 9 6843 58
rect 6843 9 6895 58
rect 6895 9 6896 58
rect 8467 122 8523 145
rect 8467 89 8469 122
rect 8469 89 8521 122
rect 8521 89 8523 122
rect 8467 58 8523 65
rect 8467 9 8469 58
rect 8469 9 8521 58
rect 8521 9 8523 58
rect 8700 122 8756 145
rect 8700 89 8701 122
rect 8701 89 8753 122
rect 8753 89 8756 122
rect 8700 58 8756 65
rect 8700 9 8701 58
rect 8701 9 8753 58
rect 8753 9 8756 58
rect 8916 122 8972 145
rect 8916 89 8918 122
rect 8918 89 8970 122
rect 8970 89 8972 122
rect 8916 58 8972 65
rect 8916 9 8918 58
rect 8918 9 8970 58
rect 8970 9 8972 58
rect 10029 122 10085 145
rect 10029 89 10031 122
rect 10031 89 10083 122
rect 10083 89 10085 122
rect 10029 58 10085 65
rect 10029 9 10031 58
rect 10031 9 10083 58
rect 10083 9 10085 58
rect 10261 122 10317 145
rect 10261 89 10263 122
rect 10263 89 10315 122
rect 10315 89 10317 122
rect 10261 58 10317 65
rect 10261 9 10263 58
rect 10263 9 10315 58
rect 10315 9 10317 58
<< metal3 >>
rect 282 38946 1423 40000
rect 282 38890 291 38946
rect 347 38890 374 38946
rect 430 38890 456 38946
rect 512 38890 538 38946
rect 594 38890 620 38946
rect 676 38890 702 38946
rect 758 38890 784 38946
rect 840 38890 866 38946
rect 922 38890 948 38946
rect 1004 38890 1030 38946
rect 1086 38890 1112 38946
rect 1168 38890 1194 38946
rect 1250 38890 1276 38946
rect 1332 38890 1358 38946
rect 1414 38890 1423 38946
rect 282 38860 1423 38890
rect 282 38804 291 38860
rect 347 38804 374 38860
rect 430 38804 456 38860
rect 512 38804 538 38860
rect 594 38804 620 38860
rect 676 38804 702 38860
rect 758 38804 784 38860
rect 840 38804 866 38860
rect 922 38804 948 38860
rect 1004 38804 1030 38860
rect 1086 38804 1112 38860
rect 1168 38804 1194 38860
rect 1250 38804 1276 38860
rect 1332 38804 1358 38860
rect 1414 38804 1423 38860
rect 282 38774 1423 38804
rect 282 38718 291 38774
rect 347 38718 374 38774
rect 430 38718 456 38774
rect 512 38718 538 38774
rect 594 38718 620 38774
rect 676 38718 702 38774
rect 758 38718 784 38774
rect 840 38718 866 38774
rect 922 38718 948 38774
rect 1004 38718 1030 38774
rect 1086 38718 1112 38774
rect 1168 38718 1194 38774
rect 1250 38718 1276 38774
rect 1332 38718 1358 38774
rect 1414 38718 1423 38774
rect 282 38688 1423 38718
rect 282 38632 291 38688
rect 347 38632 374 38688
rect 430 38632 456 38688
rect 512 38632 538 38688
rect 594 38632 620 38688
rect 676 38632 702 38688
rect 758 38632 784 38688
rect 840 38632 866 38688
rect 922 38632 948 38688
rect 1004 38632 1030 38688
rect 1086 38632 1112 38688
rect 1168 38632 1194 38688
rect 1250 38632 1276 38688
rect 1332 38632 1358 38688
rect 1414 38632 1423 38688
rect 282 38602 1423 38632
rect 282 38546 291 38602
rect 347 38546 374 38602
rect 430 38546 456 38602
rect 512 38546 538 38602
rect 594 38546 620 38602
rect 676 38546 702 38602
rect 758 38546 784 38602
rect 840 38546 866 38602
rect 922 38546 948 38602
rect 1004 38546 1030 38602
rect 1086 38546 1112 38602
rect 1168 38546 1194 38602
rect 1250 38546 1276 38602
rect 1332 38546 1358 38602
rect 1414 38546 1423 38602
rect 282 38516 1423 38546
rect 282 38460 291 38516
rect 347 38460 374 38516
rect 430 38460 456 38516
rect 512 38460 538 38516
rect 594 38460 620 38516
rect 676 38460 702 38516
rect 758 38460 784 38516
rect 840 38460 866 38516
rect 922 38460 948 38516
rect 1004 38460 1030 38516
rect 1086 38460 1112 38516
rect 1168 38460 1194 38516
rect 1250 38460 1276 38516
rect 1332 38460 1358 38516
rect 1414 38460 1423 38516
rect 282 38430 1423 38460
rect 282 38374 291 38430
rect 347 38374 374 38430
rect 430 38374 456 38430
rect 512 38374 538 38430
rect 594 38374 620 38430
rect 676 38374 702 38430
rect 758 38374 784 38430
rect 840 38374 866 38430
rect 922 38374 948 38430
rect 1004 38374 1030 38430
rect 1086 38374 1112 38430
rect 1168 38374 1194 38430
rect 1250 38374 1276 38430
rect 1332 38374 1358 38430
rect 1414 38374 1423 38430
rect 282 38344 1423 38374
rect 282 38288 291 38344
rect 347 38288 374 38344
rect 430 38288 456 38344
rect 512 38288 538 38344
rect 594 38288 620 38344
rect 676 38288 702 38344
rect 758 38288 784 38344
rect 840 38288 866 38344
rect 922 38288 948 38344
rect 1004 38288 1030 38344
rect 1086 38288 1112 38344
rect 1168 38288 1194 38344
rect 1250 38288 1276 38344
rect 1332 38288 1358 38344
rect 1414 38288 1423 38344
rect 282 38258 1423 38288
rect 282 38202 291 38258
rect 347 38202 374 38258
rect 430 38202 456 38258
rect 512 38202 538 38258
rect 594 38202 620 38258
rect 676 38202 702 38258
rect 758 38202 784 38258
rect 840 38202 866 38258
rect 922 38202 948 38258
rect 1004 38202 1030 38258
rect 1086 38202 1112 38258
rect 1168 38202 1194 38258
rect 1250 38202 1276 38258
rect 1332 38202 1358 38258
rect 1414 38202 1423 38258
rect 282 38172 1423 38202
rect 282 38116 291 38172
rect 347 38116 374 38172
rect 430 38116 456 38172
rect 512 38116 538 38172
rect 594 38116 620 38172
rect 676 38116 702 38172
rect 758 38116 784 38172
rect 840 38116 866 38172
rect 922 38116 948 38172
rect 1004 38116 1030 38172
rect 1086 38116 1112 38172
rect 1168 38116 1194 38172
rect 1250 38116 1276 38172
rect 1332 38116 1358 38172
rect 1414 38116 1423 38172
rect 282 38086 1423 38116
rect 282 38030 291 38086
rect 347 38030 374 38086
rect 430 38030 456 38086
rect 512 38030 538 38086
rect 594 38030 620 38086
rect 676 38030 702 38086
rect 758 38030 784 38086
rect 840 38030 866 38086
rect 922 38030 948 38086
rect 1004 38030 1030 38086
rect 1086 38030 1112 38086
rect 1168 38030 1194 38086
rect 1250 38030 1276 38086
rect 1332 38030 1358 38086
rect 1414 38030 1423 38086
rect 282 11131 1423 38030
rect 282 11075 632 11131
rect 688 11075 713 11131
rect 769 11075 794 11131
rect 850 11075 875 11131
rect 931 11075 956 11131
rect 1012 11075 1037 11131
rect 1093 11075 1118 11131
rect 1174 11075 1198 11131
rect 1254 11075 1278 11131
rect 1334 11075 1358 11131
rect 1414 11075 1423 11131
rect 282 10841 1423 11075
rect 282 10785 632 10841
rect 688 10785 713 10841
rect 769 10785 794 10841
rect 850 10785 875 10841
rect 931 10785 956 10841
rect 1012 10785 1037 10841
rect 1093 10785 1118 10841
rect 1174 10785 1198 10841
rect 1254 10785 1278 10841
rect 1334 10785 1358 10841
rect 1414 10785 1423 10841
rect 282 10705 1423 10785
rect 282 10649 632 10705
rect 688 10649 713 10705
rect 769 10649 794 10705
rect 850 10649 875 10705
rect 931 10649 956 10705
rect 1012 10649 1037 10705
rect 1093 10649 1118 10705
rect 1174 10649 1198 10705
rect 1254 10649 1278 10705
rect 1334 10649 1358 10705
rect 1414 10649 1423 10705
rect 282 9813 1423 10649
rect 282 9757 632 9813
rect 688 9757 713 9813
rect 769 9757 794 9813
rect 850 9757 875 9813
rect 931 9757 956 9813
rect 1012 9757 1037 9813
rect 1093 9757 1118 9813
rect 1174 9757 1198 9813
rect 1254 9757 1278 9813
rect 1334 9757 1358 9813
rect 1414 9757 1423 9813
rect 282 8153 1423 9757
rect 282 8097 637 8153
rect 693 8097 718 8153
rect 774 8097 798 8153
rect 854 8097 878 8153
rect 934 8097 958 8153
rect 1014 8097 1038 8153
rect 1094 8097 1118 8153
rect 1174 8097 1198 8153
rect 1254 8097 1278 8153
rect 1334 8097 1358 8153
rect 1414 8097 1423 8153
rect 282 8027 1423 8097
rect 282 7971 637 8027
rect 693 7971 718 8027
rect 774 7971 798 8027
rect 854 7971 878 8027
rect 934 7971 958 8027
rect 1014 7971 1038 8027
rect 1094 7971 1118 8027
rect 1174 7971 1198 8027
rect 1254 7971 1278 8027
rect 1334 7971 1358 8027
rect 1414 7971 1423 8027
rect 282 7723 1423 7971
rect 282 7667 291 7723
rect 347 7667 374 7723
rect 430 7667 456 7723
rect 512 7667 538 7723
rect 594 7667 620 7723
rect 676 7667 702 7723
rect 758 7667 784 7723
rect 840 7667 866 7723
rect 922 7667 948 7723
rect 1004 7667 1030 7723
rect 1086 7667 1112 7723
rect 1168 7667 1194 7723
rect 1250 7667 1276 7723
rect 1332 7667 1358 7723
rect 1414 7667 1423 7723
rect 282 7637 1423 7667
rect 282 7581 291 7637
rect 347 7581 374 7637
rect 430 7581 456 7637
rect 512 7581 538 7637
rect 594 7581 620 7637
rect 676 7581 702 7637
rect 758 7581 784 7637
rect 840 7581 866 7637
rect 922 7581 948 7637
rect 1004 7581 1030 7637
rect 1086 7581 1112 7637
rect 1168 7581 1194 7637
rect 1250 7581 1276 7637
rect 1332 7581 1358 7637
rect 1414 7581 1423 7637
rect 282 7551 1423 7581
rect 282 7495 291 7551
rect 347 7495 374 7551
rect 430 7495 456 7551
rect 512 7495 538 7551
rect 594 7495 620 7551
rect 676 7495 702 7551
rect 758 7495 784 7551
rect 840 7495 866 7551
rect 922 7495 948 7551
rect 1004 7495 1030 7551
rect 1086 7495 1112 7551
rect 1168 7495 1194 7551
rect 1250 7495 1276 7551
rect 1332 7495 1358 7551
rect 1414 7495 1423 7551
rect 282 7465 1423 7495
rect 282 7409 291 7465
rect 347 7409 374 7465
rect 430 7409 456 7465
rect 512 7409 538 7465
rect 594 7409 620 7465
rect 676 7409 702 7465
rect 758 7409 784 7465
rect 840 7409 866 7465
rect 922 7409 948 7465
rect 1004 7409 1030 7465
rect 1086 7409 1112 7465
rect 1168 7409 1194 7465
rect 1250 7409 1276 7465
rect 1332 7409 1358 7465
rect 1414 7409 1423 7465
rect 282 7379 1423 7409
rect 282 7323 291 7379
rect 347 7323 374 7379
rect 430 7323 456 7379
rect 512 7323 538 7379
rect 594 7323 620 7379
rect 676 7323 702 7379
rect 758 7323 784 7379
rect 840 7323 866 7379
rect 922 7323 948 7379
rect 1004 7323 1030 7379
rect 1086 7323 1112 7379
rect 1168 7323 1194 7379
rect 1250 7323 1276 7379
rect 1332 7323 1358 7379
rect 1414 7323 1423 7379
rect 282 7293 1423 7323
rect 282 7237 291 7293
rect 347 7237 374 7293
rect 430 7237 456 7293
rect 512 7237 538 7293
rect 594 7237 620 7293
rect 676 7237 702 7293
rect 758 7237 784 7293
rect 840 7237 866 7293
rect 922 7237 948 7293
rect 1004 7237 1030 7293
rect 1086 7237 1112 7293
rect 1168 7237 1194 7293
rect 1250 7237 1276 7293
rect 1332 7237 1358 7293
rect 1414 7237 1423 7293
rect 282 7207 1423 7237
rect 282 7151 291 7207
rect 347 7151 374 7207
rect 430 7151 456 7207
rect 512 7151 538 7207
rect 594 7151 620 7207
rect 676 7151 702 7207
rect 758 7151 784 7207
rect 840 7151 866 7207
rect 922 7151 948 7207
rect 1004 7151 1030 7207
rect 1086 7151 1112 7207
rect 1168 7151 1194 7207
rect 1250 7151 1276 7207
rect 1332 7151 1358 7207
rect 1414 7151 1423 7207
rect 282 7121 1423 7151
rect 282 7065 291 7121
rect 347 7065 374 7121
rect 430 7065 456 7121
rect 512 7065 538 7121
rect 594 7065 620 7121
rect 676 7065 702 7121
rect 758 7065 784 7121
rect 840 7065 866 7121
rect 922 7065 948 7121
rect 1004 7065 1030 7121
rect 1086 7065 1112 7121
rect 1168 7065 1194 7121
rect 1250 7065 1276 7121
rect 1332 7065 1358 7121
rect 1414 7065 1423 7121
rect 282 7035 1423 7065
rect 282 6979 291 7035
rect 347 6979 374 7035
rect 430 6979 456 7035
rect 512 6979 538 7035
rect 594 6979 620 7035
rect 676 6979 702 7035
rect 758 6979 784 7035
rect 840 6979 866 7035
rect 922 6979 948 7035
rect 1004 6979 1030 7035
rect 1086 6979 1112 7035
rect 1168 6979 1194 7035
rect 1250 6979 1276 7035
rect 1332 6979 1358 7035
rect 1414 6979 1423 7035
rect 282 6949 1423 6979
rect 282 6893 291 6949
rect 347 6893 374 6949
rect 430 6893 456 6949
rect 512 6893 538 6949
rect 594 6893 620 6949
rect 676 6893 702 6949
rect 758 6893 784 6949
rect 840 6893 866 6949
rect 922 6893 948 6949
rect 1004 6893 1030 6949
rect 1086 6893 1112 6949
rect 1168 6893 1194 6949
rect 1250 6893 1276 6949
rect 1332 6893 1358 6949
rect 1414 6893 1423 6949
rect 282 6863 1423 6893
rect 282 6807 291 6863
rect 347 6807 374 6863
rect 430 6807 456 6863
rect 512 6807 538 6863
rect 594 6807 620 6863
rect 676 6807 702 6863
rect 758 6807 784 6863
rect 840 6807 866 6863
rect 922 6807 948 6863
rect 1004 6807 1030 6863
rect 1086 6807 1112 6863
rect 1168 6807 1194 6863
rect 1250 6807 1276 6863
rect 1332 6807 1358 6863
rect 1414 6807 1423 6863
rect 282 821 1423 6807
rect 1583 27485 2501 40000
rect 1583 27452 2468 27485
tri 2468 27452 2501 27485 nw
rect 2661 38979 3543 40000
rect 2661 38923 2714 38979
rect 2770 38923 2794 38979
rect 2850 38923 2874 38979
rect 2930 38923 2954 38979
rect 3010 38923 3034 38979
rect 3090 38923 3114 38979
rect 3170 38923 3194 38979
rect 3250 38923 3274 38979
rect 3330 38923 3354 38979
rect 3410 38923 3434 38979
rect 3490 38923 3543 38979
rect 2661 38895 3543 38923
rect 2661 38839 2714 38895
rect 2770 38839 2794 38895
rect 2850 38839 2874 38895
rect 2930 38839 2954 38895
rect 3010 38839 3034 38895
rect 3090 38839 3114 38895
rect 3170 38839 3194 38895
rect 3250 38839 3274 38895
rect 3330 38839 3354 38895
rect 3410 38839 3434 38895
rect 3490 38839 3543 38895
rect 2661 38811 3543 38839
rect 2661 38755 2714 38811
rect 2770 38755 2794 38811
rect 2850 38755 2874 38811
rect 2930 38755 2954 38811
rect 3010 38755 3034 38811
rect 3090 38755 3114 38811
rect 3170 38755 3194 38811
rect 3250 38755 3274 38811
rect 3330 38755 3354 38811
rect 3410 38755 3434 38811
rect 3490 38755 3543 38811
rect 2661 38727 3543 38755
rect 2661 38671 2714 38727
rect 2770 38671 2794 38727
rect 2850 38671 2874 38727
rect 2930 38671 2954 38727
rect 3010 38671 3034 38727
rect 3090 38671 3114 38727
rect 3170 38671 3194 38727
rect 3250 38671 3274 38727
rect 3330 38671 3354 38727
rect 3410 38671 3434 38727
rect 3490 38671 3543 38727
rect 2661 38643 3543 38671
rect 2661 38587 2714 38643
rect 2770 38587 2794 38643
rect 2850 38587 2874 38643
rect 2930 38587 2954 38643
rect 3010 38587 3034 38643
rect 3090 38587 3114 38643
rect 3170 38587 3194 38643
rect 3250 38587 3274 38643
rect 3330 38587 3354 38643
rect 3410 38587 3434 38643
rect 3490 38587 3543 38643
rect 2661 38559 3543 38587
rect 2661 38503 2714 38559
rect 2770 38503 2794 38559
rect 2850 38503 2874 38559
rect 2930 38503 2954 38559
rect 3010 38503 3034 38559
rect 3090 38503 3114 38559
rect 3170 38503 3194 38559
rect 3250 38503 3274 38559
rect 3330 38503 3354 38559
rect 3410 38503 3434 38559
rect 3490 38503 3543 38559
rect 2661 38475 3543 38503
rect 2661 38419 2714 38475
rect 2770 38419 2794 38475
rect 2850 38419 2874 38475
rect 2930 38419 2954 38475
rect 3010 38419 3034 38475
rect 3090 38419 3114 38475
rect 3170 38419 3194 38475
rect 3250 38419 3274 38475
rect 3330 38419 3354 38475
rect 3410 38419 3434 38475
rect 3490 38419 3543 38475
rect 2661 38391 3543 38419
rect 2661 38335 2714 38391
rect 2770 38335 2794 38391
rect 2850 38335 2874 38391
rect 2930 38335 2954 38391
rect 3010 38335 3034 38391
rect 3090 38335 3114 38391
rect 3170 38335 3194 38391
rect 3250 38335 3274 38391
rect 3330 38335 3354 38391
rect 3410 38335 3434 38391
rect 3490 38335 3543 38391
rect 2661 38307 3543 38335
rect 2661 38251 2714 38307
rect 2770 38251 2794 38307
rect 2850 38251 2874 38307
rect 2930 38251 2954 38307
rect 3010 38251 3034 38307
rect 3090 38251 3114 38307
rect 3170 38251 3194 38307
rect 3250 38251 3274 38307
rect 3330 38251 3354 38307
rect 3410 38251 3434 38307
rect 3490 38251 3543 38307
rect 2661 38223 3543 38251
rect 2661 38167 2714 38223
rect 2770 38167 2794 38223
rect 2850 38167 2874 38223
rect 2930 38167 2954 38223
rect 3010 38167 3034 38223
rect 3090 38167 3114 38223
rect 3170 38167 3194 38223
rect 3250 38167 3274 38223
rect 3330 38167 3354 38223
rect 3410 38167 3434 38223
rect 3490 38167 3543 38223
rect 2661 38138 3543 38167
rect 2661 38082 2714 38138
rect 2770 38082 2794 38138
rect 2850 38082 2874 38138
rect 2930 38082 2954 38138
rect 3010 38082 3034 38138
rect 3090 38082 3114 38138
rect 3170 38082 3194 38138
rect 3250 38082 3274 38138
rect 3330 38082 3354 38138
rect 3410 38082 3434 38138
rect 3490 38082 3543 38138
rect 2661 38053 3543 38082
rect 2661 37997 2714 38053
rect 2770 37997 2794 38053
rect 2850 37997 2874 38053
rect 2930 37997 2954 38053
rect 3010 37997 3034 38053
rect 3090 37997 3114 38053
rect 3170 37997 3194 38053
rect 3250 37997 3274 38053
rect 3330 37997 3354 38053
rect 3410 37997 3434 38053
rect 3490 37997 3543 38053
rect 2661 27992 3543 37997
rect 2661 27936 2670 27992
rect 2726 27936 2759 27992
rect 2815 27936 2848 27992
rect 2904 27936 2937 27992
rect 2993 27936 3025 27992
rect 3081 27936 3113 27992
rect 3169 27936 3201 27992
rect 3257 27936 3289 27992
rect 3345 27936 3377 27992
rect 3433 27936 3543 27992
rect 2661 27902 3543 27936
rect 2661 27846 2670 27902
rect 2726 27846 2759 27902
rect 2815 27846 2848 27902
rect 2904 27846 2937 27902
rect 2993 27846 3025 27902
rect 3081 27846 3113 27902
rect 3169 27846 3201 27902
rect 3257 27846 3289 27902
rect 3345 27846 3377 27902
rect 3433 27846 3543 27902
rect 2661 27812 3543 27846
rect 2661 27756 2670 27812
rect 2726 27756 2759 27812
rect 2815 27756 2848 27812
rect 2904 27756 2937 27812
rect 2993 27756 3025 27812
rect 3081 27756 3113 27812
rect 3169 27756 3201 27812
rect 3257 27756 3289 27812
rect 3345 27756 3377 27812
rect 3433 27756 3543 27812
rect 2661 27722 3543 27756
rect 2661 27666 2670 27722
rect 2726 27666 2759 27722
rect 2815 27666 2848 27722
rect 2904 27666 2937 27722
rect 2993 27666 3025 27722
rect 3081 27666 3113 27722
rect 3169 27666 3201 27722
rect 3257 27666 3289 27722
rect 3345 27666 3377 27722
rect 3433 27666 3543 27722
rect 2661 27632 3543 27666
rect 2661 27576 2670 27632
rect 2726 27576 2759 27632
rect 2815 27576 2848 27632
rect 2904 27576 2937 27632
rect 2993 27576 3025 27632
rect 3081 27576 3113 27632
rect 3169 27576 3201 27632
rect 3257 27576 3289 27632
rect 3345 27576 3377 27632
rect 3433 27576 3543 27632
rect 2661 27542 3543 27576
rect 2661 27486 2670 27542
rect 2726 27486 2759 27542
rect 2815 27486 2848 27542
rect 2904 27486 2937 27542
rect 2993 27486 3025 27542
rect 3081 27486 3113 27542
rect 3169 27486 3201 27542
rect 3257 27486 3289 27542
rect 3345 27486 3377 27542
rect 3433 27486 3543 27542
rect 2661 27452 3543 27486
rect 1583 27396 2412 27452
tri 2412 27396 2468 27452 nw
rect 2661 27396 2670 27452
rect 2726 27396 2759 27452
rect 2815 27396 2848 27452
rect 2904 27396 2937 27452
rect 2993 27396 3025 27452
rect 3081 27396 3113 27452
rect 3169 27396 3201 27452
rect 3257 27396 3289 27452
rect 3345 27396 3377 27452
rect 3433 27396 3543 27452
rect 282 0 1423 631
rect 1583 0 2383 27396
tri 2383 27367 2412 27396 nw
rect 2483 27327 2561 27336
rect 2483 27271 2494 27327
rect 2550 27271 2561 27327
rect 2483 27247 2561 27271
rect 2483 27191 2494 27247
rect 2550 27191 2561 27247
rect 2483 145 2561 27191
rect 2483 89 2494 145
rect 2550 89 2561 145
rect 2483 65 2561 89
rect 2483 9 2494 65
rect 2550 9 2561 65
rect 2483 0 2561 9
rect 2661 24523 3543 27396
rect 2661 24467 2670 24523
rect 2726 24467 2751 24523
rect 2807 24467 2832 24523
rect 2888 24467 2913 24523
rect 2969 24467 2994 24523
rect 3050 24467 3075 24523
rect 3131 24467 3156 24523
rect 3212 24467 3237 24523
rect 3293 24467 3318 24523
rect 3374 24467 3398 24523
rect 3454 24467 3478 24523
rect 3534 24467 3543 24523
rect 2661 24397 3543 24467
rect 2661 24341 2670 24397
rect 2726 24341 2751 24397
rect 2807 24341 2832 24397
rect 2888 24341 2913 24397
rect 2969 24341 2994 24397
rect 3050 24341 3075 24397
rect 3131 24341 3156 24397
rect 3212 24341 3237 24397
rect 3293 24341 3318 24397
rect 3374 24341 3398 24397
rect 3454 24341 3478 24397
rect 3534 24341 3543 24397
rect 2661 23268 3543 24341
rect 2661 23212 2670 23268
rect 2726 23212 2751 23268
rect 2807 23212 2832 23268
rect 2888 23212 2913 23268
rect 2969 23212 2994 23268
rect 3050 23212 3075 23268
rect 3131 23212 3156 23268
rect 3212 23212 3237 23268
rect 3293 23212 3318 23268
rect 3374 23212 3398 23268
rect 3454 23212 3478 23268
rect 3534 23212 3543 23268
rect 2661 23180 3543 23212
rect 2661 23124 2670 23180
rect 2726 23124 2751 23180
rect 2807 23124 2832 23180
rect 2888 23124 2913 23180
rect 2969 23124 2994 23180
rect 3050 23124 3075 23180
rect 3131 23124 3156 23180
rect 3212 23124 3237 23180
rect 3293 23124 3318 23180
rect 3374 23124 3398 23180
rect 3454 23124 3478 23180
rect 3534 23124 3543 23180
rect 2661 23092 3543 23124
rect 2661 23036 2670 23092
rect 2726 23036 2751 23092
rect 2807 23036 2832 23092
rect 2888 23036 2913 23092
rect 2969 23036 2994 23092
rect 3050 23036 3075 23092
rect 3131 23036 3156 23092
rect 3212 23036 3237 23092
rect 3293 23036 3318 23092
rect 3374 23036 3398 23092
rect 3454 23036 3478 23092
rect 3534 23036 3543 23092
rect 2661 23004 3543 23036
rect 2661 22948 2670 23004
rect 2726 22948 2751 23004
rect 2807 22948 2832 23004
rect 2888 22948 2913 23004
rect 2969 22948 2994 23004
rect 3050 22948 3075 23004
rect 3131 22948 3156 23004
rect 3212 22948 3237 23004
rect 3293 22948 3318 23004
rect 3374 22948 3398 23004
rect 3454 22948 3478 23004
rect 3534 22948 3543 23004
rect 2661 22916 3543 22948
rect 2661 22860 2670 22916
rect 2726 22860 2751 22916
rect 2807 22860 2832 22916
rect 2888 22860 2913 22916
rect 2969 22860 2994 22916
rect 3050 22860 3075 22916
rect 3131 22860 3156 22916
rect 3212 22860 3237 22916
rect 3293 22860 3318 22916
rect 3374 22860 3398 22916
rect 3454 22860 3478 22916
rect 3534 22860 3543 22916
rect 2661 14611 3543 22860
rect 2661 14555 2670 14611
rect 2726 14555 2751 14611
rect 2807 14555 2832 14611
rect 2888 14555 2913 14611
rect 2969 14555 2994 14611
rect 3050 14555 3075 14611
rect 3131 14555 3156 14611
rect 3212 14555 3237 14611
rect 3293 14555 3318 14611
rect 3374 14555 3398 14611
rect 3454 14555 3478 14611
rect 3534 14555 3543 14611
rect 2661 14527 3543 14555
rect 2661 14471 2670 14527
rect 2726 14471 2751 14527
rect 2807 14471 2832 14527
rect 2888 14471 2913 14527
rect 2969 14471 2994 14527
rect 3050 14471 3075 14527
rect 3131 14471 3156 14527
rect 3212 14471 3237 14527
rect 3293 14471 3318 14527
rect 3374 14471 3398 14527
rect 3454 14471 3478 14527
rect 3534 14471 3543 14527
rect 2661 14443 3543 14471
rect 2661 14387 2670 14443
rect 2726 14387 2751 14443
rect 2807 14387 2832 14443
rect 2888 14387 2913 14443
rect 2969 14387 2994 14443
rect 3050 14387 3075 14443
rect 3131 14387 3156 14443
rect 3212 14387 3237 14443
rect 3293 14387 3318 14443
rect 3374 14387 3398 14443
rect 3454 14387 3478 14443
rect 3534 14387 3543 14443
rect 2661 11697 3543 14387
rect 2661 11641 2670 11697
rect 2726 11641 2751 11697
rect 2807 11641 2832 11697
rect 2888 11641 2913 11697
rect 2969 11641 2994 11697
rect 3050 11641 3075 11697
rect 3131 11641 3156 11697
rect 3212 11641 3237 11697
rect 3293 11641 3318 11697
rect 3374 11641 3398 11697
rect 3454 11641 3478 11697
rect 3534 11641 3543 11697
rect 2661 11615 3543 11641
rect 2661 11559 2670 11615
rect 2726 11559 2751 11615
rect 2807 11559 2832 11615
rect 2888 11559 2913 11615
rect 2969 11559 2994 11615
rect 3050 11559 3075 11615
rect 3131 11559 3156 11615
rect 3212 11559 3237 11615
rect 3293 11559 3318 11615
rect 3374 11559 3398 11615
rect 3454 11559 3478 11615
rect 3534 11559 3543 11615
rect 2661 7756 3543 11559
rect 2661 7700 2714 7756
rect 2770 7700 2794 7756
rect 2850 7700 2874 7756
rect 2930 7700 2954 7756
rect 3010 7700 3034 7756
rect 3090 7700 3114 7756
rect 3170 7700 3194 7756
rect 3250 7700 3274 7756
rect 3330 7700 3354 7756
rect 3410 7700 3434 7756
rect 3490 7700 3543 7756
rect 2661 7672 3543 7700
rect 2661 7616 2714 7672
rect 2770 7616 2794 7672
rect 2850 7616 2874 7672
rect 2930 7616 2954 7672
rect 3010 7616 3034 7672
rect 3090 7616 3114 7672
rect 3170 7616 3194 7672
rect 3250 7616 3274 7672
rect 3330 7616 3354 7672
rect 3410 7616 3434 7672
rect 3490 7616 3543 7672
rect 2661 7588 3543 7616
rect 2661 7532 2714 7588
rect 2770 7532 2794 7588
rect 2850 7532 2874 7588
rect 2930 7532 2954 7588
rect 3010 7532 3034 7588
rect 3090 7532 3114 7588
rect 3170 7532 3194 7588
rect 3250 7532 3274 7588
rect 3330 7532 3354 7588
rect 3410 7532 3434 7588
rect 3490 7532 3543 7588
rect 2661 7504 3543 7532
rect 2661 7448 2714 7504
rect 2770 7448 2794 7504
rect 2850 7448 2874 7504
rect 2930 7448 2954 7504
rect 3010 7448 3034 7504
rect 3090 7448 3114 7504
rect 3170 7448 3194 7504
rect 3250 7448 3274 7504
rect 3330 7448 3354 7504
rect 3410 7448 3434 7504
rect 3490 7448 3543 7504
rect 2661 7420 3543 7448
rect 2661 7364 2714 7420
rect 2770 7364 2794 7420
rect 2850 7364 2874 7420
rect 2930 7364 2954 7420
rect 3010 7364 3034 7420
rect 3090 7364 3114 7420
rect 3170 7364 3194 7420
rect 3250 7364 3274 7420
rect 3330 7364 3354 7420
rect 3410 7364 3434 7420
rect 3490 7364 3543 7420
rect 2661 7336 3543 7364
rect 2661 7280 2714 7336
rect 2770 7280 2794 7336
rect 2850 7280 2874 7336
rect 2930 7280 2954 7336
rect 3010 7280 3034 7336
rect 3090 7280 3114 7336
rect 3170 7280 3194 7336
rect 3250 7280 3274 7336
rect 3330 7280 3354 7336
rect 3410 7280 3434 7336
rect 3490 7280 3543 7336
rect 2661 7252 3543 7280
rect 2661 7196 2714 7252
rect 2770 7196 2794 7252
rect 2850 7196 2874 7252
rect 2930 7196 2954 7252
rect 3010 7196 3034 7252
rect 3090 7196 3114 7252
rect 3170 7196 3194 7252
rect 3250 7196 3274 7252
rect 3330 7196 3354 7252
rect 3410 7196 3434 7252
rect 3490 7196 3543 7252
rect 2661 7168 3543 7196
rect 2661 7112 2714 7168
rect 2770 7112 2794 7168
rect 2850 7112 2874 7168
rect 2930 7112 2954 7168
rect 3010 7112 3034 7168
rect 3090 7112 3114 7168
rect 3170 7112 3194 7168
rect 3250 7112 3274 7168
rect 3330 7112 3354 7168
rect 3410 7112 3434 7168
rect 3490 7112 3543 7168
rect 2661 7084 3543 7112
rect 2661 7028 2714 7084
rect 2770 7028 2794 7084
rect 2850 7028 2874 7084
rect 2930 7028 2954 7084
rect 3010 7028 3034 7084
rect 3090 7028 3114 7084
rect 3170 7028 3194 7084
rect 3250 7028 3274 7084
rect 3330 7028 3354 7084
rect 3410 7028 3434 7084
rect 3490 7028 3543 7084
rect 2661 7000 3543 7028
rect 2661 6944 2714 7000
rect 2770 6944 2794 7000
rect 2850 6944 2874 7000
rect 2930 6944 2954 7000
rect 3010 6944 3034 7000
rect 3090 6944 3114 7000
rect 3170 6944 3194 7000
rect 3250 6944 3274 7000
rect 3330 6944 3354 7000
rect 3410 6944 3434 7000
rect 3490 6944 3543 7000
rect 2661 6915 3543 6944
rect 2661 6859 2714 6915
rect 2770 6859 2794 6915
rect 2850 6859 2874 6915
rect 2930 6859 2954 6915
rect 3010 6859 3034 6915
rect 3090 6859 3114 6915
rect 3170 6859 3194 6915
rect 3250 6859 3274 6915
rect 3330 6859 3354 6915
rect 3410 6859 3434 6915
rect 3490 6859 3543 6915
rect 2661 6830 3543 6859
rect 2661 6774 2714 6830
rect 2770 6774 2794 6830
rect 2850 6774 2874 6830
rect 2930 6774 2954 6830
rect 3010 6774 3034 6830
rect 3090 6774 3114 6830
rect 3170 6774 3194 6830
rect 3250 6774 3274 6830
rect 3330 6774 3354 6830
rect 3410 6774 3434 6830
rect 3490 6774 3543 6830
rect 2661 0 3543 6774
rect 3703 21158 4503 40000
rect 3703 21102 3712 21158
rect 3768 21102 3793 21158
rect 3849 21102 3874 21158
rect 3930 21102 3955 21158
rect 4011 21102 4036 21158
rect 4092 21102 4117 21158
rect 4173 21102 4198 21158
rect 4254 21102 4278 21158
rect 4334 21102 4358 21158
rect 4414 21102 4438 21158
rect 4494 21102 4503 21158
rect 3703 21072 4503 21102
rect 3703 21016 3712 21072
rect 3768 21016 3793 21072
rect 3849 21016 3874 21072
rect 3930 21016 3955 21072
rect 4011 21016 4036 21072
rect 4092 21016 4117 21072
rect 4173 21016 4198 21072
rect 4254 21016 4278 21072
rect 4334 21016 4358 21072
rect 4414 21016 4438 21072
rect 4494 21016 4503 21072
rect 3703 20986 4503 21016
rect 3703 20930 3712 20986
rect 3768 20930 3793 20986
rect 3849 20930 3874 20986
rect 3930 20930 3955 20986
rect 4011 20930 4036 20986
rect 4092 20930 4117 20986
rect 4173 20930 4198 20986
rect 4254 20930 4278 20986
rect 4334 20930 4358 20986
rect 4414 20930 4438 20986
rect 4494 20930 4503 20986
rect 3703 20900 4503 20930
rect 3703 20844 3712 20900
rect 3768 20844 3793 20900
rect 3849 20844 3874 20900
rect 3930 20844 3955 20900
rect 4011 20844 4036 20900
rect 4092 20844 4117 20900
rect 4173 20844 4198 20900
rect 4254 20844 4278 20900
rect 4334 20844 4358 20900
rect 4414 20844 4438 20900
rect 4494 20844 4503 20900
rect 3703 20814 4503 20844
rect 3703 20758 3712 20814
rect 3768 20758 3793 20814
rect 3849 20758 3874 20814
rect 3930 20758 3955 20814
rect 4011 20758 4036 20814
rect 4092 20758 4117 20814
rect 4173 20758 4198 20814
rect 4254 20758 4278 20814
rect 4334 20758 4358 20814
rect 4414 20758 4438 20814
rect 4494 20758 4503 20814
rect 3703 19095 4503 20758
rect 3703 19039 3712 19095
rect 3768 19039 3793 19095
rect 3849 19039 3874 19095
rect 3930 19039 3955 19095
rect 4011 19039 4036 19095
rect 4092 19039 4117 19095
rect 4173 19039 4198 19095
rect 4254 19039 4278 19095
rect 4334 19039 4358 19095
rect 4414 19039 4438 19095
rect 4494 19039 4503 19095
rect 3703 18951 4503 19039
rect 3703 18895 3712 18951
rect 3768 18895 3793 18951
rect 3849 18895 3874 18951
rect 3930 18895 3955 18951
rect 4011 18895 4036 18951
rect 4092 18895 4117 18951
rect 4173 18895 4198 18951
rect 4254 18895 4278 18951
rect 4334 18895 4358 18951
rect 4414 18895 4438 18951
rect 4494 18895 4503 18951
rect 3703 17336 4503 18895
rect 3703 17280 3712 17336
rect 3768 17280 3793 17336
rect 3849 17280 3874 17336
rect 3930 17280 3955 17336
rect 4011 17280 4036 17336
rect 4092 17280 4117 17336
rect 4173 17280 4198 17336
rect 4254 17280 4278 17336
rect 4334 17280 4358 17336
rect 4414 17280 4438 17336
rect 4494 17280 4503 17336
rect 3703 17250 4503 17280
rect 3703 17194 3712 17250
rect 3768 17194 3793 17250
rect 3849 17194 3874 17250
rect 3930 17194 3955 17250
rect 4011 17194 4036 17250
rect 4092 17194 4117 17250
rect 4173 17194 4198 17250
rect 4254 17194 4278 17250
rect 4334 17194 4358 17250
rect 4414 17194 4438 17250
rect 4494 17194 4503 17250
rect 3703 17164 4503 17194
rect 3703 17108 3712 17164
rect 3768 17108 3793 17164
rect 3849 17108 3874 17164
rect 3930 17108 3955 17164
rect 4011 17108 4036 17164
rect 4092 17108 4117 17164
rect 4173 17108 4198 17164
rect 4254 17108 4278 17164
rect 4334 17108 4358 17164
rect 4414 17108 4438 17164
rect 4494 17108 4503 17164
rect 3703 17078 4503 17108
rect 3703 17022 3712 17078
rect 3768 17022 3793 17078
rect 3849 17022 3874 17078
rect 3930 17022 3955 17078
rect 4011 17022 4036 17078
rect 4092 17022 4117 17078
rect 4173 17022 4198 17078
rect 4254 17022 4278 17078
rect 4334 17022 4358 17078
rect 4414 17022 4438 17078
rect 4494 17022 4503 17078
rect 3703 16992 4503 17022
rect 3703 16936 3712 16992
rect 3768 16936 3793 16992
rect 3849 16936 3874 16992
rect 3930 16936 3955 16992
rect 4011 16936 4036 16992
rect 4092 16936 4117 16992
rect 4173 16936 4198 16992
rect 4254 16936 4278 16992
rect 4334 16936 4358 16992
rect 4414 16936 4438 16992
rect 4494 16936 4503 16992
rect 3703 15221 4503 16936
rect 3703 15165 3712 15221
rect 3768 15165 3793 15221
rect 3849 15165 3874 15221
rect 3930 15165 3955 15221
rect 4011 15165 4036 15221
rect 4092 15165 4117 15221
rect 4173 15165 4198 15221
rect 3703 15141 4198 15165
rect 3703 15085 3712 15141
rect 3768 15085 3793 15141
rect 3849 15085 3874 15141
rect 3930 15085 3955 15141
rect 4011 15085 4036 15141
rect 4092 15085 4117 15141
rect 4173 15085 4198 15141
rect 3703 15061 4198 15085
rect 3703 15005 3712 15061
rect 3768 15005 3793 15061
rect 3849 15005 3874 15061
rect 3930 15005 3955 15061
rect 4011 15005 4036 15061
rect 4092 15005 4117 15061
rect 4173 15005 4198 15061
rect 3703 14981 4198 15005
rect 3703 14925 3712 14981
rect 3768 14925 3793 14981
rect 3849 14925 3874 14981
rect 3930 14925 3955 14981
rect 4011 14925 4036 14981
rect 4092 14925 4117 14981
rect 4173 14925 4198 14981
rect 4494 14925 4503 15221
rect 3703 1516 4503 14925
rect 3703 1460 3712 1516
rect 3768 1460 3798 1516
rect 3854 1460 3884 1516
rect 3940 1460 3970 1516
rect 4026 1460 4056 1516
rect 4112 1460 4142 1516
rect 4198 1460 4228 1516
rect 4284 1460 4314 1516
rect 4370 1460 4399 1516
rect 4455 1460 4503 1516
rect 3703 1432 4503 1460
rect 3703 1376 3712 1432
rect 3768 1376 3798 1432
rect 3854 1376 3884 1432
rect 3940 1376 3970 1432
rect 4026 1376 4056 1432
rect 4112 1376 4142 1432
rect 4198 1376 4228 1432
rect 4284 1376 4314 1432
rect 4370 1376 4399 1432
rect 4455 1376 4503 1432
rect 3703 1348 4503 1376
rect 3703 1292 3712 1348
rect 3768 1292 3798 1348
rect 3854 1292 3884 1348
rect 3940 1292 3970 1348
rect 4026 1292 4056 1348
rect 4112 1292 4142 1348
rect 4198 1292 4228 1348
rect 4284 1292 4314 1348
rect 4370 1292 4399 1348
rect 4455 1292 4503 1348
rect 3703 1264 4503 1292
rect 3703 1208 3712 1264
rect 3768 1208 3798 1264
rect 3854 1208 3884 1264
rect 3940 1208 3970 1264
rect 4026 1208 4056 1264
rect 4112 1208 4142 1264
rect 4198 1208 4228 1264
rect 4284 1208 4314 1264
rect 4370 1208 4399 1264
rect 4455 1208 4503 1264
rect 3703 0 4503 1208
rect 4663 0 5663 40000
rect 5823 18262 6623 40000
rect 5823 18206 5832 18262
rect 5888 18206 5914 18262
rect 5970 18206 5995 18262
rect 6051 18206 6076 18262
rect 6132 18206 6157 18262
rect 6213 18206 6238 18262
rect 6294 18206 6319 18262
rect 6375 18206 6400 18262
rect 6456 18206 6481 18262
rect 6537 18206 6562 18262
rect 6618 18206 6623 18262
rect 5823 18182 6623 18206
rect 5823 18126 5832 18182
rect 5888 18126 5914 18182
rect 5970 18126 5995 18182
rect 6051 18126 6076 18182
rect 6132 18126 6157 18182
rect 6213 18126 6238 18182
rect 6294 18126 6319 18182
rect 6375 18126 6400 18182
rect 6456 18126 6481 18182
rect 6537 18126 6562 18182
rect 6618 18126 6623 18182
rect 5823 7937 6623 18126
rect 6733 26852 7908 40000
rect 6733 26796 6742 26852
rect 6798 26796 6827 26852
rect 6883 26796 6912 26852
rect 6968 26796 6997 26852
rect 7053 26796 7082 26852
rect 7138 26796 7167 26852
rect 7223 26796 7252 26852
rect 7308 26796 7337 26852
rect 7393 26796 7422 26852
rect 7478 26796 7507 26852
rect 7563 26796 7591 26852
rect 7647 26796 7675 26852
rect 7731 26796 7759 26852
rect 7815 26796 7843 26852
rect 7899 26796 7908 26852
rect 6733 26766 7908 26796
rect 6733 26710 6742 26766
rect 6798 26710 6827 26766
rect 6883 26710 6912 26766
rect 6968 26710 6997 26766
rect 7053 26710 7082 26766
rect 7138 26710 7167 26766
rect 7223 26710 7252 26766
rect 7308 26710 7337 26766
rect 7393 26710 7422 26766
rect 7478 26710 7507 26766
rect 7563 26710 7591 26766
rect 7647 26710 7675 26766
rect 7731 26710 7759 26766
rect 7815 26710 7843 26766
rect 7899 26710 7908 26766
rect 6733 26680 7908 26710
rect 6733 26624 6742 26680
rect 6798 26624 6827 26680
rect 6883 26624 6912 26680
rect 6968 26624 6997 26680
rect 7053 26624 7082 26680
rect 7138 26624 7167 26680
rect 7223 26624 7252 26680
rect 7308 26624 7337 26680
rect 7393 26624 7422 26680
rect 7478 26624 7507 26680
rect 7563 26624 7591 26680
rect 7647 26624 7675 26680
rect 7731 26624 7759 26680
rect 7815 26624 7843 26680
rect 7899 26624 7908 26680
rect 6733 26594 7908 26624
rect 6733 26538 6742 26594
rect 6798 26538 6827 26594
rect 6883 26538 6912 26594
rect 6968 26538 6997 26594
rect 7053 26538 7082 26594
rect 7138 26538 7167 26594
rect 7223 26538 7252 26594
rect 7308 26538 7337 26594
rect 7393 26538 7422 26594
rect 7478 26538 7507 26594
rect 7563 26538 7591 26594
rect 7647 26538 7675 26594
rect 7731 26538 7759 26594
rect 7815 26538 7843 26594
rect 7899 26538 7908 26594
rect 6733 26508 7908 26538
rect 6733 26452 6742 26508
rect 6798 26452 6827 26508
rect 6883 26452 6912 26508
rect 6968 26452 6997 26508
rect 7053 26452 7082 26508
rect 7138 26452 7167 26508
rect 7223 26452 7252 26508
rect 7308 26452 7337 26508
rect 7393 26452 7422 26508
rect 7478 26452 7507 26508
rect 7563 26452 7591 26508
rect 7647 26452 7675 26508
rect 7731 26452 7759 26508
rect 7815 26452 7843 26508
rect 7899 26452 7908 26508
rect 6733 12993 7908 26452
tri 6733 12726 7000 12993 ne
rect 6774 12625 6920 12630
rect 6774 12569 6779 12625
rect 6835 12569 6859 12625
rect 6915 12569 6920 12625
rect 6774 12095 6920 12569
rect 6774 12039 6779 12095
rect 6835 12039 6859 12095
rect 6915 12039 6920 12095
rect 6774 12034 6920 12039
rect 7000 12011 7908 12993
rect 7000 11622 7826 12011
tri 7826 11929 7908 12011 nw
rect 8026 36330 10856 40000
rect 8026 36274 8035 36330
rect 8091 36274 8116 36330
rect 8172 36274 8197 36330
rect 8253 36274 8277 36330
rect 8333 36274 8357 36330
rect 8413 36274 8437 36330
rect 8493 36274 8517 36330
rect 8573 36274 8597 36330
rect 8653 36274 8677 36330
rect 8733 36274 8757 36330
rect 8813 36274 8837 36330
rect 8893 36274 8917 36330
rect 8973 36274 8997 36330
rect 9053 36274 9077 36330
rect 9133 36274 9157 36330
rect 9213 36274 9237 36330
rect 9293 36274 9317 36330
rect 9373 36274 9397 36330
rect 9453 36274 9477 36330
rect 9533 36274 9557 36330
rect 9613 36274 9637 36330
rect 9693 36274 9717 36330
rect 9773 36274 9797 36330
rect 9853 36274 9877 36330
rect 9933 36274 9957 36330
rect 10013 36274 10856 36330
rect 8026 36244 10856 36274
rect 8026 36188 8035 36244
rect 8091 36188 8116 36244
rect 8172 36188 8197 36244
rect 8253 36188 8277 36244
rect 8333 36188 8357 36244
rect 8413 36188 8437 36244
rect 8493 36188 8517 36244
rect 8573 36188 8597 36244
rect 8653 36188 8677 36244
rect 8733 36188 8757 36244
rect 8813 36188 8837 36244
rect 8893 36188 8917 36244
rect 8973 36188 8997 36244
rect 9053 36188 9077 36244
rect 9133 36188 9157 36244
rect 9213 36188 9237 36244
rect 9293 36188 9317 36244
rect 9373 36188 9397 36244
rect 9453 36188 9477 36244
rect 9533 36188 9557 36244
rect 9613 36188 9637 36244
rect 9693 36188 9717 36244
rect 9773 36188 9797 36244
rect 9853 36188 9877 36244
rect 9933 36188 9957 36244
rect 10013 36188 10856 36244
rect 8026 36158 10856 36188
rect 8026 36102 8035 36158
rect 8091 36102 8116 36158
rect 8172 36102 8197 36158
rect 8253 36102 8277 36158
rect 8333 36102 8357 36158
rect 8413 36102 8437 36158
rect 8493 36102 8517 36158
rect 8573 36102 8597 36158
rect 8653 36102 8677 36158
rect 8733 36102 8757 36158
rect 8813 36102 8837 36158
rect 8893 36102 8917 36158
rect 8973 36102 8997 36158
rect 9053 36102 9077 36158
rect 9133 36102 9157 36158
rect 9213 36102 9237 36158
rect 9293 36102 9317 36158
rect 9373 36102 9397 36158
rect 9453 36102 9477 36158
rect 9533 36102 9557 36158
rect 9613 36102 9637 36158
rect 9693 36102 9717 36158
rect 9773 36102 9797 36158
rect 9853 36102 9877 36158
rect 9933 36102 9957 36158
rect 10013 36102 10856 36158
rect 8026 36072 10856 36102
rect 8026 36016 8035 36072
rect 8091 36016 8116 36072
rect 8172 36016 8197 36072
rect 8253 36016 8277 36072
rect 8333 36016 8357 36072
rect 8413 36016 8437 36072
rect 8493 36016 8517 36072
rect 8573 36016 8597 36072
rect 8653 36016 8677 36072
rect 8733 36016 8757 36072
rect 8813 36016 8837 36072
rect 8893 36016 8917 36072
rect 8973 36016 8997 36072
rect 9053 36016 9077 36072
rect 9133 36016 9157 36072
rect 9213 36016 9237 36072
rect 9293 36016 9317 36072
rect 9373 36016 9397 36072
rect 9453 36016 9477 36072
rect 9533 36016 9557 36072
rect 9613 36016 9637 36072
rect 9693 36016 9717 36072
rect 9773 36016 9797 36072
rect 9853 36016 9877 36072
rect 9933 36016 9957 36072
rect 10013 36016 10856 36072
rect 8026 35986 10856 36016
rect 8026 35930 8035 35986
rect 8091 35930 8116 35986
rect 8172 35930 8197 35986
rect 8253 35930 8277 35986
rect 8333 35930 8357 35986
rect 8413 35930 8437 35986
rect 8493 35930 8517 35986
rect 8573 35930 8597 35986
rect 8653 35930 8677 35986
rect 8733 35930 8757 35986
rect 8813 35930 8837 35986
rect 8893 35930 8917 35986
rect 8973 35930 8997 35986
rect 9053 35930 9077 35986
rect 9133 35930 9157 35986
rect 9213 35930 9237 35986
rect 9293 35930 9317 35986
rect 9373 35930 9397 35986
rect 9453 35930 9477 35986
rect 9533 35930 9557 35986
rect 9613 35930 9637 35986
rect 9693 35930 9717 35986
rect 9773 35930 9797 35986
rect 9853 35930 9877 35986
rect 9933 35930 9957 35986
rect 10013 35930 10856 35986
rect 8026 35900 10856 35930
rect 8026 35844 8035 35900
rect 8091 35844 8116 35900
rect 8172 35844 8197 35900
rect 8253 35844 8277 35900
rect 8333 35844 8357 35900
rect 8413 35844 8437 35900
rect 8493 35844 8517 35900
rect 8573 35844 8597 35900
rect 8653 35844 8677 35900
rect 8733 35844 8757 35900
rect 8813 35844 8837 35900
rect 8893 35844 8917 35900
rect 8973 35844 8997 35900
rect 9053 35844 9077 35900
rect 9133 35844 9157 35900
rect 9213 35844 9237 35900
rect 9293 35844 9317 35900
rect 9373 35844 9397 35900
rect 9453 35844 9477 35900
rect 9533 35844 9557 35900
rect 9613 35844 9637 35900
rect 9693 35844 9717 35900
rect 9773 35844 9797 35900
rect 9853 35844 9877 35900
rect 9933 35844 9957 35900
rect 10013 35844 10856 35900
rect 8026 35814 10856 35844
rect 8026 35758 8035 35814
rect 8091 35758 8116 35814
rect 8172 35758 8197 35814
rect 8253 35758 8277 35814
rect 8333 35758 8357 35814
rect 8413 35758 8437 35814
rect 8493 35758 8517 35814
rect 8573 35758 8597 35814
rect 8653 35758 8677 35814
rect 8733 35758 8757 35814
rect 8813 35758 8837 35814
rect 8893 35758 8917 35814
rect 8973 35758 8997 35814
rect 9053 35758 9077 35814
rect 9133 35758 9157 35814
rect 9213 35758 9237 35814
rect 9293 35758 9317 35814
rect 9373 35758 9397 35814
rect 9453 35758 9477 35814
rect 9533 35758 9557 35814
rect 9613 35758 9637 35814
rect 9693 35758 9717 35814
rect 9773 35758 9797 35814
rect 9853 35758 9877 35814
rect 9933 35758 9957 35814
rect 10013 35758 10856 35814
rect 8026 35728 10856 35758
rect 8026 35672 8035 35728
rect 8091 35672 8116 35728
rect 8172 35672 8197 35728
rect 8253 35672 8277 35728
rect 8333 35672 8357 35728
rect 8413 35672 8437 35728
rect 8493 35672 8517 35728
rect 8573 35672 8597 35728
rect 8653 35672 8677 35728
rect 8733 35672 8757 35728
rect 8813 35672 8837 35728
rect 8893 35672 8917 35728
rect 8973 35672 8997 35728
rect 9053 35672 9077 35728
rect 9133 35672 9157 35728
rect 9213 35672 9237 35728
rect 9293 35672 9317 35728
rect 9373 35672 9397 35728
rect 9453 35672 9477 35728
rect 9533 35672 9557 35728
rect 9613 35672 9637 35728
rect 9693 35672 9717 35728
rect 9773 35672 9797 35728
rect 9853 35672 9877 35728
rect 9933 35672 9957 35728
rect 10013 35672 10856 35728
rect 8026 35642 10856 35672
rect 8026 35586 8035 35642
rect 8091 35586 8116 35642
rect 8172 35586 8197 35642
rect 8253 35586 8277 35642
rect 8333 35586 8357 35642
rect 8413 35586 8437 35642
rect 8493 35586 8517 35642
rect 8573 35586 8597 35642
rect 8653 35586 8677 35642
rect 8733 35586 8757 35642
rect 8813 35586 8837 35642
rect 8893 35586 8917 35642
rect 8973 35586 8997 35642
rect 9053 35586 9077 35642
rect 9133 35586 9157 35642
rect 9213 35586 9237 35642
rect 9293 35586 9317 35642
rect 9373 35586 9397 35642
rect 9453 35586 9477 35642
rect 9533 35586 9557 35642
rect 9613 35586 9637 35642
rect 9693 35586 9717 35642
rect 9773 35586 9797 35642
rect 9853 35586 9877 35642
rect 9933 35586 9957 35642
rect 10013 35586 10856 35642
rect 8026 35556 10856 35586
rect 8026 35500 8035 35556
rect 8091 35500 8116 35556
rect 8172 35500 8197 35556
rect 8253 35500 8277 35556
rect 8333 35500 8357 35556
rect 8413 35500 8437 35556
rect 8493 35500 8517 35556
rect 8573 35500 8597 35556
rect 8653 35500 8677 35556
rect 8733 35500 8757 35556
rect 8813 35500 8837 35556
rect 8893 35500 8917 35556
rect 8973 35500 8997 35556
rect 9053 35500 9077 35556
rect 9133 35500 9157 35556
rect 9213 35500 9237 35556
rect 9293 35500 9317 35556
rect 9373 35500 9397 35556
rect 9453 35500 9477 35556
rect 9533 35500 9557 35556
rect 9613 35500 9637 35556
rect 9693 35500 9717 35556
rect 9773 35500 9797 35556
rect 9853 35500 9877 35556
rect 9933 35500 9957 35556
rect 10013 35500 10856 35556
rect 8026 35470 10856 35500
rect 8026 35414 8035 35470
rect 8091 35414 8116 35470
rect 8172 35414 8197 35470
rect 8253 35414 8277 35470
rect 8333 35414 8357 35470
rect 8413 35414 8437 35470
rect 8493 35414 8517 35470
rect 8573 35414 8597 35470
rect 8653 35414 8677 35470
rect 8733 35414 8757 35470
rect 8813 35414 8837 35470
rect 8893 35414 8917 35470
rect 8973 35414 8997 35470
rect 9053 35414 9077 35470
rect 9133 35414 9157 35470
rect 9213 35414 9237 35470
rect 9293 35414 9317 35470
rect 9373 35414 9397 35470
rect 9453 35414 9477 35470
rect 9533 35414 9557 35470
rect 9613 35414 9637 35470
rect 9693 35414 9717 35470
rect 9773 35414 9797 35470
rect 9853 35414 9877 35470
rect 9933 35414 9957 35470
rect 10013 35414 10856 35470
rect 8026 30338 10856 35414
rect 8026 30282 8490 30338
rect 8546 30282 8570 30338
rect 8626 30282 10856 30338
rect 8026 29462 10856 30282
rect 8026 29406 8490 29462
rect 8546 29406 8570 29462
rect 8626 29406 10856 29462
rect 8026 28927 10856 29406
rect 8026 28871 8035 28927
rect 8091 28871 8116 28927
rect 8172 28871 8197 28927
rect 8253 28871 8277 28927
rect 8333 28871 8357 28927
rect 8413 28871 8437 28927
rect 8493 28871 8517 28927
rect 8573 28871 8597 28927
rect 8653 28871 8677 28927
rect 8733 28871 8757 28927
rect 8813 28871 8837 28927
rect 8893 28871 8917 28927
rect 8973 28871 8997 28927
rect 9053 28871 9077 28927
rect 9133 28871 9157 28927
rect 9213 28871 9237 28927
rect 9293 28871 9317 28927
rect 9373 28871 9397 28927
rect 9453 28871 9477 28927
rect 9533 28871 9557 28927
rect 9613 28871 9637 28927
rect 9693 28871 9717 28927
rect 9773 28871 9797 28927
rect 9853 28871 9877 28927
rect 9933 28871 9957 28927
rect 10013 28871 10856 28927
rect 8026 28815 10856 28871
rect 8026 28759 8035 28815
rect 8091 28759 8116 28815
rect 8172 28759 8197 28815
rect 8253 28759 8277 28815
rect 8333 28759 8357 28815
rect 8413 28759 8437 28815
rect 8493 28759 8517 28815
rect 8573 28759 8597 28815
rect 8653 28759 8677 28815
rect 8733 28759 8757 28815
rect 8813 28759 8837 28815
rect 8893 28759 8917 28815
rect 8973 28759 8997 28815
rect 9053 28759 9077 28815
rect 9133 28759 9157 28815
rect 9213 28759 9237 28815
rect 9293 28759 9317 28815
rect 9373 28759 9397 28815
rect 9453 28759 9477 28815
rect 9533 28759 9557 28815
rect 9613 28759 9637 28815
rect 9693 28759 9717 28815
rect 9773 28759 9797 28815
rect 9853 28759 9877 28815
rect 9933 28759 9957 28815
rect 10013 28759 10856 28815
rect 8026 28703 10856 28759
rect 8026 28647 8035 28703
rect 8091 28647 8116 28703
rect 8172 28647 8197 28703
rect 8253 28647 8277 28703
rect 8333 28647 8357 28703
rect 8413 28647 8437 28703
rect 8493 28647 8517 28703
rect 8573 28647 8597 28703
rect 8653 28647 8677 28703
rect 8733 28647 8757 28703
rect 8813 28647 8837 28703
rect 8893 28647 8917 28703
rect 8973 28647 8997 28703
rect 9053 28647 9077 28703
rect 9133 28647 9157 28703
rect 9213 28647 9237 28703
rect 9293 28647 9317 28703
rect 9373 28647 9397 28703
rect 9453 28647 9477 28703
rect 9533 28647 9557 28703
rect 9613 28647 9637 28703
rect 9693 28647 9717 28703
rect 9773 28647 9797 28703
rect 9853 28647 9877 28703
rect 9933 28647 9957 28703
rect 10013 28647 10856 28703
rect 8026 15931 10856 28647
tri 7826 11622 7918 11714 sw
rect 5823 7881 5832 7937
rect 5888 7881 5913 7937
rect 5969 7881 5994 7937
rect 6050 7881 6075 7937
rect 6131 7881 6156 7937
rect 6212 7881 6237 7937
rect 6293 7881 6318 7937
rect 6374 7881 6398 7937
rect 6454 7881 6478 7937
rect 6534 7881 6558 7937
rect 6614 7881 6623 7937
rect 5823 7845 6623 7881
rect 5823 7789 5832 7845
rect 5888 7789 5913 7845
rect 5969 7789 5994 7845
rect 6050 7789 6075 7845
rect 6131 7789 6156 7845
rect 6212 7789 6237 7845
rect 6293 7789 6318 7845
rect 6374 7789 6398 7845
rect 6454 7789 6478 7845
rect 6534 7789 6558 7845
rect 6614 7789 6623 7845
rect 5823 6765 6623 7789
rect 6709 11274 6775 11279
rect 6709 11218 6714 11274
rect 6770 11218 6775 11274
rect 6709 11194 6775 11218
rect 6709 11138 6714 11194
rect 6770 11138 6775 11194
rect 6709 7062 6775 11138
rect 6709 7006 6714 7062
rect 6770 7006 6775 7062
rect 6709 6982 6775 7006
rect 6709 6926 6714 6982
rect 6770 6926 6775 6982
rect 6709 6917 6775 6926
rect 6835 11189 6901 11194
rect 6835 11133 6840 11189
rect 6896 11133 6901 11189
rect 6835 11109 6901 11133
rect 6835 11053 6840 11109
rect 6896 11053 6901 11109
rect 6835 7336 6901 11053
rect 6835 7280 6840 7336
rect 6896 7280 6901 7336
rect 6835 7256 6901 7280
rect 6835 7200 6840 7256
rect 6896 7200 6901 7256
tri 6623 6765 6676 6818 sw
rect 5823 6760 6676 6765
tri 6676 6760 6681 6765 sw
rect 5823 6716 6681 6760
tri 6681 6716 6725 6760 sw
rect 5823 6124 6725 6716
rect 5823 6068 6507 6124
rect 6563 6068 6587 6124
rect 6643 6068 6725 6124
rect 5823 6032 6725 6068
rect 5823 5976 6507 6032
rect 6563 5976 6587 6032
rect 6643 5976 6725 6032
rect 5823 5940 6725 5976
rect 5823 5884 6507 5940
rect 6563 5884 6587 5940
rect 6643 5884 6725 5940
rect 5823 5848 6725 5884
rect 5823 5792 6507 5848
rect 6563 5792 6587 5848
rect 6643 5792 6725 5848
rect 5823 5756 6725 5792
rect 5823 5700 6507 5756
rect 6563 5700 6587 5756
rect 6643 5700 6725 5756
rect 5823 5664 6725 5700
rect 5823 5608 6507 5664
rect 6563 5608 6587 5664
rect 6643 5608 6725 5664
rect 5823 5571 6725 5608
rect 5823 5515 6507 5571
rect 6563 5515 6587 5571
rect 6643 5515 6725 5571
rect 5823 4051 6725 5515
rect 5823 3995 6459 4051
rect 6515 3995 6561 4051
rect 6617 3995 6663 4051
rect 6719 3995 6725 4051
rect 5823 3970 6725 3995
rect 5823 3914 6459 3970
rect 6515 3914 6561 3970
rect 6617 3914 6663 3970
rect 6719 3914 6725 3970
rect 5823 3889 6725 3914
rect 5823 3833 6459 3889
rect 6515 3833 6561 3889
rect 6617 3833 6663 3889
rect 6719 3833 6725 3889
rect 5823 3807 6725 3833
rect 5823 3751 6459 3807
rect 6515 3751 6561 3807
rect 6617 3751 6663 3807
rect 6719 3751 6725 3807
rect 5823 3725 6725 3751
rect 5823 3669 6459 3725
rect 6515 3669 6561 3725
rect 6617 3669 6663 3725
rect 6719 3669 6725 3725
rect 5823 3321 6725 3669
rect 5823 3265 5832 3321
rect 5888 3265 5914 3321
rect 5970 3265 5995 3321
rect 6051 3265 6076 3321
rect 6132 3265 6157 3321
rect 6213 3265 6238 3321
rect 6294 3265 6319 3321
rect 6375 3265 6400 3321
rect 6456 3265 6481 3321
rect 6537 3265 6562 3321
rect 6618 3265 6725 3321
rect 5823 3241 6725 3265
rect 5823 3185 5832 3241
rect 5888 3185 5914 3241
rect 5970 3185 5995 3241
rect 6051 3185 6076 3241
rect 6132 3185 6157 3241
rect 6213 3185 6238 3241
rect 6294 3185 6319 3241
rect 6375 3185 6400 3241
rect 6456 3185 6481 3241
rect 6537 3185 6562 3241
rect 6618 3185 6725 3241
rect 5823 3137 6725 3185
rect 5823 3081 5832 3137
rect 5888 3081 5914 3137
rect 5970 3081 5995 3137
rect 6051 3081 6076 3137
rect 6132 3081 6157 3137
rect 6213 3081 6238 3137
rect 6294 3081 6319 3137
rect 6375 3081 6400 3137
rect 6456 3081 6481 3137
rect 6537 3081 6562 3137
rect 6618 3081 6725 3137
rect 5823 3057 6725 3081
rect 5823 3001 5832 3057
rect 5888 3001 5914 3057
rect 5970 3001 5995 3057
rect 6051 3001 6076 3057
rect 6132 3001 6157 3057
rect 6213 3001 6238 3057
rect 6294 3001 6319 3057
rect 6375 3001 6400 3057
rect 6456 3001 6481 3057
rect 6537 3001 6562 3057
rect 6618 3001 6725 3057
rect 5823 1050 6725 3001
rect 5823 994 5832 1050
rect 5888 994 5913 1050
rect 5969 994 5994 1050
rect 6050 994 6075 1050
rect 6131 994 6156 1050
rect 6212 994 6237 1050
rect 6293 994 6318 1050
rect 6374 994 6398 1050
rect 6454 994 6478 1050
rect 6534 994 6558 1050
rect 6614 994 6725 1050
rect 5823 0 6725 994
rect 6835 145 6901 7200
rect 6835 89 6840 145
rect 6896 89 6901 145
rect 6835 65 6901 89
rect 6835 9 6840 65
rect 6896 9 6901 65
rect 6835 0 6901 9
rect 7000 9927 7918 11622
rect 8026 11657 10022 15931
tri 10022 15787 10166 15931 nw
tri 10298 15787 10442 15931 ne
tri 8026 10644 9039 11657 ne
rect 9039 10644 10022 11657
rect 8548 10635 8698 10640
rect 8548 10579 8553 10635
rect 8609 10579 8633 10635
rect 8689 10579 8698 10635
rect 8548 10574 8698 10579
tri 8599 10568 8605 10574 ne
rect 8605 10568 8698 10574
tri 8605 10540 8633 10568 ne
rect 8378 10360 8528 10365
rect 8378 10304 8383 10360
rect 8439 10304 8463 10360
rect 8519 10304 8528 10360
rect 8378 10299 8528 10304
tri 8428 10265 8462 10299 ne
rect 7000 9343 7838 9927
tri 7838 9847 7918 9927 nw
rect 7938 9660 8084 9665
rect 7938 9604 7943 9660
rect 7999 9604 8023 9660
rect 8079 9604 8084 9660
rect 7938 9599 8084 9604
tri 7984 9565 8018 9599 ne
tri 7838 9343 7918 9423 sw
rect 7000 1711 7918 9343
rect 8018 3869 8084 9599
rect 8018 3813 8023 3869
rect 8079 3813 8084 3869
rect 8018 3789 8084 3813
rect 8018 3733 8023 3789
rect 8079 3733 8084 3789
rect 8018 3728 8084 3733
rect 7000 1655 7009 1711
rect 7065 1655 7137 1711
rect 7193 1655 7265 1711
rect 7321 1655 7393 1711
rect 7449 1655 7521 1711
rect 7577 1655 7649 1711
rect 7705 1655 7776 1711
rect 7832 1655 7918 1711
rect 7000 0 7918 1655
rect 8462 145 8528 10299
rect 8633 605 8698 10568
rect 8758 10639 8908 10644
rect 8758 10583 8767 10639
rect 8823 10583 8847 10639
rect 8903 10583 8908 10639
rect 8758 10578 8908 10583
tri 9039 10578 9105 10644 ne
rect 9105 10578 10022 10644
rect 8758 10568 8848 10578
tri 8848 10568 8858 10578 nw
tri 9105 10568 9115 10578 ne
rect 9115 10568 10022 10578
rect 8758 10567 8847 10568
tri 8847 10567 8848 10568 nw
tri 9115 10567 9116 10568 ne
rect 8758 1086 8824 10567
tri 8824 10544 8847 10567 nw
rect 8758 1030 8763 1086
rect 8819 1030 8824 1086
rect 8758 1006 8824 1030
rect 8758 950 8763 1006
rect 8819 950 8824 1006
rect 8758 941 8824 950
rect 8911 10156 8977 10161
rect 8911 10100 8916 10156
rect 8972 10100 8977 10156
rect 8911 10076 8977 10100
rect 8911 10020 8916 10076
rect 8972 10020 8977 10076
rect 8911 3295 8977 10020
rect 8911 3239 8916 3295
rect 8972 3239 8977 3295
rect 8911 3215 8977 3239
rect 8911 3159 8916 3215
rect 8972 3159 8977 3215
tri 8698 605 8732 639 sw
rect 8633 539 8761 605
tri 8661 505 8695 539 ne
rect 8462 89 8467 145
rect 8523 89 8528 145
rect 8462 65 8528 89
rect 8462 9 8467 65
rect 8523 9 8528 65
rect 8462 0 8528 9
rect 8695 145 8761 539
rect 8695 89 8700 145
rect 8756 89 8761 145
rect 8695 65 8761 89
rect 8695 9 8700 65
rect 8756 9 8761 65
rect 8695 0 8761 9
rect 8911 145 8977 3159
rect 8911 89 8916 145
rect 8972 89 8977 145
rect 8911 65 8977 89
rect 8911 9 8916 65
rect 8972 9 8977 65
rect 8911 0 8977 9
rect 9116 1214 10022 10568
rect 9116 0 9930 1214
tri 9930 1122 10022 1214 nw
rect 10130 15589 10196 15598
rect 10130 15533 10135 15589
rect 10191 15533 10196 15589
rect 10130 15509 10196 15533
rect 10130 15453 10135 15509
rect 10191 15453 10196 15509
rect 10130 12660 10196 15453
rect 10130 12604 10135 12660
rect 10191 12604 10196 12660
rect 10130 12536 10196 12604
rect 10130 12480 10135 12536
rect 10191 12480 10196 12536
tri 10096 904 10130 938 se
rect 10130 904 10196 12480
rect 10024 824 10196 904
rect 10256 10568 10322 10573
rect 10256 10512 10261 10568
rect 10317 10512 10322 10568
rect 10256 10488 10322 10512
rect 10256 10432 10261 10488
rect 10317 10432 10322 10488
rect 10256 5237 10322 10432
rect 10256 5181 10261 5237
rect 10317 5181 10322 5237
rect 10256 5157 10322 5181
rect 10256 5101 10261 5157
rect 10317 5101 10322 5157
rect 10024 145 10090 824
tri 10090 790 10124 824 nw
rect 10024 89 10029 145
rect 10085 89 10090 145
rect 10024 65 10090 89
rect 10024 9 10029 65
rect 10085 9 10090 65
rect 10024 0 10090 9
rect 10256 145 10322 5101
rect 10256 89 10261 145
rect 10317 89 10322 145
rect 10256 65 10322 89
rect 10256 9 10261 65
rect 10317 9 10322 65
rect 10256 0 10322 9
rect 10442 0 10856 15931
use nfet_CDNS_52468879185871  nfet_CDNS_52468879185871_0
timestamp 1701704242
transform 0 1 6880 -1 0 11037
box -79 -32 179 182
use nfet_CDNS_52468879185871  nfet_CDNS_52468879185871_1
timestamp 1701704242
transform 0 1 7467 1 0 12729
box -79 -32 179 182
use nfet_CDNS_52468879185871  nfet_CDNS_52468879185871_2
timestamp 1701704242
transform 0 1 6880 1 0 8377
box -79 -32 179 182
use nfet_CDNS_52468879185871  nfet_CDNS_52468879185871_3
timestamp 1701704242
transform 0 -1 7175 1 0 12729
box -79 -32 179 182
use nfet_CDNS_52468879185871  nfet_CDNS_52468879185871_4
timestamp 1701704242
transform 1 0 6431 0 -1 12327
box -79 -32 179 182
use nfet_CDNS_52468879185871  nfet_CDNS_52468879185871_5
timestamp 1701704242
transform 1 0 5038 0 1 10940
box -79 -32 179 182
use nfet_CDNS_52468879185872  nfet_CDNS_52468879185872_0
timestamp 1701704242
transform 0 1 6880 -1 0 10771
box -79 -32 1115 332
use nfet_CDNS_52468879185872  nfet_CDNS_52468879185872_1
timestamp 1701704242
transform 0 1 7467 1 0 12995
box -79 -32 1115 332
use nfet_CDNS_52468879185872  nfet_CDNS_52468879185872_2
timestamp 1701704242
transform 0 1 6880 1 0 8643
box -79 -32 1115 332
use nfet_CDNS_52468879185872  nfet_CDNS_52468879185872_3
timestamp 1701704242
transform 0 -1 7215 1 0 12995
box -79 -32 1115 332
use nfet_CDNS_52468879185872  nfet_CDNS_52468879185872_4
timestamp 1701704242
transform 1 0 6697 0 -1 12327
box -79 -32 1115 332
use nfet_CDNS_52468879185872  nfet_CDNS_52468879185872_5
timestamp 1701704242
transform 1 0 5304 0 1 10790
box -79 -32 1115 332
use nfet_CDNS_52468879185874  nfet_CDNS_52468879185874_0
timestamp 1701704242
transform 0 1 6472 1 0 12806
box -82 -32 650 182
use nfet_CDNS_52468879185874  nfet_CDNS_52468879185874_1
timestamp 1701704242
transform 0 1 6472 1 0 13430
box -82 -32 650 182
use nfet_CDNS_52468879185874  nfet_CDNS_52468879185874_2
timestamp 1701704242
transform 1 0 3958 0 1 10886
box -82 -32 650 182
use nfet_CDNS_52468879185874  nfet_CDNS_52468879185874_3
timestamp 1701704242
transform 1 0 3334 0 1 10886
box -82 -32 650 182
use nfet_CDNS_52468879185876  nfet_CDNS_52468879185876_0
timestamp 1701704242
transform 0 1 6472 1 0 12650
box -82 -32 182 182
use nfet_CDNS_52468879185876  nfet_CDNS_52468879185876_1
timestamp 1701704242
transform 1 0 3178 0 1 10886
box -82 -32 182 182
use pfet_CDNS_52468879185877  pfet_CDNS_52468879185877_0
timestamp 1701704242
transform 0 1 6976 -1 0 15962
box -119 -66 1779 666
use pfet_CDNS_52468879185877  pfet_CDNS_52468879185877_1
timestamp 1701704242
transform 0 1 6976 -1 0 6015
box -119 -66 1779 666
use pfet_CDNS_52468879185877  pfet_CDNS_52468879185877_2
timestamp 1701704242
transform 0 1 6976 -1 0 7841
box -119 -66 1779 666
use pfet_CDNS_52468879185877  pfet_CDNS_52468879185877_3
timestamp 1701704242
transform 0 1 6976 -1 0 4189
box -119 -66 1779 666
use pfet_CDNS_52468879185877  pfet_CDNS_52468879185877_4
timestamp 1701704242
transform 0 1 6976 -1 0 17788
box -119 -66 1779 666
use pfet_CDNS_52468879185877  pfet_CDNS_52468879185877_5
timestamp 1701704242
transform 0 1 6976 -1 0 19614
box -119 -66 1779 666
use pfet_CDNS_52468879185878  pfet_CDNS_52468879185878_0
timestamp 1701704242
transform 0 1 6025 1 0 18537
box -122 -66 222 366
use pfet_CDNS_52468879185878  pfet_CDNS_52468879185878_1
timestamp 1701704242
transform 1 0 4397 0 1 3209
box -122 -66 222 366
use pfet_CDNS_52468879185880  pfet_CDNS_52468879185880_0
timestamp 1701704242
transform 0 1 6025 1 0 18693
box -122 -66 690 366
use pfet_CDNS_52468879185880  pfet_CDNS_52468879185880_1
timestamp 1701704242
transform 0 1 6025 1 0 19317
box -122 -66 690 366
use pfet_CDNS_52468879185880  pfet_CDNS_52468879185880_2
timestamp 1701704242
transform 1 0 5177 0 1 3209
box -122 -66 690 366
use pfet_CDNS_52468879185880  pfet_CDNS_52468879185880_3
timestamp 1701704242
transform 1 0 4553 0 1 3209
box -122 -66 690 366
use PYres_CDNS_524688791856  PYres_CDNS_524688791856_0
timestamp 1701704242
transform 1 0 3386 0 1 27230
box -50 0 2090 100
use sky130_fd_io__pwrdet_lshv2hv_0_nmos  sky130_fd_io__pwrdet_lshv2hv_0_nmos_0
timestamp 1701704242
transform -1 0 6179 0 1 13304
box 39 29 3429 871
use sky130_fd_io__pwrdet_lshv2hv_0_nmos  sky130_fd_io__pwrdet_lshv2hv_0_nmos_1
timestamp 1701704242
transform -1 0 6572 0 1 9760
box 39 29 3429 871
use sky130_fd_io__pwrdet_lshv2hv_0_nmos  sky130_fd_io__pwrdet_lshv2hv_0_nmos_2
timestamp 1701704242
transform -1 0 6179 0 -1 13378
box 39 29 3429 871
use sky130_fd_io__pwrdet_lshv2hv_0_nmos  sky130_fd_io__pwrdet_lshv2hv_0_nmos_3
timestamp 1701704242
transform 1 0 3089 0 -1 9834
box 39 29 3429 871
use sky130_fd_io__pwrdet_lshv2hv_0_nmos  sky130_fd_io__pwrdet_lshv2hv_0_nmos_4
timestamp 1701704242
transform 1 0 3089 0 1 8050
box 39 29 3429 871
use sky130_fd_io__pwrdet_lshv2hv_0_nmos  sky130_fd_io__pwrdet_lshv2hv_0_nmos_5
timestamp 1701704242
transform 1 0 2928 0 1 11594
box 39 29 3429 871
use sky130_fd_io__pwrdet_lshv2hv_0_pmos1  sky130_fd_io__pwrdet_lshv2hv_0_pmos1_0
timestamp 1701704242
transform -1 0 4199 0 1 2410
box 0 0 1310 647
use sky130_fd_io__pwrdet_lshv2hv_0_pmos1  sky130_fd_io__pwrdet_lshv2hv_0_pmos1_1
timestamp 1701704242
transform -1 0 4199 0 1 263
box 0 0 1310 647
use sky130_fd_io__pwrdet_lshv2hv_0_pmos1  sky130_fd_io__pwrdet_lshv2hv_0_pmos1_2
timestamp 1701704242
transform -1 0 5509 0 1 263
box 0 0 1310 647
use sky130_fd_io__pwrdet_lshv2hv_0_pmos1  sky130_fd_io__pwrdet_lshv2hv_0_pmos1_3
timestamp 1701704242
transform -1 0 5509 0 1 2410
box 0 0 1310 647
use sky130_fd_io__pwrdet_lshv2hv_0_pmos1  sky130_fd_io__pwrdet_lshv2hv_0_pmos1_4
timestamp 1701704242
transform 1 0 5509 0 1 263
box 0 0 1310 647
use sky130_fd_io__pwrdet_lshv2hv_0_pmos1  sky130_fd_io__pwrdet_lshv2hv_0_pmos1_5
timestamp 1701704242
transform 1 0 5509 0 1 2410
box 0 0 1310 647
use sky130_fd_io__pwrdet_lshv2hv_0_pmos2  sky130_fd_io__pwrdet_lshv2hv_0_pmos2_0
timestamp 1701704242
transform -1 0 3672 0 1 1310
box 100 -32 896 391
use sky130_fd_io__pwrdet_lshv2hv_0_pmos2  sky130_fd_io__pwrdet_lshv2hv_0_pmos2_1
timestamp 1701704242
transform -1 0 3672 0 -1 2010
box 100 -32 896 391
use sky130_fd_io__pwrdet_lshv2hv_0_pmos2  sky130_fd_io__pwrdet_lshv2hv_0_pmos2_2
timestamp 1701704242
transform -1 0 5588 0 -1 2010
box 100 -32 896 391
use sky130_fd_io__pwrdet_lshv2hv_0_pmos2  sky130_fd_io__pwrdet_lshv2hv_0_pmos2_3
timestamp 1701704242
transform -1 0 7020 0 -1 2010
box 100 -32 896 391
use sky130_fd_io__pwrdet_lshv2hv_0_pmos2  sky130_fd_io__pwrdet_lshv2hv_0_pmos2_4
timestamp 1701704242
transform -1 0 6304 0 -1 2010
box 100 -32 896 391
use sky130_fd_io__pwrdet_lshv2hv_0_pmos2  sky130_fd_io__pwrdet_lshv2hv_0_pmos2_5
timestamp 1701704242
transform -1 0 4388 0 -1 2010
box 100 -32 896 391
use sky130_fd_io__pwrdet_vddd  sky130_fd_io__pwrdet_vddd_0
timestamp 1701704242
transform 1 0 0 0 1 0
box 348 14 10846 40000
use sky130_fd_io__pwrdet_vddio  sky130_fd_io__pwrdet_vddio_0
timestamp 1701704242
transform 1 0 0 0 1 0
box 908 0 9619 40000
<< labels >>
flabel comment s 4474 27292 4474 27292 0 FreeSans 400 0 0 0 leaker
flabel comment s 4651 8047 4651 8047 0 FreeSans 600 0 0 0 condiode
flabel metal1 s 9232 0 9284 128 3 FreeSans 200 90 0 0 in1_vddd_hv
port 2 nsew signal input
flabel metal1 s 9572 0 9624 128 3 FreeSans 200 90 0 0 in2_vddd_hv
port 3 nsew signal input
flabel metal1 s 6843 0 6895 128 3 FreeSans 200 90 0 0 out3_vddio_hv
port 4 nsew signal output
flabel metal1 s 8918 0 8970 128 3 FreeSans 200 90 0 0 out1_vddio_hv
port 5 nsew signal output
flabel metal1 s 10263 0 10315 128 3 FreeSans 200 90 0 0 out2_vddio_hv
port 6 nsew signal output
flabel metal1 s 8701 0 8753 128 3 FreeSans 200 90 0 0 out2_vddd_hv
port 7 nsew signal output
flabel metal1 s 10031 0 10083 128 3 FreeSans 200 90 0 0 out1_vddd_hv
port 8 nsew signal output
flabel metal1 s 8176 0 8228 128 3 FreeSans 200 90 0 0 vddio_present_vddd_hv
port 10 nsew signal output
flabel metal1 s 2483 0 2561 128 3 FreeSans 520 90 0 0 tie_lo_esd
port 12 nsew signal output
flabel metal1 s 282 0 334 128 3 FreeSans 200 90 0 0 rst_por_hv_n
port 13 nsew signal input
flabel metal1 s 8469 0 8521 128 3 FreeSans 200 90 0 0 out3_vddd_hv
port 14 nsew signal output
flabel metal1 s 1415 0 1467 128 3 FreeSans 200 90 0 0 in3_vddio_hv
port 15 nsew signal input
flabel metal1 s 1652 0 1704 128 3 FreeSans 200 90 0 0 in2_vddio_hv
port 16 nsew signal input
flabel metal1 s 1909 0 1961 128 3 FreeSans 200 90 0 0 vddd_present_vddio_hv
port 11 nsew signal output
flabel metal1 s 2163 0 2215 128 3 FreeSans 200 90 0 0 in3_vddd_hv
port 17 nsew signal input
flabel metal1 s 9784 0 9836 128 3 FreeSans 200 90 0 0 in1_vddio_hv
port 9 nsew signal input
flabel metal3 s 282 0 1423 242 3 FreeSans 520 0 0 0 vssio_q
port 18 nsew ground bidirectional
flabel metal3 s 1583 0 2383 242 3 FreeSans 520 0 0 0 vccd
port 19 nsew power bidirectional
flabel metal3 s 3703 0 4503 242 3 FreeSans 520 0 0 0 vddd1
port 20 nsew power bidirectional
flabel metal3 s 4663 0 5663 242 3 FreeSans 520 0 0 0 vssa
port 21 nsew ground bidirectional
flabel metal3 s 5823 0 6725 242 3 FreeSans 520 0 0 0 vddio_q
port 22 nsew power bidirectional
flabel metal3 s 7001 0 7918 242 3 FreeSans 520 0 0 0 vddd2
port 23 nsew power bidirectional
flabel metal3 s 2661 0 3543 242 3 FreeSans 520 0 0 0 vssd
port 24 nsew ground bidirectional
flabel metal3 s 2661 39758 3543 40000 3 FreeSans 520 0 0 0 vssd
port 24 nsew ground bidirectional
flabel metal3 s 3703 39758 4503 40000 3 FreeSans 520 0 0 0 vddd1
port 20 nsew power bidirectional
flabel metal3 s 6733 39758 7908 40000 3 FreeSans 520 0 0 0 vddd2
port 23 nsew power bidirectional
flabel metal3 s 4663 39758 5663 40000 3 FreeSans 520 0 0 0 vssa
port 21 nsew ground bidirectional
flabel metal3 s 5823 39758 6623 40000 3 FreeSans 520 0 0 0 vddio_q
port 22 nsew power bidirectional
flabel metal3 s 1583 39758 2501 40000 3 FreeSans 520 0 0 0 vccd
port 19 nsew power bidirectional
flabel metal2 s 2483 0 2561 128 3 FreeSans 520 90 0 0 tie_lo_esd
port 12 nsew signal output
flabel metal2 s 8176 0 8228 128 3 FreeSans 200 90 0 0 vddio_present_vddd_hv
port 10 nsew signal output
flabel metal2 s 9784 0 9836 128 3 FreeSans 200 90 0 0 in1_vddio_hv
port 9 nsew signal input
flabel metal2 s 10031 0 10083 128 3 FreeSans 200 90 0 0 out1_vddd_hv
port 8 nsew signal output
flabel metal2 s 9572 0 9624 128 3 FreeSans 200 90 0 0 in2_vddd_hv
port 3 nsew signal input
flabel metal2 s 10263 0 10315 128 3 FreeSans 200 90 0 0 out2_vddio_hv
port 6 nsew signal output
flabel metal2 s 9232 0 9284 128 3 FreeSans 200 90 0 0 in1_vddd_hv
port 2 nsew signal input
flabel metal2 s 8918 0 8970 128 3 FreeSans 200 90 0 0 out1_vddio_hv
port 5 nsew signal output
flabel metal2 s 6843 0 6895 128 3 FreeSans 200 90 0 0 out3_vddio_hv
port 4 nsew signal output
flabel metal2 s 2163 0 2215 128 3 FreeSans 200 90 0 0 in3_vddd_hv
port 17 nsew signal input
flabel metal2 s 1909 0 1961 128 3 FreeSans 200 90 0 0 vddd_present_vddio_hv
port 11 nsew signal output
flabel metal2 s 1652 0 1704 128 3 FreeSans 200 90 0 0 in2_vddio_hv
port 16 nsew signal input
flabel metal2 s 1415 0 1467 128 3 FreeSans 200 90 0 0 in3_vddio_hv
port 15 nsew signal input
flabel metal2 s 8701 0 8753 128 3 FreeSans 200 90 0 0 out2_vddd_hv
port 7 nsew signal output
flabel metal2 s 8469 0 8521 128 3 FreeSans 200 90 0 0 out3_vddd_hv
port 14 nsew signal output
flabel metal2 s 282 0 334 128 3 FreeSans 200 90 0 0 rst_por_hv_n
port 13 nsew signal input
rlabel metal1 s 2483 0 2561 164 1 tie_lo_esd
port 12 nsew signal output
rlabel metal1 s 8388 872 8440 878 1 vddio_present_vddd_hv
port 10 nsew signal output
rlabel metal1 s 8382 858 8440 872 1 vddio_present_vddd_hv
port 10 nsew signal output
rlabel metal1 s 8368 844 8440 858 1 vddio_present_vddd_hv
port 10 nsew signal output
rlabel metal1 s 8388 878 8440 1095 1 vddio_present_vddd_hv
port 10 nsew signal output
rlabel metal1 s 8176 0 8228 758 1 vddio_present_vddd_hv
port 10 nsew signal output
rlabel metal1 s 8176 786 8256 792 1 vddio_present_vddd_hv
port 10 nsew signal output
rlabel metal1 s 8176 772 8242 786 1 vddio_present_vddd_hv
port 10 nsew signal output
rlabel metal1 s 8176 758 8228 772 1 vddio_present_vddd_hv
port 10 nsew signal output
rlabel metal1 s 8176 792 8440 844 1 vddio_present_vddd_hv
port 10 nsew signal output
rlabel metal1 s 9652 377 9704 12268 1 in1_vddio_hv
port 9 nsew signal input
rlabel metal1 s 9652 371 9704 377 1 in1_vddio_hv
port 9 nsew signal input
rlabel metal1 s 9652 357 9710 371 1 in1_vddio_hv
port 9 nsew signal input
rlabel metal1 s 9652 343 9724 357 1 in1_vddio_hv
port 9 nsew signal input
rlabel metal1 s 9784 0 9836 257 1 in1_vddio_hv
port 9 nsew signal input
rlabel metal1 s 9756 285 9836 291 1 in1_vddio_hv
port 9 nsew signal input
rlabel metal1 s 9770 271 9836 285 1 in1_vddio_hv
port 9 nsew signal input
rlabel metal1 s 9784 257 9836 271 1 in1_vddio_hv
port 9 nsew signal input
rlabel metal1 s 9652 291 9836 343 1 in1_vddio_hv
port 9 nsew signal input
rlabel metal1 s 10031 0 10083 128 1 out1_vddd_hv
port 8 nsew signal output
rlabel metal1 s 9572 0 9624 1086 1 in2_vddd_hv
port 3 nsew signal input
rlabel metal1 s 10263 0 10315 128 1 out2_vddio_hv
port 6 nsew signal output
rlabel metal1 s 9492 386 9544 952 1 in1_vddd_hv
port 2 nsew signal input
rlabel metal1 s 9492 380 9544 386 1 in1_vddd_hv
port 2 nsew signal input
rlabel metal1 s 9486 366 9544 380 1 in1_vddd_hv
port 2 nsew signal input
rlabel metal1 s 9472 352 9544 366 1 in1_vddd_hv
port 2 nsew signal input
rlabel metal1 s 9232 0 9284 266 1 in1_vddd_hv
port 2 nsew signal input
rlabel metal1 s 9232 294 9312 300 1 in1_vddd_hv
port 2 nsew signal input
rlabel metal1 s 9232 280 9298 294 1 in1_vddd_hv
port 2 nsew signal input
rlabel metal1 s 9232 266 9284 280 1 in1_vddd_hv
port 2 nsew signal input
rlabel metal1 s 9232 300 9544 352 1 in1_vddd_hv
port 2 nsew signal input
rlabel metal1 s 8918 0 8970 128 1 out1_vddio_hv
port 5 nsew signal output
rlabel metal1 s 6843 0 6895 128 1 out3_vddio_hv
port 4 nsew signal output
rlabel metal1 s 1813 2076 1865 2082 1 in3_vddd_hv
port 17 nsew signal input
rlabel metal1 s 1813 2062 1871 2076 1 in3_vddd_hv
port 17 nsew signal input
rlabel metal1 s 1813 2048 1885 2062 1 in3_vddd_hv
port 17 nsew signal input
rlabel metal1 s 1813 2082 1865 10358 1 in3_vddd_hv
port 17 nsew signal input
rlabel metal1 s 2135 2159 2215 2165 1 in3_vddd_hv
port 17 nsew signal input
rlabel metal1 s 2149 2145 2215 2159 1 in3_vddd_hv
port 17 nsew signal input
rlabel metal1 s 2163 2131 2215 2145 1 in3_vddd_hv
port 17 nsew signal input
rlabel metal1 s 2163 2082 2215 2131 1 in3_vddd_hv
port 17 nsew signal input
rlabel metal1 s 2163 2076 2215 2082 1 in3_vddd_hv
port 17 nsew signal input
rlabel metal1 s 2157 2062 2215 2076 1 in3_vddd_hv
port 17 nsew signal input
rlabel metal1 s 2143 2048 2215 2062 1 in3_vddd_hv
port 17 nsew signal input
rlabel metal1 s 2135 1990 2215 1996 1 in3_vddd_hv
port 17 nsew signal input
rlabel metal1 s 2149 1976 2215 1990 1 in3_vddd_hv
port 17 nsew signal input
rlabel metal1 s 2163 1962 2215 1976 1 in3_vddd_hv
port 17 nsew signal input
rlabel metal1 s 2163 0 2215 1962 1 in3_vddd_hv
port 17 nsew signal input
rlabel metal1 s 1813 1996 2215 2048 1 in3_vddd_hv
port 17 nsew signal input
rlabel metal1 s 2087 2165 2215 2217 1 in3_vddd_hv
port 17 nsew signal input
rlabel metal1 s 1733 1900 1785 11043 1 vddd_present_vddio_hv
port 11 nsew signal output
rlabel metal1 s 1733 1894 1785 1900 1 vddd_present_vddio_hv
port 11 nsew signal output
rlabel metal1 s 1733 1880 1791 1894 1 vddd_present_vddio_hv
port 11 nsew signal output
rlabel metal1 s 1733 1866 1805 1880 1 vddd_present_vddio_hv
port 11 nsew signal output
rlabel metal1 s 1881 1808 1961 1814 1 vddd_present_vddio_hv
port 11 nsew signal output
rlabel metal1 s 1895 1794 1961 1808 1 vddd_present_vddio_hv
port 11 nsew signal output
rlabel metal1 s 1909 1780 1961 1794 1 vddd_present_vddio_hv
port 11 nsew signal output
rlabel metal1 s 1909 0 1961 1780 1 vddd_present_vddio_hv
port 11 nsew signal output
rlabel metal1 s 1733 1814 1961 1866 1 vddd_present_vddio_hv
port 11 nsew signal output
rlabel metal1 s 1859 12829 1915 12835 1 in2_vddio_hv
port 16 nsew signal input
rlabel metal1 s 1859 12815 1901 12829 1 in2_vddio_hv
port 16 nsew signal input
rlabel metal1 s 1859 12801 1887 12815 1 in2_vddio_hv
port 16 nsew signal input
rlabel metal1 s 1859 11502 1887 12801 1 in2_vddio_hv
port 16 nsew signal input
rlabel metal1 s 1859 11496 1887 11502 1 in2_vddio_hv
port 16 nsew signal input
rlabel metal1 s 1853 11482 1887 11496 1 in2_vddio_hv
port 16 nsew signal input
rlabel metal1 s 1839 11468 1887 11482 1 in2_vddio_hv
port 16 nsew signal input
rlabel metal1 s 1576 11434 1632 11440 1 in2_vddio_hv
port 16 nsew signal input
rlabel metal1 s 1576 11420 1618 11434 1 in2_vddio_hv
port 16 nsew signal input
rlabel metal1 s 1576 11406 1604 11420 1 in2_vddio_hv
port 16 nsew signal input
rlabel metal1 s 1576 2171 1604 11406 1 in2_vddio_hv
port 16 nsew signal input
rlabel metal1 s 1576 2165 1604 2171 1 in2_vddio_hv
port 16 nsew signal input
rlabel metal1 s 1576 2151 1610 2165 1 in2_vddio_hv
port 16 nsew signal input
rlabel metal1 s 1576 2137 1624 2151 1 in2_vddio_hv
port 16 nsew signal input
rlabel metal1 s 1624 2079 1704 2085 1 in2_vddio_hv
port 16 nsew signal input
rlabel metal1 s 1638 2065 1704 2079 1 in2_vddio_hv
port 16 nsew signal input
rlabel metal1 s 1652 2051 1704 2065 1 in2_vddio_hv
port 16 nsew signal input
rlabel metal1 s 1652 0 1704 2051 1 in2_vddio_hv
port 16 nsew signal input
rlabel metal1 s 1859 12835 1987 12887 1 in2_vddio_hv
port 16 nsew signal input
rlabel metal1 s 1576 11440 1887 11468 1 in2_vddio_hv
port 16 nsew signal input
rlabel metal1 s 1576 2085 1704 2137 1 in2_vddio_hv
port 16 nsew signal input
rlabel metal1 s 1579 13789 1635 13795 1 in3_vddio_hv
port 15 nsew signal input
rlabel metal1 s 1579 13775 1621 13789 1 in3_vddio_hv
port 15 nsew signal input
rlabel metal1 s 1579 13761 1607 13775 1 in3_vddio_hv
port 15 nsew signal input
rlabel metal1 s 1579 11954 1607 13761 1 in3_vddio_hv
port 15 nsew signal input
rlabel metal1 s 1579 11948 1607 11954 1 in3_vddio_hv
port 15 nsew signal input
rlabel metal1 s 1573 11934 1607 11948 1 in3_vddio_hv
port 15 nsew signal input
rlabel metal1 s 1559 11920 1607 11934 1 in3_vddio_hv
port 15 nsew signal input
rlabel metal1 s 1296 11886 1352 11892 1 in3_vddio_hv
port 15 nsew signal input
rlabel metal1 s 1296 11872 1338 11886 1 in3_vddio_hv
port 15 nsew signal input
rlabel metal1 s 1296 11858 1324 11872 1 in3_vddio_hv
port 15 nsew signal input
rlabel metal1 s 1296 1286 1324 11858 1 in3_vddio_hv
port 15 nsew signal input
rlabel metal1 s 1296 1280 1324 1286 1 in3_vddio_hv
port 15 nsew signal input
rlabel metal1 s 1296 1266 1330 1280 1 in3_vddio_hv
port 15 nsew signal input
rlabel metal1 s 1296 1252 1344 1266 1 in3_vddio_hv
port 15 nsew signal input
rlabel metal1 s 1387 1194 1467 1200 1 in3_vddio_hv
port 15 nsew signal input
rlabel metal1 s 1401 1180 1467 1194 1 in3_vddio_hv
port 15 nsew signal input
rlabel metal1 s 1415 1166 1467 1180 1 in3_vddio_hv
port 15 nsew signal input
rlabel metal1 s 1415 0 1467 1166 1 in3_vddio_hv
port 15 nsew signal input
rlabel metal1 s 1296 1200 1467 1252 1 in3_vddio_hv
port 15 nsew signal input
rlabel metal1 s 1579 13795 1707 13847 1 in3_vddio_hv
port 15 nsew signal input
rlabel metal1 s 1296 11892 1607 11920 1 in3_vddio_hv
port 15 nsew signal input
rlabel metal1 s 8701 0 8753 128 1 out2_vddd_hv
port 7 nsew signal output
rlabel metal1 s 8469 0 8521 128 1 out3_vddd_hv
port 14 nsew signal output
rlabel metal1 s 282 0 334 22755 1 rst_por_hv_n
port 13 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 11200 40000
string GDS_END 8293100
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 7616778
string LEFclass BLOCK
string LEFsymmetry R90
string path 15.675 277.575 35.475 277.575 
<< end >>
