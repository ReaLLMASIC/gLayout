magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< pwell >>
rect -68 -26 3543 106
<< ndiff >>
rect -42 57 0 80
rect -42 23 -34 57
rect -42 0 0 23
rect 3475 57 3517 80
rect 3509 23 3517 57
rect 3475 0 3517 23
<< ndiffc >>
rect -34 23 0 57
rect 3475 23 3509 57
<< ndiffres >>
rect 0 0 3475 80
<< locali >>
rect -34 57 0 73
rect -34 7 0 23
rect 3475 57 3509 73
rect 3475 7 3509 23
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_0
timestamp 1701704242
transform -1 0 8 0 1 11
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_1
timestamp 1701704242
transform 1 0 3467 0 1 11
box 0 0 1 1
<< properties >>
string GDS_END 78949142
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 78948640
<< end >>
