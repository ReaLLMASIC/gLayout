magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -119 -66 319 1466
<< mvpmos >>
rect 0 0 200 1400
<< mvpdiff >>
rect -50 0 0 1400
rect 200 0 250 1400
<< poly >>
rect 0 1400 200 1452
rect 0 -52 200 0
<< locali >>
rect -45 -4 -11 1354
rect 211 -4 245 1354
use DFL1sd_CDNS_52468879185620  DFL1sd_CDNS_52468879185620_0
timestamp 1701704242
transform 1 0 200 0 1 0
box -36 -36 89 1436
use hvDFL1sd_CDNS_5246887918573  hvDFL1sd_CDNS_5246887918573_0
timestamp 1701704242
transform -1 0 0 0 1 0
box -36 -36 89 1436
<< labels >>
flabel comment s -28 675 -28 675 0 FreeSans 300 0 0 0 S
flabel comment s 228 675 228 675 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 79931096
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 79930080
<< end >>
