magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< metal3 >>
rect 106 11282 4879 11346
rect 10078 11282 14858 11346
rect 10048 10564 10284 10565
rect 10380 10564 10616 10565
rect 10711 10564 10947 10565
rect 11048 10564 11284 10565
rect 11380 10564 11616 10565
rect 11711 10564 11947 10565
rect 12048 10564 12284 10565
rect 12380 10564 12616 10565
rect 12711 10564 12947 10565
rect 13048 10564 13284 10565
rect 13380 10564 13616 10565
rect 13711 10564 13947 10565
rect 14048 10564 14284 10565
rect 14380 10564 14616 10565
rect 10048 10330 14858 10564
rect 10048 10329 10284 10330
rect 10380 10329 10616 10330
rect 10711 10329 10947 10330
rect 11048 10329 11284 10330
rect 11380 10329 11616 10330
rect 11711 10329 11947 10330
rect 12048 10329 12284 10330
rect 12380 10329 12616 10330
rect 12711 10329 12947 10330
rect 13048 10329 13284 10330
rect 13380 10329 13616 10330
rect 13711 10329 13947 10330
rect 14048 10329 14284 10330
rect 14380 10329 14616 10330
rect 106 9548 4879 9612
rect 10078 9548 14858 9612
rect 194 7993 4879 8036
rect 194 7757 4887 7993
rect 194 7627 4879 7757
rect 194 7391 4887 7627
rect 194 7348 4879 7391
rect 10078 7348 14858 8036
<< obsm3 >>
rect 99 10330 4879 10564
<< metal4 >>
rect 0 35157 254 40000
rect 14746 35157 15000 40000
rect 0 14007 254 19000
rect 14746 14007 15000 19000
rect 0 12817 254 13707
rect 14746 12817 15000 13707
rect 0 11647 254 12537
rect 14746 11647 15000 12537
rect 0 11281 254 11347
rect 14746 11281 15000 11347
rect 0 10625 15000 11221
rect 0 10329 254 10565
rect 269 10499 333 10563
rect 351 10499 415 10563
rect 433 10499 497 10563
rect 515 10499 579 10563
rect 597 10499 661 10563
rect 678 10499 742 10563
rect 759 10499 823 10563
rect 840 10499 904 10563
rect 921 10499 985 10563
rect 1002 10499 1066 10563
rect 1083 10499 1147 10563
rect 1164 10499 1228 10563
rect 1245 10499 1309 10563
rect 1326 10499 1390 10563
rect 1407 10499 1471 10563
rect 1488 10499 1552 10563
rect 1569 10499 1633 10563
rect 1650 10499 1714 10563
rect 1731 10499 1795 10563
rect 1812 10499 1876 10563
rect 1893 10499 1957 10563
rect 1974 10499 2038 10563
rect 2055 10499 2119 10563
rect 2136 10499 2200 10563
rect 2217 10499 2281 10563
rect 2298 10499 2362 10563
rect 2379 10499 2443 10563
rect 2460 10499 2524 10563
rect 2541 10499 2605 10563
rect 2622 10499 2686 10563
rect 2703 10499 2767 10563
rect 2784 10499 2848 10563
rect 2865 10499 2929 10563
rect 2946 10499 3010 10563
rect 3027 10499 3091 10563
rect 3108 10499 3172 10563
rect 3189 10499 3253 10563
rect 3270 10499 3334 10563
rect 3351 10499 3415 10563
rect 3432 10499 3496 10563
rect 3513 10499 3577 10563
rect 3594 10499 3658 10563
rect 3675 10499 3739 10563
rect 3756 10499 3820 10563
rect 3837 10499 3901 10563
rect 3918 10499 3982 10563
rect 3999 10499 4063 10563
rect 4080 10499 4144 10563
rect 4161 10499 4225 10563
rect 4242 10499 4306 10563
rect 4323 10499 4387 10563
rect 4404 10499 4468 10563
rect 4485 10499 4549 10563
rect 4566 10499 4630 10563
rect 4647 10499 4711 10563
rect 4728 10499 4792 10563
rect 4809 10499 4873 10563
rect 269 10415 333 10479
rect 351 10415 415 10479
rect 433 10415 497 10479
rect 515 10415 579 10479
rect 597 10415 661 10479
rect 678 10415 742 10479
rect 759 10415 823 10479
rect 840 10415 904 10479
rect 921 10415 985 10479
rect 1002 10415 1066 10479
rect 1083 10415 1147 10479
rect 1164 10415 1228 10479
rect 1245 10415 1309 10479
rect 1326 10415 1390 10479
rect 1407 10415 1471 10479
rect 1488 10415 1552 10479
rect 1569 10415 1633 10479
rect 1650 10415 1714 10479
rect 1731 10415 1795 10479
rect 1812 10415 1876 10479
rect 1893 10415 1957 10479
rect 1974 10415 2038 10479
rect 2055 10415 2119 10479
rect 2136 10415 2200 10479
rect 2217 10415 2281 10479
rect 2298 10415 2362 10479
rect 2379 10415 2443 10479
rect 2460 10415 2524 10479
rect 2541 10415 2605 10479
rect 2622 10415 2686 10479
rect 2703 10415 2767 10479
rect 2784 10415 2848 10479
rect 2865 10415 2929 10479
rect 2946 10415 3010 10479
rect 3027 10415 3091 10479
rect 3108 10415 3172 10479
rect 3189 10415 3253 10479
rect 3270 10415 3334 10479
rect 3351 10415 3415 10479
rect 3432 10415 3496 10479
rect 3513 10415 3577 10479
rect 3594 10415 3658 10479
rect 3675 10415 3739 10479
rect 3756 10415 3820 10479
rect 3837 10415 3901 10479
rect 3918 10415 3982 10479
rect 3999 10415 4063 10479
rect 4080 10415 4144 10479
rect 4161 10415 4225 10479
rect 4242 10415 4306 10479
rect 4323 10415 4387 10479
rect 4404 10415 4468 10479
rect 4485 10415 4549 10479
rect 4566 10415 4630 10479
rect 4647 10415 4711 10479
rect 4728 10415 4792 10479
rect 4809 10415 4873 10479
rect 269 10331 333 10395
rect 351 10331 415 10395
rect 433 10331 497 10395
rect 515 10331 579 10395
rect 597 10331 661 10395
rect 678 10331 742 10395
rect 759 10331 823 10395
rect 840 10331 904 10395
rect 921 10331 985 10395
rect 1002 10331 1066 10395
rect 1083 10331 1147 10395
rect 1164 10331 1228 10395
rect 1245 10331 1309 10395
rect 1326 10331 1390 10395
rect 1407 10331 1471 10395
rect 1488 10331 1552 10395
rect 1569 10331 1633 10395
rect 1650 10331 1714 10395
rect 1731 10331 1795 10395
rect 1812 10331 1876 10395
rect 1893 10331 1957 10395
rect 1974 10331 2038 10395
rect 2055 10331 2119 10395
rect 2136 10331 2200 10395
rect 2217 10331 2281 10395
rect 2298 10331 2362 10395
rect 2379 10331 2443 10395
rect 2460 10331 2524 10395
rect 2541 10331 2605 10395
rect 2622 10331 2686 10395
rect 2703 10331 2767 10395
rect 2784 10331 2848 10395
rect 2865 10331 2929 10395
rect 2946 10331 3010 10395
rect 3027 10331 3091 10395
rect 3108 10331 3172 10395
rect 3189 10331 3253 10395
rect 3270 10331 3334 10395
rect 3351 10331 3415 10395
rect 3432 10331 3496 10395
rect 3513 10331 3577 10395
rect 3594 10331 3658 10395
rect 3675 10331 3739 10395
rect 3756 10331 3820 10395
rect 3837 10331 3901 10395
rect 3918 10331 3982 10395
rect 3999 10331 4063 10395
rect 4080 10331 4144 10395
rect 4161 10331 4225 10395
rect 4242 10331 4306 10395
rect 4323 10331 4387 10395
rect 4404 10331 4468 10395
rect 4485 10331 4549 10395
rect 4566 10331 4630 10395
rect 4647 10331 4711 10395
rect 4728 10331 4792 10395
rect 4809 10331 4873 10395
rect 10048 10329 10284 10565
rect 10380 10329 10616 10565
rect 10711 10329 10947 10565
rect 11048 10329 11284 10565
rect 11380 10329 11616 10565
rect 11711 10329 11947 10565
rect 12048 10329 12284 10565
rect 12380 10329 12616 10565
rect 12711 10329 12947 10565
rect 13048 10329 13284 10565
rect 13380 10329 13616 10565
rect 13711 10329 13947 10565
rect 14048 10329 14284 10565
rect 14380 10329 14616 10565
rect 14746 10329 15000 10565
rect 0 9673 15000 10269
rect 0 9547 254 9613
rect 14746 9547 15000 9613
rect 0 8317 254 9247
rect 14746 8317 15000 9247
rect 0 7993 254 8037
rect 14746 7993 15000 8037
rect 0 7757 379 7993
rect 465 7757 701 7993
rect 787 7757 1023 7993
rect 1109 7757 1345 7993
rect 1431 7757 1667 7993
rect 1753 7757 1989 7993
rect 2075 7757 2311 7993
rect 2397 7757 2633 7993
rect 2719 7757 2955 7993
rect 3041 7757 3277 7993
rect 3363 7757 3599 7993
rect 3685 7757 3921 7993
rect 4007 7757 4243 7993
rect 4329 7757 4565 7993
rect 4651 7757 4887 7993
rect 10111 7757 10347 7993
rect 10432 7757 10668 7993
rect 10753 7757 10989 7993
rect 11074 7757 11310 7993
rect 11395 7757 11631 7993
rect 11716 7757 11952 7993
rect 12037 7757 12273 7993
rect 12358 7757 12594 7993
rect 12679 7757 12915 7993
rect 13000 7757 13236 7993
rect 13321 7757 13557 7993
rect 13642 7757 13878 7993
rect 13963 7757 14199 7993
rect 14284 7757 14520 7993
rect 14605 7757 15000 7993
rect 0 7627 254 7757
rect 14746 7627 15000 7757
rect 0 7391 379 7627
rect 465 7391 701 7627
rect 787 7391 1023 7627
rect 1109 7391 1345 7627
rect 1431 7391 1667 7627
rect 1753 7391 1989 7627
rect 2075 7391 2311 7627
rect 2397 7391 2633 7627
rect 2719 7391 2955 7627
rect 3041 7391 3277 7627
rect 3363 7391 3599 7627
rect 3685 7391 3921 7627
rect 4007 7391 4243 7627
rect 4329 7391 4565 7627
rect 4651 7391 4887 7627
rect 10111 7391 10347 7627
rect 10432 7391 10668 7627
rect 10753 7391 10989 7627
rect 11074 7391 11310 7627
rect 11395 7391 11631 7627
rect 11716 7391 11952 7627
rect 12037 7391 12273 7627
rect 12358 7391 12594 7627
rect 12679 7391 12915 7627
rect 13000 7391 13236 7627
rect 13321 7391 13557 7627
rect 13642 7391 13878 7627
rect 13963 7391 14199 7627
rect 14284 7391 14520 7627
rect 14605 7391 15000 7627
rect 0 7347 254 7391
rect 14746 7347 15000 7391
rect 0 6377 254 7067
rect 14746 6377 15000 7067
rect 0 5167 254 6097
rect 14746 5167 15000 6097
rect 0 3957 254 4887
rect 14746 3957 15000 4887
rect 0 2987 193 3677
rect 14807 2987 15000 3677
rect 0 1777 254 2707
rect 14746 1777 15000 2707
rect 0 407 254 1497
rect 14746 407 15000 1497
<< obsm4 >>
rect 334 35077 14666 40000
rect 193 19080 14807 35077
rect 334 13927 14666 19080
rect 193 13787 14807 13927
rect 334 12737 14666 13787
rect 193 12617 14807 12737
rect 334 11567 14666 12617
rect 193 11427 14807 11567
rect 334 11301 14666 11427
rect 334 10499 351 10545
rect 415 10499 433 10545
rect 497 10499 515 10545
rect 579 10499 597 10545
rect 661 10499 678 10545
rect 742 10499 759 10545
rect 823 10499 840 10545
rect 904 10499 921 10545
rect 985 10499 1002 10545
rect 1066 10499 1083 10545
rect 1147 10499 1164 10545
rect 1228 10499 1245 10545
rect 1309 10499 1326 10545
rect 1390 10499 1407 10545
rect 1471 10499 1488 10545
rect 1552 10499 1569 10545
rect 1633 10499 1650 10545
rect 1714 10499 1731 10545
rect 1795 10499 1812 10545
rect 1876 10499 1893 10545
rect 1957 10499 1974 10545
rect 2038 10499 2055 10545
rect 2119 10499 2136 10545
rect 2200 10499 2217 10545
rect 2281 10499 2298 10545
rect 2362 10499 2379 10545
rect 2443 10499 2460 10545
rect 2524 10499 2541 10545
rect 2605 10499 2622 10545
rect 2686 10499 2703 10545
rect 2767 10499 2784 10545
rect 2848 10499 2865 10545
rect 2929 10499 2946 10545
rect 3010 10499 3027 10545
rect 3091 10499 3108 10545
rect 3172 10499 3189 10545
rect 3253 10499 3270 10545
rect 3334 10499 3351 10545
rect 3415 10499 3432 10545
rect 3496 10499 3513 10545
rect 3577 10499 3594 10545
rect 3658 10499 3675 10545
rect 3739 10499 3756 10545
rect 3820 10499 3837 10545
rect 3901 10499 3918 10545
rect 3982 10499 3999 10545
rect 4063 10499 4080 10545
rect 4144 10499 4161 10545
rect 4225 10499 4242 10545
rect 4306 10499 4323 10545
rect 4387 10499 4404 10545
rect 4468 10499 4485 10545
rect 4549 10499 4566 10545
rect 4630 10499 4647 10545
rect 4711 10499 4728 10545
rect 4792 10499 4809 10545
rect 4873 10499 10048 10545
rect 334 10479 10048 10499
rect 334 10415 351 10479
rect 415 10415 433 10479
rect 497 10415 515 10479
rect 579 10415 597 10479
rect 661 10415 678 10479
rect 742 10415 759 10479
rect 823 10415 840 10479
rect 904 10415 921 10479
rect 985 10415 1002 10479
rect 1066 10415 1083 10479
rect 1147 10415 1164 10479
rect 1228 10415 1245 10479
rect 1309 10415 1326 10479
rect 1390 10415 1407 10479
rect 1471 10415 1488 10479
rect 1552 10415 1569 10479
rect 1633 10415 1650 10479
rect 1714 10415 1731 10479
rect 1795 10415 1812 10479
rect 1876 10415 1893 10479
rect 1957 10415 1974 10479
rect 2038 10415 2055 10479
rect 2119 10415 2136 10479
rect 2200 10415 2217 10479
rect 2281 10415 2298 10479
rect 2362 10415 2379 10479
rect 2443 10415 2460 10479
rect 2524 10415 2541 10479
rect 2605 10415 2622 10479
rect 2686 10415 2703 10479
rect 2767 10415 2784 10479
rect 2848 10415 2865 10479
rect 2929 10415 2946 10479
rect 3010 10415 3027 10479
rect 3091 10415 3108 10479
rect 3172 10415 3189 10479
rect 3253 10415 3270 10479
rect 3334 10415 3351 10479
rect 3415 10415 3432 10479
rect 3496 10415 3513 10479
rect 3577 10415 3594 10479
rect 3658 10415 3675 10479
rect 3739 10415 3756 10479
rect 3820 10415 3837 10479
rect 3901 10415 3918 10479
rect 3982 10415 3999 10479
rect 4063 10415 4080 10479
rect 4144 10415 4161 10479
rect 4225 10415 4242 10479
rect 4306 10415 4323 10479
rect 4387 10415 4404 10479
rect 4468 10415 4485 10479
rect 4549 10415 4566 10479
rect 4630 10415 4647 10479
rect 4711 10415 4728 10479
rect 4792 10415 4809 10479
rect 4873 10415 10048 10479
rect 334 10395 10048 10415
rect 334 10349 351 10395
rect 415 10349 433 10395
rect 497 10349 515 10395
rect 579 10349 597 10395
rect 661 10349 678 10395
rect 742 10349 759 10395
rect 823 10349 840 10395
rect 904 10349 921 10395
rect 985 10349 1002 10395
rect 1066 10349 1083 10395
rect 1147 10349 1164 10395
rect 1228 10349 1245 10395
rect 1309 10349 1326 10395
rect 1390 10349 1407 10395
rect 1471 10349 1488 10395
rect 1552 10349 1569 10395
rect 1633 10349 1650 10395
rect 1714 10349 1731 10395
rect 1795 10349 1812 10395
rect 1876 10349 1893 10395
rect 1957 10349 1974 10395
rect 2038 10349 2055 10395
rect 2119 10349 2136 10395
rect 2200 10349 2217 10395
rect 2281 10349 2298 10395
rect 2362 10349 2379 10395
rect 2443 10349 2460 10395
rect 2524 10349 2541 10395
rect 2605 10349 2622 10395
rect 2686 10349 2703 10395
rect 2767 10349 2784 10395
rect 2848 10349 2865 10395
rect 2929 10349 2946 10395
rect 3010 10349 3027 10395
rect 3091 10349 3108 10395
rect 3172 10349 3189 10395
rect 3253 10349 3270 10395
rect 3334 10349 3351 10395
rect 3415 10349 3432 10395
rect 3496 10349 3513 10395
rect 3577 10349 3594 10395
rect 3658 10349 3675 10395
rect 3739 10349 3756 10395
rect 3820 10349 3837 10395
rect 3901 10349 3918 10395
rect 3982 10349 3999 10395
rect 4063 10349 4080 10395
rect 4144 10349 4161 10395
rect 4225 10349 4242 10395
rect 4306 10349 4323 10395
rect 4387 10349 4404 10395
rect 4468 10349 4485 10395
rect 4549 10349 4566 10395
rect 4630 10349 4647 10395
rect 4711 10349 4728 10395
rect 4792 10349 4809 10395
rect 4873 10349 10048 10395
rect 10284 10349 10380 10545
rect 10616 10349 10711 10545
rect 10947 10349 11048 10545
rect 11284 10349 11380 10545
rect 11616 10349 11711 10545
rect 11947 10349 12048 10545
rect 12284 10349 12380 10545
rect 12616 10349 12711 10545
rect 12947 10349 13048 10545
rect 13284 10349 13380 10545
rect 13616 10349 13711 10545
rect 13947 10349 14048 10545
rect 14284 10349 14380 10545
rect 14616 10349 14666 10545
rect 334 9467 14666 9593
rect 193 9327 14807 9467
rect 334 8237 14666 9327
rect 193 8117 14807 8237
rect 334 7993 14666 8117
rect 379 7757 465 7993
rect 701 7757 787 7993
rect 1023 7757 1109 7993
rect 1345 7757 1431 7993
rect 1667 7757 1753 7993
rect 1989 7757 2075 7993
rect 2311 7757 2397 7993
rect 2633 7757 2719 7993
rect 2955 7757 3041 7993
rect 3277 7757 3363 7993
rect 3599 7757 3685 7993
rect 3921 7757 4007 7993
rect 4243 7757 4329 7993
rect 4565 7757 4651 7993
rect 4887 7757 10111 7993
rect 10347 7757 10432 7993
rect 10668 7757 10753 7993
rect 10989 7757 11074 7993
rect 11310 7757 11395 7993
rect 11631 7757 11716 7993
rect 11952 7757 12037 7993
rect 12273 7757 12358 7993
rect 12594 7757 12679 7993
rect 12915 7757 13000 7993
rect 13236 7757 13321 7993
rect 13557 7757 13642 7993
rect 13878 7757 13963 7993
rect 14199 7757 14284 7993
rect 14520 7757 14605 7993
rect 334 7627 14666 7757
rect 379 7391 465 7627
rect 701 7391 787 7627
rect 1023 7391 1109 7627
rect 1345 7391 1431 7627
rect 1667 7391 1753 7627
rect 1989 7391 2075 7627
rect 2311 7391 2397 7627
rect 2633 7391 2719 7627
rect 2955 7391 3041 7627
rect 3277 7391 3363 7627
rect 3599 7391 3685 7627
rect 3921 7391 4007 7627
rect 4243 7391 4329 7627
rect 4565 7391 4651 7627
rect 4887 7391 10111 7627
rect 10347 7391 10432 7627
rect 10668 7391 10753 7627
rect 10989 7391 11074 7627
rect 11310 7391 11395 7627
rect 11631 7391 11716 7627
rect 11952 7391 12037 7627
rect 12273 7391 12358 7627
rect 12594 7391 12679 7627
rect 12915 7391 13000 7627
rect 13236 7391 13321 7627
rect 13557 7391 13642 7627
rect 13878 7391 13963 7627
rect 14199 7391 14284 7627
rect 14520 7391 14605 7627
rect 334 7267 14666 7391
rect 193 7147 14807 7267
rect 334 6297 14666 7147
rect 193 6177 14807 6297
rect 334 5087 14666 6177
rect 193 4967 14807 5087
rect 334 3877 14666 4967
rect 193 3757 14807 3877
rect 273 2907 14727 3757
rect 193 2787 14807 2907
rect 334 1697 14666 2787
rect 193 1577 14807 1697
rect 334 407 14666 1577
<< metal5 >>
rect 0 35157 254 40000
rect 14746 35157 15000 40000
rect 0 14007 254 18997
rect 0 12837 254 13687
rect 0 11667 254 12517
rect 0 9547 254 11347
rect 14746 14007 15000 18997
rect 14746 12837 15000 13687
rect 14746 11667 15000 12517
rect 10048 10329 10284 10565
rect 10380 10329 10616 10565
rect 10711 10329 10947 10565
rect 11048 10329 11284 10565
rect 11380 10329 11616 10565
rect 11711 10329 11947 10565
rect 12048 10329 12284 10565
rect 12380 10329 12616 10565
rect 12711 10329 12947 10565
rect 13048 10329 13284 10565
rect 13380 10329 13616 10565
rect 13711 10329 13947 10565
rect 14048 10329 14284 10565
rect 14380 10329 14616 10565
rect 0 8337 254 9227
rect 0 7993 254 8017
rect 14746 9547 15000 11347
rect 14746 8337 15000 9227
rect 14746 7993 15000 8017
rect 0 7757 379 7993
rect 465 7757 701 7993
rect 787 7757 1023 7993
rect 1109 7757 1345 7993
rect 1431 7757 1667 7993
rect 1753 7757 1989 7993
rect 2075 7757 2311 7993
rect 2397 7757 2633 7993
rect 2719 7757 2955 7993
rect 3041 7757 3277 7993
rect 3363 7757 3599 7993
rect 3685 7757 3921 7993
rect 4007 7757 4243 7993
rect 4329 7757 4565 7993
rect 4651 7757 4887 7993
rect 10111 7757 10347 7993
rect 10432 7757 10668 7993
rect 10753 7757 10989 7993
rect 11074 7757 11310 7993
rect 11395 7757 11631 7993
rect 11716 7757 11952 7993
rect 12037 7757 12273 7993
rect 12358 7757 12594 7993
rect 12679 7757 12915 7993
rect 13000 7757 13236 7993
rect 13321 7757 13557 7993
rect 13642 7757 13878 7993
rect 13963 7757 14199 7993
rect 14284 7757 14520 7993
rect 14605 7757 15000 7993
rect 0 7627 254 7757
rect 14746 7627 15000 7757
rect 0 7391 379 7627
rect 465 7391 701 7627
rect 787 7391 1023 7627
rect 1109 7391 1345 7627
rect 1431 7391 1667 7627
rect 1753 7391 1989 7627
rect 2075 7391 2311 7627
rect 2397 7391 2633 7627
rect 2719 7391 2955 7627
rect 3041 7391 3277 7627
rect 3363 7391 3599 7627
rect 3685 7391 3921 7627
rect 4007 7391 4243 7627
rect 4329 7391 4565 7627
rect 4651 7391 4887 7627
rect 10111 7391 10347 7627
rect 10432 7391 10668 7627
rect 10753 7391 10989 7627
rect 11074 7391 11310 7627
rect 11395 7391 11631 7627
rect 11716 7391 11952 7627
rect 12037 7391 12273 7627
rect 12358 7391 12594 7627
rect 12679 7391 12915 7627
rect 13000 7391 13236 7627
rect 13321 7391 13557 7627
rect 13642 7391 13878 7627
rect 13963 7391 14199 7627
rect 14284 7391 14520 7627
rect 14605 7391 15000 7627
rect 0 7368 254 7391
rect 14746 7368 15000 7391
rect 0 6397 254 7047
rect 0 5187 254 6077
rect 0 3977 254 4867
rect 14746 6397 15000 7047
rect 14746 5187 15000 6077
rect 14746 3977 15000 4867
rect 0 3007 193 3657
rect 14807 3007 15000 3657
rect 0 1797 254 2687
rect 0 427 254 1477
rect 14746 1797 15000 2687
rect 14746 427 15000 1477
<< obsm5 >>
rect 574 34837 14426 40000
rect 0 19317 15000 34837
rect 574 10565 14426 19317
rect 574 10329 10048 10565
rect 10284 10329 10380 10565
rect 10616 10329 10711 10565
rect 10947 10329 11048 10565
rect 11284 10329 11380 10565
rect 11616 10329 11711 10565
rect 11947 10329 12048 10565
rect 12284 10329 12380 10565
rect 12616 10329 12711 10565
rect 12947 10329 13048 10565
rect 13284 10329 13380 10565
rect 13616 10329 13711 10565
rect 13947 10329 14048 10565
rect 14284 10329 14380 10565
rect 574 7993 14426 10329
rect 701 7757 787 7993
rect 1023 7757 1109 7993
rect 1345 7757 1431 7993
rect 1667 7757 1753 7993
rect 1989 7757 2075 7993
rect 2311 7757 2397 7993
rect 2633 7757 2719 7993
rect 2955 7757 3041 7993
rect 3277 7757 3363 7993
rect 3599 7757 3685 7993
rect 3921 7757 4007 7993
rect 4243 7757 4329 7993
rect 4565 7757 4651 7993
rect 4887 7757 10111 7993
rect 10347 7757 10432 7993
rect 10668 7757 10753 7993
rect 10989 7757 11074 7993
rect 11310 7757 11395 7993
rect 11631 7757 11716 7993
rect 11952 7757 12037 7993
rect 12273 7757 12358 7993
rect 12594 7757 12679 7993
rect 12915 7757 13000 7993
rect 13236 7757 13321 7993
rect 13557 7757 13642 7993
rect 13878 7757 13963 7993
rect 14199 7757 14284 7993
rect 574 7627 14426 7757
rect 701 7391 787 7627
rect 1023 7391 1109 7627
rect 1345 7391 1431 7627
rect 1667 7391 1753 7627
rect 1989 7391 2075 7627
rect 2311 7391 2397 7627
rect 2633 7391 2719 7627
rect 2955 7391 3041 7627
rect 3277 7391 3363 7627
rect 3599 7391 3685 7627
rect 3921 7391 4007 7627
rect 4243 7391 4329 7627
rect 4565 7391 4651 7627
rect 4887 7391 10111 7627
rect 10347 7391 10432 7627
rect 10668 7391 10753 7627
rect 10989 7391 11074 7627
rect 11310 7391 11395 7627
rect 11631 7391 11716 7627
rect 11952 7391 12037 7627
rect 12273 7391 12358 7627
rect 12594 7391 12679 7627
rect 12915 7391 13000 7627
rect 13236 7391 13321 7627
rect 13557 7391 13642 7627
rect 13878 7391 13963 7627
rect 14199 7391 14284 7627
rect 574 7368 14426 7391
rect 0 7367 15000 7368
rect 574 3657 14426 7367
rect 513 3007 14487 3657
rect 574 427 14426 3007
<< labels >>
rlabel metal5 s 0 3007 193 3657 6 VDDA
port 1 nsew power bidirectional
rlabel metal5 s 14807 3007 15000 3657 6 VDDA
port 1 nsew power bidirectional
rlabel metal4 s 14807 2987 15000 3677 6 VDDA
port 1 nsew power bidirectional
rlabel metal4 s 0 2987 193 3677 6 VDDA
port 1 nsew power bidirectional
rlabel metal5 s 14746 1797 15000 2687 6 VCCD
port 2 nsew power bidirectional
rlabel metal5 s 0 1797 254 2687 6 VCCD
port 2 nsew power bidirectional
rlabel metal4 s 0 1777 254 2707 6 VCCD
port 2 nsew power bidirectional
rlabel metal4 s 14746 1777 15000 2707 6 VCCD
port 2 nsew power bidirectional
rlabel metal5 s 14746 14007 15000 18997 6 VDDIO
port 3 nsew power bidirectional
rlabel metal5 s 14746 3977 15000 4867 6 VDDIO
port 3 nsew power bidirectional
rlabel metal5 s 0 14007 254 18997 6 VDDIO
port 3 nsew power bidirectional
rlabel metal5 s 0 3977 254 4867 6 VDDIO
port 3 nsew power bidirectional
rlabel metal4 s 14746 3957 15000 4887 6 VDDIO
port 3 nsew power bidirectional
rlabel metal4 s 14746 14007 15000 19000 6 VDDIO
port 3 nsew power bidirectional
rlabel metal4 s 0 3957 254 4887 6 VDDIO
port 3 nsew power bidirectional
rlabel metal4 s 0 14007 254 19000 6 VDDIO
port 3 nsew power bidirectional
rlabel metal5 s 14746 12837 15000 13687 6 VDDIO_Q
port 4 nsew power bidirectional
rlabel metal5 s 0 12837 254 13687 6 VDDIO_Q
port 4 nsew power bidirectional
rlabel metal4 s 14746 12817 15000 13707 6 VDDIO_Q
port 4 nsew power bidirectional
rlabel metal4 s 0 12817 254 13707 6 VDDIO_Q
port 4 nsew power bidirectional
rlabel metal5 s 14746 35157 15000 40000 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 14746 5187 15000 6077 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 0 35157 254 40000 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 0 5187 254 6077 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14746 35157 15000 40000 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14746 5167 15000 6097 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 0 35157 254 40000 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 0 5167 254 6097 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 14746 11667 15000 12517 6 VSSIO_Q
port 6 nsew ground bidirectional
rlabel metal5 s 0 11667 254 12517 6 VSSIO_Q
port 6 nsew ground bidirectional
rlabel metal4 s 14746 11647 15000 12537 6 VSSIO_Q
port 6 nsew ground bidirectional
rlabel metal4 s 0 11647 254 12537 6 VSSIO_Q
port 6 nsew ground bidirectional
rlabel metal5 s 14746 6397 15000 7047 6 VSWITCH
port 7 nsew power bidirectional
rlabel metal5 s 0 6397 254 7047 6 VSWITCH
port 7 nsew power bidirectional
rlabel metal4 s 14746 6377 15000 7067 6 VSWITCH
port 7 nsew power bidirectional
rlabel metal4 s 0 6377 254 7067 6 VSWITCH
port 7 nsew power bidirectional
rlabel metal5 s 0 427 254 1477 6 VCCHIB
port 8 nsew power bidirectional
rlabel metal5 s 14746 427 15000 1477 6 VCCHIB
port 8 nsew power bidirectional
rlabel metal4 s 14746 407 15000 1497 6 VCCHIB
port 8 nsew power bidirectional
rlabel metal4 s 0 407 254 1497 6 VCCHIB
port 8 nsew power bidirectional
rlabel metal5 s 14746 9547 15000 11347 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 14746 7368 15000 8017 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 0 9547 254 11347 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 0 7368 254 8017 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 14746 7347 15000 8037 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 0 9547 254 9613 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 0 10329 254 10565 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 0 11281 254 11347 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 0 7347 254 8037 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 14746 9547 15000 9613 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 14746 11281 15000 11347 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 14746 10329 15000 10565 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 106 9548 4879 9612 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 106 11282 4879 11346 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 194 7348 4879 8036 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10078 7348 14858 8036 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10078 9548 14858 9612 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10078 10330 14858 10564 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10078 11282 14858 11346 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14800 11294 14840 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14800 10511 14840 10551 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14800 10427 14840 10467 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14800 10343 14840 10383 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14800 9560 14840 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14800 7980 14840 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14800 7892 14840 7932 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14800 7804 14840 7844 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14800 7716 14840 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14800 7628 14840 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14800 7540 14840 7580 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14800 7452 14840 7492 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14800 7364 14840 7404 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14719 10511 14759 10551 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14719 10427 14759 10467 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14719 10343 14759 10383 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14719 7980 14759 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14719 7892 14759 7932 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14719 7804 14759 7844 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14719 7716 14759 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14719 7628 14759 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14719 7540 14759 7580 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14719 7452 14759 7492 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14719 7364 14759 7404 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14718 11294 14758 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14718 9560 14758 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14638 10511 14678 10551 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14638 10427 14678 10467 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14638 10343 14678 10383 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14638 7980 14678 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 14605 7757 14746 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 14605 7757 14746 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14605 7757 14746 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14638 7716 14678 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14638 7628 14678 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 14605 7391 14746 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 14605 7391 14746 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14605 7391 14746 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14636 11294 14676 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14636 9560 14676 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 14380 10329 14616 10565 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 14380 10329 14616 10565 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14380 10329 14616 10565 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14557 7980 14597 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14557 7892 14597 7932 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14557 7804 14597 7844 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14557 7716 14597 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14557 7628 14597 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14557 7540 14597 7580 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14557 7452 14597 7492 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14557 7364 14597 7404 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14554 11294 14594 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14554 9560 14594 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14476 7980 14516 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 14284 7757 14520 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 14284 7757 14520 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14284 7757 14520 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14476 7716 14516 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14476 7628 14516 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 14284 7391 14520 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 14284 7391 14520 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14284 7391 14520 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14472 11294 14512 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14472 9560 14512 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14395 7716 14435 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14395 7628 14435 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14390 11294 14430 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14390 9560 14430 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14314 10511 14354 10551 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14314 10427 14354 10467 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14314 10343 14354 10383 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14314 7716 14354 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14314 7628 14354 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14308 11294 14348 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14308 9560 14348 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 14048 10329 14284 10565 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 14048 10329 14284 10565 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14048 10329 14284 10565 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14233 7980 14273 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14233 7892 14273 7932 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14233 7804 14273 7844 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14233 7716 14273 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14233 7628 14273 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14233 7540 14273 7580 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14233 7452 14273 7492 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14233 7364 14273 7404 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14227 11294 14267 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14227 9560 14267 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14152 7980 14192 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 13963 7757 14199 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 13963 7757 14199 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13963 7757 14199 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14152 7716 14192 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14152 7628 14192 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 13963 7391 14199 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 13963 7391 14199 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13963 7391 14199 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14146 11294 14186 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14146 9560 14186 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14071 7716 14111 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14071 7628 14111 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14065 11294 14105 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 14065 9560 14105 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13990 10511 14030 10551 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13990 10427 14030 10467 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13990 10343 14030 10383 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13990 7716 14030 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13990 7628 14030 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13984 11294 14024 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13984 9560 14024 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13909 10511 13949 10551 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13909 10427 13949 10467 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13909 10343 13949 10383 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13909 7980 13949 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13909 7892 13949 7932 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13909 7804 13949 7844 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13909 7716 13949 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13909 7628 13949 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13909 7540 13949 7580 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13909 7452 13949 7492 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13909 7364 13949 7404 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13903 11294 13943 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13903 9560 13943 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 13711 10329 13947 10565 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 13711 10329 13947 10565 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13711 10329 13947 10565 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13828 7980 13868 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 13642 7757 13878 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 13642 7757 13878 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13642 7757 13878 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13828 7716 13868 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13828 7628 13868 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 13642 7391 13878 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 13642 7391 13878 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13642 7391 13878 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13822 11294 13862 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13822 9560 13862 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13747 7716 13787 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13747 7628 13787 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13741 11294 13781 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13741 9560 13781 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13666 10511 13706 10551 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13666 10427 13706 10467 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13666 10343 13706 10383 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13666 7716 13706 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13666 7628 13706 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13660 11294 13700 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13660 9560 13700 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13585 10511 13625 10551 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13585 10427 13625 10467 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13585 10343 13625 10383 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13585 7980 13625 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13585 7892 13625 7932 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13585 7804 13625 7844 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13585 7716 13625 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13585 7628 13625 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13585 7540 13625 7580 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13585 7452 13625 7492 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13585 7364 13625 7404 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13579 11294 13619 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13579 9560 13619 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 13380 10329 13616 10565 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 13380 10329 13616 10565 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13380 10329 13616 10565 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13504 7980 13544 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 13321 7757 13557 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 13321 7757 13557 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13321 7757 13557 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13504 7716 13544 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13504 7628 13544 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 13321 7391 13557 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 13321 7391 13557 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13321 7391 13557 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13498 11294 13538 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13498 9560 13538 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13423 7716 13463 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13423 7628 13463 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13417 11294 13457 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13417 9560 13457 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13342 7716 13382 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13342 7628 13382 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13336 11294 13376 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13336 9560 13376 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13261 10511 13301 10551 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13261 10427 13301 10467 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13261 10343 13301 10383 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13261 7980 13301 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13261 7892 13301 7932 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13261 7804 13301 7844 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13261 7716 13301 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13261 7628 13301 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13261 7540 13301 7580 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13261 7452 13301 7492 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13261 7364 13301 7404 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13255 11294 13295 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13255 9560 13295 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 13048 10329 13284 10565 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 13048 10329 13284 10565 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13048 10329 13284 10565 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13180 7980 13220 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 13000 7757 13236 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 13000 7757 13236 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13000 7757 13236 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13180 7716 13220 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13180 7628 13220 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 13000 7391 13236 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 13000 7391 13236 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13000 7391 13236 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13174 11294 13214 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13174 9560 13214 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13099 7716 13139 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13099 7628 13139 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13093 11294 13133 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13093 9560 13133 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13018 7716 13058 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13018 7628 13058 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13012 11294 13052 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 13012 9560 13052 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12937 10511 12977 10551 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12937 10427 12977 10467 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12937 10343 12977 10383 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12937 7980 12977 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12937 7892 12977 7932 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12937 7804 12977 7844 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12937 7716 12977 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12937 7628 12977 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12937 7540 12977 7580 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12937 7452 12977 7492 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12937 7364 12977 7404 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12931 11294 12971 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12931 9560 12971 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 12711 10329 12947 10565 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 12711 10329 12947 10565 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12711 10329 12947 10565 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12856 7980 12896 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 12679 7757 12915 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 12679 7757 12915 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12679 7757 12915 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12856 7716 12896 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12856 7628 12896 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 12679 7391 12915 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 12679 7391 12915 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12679 7391 12915 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12850 11294 12890 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12850 9560 12890 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12775 7716 12815 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12775 7628 12815 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12769 11294 12809 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12769 9560 12809 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12694 7716 12734 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12694 7628 12734 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12688 11294 12728 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12688 9560 12728 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12613 10511 12653 10551 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12613 10427 12653 10467 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12613 10343 12653 10383 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12613 7980 12653 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12613 7892 12653 7932 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12613 7804 12653 7844 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12613 7716 12653 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12613 7628 12653 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12613 7540 12653 7580 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12613 7452 12653 7492 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12613 7364 12653 7404 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12607 11294 12647 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12607 9560 12647 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 12380 10329 12616 10565 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 12380 10329 12616 10565 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12380 10329 12616 10565 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12532 7980 12572 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 12358 7757 12594 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 12358 7757 12594 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12358 7757 12594 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12532 7716 12572 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12532 7628 12572 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 12358 7391 12594 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 12358 7391 12594 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12358 7391 12594 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12526 11294 12566 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12526 9560 12566 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12451 7716 12491 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12451 7628 12491 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12445 11294 12485 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12445 9560 12485 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12370 7716 12410 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12370 7628 12410 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12364 11294 12404 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12364 9560 12404 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12289 10511 12329 10551 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12289 10427 12329 10467 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12289 10343 12329 10383 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12289 7980 12329 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12289 7892 12329 7932 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12289 7804 12329 7844 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12289 7716 12329 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12289 7628 12329 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12289 7540 12329 7580 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12289 7452 12329 7492 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12289 7364 12329 7404 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12283 11294 12323 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12283 9560 12323 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 12048 10329 12284 10565 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 12048 10329 12284 10565 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12048 10329 12284 10565 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12208 7980 12248 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 12037 7757 12273 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 12037 7757 12273 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12037 7757 12273 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12208 7716 12248 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12208 7628 12248 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 12037 7391 12273 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 12037 7391 12273 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12037 7391 12273 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12202 11294 12242 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12202 9560 12242 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12127 7716 12167 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12127 7628 12167 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12121 11294 12161 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12121 9560 12161 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12046 7716 12086 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12046 7628 12086 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12040 11294 12080 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 12040 9560 12080 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11965 10511 12005 10551 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11965 10427 12005 10467 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11965 10343 12005 10383 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11965 7980 12005 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11965 7892 12005 7932 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11965 7804 12005 7844 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11965 7716 12005 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11965 7628 12005 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11965 7540 12005 7580 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11965 7452 12005 7492 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11965 7364 12005 7404 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11959 11294 11999 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11959 9560 11999 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 11711 10329 11947 10565 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 11711 10329 11947 10565 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11711 10329 11947 10565 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11884 7980 11924 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 11716 7757 11952 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 11716 7757 11952 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11716 7757 11952 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11884 7716 11924 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11884 7628 11924 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 11716 7391 11952 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 11716 7391 11952 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11716 7391 11952 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11878 11294 11918 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11878 9560 11918 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11803 7716 11843 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11803 7628 11843 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11797 11294 11837 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11797 9560 11837 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11722 7716 11762 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11722 7628 11762 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11716 11294 11756 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11716 9560 11756 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11641 10511 11681 10551 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11641 10427 11681 10467 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11641 10343 11681 10383 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11641 7980 11681 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11641 7892 11681 7932 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11641 7804 11681 7844 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11641 7716 11681 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11641 7628 11681 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11641 7540 11681 7580 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11641 7452 11681 7492 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11641 7364 11681 7404 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11635 11294 11675 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11635 9560 11675 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 11380 10329 11616 10565 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 11380 10329 11616 10565 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11380 10329 11616 10565 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11560 7980 11600 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 11395 7757 11631 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 11395 7757 11631 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11395 7757 11631 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11560 7716 11600 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11560 7628 11600 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 11395 7391 11631 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 11395 7391 11631 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11395 7391 11631 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11554 11294 11594 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11554 9560 11594 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11479 7716 11519 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11479 7628 11519 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11473 11294 11513 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11473 9560 11513 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11398 7716 11438 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11398 7628 11438 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11392 11294 11432 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11392 9560 11432 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11317 10511 11357 10551 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11317 10427 11357 10467 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11317 10343 11357 10383 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11317 7980 11357 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11317 7892 11357 7932 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11317 7804 11357 7844 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11317 7716 11357 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11317 7628 11357 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11317 7540 11357 7580 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11317 7452 11357 7492 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11317 7364 11357 7404 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11311 11294 11351 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11311 9560 11351 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 11048 10329 11284 10565 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 11048 10329 11284 10565 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11048 10329 11284 10565 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11236 7980 11276 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 11074 7757 11310 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 11074 7757 11310 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11074 7757 11310 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11236 7716 11276 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11236 7628 11276 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 11074 7391 11310 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 11074 7391 11310 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11074 7391 11310 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11230 11294 11270 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11230 9560 11270 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11155 7716 11195 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11155 7628 11195 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11149 11294 11189 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11149 9560 11189 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11074 7716 11114 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11074 7628 11114 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11068 11294 11108 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 11068 9560 11108 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10993 10511 11033 10551 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10993 10427 11033 10467 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10993 10343 11033 10383 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10993 7980 11033 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10993 7892 11033 7932 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10993 7804 11033 7844 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10993 7716 11033 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10993 7628 11033 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10993 7540 11033 7580 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10993 7452 11033 7492 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10993 7364 11033 7404 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10987 11294 11027 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10987 9560 11027 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10912 10511 10952 10551 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10912 10427 10952 10467 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10912 10343 10952 10383 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10912 7980 10952 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 10753 7757 10989 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 10753 7757 10989 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10753 7757 10989 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10912 7716 10952 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10912 7628 10952 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 10753 7391 10989 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 10753 7391 10989 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10753 7391 10989 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10906 11294 10946 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10906 9560 10946 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 10711 10329 10947 10565 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 10711 10329 10947 10565 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10711 10329 10947 10565 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10831 7716 10871 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10831 7628 10871 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10825 11294 10865 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10825 9560 10865 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10750 7716 10790 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10750 7628 10790 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10744 11294 10784 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10744 9560 10784 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10669 10511 10709 10551 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10669 10427 10709 10467 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10669 10343 10709 10383 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10669 7980 10709 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10669 7892 10709 7932 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10669 7804 10709 7844 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10669 7716 10709 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10669 7628 10709 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10669 7540 10709 7580 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10669 7452 10709 7492 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10669 7364 10709 7404 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10663 11294 10703 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10663 9560 10703 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10588 10511 10628 10551 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10588 10427 10628 10467 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10588 10343 10628 10383 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10588 7980 10628 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 10432 7757 10668 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 10432 7757 10668 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10432 7757 10668 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10588 7716 10628 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10588 7628 10628 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 10432 7391 10668 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 10432 7391 10668 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10432 7391 10668 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10582 11294 10622 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10582 9560 10622 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 10380 10329 10616 10565 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 10380 10329 10616 10565 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10380 10329 10616 10565 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10506 7716 10546 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10506 7628 10546 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10501 11294 10541 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10501 9560 10541 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10424 7716 10464 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10424 7628 10464 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10420 11294 10460 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10420 9560 10460 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10342 7980 10382 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10342 7892 10382 7932 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10342 7804 10382 7844 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10342 7716 10382 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10342 7628 10382 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10342 7540 10382 7580 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10342 7452 10382 7492 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10342 7364 10382 7404 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10339 11294 10379 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10339 9560 10379 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10260 10511 10300 10551 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10260 10427 10300 10467 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10260 10343 10300 10383 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10260 7980 10300 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 10111 7757 10347 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 10111 7757 10347 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10111 7757 10347 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10260 7716 10300 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10260 7628 10300 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 10111 7391 10347 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 10111 7391 10347 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10111 7391 10347 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10258 11294 10298 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10258 9560 10298 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 10048 10329 10284 10565 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 10048 10329 10284 10565 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10048 10329 10284 10565 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10178 7716 10218 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10178 7628 10218 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10177 11294 10217 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10177 9560 10217 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10096 11294 10136 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10096 9560 10136 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10096 7716 10136 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 10096 7628 10136 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4821 11294 4861 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 4809 10499 4873 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4809 10499 4873 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 4809 10415 4873 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4809 10415 4873 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 4809 10331 4873 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4809 10331 4873 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4821 9560 4861 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4821 7980 4861 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 4651 7757 4887 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 4651 7757 4887 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4651 7757 4887 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4821 7716 4861 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4821 7628 4861 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 4651 7391 4887 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 4651 7391 4887 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4651 7391 4887 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4741 11294 4781 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4741 9560 4781 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4741 7716 4781 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4741 7628 4781 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 4728 10499 4792 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4728 10499 4792 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 4728 10415 4792 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4728 10415 4792 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 4728 10331 4792 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4728 10331 4792 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4661 7716 4701 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4661 7628 4701 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4660 11294 4700 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4660 9560 4700 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 4647 10499 4711 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4647 10499 4711 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 4647 10415 4711 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4647 10415 4711 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 4647 10331 4711 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4647 10331 4711 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4581 7980 4621 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4581 7892 4621 7932 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4581 7804 4621 7844 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4581 7716 4621 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4581 7628 4621 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4581 7540 4621 7580 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4581 7452 4621 7492 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4581 7364 4621 7404 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4579 11294 4619 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4579 9560 4619 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 4566 10499 4630 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4566 10499 4630 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 4566 10415 4630 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4566 10415 4630 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 4566 10331 4630 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4566 10331 4630 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4501 7980 4541 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 4329 7757 4565 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 4329 7757 4565 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4329 7757 4565 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4501 7716 4541 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4501 7628 4541 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 4329 7391 4565 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 4329 7391 4565 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4329 7391 4565 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4498 11294 4538 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4498 9560 4538 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 4485 10499 4549 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4485 10499 4549 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 4485 10415 4549 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4485 10415 4549 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 4485 10331 4549 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4485 10331 4549 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4421 7716 4461 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4421 7628 4461 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4417 11294 4457 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4417 9560 4457 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 4404 10499 4468 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4404 10499 4468 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 4404 10415 4468 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4404 10415 4468 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 4404 10331 4468 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4404 10331 4468 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4341 7716 4381 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4341 7628 4381 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4336 11294 4376 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4336 9560 4376 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 4323 10499 4387 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4323 10499 4387 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 4323 10415 4387 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4323 10415 4387 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 4323 10331 4387 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4323 10331 4387 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4261 7980 4301 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4261 7892 4301 7932 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4261 7804 4301 7844 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4261 7716 4301 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4261 7628 4301 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4261 7540 4301 7580 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4261 7452 4301 7492 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4261 7364 4301 7404 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4255 11294 4295 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4255 9560 4295 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 4242 10499 4306 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4242 10499 4306 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 4242 10415 4306 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4242 10415 4306 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 4242 10331 4306 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4242 10331 4306 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4181 7980 4221 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 4007 7757 4243 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 4007 7757 4243 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4007 7757 4243 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4181 7716 4221 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4181 7628 4221 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 4007 7391 4243 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 4007 7391 4243 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4007 7391 4243 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4174 11294 4214 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4174 9560 4214 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 4161 10499 4225 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4161 10499 4225 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 4161 10415 4225 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4161 10415 4225 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 4161 10331 4225 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4161 10331 4225 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4100 7716 4140 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4100 7628 4140 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4093 11294 4133 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4093 9560 4133 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 4080 10499 4144 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4080 10499 4144 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 4080 10415 4144 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4080 10415 4144 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 4080 10331 4144 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4080 10331 4144 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4019 7716 4059 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4019 7628 4059 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4012 11294 4052 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 4012 9560 4052 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 3999 10499 4063 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3999 10499 4063 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 3999 10415 4063 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3999 10415 4063 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 3999 10331 4063 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3999 10331 4063 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3938 7980 3978 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3938 7892 3978 7932 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3938 7804 3978 7844 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3938 7716 3978 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3938 7628 3978 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3938 7540 3978 7580 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3938 7452 3978 7492 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3938 7364 3978 7404 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3931 11294 3971 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3931 9560 3971 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 3918 10499 3982 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3918 10499 3982 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 3918 10415 3982 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3918 10415 3982 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 3918 10331 3982 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3918 10331 3982 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3857 7980 3897 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 3685 7757 3921 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 3685 7757 3921 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3685 7757 3921 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3857 7716 3897 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3857 7628 3897 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 3685 7391 3921 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 3685 7391 3921 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3685 7391 3921 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3850 11294 3890 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3850 9560 3890 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 3837 10499 3901 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3837 10499 3901 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 3837 10415 3901 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3837 10415 3901 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 3837 10331 3901 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3837 10331 3901 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3776 7716 3816 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3776 7628 3816 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3769 11294 3809 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3769 9560 3809 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 3756 10499 3820 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3756 10499 3820 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 3756 10415 3820 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3756 10415 3820 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 3756 10331 3820 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3756 10331 3820 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3695 7716 3735 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3695 7628 3735 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3688 11294 3728 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3688 9560 3728 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 3675 10499 3739 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3675 10499 3739 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 3675 10415 3739 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3675 10415 3739 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 3675 10331 3739 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3675 10331 3739 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3614 7980 3654 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3614 7892 3654 7932 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3614 7804 3654 7844 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3614 7716 3654 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3614 7628 3654 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3614 7540 3654 7580 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3614 7452 3654 7492 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3614 7364 3654 7404 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3607 11294 3647 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3607 9560 3647 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 3594 10499 3658 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3594 10499 3658 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 3594 10415 3658 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3594 10415 3658 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 3594 10331 3658 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3594 10331 3658 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3533 7980 3573 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 3363 7757 3599 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 3363 7757 3599 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3363 7757 3599 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3533 7716 3573 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3533 7628 3573 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 3363 7391 3599 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 3363 7391 3599 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3363 7391 3599 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3526 11294 3566 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3526 9560 3566 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 3513 10499 3577 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3513 10499 3577 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 3513 10415 3577 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3513 10415 3577 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 3513 10331 3577 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3513 10331 3577 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3452 7716 3492 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3452 7628 3492 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3445 11294 3485 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3445 9560 3485 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 3432 10499 3496 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3432 10499 3496 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 3432 10415 3496 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3432 10415 3496 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 3432 10331 3496 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3432 10331 3496 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3371 7716 3411 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3371 7628 3411 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3364 11294 3404 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3364 9560 3404 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 3351 10499 3415 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3351 10499 3415 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 3351 10415 3415 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3351 10415 3415 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 3351 10331 3415 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3351 10331 3415 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3290 7980 3330 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3290 7892 3330 7932 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3290 7804 3330 7844 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3290 7716 3330 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3290 7628 3330 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3290 7540 3330 7580 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3290 7452 3330 7492 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3290 7364 3330 7404 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3283 11294 3323 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3283 9560 3323 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 3270 10499 3334 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3270 10499 3334 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 3270 10415 3334 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3270 10415 3334 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 3270 10331 3334 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3270 10331 3334 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3209 7980 3249 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 3041 7757 3277 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 3041 7757 3277 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3041 7757 3277 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3209 7716 3249 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3209 7628 3249 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 3041 7391 3277 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 3041 7391 3277 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3041 7391 3277 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3202 11294 3242 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3202 9560 3242 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 3189 10499 3253 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3189 10499 3253 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 3189 10415 3253 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3189 10415 3253 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 3189 10331 3253 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3189 10331 3253 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3128 7716 3168 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3128 7628 3168 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3121 11294 3161 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3121 9560 3161 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 3108 10499 3172 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3108 10499 3172 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 3108 10415 3172 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3108 10415 3172 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 3108 10331 3172 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3108 10331 3172 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3047 7716 3087 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3047 7628 3087 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3040 11294 3080 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3040 9560 3080 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 3027 10499 3091 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3027 10499 3091 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 3027 10415 3091 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3027 10415 3091 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 3027 10331 3091 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 3027 10331 3091 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2966 7980 3006 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2966 7892 3006 7932 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2966 7804 3006 7844 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2966 7716 3006 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2966 7628 3006 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2966 7540 3006 7580 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2966 7452 3006 7492 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2966 7364 3006 7404 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2959 11294 2999 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2959 9560 2999 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 2946 10499 3010 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2946 10499 3010 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 2946 10415 3010 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2946 10415 3010 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 2946 10331 3010 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2946 10331 3010 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2885 7980 2925 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 2719 7757 2955 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 2719 7757 2955 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2719 7757 2955 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2885 7716 2925 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2885 7628 2925 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 2719 7391 2955 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 2719 7391 2955 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2719 7391 2955 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2878 11294 2918 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2878 9560 2918 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 2865 10499 2929 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2865 10499 2929 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 2865 10415 2929 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2865 10415 2929 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 2865 10331 2929 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2865 10331 2929 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2804 7716 2844 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2804 7628 2844 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2797 11294 2837 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2797 9560 2837 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 2784 10499 2848 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2784 10499 2848 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 2784 10415 2848 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2784 10415 2848 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 2784 10331 2848 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2784 10331 2848 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2723 7716 2763 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2723 7628 2763 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2716 11294 2756 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2716 9560 2756 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 2703 10499 2767 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2703 10499 2767 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 2703 10415 2767 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2703 10415 2767 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 2703 10331 2767 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2703 10331 2767 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2642 7980 2682 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2642 7892 2682 7932 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2642 7804 2682 7844 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2642 7716 2682 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2642 7628 2682 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2642 7540 2682 7580 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2642 7452 2682 7492 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2642 7364 2682 7404 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2635 11294 2675 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2635 9560 2675 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 2622 10499 2686 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2622 10499 2686 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 2622 10415 2686 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2622 10415 2686 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 2622 10331 2686 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2622 10331 2686 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2561 7980 2601 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 2397 7757 2633 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 2397 7757 2633 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2397 7757 2633 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2561 7716 2601 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2561 7628 2601 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 2397 7391 2633 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 2397 7391 2633 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2397 7391 2633 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2554 11294 2594 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2554 9560 2594 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 2541 10499 2605 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2541 10499 2605 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 2541 10415 2605 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2541 10415 2605 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 2541 10331 2605 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2541 10331 2605 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2480 7716 2520 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2480 7628 2520 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2473 11294 2513 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2473 9560 2513 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 2460 10499 2524 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2460 10499 2524 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 2460 10415 2524 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2460 10415 2524 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 2460 10331 2524 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2460 10331 2524 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2399 7716 2439 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2399 7628 2439 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2392 11294 2432 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2392 9560 2432 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 2379 10499 2443 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2379 10499 2443 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 2379 10415 2443 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2379 10415 2443 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 2379 10331 2443 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2379 10331 2443 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2318 7980 2358 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2318 7892 2358 7932 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2318 7804 2358 7844 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2318 7716 2358 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2318 7628 2358 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2318 7540 2358 7580 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2318 7452 2358 7492 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2318 7364 2358 7404 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2311 11294 2351 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2311 9560 2351 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 2298 10499 2362 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2298 10499 2362 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 2298 10415 2362 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2298 10415 2362 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 2298 10331 2362 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2298 10331 2362 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2237 7980 2277 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 2075 7757 2311 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 2075 7757 2311 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2075 7757 2311 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2237 7716 2277 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2237 7628 2277 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 2075 7391 2311 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 2075 7391 2311 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2075 7391 2311 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2230 11294 2270 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2230 9560 2270 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 2217 10499 2281 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2217 10499 2281 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 2217 10415 2281 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2217 10415 2281 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 2217 10331 2281 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2217 10331 2281 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2156 7716 2196 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2156 7628 2196 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2149 11294 2189 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2149 9560 2189 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 2136 10499 2200 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2136 10499 2200 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 2136 10415 2200 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2136 10415 2200 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 2136 10331 2200 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2136 10331 2200 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2075 7716 2115 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2075 7628 2115 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2068 11294 2108 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2068 9560 2108 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 2055 10499 2119 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2055 10499 2119 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 2055 10415 2119 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2055 10415 2119 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 2055 10331 2119 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 2055 10331 2119 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1994 7980 2034 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1994 7892 2034 7932 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1994 7804 2034 7844 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1994 7716 2034 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1994 7628 2034 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1994 7540 2034 7580 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1994 7452 2034 7492 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1994 7364 2034 7404 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1987 11294 2027 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1987 9560 2027 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 1974 10499 2038 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1974 10499 2038 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 1974 10415 2038 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1974 10415 2038 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 1974 10331 2038 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1974 10331 2038 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1913 7980 1953 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 1753 7757 1989 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 1753 7757 1989 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1753 7757 1989 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1913 7716 1953 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1913 7628 1953 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 1753 7391 1989 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 1753 7391 1989 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1753 7391 1989 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1906 11294 1946 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1906 9560 1946 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 1893 10499 1957 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1893 10499 1957 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 1893 10415 1957 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1893 10415 1957 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 1893 10331 1957 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1893 10331 1957 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1832 7716 1872 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1832 7628 1872 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1825 11294 1865 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1825 9560 1865 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 1812 10499 1876 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1812 10499 1876 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 1812 10415 1876 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1812 10415 1876 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 1812 10331 1876 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1812 10331 1876 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1751 7716 1791 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1751 7628 1791 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1744 11294 1784 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1744 9560 1784 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 1731 10499 1795 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1731 10499 1795 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 1731 10415 1795 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1731 10415 1795 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 1731 10331 1795 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1731 10331 1795 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1670 7980 1710 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1670 7892 1710 7932 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1670 7804 1710 7844 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1670 7716 1710 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1670 7628 1710 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1670 7540 1710 7580 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1670 7452 1710 7492 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1670 7364 1710 7404 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1663 11294 1703 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1663 9560 1703 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 1650 10499 1714 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1650 10499 1714 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 1650 10415 1714 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1650 10415 1714 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 1650 10331 1714 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1650 10331 1714 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1589 7980 1629 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 1431 7757 1667 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 1431 7757 1667 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1431 7757 1667 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1589 7716 1629 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1589 7628 1629 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 1431 7391 1667 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 1431 7391 1667 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1431 7391 1667 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1582 11294 1622 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1582 9560 1622 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 1569 10499 1633 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1569 10499 1633 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 1569 10415 1633 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1569 10415 1633 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 1569 10331 1633 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1569 10331 1633 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1508 7716 1548 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1508 7628 1548 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1501 11294 1541 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1501 9560 1541 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 1488 10499 1552 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1488 10499 1552 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 1488 10415 1552 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1488 10415 1552 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 1488 10331 1552 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1488 10331 1552 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1427 7716 1467 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1427 7628 1467 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1420 11294 1460 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1420 9560 1460 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 1407 10499 1471 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1407 10499 1471 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 1407 10415 1471 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1407 10415 1471 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 1407 10331 1471 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1407 10331 1471 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1346 7980 1386 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1346 7892 1386 7932 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1346 7804 1386 7844 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1346 7716 1386 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1346 7628 1386 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1346 7540 1386 7580 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1346 7452 1386 7492 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1346 7364 1386 7404 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1339 11294 1379 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1339 9560 1379 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 1326 10499 1390 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1326 10499 1390 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 1326 10415 1390 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1326 10415 1390 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 1326 10331 1390 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1326 10331 1390 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1265 7980 1305 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 1109 7757 1345 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 1109 7757 1345 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1109 7757 1345 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1265 7716 1305 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1265 7628 1305 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 1109 7391 1345 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 1109 7391 1345 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1109 7391 1345 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1258 11294 1298 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1258 9560 1298 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 1245 10499 1309 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1245 10499 1309 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 1245 10415 1309 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1245 10415 1309 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 1245 10331 1309 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1245 10331 1309 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1184 7716 1224 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1184 7628 1224 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1177 11294 1217 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1177 9560 1217 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 1164 10499 1228 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1164 10499 1228 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 1164 10415 1228 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1164 10415 1228 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 1164 10331 1228 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1164 10331 1228 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1103 7716 1143 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1103 7628 1143 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1096 11294 1136 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1096 9560 1136 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 1083 10499 1147 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1083 10499 1147 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 1083 10415 1147 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1083 10415 1147 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 1083 10331 1147 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1083 10331 1147 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1022 7980 1062 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1022 7892 1062 7932 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1022 7804 1062 7844 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1022 7716 1062 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1022 7628 1062 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1022 7540 1062 7580 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1022 7452 1062 7492 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1022 7364 1062 7404 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1015 11294 1055 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1015 9560 1055 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 1002 10499 1066 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1002 10499 1066 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 1002 10415 1066 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1002 10415 1066 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 1002 10331 1066 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 1002 10331 1066 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 941 7980 981 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 787 7757 1023 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 787 7757 1023 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 787 7757 1023 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 941 7716 981 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 941 7628 981 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 787 7391 1023 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 787 7391 1023 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 787 7391 1023 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 934 11294 974 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 934 9560 974 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 921 10499 985 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 921 10499 985 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 921 10415 985 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 921 10415 985 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 921 10331 985 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 921 10331 985 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 860 7716 900 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 860 7628 900 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 853 11294 893 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 853 9560 893 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 840 10499 904 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 840 10499 904 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 840 10415 904 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 840 10415 904 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 840 10331 904 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 840 10331 904 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 779 7716 819 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 779 7628 819 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 772 11294 812 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 772 9560 812 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 759 10499 823 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 759 10499 823 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 759 10415 823 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 759 10415 823 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 759 10331 823 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 759 10331 823 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 698 7980 738 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 698 7892 738 7932 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 698 7804 738 7844 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 698 7716 738 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 698 7628 738 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 698 7540 738 7580 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 698 7452 738 7492 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 698 7364 738 7404 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 691 11294 731 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 691 9560 731 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 678 10499 742 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 678 10499 742 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 678 10415 742 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 678 10415 742 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 678 10331 742 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 678 10331 742 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 617 7980 657 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 465 7757 701 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 465 7757 701 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 465 7757 701 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 617 7716 657 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 617 7628 657 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 465 7391 701 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 465 7391 701 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 465 7391 701 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 610 11294 650 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 610 9560 650 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 597 10499 661 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 597 10499 661 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 597 10415 661 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 597 10415 661 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 597 10331 661 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 597 10331 661 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 536 7716 576 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 536 7628 576 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 529 11294 569 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 529 9560 569 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 515 10499 579 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 515 10499 579 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 515 10415 579 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 515 10415 579 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 515 10331 579 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 515 10331 579 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 455 7716 495 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 455 7628 495 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 448 11294 488 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 448 9560 488 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 433 10499 497 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 433 10499 497 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 433 10415 497 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 433 10415 497 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 433 10331 497 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 433 10331 497 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 374 7980 414 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 374 7892 414 7932 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 374 7804 414 7844 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 374 7716 414 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 374 7628 414 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 374 7540 414 7580 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 374 7452 414 7492 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 374 7364 414 7404 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 367 11294 407 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 367 9560 407 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 351 10499 415 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 351 10499 415 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 351 10415 415 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 351 10415 415 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 351 10331 415 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 351 10331 415 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 293 7980 333 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 254 7757 379 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 254 7757 379 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 254 7757 379 7993 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 293 7716 333 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 293 7628 333 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 254 7391 379 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 254 7391 379 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 254 7391 379 7627 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 286 11294 326 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 286 9560 326 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 269 10499 333 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 269 10499 333 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 269 10415 333 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 269 10415 333 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal4 s 269 10331 333 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 269 10331 333 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 212 7980 252 8020 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 212 7892 252 7932 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 212 7804 252 7844 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 212 7716 252 7756 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 212 7628 252 7668 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 212 7540 252 7580 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 212 7452 252 7492 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 212 7364 252 7404 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 205 11294 245 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 205 9560 245 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 187 10499 251 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 187 10415 251 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 187 10331 251 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 124 11294 164 11334 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 124 9560 164 9600 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 105 10499 169 10563 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 105 10415 169 10479 6 VSSA
port 9 nsew ground bidirectional
rlabel metal3 s 105 10331 169 10395 6 VSSA
port 9 nsew ground bidirectional
rlabel metal5 s 14746 8337 15000 9227 6 VSSD
port 10 nsew ground bidirectional
rlabel metal5 s 0 8337 254 9227 6 VSSD
port 10 nsew ground bidirectional
rlabel metal4 s 14746 8317 15000 9247 6 VSSD
port 10 nsew ground bidirectional
rlabel metal4 s 0 8317 254 9247 6 VSSD
port 10 nsew ground bidirectional
rlabel metal4 s 0 9673 15000 10269 6 AMUXBUS_B
port 11 nsew signal bidirectional
rlabel metal4 s 0 10625 15000 11221 6 AMUXBUS_A
port 12 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 15000 40000
string LEFclass PAD
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 11658086
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 11551190
<< end >>
