magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< obsli1 >>
rect 385 44 15623 39966
<< metal1 >>
rect 11512 668 12080 720
rect 12058 646 12080 668
rect 12099 646 12151 649
rect 12080 627 12151 646
rect 5983 547 6111 599
rect 6025 513 6111 547
rect 979 0 1031 128
rect 1231 0 1283 128
rect 6059 0 6111 513
rect 6347 0 6399 128
rect 6547 0 6599 128
rect 6745 0 6797 128
rect 7497 0 7625 128
rect 12099 0 12151 627
rect 13080 0 13132 128
<< obsm1 >>
rect 385 776 15623 40000
rect 385 655 11456 776
rect 12136 705 15623 776
rect 385 491 5927 655
rect 6167 612 11456 655
rect 385 457 5969 491
rect 385 184 6003 457
rect 385 38 923 184
rect 1087 38 1175 184
rect 1339 38 6003 184
rect 6167 590 12002 612
rect 6167 571 12024 590
rect 6167 184 12043 571
rect 6167 38 6291 184
rect 6455 38 6491 184
rect 6655 38 6689 184
rect 6853 38 7441 184
rect 7681 38 12043 184
rect 12207 184 15623 705
rect 12207 38 13024 184
rect 13188 38 15623 184
<< metal2 >>
rect 979 0 1031 128
rect 1231 0 1283 128
rect 6059 0 6111 128
rect 6347 0 6399 128
rect 6547 0 6599 128
rect 6745 0 6797 128
rect 7497 0 7625 128
rect 12099 0 12151 128
rect 13080 0 13132 128
<< obsm2 >>
rect 385 184 15623 39934
rect 385 0 923 184
rect 1087 0 1175 184
rect 1339 0 6003 184
rect 6167 0 6291 184
rect 6455 0 6491 184
rect 6655 0 6689 184
rect 6853 0 7441 184
rect 7681 0 12043 184
rect 12207 0 13024 184
rect 13188 0 15623 184
<< obsm3 >>
rect 391 0 15623 40000
<< metal4 >>
rect 0 35157 254 39999
rect 15556 35157 16000 40000
rect 0 14007 254 19000
rect 15603 14007 16000 19000
rect 0 12817 254 13707
rect 15557 12817 16000 13707
rect 0 11647 254 12537
rect 15556 11647 16000 12537
rect 0 11281 16000 11347
rect 0 10625 16000 11221
rect 0 10329 254 10565
rect 15556 10329 16000 10565
rect 0 9673 16000 10269
rect 0 9547 16000 9613
rect 0 8317 254 9247
rect 15617 8317 16000 9247
rect 0 7347 254 8037
rect 15556 7347 16000 8037
rect 0 6377 254 7067
rect 15556 6377 16000 7067
rect 0 5167 254 6097
rect 15556 5167 16000 6097
rect 0 3957 254 4887
rect 15556 3957 16000 4887
rect 0 2987 215 3677
rect 15556 2987 16000 3677
rect 0 1777 254 2707
rect 15556 1777 16000 2707
rect 0 407 254 1497
rect 15556 407 16000 1497
<< obsm4 >>
rect 0 39999 15556 40000
rect 334 35077 15476 39999
rect 0 19080 15617 35077
rect 334 13927 15523 19080
rect 0 13787 15617 13927
rect 334 12737 15477 13787
rect 0 12617 15617 12737
rect 334 11567 15476 12617
rect 0 11427 15617 11567
rect 334 10349 15476 10545
rect 0 9327 15617 9467
rect 334 8237 15537 9327
rect 0 8117 15617 8237
rect 334 7267 15476 8117
rect 0 7147 15617 7267
rect 334 6297 15476 7147
rect 0 6177 15617 6297
rect 334 5087 15476 6177
rect 0 4967 15617 5087
rect 334 3877 15476 4967
rect 0 3757 15617 3877
rect 295 2907 15476 3757
rect 0 2787 15617 2907
rect 334 1697 15476 2787
rect 0 1577 15617 1697
rect 334 407 15476 1577
<< metal5 >>
rect 0 35157 254 40000
rect 15556 35157 16000 40000
rect 0 14007 254 18997
rect 15603 14007 16000 18997
rect 0 12837 254 13687
rect 15557 12837 16000 13687
rect 0 11667 254 12517
rect 0 9547 254 11347
rect 15556 11667 16000 12517
rect 15556 9547 16000 11347
rect 0 8337 254 9227
rect 15557 8337 16000 9227
rect 0 7367 254 8017
rect 0 6397 254 7047
rect 0 5187 254 6077
rect 0 3977 254 4867
rect 15556 7367 16000 8017
rect 15556 6397 16000 7047
rect 15556 5187 16000 6077
rect 15556 3977 16000 4867
rect 0 3007 215 3657
rect 15556 3007 16000 3657
rect 0 1797 254 2687
rect 0 427 254 1477
rect 15556 1797 16000 2687
rect 15556 427 16000 1477
<< obsm5 >>
rect 574 34837 15236 40000
rect 215 19317 15603 34837
rect 574 14007 15283 19317
rect 574 12837 15237 14007
rect 574 9227 15236 12837
rect 574 8337 15237 9227
rect 574 3657 15236 8337
rect 535 3007 15236 3657
rect 574 427 15236 3007
<< labels >>
rlabel metal1 s 1231 0 1283 128 6 ref_sel<4>
port 1 nsew signal input
rlabel metal2 s 1231 0 1283 128 6 ref_sel<4>
port 1 nsew signal input
rlabel metal1 s 979 0 1031 128 6 ref_sel<3>
port 2 nsew signal input
rlabel metal2 s 979 0 1031 128 6 ref_sel<3>
port 2 nsew signal input
rlabel metal1 s 13080 0 13132 128 6 ref_sel<1>
port 3 nsew signal input
rlabel metal2 s 13080 0 13132 128 6 ref_sel<1>
port 3 nsew signal input
rlabel metal1 s 6059 0 6111 128 6 vrefgen_en
port 4 nsew signal input
rlabel metal2 s 6059 0 6111 128 6 vrefgen_en
port 4 nsew signal input
rlabel metal1 s 5983 547 6111 599 6 vrefgen_en
port 4 nsew signal input
rlabel metal1 s 6025 513 6059 547 6 vrefgen_en
port 4 nsew signal input
rlabel metal1 s 6059 128 6111 547 6 vrefgen_en
port 4 nsew signal input
rlabel metal1 s 6347 0 6399 128 6 hld_h_n
port 5 nsew signal input
rlabel metal2 s 6347 0 6399 128 6 hld_h_n
port 5 nsew signal input
rlabel metal1 s 6547 0 6599 128 6 enable_h
port 6 nsew signal input
rlabel metal2 s 6547 0 6599 128 6 enable_h
port 6 nsew signal input
rlabel metal1 s 6745 0 6797 128 6 ref_sel<2>
port 7 nsew signal input
rlabel metal2 s 6745 0 6797 128 6 ref_sel<2>
port 7 nsew signal input
rlabel metal1 s 12099 0 12151 128 6 ref_sel<0>
port 8 nsew signal input
rlabel metal2 s 12099 0 12151 128 6 ref_sel<0>
port 8 nsew signal input
rlabel metal1 s 11512 668 12080 720 6 ref_sel<0>
port 8 nsew signal input
rlabel metal1 s 12058 646 12080 668 6 ref_sel<0>
port 8 nsew signal input
rlabel metal1 s 12080 627 12099 646 6 ref_sel<0>
port 8 nsew signal input
rlabel metal1 s 12099 128 12151 649 6 ref_sel<0>
port 8 nsew signal input
rlabel metal1 s 7497 0 7625 128 6 vinref
port 9 nsew signal bidirectional
rlabel metal2 s 7497 0 7625 128 6 vinref
port 9 nsew signal bidirectional
rlabel metal5 s 0 12837 254 13687 6 vddio_q
port 10 nsew power bidirectional
rlabel metal5 s 15557 12837 16000 13687 6 vddio_q
port 10 nsew power bidirectional
rlabel metal4 s 0 12817 254 13707 6 vddio_q
port 10 nsew power bidirectional
rlabel metal4 s 15557 12817 16000 13707 6 vddio_q
port 10 nsew power bidirectional
rlabel metal5 s 0 14007 254 18997 6 vddio
port 11 nsew power bidirectional
rlabel metal5 s 0 3977 254 4867 6 vddio
port 11 nsew power bidirectional
rlabel metal5 s 15556 3977 16000 4867 6 vddio
port 11 nsew power bidirectional
rlabel metal5 s 15603 14007 16000 18997 6 vddio
port 11 nsew power bidirectional
rlabel metal4 s 0 14007 254 19000 6 vddio
port 11 nsew power bidirectional
rlabel metal4 s 0 3957 254 4887 6 vddio
port 11 nsew power bidirectional
rlabel metal4 s 15556 3957 16000 4887 6 vddio
port 11 nsew power bidirectional
rlabel metal4 s 15603 14007 16000 19000 6 vddio
port 11 nsew power bidirectional
rlabel metal5 s 0 35157 254 40000 6 vssio
port 12 nsew ground bidirectional
rlabel metal5 s 0 5187 254 6077 6 vssio
port 12 nsew ground bidirectional
rlabel metal5 s 15556 5187 16000 6077 6 vssio
port 12 nsew ground bidirectional
rlabel metal5 s 15556 35157 16000 40000 6 vssio
port 12 nsew ground bidirectional
rlabel metal4 s 0 35157 254 39999 6 vssio
port 12 nsew ground bidirectional
rlabel metal4 s 0 5167 254 6097 6 vssio
port 12 nsew ground bidirectional
rlabel metal4 s 15556 5167 16000 6097 6 vssio
port 12 nsew ground bidirectional
rlabel metal4 s 15556 35157 16000 40000 6 vssio
port 12 nsew ground bidirectional
rlabel metal5 s 0 9547 254 11347 6 vssa
port 13 nsew ground bidirectional
rlabel metal5 s 0 7367 254 8017 6 vssa
port 13 nsew ground bidirectional
rlabel metal5 s 15556 9547 16000 11347 6 vssa
port 13 nsew ground bidirectional
rlabel metal5 s 15556 7367 16000 8017 6 vssa
port 13 nsew ground bidirectional
rlabel metal4 s 0 7347 254 8037 6 vssa
port 13 nsew ground bidirectional
rlabel metal4 s 0 11281 16000 11347 6 vssa
port 13 nsew ground bidirectional
rlabel metal4 s 0 10329 254 10565 6 vssa
port 13 nsew ground bidirectional
rlabel metal4 s 0 9547 16000 9613 6 vssa
port 13 nsew ground bidirectional
rlabel metal4 s 15556 10329 16000 10565 6 vssa
port 13 nsew ground bidirectional
rlabel metal4 s 15556 7347 16000 8037 6 vssa
port 13 nsew ground bidirectional
rlabel metal5 s 0 1797 254 2687 6 vccd
port 14 nsew power bidirectional
rlabel metal5 s 15556 1797 16000 2687 6 vccd
port 14 nsew power bidirectional
rlabel metal4 s 0 1777 254 2707 6 vccd
port 14 nsew power bidirectional
rlabel metal4 s 15556 1777 16000 2707 6 vccd
port 14 nsew power bidirectional
rlabel metal5 s 0 427 254 1477 6 vcchib
port 15 nsew power bidirectional
rlabel metal5 s 15556 427 16000 1477 6 vcchib
port 15 nsew power bidirectional
rlabel metal4 s 0 407 254 1497 6 vcchib
port 15 nsew power bidirectional
rlabel metal4 s 15556 407 16000 1497 6 vcchib
port 15 nsew power bidirectional
rlabel metal5 s 0 6397 254 7047 6 vswitch
port 16 nsew power bidirectional
rlabel metal5 s 15556 6397 16000 7047 6 vswitch
port 16 nsew power bidirectional
rlabel metal4 s 0 6377 254 7067 6 vswitch
port 16 nsew power bidirectional
rlabel metal4 s 15556 6377 16000 7067 6 vswitch
port 16 nsew power bidirectional
rlabel metal5 s 0 11667 254 12517 6 vssio_q
port 17 nsew ground bidirectional
rlabel metal5 s 15556 11667 16000 12517 6 vssio_q
port 17 nsew ground bidirectional
rlabel metal4 s 0 11647 254 12537 6 vssio_q
port 17 nsew ground bidirectional
rlabel metal4 s 15556 11647 16000 12537 6 vssio_q
port 17 nsew ground bidirectional
rlabel metal5 s 0 3007 215 3657 6 vdda
port 18 nsew power bidirectional
rlabel metal5 s 15556 3007 16000 3657 6 vdda
port 18 nsew power bidirectional
rlabel metal4 s 0 2987 215 3677 6 vdda
port 18 nsew power bidirectional
rlabel metal4 s 15556 2987 16000 3677 6 vdda
port 18 nsew power bidirectional
rlabel metal5 s 0 8337 254 9227 6 vssd
port 19 nsew ground bidirectional
rlabel metal5 s 15557 8337 16000 9227 6 vssd
port 19 nsew ground bidirectional
rlabel metal4 s 0 8317 254 9247 6 vssd
port 19 nsew ground bidirectional
rlabel metal4 s 15617 8317 16000 9247 6 vssd
port 19 nsew ground bidirectional
rlabel metal4 s 0 9673 16000 10269 6 amuxbus_b
port 20 nsew signal bidirectional
rlabel metal4 s 0 10625 16000 11221 6 amuxbus_a
port 21 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 16000 40000
string LEFclass BLOCK
string LEFsymmetry R90
string LEFview TRUE
string GDS_END 26381912
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 25924122
<< end >>
