magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< nwell >>
rect 97 1268 551 1540
rect 611 1268 717 1540
<< pwell >>
rect 887 374 973 790
<< nsubdiff >>
rect 133 1470 167 1504
rect 133 1372 167 1436
rect 133 1304 167 1338
rect 647 1470 681 1504
rect 647 1372 681 1436
rect 647 1304 681 1338
<< mvpsubdiff >>
rect 913 740 947 764
rect 913 672 947 706
rect 913 604 947 638
rect 913 536 947 570
rect 913 468 947 502
rect 913 400 947 434
<< nsubdiffcont >>
rect 133 1436 167 1470
rect 133 1338 167 1372
rect 647 1436 681 1470
rect 647 1338 681 1372
<< mvpsubdiffcont >>
rect 913 706 947 740
rect 913 638 947 672
rect 913 570 947 604
rect 913 502 947 536
rect 913 434 947 468
<< poly >>
rect 274 1248 324 1278
rect 167 1232 324 1248
rect 167 1198 183 1232
rect 217 1198 251 1232
rect 285 1198 324 1232
rect 167 1182 324 1198
rect 490 1226 540 1278
rect 490 1210 667 1226
rect 490 1176 549 1210
rect 583 1176 617 1210
rect 651 1176 667 1210
rect 490 1160 667 1176
rect 14 50 148 66
rect 14 16 30 50
rect 64 16 98 50
rect 132 16 148 50
rect 14 0 148 16
rect 204 50 338 66
rect 204 16 220 50
rect 254 16 288 50
rect 322 16 338 50
rect 204 0 338 16
rect 476 50 610 66
rect 476 16 492 50
rect 526 16 560 50
rect 594 16 610 50
rect 476 0 610 16
rect 666 50 800 66
rect 666 16 682 50
rect 716 16 750 50
rect 784 16 800 50
rect 666 0 800 16
<< polycont >>
rect 183 1198 217 1232
rect 251 1198 285 1232
rect 549 1176 583 1210
rect 617 1176 651 1210
rect 30 16 64 50
rect 98 16 132 50
rect 220 16 254 50
rect 288 16 322 50
rect 492 16 526 50
rect 560 16 594 50
rect 682 16 716 50
rect 750 16 784 50
<< locali >>
rect 133 1470 167 1504
rect 133 1372 167 1436
rect 229 1490 263 1528
rect 229 1418 263 1456
rect 551 1418 585 1456
rect 647 1470 681 1504
rect 133 1304 167 1338
rect 647 1372 681 1436
rect 647 1304 681 1338
rect 229 1232 267 1238
rect 167 1198 183 1232
rect 229 1204 251 1232
rect 217 1198 251 1204
rect 285 1198 301 1204
rect 335 1164 369 1300
rect 445 1238 479 1300
rect 443 1204 481 1238
rect 549 1210 651 1226
rect 333 1130 371 1164
rect -17 1012 17 1050
rect 335 988 369 1130
rect 445 1012 479 1204
rect 583 1176 617 1210
rect 549 1164 651 1176
rect 581 1130 619 1164
rect 797 1012 831 1050
rect -17 940 17 978
rect 797 940 831 978
rect 913 740 947 764
rect 913 672 947 706
rect 913 604 947 638
rect 913 536 947 570
rect 913 468 947 502
rect 913 400 947 434
rect 157 342 195 376
rect 619 342 657 376
rect 78 50 116 60
rect 700 50 738 58
rect 14 16 30 50
rect 78 26 98 50
rect 64 16 98 26
rect 132 16 148 26
rect 204 16 220 50
rect 254 16 288 50
rect 322 16 338 50
rect 476 16 492 50
rect 526 16 560 50
rect 594 16 610 50
rect 716 24 738 50
rect 666 16 682 24
rect 716 16 750 24
rect 784 16 800 50
<< viali >>
rect 229 1528 263 1562
rect 229 1456 263 1490
rect 229 1384 263 1418
rect 551 1456 585 1490
rect 551 1384 585 1418
rect 195 1232 229 1238
rect 267 1232 301 1238
rect 195 1204 217 1232
rect 217 1204 229 1232
rect 267 1204 285 1232
rect 285 1204 301 1232
rect 409 1204 443 1238
rect 481 1204 515 1238
rect 299 1130 333 1164
rect 371 1130 405 1164
rect -17 1050 17 1084
rect -17 978 17 1012
rect 547 1130 581 1164
rect 619 1130 653 1164
rect 797 1050 831 1084
rect -17 906 17 940
rect 797 978 831 1012
rect 797 906 831 940
rect 123 342 157 376
rect 195 342 229 376
rect 585 342 619 376
rect 657 342 691 376
rect 44 50 78 60
rect 116 50 150 60
rect 666 50 700 58
rect 738 50 772 58
rect 44 26 64 50
rect 64 26 78 50
rect 116 26 132 50
rect 132 26 150 50
rect 666 24 682 50
rect 682 24 700 50
rect 738 24 750 50
rect 750 24 772 50
<< metal1 >>
rect 223 1562 605 1574
rect 223 1528 229 1562
rect 263 1528 605 1562
rect 223 1490 605 1528
rect 223 1456 229 1490
rect 263 1456 551 1490
rect 585 1456 605 1490
rect 223 1418 605 1456
rect 223 1384 229 1418
rect 263 1384 551 1418
rect 585 1384 605 1418
rect 223 1372 605 1384
rect 183 1238 527 1244
rect 183 1204 195 1238
rect 229 1204 267 1238
rect 301 1204 409 1238
rect 443 1204 481 1238
rect 515 1204 527 1238
rect 183 1198 527 1204
rect 287 1164 665 1170
rect 287 1130 299 1164
rect 333 1130 371 1164
rect 405 1130 547 1164
rect 581 1130 619 1164
rect 653 1130 665 1164
rect 287 1124 665 1130
rect -25 1084 853 1096
rect -25 1050 -17 1084
rect 17 1050 797 1084
rect 831 1050 853 1084
rect -25 1012 853 1050
rect -25 978 -17 1012
rect 17 978 797 1012
rect 831 978 853 1012
rect -25 940 853 978
rect -25 906 -17 940
rect 17 906 797 940
rect 831 906 853 940
rect -25 894 853 906
rect 111 376 703 382
rect 111 342 123 376
rect 157 342 195 376
rect 229 342 585 376
rect 619 342 657 376
rect 691 342 703 376
rect 111 336 703 342
tri 32 66 40 74 se
rect 40 66 774 74
tri 774 66 782 74 sw
rect 32 64 782 66
tri 782 64 784 66 sw
rect 32 60 784 64
rect 32 26 44 60
rect 78 26 116 60
rect 150 58 784 60
rect 150 44 666 58
rect 150 26 162 44
rect 32 20 162 26
rect 654 24 666 44
rect 700 24 738 58
rect 772 24 784 58
rect 654 18 784 24
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1701704242
transform 0 -1 585 -1 0 1490
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1701704242
transform -1 0 150 0 1 26
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1701704242
transform -1 0 772 0 1 24
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_3
timestamp 1701704242
transform -1 0 229 0 -1 376
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_4
timestamp 1701704242
transform -1 0 691 0 -1 376
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_5
timestamp 1701704242
transform 1 0 547 0 1 1130
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_6
timestamp 1701704242
transform 1 0 195 0 1 1204
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_7
timestamp 1701704242
transform 1 0 409 0 1 1204
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_8
timestamp 1701704242
transform 1 0 299 0 1 1130
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_0
timestamp 1701704242
transform 0 1 797 -1 0 1084
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_1
timestamp 1701704242
transform 0 1 -17 1 0 906
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_2
timestamp 1701704242
transform 0 -1 263 1 0 1384
box 0 0 1 1
use nfet_CDNS_5246887918591  nfet_CDNS_5246887918591_0
timestamp 1701704242
transform 1 0 204 0 -1 1092
box -79 -26 199 1026
use nfet_CDNS_5246887918594  nfet_CDNS_5246887918594_0
timestamp 1701704242
transform -1 0 610 0 -1 1092
box -79 -26 199 1026
use nfet_CDNS_52468879185124  nfet_CDNS_52468879185124_0
timestamp 1701704242
transform -1 0 786 0 -1 1092
box -79 -26 199 1026
use nfet_CDNS_52468879185124  nfet_CDNS_52468879185124_1
timestamp 1701704242
transform 1 0 28 0 -1 1092
box -79 -26 199 1026
use pfet_CDNS_5246887918595  pfet_CDNS_5246887918595_0
timestamp 1701704242
transform -1 0 540 0 1 1304
box -89 -36 139 236
use pfet_CDNS_5246887918595  pfet_CDNS_5246887918595_1
timestamp 1701704242
transform 1 0 274 0 1 1304
box -89 -36 139 236
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_0
timestamp 1701704242
transform 1 0 533 0 1 1160
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_0
timestamp 1701704242
transform 0 1 204 1 0 0
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_1
timestamp 1701704242
transform 0 1 476 1 0 0
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_2
timestamp 1701704242
transform 0 1 666 1 0 0
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_3
timestamp 1701704242
transform 0 1 167 1 0 1182
box 0 0 1 1
use PYL1_CDNS_52468879185123  PYL1_CDNS_52468879185123_0
timestamp 1701704242
transform 1 0 14 0 1 0
box 0 0 1 1
<< labels >>
flabel metal1 s 0 894 25 1096 3 FreeSans 400 0 0 0 vgnd
port 1 nsew
flabel metal1 s 223 1372 246 1574 3 FreeSans 400 0 0 0 vpwr
port 2 nsew
flabel metal1 s 403 378 403 378 0 FreeSans 400 0 0 0 vgnd_en
flabel metal1 s 299 1130 332 1164 0 FreeSans 200 0 0 0 out_c
port 4 nsew
flabel metal1 s 481 1204 515 1238 0 FreeSans 200 0 0 0 out_t
port 3 nsew
flabel locali s 647 1387 681 1421 0 FreeSans 200 0 0 0 vpb
port 6 nsew
flabel locali s 716 16 750 50 0 FreeSans 600 0 0 0 en_h
port 7 nsew
flabel locali s 526 16 560 50 0 FreeSans 600 0 0 0 in_c
port 8 nsew
flabel locali s 254 16 288 50 0 FreeSans 600 0 0 0 in_t
port 9 nsew
flabel locali s 64 16 98 50 0 FreeSans 600 0 0 0 en_h
port 7 nsew
<< properties >>
string GDS_END 85564804
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85559532
string path 3.750 38.250 3.750 31.950 
<< end >>
