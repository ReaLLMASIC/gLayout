magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -119 -66 375 216
<< mvpmos >>
rect 0 0 100 150
rect 156 0 256 150
<< mvpdiff >>
rect -53 114 0 150
rect -53 80 -45 114
rect -11 80 0 114
rect -53 46 0 80
rect -53 12 -45 46
rect -11 12 0 46
rect -53 0 0 12
rect 100 114 156 150
rect 100 80 111 114
rect 145 80 156 114
rect 100 46 156 80
rect 100 12 111 46
rect 145 12 156 46
rect 100 0 156 12
rect 256 114 309 150
rect 256 80 267 114
rect 301 80 309 114
rect 256 46 309 80
rect 256 12 267 46
rect 301 12 309 46
rect 256 0 309 12
<< mvpdiffc >>
rect -45 80 -11 114
rect -45 12 -11 46
rect 111 80 145 114
rect 111 12 145 46
rect 267 80 301 114
rect 267 12 301 46
<< poly >>
rect 0 150 100 182
rect 156 150 256 182
rect 0 -32 100 0
rect 156 -32 256 0
<< locali >>
rect -45 114 -11 130
rect -45 46 -11 68
rect 111 114 145 130
rect 111 46 145 80
rect 111 -4 145 12
rect 267 114 301 130
rect 267 46 301 68
<< viali >>
rect -45 80 -11 102
rect -45 68 -11 80
rect -45 12 -11 30
rect -45 -4 -11 12
rect 267 80 301 102
rect 267 68 301 80
rect 267 12 301 30
rect 267 -4 301 12
<< metal1 >>
rect -51 102 -5 114
rect -51 68 -45 102
rect -11 68 -5 102
rect -51 30 -5 68
rect -51 -4 -45 30
rect -11 -4 -5 30
rect -51 -16 -5 -4
rect 261 102 307 114
rect 261 68 267 102
rect 301 68 307 102
rect 261 30 307 68
rect 261 -4 267 30
rect 301 -4 307 30
rect 261 -16 307 -4
use hvDFL1sd2_CDNS_52468879185654  hvDFL1sd2_CDNS_52468879185654_0
timestamp 1701704242
transform 1 0 100 0 1 0
box 0 0 1 1
use hvDFM1sd_CDNS_52468879185172  hvDFM1sd_CDNS_52468879185172_0
timestamp 1701704242
transform -1 0 0 0 1 0
box 0 0 1 1
use hvDFM1sd_CDNS_52468879185172  hvDFM1sd_CDNS_52468879185172_1
timestamp 1701704242
transform 1 0 256 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s -28 49 -28 49 0 FreeSans 300 0 0 0 D
flabel comment s 128 63 128 63 0 FreeSans 300 0 0 0 S
flabel comment s 284 49 284 49 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 85607732
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85606214
<< end >>
