magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< mvpmosesd >>
tri 579 2604 599 2624 sw
tri 3659 2604 3679 2624 se
rect 579 2494 3679 2604
tri 3821 2604 3841 2624 sw
tri 6901 2604 6921 2624 se
tri 579 2474 599 2494 nw
tri 3659 2474 3679 2494 ne
rect 3821 2494 6921 2604
tri 7063 2604 7083 2624 sw
tri 10143 2604 10163 2624 se
tri 3821 2474 3841 2494 nw
tri 6901 2474 6921 2494 ne
rect 7063 2494 10163 2604
tri 10305 2604 10325 2624 sw
tri 13385 2604 13405 2624 se
tri 7063 2474 7083 2494 nw
tri 10143 2474 10163 2494 ne
rect 10305 2494 13405 2604
tri 13547 2604 13567 2624 sw
tri 16627 2604 16647 2624 se
tri 10305 2474 10325 2494 nw
tri 13385 2474 13405 2494 ne
rect 13547 2494 16647 2604
tri 13547 2474 13567 2494 nw
tri 16627 2474 16647 2494 ne
tri 16789 2604 16809 2624 sw
tri 19869 2604 19889 2624 se
rect 16789 2494 19889 2604
tri 16789 2474 16809 2494 nw
tri 19869 2474 19889 2494 ne
tri 579 2192 599 2212 sw
tri 3659 2192 3679 2212 se
rect 579 2082 3679 2192
tri 3821 2192 3841 2212 sw
tri 6901 2192 6921 2212 se
tri 579 2062 599 2082 nw
tri 3659 2062 3679 2082 ne
rect 3821 2082 6921 2192
tri 7063 2192 7083 2212 sw
tri 10143 2192 10163 2212 se
tri 3821 2062 3841 2082 nw
tri 6901 2062 6921 2082 ne
rect 7063 2082 10163 2192
tri 10305 2192 10325 2212 sw
tri 13385 2192 13405 2212 se
tri 7063 2062 7083 2082 nw
tri 10143 2062 10163 2082 ne
rect 10305 2082 13405 2192
tri 13547 2192 13567 2212 sw
tri 16627 2192 16647 2212 se
tri 10305 2062 10325 2082 nw
tri 13385 2062 13405 2082 ne
rect 13547 2082 16647 2192
tri 13547 2062 13567 2082 nw
tri 16627 2062 16647 2082 ne
tri 16789 2192 16809 2212 sw
tri 19869 2192 19889 2212 se
rect 16789 2082 19889 2192
tri 16789 2062 16809 2082 nw
tri 19869 2062 19889 2082 ne
<< poly >>
rect 481 2624 559 2644
tri 559 2624 579 2644 sw
tri 3679 2624 3699 2644 se
rect 3699 2624 3801 2644
tri 3801 2624 3821 2644 sw
tri 6921 2624 6941 2644 se
rect 6941 2624 7043 2644
tri 7043 2624 7063 2644 sw
tri 10163 2624 10183 2644 se
rect 10183 2624 10285 2644
tri 10285 2624 10305 2644 sw
tri 13405 2624 13425 2644 se
rect 13425 2624 13527 2644
tri 13527 2624 13547 2644 sw
tri 16647 2624 16667 2644 se
rect 16667 2624 16697 2644
rect 481 2598 579 2624
rect 481 2564 497 2598
rect 531 2564 579 2598
rect 481 2530 579 2564
rect 481 2496 497 2530
rect 531 2496 579 2530
rect 481 2474 579 2496
rect 3679 2600 3821 2624
rect 3679 2566 3738 2600
rect 3772 2566 3821 2600
rect 3679 2532 3821 2566
rect 3679 2498 3738 2532
rect 3772 2498 3821 2532
rect 3679 2474 3821 2498
rect 6921 2600 7063 2624
rect 6921 2566 6980 2600
rect 7014 2566 7063 2600
rect 6921 2532 7063 2566
rect 6921 2498 6980 2532
rect 7014 2498 7063 2532
rect 6921 2474 7063 2498
rect 10163 2598 10305 2624
rect 10163 2564 10222 2598
rect 10256 2564 10305 2598
rect 10163 2530 10305 2564
rect 10163 2496 10222 2530
rect 10256 2496 10305 2530
rect 10163 2474 10305 2496
rect 13405 2598 13547 2624
rect 13405 2564 13465 2598
rect 13499 2564 13547 2598
rect 13405 2530 13547 2564
rect 13405 2496 13465 2530
rect 13499 2496 13547 2530
rect 13405 2474 13547 2496
rect 16647 2474 16697 2624
rect 481 2454 559 2474
tri 559 2454 579 2474 nw
tri 3679 2454 3699 2474 ne
rect 3699 2454 3801 2474
tri 3801 2454 3821 2474 nw
tri 6921 2454 6941 2474 ne
rect 6941 2454 7043 2474
tri 7043 2454 7063 2474 nw
tri 10163 2454 10183 2474 ne
rect 10183 2454 10285 2474
tri 10285 2454 10305 2474 nw
tri 13405 2454 13425 2474 ne
rect 13425 2454 13527 2474
tri 13527 2454 13547 2474 nw
tri 16647 2454 16667 2474 ne
rect 16667 2454 16697 2474
rect 16739 2624 16769 2644
tri 16769 2624 16789 2644 sw
tri 19889 2624 19909 2644 se
rect 19909 2624 19987 2644
rect 16739 2474 16789 2624
rect 19889 2600 19987 2624
rect 19889 2566 19937 2600
rect 19971 2566 19987 2600
rect 19889 2532 19987 2566
rect 19889 2498 19937 2532
rect 19971 2498 19987 2532
rect 19889 2474 19987 2498
rect 16739 2454 16769 2474
tri 16769 2454 16789 2474 nw
tri 19889 2454 19909 2474 ne
rect 19909 2454 19987 2474
rect 481 2212 559 2232
tri 559 2212 579 2232 sw
tri 3679 2212 3699 2232 se
rect 3699 2212 3801 2232
tri 3801 2212 3821 2232 sw
tri 6921 2212 6941 2232 se
rect 6941 2212 7043 2232
tri 7043 2212 7063 2232 sw
tri 10163 2212 10183 2232 se
rect 10183 2212 10285 2232
tri 10285 2212 10305 2232 sw
tri 13405 2212 13425 2232 se
rect 13425 2212 13527 2232
tri 13527 2212 13547 2232 sw
tri 16647 2212 16667 2232 se
rect 16667 2212 16697 2232
rect 481 2188 579 2212
rect 481 2154 497 2188
rect 531 2154 579 2188
rect 481 2120 579 2154
rect 481 2086 497 2120
rect 531 2086 579 2120
rect 481 2062 579 2086
rect 3679 2188 3821 2212
rect 3679 2154 3738 2188
rect 3772 2154 3821 2188
rect 3679 2120 3821 2154
rect 3679 2086 3738 2120
rect 3772 2086 3821 2120
rect 3679 2062 3821 2086
rect 6921 2188 7063 2212
rect 6921 2154 6980 2188
rect 7014 2154 7063 2188
rect 6921 2120 7063 2154
rect 6921 2086 6980 2120
rect 7014 2086 7063 2120
rect 6921 2062 7063 2086
rect 10163 2190 10305 2212
rect 10163 2156 10222 2190
rect 10256 2156 10305 2190
rect 10163 2122 10305 2156
rect 10163 2088 10222 2122
rect 10256 2088 10305 2122
rect 10163 2062 10305 2088
rect 13405 2188 13547 2212
rect 13405 2154 13465 2188
rect 13499 2154 13547 2188
rect 13405 2120 13547 2154
rect 13405 2086 13465 2120
rect 13499 2086 13547 2120
rect 13405 2062 13547 2086
rect 16647 2062 16697 2212
rect 481 2042 559 2062
tri 559 2042 579 2062 nw
tri 3679 2042 3699 2062 ne
rect 3699 2042 3801 2062
tri 3801 2042 3821 2062 nw
tri 6921 2042 6941 2062 ne
rect 6941 2042 7043 2062
tri 7043 2042 7063 2062 nw
tri 10163 2042 10183 2062 ne
rect 10183 2042 10285 2062
tri 10285 2042 10305 2062 nw
tri 13405 2042 13425 2062 ne
rect 13425 2042 13527 2062
tri 13527 2042 13547 2062 nw
tri 16647 2042 16667 2062 ne
rect 16667 2042 16697 2062
rect 16739 2212 16769 2232
tri 16769 2212 16789 2232 sw
tri 19889 2212 19909 2232 se
rect 19909 2212 19987 2232
rect 16739 2062 16789 2212
rect 19889 2188 19987 2212
rect 19889 2154 19937 2188
rect 19971 2154 19987 2188
rect 19889 2120 19987 2154
rect 19889 2086 19937 2120
rect 19971 2086 19987 2120
rect 19889 2062 19987 2086
rect 16739 2042 16769 2062
tri 16769 2042 16789 2062 nw
tri 19889 2042 19909 2062 ne
rect 19909 2042 19987 2062
<< polycont >>
rect 497 2564 531 2598
rect 497 2496 531 2530
rect 3738 2566 3772 2600
rect 3738 2498 3772 2532
rect 6980 2566 7014 2600
rect 6980 2498 7014 2532
rect 10222 2564 10256 2598
rect 10222 2496 10256 2530
rect 13465 2564 13499 2598
rect 13465 2496 13499 2530
rect 19937 2566 19971 2600
rect 19937 2498 19971 2532
rect 497 2154 531 2188
rect 497 2086 531 2120
rect 3738 2154 3772 2188
rect 3738 2086 3772 2120
rect 6980 2154 7014 2188
rect 6980 2086 7014 2120
rect 10222 2156 10256 2190
rect 10222 2088 10256 2122
rect 13465 2154 13499 2188
rect 13465 2086 13499 2120
rect 19937 2154 19971 2188
rect 19937 2086 19971 2120
<< locali >>
rect 579 2774 679 2808
rect 713 2774 752 2808
rect 786 2774 825 2808
rect 859 2774 898 2808
rect 932 2774 971 2808
rect 1005 2774 1044 2808
rect 1078 2774 1117 2808
rect 1151 2774 1190 2808
rect 1224 2774 1263 2808
rect 1297 2774 1336 2808
rect 1370 2774 1409 2808
rect 1443 2774 1482 2808
rect 1516 2774 1555 2808
rect 1589 2774 1628 2808
rect 1662 2774 1701 2808
rect 1735 2774 1774 2808
rect 1808 2774 1847 2808
rect 1881 2774 1920 2808
rect 1954 2774 1993 2808
rect 2027 2774 2066 2808
rect 2100 2774 2139 2808
rect 2173 2774 2213 2808
rect 2247 2774 2287 2808
rect 2321 2774 2361 2808
rect 2395 2774 2435 2808
rect 2469 2774 2509 2808
rect 2543 2774 2583 2808
rect 2617 2774 2657 2808
rect 2691 2774 2731 2808
rect 2765 2774 2805 2808
rect 2839 2774 2879 2808
rect 2913 2774 2953 2808
rect 2987 2774 3027 2808
rect 3061 2774 3101 2808
rect 3135 2774 3175 2808
rect 3209 2774 3249 2808
rect 3283 2774 3323 2808
rect 3357 2774 3397 2808
rect 3431 2774 3471 2808
rect 3505 2774 3545 2808
rect 3579 2774 3679 2808
rect 579 2736 3679 2774
rect 579 2702 679 2736
rect 713 2702 752 2736
rect 786 2702 825 2736
rect 859 2702 898 2736
rect 932 2702 971 2736
rect 1005 2702 1044 2736
rect 1078 2702 1117 2736
rect 1151 2702 1190 2736
rect 1224 2702 1263 2736
rect 1297 2702 1336 2736
rect 1370 2702 1409 2736
rect 1443 2702 1482 2736
rect 1516 2702 1555 2736
rect 1589 2702 1628 2736
rect 1662 2702 1701 2736
rect 1735 2702 1774 2736
rect 1808 2702 1847 2736
rect 1881 2702 1920 2736
rect 1954 2702 1993 2736
rect 2027 2702 2066 2736
rect 2100 2702 2139 2736
rect 2173 2702 2213 2736
rect 2247 2702 2287 2736
rect 2321 2702 2361 2736
rect 2395 2702 2435 2736
rect 2469 2702 2509 2736
rect 2543 2702 2583 2736
rect 2617 2702 2657 2736
rect 2691 2702 2731 2736
rect 2765 2702 2805 2736
rect 2839 2702 2879 2736
rect 2913 2702 2953 2736
rect 2987 2702 3027 2736
rect 3061 2702 3101 2736
rect 3135 2702 3175 2736
rect 3209 2702 3249 2736
rect 3283 2702 3323 2736
rect 3357 2702 3397 2736
rect 3431 2702 3471 2736
rect 3505 2702 3545 2736
rect 3579 2702 3679 2736
rect 3821 2774 3921 2808
rect 3955 2774 3995 2808
rect 4029 2774 4069 2808
rect 4103 2774 4143 2808
rect 4177 2774 4217 2808
rect 4251 2774 4291 2808
rect 4325 2774 4365 2808
rect 4399 2774 4439 2808
rect 4473 2774 4513 2808
rect 4547 2774 4587 2808
rect 4621 2774 4661 2808
rect 4695 2774 4735 2808
rect 4769 2774 4809 2808
rect 4843 2774 4883 2808
rect 4917 2774 4957 2808
rect 4991 2774 5031 2808
rect 5065 2774 5105 2808
rect 5139 2774 5179 2808
rect 5213 2774 5253 2808
rect 5287 2774 5327 2808
rect 5361 2774 5400 2808
rect 5434 2774 5473 2808
rect 5507 2774 5546 2808
rect 5580 2774 5619 2808
rect 5653 2774 5692 2808
rect 5726 2774 5765 2808
rect 5799 2774 5838 2808
rect 5872 2774 5911 2808
rect 5945 2774 5984 2808
rect 6018 2774 6057 2808
rect 6091 2774 6130 2808
rect 6164 2774 6203 2808
rect 6237 2774 6276 2808
rect 6310 2774 6349 2808
rect 6383 2774 6422 2808
rect 6456 2774 6495 2808
rect 6529 2774 6568 2808
rect 6602 2774 6641 2808
rect 6675 2774 6714 2808
rect 6748 2774 6787 2808
rect 6821 2774 6921 2808
rect 3821 2736 6921 2774
rect 3821 2702 3921 2736
rect 3955 2702 3995 2736
rect 4029 2702 4069 2736
rect 4103 2702 4143 2736
rect 4177 2702 4217 2736
rect 4251 2702 4291 2736
rect 4325 2702 4365 2736
rect 4399 2702 4439 2736
rect 4473 2702 4513 2736
rect 4547 2702 4587 2736
rect 4621 2702 4661 2736
rect 4695 2702 4735 2736
rect 4769 2702 4809 2736
rect 4843 2702 4883 2736
rect 4917 2702 4957 2736
rect 4991 2702 5031 2736
rect 5065 2702 5105 2736
rect 5139 2702 5179 2736
rect 5213 2702 5253 2736
rect 5287 2702 5327 2736
rect 5361 2702 5400 2736
rect 5434 2702 5473 2736
rect 5507 2702 5546 2736
rect 5580 2702 5619 2736
rect 5653 2702 5692 2736
rect 5726 2702 5765 2736
rect 5799 2702 5838 2736
rect 5872 2702 5911 2736
rect 5945 2702 5984 2736
rect 6018 2702 6057 2736
rect 6091 2702 6130 2736
rect 6164 2702 6203 2736
rect 6237 2702 6276 2736
rect 6310 2702 6349 2736
rect 6383 2702 6422 2736
rect 6456 2702 6495 2736
rect 6529 2702 6568 2736
rect 6602 2702 6641 2736
rect 6675 2702 6714 2736
rect 6748 2702 6787 2736
rect 6821 2702 6921 2736
rect 7063 2774 7163 2808
rect 7197 2774 7236 2808
rect 7270 2774 7309 2808
rect 7343 2774 7382 2808
rect 7416 2774 7455 2808
rect 7489 2774 7528 2808
rect 7562 2774 7601 2808
rect 7635 2774 7674 2808
rect 7708 2774 7747 2808
rect 7781 2774 7820 2808
rect 7854 2774 7893 2808
rect 7927 2774 7966 2808
rect 8000 2774 8039 2808
rect 8073 2774 8112 2808
rect 8146 2774 8185 2808
rect 8219 2774 8258 2808
rect 8292 2774 8331 2808
rect 8365 2774 8404 2808
rect 8438 2774 8477 2808
rect 8511 2774 8550 2808
rect 8584 2774 8623 2808
rect 8657 2774 8697 2808
rect 8731 2774 8771 2808
rect 8805 2774 8845 2808
rect 8879 2774 8919 2808
rect 8953 2774 8993 2808
rect 9027 2774 9067 2808
rect 9101 2774 9141 2808
rect 9175 2774 9215 2808
rect 9249 2774 9289 2808
rect 9323 2774 9363 2808
rect 9397 2774 9437 2808
rect 9471 2774 9511 2808
rect 9545 2774 9585 2808
rect 9619 2774 9659 2808
rect 9693 2774 9733 2808
rect 9767 2774 9807 2808
rect 9841 2774 9881 2808
rect 9915 2774 9955 2808
rect 9989 2774 10029 2808
rect 10063 2774 10163 2808
rect 7063 2736 10163 2774
rect 7063 2702 7163 2736
rect 7197 2702 7236 2736
rect 7270 2702 7309 2736
rect 7343 2702 7382 2736
rect 7416 2702 7455 2736
rect 7489 2702 7528 2736
rect 7562 2702 7601 2736
rect 7635 2702 7674 2736
rect 7708 2702 7747 2736
rect 7781 2702 7820 2736
rect 7854 2702 7893 2736
rect 7927 2702 7966 2736
rect 8000 2702 8039 2736
rect 8073 2702 8112 2736
rect 8146 2702 8185 2736
rect 8219 2702 8258 2736
rect 8292 2702 8331 2736
rect 8365 2702 8404 2736
rect 8438 2702 8477 2736
rect 8511 2702 8550 2736
rect 8584 2702 8623 2736
rect 8657 2702 8697 2736
rect 8731 2702 8771 2736
rect 8805 2702 8845 2736
rect 8879 2702 8919 2736
rect 8953 2702 8993 2736
rect 9027 2702 9067 2736
rect 9101 2702 9141 2736
rect 9175 2702 9215 2736
rect 9249 2702 9289 2736
rect 9323 2702 9363 2736
rect 9397 2702 9437 2736
rect 9471 2702 9511 2736
rect 9545 2702 9585 2736
rect 9619 2702 9659 2736
rect 9693 2702 9733 2736
rect 9767 2702 9807 2736
rect 9841 2702 9881 2736
rect 9915 2702 9955 2736
rect 9989 2702 10029 2736
rect 10063 2702 10163 2736
rect 10305 2774 10405 2808
rect 10439 2774 10479 2808
rect 10513 2774 10553 2808
rect 10587 2774 10627 2808
rect 10661 2774 10701 2808
rect 10735 2774 10775 2808
rect 10809 2774 10849 2808
rect 10883 2774 10923 2808
rect 10957 2774 10997 2808
rect 11031 2774 11071 2808
rect 11105 2774 11145 2808
rect 11179 2774 11219 2808
rect 11253 2774 11293 2808
rect 11327 2774 11367 2808
rect 11401 2774 11441 2808
rect 11475 2774 11515 2808
rect 11549 2774 11589 2808
rect 11623 2774 11663 2808
rect 11697 2774 11737 2808
rect 11771 2774 11811 2808
rect 11845 2774 11884 2808
rect 11918 2774 11957 2808
rect 11991 2774 12030 2808
rect 12064 2774 12103 2808
rect 12137 2774 12176 2808
rect 12210 2774 12249 2808
rect 12283 2774 12322 2808
rect 12356 2774 12395 2808
rect 12429 2774 12468 2808
rect 12502 2774 12541 2808
rect 12575 2774 12614 2808
rect 12648 2774 12687 2808
rect 12721 2774 12760 2808
rect 12794 2774 12833 2808
rect 12867 2774 12906 2808
rect 12940 2774 12979 2808
rect 13013 2774 13052 2808
rect 13086 2774 13125 2808
rect 13159 2774 13198 2808
rect 13232 2774 13271 2808
rect 13305 2774 13405 2808
rect 10305 2736 13405 2774
rect 10305 2702 10405 2736
rect 10439 2702 10479 2736
rect 10513 2702 10553 2736
rect 10587 2702 10627 2736
rect 10661 2702 10701 2736
rect 10735 2702 10775 2736
rect 10809 2702 10849 2736
rect 10883 2702 10923 2736
rect 10957 2702 10997 2736
rect 11031 2702 11071 2736
rect 11105 2702 11145 2736
rect 11179 2702 11219 2736
rect 11253 2702 11293 2736
rect 11327 2702 11367 2736
rect 11401 2702 11441 2736
rect 11475 2702 11515 2736
rect 11549 2702 11589 2736
rect 11623 2702 11663 2736
rect 11697 2702 11737 2736
rect 11771 2702 11811 2736
rect 11845 2702 11884 2736
rect 11918 2702 11957 2736
rect 11991 2702 12030 2736
rect 12064 2702 12103 2736
rect 12137 2702 12176 2736
rect 12210 2702 12249 2736
rect 12283 2702 12322 2736
rect 12356 2702 12395 2736
rect 12429 2702 12468 2736
rect 12502 2702 12541 2736
rect 12575 2702 12614 2736
rect 12648 2702 12687 2736
rect 12721 2702 12760 2736
rect 12794 2702 12833 2736
rect 12867 2702 12906 2736
rect 12940 2702 12979 2736
rect 13013 2702 13052 2736
rect 13086 2702 13125 2736
rect 13159 2702 13198 2736
rect 13232 2702 13271 2736
rect 13305 2702 13405 2736
rect 13547 2774 13647 2808
rect 13681 2774 13720 2808
rect 13754 2774 13793 2808
rect 13827 2774 13866 2808
rect 13900 2774 13939 2808
rect 13973 2774 14012 2808
rect 14046 2774 14085 2808
rect 14119 2774 14158 2808
rect 14192 2774 14231 2808
rect 14265 2774 14304 2808
rect 14338 2774 14377 2808
rect 14411 2774 14450 2808
rect 14484 2774 14523 2808
rect 14557 2774 14596 2808
rect 14630 2774 14669 2808
rect 14703 2774 14742 2808
rect 14776 2774 14815 2808
rect 14849 2774 14888 2808
rect 14922 2774 14961 2808
rect 14995 2774 15034 2808
rect 15068 2774 15107 2808
rect 15141 2774 15181 2808
rect 15215 2774 15255 2808
rect 15289 2774 15329 2808
rect 15363 2774 15403 2808
rect 15437 2774 15477 2808
rect 15511 2774 15551 2808
rect 15585 2774 15625 2808
rect 15659 2774 15699 2808
rect 15733 2774 15773 2808
rect 15807 2774 15847 2808
rect 15881 2774 15921 2808
rect 15955 2774 15995 2808
rect 16029 2774 16069 2808
rect 16103 2774 16143 2808
rect 16177 2774 16217 2808
rect 16251 2774 16291 2808
rect 16325 2774 16365 2808
rect 16399 2774 16439 2808
rect 16473 2774 16513 2808
rect 16547 2774 16647 2808
rect 13547 2736 16647 2774
rect 13547 2702 13647 2736
rect 13681 2702 13720 2736
rect 13754 2702 13793 2736
rect 13827 2702 13866 2736
rect 13900 2702 13939 2736
rect 13973 2702 14012 2736
rect 14046 2702 14085 2736
rect 14119 2702 14158 2736
rect 14192 2702 14231 2736
rect 14265 2702 14304 2736
rect 14338 2702 14377 2736
rect 14411 2702 14450 2736
rect 14484 2702 14523 2736
rect 14557 2702 14596 2736
rect 14630 2702 14669 2736
rect 14703 2702 14742 2736
rect 14776 2702 14815 2736
rect 14849 2702 14888 2736
rect 14922 2702 14961 2736
rect 14995 2702 15034 2736
rect 15068 2702 15107 2736
rect 15141 2702 15181 2736
rect 15215 2702 15255 2736
rect 15289 2702 15329 2736
rect 15363 2702 15403 2736
rect 15437 2702 15477 2736
rect 15511 2702 15551 2736
rect 15585 2702 15625 2736
rect 15659 2702 15699 2736
rect 15733 2702 15773 2736
rect 15807 2702 15847 2736
rect 15881 2702 15921 2736
rect 15955 2702 15995 2736
rect 16029 2702 16069 2736
rect 16103 2702 16143 2736
rect 16177 2702 16217 2736
rect 16251 2702 16291 2736
rect 16325 2702 16365 2736
rect 16399 2702 16439 2736
rect 16473 2702 16513 2736
rect 16547 2702 16647 2736
rect 16789 2774 16889 2808
rect 16923 2774 16963 2808
rect 16997 2774 17037 2808
rect 17071 2774 17111 2808
rect 17145 2774 17185 2808
rect 17219 2774 17259 2808
rect 17293 2774 17333 2808
rect 17367 2774 17407 2808
rect 17441 2774 17481 2808
rect 17515 2774 17555 2808
rect 17589 2774 17629 2808
rect 17663 2774 17703 2808
rect 17737 2774 17777 2808
rect 17811 2774 17851 2808
rect 17885 2774 17925 2808
rect 17959 2774 17999 2808
rect 18033 2774 18073 2808
rect 18107 2774 18147 2808
rect 18181 2774 18221 2808
rect 18255 2774 18295 2808
rect 18329 2774 18368 2808
rect 18402 2774 18441 2808
rect 18475 2774 18514 2808
rect 18548 2774 18587 2808
rect 18621 2774 18660 2808
rect 18694 2774 18733 2808
rect 18767 2774 18806 2808
rect 18840 2774 18879 2808
rect 18913 2774 18952 2808
rect 18986 2774 19025 2808
rect 19059 2774 19098 2808
rect 19132 2774 19171 2808
rect 19205 2774 19244 2808
rect 19278 2774 19317 2808
rect 19351 2774 19390 2808
rect 19424 2774 19463 2808
rect 19497 2774 19536 2808
rect 19570 2774 19609 2808
rect 19643 2774 19682 2808
rect 19716 2774 19755 2808
rect 19789 2774 19889 2808
rect 16789 2736 19889 2774
rect 16789 2702 16889 2736
rect 16923 2702 16963 2736
rect 16997 2702 17037 2736
rect 17071 2702 17111 2736
rect 17145 2702 17185 2736
rect 17219 2702 17259 2736
rect 17293 2702 17333 2736
rect 17367 2702 17407 2736
rect 17441 2702 17481 2736
rect 17515 2702 17555 2736
rect 17589 2702 17629 2736
rect 17663 2702 17703 2736
rect 17737 2702 17777 2736
rect 17811 2702 17851 2736
rect 17885 2702 17925 2736
rect 17959 2702 17999 2736
rect 18033 2702 18073 2736
rect 18107 2702 18147 2736
rect 18181 2702 18221 2736
rect 18255 2702 18295 2736
rect 18329 2702 18368 2736
rect 18402 2702 18441 2736
rect 18475 2702 18514 2736
rect 18548 2702 18587 2736
rect 18621 2702 18660 2736
rect 18694 2702 18733 2736
rect 18767 2702 18806 2736
rect 18840 2702 18879 2736
rect 18913 2702 18952 2736
rect 18986 2702 19025 2736
rect 19059 2702 19098 2736
rect 19132 2702 19171 2736
rect 19205 2702 19244 2736
rect 19278 2702 19317 2736
rect 19351 2702 19390 2736
rect 19424 2702 19463 2736
rect 19497 2702 19536 2736
rect 19570 2702 19609 2736
rect 19643 2702 19682 2736
rect 19716 2702 19755 2736
rect 19789 2702 19889 2736
rect 3738 2614 3772 2616
rect 6980 2614 7014 2616
rect 517 2598 555 2614
rect 531 2580 555 2598
rect 3735 2600 3773 2614
rect 3735 2580 3738 2600
rect 497 2530 531 2564
rect 497 2480 531 2496
rect 3772 2580 3773 2600
rect 6977 2600 7015 2614
rect 6977 2580 6980 2600
rect 3738 2532 3772 2566
rect 3738 2482 3772 2498
rect 7014 2580 7015 2600
rect 10219 2598 10257 2614
rect 10219 2580 10222 2598
rect 6980 2532 7014 2566
rect 6980 2482 7014 2498
rect 10256 2580 10257 2598
rect 13485 2598 13523 2614
rect 13499 2580 13523 2598
rect 19937 2603 19971 2616
rect 10222 2530 10256 2564
rect 10222 2480 10256 2496
rect 13465 2530 13499 2564
rect 13465 2480 13499 2496
rect 19937 2532 19971 2566
rect 19937 2482 19971 2497
rect 579 2362 679 2396
rect 713 2362 752 2396
rect 786 2362 825 2396
rect 859 2362 898 2396
rect 932 2362 971 2396
rect 1005 2362 1044 2396
rect 1078 2362 1117 2396
rect 1151 2362 1190 2396
rect 1224 2362 1263 2396
rect 1297 2362 1336 2396
rect 1370 2362 1409 2396
rect 1443 2362 1482 2396
rect 1516 2362 1555 2396
rect 1589 2362 1628 2396
rect 1662 2362 1701 2396
rect 1735 2362 1774 2396
rect 1808 2362 1847 2396
rect 1881 2362 1920 2396
rect 1954 2362 1993 2396
rect 2027 2362 2066 2396
rect 2100 2362 2139 2396
rect 2173 2362 2213 2396
rect 2247 2362 2287 2396
rect 2321 2362 2361 2396
rect 2395 2362 2435 2396
rect 2469 2362 2509 2396
rect 2543 2362 2583 2396
rect 2617 2362 2657 2396
rect 2691 2362 2731 2396
rect 2765 2362 2805 2396
rect 2839 2362 2879 2396
rect 2913 2362 2953 2396
rect 2987 2362 3027 2396
rect 3061 2362 3101 2396
rect 3135 2362 3175 2396
rect 3209 2362 3249 2396
rect 3283 2362 3323 2396
rect 3357 2362 3397 2396
rect 3431 2362 3471 2396
rect 3505 2362 3545 2396
rect 3579 2362 3679 2396
rect 579 2324 3679 2362
rect 579 2290 679 2324
rect 713 2290 752 2324
rect 786 2290 825 2324
rect 859 2290 898 2324
rect 932 2290 971 2324
rect 1005 2290 1044 2324
rect 1078 2290 1117 2324
rect 1151 2290 1190 2324
rect 1224 2290 1263 2324
rect 1297 2290 1336 2324
rect 1370 2290 1409 2324
rect 1443 2290 1482 2324
rect 1516 2290 1555 2324
rect 1589 2290 1628 2324
rect 1662 2290 1701 2324
rect 1735 2290 1774 2324
rect 1808 2290 1847 2324
rect 1881 2290 1920 2324
rect 1954 2290 1993 2324
rect 2027 2290 2066 2324
rect 2100 2290 2139 2324
rect 2173 2290 2213 2324
rect 2247 2290 2287 2324
rect 2321 2290 2361 2324
rect 2395 2290 2435 2324
rect 2469 2290 2509 2324
rect 2543 2290 2583 2324
rect 2617 2290 2657 2324
rect 2691 2290 2731 2324
rect 2765 2290 2805 2324
rect 2839 2290 2879 2324
rect 2913 2290 2953 2324
rect 2987 2290 3027 2324
rect 3061 2290 3101 2324
rect 3135 2290 3175 2324
rect 3209 2290 3249 2324
rect 3283 2290 3323 2324
rect 3357 2290 3397 2324
rect 3431 2290 3471 2324
rect 3505 2290 3545 2324
rect 3579 2290 3679 2324
rect 3821 2362 3921 2396
rect 3955 2362 3995 2396
rect 4029 2362 4069 2396
rect 4103 2362 4143 2396
rect 4177 2362 4217 2396
rect 4251 2362 4291 2396
rect 4325 2362 4365 2396
rect 4399 2362 4439 2396
rect 4473 2362 4513 2396
rect 4547 2362 4587 2396
rect 4621 2362 4661 2396
rect 4695 2362 4735 2396
rect 4769 2362 4809 2396
rect 4843 2362 4883 2396
rect 4917 2362 4957 2396
rect 4991 2362 5031 2396
rect 5065 2362 5105 2396
rect 5139 2362 5179 2396
rect 5213 2362 5253 2396
rect 5287 2362 5327 2396
rect 5361 2362 5400 2396
rect 5434 2362 5473 2396
rect 5507 2362 5546 2396
rect 5580 2362 5619 2396
rect 5653 2362 5692 2396
rect 5726 2362 5765 2396
rect 5799 2362 5838 2396
rect 5872 2362 5911 2396
rect 5945 2362 5984 2396
rect 6018 2362 6057 2396
rect 6091 2362 6130 2396
rect 6164 2362 6203 2396
rect 6237 2362 6276 2396
rect 6310 2362 6349 2396
rect 6383 2362 6422 2396
rect 6456 2362 6495 2396
rect 6529 2362 6568 2396
rect 6602 2362 6641 2396
rect 6675 2362 6714 2396
rect 6748 2362 6787 2396
rect 6821 2362 6921 2396
rect 3821 2324 6921 2362
rect 3821 2290 3921 2324
rect 3955 2290 3995 2324
rect 4029 2290 4069 2324
rect 4103 2290 4143 2324
rect 4177 2290 4217 2324
rect 4251 2290 4291 2324
rect 4325 2290 4365 2324
rect 4399 2290 4439 2324
rect 4473 2290 4513 2324
rect 4547 2290 4587 2324
rect 4621 2290 4661 2324
rect 4695 2290 4735 2324
rect 4769 2290 4809 2324
rect 4843 2290 4883 2324
rect 4917 2290 4957 2324
rect 4991 2290 5031 2324
rect 5065 2290 5105 2324
rect 5139 2290 5179 2324
rect 5213 2290 5253 2324
rect 5287 2290 5327 2324
rect 5361 2290 5400 2324
rect 5434 2290 5473 2324
rect 5507 2290 5546 2324
rect 5580 2290 5619 2324
rect 5653 2290 5692 2324
rect 5726 2290 5765 2324
rect 5799 2290 5838 2324
rect 5872 2290 5911 2324
rect 5945 2290 5984 2324
rect 6018 2290 6057 2324
rect 6091 2290 6130 2324
rect 6164 2290 6203 2324
rect 6237 2290 6276 2324
rect 6310 2290 6349 2324
rect 6383 2290 6422 2324
rect 6456 2290 6495 2324
rect 6529 2290 6568 2324
rect 6602 2290 6641 2324
rect 6675 2290 6714 2324
rect 6748 2290 6787 2324
rect 6821 2290 6921 2324
rect 7063 2362 7163 2396
rect 7197 2362 7236 2396
rect 7270 2362 7309 2396
rect 7343 2362 7382 2396
rect 7416 2362 7455 2396
rect 7489 2362 7528 2396
rect 7562 2362 7601 2396
rect 7635 2362 7674 2396
rect 7708 2362 7747 2396
rect 7781 2362 7820 2396
rect 7854 2362 7893 2396
rect 7927 2362 7966 2396
rect 8000 2362 8039 2396
rect 8073 2362 8112 2396
rect 8146 2362 8185 2396
rect 8219 2362 8258 2396
rect 8292 2362 8331 2396
rect 8365 2362 8404 2396
rect 8438 2362 8477 2396
rect 8511 2362 8550 2396
rect 8584 2362 8623 2396
rect 8657 2362 8697 2396
rect 8731 2362 8771 2396
rect 8805 2362 8845 2396
rect 8879 2362 8919 2396
rect 8953 2362 8993 2396
rect 9027 2362 9067 2396
rect 9101 2362 9141 2396
rect 9175 2362 9215 2396
rect 9249 2362 9289 2396
rect 9323 2362 9363 2396
rect 9397 2362 9437 2396
rect 9471 2362 9511 2396
rect 9545 2362 9585 2396
rect 9619 2362 9659 2396
rect 9693 2362 9733 2396
rect 9767 2362 9807 2396
rect 9841 2362 9881 2396
rect 9915 2362 9955 2396
rect 9989 2362 10029 2396
rect 10063 2362 10163 2396
rect 7063 2324 10163 2362
rect 7063 2290 7163 2324
rect 7197 2290 7236 2324
rect 7270 2290 7309 2324
rect 7343 2290 7382 2324
rect 7416 2290 7455 2324
rect 7489 2290 7528 2324
rect 7562 2290 7601 2324
rect 7635 2290 7674 2324
rect 7708 2290 7747 2324
rect 7781 2290 7820 2324
rect 7854 2290 7893 2324
rect 7927 2290 7966 2324
rect 8000 2290 8039 2324
rect 8073 2290 8112 2324
rect 8146 2290 8185 2324
rect 8219 2290 8258 2324
rect 8292 2290 8331 2324
rect 8365 2290 8404 2324
rect 8438 2290 8477 2324
rect 8511 2290 8550 2324
rect 8584 2290 8623 2324
rect 8657 2290 8697 2324
rect 8731 2290 8771 2324
rect 8805 2290 8845 2324
rect 8879 2290 8919 2324
rect 8953 2290 8993 2324
rect 9027 2290 9067 2324
rect 9101 2290 9141 2324
rect 9175 2290 9215 2324
rect 9249 2290 9289 2324
rect 9323 2290 9363 2324
rect 9397 2290 9437 2324
rect 9471 2290 9511 2324
rect 9545 2290 9585 2324
rect 9619 2290 9659 2324
rect 9693 2290 9733 2324
rect 9767 2290 9807 2324
rect 9841 2290 9881 2324
rect 9915 2290 9955 2324
rect 9989 2290 10029 2324
rect 10063 2290 10163 2324
rect 10305 2362 10405 2396
rect 10439 2362 10479 2396
rect 10513 2362 10553 2396
rect 10587 2362 10627 2396
rect 10661 2362 10701 2396
rect 10735 2362 10775 2396
rect 10809 2362 10849 2396
rect 10883 2362 10923 2396
rect 10957 2362 10997 2396
rect 11031 2362 11071 2396
rect 11105 2362 11145 2396
rect 11179 2362 11219 2396
rect 11253 2362 11293 2396
rect 11327 2362 11367 2396
rect 11401 2362 11441 2396
rect 11475 2362 11515 2396
rect 11549 2362 11589 2396
rect 11623 2362 11663 2396
rect 11697 2362 11737 2396
rect 11771 2362 11811 2396
rect 11845 2362 11884 2396
rect 11918 2362 11957 2396
rect 11991 2362 12030 2396
rect 12064 2362 12103 2396
rect 12137 2362 12176 2396
rect 12210 2362 12249 2396
rect 12283 2362 12322 2396
rect 12356 2362 12395 2396
rect 12429 2362 12468 2396
rect 12502 2362 12541 2396
rect 12575 2362 12614 2396
rect 12648 2362 12687 2396
rect 12721 2362 12760 2396
rect 12794 2362 12833 2396
rect 12867 2362 12906 2396
rect 12940 2362 12979 2396
rect 13013 2362 13052 2396
rect 13086 2362 13125 2396
rect 13159 2362 13198 2396
rect 13232 2362 13271 2396
rect 13305 2362 13405 2396
rect 10305 2324 13405 2362
rect 10305 2290 10405 2324
rect 10439 2290 10479 2324
rect 10513 2290 10553 2324
rect 10587 2290 10627 2324
rect 10661 2290 10701 2324
rect 10735 2290 10775 2324
rect 10809 2290 10849 2324
rect 10883 2290 10923 2324
rect 10957 2290 10997 2324
rect 11031 2290 11071 2324
rect 11105 2290 11145 2324
rect 11179 2290 11219 2324
rect 11253 2290 11293 2324
rect 11327 2290 11367 2324
rect 11401 2290 11441 2324
rect 11475 2290 11515 2324
rect 11549 2290 11589 2324
rect 11623 2290 11663 2324
rect 11697 2290 11737 2324
rect 11771 2290 11811 2324
rect 11845 2290 11884 2324
rect 11918 2290 11957 2324
rect 11991 2290 12030 2324
rect 12064 2290 12103 2324
rect 12137 2290 12176 2324
rect 12210 2290 12249 2324
rect 12283 2290 12322 2324
rect 12356 2290 12395 2324
rect 12429 2290 12468 2324
rect 12502 2290 12541 2324
rect 12575 2290 12614 2324
rect 12648 2290 12687 2324
rect 12721 2290 12760 2324
rect 12794 2290 12833 2324
rect 12867 2290 12906 2324
rect 12940 2290 12979 2324
rect 13013 2290 13052 2324
rect 13086 2290 13125 2324
rect 13159 2290 13198 2324
rect 13232 2290 13271 2324
rect 13305 2290 13405 2324
rect 13547 2362 13647 2396
rect 13681 2362 13720 2396
rect 13754 2362 13793 2396
rect 13827 2362 13866 2396
rect 13900 2362 13939 2396
rect 13973 2362 14012 2396
rect 14046 2362 14085 2396
rect 14119 2362 14158 2396
rect 14192 2362 14231 2396
rect 14265 2362 14304 2396
rect 14338 2362 14377 2396
rect 14411 2362 14450 2396
rect 14484 2362 14523 2396
rect 14557 2362 14596 2396
rect 14630 2362 14669 2396
rect 14703 2362 14742 2396
rect 14776 2362 14815 2396
rect 14849 2362 14888 2396
rect 14922 2362 14961 2396
rect 14995 2362 15034 2396
rect 15068 2362 15107 2396
rect 15141 2362 15181 2396
rect 15215 2362 15255 2396
rect 15289 2362 15329 2396
rect 15363 2362 15403 2396
rect 15437 2362 15477 2396
rect 15511 2362 15551 2396
rect 15585 2362 15625 2396
rect 15659 2362 15699 2396
rect 15733 2362 15773 2396
rect 15807 2362 15847 2396
rect 15881 2362 15921 2396
rect 15955 2362 15995 2396
rect 16029 2362 16069 2396
rect 16103 2362 16143 2396
rect 16177 2362 16217 2396
rect 16251 2362 16291 2396
rect 16325 2362 16365 2396
rect 16399 2362 16439 2396
rect 16473 2362 16513 2396
rect 16547 2362 16647 2396
rect 13547 2324 16647 2362
rect 13547 2290 13647 2324
rect 13681 2290 13720 2324
rect 13754 2290 13793 2324
rect 13827 2290 13866 2324
rect 13900 2290 13939 2324
rect 13973 2290 14012 2324
rect 14046 2290 14085 2324
rect 14119 2290 14158 2324
rect 14192 2290 14231 2324
rect 14265 2290 14304 2324
rect 14338 2290 14377 2324
rect 14411 2290 14450 2324
rect 14484 2290 14523 2324
rect 14557 2290 14596 2324
rect 14630 2290 14669 2324
rect 14703 2290 14742 2324
rect 14776 2290 14815 2324
rect 14849 2290 14888 2324
rect 14922 2290 14961 2324
rect 14995 2290 15034 2324
rect 15068 2290 15107 2324
rect 15141 2290 15181 2324
rect 15215 2290 15255 2324
rect 15289 2290 15329 2324
rect 15363 2290 15403 2324
rect 15437 2290 15477 2324
rect 15511 2290 15551 2324
rect 15585 2290 15625 2324
rect 15659 2290 15699 2324
rect 15733 2290 15773 2324
rect 15807 2290 15847 2324
rect 15881 2290 15921 2324
rect 15955 2290 15995 2324
rect 16029 2290 16069 2324
rect 16103 2290 16143 2324
rect 16177 2290 16217 2324
rect 16251 2290 16291 2324
rect 16325 2290 16365 2324
rect 16399 2290 16439 2324
rect 16473 2290 16513 2324
rect 16547 2290 16647 2324
rect 16789 2362 16889 2396
rect 16923 2362 16963 2396
rect 16997 2362 17037 2396
rect 17071 2362 17111 2396
rect 17145 2362 17185 2396
rect 17219 2362 17259 2396
rect 17293 2362 17333 2396
rect 17367 2362 17407 2396
rect 17441 2362 17481 2396
rect 17515 2362 17555 2396
rect 17589 2362 17629 2396
rect 17663 2362 17703 2396
rect 17737 2362 17777 2396
rect 17811 2362 17851 2396
rect 17885 2362 17925 2396
rect 17959 2362 17999 2396
rect 18033 2362 18073 2396
rect 18107 2362 18147 2396
rect 18181 2362 18221 2396
rect 18255 2362 18295 2396
rect 18329 2362 18368 2396
rect 18402 2362 18441 2396
rect 18475 2362 18514 2396
rect 18548 2362 18587 2396
rect 18621 2362 18660 2396
rect 18694 2362 18733 2396
rect 18767 2362 18806 2396
rect 18840 2362 18879 2396
rect 18913 2362 18952 2396
rect 18986 2362 19025 2396
rect 19059 2362 19098 2396
rect 19132 2362 19171 2396
rect 19205 2362 19244 2396
rect 19278 2362 19317 2396
rect 19351 2362 19390 2396
rect 19424 2362 19463 2396
rect 19497 2362 19536 2396
rect 19570 2362 19609 2396
rect 19643 2362 19682 2396
rect 19716 2362 19755 2396
rect 19789 2362 19889 2396
rect 16789 2324 19889 2362
rect 16789 2290 16889 2324
rect 16923 2290 16963 2324
rect 16997 2290 17037 2324
rect 17071 2290 17111 2324
rect 17145 2290 17185 2324
rect 17219 2290 17259 2324
rect 17293 2290 17333 2324
rect 17367 2290 17407 2324
rect 17441 2290 17481 2324
rect 17515 2290 17555 2324
rect 17589 2290 17629 2324
rect 17663 2290 17703 2324
rect 17737 2290 17777 2324
rect 17811 2290 17851 2324
rect 17885 2290 17925 2324
rect 17959 2290 17999 2324
rect 18033 2290 18073 2324
rect 18107 2290 18147 2324
rect 18181 2290 18221 2324
rect 18255 2290 18295 2324
rect 18329 2290 18368 2324
rect 18402 2290 18441 2324
rect 18475 2290 18514 2324
rect 18548 2290 18587 2324
rect 18621 2290 18660 2324
rect 18694 2290 18733 2324
rect 18767 2290 18806 2324
rect 18840 2290 18879 2324
rect 18913 2290 18952 2324
rect 18986 2290 19025 2324
rect 19059 2290 19098 2324
rect 19132 2290 19171 2324
rect 19205 2290 19244 2324
rect 19278 2290 19317 2324
rect 19351 2290 19390 2324
rect 19424 2290 19463 2324
rect 19497 2290 19536 2324
rect 19570 2290 19609 2324
rect 19643 2290 19682 2324
rect 19716 2290 19755 2324
rect 19789 2290 19889 2324
rect 497 2188 531 2204
rect 497 2120 531 2154
rect 3738 2188 3772 2204
rect 3738 2120 3772 2154
rect 531 2086 555 2106
rect 517 2072 555 2086
rect 3735 2086 3738 2106
rect 6980 2188 7014 2204
rect 6980 2120 7014 2154
rect 3772 2086 3773 2106
rect 3735 2072 3773 2086
rect 6977 2086 6980 2106
rect 10222 2190 10256 2206
rect 10222 2122 10256 2156
rect 7014 2086 7015 2106
rect 6977 2072 7015 2086
rect 10219 2088 10222 2106
rect 13465 2188 13499 2204
rect 13465 2120 13499 2154
rect 19937 2191 19971 2204
rect 19937 2120 19971 2154
rect 10256 2088 10257 2106
rect 10219 2072 10257 2088
rect 13499 2086 13523 2106
rect 13485 2072 13523 2086
rect 497 2070 531 2072
rect 3738 2070 3772 2072
rect 6980 2070 7014 2072
rect 13465 2070 13499 2072
rect 19937 2070 19971 2085
rect 579 1950 679 1984
rect 713 1950 752 1984
rect 786 1950 825 1984
rect 859 1950 898 1984
rect 932 1950 971 1984
rect 1005 1950 1044 1984
rect 1078 1950 1117 1984
rect 1151 1950 1190 1984
rect 1224 1950 1263 1984
rect 1297 1950 1336 1984
rect 1370 1950 1409 1984
rect 1443 1950 1482 1984
rect 1516 1950 1555 1984
rect 1589 1950 1628 1984
rect 1662 1950 1701 1984
rect 1735 1950 1774 1984
rect 1808 1950 1847 1984
rect 1881 1950 1920 1984
rect 1954 1950 1993 1984
rect 2027 1950 2066 1984
rect 2100 1950 2139 1984
rect 2173 1950 2213 1984
rect 2247 1950 2287 1984
rect 2321 1950 2361 1984
rect 2395 1950 2435 1984
rect 2469 1950 2509 1984
rect 2543 1950 2583 1984
rect 2617 1950 2657 1984
rect 2691 1950 2731 1984
rect 2765 1950 2805 1984
rect 2839 1950 2879 1984
rect 2913 1950 2953 1984
rect 2987 1950 3027 1984
rect 3061 1950 3101 1984
rect 3135 1950 3175 1984
rect 3209 1950 3249 1984
rect 3283 1950 3323 1984
rect 3357 1950 3397 1984
rect 3431 1950 3471 1984
rect 3505 1950 3545 1984
rect 3579 1950 3679 1984
rect 579 1912 3679 1950
rect 579 1878 679 1912
rect 713 1878 752 1912
rect 786 1878 825 1912
rect 859 1878 898 1912
rect 932 1878 971 1912
rect 1005 1878 1044 1912
rect 1078 1878 1117 1912
rect 1151 1878 1190 1912
rect 1224 1878 1263 1912
rect 1297 1878 1336 1912
rect 1370 1878 1409 1912
rect 1443 1878 1482 1912
rect 1516 1878 1555 1912
rect 1589 1878 1628 1912
rect 1662 1878 1701 1912
rect 1735 1878 1774 1912
rect 1808 1878 1847 1912
rect 1881 1878 1920 1912
rect 1954 1878 1993 1912
rect 2027 1878 2066 1912
rect 2100 1878 2139 1912
rect 2173 1878 2213 1912
rect 2247 1878 2287 1912
rect 2321 1878 2361 1912
rect 2395 1878 2435 1912
rect 2469 1878 2509 1912
rect 2543 1878 2583 1912
rect 2617 1878 2657 1912
rect 2691 1878 2731 1912
rect 2765 1878 2805 1912
rect 2839 1878 2879 1912
rect 2913 1878 2953 1912
rect 2987 1878 3027 1912
rect 3061 1878 3101 1912
rect 3135 1878 3175 1912
rect 3209 1878 3249 1912
rect 3283 1878 3323 1912
rect 3357 1878 3397 1912
rect 3431 1878 3471 1912
rect 3505 1878 3545 1912
rect 3579 1878 3679 1912
rect 3821 1950 3921 1984
rect 3955 1950 3995 1984
rect 4029 1950 4069 1984
rect 4103 1950 4143 1984
rect 4177 1950 4217 1984
rect 4251 1950 4291 1984
rect 4325 1950 4365 1984
rect 4399 1950 4439 1984
rect 4473 1950 4513 1984
rect 4547 1950 4587 1984
rect 4621 1950 4661 1984
rect 4695 1950 4735 1984
rect 4769 1950 4809 1984
rect 4843 1950 4883 1984
rect 4917 1950 4957 1984
rect 4991 1950 5031 1984
rect 5065 1950 5105 1984
rect 5139 1950 5179 1984
rect 5213 1950 5253 1984
rect 5287 1950 5327 1984
rect 5361 1950 5400 1984
rect 5434 1950 5473 1984
rect 5507 1950 5546 1984
rect 5580 1950 5619 1984
rect 5653 1950 5692 1984
rect 5726 1950 5765 1984
rect 5799 1950 5838 1984
rect 5872 1950 5911 1984
rect 5945 1950 5984 1984
rect 6018 1950 6057 1984
rect 6091 1950 6130 1984
rect 6164 1950 6203 1984
rect 6237 1950 6276 1984
rect 6310 1950 6349 1984
rect 6383 1950 6422 1984
rect 6456 1950 6495 1984
rect 6529 1950 6568 1984
rect 6602 1950 6641 1984
rect 6675 1950 6714 1984
rect 6748 1950 6787 1984
rect 6821 1950 6921 1984
rect 3821 1912 6921 1950
rect 3821 1878 3921 1912
rect 3955 1878 3995 1912
rect 4029 1878 4069 1912
rect 4103 1878 4143 1912
rect 4177 1878 4217 1912
rect 4251 1878 4291 1912
rect 4325 1878 4365 1912
rect 4399 1878 4439 1912
rect 4473 1878 4513 1912
rect 4547 1878 4587 1912
rect 4621 1878 4661 1912
rect 4695 1878 4735 1912
rect 4769 1878 4809 1912
rect 4843 1878 4883 1912
rect 4917 1878 4957 1912
rect 4991 1878 5031 1912
rect 5065 1878 5105 1912
rect 5139 1878 5179 1912
rect 5213 1878 5253 1912
rect 5287 1878 5327 1912
rect 5361 1878 5400 1912
rect 5434 1878 5473 1912
rect 5507 1878 5546 1912
rect 5580 1878 5619 1912
rect 5653 1878 5692 1912
rect 5726 1878 5765 1912
rect 5799 1878 5838 1912
rect 5872 1878 5911 1912
rect 5945 1878 5984 1912
rect 6018 1878 6057 1912
rect 6091 1878 6130 1912
rect 6164 1878 6203 1912
rect 6237 1878 6276 1912
rect 6310 1878 6349 1912
rect 6383 1878 6422 1912
rect 6456 1878 6495 1912
rect 6529 1878 6568 1912
rect 6602 1878 6641 1912
rect 6675 1878 6714 1912
rect 6748 1878 6787 1912
rect 6821 1878 6921 1912
rect 7063 1950 7163 1984
rect 7197 1950 7236 1984
rect 7270 1950 7309 1984
rect 7343 1950 7382 1984
rect 7416 1950 7455 1984
rect 7489 1950 7528 1984
rect 7562 1950 7601 1984
rect 7635 1950 7674 1984
rect 7708 1950 7747 1984
rect 7781 1950 7820 1984
rect 7854 1950 7893 1984
rect 7927 1950 7966 1984
rect 8000 1950 8039 1984
rect 8073 1950 8112 1984
rect 8146 1950 8185 1984
rect 8219 1950 8258 1984
rect 8292 1950 8331 1984
rect 8365 1950 8404 1984
rect 8438 1950 8477 1984
rect 8511 1950 8550 1984
rect 8584 1950 8623 1984
rect 8657 1950 8697 1984
rect 8731 1950 8771 1984
rect 8805 1950 8845 1984
rect 8879 1950 8919 1984
rect 8953 1950 8993 1984
rect 9027 1950 9067 1984
rect 9101 1950 9141 1984
rect 9175 1950 9215 1984
rect 9249 1950 9289 1984
rect 9323 1950 9363 1984
rect 9397 1950 9437 1984
rect 9471 1950 9511 1984
rect 9545 1950 9585 1984
rect 9619 1950 9659 1984
rect 9693 1950 9733 1984
rect 9767 1950 9807 1984
rect 9841 1950 9881 1984
rect 9915 1950 9955 1984
rect 9989 1950 10029 1984
rect 10063 1950 10163 1984
rect 7063 1912 10163 1950
rect 7063 1878 7163 1912
rect 7197 1878 7236 1912
rect 7270 1878 7309 1912
rect 7343 1878 7382 1912
rect 7416 1878 7455 1912
rect 7489 1878 7528 1912
rect 7562 1878 7601 1912
rect 7635 1878 7674 1912
rect 7708 1878 7747 1912
rect 7781 1878 7820 1912
rect 7854 1878 7893 1912
rect 7927 1878 7966 1912
rect 8000 1878 8039 1912
rect 8073 1878 8112 1912
rect 8146 1878 8185 1912
rect 8219 1878 8258 1912
rect 8292 1878 8331 1912
rect 8365 1878 8404 1912
rect 8438 1878 8477 1912
rect 8511 1878 8550 1912
rect 8584 1878 8623 1912
rect 8657 1878 8697 1912
rect 8731 1878 8771 1912
rect 8805 1878 8845 1912
rect 8879 1878 8919 1912
rect 8953 1878 8993 1912
rect 9027 1878 9067 1912
rect 9101 1878 9141 1912
rect 9175 1878 9215 1912
rect 9249 1878 9289 1912
rect 9323 1878 9363 1912
rect 9397 1878 9437 1912
rect 9471 1878 9511 1912
rect 9545 1878 9585 1912
rect 9619 1878 9659 1912
rect 9693 1878 9733 1912
rect 9767 1878 9807 1912
rect 9841 1878 9881 1912
rect 9915 1878 9955 1912
rect 9989 1878 10029 1912
rect 10063 1878 10163 1912
rect 10305 1950 10405 1984
rect 10439 1950 10479 1984
rect 10513 1950 10553 1984
rect 10587 1950 10627 1984
rect 10661 1950 10701 1984
rect 10735 1950 10775 1984
rect 10809 1950 10849 1984
rect 10883 1950 10923 1984
rect 10957 1950 10997 1984
rect 11031 1950 11071 1984
rect 11105 1950 11145 1984
rect 11179 1950 11219 1984
rect 11253 1950 11293 1984
rect 11327 1950 11367 1984
rect 11401 1950 11441 1984
rect 11475 1950 11515 1984
rect 11549 1950 11589 1984
rect 11623 1950 11663 1984
rect 11697 1950 11737 1984
rect 11771 1950 11811 1984
rect 11845 1950 11884 1984
rect 11918 1950 11957 1984
rect 11991 1950 12030 1984
rect 12064 1950 12103 1984
rect 12137 1950 12176 1984
rect 12210 1950 12249 1984
rect 12283 1950 12322 1984
rect 12356 1950 12395 1984
rect 12429 1950 12468 1984
rect 12502 1950 12541 1984
rect 12575 1950 12614 1984
rect 12648 1950 12687 1984
rect 12721 1950 12760 1984
rect 12794 1950 12833 1984
rect 12867 1950 12906 1984
rect 12940 1950 12979 1984
rect 13013 1950 13052 1984
rect 13086 1950 13125 1984
rect 13159 1950 13198 1984
rect 13232 1950 13271 1984
rect 13305 1950 13405 1984
rect 10305 1912 13405 1950
rect 10305 1878 10405 1912
rect 10439 1878 10479 1912
rect 10513 1878 10553 1912
rect 10587 1878 10627 1912
rect 10661 1878 10701 1912
rect 10735 1878 10775 1912
rect 10809 1878 10849 1912
rect 10883 1878 10923 1912
rect 10957 1878 10997 1912
rect 11031 1878 11071 1912
rect 11105 1878 11145 1912
rect 11179 1878 11219 1912
rect 11253 1878 11293 1912
rect 11327 1878 11367 1912
rect 11401 1878 11441 1912
rect 11475 1878 11515 1912
rect 11549 1878 11589 1912
rect 11623 1878 11663 1912
rect 11697 1878 11737 1912
rect 11771 1878 11811 1912
rect 11845 1878 11884 1912
rect 11918 1878 11957 1912
rect 11991 1878 12030 1912
rect 12064 1878 12103 1912
rect 12137 1878 12176 1912
rect 12210 1878 12249 1912
rect 12283 1878 12322 1912
rect 12356 1878 12395 1912
rect 12429 1878 12468 1912
rect 12502 1878 12541 1912
rect 12575 1878 12614 1912
rect 12648 1878 12687 1912
rect 12721 1878 12760 1912
rect 12794 1878 12833 1912
rect 12867 1878 12906 1912
rect 12940 1878 12979 1912
rect 13013 1878 13052 1912
rect 13086 1878 13125 1912
rect 13159 1878 13198 1912
rect 13232 1878 13271 1912
rect 13305 1878 13405 1912
rect 13547 1950 13647 1984
rect 13681 1950 13720 1984
rect 13754 1950 13793 1984
rect 13827 1950 13866 1984
rect 13900 1950 13939 1984
rect 13973 1950 14012 1984
rect 14046 1950 14085 1984
rect 14119 1950 14158 1984
rect 14192 1950 14231 1984
rect 14265 1950 14304 1984
rect 14338 1950 14377 1984
rect 14411 1950 14450 1984
rect 14484 1950 14523 1984
rect 14557 1950 14596 1984
rect 14630 1950 14669 1984
rect 14703 1950 14742 1984
rect 14776 1950 14815 1984
rect 14849 1950 14888 1984
rect 14922 1950 14961 1984
rect 14995 1950 15034 1984
rect 15068 1950 15107 1984
rect 15141 1950 15181 1984
rect 15215 1950 15255 1984
rect 15289 1950 15329 1984
rect 15363 1950 15403 1984
rect 15437 1950 15477 1984
rect 15511 1950 15551 1984
rect 15585 1950 15625 1984
rect 15659 1950 15699 1984
rect 15733 1950 15773 1984
rect 15807 1950 15847 1984
rect 15881 1950 15921 1984
rect 15955 1950 15995 1984
rect 16029 1950 16069 1984
rect 16103 1950 16143 1984
rect 16177 1950 16217 1984
rect 16251 1950 16291 1984
rect 16325 1950 16365 1984
rect 16399 1950 16439 1984
rect 16473 1950 16513 1984
rect 16547 1950 16647 1984
rect 13547 1912 16647 1950
rect 13547 1878 13647 1912
rect 13681 1878 13720 1912
rect 13754 1878 13793 1912
rect 13827 1878 13866 1912
rect 13900 1878 13939 1912
rect 13973 1878 14012 1912
rect 14046 1878 14085 1912
rect 14119 1878 14158 1912
rect 14192 1878 14231 1912
rect 14265 1878 14304 1912
rect 14338 1878 14377 1912
rect 14411 1878 14450 1912
rect 14484 1878 14523 1912
rect 14557 1878 14596 1912
rect 14630 1878 14669 1912
rect 14703 1878 14742 1912
rect 14776 1878 14815 1912
rect 14849 1878 14888 1912
rect 14922 1878 14961 1912
rect 14995 1878 15034 1912
rect 15068 1878 15107 1912
rect 15141 1878 15181 1912
rect 15215 1878 15255 1912
rect 15289 1878 15329 1912
rect 15363 1878 15403 1912
rect 15437 1878 15477 1912
rect 15511 1878 15551 1912
rect 15585 1878 15625 1912
rect 15659 1878 15699 1912
rect 15733 1878 15773 1912
rect 15807 1878 15847 1912
rect 15881 1878 15921 1912
rect 15955 1878 15995 1912
rect 16029 1878 16069 1912
rect 16103 1878 16143 1912
rect 16177 1878 16217 1912
rect 16251 1878 16291 1912
rect 16325 1878 16365 1912
rect 16399 1878 16439 1912
rect 16473 1878 16513 1912
rect 16547 1878 16647 1912
rect 16789 1950 16889 1984
rect 16923 1950 16963 1984
rect 16997 1950 17037 1984
rect 17071 1950 17111 1984
rect 17145 1950 17185 1984
rect 17219 1950 17259 1984
rect 17293 1950 17333 1984
rect 17367 1950 17407 1984
rect 17441 1950 17481 1984
rect 17515 1950 17555 1984
rect 17589 1950 17629 1984
rect 17663 1950 17703 1984
rect 17737 1950 17777 1984
rect 17811 1950 17851 1984
rect 17885 1950 17925 1984
rect 17959 1950 17999 1984
rect 18033 1950 18073 1984
rect 18107 1950 18147 1984
rect 18181 1950 18221 1984
rect 18255 1950 18295 1984
rect 18329 1950 18368 1984
rect 18402 1950 18441 1984
rect 18475 1950 18514 1984
rect 18548 1950 18587 1984
rect 18621 1950 18660 1984
rect 18694 1950 18733 1984
rect 18767 1950 18806 1984
rect 18840 1950 18879 1984
rect 18913 1950 18952 1984
rect 18986 1950 19025 1984
rect 19059 1950 19098 1984
rect 19132 1950 19171 1984
rect 19205 1950 19244 1984
rect 19278 1950 19317 1984
rect 19351 1950 19390 1984
rect 19424 1950 19463 1984
rect 19497 1950 19536 1984
rect 19570 1950 19609 1984
rect 19643 1950 19682 1984
rect 19716 1950 19755 1984
rect 19789 1950 19889 1984
rect 16789 1912 19889 1950
rect 16789 1878 16889 1912
rect 16923 1878 16963 1912
rect 16997 1878 17037 1912
rect 17071 1878 17111 1912
rect 17145 1878 17185 1912
rect 17219 1878 17259 1912
rect 17293 1878 17333 1912
rect 17367 1878 17407 1912
rect 17441 1878 17481 1912
rect 17515 1878 17555 1912
rect 17589 1878 17629 1912
rect 17663 1878 17703 1912
rect 17737 1878 17777 1912
rect 17811 1878 17851 1912
rect 17885 1878 17925 1912
rect 17959 1878 17999 1912
rect 18033 1878 18073 1912
rect 18107 1878 18147 1912
rect 18181 1878 18221 1912
rect 18255 1878 18295 1912
rect 18329 1878 18368 1912
rect 18402 1878 18441 1912
rect 18475 1878 18514 1912
rect 18548 1878 18587 1912
rect 18621 1878 18660 1912
rect 18694 1878 18733 1912
rect 18767 1878 18806 1912
rect 18840 1878 18879 1912
rect 18913 1878 18952 1912
rect 18986 1878 19025 1912
rect 19059 1878 19098 1912
rect 19132 1878 19171 1912
rect 19205 1878 19244 1912
rect 19278 1878 19317 1912
rect 19351 1878 19390 1912
rect 19424 1878 19463 1912
rect 19497 1878 19536 1912
rect 19570 1878 19609 1912
rect 19643 1878 19682 1912
rect 19716 1878 19755 1912
rect 19789 1878 19889 1912
<< viali >>
rect 679 2774 713 2808
rect 752 2774 786 2808
rect 825 2774 859 2808
rect 898 2774 932 2808
rect 971 2774 1005 2808
rect 1044 2774 1078 2808
rect 1117 2774 1151 2808
rect 1190 2774 1224 2808
rect 1263 2774 1297 2808
rect 1336 2774 1370 2808
rect 1409 2774 1443 2808
rect 1482 2774 1516 2808
rect 1555 2774 1589 2808
rect 1628 2774 1662 2808
rect 1701 2774 1735 2808
rect 1774 2774 1808 2808
rect 1847 2774 1881 2808
rect 1920 2774 1954 2808
rect 1993 2774 2027 2808
rect 2066 2774 2100 2808
rect 2139 2774 2173 2808
rect 2213 2774 2247 2808
rect 2287 2774 2321 2808
rect 2361 2774 2395 2808
rect 2435 2774 2469 2808
rect 2509 2774 2543 2808
rect 2583 2774 2617 2808
rect 2657 2774 2691 2808
rect 2731 2774 2765 2808
rect 2805 2774 2839 2808
rect 2879 2774 2913 2808
rect 2953 2774 2987 2808
rect 3027 2774 3061 2808
rect 3101 2774 3135 2808
rect 3175 2774 3209 2808
rect 3249 2774 3283 2808
rect 3323 2774 3357 2808
rect 3397 2774 3431 2808
rect 3471 2774 3505 2808
rect 3545 2774 3579 2808
rect 679 2702 713 2736
rect 752 2702 786 2736
rect 825 2702 859 2736
rect 898 2702 932 2736
rect 971 2702 1005 2736
rect 1044 2702 1078 2736
rect 1117 2702 1151 2736
rect 1190 2702 1224 2736
rect 1263 2702 1297 2736
rect 1336 2702 1370 2736
rect 1409 2702 1443 2736
rect 1482 2702 1516 2736
rect 1555 2702 1589 2736
rect 1628 2702 1662 2736
rect 1701 2702 1735 2736
rect 1774 2702 1808 2736
rect 1847 2702 1881 2736
rect 1920 2702 1954 2736
rect 1993 2702 2027 2736
rect 2066 2702 2100 2736
rect 2139 2702 2173 2736
rect 2213 2702 2247 2736
rect 2287 2702 2321 2736
rect 2361 2702 2395 2736
rect 2435 2702 2469 2736
rect 2509 2702 2543 2736
rect 2583 2702 2617 2736
rect 2657 2702 2691 2736
rect 2731 2702 2765 2736
rect 2805 2702 2839 2736
rect 2879 2702 2913 2736
rect 2953 2702 2987 2736
rect 3027 2702 3061 2736
rect 3101 2702 3135 2736
rect 3175 2702 3209 2736
rect 3249 2702 3283 2736
rect 3323 2702 3357 2736
rect 3397 2702 3431 2736
rect 3471 2702 3505 2736
rect 3545 2702 3579 2736
rect 3921 2774 3955 2808
rect 3995 2774 4029 2808
rect 4069 2774 4103 2808
rect 4143 2774 4177 2808
rect 4217 2774 4251 2808
rect 4291 2774 4325 2808
rect 4365 2774 4399 2808
rect 4439 2774 4473 2808
rect 4513 2774 4547 2808
rect 4587 2774 4621 2808
rect 4661 2774 4695 2808
rect 4735 2774 4769 2808
rect 4809 2774 4843 2808
rect 4883 2774 4917 2808
rect 4957 2774 4991 2808
rect 5031 2774 5065 2808
rect 5105 2774 5139 2808
rect 5179 2774 5213 2808
rect 5253 2774 5287 2808
rect 5327 2774 5361 2808
rect 5400 2774 5434 2808
rect 5473 2774 5507 2808
rect 5546 2774 5580 2808
rect 5619 2774 5653 2808
rect 5692 2774 5726 2808
rect 5765 2774 5799 2808
rect 5838 2774 5872 2808
rect 5911 2774 5945 2808
rect 5984 2774 6018 2808
rect 6057 2774 6091 2808
rect 6130 2774 6164 2808
rect 6203 2774 6237 2808
rect 6276 2774 6310 2808
rect 6349 2774 6383 2808
rect 6422 2774 6456 2808
rect 6495 2774 6529 2808
rect 6568 2774 6602 2808
rect 6641 2774 6675 2808
rect 6714 2774 6748 2808
rect 6787 2774 6821 2808
rect 3921 2702 3955 2736
rect 3995 2702 4029 2736
rect 4069 2702 4103 2736
rect 4143 2702 4177 2736
rect 4217 2702 4251 2736
rect 4291 2702 4325 2736
rect 4365 2702 4399 2736
rect 4439 2702 4473 2736
rect 4513 2702 4547 2736
rect 4587 2702 4621 2736
rect 4661 2702 4695 2736
rect 4735 2702 4769 2736
rect 4809 2702 4843 2736
rect 4883 2702 4917 2736
rect 4957 2702 4991 2736
rect 5031 2702 5065 2736
rect 5105 2702 5139 2736
rect 5179 2702 5213 2736
rect 5253 2702 5287 2736
rect 5327 2702 5361 2736
rect 5400 2702 5434 2736
rect 5473 2702 5507 2736
rect 5546 2702 5580 2736
rect 5619 2702 5653 2736
rect 5692 2702 5726 2736
rect 5765 2702 5799 2736
rect 5838 2702 5872 2736
rect 5911 2702 5945 2736
rect 5984 2702 6018 2736
rect 6057 2702 6091 2736
rect 6130 2702 6164 2736
rect 6203 2702 6237 2736
rect 6276 2702 6310 2736
rect 6349 2702 6383 2736
rect 6422 2702 6456 2736
rect 6495 2702 6529 2736
rect 6568 2702 6602 2736
rect 6641 2702 6675 2736
rect 6714 2702 6748 2736
rect 6787 2702 6821 2736
rect 7163 2774 7197 2808
rect 7236 2774 7270 2808
rect 7309 2774 7343 2808
rect 7382 2774 7416 2808
rect 7455 2774 7489 2808
rect 7528 2774 7562 2808
rect 7601 2774 7635 2808
rect 7674 2774 7708 2808
rect 7747 2774 7781 2808
rect 7820 2774 7854 2808
rect 7893 2774 7927 2808
rect 7966 2774 8000 2808
rect 8039 2774 8073 2808
rect 8112 2774 8146 2808
rect 8185 2774 8219 2808
rect 8258 2774 8292 2808
rect 8331 2774 8365 2808
rect 8404 2774 8438 2808
rect 8477 2774 8511 2808
rect 8550 2774 8584 2808
rect 8623 2774 8657 2808
rect 8697 2774 8731 2808
rect 8771 2774 8805 2808
rect 8845 2774 8879 2808
rect 8919 2774 8953 2808
rect 8993 2774 9027 2808
rect 9067 2774 9101 2808
rect 9141 2774 9175 2808
rect 9215 2774 9249 2808
rect 9289 2774 9323 2808
rect 9363 2774 9397 2808
rect 9437 2774 9471 2808
rect 9511 2774 9545 2808
rect 9585 2774 9619 2808
rect 9659 2774 9693 2808
rect 9733 2774 9767 2808
rect 9807 2774 9841 2808
rect 9881 2774 9915 2808
rect 9955 2774 9989 2808
rect 10029 2774 10063 2808
rect 7163 2702 7197 2736
rect 7236 2702 7270 2736
rect 7309 2702 7343 2736
rect 7382 2702 7416 2736
rect 7455 2702 7489 2736
rect 7528 2702 7562 2736
rect 7601 2702 7635 2736
rect 7674 2702 7708 2736
rect 7747 2702 7781 2736
rect 7820 2702 7854 2736
rect 7893 2702 7927 2736
rect 7966 2702 8000 2736
rect 8039 2702 8073 2736
rect 8112 2702 8146 2736
rect 8185 2702 8219 2736
rect 8258 2702 8292 2736
rect 8331 2702 8365 2736
rect 8404 2702 8438 2736
rect 8477 2702 8511 2736
rect 8550 2702 8584 2736
rect 8623 2702 8657 2736
rect 8697 2702 8731 2736
rect 8771 2702 8805 2736
rect 8845 2702 8879 2736
rect 8919 2702 8953 2736
rect 8993 2702 9027 2736
rect 9067 2702 9101 2736
rect 9141 2702 9175 2736
rect 9215 2702 9249 2736
rect 9289 2702 9323 2736
rect 9363 2702 9397 2736
rect 9437 2702 9471 2736
rect 9511 2702 9545 2736
rect 9585 2702 9619 2736
rect 9659 2702 9693 2736
rect 9733 2702 9767 2736
rect 9807 2702 9841 2736
rect 9881 2702 9915 2736
rect 9955 2702 9989 2736
rect 10029 2702 10063 2736
rect 10405 2774 10439 2808
rect 10479 2774 10513 2808
rect 10553 2774 10587 2808
rect 10627 2774 10661 2808
rect 10701 2774 10735 2808
rect 10775 2774 10809 2808
rect 10849 2774 10883 2808
rect 10923 2774 10957 2808
rect 10997 2774 11031 2808
rect 11071 2774 11105 2808
rect 11145 2774 11179 2808
rect 11219 2774 11253 2808
rect 11293 2774 11327 2808
rect 11367 2774 11401 2808
rect 11441 2774 11475 2808
rect 11515 2774 11549 2808
rect 11589 2774 11623 2808
rect 11663 2774 11697 2808
rect 11737 2774 11771 2808
rect 11811 2774 11845 2808
rect 11884 2774 11918 2808
rect 11957 2774 11991 2808
rect 12030 2774 12064 2808
rect 12103 2774 12137 2808
rect 12176 2774 12210 2808
rect 12249 2774 12283 2808
rect 12322 2774 12356 2808
rect 12395 2774 12429 2808
rect 12468 2774 12502 2808
rect 12541 2774 12575 2808
rect 12614 2774 12648 2808
rect 12687 2774 12721 2808
rect 12760 2774 12794 2808
rect 12833 2774 12867 2808
rect 12906 2774 12940 2808
rect 12979 2774 13013 2808
rect 13052 2774 13086 2808
rect 13125 2774 13159 2808
rect 13198 2774 13232 2808
rect 13271 2774 13305 2808
rect 10405 2702 10439 2736
rect 10479 2702 10513 2736
rect 10553 2702 10587 2736
rect 10627 2702 10661 2736
rect 10701 2702 10735 2736
rect 10775 2702 10809 2736
rect 10849 2702 10883 2736
rect 10923 2702 10957 2736
rect 10997 2702 11031 2736
rect 11071 2702 11105 2736
rect 11145 2702 11179 2736
rect 11219 2702 11253 2736
rect 11293 2702 11327 2736
rect 11367 2702 11401 2736
rect 11441 2702 11475 2736
rect 11515 2702 11549 2736
rect 11589 2702 11623 2736
rect 11663 2702 11697 2736
rect 11737 2702 11771 2736
rect 11811 2702 11845 2736
rect 11884 2702 11918 2736
rect 11957 2702 11991 2736
rect 12030 2702 12064 2736
rect 12103 2702 12137 2736
rect 12176 2702 12210 2736
rect 12249 2702 12283 2736
rect 12322 2702 12356 2736
rect 12395 2702 12429 2736
rect 12468 2702 12502 2736
rect 12541 2702 12575 2736
rect 12614 2702 12648 2736
rect 12687 2702 12721 2736
rect 12760 2702 12794 2736
rect 12833 2702 12867 2736
rect 12906 2702 12940 2736
rect 12979 2702 13013 2736
rect 13052 2702 13086 2736
rect 13125 2702 13159 2736
rect 13198 2702 13232 2736
rect 13271 2702 13305 2736
rect 13647 2774 13681 2808
rect 13720 2774 13754 2808
rect 13793 2774 13827 2808
rect 13866 2774 13900 2808
rect 13939 2774 13973 2808
rect 14012 2774 14046 2808
rect 14085 2774 14119 2808
rect 14158 2774 14192 2808
rect 14231 2774 14265 2808
rect 14304 2774 14338 2808
rect 14377 2774 14411 2808
rect 14450 2774 14484 2808
rect 14523 2774 14557 2808
rect 14596 2774 14630 2808
rect 14669 2774 14703 2808
rect 14742 2774 14776 2808
rect 14815 2774 14849 2808
rect 14888 2774 14922 2808
rect 14961 2774 14995 2808
rect 15034 2774 15068 2808
rect 15107 2774 15141 2808
rect 15181 2774 15215 2808
rect 15255 2774 15289 2808
rect 15329 2774 15363 2808
rect 15403 2774 15437 2808
rect 15477 2774 15511 2808
rect 15551 2774 15585 2808
rect 15625 2774 15659 2808
rect 15699 2774 15733 2808
rect 15773 2774 15807 2808
rect 15847 2774 15881 2808
rect 15921 2774 15955 2808
rect 15995 2774 16029 2808
rect 16069 2774 16103 2808
rect 16143 2774 16177 2808
rect 16217 2774 16251 2808
rect 16291 2774 16325 2808
rect 16365 2774 16399 2808
rect 16439 2774 16473 2808
rect 16513 2774 16547 2808
rect 13647 2702 13681 2736
rect 13720 2702 13754 2736
rect 13793 2702 13827 2736
rect 13866 2702 13900 2736
rect 13939 2702 13973 2736
rect 14012 2702 14046 2736
rect 14085 2702 14119 2736
rect 14158 2702 14192 2736
rect 14231 2702 14265 2736
rect 14304 2702 14338 2736
rect 14377 2702 14411 2736
rect 14450 2702 14484 2736
rect 14523 2702 14557 2736
rect 14596 2702 14630 2736
rect 14669 2702 14703 2736
rect 14742 2702 14776 2736
rect 14815 2702 14849 2736
rect 14888 2702 14922 2736
rect 14961 2702 14995 2736
rect 15034 2702 15068 2736
rect 15107 2702 15141 2736
rect 15181 2702 15215 2736
rect 15255 2702 15289 2736
rect 15329 2702 15363 2736
rect 15403 2702 15437 2736
rect 15477 2702 15511 2736
rect 15551 2702 15585 2736
rect 15625 2702 15659 2736
rect 15699 2702 15733 2736
rect 15773 2702 15807 2736
rect 15847 2702 15881 2736
rect 15921 2702 15955 2736
rect 15995 2702 16029 2736
rect 16069 2702 16103 2736
rect 16143 2702 16177 2736
rect 16217 2702 16251 2736
rect 16291 2702 16325 2736
rect 16365 2702 16399 2736
rect 16439 2702 16473 2736
rect 16513 2702 16547 2736
rect 16889 2774 16923 2808
rect 16963 2774 16997 2808
rect 17037 2774 17071 2808
rect 17111 2774 17145 2808
rect 17185 2774 17219 2808
rect 17259 2774 17293 2808
rect 17333 2774 17367 2808
rect 17407 2774 17441 2808
rect 17481 2774 17515 2808
rect 17555 2774 17589 2808
rect 17629 2774 17663 2808
rect 17703 2774 17737 2808
rect 17777 2774 17811 2808
rect 17851 2774 17885 2808
rect 17925 2774 17959 2808
rect 17999 2774 18033 2808
rect 18073 2774 18107 2808
rect 18147 2774 18181 2808
rect 18221 2774 18255 2808
rect 18295 2774 18329 2808
rect 18368 2774 18402 2808
rect 18441 2774 18475 2808
rect 18514 2774 18548 2808
rect 18587 2774 18621 2808
rect 18660 2774 18694 2808
rect 18733 2774 18767 2808
rect 18806 2774 18840 2808
rect 18879 2774 18913 2808
rect 18952 2774 18986 2808
rect 19025 2774 19059 2808
rect 19098 2774 19132 2808
rect 19171 2774 19205 2808
rect 19244 2774 19278 2808
rect 19317 2774 19351 2808
rect 19390 2774 19424 2808
rect 19463 2774 19497 2808
rect 19536 2774 19570 2808
rect 19609 2774 19643 2808
rect 19682 2774 19716 2808
rect 19755 2774 19789 2808
rect 16889 2702 16923 2736
rect 16963 2702 16997 2736
rect 17037 2702 17071 2736
rect 17111 2702 17145 2736
rect 17185 2702 17219 2736
rect 17259 2702 17293 2736
rect 17333 2702 17367 2736
rect 17407 2702 17441 2736
rect 17481 2702 17515 2736
rect 17555 2702 17589 2736
rect 17629 2702 17663 2736
rect 17703 2702 17737 2736
rect 17777 2702 17811 2736
rect 17851 2702 17885 2736
rect 17925 2702 17959 2736
rect 17999 2702 18033 2736
rect 18073 2702 18107 2736
rect 18147 2702 18181 2736
rect 18221 2702 18255 2736
rect 18295 2702 18329 2736
rect 18368 2702 18402 2736
rect 18441 2702 18475 2736
rect 18514 2702 18548 2736
rect 18587 2702 18621 2736
rect 18660 2702 18694 2736
rect 18733 2702 18767 2736
rect 18806 2702 18840 2736
rect 18879 2702 18913 2736
rect 18952 2702 18986 2736
rect 19025 2702 19059 2736
rect 19098 2702 19132 2736
rect 19171 2702 19205 2736
rect 19244 2702 19278 2736
rect 19317 2702 19351 2736
rect 19390 2702 19424 2736
rect 19463 2702 19497 2736
rect 19536 2702 19570 2736
rect 19609 2702 19643 2736
rect 19682 2702 19716 2736
rect 19755 2702 19789 2736
rect 483 2598 517 2614
rect 483 2580 497 2598
rect 497 2580 517 2598
rect 555 2580 589 2614
rect 3701 2580 3735 2614
rect 3773 2580 3807 2614
rect 6943 2580 6977 2614
rect 7015 2580 7049 2614
rect 10185 2580 10219 2614
rect 10257 2580 10291 2614
rect 13451 2598 13485 2614
rect 13451 2580 13465 2598
rect 13465 2580 13485 2598
rect 13523 2580 13557 2614
rect 19937 2600 19971 2603
rect 19937 2569 19971 2600
rect 19937 2498 19971 2531
rect 19937 2497 19971 2498
rect 679 2362 713 2396
rect 752 2362 786 2396
rect 825 2362 859 2396
rect 898 2362 932 2396
rect 971 2362 1005 2396
rect 1044 2362 1078 2396
rect 1117 2362 1151 2396
rect 1190 2362 1224 2396
rect 1263 2362 1297 2396
rect 1336 2362 1370 2396
rect 1409 2362 1443 2396
rect 1482 2362 1516 2396
rect 1555 2362 1589 2396
rect 1628 2362 1662 2396
rect 1701 2362 1735 2396
rect 1774 2362 1808 2396
rect 1847 2362 1881 2396
rect 1920 2362 1954 2396
rect 1993 2362 2027 2396
rect 2066 2362 2100 2396
rect 2139 2362 2173 2396
rect 2213 2362 2247 2396
rect 2287 2362 2321 2396
rect 2361 2362 2395 2396
rect 2435 2362 2469 2396
rect 2509 2362 2543 2396
rect 2583 2362 2617 2396
rect 2657 2362 2691 2396
rect 2731 2362 2765 2396
rect 2805 2362 2839 2396
rect 2879 2362 2913 2396
rect 2953 2362 2987 2396
rect 3027 2362 3061 2396
rect 3101 2362 3135 2396
rect 3175 2362 3209 2396
rect 3249 2362 3283 2396
rect 3323 2362 3357 2396
rect 3397 2362 3431 2396
rect 3471 2362 3505 2396
rect 3545 2362 3579 2396
rect 679 2290 713 2324
rect 752 2290 786 2324
rect 825 2290 859 2324
rect 898 2290 932 2324
rect 971 2290 1005 2324
rect 1044 2290 1078 2324
rect 1117 2290 1151 2324
rect 1190 2290 1224 2324
rect 1263 2290 1297 2324
rect 1336 2290 1370 2324
rect 1409 2290 1443 2324
rect 1482 2290 1516 2324
rect 1555 2290 1589 2324
rect 1628 2290 1662 2324
rect 1701 2290 1735 2324
rect 1774 2290 1808 2324
rect 1847 2290 1881 2324
rect 1920 2290 1954 2324
rect 1993 2290 2027 2324
rect 2066 2290 2100 2324
rect 2139 2290 2173 2324
rect 2213 2290 2247 2324
rect 2287 2290 2321 2324
rect 2361 2290 2395 2324
rect 2435 2290 2469 2324
rect 2509 2290 2543 2324
rect 2583 2290 2617 2324
rect 2657 2290 2691 2324
rect 2731 2290 2765 2324
rect 2805 2290 2839 2324
rect 2879 2290 2913 2324
rect 2953 2290 2987 2324
rect 3027 2290 3061 2324
rect 3101 2290 3135 2324
rect 3175 2290 3209 2324
rect 3249 2290 3283 2324
rect 3323 2290 3357 2324
rect 3397 2290 3431 2324
rect 3471 2290 3505 2324
rect 3545 2290 3579 2324
rect 3921 2362 3955 2396
rect 3995 2362 4029 2396
rect 4069 2362 4103 2396
rect 4143 2362 4177 2396
rect 4217 2362 4251 2396
rect 4291 2362 4325 2396
rect 4365 2362 4399 2396
rect 4439 2362 4473 2396
rect 4513 2362 4547 2396
rect 4587 2362 4621 2396
rect 4661 2362 4695 2396
rect 4735 2362 4769 2396
rect 4809 2362 4843 2396
rect 4883 2362 4917 2396
rect 4957 2362 4991 2396
rect 5031 2362 5065 2396
rect 5105 2362 5139 2396
rect 5179 2362 5213 2396
rect 5253 2362 5287 2396
rect 5327 2362 5361 2396
rect 5400 2362 5434 2396
rect 5473 2362 5507 2396
rect 5546 2362 5580 2396
rect 5619 2362 5653 2396
rect 5692 2362 5726 2396
rect 5765 2362 5799 2396
rect 5838 2362 5872 2396
rect 5911 2362 5945 2396
rect 5984 2362 6018 2396
rect 6057 2362 6091 2396
rect 6130 2362 6164 2396
rect 6203 2362 6237 2396
rect 6276 2362 6310 2396
rect 6349 2362 6383 2396
rect 6422 2362 6456 2396
rect 6495 2362 6529 2396
rect 6568 2362 6602 2396
rect 6641 2362 6675 2396
rect 6714 2362 6748 2396
rect 6787 2362 6821 2396
rect 3921 2290 3955 2324
rect 3995 2290 4029 2324
rect 4069 2290 4103 2324
rect 4143 2290 4177 2324
rect 4217 2290 4251 2324
rect 4291 2290 4325 2324
rect 4365 2290 4399 2324
rect 4439 2290 4473 2324
rect 4513 2290 4547 2324
rect 4587 2290 4621 2324
rect 4661 2290 4695 2324
rect 4735 2290 4769 2324
rect 4809 2290 4843 2324
rect 4883 2290 4917 2324
rect 4957 2290 4991 2324
rect 5031 2290 5065 2324
rect 5105 2290 5139 2324
rect 5179 2290 5213 2324
rect 5253 2290 5287 2324
rect 5327 2290 5361 2324
rect 5400 2290 5434 2324
rect 5473 2290 5507 2324
rect 5546 2290 5580 2324
rect 5619 2290 5653 2324
rect 5692 2290 5726 2324
rect 5765 2290 5799 2324
rect 5838 2290 5872 2324
rect 5911 2290 5945 2324
rect 5984 2290 6018 2324
rect 6057 2290 6091 2324
rect 6130 2290 6164 2324
rect 6203 2290 6237 2324
rect 6276 2290 6310 2324
rect 6349 2290 6383 2324
rect 6422 2290 6456 2324
rect 6495 2290 6529 2324
rect 6568 2290 6602 2324
rect 6641 2290 6675 2324
rect 6714 2290 6748 2324
rect 6787 2290 6821 2324
rect 7163 2362 7197 2396
rect 7236 2362 7270 2396
rect 7309 2362 7343 2396
rect 7382 2362 7416 2396
rect 7455 2362 7489 2396
rect 7528 2362 7562 2396
rect 7601 2362 7635 2396
rect 7674 2362 7708 2396
rect 7747 2362 7781 2396
rect 7820 2362 7854 2396
rect 7893 2362 7927 2396
rect 7966 2362 8000 2396
rect 8039 2362 8073 2396
rect 8112 2362 8146 2396
rect 8185 2362 8219 2396
rect 8258 2362 8292 2396
rect 8331 2362 8365 2396
rect 8404 2362 8438 2396
rect 8477 2362 8511 2396
rect 8550 2362 8584 2396
rect 8623 2362 8657 2396
rect 8697 2362 8731 2396
rect 8771 2362 8805 2396
rect 8845 2362 8879 2396
rect 8919 2362 8953 2396
rect 8993 2362 9027 2396
rect 9067 2362 9101 2396
rect 9141 2362 9175 2396
rect 9215 2362 9249 2396
rect 9289 2362 9323 2396
rect 9363 2362 9397 2396
rect 9437 2362 9471 2396
rect 9511 2362 9545 2396
rect 9585 2362 9619 2396
rect 9659 2362 9693 2396
rect 9733 2362 9767 2396
rect 9807 2362 9841 2396
rect 9881 2362 9915 2396
rect 9955 2362 9989 2396
rect 10029 2362 10063 2396
rect 7163 2290 7197 2324
rect 7236 2290 7270 2324
rect 7309 2290 7343 2324
rect 7382 2290 7416 2324
rect 7455 2290 7489 2324
rect 7528 2290 7562 2324
rect 7601 2290 7635 2324
rect 7674 2290 7708 2324
rect 7747 2290 7781 2324
rect 7820 2290 7854 2324
rect 7893 2290 7927 2324
rect 7966 2290 8000 2324
rect 8039 2290 8073 2324
rect 8112 2290 8146 2324
rect 8185 2290 8219 2324
rect 8258 2290 8292 2324
rect 8331 2290 8365 2324
rect 8404 2290 8438 2324
rect 8477 2290 8511 2324
rect 8550 2290 8584 2324
rect 8623 2290 8657 2324
rect 8697 2290 8731 2324
rect 8771 2290 8805 2324
rect 8845 2290 8879 2324
rect 8919 2290 8953 2324
rect 8993 2290 9027 2324
rect 9067 2290 9101 2324
rect 9141 2290 9175 2324
rect 9215 2290 9249 2324
rect 9289 2290 9323 2324
rect 9363 2290 9397 2324
rect 9437 2290 9471 2324
rect 9511 2290 9545 2324
rect 9585 2290 9619 2324
rect 9659 2290 9693 2324
rect 9733 2290 9767 2324
rect 9807 2290 9841 2324
rect 9881 2290 9915 2324
rect 9955 2290 9989 2324
rect 10029 2290 10063 2324
rect 10405 2362 10439 2396
rect 10479 2362 10513 2396
rect 10553 2362 10587 2396
rect 10627 2362 10661 2396
rect 10701 2362 10735 2396
rect 10775 2362 10809 2396
rect 10849 2362 10883 2396
rect 10923 2362 10957 2396
rect 10997 2362 11031 2396
rect 11071 2362 11105 2396
rect 11145 2362 11179 2396
rect 11219 2362 11253 2396
rect 11293 2362 11327 2396
rect 11367 2362 11401 2396
rect 11441 2362 11475 2396
rect 11515 2362 11549 2396
rect 11589 2362 11623 2396
rect 11663 2362 11697 2396
rect 11737 2362 11771 2396
rect 11811 2362 11845 2396
rect 11884 2362 11918 2396
rect 11957 2362 11991 2396
rect 12030 2362 12064 2396
rect 12103 2362 12137 2396
rect 12176 2362 12210 2396
rect 12249 2362 12283 2396
rect 12322 2362 12356 2396
rect 12395 2362 12429 2396
rect 12468 2362 12502 2396
rect 12541 2362 12575 2396
rect 12614 2362 12648 2396
rect 12687 2362 12721 2396
rect 12760 2362 12794 2396
rect 12833 2362 12867 2396
rect 12906 2362 12940 2396
rect 12979 2362 13013 2396
rect 13052 2362 13086 2396
rect 13125 2362 13159 2396
rect 13198 2362 13232 2396
rect 13271 2362 13305 2396
rect 10405 2290 10439 2324
rect 10479 2290 10513 2324
rect 10553 2290 10587 2324
rect 10627 2290 10661 2324
rect 10701 2290 10735 2324
rect 10775 2290 10809 2324
rect 10849 2290 10883 2324
rect 10923 2290 10957 2324
rect 10997 2290 11031 2324
rect 11071 2290 11105 2324
rect 11145 2290 11179 2324
rect 11219 2290 11253 2324
rect 11293 2290 11327 2324
rect 11367 2290 11401 2324
rect 11441 2290 11475 2324
rect 11515 2290 11549 2324
rect 11589 2290 11623 2324
rect 11663 2290 11697 2324
rect 11737 2290 11771 2324
rect 11811 2290 11845 2324
rect 11884 2290 11918 2324
rect 11957 2290 11991 2324
rect 12030 2290 12064 2324
rect 12103 2290 12137 2324
rect 12176 2290 12210 2324
rect 12249 2290 12283 2324
rect 12322 2290 12356 2324
rect 12395 2290 12429 2324
rect 12468 2290 12502 2324
rect 12541 2290 12575 2324
rect 12614 2290 12648 2324
rect 12687 2290 12721 2324
rect 12760 2290 12794 2324
rect 12833 2290 12867 2324
rect 12906 2290 12940 2324
rect 12979 2290 13013 2324
rect 13052 2290 13086 2324
rect 13125 2290 13159 2324
rect 13198 2290 13232 2324
rect 13271 2290 13305 2324
rect 13647 2362 13681 2396
rect 13720 2362 13754 2396
rect 13793 2362 13827 2396
rect 13866 2362 13900 2396
rect 13939 2362 13973 2396
rect 14012 2362 14046 2396
rect 14085 2362 14119 2396
rect 14158 2362 14192 2396
rect 14231 2362 14265 2396
rect 14304 2362 14338 2396
rect 14377 2362 14411 2396
rect 14450 2362 14484 2396
rect 14523 2362 14557 2396
rect 14596 2362 14630 2396
rect 14669 2362 14703 2396
rect 14742 2362 14776 2396
rect 14815 2362 14849 2396
rect 14888 2362 14922 2396
rect 14961 2362 14995 2396
rect 15034 2362 15068 2396
rect 15107 2362 15141 2396
rect 15181 2362 15215 2396
rect 15255 2362 15289 2396
rect 15329 2362 15363 2396
rect 15403 2362 15437 2396
rect 15477 2362 15511 2396
rect 15551 2362 15585 2396
rect 15625 2362 15659 2396
rect 15699 2362 15733 2396
rect 15773 2362 15807 2396
rect 15847 2362 15881 2396
rect 15921 2362 15955 2396
rect 15995 2362 16029 2396
rect 16069 2362 16103 2396
rect 16143 2362 16177 2396
rect 16217 2362 16251 2396
rect 16291 2362 16325 2396
rect 16365 2362 16399 2396
rect 16439 2362 16473 2396
rect 16513 2362 16547 2396
rect 13647 2290 13681 2324
rect 13720 2290 13754 2324
rect 13793 2290 13827 2324
rect 13866 2290 13900 2324
rect 13939 2290 13973 2324
rect 14012 2290 14046 2324
rect 14085 2290 14119 2324
rect 14158 2290 14192 2324
rect 14231 2290 14265 2324
rect 14304 2290 14338 2324
rect 14377 2290 14411 2324
rect 14450 2290 14484 2324
rect 14523 2290 14557 2324
rect 14596 2290 14630 2324
rect 14669 2290 14703 2324
rect 14742 2290 14776 2324
rect 14815 2290 14849 2324
rect 14888 2290 14922 2324
rect 14961 2290 14995 2324
rect 15034 2290 15068 2324
rect 15107 2290 15141 2324
rect 15181 2290 15215 2324
rect 15255 2290 15289 2324
rect 15329 2290 15363 2324
rect 15403 2290 15437 2324
rect 15477 2290 15511 2324
rect 15551 2290 15585 2324
rect 15625 2290 15659 2324
rect 15699 2290 15733 2324
rect 15773 2290 15807 2324
rect 15847 2290 15881 2324
rect 15921 2290 15955 2324
rect 15995 2290 16029 2324
rect 16069 2290 16103 2324
rect 16143 2290 16177 2324
rect 16217 2290 16251 2324
rect 16291 2290 16325 2324
rect 16365 2290 16399 2324
rect 16439 2290 16473 2324
rect 16513 2290 16547 2324
rect 16889 2362 16923 2396
rect 16963 2362 16997 2396
rect 17037 2362 17071 2396
rect 17111 2362 17145 2396
rect 17185 2362 17219 2396
rect 17259 2362 17293 2396
rect 17333 2362 17367 2396
rect 17407 2362 17441 2396
rect 17481 2362 17515 2396
rect 17555 2362 17589 2396
rect 17629 2362 17663 2396
rect 17703 2362 17737 2396
rect 17777 2362 17811 2396
rect 17851 2362 17885 2396
rect 17925 2362 17959 2396
rect 17999 2362 18033 2396
rect 18073 2362 18107 2396
rect 18147 2362 18181 2396
rect 18221 2362 18255 2396
rect 18295 2362 18329 2396
rect 18368 2362 18402 2396
rect 18441 2362 18475 2396
rect 18514 2362 18548 2396
rect 18587 2362 18621 2396
rect 18660 2362 18694 2396
rect 18733 2362 18767 2396
rect 18806 2362 18840 2396
rect 18879 2362 18913 2396
rect 18952 2362 18986 2396
rect 19025 2362 19059 2396
rect 19098 2362 19132 2396
rect 19171 2362 19205 2396
rect 19244 2362 19278 2396
rect 19317 2362 19351 2396
rect 19390 2362 19424 2396
rect 19463 2362 19497 2396
rect 19536 2362 19570 2396
rect 19609 2362 19643 2396
rect 19682 2362 19716 2396
rect 19755 2362 19789 2396
rect 16889 2290 16923 2324
rect 16963 2290 16997 2324
rect 17037 2290 17071 2324
rect 17111 2290 17145 2324
rect 17185 2290 17219 2324
rect 17259 2290 17293 2324
rect 17333 2290 17367 2324
rect 17407 2290 17441 2324
rect 17481 2290 17515 2324
rect 17555 2290 17589 2324
rect 17629 2290 17663 2324
rect 17703 2290 17737 2324
rect 17777 2290 17811 2324
rect 17851 2290 17885 2324
rect 17925 2290 17959 2324
rect 17999 2290 18033 2324
rect 18073 2290 18107 2324
rect 18147 2290 18181 2324
rect 18221 2290 18255 2324
rect 18295 2290 18329 2324
rect 18368 2290 18402 2324
rect 18441 2290 18475 2324
rect 18514 2290 18548 2324
rect 18587 2290 18621 2324
rect 18660 2290 18694 2324
rect 18733 2290 18767 2324
rect 18806 2290 18840 2324
rect 18879 2290 18913 2324
rect 18952 2290 18986 2324
rect 19025 2290 19059 2324
rect 19098 2290 19132 2324
rect 19171 2290 19205 2324
rect 19244 2290 19278 2324
rect 19317 2290 19351 2324
rect 19390 2290 19424 2324
rect 19463 2290 19497 2324
rect 19536 2290 19570 2324
rect 19609 2290 19643 2324
rect 19682 2290 19716 2324
rect 19755 2290 19789 2324
rect 483 2086 497 2106
rect 497 2086 517 2106
rect 483 2072 517 2086
rect 555 2072 589 2106
rect 3701 2072 3735 2106
rect 3773 2072 3807 2106
rect 6943 2072 6977 2106
rect 7015 2072 7049 2106
rect 10185 2072 10219 2106
rect 19937 2188 19971 2191
rect 19937 2157 19971 2188
rect 10257 2072 10291 2106
rect 13451 2086 13465 2106
rect 13465 2086 13485 2106
rect 13451 2072 13485 2086
rect 13523 2072 13557 2106
rect 19937 2086 19971 2119
rect 19937 2085 19971 2086
rect 679 1950 713 1984
rect 752 1950 786 1984
rect 825 1950 859 1984
rect 898 1950 932 1984
rect 971 1950 1005 1984
rect 1044 1950 1078 1984
rect 1117 1950 1151 1984
rect 1190 1950 1224 1984
rect 1263 1950 1297 1984
rect 1336 1950 1370 1984
rect 1409 1950 1443 1984
rect 1482 1950 1516 1984
rect 1555 1950 1589 1984
rect 1628 1950 1662 1984
rect 1701 1950 1735 1984
rect 1774 1950 1808 1984
rect 1847 1950 1881 1984
rect 1920 1950 1954 1984
rect 1993 1950 2027 1984
rect 2066 1950 2100 1984
rect 2139 1950 2173 1984
rect 2213 1950 2247 1984
rect 2287 1950 2321 1984
rect 2361 1950 2395 1984
rect 2435 1950 2469 1984
rect 2509 1950 2543 1984
rect 2583 1950 2617 1984
rect 2657 1950 2691 1984
rect 2731 1950 2765 1984
rect 2805 1950 2839 1984
rect 2879 1950 2913 1984
rect 2953 1950 2987 1984
rect 3027 1950 3061 1984
rect 3101 1950 3135 1984
rect 3175 1950 3209 1984
rect 3249 1950 3283 1984
rect 3323 1950 3357 1984
rect 3397 1950 3431 1984
rect 3471 1950 3505 1984
rect 3545 1950 3579 1984
rect 679 1878 713 1912
rect 752 1878 786 1912
rect 825 1878 859 1912
rect 898 1878 932 1912
rect 971 1878 1005 1912
rect 1044 1878 1078 1912
rect 1117 1878 1151 1912
rect 1190 1878 1224 1912
rect 1263 1878 1297 1912
rect 1336 1878 1370 1912
rect 1409 1878 1443 1912
rect 1482 1878 1516 1912
rect 1555 1878 1589 1912
rect 1628 1878 1662 1912
rect 1701 1878 1735 1912
rect 1774 1878 1808 1912
rect 1847 1878 1881 1912
rect 1920 1878 1954 1912
rect 1993 1878 2027 1912
rect 2066 1878 2100 1912
rect 2139 1878 2173 1912
rect 2213 1878 2247 1912
rect 2287 1878 2321 1912
rect 2361 1878 2395 1912
rect 2435 1878 2469 1912
rect 2509 1878 2543 1912
rect 2583 1878 2617 1912
rect 2657 1878 2691 1912
rect 2731 1878 2765 1912
rect 2805 1878 2839 1912
rect 2879 1878 2913 1912
rect 2953 1878 2987 1912
rect 3027 1878 3061 1912
rect 3101 1878 3135 1912
rect 3175 1878 3209 1912
rect 3249 1878 3283 1912
rect 3323 1878 3357 1912
rect 3397 1878 3431 1912
rect 3471 1878 3505 1912
rect 3545 1878 3579 1912
rect 3921 1950 3955 1984
rect 3995 1950 4029 1984
rect 4069 1950 4103 1984
rect 4143 1950 4177 1984
rect 4217 1950 4251 1984
rect 4291 1950 4325 1984
rect 4365 1950 4399 1984
rect 4439 1950 4473 1984
rect 4513 1950 4547 1984
rect 4587 1950 4621 1984
rect 4661 1950 4695 1984
rect 4735 1950 4769 1984
rect 4809 1950 4843 1984
rect 4883 1950 4917 1984
rect 4957 1950 4991 1984
rect 5031 1950 5065 1984
rect 5105 1950 5139 1984
rect 5179 1950 5213 1984
rect 5253 1950 5287 1984
rect 5327 1950 5361 1984
rect 5400 1950 5434 1984
rect 5473 1950 5507 1984
rect 5546 1950 5580 1984
rect 5619 1950 5653 1984
rect 5692 1950 5726 1984
rect 5765 1950 5799 1984
rect 5838 1950 5872 1984
rect 5911 1950 5945 1984
rect 5984 1950 6018 1984
rect 6057 1950 6091 1984
rect 6130 1950 6164 1984
rect 6203 1950 6237 1984
rect 6276 1950 6310 1984
rect 6349 1950 6383 1984
rect 6422 1950 6456 1984
rect 6495 1950 6529 1984
rect 6568 1950 6602 1984
rect 6641 1950 6675 1984
rect 6714 1950 6748 1984
rect 6787 1950 6821 1984
rect 3921 1878 3955 1912
rect 3995 1878 4029 1912
rect 4069 1878 4103 1912
rect 4143 1878 4177 1912
rect 4217 1878 4251 1912
rect 4291 1878 4325 1912
rect 4365 1878 4399 1912
rect 4439 1878 4473 1912
rect 4513 1878 4547 1912
rect 4587 1878 4621 1912
rect 4661 1878 4695 1912
rect 4735 1878 4769 1912
rect 4809 1878 4843 1912
rect 4883 1878 4917 1912
rect 4957 1878 4991 1912
rect 5031 1878 5065 1912
rect 5105 1878 5139 1912
rect 5179 1878 5213 1912
rect 5253 1878 5287 1912
rect 5327 1878 5361 1912
rect 5400 1878 5434 1912
rect 5473 1878 5507 1912
rect 5546 1878 5580 1912
rect 5619 1878 5653 1912
rect 5692 1878 5726 1912
rect 5765 1878 5799 1912
rect 5838 1878 5872 1912
rect 5911 1878 5945 1912
rect 5984 1878 6018 1912
rect 6057 1878 6091 1912
rect 6130 1878 6164 1912
rect 6203 1878 6237 1912
rect 6276 1878 6310 1912
rect 6349 1878 6383 1912
rect 6422 1878 6456 1912
rect 6495 1878 6529 1912
rect 6568 1878 6602 1912
rect 6641 1878 6675 1912
rect 6714 1878 6748 1912
rect 6787 1878 6821 1912
rect 7163 1950 7197 1984
rect 7236 1950 7270 1984
rect 7309 1950 7343 1984
rect 7382 1950 7416 1984
rect 7455 1950 7489 1984
rect 7528 1950 7562 1984
rect 7601 1950 7635 1984
rect 7674 1950 7708 1984
rect 7747 1950 7781 1984
rect 7820 1950 7854 1984
rect 7893 1950 7927 1984
rect 7966 1950 8000 1984
rect 8039 1950 8073 1984
rect 8112 1950 8146 1984
rect 8185 1950 8219 1984
rect 8258 1950 8292 1984
rect 8331 1950 8365 1984
rect 8404 1950 8438 1984
rect 8477 1950 8511 1984
rect 8550 1950 8584 1984
rect 8623 1950 8657 1984
rect 8697 1950 8731 1984
rect 8771 1950 8805 1984
rect 8845 1950 8879 1984
rect 8919 1950 8953 1984
rect 8993 1950 9027 1984
rect 9067 1950 9101 1984
rect 9141 1950 9175 1984
rect 9215 1950 9249 1984
rect 9289 1950 9323 1984
rect 9363 1950 9397 1984
rect 9437 1950 9471 1984
rect 9511 1950 9545 1984
rect 9585 1950 9619 1984
rect 9659 1950 9693 1984
rect 9733 1950 9767 1984
rect 9807 1950 9841 1984
rect 9881 1950 9915 1984
rect 9955 1950 9989 1984
rect 10029 1950 10063 1984
rect 7163 1878 7197 1912
rect 7236 1878 7270 1912
rect 7309 1878 7343 1912
rect 7382 1878 7416 1912
rect 7455 1878 7489 1912
rect 7528 1878 7562 1912
rect 7601 1878 7635 1912
rect 7674 1878 7708 1912
rect 7747 1878 7781 1912
rect 7820 1878 7854 1912
rect 7893 1878 7927 1912
rect 7966 1878 8000 1912
rect 8039 1878 8073 1912
rect 8112 1878 8146 1912
rect 8185 1878 8219 1912
rect 8258 1878 8292 1912
rect 8331 1878 8365 1912
rect 8404 1878 8438 1912
rect 8477 1878 8511 1912
rect 8550 1878 8584 1912
rect 8623 1878 8657 1912
rect 8697 1878 8731 1912
rect 8771 1878 8805 1912
rect 8845 1878 8879 1912
rect 8919 1878 8953 1912
rect 8993 1878 9027 1912
rect 9067 1878 9101 1912
rect 9141 1878 9175 1912
rect 9215 1878 9249 1912
rect 9289 1878 9323 1912
rect 9363 1878 9397 1912
rect 9437 1878 9471 1912
rect 9511 1878 9545 1912
rect 9585 1878 9619 1912
rect 9659 1878 9693 1912
rect 9733 1878 9767 1912
rect 9807 1878 9841 1912
rect 9881 1878 9915 1912
rect 9955 1878 9989 1912
rect 10029 1878 10063 1912
rect 10405 1950 10439 1984
rect 10479 1950 10513 1984
rect 10553 1950 10587 1984
rect 10627 1950 10661 1984
rect 10701 1950 10735 1984
rect 10775 1950 10809 1984
rect 10849 1950 10883 1984
rect 10923 1950 10957 1984
rect 10997 1950 11031 1984
rect 11071 1950 11105 1984
rect 11145 1950 11179 1984
rect 11219 1950 11253 1984
rect 11293 1950 11327 1984
rect 11367 1950 11401 1984
rect 11441 1950 11475 1984
rect 11515 1950 11549 1984
rect 11589 1950 11623 1984
rect 11663 1950 11697 1984
rect 11737 1950 11771 1984
rect 11811 1950 11845 1984
rect 11884 1950 11918 1984
rect 11957 1950 11991 1984
rect 12030 1950 12064 1984
rect 12103 1950 12137 1984
rect 12176 1950 12210 1984
rect 12249 1950 12283 1984
rect 12322 1950 12356 1984
rect 12395 1950 12429 1984
rect 12468 1950 12502 1984
rect 12541 1950 12575 1984
rect 12614 1950 12648 1984
rect 12687 1950 12721 1984
rect 12760 1950 12794 1984
rect 12833 1950 12867 1984
rect 12906 1950 12940 1984
rect 12979 1950 13013 1984
rect 13052 1950 13086 1984
rect 13125 1950 13159 1984
rect 13198 1950 13232 1984
rect 13271 1950 13305 1984
rect 10405 1878 10439 1912
rect 10479 1878 10513 1912
rect 10553 1878 10587 1912
rect 10627 1878 10661 1912
rect 10701 1878 10735 1912
rect 10775 1878 10809 1912
rect 10849 1878 10883 1912
rect 10923 1878 10957 1912
rect 10997 1878 11031 1912
rect 11071 1878 11105 1912
rect 11145 1878 11179 1912
rect 11219 1878 11253 1912
rect 11293 1878 11327 1912
rect 11367 1878 11401 1912
rect 11441 1878 11475 1912
rect 11515 1878 11549 1912
rect 11589 1878 11623 1912
rect 11663 1878 11697 1912
rect 11737 1878 11771 1912
rect 11811 1878 11845 1912
rect 11884 1878 11918 1912
rect 11957 1878 11991 1912
rect 12030 1878 12064 1912
rect 12103 1878 12137 1912
rect 12176 1878 12210 1912
rect 12249 1878 12283 1912
rect 12322 1878 12356 1912
rect 12395 1878 12429 1912
rect 12468 1878 12502 1912
rect 12541 1878 12575 1912
rect 12614 1878 12648 1912
rect 12687 1878 12721 1912
rect 12760 1878 12794 1912
rect 12833 1878 12867 1912
rect 12906 1878 12940 1912
rect 12979 1878 13013 1912
rect 13052 1878 13086 1912
rect 13125 1878 13159 1912
rect 13198 1878 13232 1912
rect 13271 1878 13305 1912
rect 13647 1950 13681 1984
rect 13720 1950 13754 1984
rect 13793 1950 13827 1984
rect 13866 1950 13900 1984
rect 13939 1950 13973 1984
rect 14012 1950 14046 1984
rect 14085 1950 14119 1984
rect 14158 1950 14192 1984
rect 14231 1950 14265 1984
rect 14304 1950 14338 1984
rect 14377 1950 14411 1984
rect 14450 1950 14484 1984
rect 14523 1950 14557 1984
rect 14596 1950 14630 1984
rect 14669 1950 14703 1984
rect 14742 1950 14776 1984
rect 14815 1950 14849 1984
rect 14888 1950 14922 1984
rect 14961 1950 14995 1984
rect 15034 1950 15068 1984
rect 15107 1950 15141 1984
rect 15181 1950 15215 1984
rect 15255 1950 15289 1984
rect 15329 1950 15363 1984
rect 15403 1950 15437 1984
rect 15477 1950 15511 1984
rect 15551 1950 15585 1984
rect 15625 1950 15659 1984
rect 15699 1950 15733 1984
rect 15773 1950 15807 1984
rect 15847 1950 15881 1984
rect 15921 1950 15955 1984
rect 15995 1950 16029 1984
rect 16069 1950 16103 1984
rect 16143 1950 16177 1984
rect 16217 1950 16251 1984
rect 16291 1950 16325 1984
rect 16365 1950 16399 1984
rect 16439 1950 16473 1984
rect 16513 1950 16547 1984
rect 13647 1878 13681 1912
rect 13720 1878 13754 1912
rect 13793 1878 13827 1912
rect 13866 1878 13900 1912
rect 13939 1878 13973 1912
rect 14012 1878 14046 1912
rect 14085 1878 14119 1912
rect 14158 1878 14192 1912
rect 14231 1878 14265 1912
rect 14304 1878 14338 1912
rect 14377 1878 14411 1912
rect 14450 1878 14484 1912
rect 14523 1878 14557 1912
rect 14596 1878 14630 1912
rect 14669 1878 14703 1912
rect 14742 1878 14776 1912
rect 14815 1878 14849 1912
rect 14888 1878 14922 1912
rect 14961 1878 14995 1912
rect 15034 1878 15068 1912
rect 15107 1878 15141 1912
rect 15181 1878 15215 1912
rect 15255 1878 15289 1912
rect 15329 1878 15363 1912
rect 15403 1878 15437 1912
rect 15477 1878 15511 1912
rect 15551 1878 15585 1912
rect 15625 1878 15659 1912
rect 15699 1878 15733 1912
rect 15773 1878 15807 1912
rect 15847 1878 15881 1912
rect 15921 1878 15955 1912
rect 15995 1878 16029 1912
rect 16069 1878 16103 1912
rect 16143 1878 16177 1912
rect 16217 1878 16251 1912
rect 16291 1878 16325 1912
rect 16365 1878 16399 1912
rect 16439 1878 16473 1912
rect 16513 1878 16547 1912
rect 16889 1950 16923 1984
rect 16963 1950 16997 1984
rect 17037 1950 17071 1984
rect 17111 1950 17145 1984
rect 17185 1950 17219 1984
rect 17259 1950 17293 1984
rect 17333 1950 17367 1984
rect 17407 1950 17441 1984
rect 17481 1950 17515 1984
rect 17555 1950 17589 1984
rect 17629 1950 17663 1984
rect 17703 1950 17737 1984
rect 17777 1950 17811 1984
rect 17851 1950 17885 1984
rect 17925 1950 17959 1984
rect 17999 1950 18033 1984
rect 18073 1950 18107 1984
rect 18147 1950 18181 1984
rect 18221 1950 18255 1984
rect 18295 1950 18329 1984
rect 18368 1950 18402 1984
rect 18441 1950 18475 1984
rect 18514 1950 18548 1984
rect 18587 1950 18621 1984
rect 18660 1950 18694 1984
rect 18733 1950 18767 1984
rect 18806 1950 18840 1984
rect 18879 1950 18913 1984
rect 18952 1950 18986 1984
rect 19025 1950 19059 1984
rect 19098 1950 19132 1984
rect 19171 1950 19205 1984
rect 19244 1950 19278 1984
rect 19317 1950 19351 1984
rect 19390 1950 19424 1984
rect 19463 1950 19497 1984
rect 19536 1950 19570 1984
rect 19609 1950 19643 1984
rect 19682 1950 19716 1984
rect 19755 1950 19789 1984
rect 16889 1878 16923 1912
rect 16963 1878 16997 1912
rect 17037 1878 17071 1912
rect 17111 1878 17145 1912
rect 17185 1878 17219 1912
rect 17259 1878 17293 1912
rect 17333 1878 17367 1912
rect 17407 1878 17441 1912
rect 17481 1878 17515 1912
rect 17555 1878 17589 1912
rect 17629 1878 17663 1912
rect 17703 1878 17737 1912
rect 17777 1878 17811 1912
rect 17851 1878 17885 1912
rect 17925 1878 17959 1912
rect 17999 1878 18033 1912
rect 18073 1878 18107 1912
rect 18147 1878 18181 1912
rect 18221 1878 18255 1912
rect 18295 1878 18329 1912
rect 18368 1878 18402 1912
rect 18441 1878 18475 1912
rect 18514 1878 18548 1912
rect 18587 1878 18621 1912
rect 18660 1878 18694 1912
rect 18733 1878 18767 1912
rect 18806 1878 18840 1912
rect 18879 1878 18913 1912
rect 18952 1878 18986 1912
rect 19025 1878 19059 1912
rect 19098 1878 19132 1912
rect 19171 1878 19205 1912
rect 19244 1878 19278 1912
rect 19317 1878 19351 1912
rect 19390 1878 19424 1912
rect 19463 1878 19497 1912
rect 19536 1878 19570 1912
rect 19609 1878 19643 1912
rect 19682 1878 19716 1912
rect 19755 1878 19789 1912
<< metal1 >>
rect 1109 4397 1115 4449
rect 1167 4397 6333 4449
rect 6385 4397 6400 4449
rect 6452 4397 6467 4449
rect 6519 4397 6534 4449
rect 6586 4397 6601 4449
rect 6653 4397 6668 4449
rect 6720 4397 7264 4449
rect 7316 4397 7331 4449
rect 7383 4397 7398 4449
rect 7450 4397 7465 4449
rect 7517 4397 7532 4449
rect 7584 4397 7599 4449
rect 7651 4397 12817 4449
rect 12869 4397 12884 4449
rect 12936 4397 12951 4449
rect 13003 4397 13018 4449
rect 13070 4397 13085 4449
rect 13137 4397 13152 4449
rect 13204 4397 13748 4449
rect 13800 4397 13815 4449
rect 13867 4397 13882 4449
rect 13934 4397 13949 4449
rect 14001 4397 14016 4449
rect 14068 4397 14083 4449
rect 14135 4397 19382 4449
rect 19434 4397 19467 4449
rect 19519 4397 19552 4449
rect 19604 4397 19636 4449
rect 19688 4397 19694 4449
rect 1109 4369 19694 4397
rect 1109 4317 1115 4369
rect 1167 4317 6333 4369
rect 6385 4317 6400 4369
rect 6452 4317 6467 4369
rect 6519 4317 6534 4369
rect 6586 4317 6601 4369
rect 6653 4317 6668 4369
rect 6720 4317 7264 4369
rect 7316 4317 7331 4369
rect 7383 4317 7398 4369
rect 7450 4317 7465 4369
rect 7517 4317 7532 4369
rect 7584 4317 7599 4369
rect 7651 4317 12817 4369
rect 12869 4317 12884 4369
rect 12936 4317 12951 4369
rect 13003 4317 13018 4369
rect 13070 4317 13085 4369
rect 13137 4317 13152 4369
rect 13204 4317 13748 4369
rect 13800 4317 13815 4369
rect 13867 4317 13882 4369
rect 13934 4317 13949 4369
rect 14001 4317 14016 4369
rect 14068 4317 14083 4369
rect 14135 4317 19382 4369
rect 19434 4317 19467 4369
rect 19519 4317 19552 4369
rect 19604 4317 19636 4369
rect 19688 4317 19694 4369
rect 6327 3009 6333 3061
rect 6385 3009 6400 3061
rect 6452 3009 6467 3061
rect 6519 3009 6534 3061
rect 6586 3009 6601 3061
rect 6653 3009 6668 3061
rect 6720 3009 6726 3061
rect 6327 2981 6726 3009
rect 6327 2929 6333 2981
rect 6385 2929 6400 2981
rect 6452 2929 6467 2981
rect 6519 2929 6534 2981
rect 6586 2929 6601 2981
rect 6653 2929 6668 2981
rect 6720 2929 6726 2981
rect 7258 3009 7264 3061
rect 7316 3009 7331 3061
rect 7383 3009 7398 3061
rect 7450 3009 7465 3061
rect 7517 3009 7532 3061
rect 7584 3009 7599 3061
rect 7651 3009 7657 3061
rect 7258 2981 7657 3009
rect 7258 2929 7264 2981
rect 7316 2929 7331 2981
rect 7383 2929 7398 2981
rect 7450 2929 7465 2981
rect 7517 2929 7532 2981
rect 7584 2929 7599 2981
rect 7651 2929 7657 2981
rect 12811 3009 12817 3061
rect 12869 3009 12884 3061
rect 12936 3009 12951 3061
rect 13003 3009 13018 3061
rect 13070 3009 13085 3061
rect 13137 3009 13152 3061
rect 13204 3009 13210 3061
rect 12811 2981 13210 3009
rect 12811 2929 12817 2981
rect 12869 2929 12884 2981
rect 12936 2929 12951 2981
rect 13003 2929 13018 2981
rect 13070 2929 13085 2981
rect 13137 2929 13152 2981
rect 13204 2929 13210 2981
rect 13742 3009 13748 3061
rect 13800 3009 13815 3061
rect 13867 3009 13882 3061
rect 13934 3009 13949 3061
rect 14001 3009 14016 3061
rect 14068 3009 14083 3061
rect 14135 3009 14141 3061
rect 13742 2981 14141 3009
rect 13742 2929 13748 2981
rect 13800 2929 13815 2981
rect 13867 2929 13882 2981
rect 13934 2929 13949 2981
rect 14001 2929 14016 2981
rect 14068 2929 14083 2981
rect 14135 2929 14141 2981
rect 19380 3009 19386 3061
rect 19438 3009 19470 3061
rect 19522 3009 19553 3061
rect 19605 3009 19636 3061
rect 19688 3009 19694 3061
rect 19380 2981 19694 3009
rect 19380 2929 19386 2981
rect 19438 2929 19470 2981
rect 19522 2929 19553 2981
rect 19605 2929 19636 2981
rect 19688 2929 19694 2981
tri 579 2808 626 2855 se
rect 626 2840 3632 2855
rect 626 2808 959 2840
rect 579 2774 679 2808
rect 713 2774 752 2808
rect 786 2774 825 2808
rect 859 2774 898 2808
rect 932 2788 959 2808
rect 1011 2788 1043 2840
rect 1095 2808 1127 2840
rect 1179 2808 1210 2840
rect 1262 2808 3632 2840
tri 3632 2808 3679 2855 sw
tri 3821 2808 3868 2855 se
rect 3868 2840 6874 2855
tri 6874 2840 6889 2855 sw
tri 7095 2840 7110 2855 se
rect 7110 2840 10116 2855
tri 10116 2840 10131 2855 sw
tri 10337 2840 10352 2855 se
rect 10352 2840 13358 2855
tri 13358 2840 13373 2855 sw
tri 13579 2840 13594 2855 se
rect 13594 2840 16600 2855
rect 3868 2808 6333 2840
rect 1095 2788 1117 2808
rect 1179 2788 1190 2808
rect 1262 2788 1263 2808
rect 932 2776 971 2788
rect 1005 2776 1044 2788
rect 1078 2776 1117 2788
rect 1151 2776 1190 2788
rect 1224 2776 1263 2788
rect 932 2774 959 2776
rect 579 2736 959 2774
rect 579 2702 679 2736
rect 713 2702 752 2736
rect 786 2702 825 2736
rect 859 2702 898 2736
rect 932 2724 959 2736
rect 1011 2724 1043 2776
rect 1095 2774 1117 2776
rect 1179 2774 1190 2776
rect 1262 2774 1263 2776
rect 1297 2774 1336 2808
rect 1370 2774 1409 2808
rect 1443 2774 1482 2808
rect 1516 2774 1555 2808
rect 1589 2774 1628 2808
rect 1662 2774 1701 2808
rect 1735 2774 1774 2808
rect 1808 2774 1847 2808
rect 1881 2774 1920 2808
rect 1954 2774 1993 2808
rect 2027 2774 2066 2808
rect 2100 2774 2139 2808
rect 2173 2774 2213 2808
rect 2247 2774 2287 2808
rect 2321 2774 2361 2808
rect 2395 2774 2435 2808
rect 2469 2774 2509 2808
rect 2543 2774 2583 2808
rect 2617 2774 2657 2808
rect 2691 2774 2731 2808
rect 2765 2774 2805 2808
rect 2839 2774 2879 2808
rect 2913 2774 2953 2808
rect 2987 2774 3027 2808
rect 3061 2774 3101 2808
rect 3135 2774 3175 2808
rect 3209 2774 3249 2808
rect 3283 2774 3323 2808
rect 3357 2774 3397 2808
rect 3431 2774 3471 2808
rect 3505 2774 3545 2808
rect 3579 2774 3921 2808
rect 3955 2774 3995 2808
rect 4029 2774 4069 2808
rect 4103 2774 4143 2808
rect 4177 2774 4217 2808
rect 4251 2774 4291 2808
rect 4325 2774 4365 2808
rect 4399 2774 4439 2808
rect 4473 2774 4513 2808
rect 4547 2774 4587 2808
rect 4621 2774 4661 2808
rect 4695 2774 4735 2808
rect 4769 2774 4809 2808
rect 4843 2774 4883 2808
rect 4917 2774 4957 2808
rect 4991 2774 5031 2808
rect 5065 2774 5105 2808
rect 5139 2774 5179 2808
rect 5213 2774 5253 2808
rect 5287 2774 5327 2808
rect 5361 2774 5400 2808
rect 5434 2774 5473 2808
rect 5507 2774 5546 2808
rect 5580 2774 5619 2808
rect 5653 2774 5692 2808
rect 5726 2774 5765 2808
rect 5799 2774 5838 2808
rect 5872 2774 5911 2808
rect 5945 2774 5984 2808
rect 6018 2774 6057 2808
rect 6091 2774 6130 2808
rect 6164 2774 6203 2808
rect 6237 2774 6276 2808
rect 6310 2788 6333 2808
rect 6385 2788 6400 2840
rect 6452 2808 6467 2840
rect 6519 2808 6534 2840
rect 6586 2808 6601 2840
rect 6653 2808 6668 2840
rect 6720 2808 6889 2840
tri 6889 2808 6921 2840 sw
tri 7063 2808 7095 2840 se
rect 7095 2808 7264 2840
rect 7316 2808 7331 2840
rect 7383 2808 7398 2840
rect 7450 2808 7465 2840
rect 7517 2808 7532 2840
rect 6456 2788 6467 2808
rect 6529 2788 6534 2808
rect 6310 2776 6349 2788
rect 6383 2776 6422 2788
rect 6456 2776 6495 2788
rect 6529 2776 6568 2788
rect 6602 2776 6641 2788
rect 6675 2776 6714 2788
rect 6310 2774 6333 2776
rect 1095 2736 1127 2774
rect 1179 2736 1210 2774
rect 1262 2736 6333 2774
rect 1095 2724 1117 2736
rect 1179 2724 1190 2736
rect 1262 2724 1263 2736
rect 932 2712 971 2724
rect 1005 2712 1044 2724
rect 1078 2712 1117 2724
rect 1151 2712 1190 2724
rect 1224 2712 1263 2724
rect 932 2702 959 2712
tri 579 2655 626 2702 ne
rect 626 2660 959 2702
rect 1011 2660 1043 2712
rect 1095 2702 1117 2712
rect 1179 2702 1190 2712
rect 1262 2702 1263 2712
rect 1297 2702 1336 2736
rect 1370 2702 1409 2736
rect 1443 2702 1482 2736
rect 1516 2702 1555 2736
rect 1589 2702 1628 2736
rect 1662 2702 1701 2736
rect 1735 2702 1774 2736
rect 1808 2702 1847 2736
rect 1881 2702 1920 2736
rect 1954 2702 1993 2736
rect 2027 2702 2066 2736
rect 2100 2702 2139 2736
rect 2173 2702 2213 2736
rect 2247 2702 2287 2736
rect 2321 2702 2361 2736
rect 2395 2702 2435 2736
rect 2469 2702 2509 2736
rect 2543 2702 2583 2736
rect 2617 2702 2657 2736
rect 2691 2702 2731 2736
rect 2765 2702 2805 2736
rect 2839 2702 2879 2736
rect 2913 2702 2953 2736
rect 2987 2702 3027 2736
rect 3061 2702 3101 2736
rect 3135 2702 3175 2736
rect 3209 2702 3249 2736
rect 3283 2702 3323 2736
rect 3357 2702 3397 2736
rect 3431 2702 3471 2736
rect 3505 2702 3545 2736
rect 3579 2702 3921 2736
rect 3955 2702 3995 2736
rect 4029 2702 4069 2736
rect 4103 2702 4143 2736
rect 4177 2702 4217 2736
rect 4251 2702 4291 2736
rect 4325 2702 4365 2736
rect 4399 2702 4439 2736
rect 4473 2702 4513 2736
rect 4547 2702 4587 2736
rect 4621 2702 4661 2736
rect 4695 2702 4735 2736
rect 4769 2702 4809 2736
rect 4843 2702 4883 2736
rect 4917 2702 4957 2736
rect 4991 2702 5031 2736
rect 5065 2702 5105 2736
rect 5139 2702 5179 2736
rect 5213 2702 5253 2736
rect 5287 2702 5327 2736
rect 5361 2702 5400 2736
rect 5434 2702 5473 2736
rect 5507 2702 5546 2736
rect 5580 2702 5619 2736
rect 5653 2702 5692 2736
rect 5726 2702 5765 2736
rect 5799 2702 5838 2736
rect 5872 2702 5911 2736
rect 5945 2702 5984 2736
rect 6018 2702 6057 2736
rect 6091 2702 6130 2736
rect 6164 2702 6203 2736
rect 6237 2702 6276 2736
rect 6310 2724 6333 2736
rect 6385 2724 6400 2776
rect 6456 2774 6467 2776
rect 6529 2774 6534 2776
rect 6748 2774 6787 2808
rect 6821 2774 7163 2808
rect 7197 2774 7236 2808
rect 7450 2788 7455 2808
rect 7517 2788 7528 2808
rect 7584 2788 7599 2840
rect 7651 2808 10131 2840
tri 10131 2808 10163 2840 sw
tri 10305 2808 10337 2840 se
rect 10337 2808 12817 2840
rect 7651 2788 7674 2808
rect 7270 2776 7309 2788
rect 7343 2776 7382 2788
rect 7416 2776 7455 2788
rect 7489 2776 7528 2788
rect 7562 2776 7601 2788
rect 7635 2776 7674 2788
rect 7450 2774 7455 2776
rect 7517 2774 7528 2776
rect 6452 2736 6467 2774
rect 6519 2736 6534 2774
rect 6586 2736 6601 2774
rect 6653 2736 6668 2774
rect 6720 2736 7264 2774
rect 7316 2736 7331 2774
rect 7383 2736 7398 2774
rect 7450 2736 7465 2774
rect 7517 2736 7532 2774
rect 6456 2724 6467 2736
rect 6529 2724 6534 2736
rect 6310 2712 6349 2724
rect 6383 2712 6422 2724
rect 6456 2712 6495 2724
rect 6529 2712 6568 2724
rect 6602 2712 6641 2724
rect 6675 2712 6714 2724
rect 6310 2702 6333 2712
rect 1095 2660 1127 2702
rect 1179 2660 1210 2702
rect 1262 2660 3632 2702
rect 626 2655 3632 2660
tri 3632 2655 3679 2702 nw
tri 3821 2655 3868 2702 ne
rect 3868 2660 6333 2702
rect 6385 2660 6400 2712
rect 6456 2702 6467 2712
rect 6529 2702 6534 2712
rect 6748 2702 6787 2736
rect 6821 2702 7163 2736
rect 7197 2702 7236 2736
rect 7450 2724 7455 2736
rect 7517 2724 7528 2736
rect 7584 2724 7599 2776
rect 7651 2774 7674 2776
rect 7708 2774 7747 2808
rect 7781 2774 7820 2808
rect 7854 2774 7893 2808
rect 7927 2774 7966 2808
rect 8000 2774 8039 2808
rect 8073 2774 8112 2808
rect 8146 2774 8185 2808
rect 8219 2774 8258 2808
rect 8292 2774 8331 2808
rect 8365 2774 8404 2808
rect 8438 2774 8477 2808
rect 8511 2774 8550 2808
rect 8584 2774 8623 2808
rect 8657 2774 8697 2808
rect 8731 2774 8771 2808
rect 8805 2774 8845 2808
rect 8879 2774 8919 2808
rect 8953 2774 8993 2808
rect 9027 2774 9067 2808
rect 9101 2774 9141 2808
rect 9175 2774 9215 2808
rect 9249 2774 9289 2808
rect 9323 2774 9363 2808
rect 9397 2774 9437 2808
rect 9471 2774 9511 2808
rect 9545 2774 9585 2808
rect 9619 2774 9659 2808
rect 9693 2774 9733 2808
rect 9767 2774 9807 2808
rect 9841 2774 9881 2808
rect 9915 2774 9955 2808
rect 9989 2774 10029 2808
rect 10063 2774 10405 2808
rect 10439 2774 10479 2808
rect 10513 2774 10553 2808
rect 10587 2774 10627 2808
rect 10661 2774 10701 2808
rect 10735 2774 10775 2808
rect 10809 2774 10849 2808
rect 10883 2774 10923 2808
rect 10957 2774 10997 2808
rect 11031 2774 11071 2808
rect 11105 2774 11145 2808
rect 11179 2774 11219 2808
rect 11253 2774 11293 2808
rect 11327 2774 11367 2808
rect 11401 2774 11441 2808
rect 11475 2774 11515 2808
rect 11549 2774 11589 2808
rect 11623 2774 11663 2808
rect 11697 2774 11737 2808
rect 11771 2774 11811 2808
rect 11845 2774 11884 2808
rect 11918 2774 11957 2808
rect 11991 2774 12030 2808
rect 12064 2774 12103 2808
rect 12137 2774 12176 2808
rect 12210 2774 12249 2808
rect 12283 2774 12322 2808
rect 12356 2774 12395 2808
rect 12429 2774 12468 2808
rect 12502 2774 12541 2808
rect 12575 2774 12614 2808
rect 12648 2774 12687 2808
rect 12721 2774 12760 2808
rect 12794 2788 12817 2808
rect 12869 2788 12884 2840
rect 12936 2808 12951 2840
rect 13003 2808 13018 2840
rect 13070 2808 13085 2840
rect 13137 2808 13152 2840
rect 13204 2808 13373 2840
tri 13373 2808 13405 2840 sw
tri 13547 2808 13579 2840 se
rect 13579 2808 13748 2840
rect 13800 2808 13815 2840
rect 13867 2808 13882 2840
rect 13934 2808 13949 2840
rect 14001 2808 14016 2840
rect 12940 2788 12951 2808
rect 13013 2788 13018 2808
rect 12794 2776 12833 2788
rect 12867 2776 12906 2788
rect 12940 2776 12979 2788
rect 13013 2776 13052 2788
rect 13086 2776 13125 2788
rect 13159 2776 13198 2788
rect 12794 2774 12817 2776
rect 7651 2736 12817 2774
rect 7651 2724 7674 2736
rect 7270 2712 7309 2724
rect 7343 2712 7382 2724
rect 7416 2712 7455 2724
rect 7489 2712 7528 2724
rect 7562 2712 7601 2724
rect 7635 2712 7674 2724
rect 7450 2702 7455 2712
rect 7517 2702 7528 2712
rect 6452 2660 6467 2702
rect 6519 2660 6534 2702
rect 6586 2660 6601 2702
rect 6653 2660 6668 2702
rect 6720 2660 6879 2702
tri 6879 2660 6921 2702 nw
tri 7063 2660 7105 2702 ne
rect 7105 2660 7264 2702
rect 7316 2660 7331 2702
rect 7383 2660 7398 2702
rect 7450 2660 7465 2702
rect 7517 2660 7532 2702
rect 7584 2660 7599 2712
rect 7651 2702 7674 2712
rect 7708 2702 7747 2736
rect 7781 2702 7820 2736
rect 7854 2702 7893 2736
rect 7927 2702 7966 2736
rect 8000 2702 8039 2736
rect 8073 2702 8112 2736
rect 8146 2702 8185 2736
rect 8219 2702 8258 2736
rect 8292 2702 8331 2736
rect 8365 2702 8404 2736
rect 8438 2702 8477 2736
rect 8511 2702 8550 2736
rect 8584 2702 8623 2736
rect 8657 2702 8697 2736
rect 8731 2702 8771 2736
rect 8805 2702 8845 2736
rect 8879 2702 8919 2736
rect 8953 2702 8993 2736
rect 9027 2702 9067 2736
rect 9101 2702 9141 2736
rect 9175 2702 9215 2736
rect 9249 2702 9289 2736
rect 9323 2702 9363 2736
rect 9397 2702 9437 2736
rect 9471 2702 9511 2736
rect 9545 2702 9585 2736
rect 9619 2702 9659 2736
rect 9693 2702 9733 2736
rect 9767 2702 9807 2736
rect 9841 2702 9881 2736
rect 9915 2702 9955 2736
rect 9989 2702 10029 2736
rect 10063 2702 10405 2736
rect 10439 2702 10479 2736
rect 10513 2702 10553 2736
rect 10587 2702 10627 2736
rect 10661 2702 10701 2736
rect 10735 2702 10775 2736
rect 10809 2702 10849 2736
rect 10883 2702 10923 2736
rect 10957 2702 10997 2736
rect 11031 2702 11071 2736
rect 11105 2702 11145 2736
rect 11179 2702 11219 2736
rect 11253 2702 11293 2736
rect 11327 2702 11367 2736
rect 11401 2702 11441 2736
rect 11475 2702 11515 2736
rect 11549 2702 11589 2736
rect 11623 2702 11663 2736
rect 11697 2702 11737 2736
rect 11771 2702 11811 2736
rect 11845 2702 11884 2736
rect 11918 2702 11957 2736
rect 11991 2702 12030 2736
rect 12064 2702 12103 2736
rect 12137 2702 12176 2736
rect 12210 2702 12249 2736
rect 12283 2702 12322 2736
rect 12356 2702 12395 2736
rect 12429 2702 12468 2736
rect 12502 2702 12541 2736
rect 12575 2702 12614 2736
rect 12648 2702 12687 2736
rect 12721 2702 12760 2736
rect 12794 2724 12817 2736
rect 12869 2724 12884 2776
rect 12940 2774 12951 2776
rect 13013 2774 13018 2776
rect 13232 2774 13271 2808
rect 13305 2774 13647 2808
rect 13681 2774 13720 2808
rect 13934 2788 13939 2808
rect 14001 2788 14012 2808
rect 14068 2788 14083 2840
rect 14135 2808 16600 2840
tri 16600 2808 16647 2855 sw
tri 16821 2840 16836 2855 se
rect 16836 2840 19842 2855
tri 19842 2840 19857 2855 sw
tri 16789 2808 16821 2840 se
rect 16821 2808 19386 2840
rect 19438 2808 19469 2840
rect 19521 2808 19552 2840
rect 19604 2808 19636 2840
rect 19688 2808 19857 2840
tri 19857 2808 19889 2840 sw
rect 14135 2788 14158 2808
rect 13754 2776 13793 2788
rect 13827 2776 13866 2788
rect 13900 2776 13939 2788
rect 13973 2776 14012 2788
rect 14046 2776 14085 2788
rect 14119 2776 14158 2788
rect 13934 2774 13939 2776
rect 14001 2774 14012 2776
rect 12936 2736 12951 2774
rect 13003 2736 13018 2774
rect 13070 2736 13085 2774
rect 13137 2736 13152 2774
rect 13204 2736 13748 2774
rect 13800 2736 13815 2774
rect 13867 2736 13882 2774
rect 13934 2736 13949 2774
rect 14001 2736 14016 2774
rect 12940 2724 12951 2736
rect 13013 2724 13018 2736
rect 12794 2712 12833 2724
rect 12867 2712 12906 2724
rect 12940 2712 12979 2724
rect 13013 2712 13052 2724
rect 13086 2712 13125 2724
rect 13159 2712 13198 2724
rect 12794 2702 12817 2712
rect 7651 2660 10121 2702
tri 10121 2660 10163 2702 nw
tri 10305 2660 10347 2702 ne
rect 10347 2660 12817 2702
rect 12869 2660 12884 2712
rect 12940 2702 12951 2712
rect 13013 2702 13018 2712
rect 13232 2702 13271 2736
rect 13305 2702 13647 2736
rect 13681 2702 13720 2736
rect 13934 2724 13939 2736
rect 14001 2724 14012 2736
rect 14068 2724 14083 2776
rect 14135 2774 14158 2776
rect 14192 2774 14231 2808
rect 14265 2774 14304 2808
rect 14338 2774 14377 2808
rect 14411 2774 14450 2808
rect 14484 2774 14523 2808
rect 14557 2774 14596 2808
rect 14630 2774 14669 2808
rect 14703 2774 14742 2808
rect 14776 2774 14815 2808
rect 14849 2774 14888 2808
rect 14922 2774 14961 2808
rect 14995 2774 15034 2808
rect 15068 2774 15107 2808
rect 15141 2774 15181 2808
rect 15215 2774 15255 2808
rect 15289 2774 15329 2808
rect 15363 2774 15403 2808
rect 15437 2774 15477 2808
rect 15511 2774 15551 2808
rect 15585 2774 15625 2808
rect 15659 2774 15699 2808
rect 15733 2774 15773 2808
rect 15807 2774 15847 2808
rect 15881 2774 15921 2808
rect 15955 2774 15995 2808
rect 16029 2774 16069 2808
rect 16103 2774 16143 2808
rect 16177 2774 16217 2808
rect 16251 2774 16291 2808
rect 16325 2774 16365 2808
rect 16399 2774 16439 2808
rect 16473 2774 16513 2808
rect 16547 2774 16889 2808
rect 16923 2774 16963 2808
rect 16997 2774 17037 2808
rect 17071 2774 17111 2808
rect 17145 2774 17185 2808
rect 17219 2774 17259 2808
rect 17293 2774 17333 2808
rect 17367 2774 17407 2808
rect 17441 2774 17481 2808
rect 17515 2774 17555 2808
rect 17589 2774 17629 2808
rect 17663 2774 17703 2808
rect 17737 2774 17777 2808
rect 17811 2774 17851 2808
rect 17885 2774 17925 2808
rect 17959 2774 17999 2808
rect 18033 2774 18073 2808
rect 18107 2774 18147 2808
rect 18181 2774 18221 2808
rect 18255 2774 18295 2808
rect 18329 2774 18368 2808
rect 18402 2774 18441 2808
rect 18475 2774 18514 2808
rect 18548 2774 18587 2808
rect 18621 2774 18660 2808
rect 18694 2774 18733 2808
rect 18767 2774 18806 2808
rect 18840 2774 18879 2808
rect 18913 2774 18952 2808
rect 18986 2774 19025 2808
rect 19059 2774 19098 2808
rect 19132 2774 19171 2808
rect 19205 2774 19244 2808
rect 19278 2774 19317 2808
rect 19351 2788 19386 2808
rect 19438 2788 19463 2808
rect 19521 2788 19536 2808
rect 19604 2788 19609 2808
rect 19351 2776 19390 2788
rect 19424 2776 19463 2788
rect 19497 2776 19536 2788
rect 19570 2776 19609 2788
rect 19643 2776 19682 2788
rect 19351 2774 19386 2776
rect 19438 2774 19463 2776
rect 19521 2774 19536 2776
rect 19604 2774 19609 2776
rect 19716 2774 19755 2808
rect 19789 2774 19889 2808
rect 14135 2736 19386 2774
rect 19438 2736 19469 2774
rect 19521 2736 19552 2774
rect 19604 2736 19636 2774
rect 19688 2736 19889 2774
rect 14135 2724 14158 2736
rect 13754 2712 13793 2724
rect 13827 2712 13866 2724
rect 13900 2712 13939 2724
rect 13973 2712 14012 2724
rect 14046 2712 14085 2724
rect 14119 2712 14158 2724
rect 13934 2702 13939 2712
rect 14001 2702 14012 2712
rect 12936 2660 12951 2702
rect 13003 2660 13018 2702
rect 13070 2660 13085 2702
rect 13137 2660 13152 2702
rect 13204 2660 13363 2702
tri 13363 2660 13405 2702 nw
tri 13547 2660 13589 2702 ne
rect 13589 2660 13748 2702
rect 13800 2660 13815 2702
rect 13867 2660 13882 2702
rect 13934 2660 13949 2702
rect 14001 2660 14016 2702
rect 14068 2660 14083 2712
rect 14135 2702 14158 2712
rect 14192 2702 14231 2736
rect 14265 2702 14304 2736
rect 14338 2702 14377 2736
rect 14411 2702 14450 2736
rect 14484 2702 14523 2736
rect 14557 2702 14596 2736
rect 14630 2702 14669 2736
rect 14703 2702 14742 2736
rect 14776 2702 14815 2736
rect 14849 2702 14888 2736
rect 14922 2702 14961 2736
rect 14995 2702 15034 2736
rect 15068 2702 15107 2736
rect 15141 2702 15181 2736
rect 15215 2702 15255 2736
rect 15289 2702 15329 2736
rect 15363 2702 15403 2736
rect 15437 2702 15477 2736
rect 15511 2702 15551 2736
rect 15585 2702 15625 2736
rect 15659 2702 15699 2736
rect 15733 2702 15773 2736
rect 15807 2702 15847 2736
rect 15881 2702 15921 2736
rect 15955 2702 15995 2736
rect 16029 2702 16069 2736
rect 16103 2702 16143 2736
rect 16177 2702 16217 2736
rect 16251 2702 16291 2736
rect 16325 2702 16365 2736
rect 16399 2702 16439 2736
rect 16473 2702 16513 2736
rect 16547 2702 16889 2736
rect 16923 2702 16963 2736
rect 16997 2702 17037 2736
rect 17071 2702 17111 2736
rect 17145 2702 17185 2736
rect 17219 2702 17259 2736
rect 17293 2702 17333 2736
rect 17367 2702 17407 2736
rect 17441 2702 17481 2736
rect 17515 2702 17555 2736
rect 17589 2702 17629 2736
rect 17663 2702 17703 2736
rect 17737 2702 17777 2736
rect 17811 2702 17851 2736
rect 17885 2702 17925 2736
rect 17959 2702 17999 2736
rect 18033 2702 18073 2736
rect 18107 2702 18147 2736
rect 18181 2702 18221 2736
rect 18255 2702 18295 2736
rect 18329 2702 18368 2736
rect 18402 2702 18441 2736
rect 18475 2702 18514 2736
rect 18548 2702 18587 2736
rect 18621 2702 18660 2736
rect 18694 2702 18733 2736
rect 18767 2702 18806 2736
rect 18840 2702 18879 2736
rect 18913 2702 18952 2736
rect 18986 2702 19025 2736
rect 19059 2702 19098 2736
rect 19132 2702 19171 2736
rect 19205 2702 19244 2736
rect 19278 2702 19317 2736
rect 19351 2724 19386 2736
rect 19438 2724 19463 2736
rect 19521 2724 19536 2736
rect 19604 2724 19609 2736
rect 19351 2712 19390 2724
rect 19424 2712 19463 2724
rect 19497 2712 19536 2724
rect 19570 2712 19609 2724
rect 19643 2712 19682 2724
rect 19351 2702 19386 2712
rect 19438 2702 19463 2712
rect 19521 2702 19536 2712
rect 19604 2702 19609 2712
rect 19716 2702 19755 2736
rect 19789 2702 19889 2736
rect 14135 2660 16600 2702
rect 3868 2655 6874 2660
tri 6874 2655 6879 2660 nw
tri 7105 2655 7110 2660 ne
rect 7110 2655 10116 2660
tri 10116 2655 10121 2660 nw
tri 10347 2655 10352 2660 ne
rect 10352 2655 13358 2660
tri 13358 2655 13363 2660 nw
tri 13589 2655 13594 2660 ne
rect 13594 2655 16600 2660
tri 16600 2655 16647 2702 nw
tri 16789 2660 16831 2702 ne
rect 16831 2660 19386 2702
rect 19438 2660 19469 2702
rect 19521 2660 19552 2702
rect 19604 2660 19636 2702
rect 19688 2660 19847 2702
tri 19847 2660 19889 2702 nw
tri 16831 2655 16836 2660 ne
rect 16836 2655 19842 2660
tri 19842 2655 19847 2660 nw
rect 471 2614 16697 2620
rect 471 2580 483 2614
rect 517 2580 555 2614
rect 589 2580 3701 2614
rect 3735 2580 3773 2614
rect 3807 2580 6943 2614
rect 6977 2580 7015 2614
rect 7049 2580 10185 2614
rect 10219 2580 10257 2614
rect 10291 2580 13451 2614
rect 13485 2580 13523 2614
rect 13557 2580 16697 2614
rect 19931 2613 19977 2615
rect 471 2574 16697 2580
rect 19925 2607 19977 2613
rect 471 2569 552 2574
tri 552 2569 557 2574 nw
rect 471 2194 532 2569
tri 532 2549 552 2569 nw
rect 19925 2543 19977 2555
tri 614 2531 626 2543 se
rect 626 2539 3604 2543
rect 626 2531 1342 2539
tri 580 2497 614 2531 se
rect 614 2497 1342 2531
rect 0 2188 230 2194
rect 52 2136 178 2188
rect 0 2124 230 2136
rect 52 2072 178 2124
rect 0 2066 230 2072
rect 459 2188 532 2194
rect 511 2143 532 2188
tri 579 2496 580 2497 se
rect 580 2496 1342 2497
rect 579 2487 1342 2496
rect 1394 2487 1407 2539
rect 1459 2487 1472 2539
rect 1524 2487 1537 2539
rect 1589 2487 1601 2539
rect 1653 2487 1665 2539
rect 1717 2487 1729 2539
rect 1781 2487 1793 2539
rect 1845 2487 1857 2539
rect 1909 2487 1921 2539
rect 1973 2487 1985 2539
rect 2037 2487 2049 2539
rect 2101 2487 2113 2539
rect 2165 2487 2177 2539
rect 2229 2531 3604 2539
tri 3604 2531 3616 2543 sw
tri 3888 2531 3900 2543 se
rect 3900 2539 6842 2543
rect 3900 2531 5271 2539
rect 2229 2497 3616 2531
tri 3616 2497 3650 2531 sw
tri 3854 2497 3888 2531 se
rect 3888 2497 5271 2531
rect 2229 2496 3650 2497
tri 3650 2496 3651 2497 sw
tri 3853 2496 3854 2497 se
rect 3854 2496 5271 2497
rect 2229 2487 5271 2496
rect 5323 2487 5335 2539
rect 5387 2487 5399 2539
rect 5451 2487 5463 2539
rect 5515 2487 5527 2539
rect 5579 2487 5591 2539
rect 5643 2487 5655 2539
rect 5707 2487 5719 2539
rect 5771 2487 5783 2539
rect 5835 2487 5847 2539
rect 5899 2487 5911 2539
rect 5963 2487 5976 2539
rect 6028 2487 6041 2539
rect 6093 2487 6106 2539
rect 6158 2531 6842 2539
tri 6842 2531 6854 2543 sw
tri 7124 2531 7136 2543 se
rect 7136 2539 10075 2543
rect 7136 2531 7826 2539
rect 6158 2497 6854 2531
tri 6854 2497 6888 2531 sw
tri 7090 2497 7124 2531 se
rect 7124 2497 7826 2531
rect 6158 2496 6888 2497
tri 6888 2496 6889 2497 sw
tri 7089 2496 7090 2497 se
rect 7090 2496 7826 2497
rect 6158 2487 7826 2496
rect 7878 2487 7891 2539
rect 7943 2487 7956 2539
rect 8008 2487 8021 2539
rect 8073 2487 8085 2539
rect 8137 2487 8149 2539
rect 8201 2487 8213 2539
rect 8265 2487 8277 2539
rect 8329 2487 8341 2539
rect 8393 2487 8405 2539
rect 8457 2487 8469 2539
rect 8521 2487 8533 2539
rect 8585 2487 8597 2539
rect 8649 2487 8661 2539
rect 8713 2531 10075 2539
tri 10075 2531 10087 2543 sw
tri 10357 2531 10369 2543 se
rect 10369 2539 13329 2543
rect 10369 2531 11755 2539
rect 8713 2497 10087 2531
tri 10087 2497 10121 2531 sw
tri 10323 2497 10357 2531 se
rect 10357 2497 11755 2531
rect 8713 2496 10121 2497
tri 10121 2496 10122 2497 sw
tri 10322 2496 10323 2497 se
rect 10323 2496 11755 2497
rect 8713 2487 11755 2496
rect 11807 2487 11819 2539
rect 11871 2487 11883 2539
rect 11935 2487 11947 2539
rect 11999 2487 12011 2539
rect 12063 2487 12075 2539
rect 12127 2487 12139 2539
rect 12191 2487 12203 2539
rect 12255 2487 12267 2539
rect 12319 2487 12331 2539
rect 12383 2487 12395 2539
rect 12447 2487 12460 2539
rect 12512 2487 12525 2539
rect 12577 2487 12590 2539
rect 12642 2531 13329 2539
tri 13329 2531 13341 2543 sw
tri 13612 2531 13624 2543 se
rect 13624 2539 16566 2543
rect 13624 2531 14310 2539
rect 12642 2497 13341 2531
tri 13341 2497 13375 2531 sw
tri 13578 2497 13612 2531 se
rect 13612 2497 14310 2531
rect 12642 2496 13375 2497
tri 13375 2496 13376 2497 sw
tri 13577 2496 13578 2497 se
rect 13578 2496 14310 2497
rect 12642 2487 14310 2496
rect 14362 2487 14375 2539
rect 14427 2487 14440 2539
rect 14492 2487 14505 2539
rect 14557 2487 14569 2539
rect 14621 2487 14633 2539
rect 14685 2487 14697 2539
rect 14749 2487 14761 2539
rect 14813 2487 14825 2539
rect 14877 2487 14889 2539
rect 14941 2487 14953 2539
rect 15005 2487 15017 2539
rect 15069 2487 15081 2539
rect 15133 2487 15145 2539
rect 15197 2531 16566 2539
tri 16566 2531 16578 2543 sw
tri 16848 2531 16860 2543 se
rect 16860 2539 19842 2543
rect 16860 2531 18239 2539
rect 15197 2497 16578 2531
tri 16578 2497 16612 2531 sw
tri 16814 2497 16848 2531 se
rect 16848 2497 18239 2531
rect 15197 2496 16612 2497
tri 16612 2496 16613 2497 sw
tri 16813 2496 16814 2497 se
rect 16814 2496 18239 2497
rect 15197 2487 18239 2496
rect 18291 2487 18303 2539
rect 18355 2487 18367 2539
rect 18419 2487 18431 2539
rect 18483 2487 18495 2539
rect 18547 2487 18559 2539
rect 18611 2487 18623 2539
rect 18675 2487 18687 2539
rect 18739 2487 18751 2539
rect 18803 2487 18815 2539
rect 18867 2487 18879 2539
rect 18931 2487 18944 2539
rect 18996 2487 19009 2539
rect 19061 2487 19074 2539
rect 19126 2531 19842 2539
tri 19842 2531 19854 2543 sw
rect 19126 2497 19854 2531
tri 19854 2497 19888 2531 sw
rect 19126 2496 19888 2497
tri 19888 2496 19889 2497 sw
rect 19126 2487 19889 2496
rect 579 2471 19889 2487
rect 579 2419 1342 2471
rect 1394 2419 1407 2471
rect 1459 2419 1472 2471
rect 1524 2419 1537 2471
rect 1589 2419 1601 2471
rect 1653 2419 1665 2471
rect 1717 2419 1729 2471
rect 1781 2419 1793 2471
rect 1845 2419 1857 2471
rect 1909 2419 1921 2471
rect 1973 2419 1985 2471
rect 2037 2419 2049 2471
rect 2101 2419 2113 2471
rect 2165 2419 2177 2471
rect 2229 2419 5271 2471
rect 5323 2419 5335 2471
rect 5387 2419 5399 2471
rect 5451 2419 5463 2471
rect 5515 2419 5527 2471
rect 5579 2419 5591 2471
rect 5643 2419 5655 2471
rect 5707 2419 5719 2471
rect 5771 2419 5783 2471
rect 5835 2419 5847 2471
rect 5899 2419 5911 2471
rect 5963 2419 5976 2471
rect 6028 2419 6041 2471
rect 6093 2419 6106 2471
rect 6158 2419 7826 2471
rect 7878 2419 7891 2471
rect 7943 2419 7956 2471
rect 8008 2419 8021 2471
rect 8073 2419 8085 2471
rect 8137 2419 8149 2471
rect 8201 2419 8213 2471
rect 8265 2419 8277 2471
rect 8329 2419 8341 2471
rect 8393 2419 8405 2471
rect 8457 2419 8469 2471
rect 8521 2419 8533 2471
rect 8585 2419 8597 2471
rect 8649 2419 8661 2471
rect 8713 2419 11755 2471
rect 11807 2419 11819 2471
rect 11871 2419 11883 2471
rect 11935 2419 11947 2471
rect 11999 2419 12011 2471
rect 12063 2419 12075 2471
rect 12127 2419 12139 2471
rect 12191 2419 12203 2471
rect 12255 2419 12267 2471
rect 12319 2419 12331 2471
rect 12383 2419 12395 2471
rect 12447 2419 12460 2471
rect 12512 2419 12525 2471
rect 12577 2419 12590 2471
rect 12642 2419 14310 2471
rect 14362 2419 14375 2471
rect 14427 2419 14440 2471
rect 14492 2419 14505 2471
rect 14557 2419 14569 2471
rect 14621 2419 14633 2471
rect 14685 2419 14697 2471
rect 14749 2419 14761 2471
rect 14813 2419 14825 2471
rect 14877 2419 14889 2471
rect 14941 2419 14953 2471
rect 15005 2419 15017 2471
rect 15069 2419 15081 2471
rect 15133 2419 15145 2471
rect 15197 2419 18239 2471
rect 18291 2419 18303 2471
rect 18355 2419 18367 2471
rect 18419 2419 18431 2471
rect 18483 2419 18495 2471
rect 18547 2419 18559 2471
rect 18611 2419 18623 2471
rect 18675 2419 18687 2471
rect 18739 2419 18751 2471
rect 18803 2419 18815 2471
rect 18867 2419 18879 2471
rect 18931 2419 18944 2471
rect 18996 2419 19009 2471
rect 19061 2419 19074 2471
rect 19126 2419 19889 2471
rect 579 2403 19889 2419
rect 579 2396 1342 2403
rect 579 2362 679 2396
rect 713 2362 752 2396
rect 786 2362 825 2396
rect 859 2362 898 2396
rect 932 2362 971 2396
rect 1005 2362 1044 2396
rect 1078 2362 1117 2396
rect 1151 2362 1190 2396
rect 1224 2362 1263 2396
rect 1297 2362 1336 2396
rect 579 2351 1342 2362
rect 1394 2351 1407 2403
rect 1459 2351 1472 2403
rect 1524 2351 1537 2403
rect 1589 2351 1601 2403
rect 1653 2396 1665 2403
rect 1717 2396 1729 2403
rect 1781 2396 1793 2403
rect 1845 2396 1857 2403
rect 1909 2396 1921 2403
rect 1662 2362 1665 2396
rect 1845 2362 1847 2396
rect 1909 2362 1920 2396
rect 1653 2351 1665 2362
rect 1717 2351 1729 2362
rect 1781 2351 1793 2362
rect 1845 2351 1857 2362
rect 1909 2351 1921 2362
rect 1973 2351 1985 2403
rect 2037 2351 2049 2403
rect 2101 2351 2113 2403
rect 2165 2396 2177 2403
rect 2229 2396 5271 2403
rect 5323 2396 5335 2403
rect 2173 2362 2177 2396
rect 2247 2362 2287 2396
rect 2321 2362 2361 2396
rect 2395 2362 2435 2396
rect 2469 2362 2509 2396
rect 2543 2362 2583 2396
rect 2617 2362 2657 2396
rect 2691 2362 2731 2396
rect 2765 2362 2805 2396
rect 2839 2362 2879 2396
rect 2913 2362 2953 2396
rect 2987 2362 3027 2396
rect 3061 2362 3101 2396
rect 3135 2362 3175 2396
rect 3209 2362 3249 2396
rect 3283 2362 3323 2396
rect 3357 2362 3397 2396
rect 3431 2362 3471 2396
rect 3505 2362 3545 2396
rect 3579 2362 3921 2396
rect 3955 2362 3995 2396
rect 4029 2362 4069 2396
rect 4103 2362 4143 2396
rect 4177 2362 4217 2396
rect 4251 2362 4291 2396
rect 4325 2362 4365 2396
rect 4399 2362 4439 2396
rect 4473 2362 4513 2396
rect 4547 2362 4587 2396
rect 4621 2362 4661 2396
rect 4695 2362 4735 2396
rect 4769 2362 4809 2396
rect 4843 2362 4883 2396
rect 4917 2362 4957 2396
rect 4991 2362 5031 2396
rect 5065 2362 5105 2396
rect 5139 2362 5179 2396
rect 5213 2362 5253 2396
rect 5323 2362 5327 2396
rect 2165 2351 2177 2362
rect 2229 2351 5271 2362
rect 5323 2351 5335 2362
rect 5387 2351 5399 2403
rect 5451 2351 5463 2403
rect 5515 2351 5527 2403
rect 5579 2396 5591 2403
rect 5643 2396 5655 2403
rect 5707 2396 5719 2403
rect 5771 2396 5783 2403
rect 5835 2396 5847 2403
rect 5580 2362 5591 2396
rect 5653 2362 5655 2396
rect 5835 2362 5838 2396
rect 5579 2351 5591 2362
rect 5643 2351 5655 2362
rect 5707 2351 5719 2362
rect 5771 2351 5783 2362
rect 5835 2351 5847 2362
rect 5899 2351 5911 2403
rect 5963 2351 5976 2403
rect 6028 2351 6041 2403
rect 6093 2351 6106 2403
rect 6158 2396 7826 2403
rect 6164 2362 6203 2396
rect 6237 2362 6276 2396
rect 6310 2362 6349 2396
rect 6383 2362 6422 2396
rect 6456 2362 6495 2396
rect 6529 2362 6568 2396
rect 6602 2362 6641 2396
rect 6675 2362 6714 2396
rect 6748 2362 6787 2396
rect 6821 2362 7163 2396
rect 7197 2362 7236 2396
rect 7270 2362 7309 2396
rect 7343 2362 7382 2396
rect 7416 2362 7455 2396
rect 7489 2362 7528 2396
rect 7562 2362 7601 2396
rect 7635 2362 7674 2396
rect 7708 2362 7747 2396
rect 7781 2362 7820 2396
rect 6158 2351 7826 2362
rect 7878 2351 7891 2403
rect 7943 2351 7956 2403
rect 8008 2351 8021 2403
rect 8073 2351 8085 2403
rect 8137 2396 8149 2403
rect 8201 2396 8213 2403
rect 8265 2396 8277 2403
rect 8329 2396 8341 2403
rect 8393 2396 8405 2403
rect 8146 2362 8149 2396
rect 8329 2362 8331 2396
rect 8393 2362 8404 2396
rect 8137 2351 8149 2362
rect 8201 2351 8213 2362
rect 8265 2351 8277 2362
rect 8329 2351 8341 2362
rect 8393 2351 8405 2362
rect 8457 2351 8469 2403
rect 8521 2351 8533 2403
rect 8585 2351 8597 2403
rect 8649 2396 8661 2403
rect 8713 2396 11755 2403
rect 11807 2396 11819 2403
rect 8657 2362 8661 2396
rect 8731 2362 8771 2396
rect 8805 2362 8845 2396
rect 8879 2362 8919 2396
rect 8953 2362 8993 2396
rect 9027 2362 9067 2396
rect 9101 2362 9141 2396
rect 9175 2362 9215 2396
rect 9249 2362 9289 2396
rect 9323 2362 9363 2396
rect 9397 2362 9437 2396
rect 9471 2362 9511 2396
rect 9545 2362 9585 2396
rect 9619 2362 9659 2396
rect 9693 2362 9733 2396
rect 9767 2362 9807 2396
rect 9841 2362 9881 2396
rect 9915 2362 9955 2396
rect 9989 2362 10029 2396
rect 10063 2362 10405 2396
rect 10439 2362 10479 2396
rect 10513 2362 10553 2396
rect 10587 2362 10627 2396
rect 10661 2362 10701 2396
rect 10735 2362 10775 2396
rect 10809 2362 10849 2396
rect 10883 2362 10923 2396
rect 10957 2362 10997 2396
rect 11031 2362 11071 2396
rect 11105 2362 11145 2396
rect 11179 2362 11219 2396
rect 11253 2362 11293 2396
rect 11327 2362 11367 2396
rect 11401 2362 11441 2396
rect 11475 2362 11515 2396
rect 11549 2362 11589 2396
rect 11623 2362 11663 2396
rect 11697 2362 11737 2396
rect 11807 2362 11811 2396
rect 8649 2351 8661 2362
rect 8713 2351 11755 2362
rect 11807 2351 11819 2362
rect 11871 2351 11883 2403
rect 11935 2351 11947 2403
rect 11999 2351 12011 2403
rect 12063 2396 12075 2403
rect 12127 2396 12139 2403
rect 12191 2396 12203 2403
rect 12255 2396 12267 2403
rect 12319 2396 12331 2403
rect 12064 2362 12075 2396
rect 12137 2362 12139 2396
rect 12319 2362 12322 2396
rect 12063 2351 12075 2362
rect 12127 2351 12139 2362
rect 12191 2351 12203 2362
rect 12255 2351 12267 2362
rect 12319 2351 12331 2362
rect 12383 2351 12395 2403
rect 12447 2351 12460 2403
rect 12512 2351 12525 2403
rect 12577 2351 12590 2403
rect 12642 2396 14310 2403
rect 12648 2362 12687 2396
rect 12721 2362 12760 2396
rect 12794 2362 12833 2396
rect 12867 2362 12906 2396
rect 12940 2362 12979 2396
rect 13013 2362 13052 2396
rect 13086 2362 13125 2396
rect 13159 2362 13198 2396
rect 13232 2362 13271 2396
rect 13305 2362 13647 2396
rect 13681 2362 13720 2396
rect 13754 2362 13793 2396
rect 13827 2362 13866 2396
rect 13900 2362 13939 2396
rect 13973 2362 14012 2396
rect 14046 2362 14085 2396
rect 14119 2362 14158 2396
rect 14192 2362 14231 2396
rect 14265 2362 14304 2396
rect 12642 2351 14310 2362
rect 14362 2351 14375 2403
rect 14427 2351 14440 2403
rect 14492 2351 14505 2403
rect 14557 2351 14569 2403
rect 14621 2396 14633 2403
rect 14685 2396 14697 2403
rect 14749 2396 14761 2403
rect 14813 2396 14825 2403
rect 14877 2396 14889 2403
rect 14630 2362 14633 2396
rect 14813 2362 14815 2396
rect 14877 2362 14888 2396
rect 14621 2351 14633 2362
rect 14685 2351 14697 2362
rect 14749 2351 14761 2362
rect 14813 2351 14825 2362
rect 14877 2351 14889 2362
rect 14941 2351 14953 2403
rect 15005 2351 15017 2403
rect 15069 2351 15081 2403
rect 15133 2396 15145 2403
rect 15197 2396 18239 2403
rect 18291 2396 18303 2403
rect 15141 2362 15145 2396
rect 15215 2362 15255 2396
rect 15289 2362 15329 2396
rect 15363 2362 15403 2396
rect 15437 2362 15477 2396
rect 15511 2362 15551 2396
rect 15585 2362 15625 2396
rect 15659 2362 15699 2396
rect 15733 2362 15773 2396
rect 15807 2362 15847 2396
rect 15881 2362 15921 2396
rect 15955 2362 15995 2396
rect 16029 2362 16069 2396
rect 16103 2362 16143 2396
rect 16177 2362 16217 2396
rect 16251 2362 16291 2396
rect 16325 2362 16365 2396
rect 16399 2362 16439 2396
rect 16473 2362 16513 2396
rect 16547 2362 16889 2396
rect 16923 2362 16963 2396
rect 16997 2362 17037 2396
rect 17071 2362 17111 2396
rect 17145 2362 17185 2396
rect 17219 2362 17259 2396
rect 17293 2362 17333 2396
rect 17367 2362 17407 2396
rect 17441 2362 17481 2396
rect 17515 2362 17555 2396
rect 17589 2362 17629 2396
rect 17663 2362 17703 2396
rect 17737 2362 17777 2396
rect 17811 2362 17851 2396
rect 17885 2362 17925 2396
rect 17959 2362 17999 2396
rect 18033 2362 18073 2396
rect 18107 2362 18147 2396
rect 18181 2362 18221 2396
rect 18291 2362 18295 2396
rect 15133 2351 15145 2362
rect 15197 2351 18239 2362
rect 18291 2351 18303 2362
rect 18355 2351 18367 2403
rect 18419 2351 18431 2403
rect 18483 2351 18495 2403
rect 18547 2396 18559 2403
rect 18611 2396 18623 2403
rect 18675 2396 18687 2403
rect 18739 2396 18751 2403
rect 18803 2396 18815 2403
rect 18548 2362 18559 2396
rect 18621 2362 18623 2396
rect 18803 2362 18806 2396
rect 18547 2351 18559 2362
rect 18611 2351 18623 2362
rect 18675 2351 18687 2362
rect 18739 2351 18751 2362
rect 18803 2351 18815 2362
rect 18867 2351 18879 2403
rect 18931 2351 18944 2403
rect 18996 2351 19009 2403
rect 19061 2351 19074 2403
rect 19126 2396 19889 2403
rect 19132 2362 19171 2396
rect 19205 2362 19244 2396
rect 19278 2362 19317 2396
rect 19351 2362 19390 2396
rect 19424 2362 19463 2396
rect 19497 2362 19536 2396
rect 19570 2362 19609 2396
rect 19643 2362 19682 2396
rect 19716 2362 19755 2396
rect 19789 2362 19889 2396
rect 19126 2351 19889 2362
rect 579 2335 19889 2351
rect 579 2324 1342 2335
rect 579 2290 679 2324
rect 713 2290 752 2324
rect 786 2290 825 2324
rect 859 2290 898 2324
rect 932 2290 971 2324
rect 1005 2290 1044 2324
rect 1078 2290 1117 2324
rect 1151 2290 1190 2324
rect 1224 2290 1263 2324
rect 1297 2290 1336 2324
rect 579 2283 1342 2290
rect 1394 2283 1407 2335
rect 1459 2283 1472 2335
rect 1524 2283 1537 2335
rect 1589 2283 1601 2335
rect 1653 2324 1665 2335
rect 1717 2324 1729 2335
rect 1781 2324 1793 2335
rect 1845 2324 1857 2335
rect 1909 2324 1921 2335
rect 1662 2290 1665 2324
rect 1845 2290 1847 2324
rect 1909 2290 1920 2324
rect 1653 2283 1665 2290
rect 1717 2283 1729 2290
rect 1781 2283 1793 2290
rect 1845 2283 1857 2290
rect 1909 2283 1921 2290
rect 1973 2283 1985 2335
rect 2037 2283 2049 2335
rect 2101 2283 2113 2335
rect 2165 2324 2177 2335
rect 2229 2324 5271 2335
rect 5323 2324 5335 2335
rect 2173 2290 2177 2324
rect 2247 2290 2287 2324
rect 2321 2290 2361 2324
rect 2395 2290 2435 2324
rect 2469 2290 2509 2324
rect 2543 2290 2583 2324
rect 2617 2290 2657 2324
rect 2691 2290 2731 2324
rect 2765 2290 2805 2324
rect 2839 2290 2879 2324
rect 2913 2290 2953 2324
rect 2987 2290 3027 2324
rect 3061 2290 3101 2324
rect 3135 2290 3175 2324
rect 3209 2290 3249 2324
rect 3283 2290 3323 2324
rect 3357 2290 3397 2324
rect 3431 2290 3471 2324
rect 3505 2290 3545 2324
rect 3579 2290 3921 2324
rect 3955 2290 3995 2324
rect 4029 2290 4069 2324
rect 4103 2290 4143 2324
rect 4177 2290 4217 2324
rect 4251 2290 4291 2324
rect 4325 2290 4365 2324
rect 4399 2290 4439 2324
rect 4473 2290 4513 2324
rect 4547 2290 4587 2324
rect 4621 2290 4661 2324
rect 4695 2290 4735 2324
rect 4769 2290 4809 2324
rect 4843 2290 4883 2324
rect 4917 2290 4957 2324
rect 4991 2290 5031 2324
rect 5065 2290 5105 2324
rect 5139 2290 5179 2324
rect 5213 2290 5253 2324
rect 5323 2290 5327 2324
rect 2165 2283 2177 2290
rect 2229 2283 5271 2290
rect 5323 2283 5335 2290
rect 5387 2283 5399 2335
rect 5451 2283 5463 2335
rect 5515 2283 5527 2335
rect 5579 2324 5591 2335
rect 5643 2324 5655 2335
rect 5707 2324 5719 2335
rect 5771 2324 5783 2335
rect 5835 2324 5847 2335
rect 5580 2290 5591 2324
rect 5653 2290 5655 2324
rect 5835 2290 5838 2324
rect 5579 2283 5591 2290
rect 5643 2283 5655 2290
rect 5707 2283 5719 2290
rect 5771 2283 5783 2290
rect 5835 2283 5847 2290
rect 5899 2283 5911 2335
rect 5963 2283 5976 2335
rect 6028 2283 6041 2335
rect 6093 2283 6106 2335
rect 6158 2324 7826 2335
rect 6164 2290 6203 2324
rect 6237 2290 6276 2324
rect 6310 2290 6349 2324
rect 6383 2290 6422 2324
rect 6456 2290 6495 2324
rect 6529 2290 6568 2324
rect 6602 2290 6641 2324
rect 6675 2290 6714 2324
rect 6748 2290 6787 2324
rect 6821 2290 7163 2324
rect 7197 2290 7236 2324
rect 7270 2290 7309 2324
rect 7343 2290 7382 2324
rect 7416 2290 7455 2324
rect 7489 2290 7528 2324
rect 7562 2290 7601 2324
rect 7635 2290 7674 2324
rect 7708 2290 7747 2324
rect 7781 2290 7820 2324
rect 6158 2283 7826 2290
rect 7878 2283 7891 2335
rect 7943 2283 7956 2335
rect 8008 2283 8021 2335
rect 8073 2283 8085 2335
rect 8137 2324 8149 2335
rect 8201 2324 8213 2335
rect 8265 2324 8277 2335
rect 8329 2324 8341 2335
rect 8393 2324 8405 2335
rect 8146 2290 8149 2324
rect 8329 2290 8331 2324
rect 8393 2290 8404 2324
rect 8137 2283 8149 2290
rect 8201 2283 8213 2290
rect 8265 2283 8277 2290
rect 8329 2283 8341 2290
rect 8393 2283 8405 2290
rect 8457 2283 8469 2335
rect 8521 2283 8533 2335
rect 8585 2283 8597 2335
rect 8649 2324 8661 2335
rect 8713 2324 11755 2335
rect 11807 2324 11819 2335
rect 8657 2290 8661 2324
rect 8731 2290 8771 2324
rect 8805 2290 8845 2324
rect 8879 2290 8919 2324
rect 8953 2290 8993 2324
rect 9027 2290 9067 2324
rect 9101 2290 9141 2324
rect 9175 2290 9215 2324
rect 9249 2290 9289 2324
rect 9323 2290 9363 2324
rect 9397 2290 9437 2324
rect 9471 2290 9511 2324
rect 9545 2290 9585 2324
rect 9619 2290 9659 2324
rect 9693 2290 9733 2324
rect 9767 2290 9807 2324
rect 9841 2290 9881 2324
rect 9915 2290 9955 2324
rect 9989 2290 10029 2324
rect 10063 2290 10405 2324
rect 10439 2290 10479 2324
rect 10513 2290 10553 2324
rect 10587 2290 10627 2324
rect 10661 2290 10701 2324
rect 10735 2290 10775 2324
rect 10809 2290 10849 2324
rect 10883 2290 10923 2324
rect 10957 2290 10997 2324
rect 11031 2290 11071 2324
rect 11105 2290 11145 2324
rect 11179 2290 11219 2324
rect 11253 2290 11293 2324
rect 11327 2290 11367 2324
rect 11401 2290 11441 2324
rect 11475 2290 11515 2324
rect 11549 2290 11589 2324
rect 11623 2290 11663 2324
rect 11697 2290 11737 2324
rect 11807 2290 11811 2324
rect 8649 2283 8661 2290
rect 8713 2283 11755 2290
rect 11807 2283 11819 2290
rect 11871 2283 11883 2335
rect 11935 2283 11947 2335
rect 11999 2283 12011 2335
rect 12063 2324 12075 2335
rect 12127 2324 12139 2335
rect 12191 2324 12203 2335
rect 12255 2324 12267 2335
rect 12319 2324 12331 2335
rect 12064 2290 12075 2324
rect 12137 2290 12139 2324
rect 12319 2290 12322 2324
rect 12063 2283 12075 2290
rect 12127 2283 12139 2290
rect 12191 2283 12203 2290
rect 12255 2283 12267 2290
rect 12319 2283 12331 2290
rect 12383 2283 12395 2335
rect 12447 2283 12460 2335
rect 12512 2283 12525 2335
rect 12577 2283 12590 2335
rect 12642 2324 14310 2335
rect 12648 2290 12687 2324
rect 12721 2290 12760 2324
rect 12794 2290 12833 2324
rect 12867 2290 12906 2324
rect 12940 2290 12979 2324
rect 13013 2290 13052 2324
rect 13086 2290 13125 2324
rect 13159 2290 13198 2324
rect 13232 2290 13271 2324
rect 13305 2290 13647 2324
rect 13681 2290 13720 2324
rect 13754 2290 13793 2324
rect 13827 2290 13866 2324
rect 13900 2290 13939 2324
rect 13973 2290 14012 2324
rect 14046 2290 14085 2324
rect 14119 2290 14158 2324
rect 14192 2290 14231 2324
rect 14265 2290 14304 2324
rect 12642 2283 14310 2290
rect 14362 2283 14375 2335
rect 14427 2283 14440 2335
rect 14492 2283 14505 2335
rect 14557 2283 14569 2335
rect 14621 2324 14633 2335
rect 14685 2324 14697 2335
rect 14749 2324 14761 2335
rect 14813 2324 14825 2335
rect 14877 2324 14889 2335
rect 14630 2290 14633 2324
rect 14813 2290 14815 2324
rect 14877 2290 14888 2324
rect 14621 2283 14633 2290
rect 14685 2283 14697 2290
rect 14749 2283 14761 2290
rect 14813 2283 14825 2290
rect 14877 2283 14889 2290
rect 14941 2283 14953 2335
rect 15005 2283 15017 2335
rect 15069 2283 15081 2335
rect 15133 2324 15145 2335
rect 15197 2324 18239 2335
rect 18291 2324 18303 2335
rect 15141 2290 15145 2324
rect 15215 2290 15255 2324
rect 15289 2290 15329 2324
rect 15363 2290 15403 2324
rect 15437 2290 15477 2324
rect 15511 2290 15551 2324
rect 15585 2290 15625 2324
rect 15659 2290 15699 2324
rect 15733 2290 15773 2324
rect 15807 2290 15847 2324
rect 15881 2290 15921 2324
rect 15955 2290 15995 2324
rect 16029 2290 16069 2324
rect 16103 2290 16143 2324
rect 16177 2290 16217 2324
rect 16251 2290 16291 2324
rect 16325 2290 16365 2324
rect 16399 2290 16439 2324
rect 16473 2290 16513 2324
rect 16547 2290 16889 2324
rect 16923 2290 16963 2324
rect 16997 2290 17037 2324
rect 17071 2290 17111 2324
rect 17145 2290 17185 2324
rect 17219 2290 17259 2324
rect 17293 2290 17333 2324
rect 17367 2290 17407 2324
rect 17441 2290 17481 2324
rect 17515 2290 17555 2324
rect 17589 2290 17629 2324
rect 17663 2290 17703 2324
rect 17737 2290 17777 2324
rect 17811 2290 17851 2324
rect 17885 2290 17925 2324
rect 17959 2290 17999 2324
rect 18033 2290 18073 2324
rect 18107 2290 18147 2324
rect 18181 2290 18221 2324
rect 18291 2290 18295 2324
rect 15133 2283 15145 2290
rect 15197 2283 18239 2290
rect 18291 2283 18303 2290
rect 18355 2283 18367 2335
rect 18419 2283 18431 2335
rect 18483 2283 18495 2335
rect 18547 2324 18559 2335
rect 18611 2324 18623 2335
rect 18675 2324 18687 2335
rect 18739 2324 18751 2335
rect 18803 2324 18815 2335
rect 18548 2290 18559 2324
rect 18621 2290 18623 2324
rect 18803 2290 18806 2324
rect 18547 2283 18559 2290
rect 18611 2283 18623 2290
rect 18675 2283 18687 2290
rect 18739 2283 18751 2290
rect 18803 2283 18815 2290
rect 18867 2283 18879 2335
rect 18931 2283 18944 2335
rect 18996 2283 19009 2335
rect 19061 2283 19074 2335
rect 19126 2324 19889 2335
rect 19132 2290 19171 2324
rect 19205 2290 19244 2324
rect 19278 2290 19317 2324
rect 19351 2290 19390 2324
rect 19424 2290 19463 2324
rect 19497 2290 19536 2324
rect 19570 2290 19609 2324
rect 19643 2290 19682 2324
rect 19716 2290 19755 2324
rect 19789 2290 19889 2324
rect 19126 2283 19889 2290
rect 579 2267 19889 2283
rect 579 2215 1342 2267
rect 1394 2215 1407 2267
rect 1459 2215 1472 2267
rect 1524 2215 1537 2267
rect 1589 2215 1601 2267
rect 1653 2215 1665 2267
rect 1717 2215 1729 2267
rect 1781 2215 1793 2267
rect 1845 2215 1857 2267
rect 1909 2215 1921 2267
rect 1973 2215 1985 2267
rect 2037 2215 2049 2267
rect 2101 2215 2113 2267
rect 2165 2215 2177 2267
rect 2229 2215 5271 2267
rect 5323 2215 5335 2267
rect 5387 2215 5399 2267
rect 5451 2215 5463 2267
rect 5515 2215 5527 2267
rect 5579 2215 5591 2267
rect 5643 2215 5655 2267
rect 5707 2215 5719 2267
rect 5771 2215 5783 2267
rect 5835 2215 5847 2267
rect 5899 2215 5911 2267
rect 5963 2215 5976 2267
rect 6028 2215 6041 2267
rect 6093 2215 6106 2267
rect 6158 2215 7826 2267
rect 7878 2215 7891 2267
rect 7943 2215 7956 2267
rect 8008 2215 8021 2267
rect 8073 2215 8085 2267
rect 8137 2215 8149 2267
rect 8201 2215 8213 2267
rect 8265 2215 8277 2267
rect 8329 2215 8341 2267
rect 8393 2215 8405 2267
rect 8457 2215 8469 2267
rect 8521 2215 8533 2267
rect 8585 2215 8597 2267
rect 8649 2215 8661 2267
rect 8713 2215 11755 2267
rect 11807 2215 11819 2267
rect 11871 2215 11883 2267
rect 11935 2215 11947 2267
rect 11999 2215 12011 2267
rect 12063 2215 12075 2267
rect 12127 2215 12139 2267
rect 12191 2215 12203 2267
rect 12255 2215 12267 2267
rect 12319 2215 12331 2267
rect 12383 2215 12395 2267
rect 12447 2215 12460 2267
rect 12512 2215 12525 2267
rect 12577 2215 12590 2267
rect 12642 2215 14310 2267
rect 14362 2215 14375 2267
rect 14427 2215 14440 2267
rect 14492 2215 14505 2267
rect 14557 2215 14569 2267
rect 14621 2215 14633 2267
rect 14685 2215 14697 2267
rect 14749 2215 14761 2267
rect 14813 2215 14825 2267
rect 14877 2215 14889 2267
rect 14941 2215 14953 2267
rect 15005 2215 15017 2267
rect 15069 2215 15081 2267
rect 15133 2215 15145 2267
rect 15197 2215 18239 2267
rect 18291 2215 18303 2267
rect 18355 2215 18367 2267
rect 18419 2215 18431 2267
rect 18483 2215 18495 2267
rect 18547 2215 18559 2267
rect 18611 2215 18623 2267
rect 18675 2215 18687 2267
rect 18739 2215 18751 2267
rect 18803 2215 18815 2267
rect 18867 2215 18879 2267
rect 18931 2215 18944 2267
rect 18996 2215 19009 2267
rect 19061 2215 19074 2267
rect 19126 2215 19889 2267
rect 579 2199 19889 2215
rect 579 2190 1342 2199
tri 579 2157 612 2190 ne
rect 612 2157 1342 2190
tri 612 2150 619 2157 ne
rect 619 2150 1342 2157
tri 532 2143 539 2150 sw
tri 619 2143 626 2150 ne
rect 626 2147 1342 2150
rect 1394 2147 1407 2199
rect 1459 2147 1472 2199
rect 1524 2147 1537 2199
rect 1589 2147 1601 2199
rect 1653 2147 1665 2199
rect 1717 2147 1729 2199
rect 1781 2147 1793 2199
rect 1845 2147 1857 2199
rect 1909 2147 1921 2199
rect 1973 2147 1985 2199
rect 2037 2147 2049 2199
rect 2101 2147 2113 2199
rect 2165 2147 2177 2199
rect 2229 2190 5271 2199
rect 2229 2157 3618 2190
tri 3618 2157 3651 2190 nw
tri 3852 2157 3885 2190 ne
rect 3885 2157 5271 2190
rect 2229 2147 3604 2157
rect 626 2143 3604 2147
tri 3604 2143 3618 2157 nw
tri 3885 2143 3899 2157 ne
rect 3899 2147 5271 2157
rect 5323 2147 5335 2199
rect 5387 2147 5399 2199
rect 5451 2147 5463 2199
rect 5515 2147 5527 2199
rect 5579 2147 5591 2199
rect 5643 2147 5655 2199
rect 5707 2147 5719 2199
rect 5771 2147 5783 2199
rect 5835 2147 5847 2199
rect 5899 2147 5911 2199
rect 5963 2147 5976 2199
rect 6028 2147 6041 2199
rect 6093 2147 6106 2199
rect 6158 2190 7826 2199
rect 6158 2157 6856 2190
tri 6856 2157 6889 2190 nw
tri 7091 2157 7124 2190 ne
rect 7124 2157 7826 2190
rect 6158 2147 6842 2157
rect 3899 2143 6842 2147
tri 6842 2143 6856 2157 nw
tri 7124 2143 7138 2157 ne
rect 7138 2147 7826 2157
rect 7878 2147 7891 2199
rect 7943 2147 7956 2199
rect 8008 2147 8021 2199
rect 8073 2147 8085 2199
rect 8137 2147 8149 2199
rect 8201 2147 8213 2199
rect 8265 2147 8277 2199
rect 8329 2147 8341 2199
rect 8393 2147 8405 2199
rect 8457 2147 8469 2199
rect 8521 2147 8533 2199
rect 8585 2147 8597 2199
rect 8649 2147 8661 2199
rect 8713 2190 11755 2199
rect 8713 2157 10089 2190
tri 10089 2157 10122 2190 nw
tri 10323 2157 10356 2190 ne
rect 10356 2157 11755 2190
rect 8713 2147 10075 2157
rect 7138 2143 10075 2147
tri 10075 2143 10089 2157 nw
tri 10356 2143 10370 2157 ne
rect 10370 2147 11755 2157
rect 11807 2147 11819 2199
rect 11871 2147 11883 2199
rect 11935 2147 11947 2199
rect 11999 2147 12011 2199
rect 12063 2147 12075 2199
rect 12127 2147 12139 2199
rect 12191 2147 12203 2199
rect 12255 2147 12267 2199
rect 12319 2147 12331 2199
rect 12383 2147 12395 2199
rect 12447 2147 12460 2199
rect 12512 2147 12525 2199
rect 12577 2147 12590 2199
rect 12642 2190 14310 2199
rect 12642 2157 13343 2190
tri 13343 2157 13376 2190 nw
tri 13577 2157 13610 2190 ne
rect 13610 2157 14310 2190
rect 12642 2147 13329 2157
rect 10370 2143 13329 2147
tri 13329 2143 13343 2157 nw
tri 13610 2143 13624 2157 ne
rect 13624 2147 14310 2157
rect 14362 2147 14375 2199
rect 14427 2147 14440 2199
rect 14492 2147 14505 2199
rect 14557 2147 14569 2199
rect 14621 2147 14633 2199
rect 14685 2147 14697 2199
rect 14749 2147 14761 2199
rect 14813 2147 14825 2199
rect 14877 2147 14889 2199
rect 14941 2147 14953 2199
rect 15005 2147 15017 2199
rect 15069 2147 15081 2199
rect 15133 2147 15145 2199
rect 15197 2190 18239 2199
rect 15197 2157 16580 2190
tri 16580 2157 16613 2190 nw
tri 16813 2157 16846 2190 ne
rect 16846 2157 18239 2190
rect 15197 2147 16566 2157
rect 13624 2143 16566 2147
tri 16566 2143 16580 2157 nw
tri 16846 2143 16860 2157 ne
rect 16860 2147 18239 2157
rect 18291 2147 18303 2199
rect 18355 2147 18367 2199
rect 18419 2147 18431 2199
rect 18483 2147 18495 2199
rect 18547 2147 18559 2199
rect 18611 2147 18623 2199
rect 18675 2147 18687 2199
rect 18739 2147 18751 2199
rect 18803 2147 18815 2199
rect 18867 2147 18879 2199
rect 18931 2147 18944 2199
rect 18996 2147 19009 2199
rect 19061 2147 19074 2199
rect 19126 2190 19889 2199
rect 19126 2157 19856 2190
tri 19856 2157 19889 2190 nw
rect 19925 2195 19977 2491
rect 19126 2147 19842 2157
rect 16860 2143 19842 2147
tri 19842 2143 19856 2157 nw
rect 511 2136 539 2143
rect 459 2124 539 2136
rect 511 2119 539 2124
tri 539 2119 563 2143 sw
rect 19925 2131 19977 2143
rect 511 2112 563 2119
tri 563 2112 570 2119 sw
rect 511 2106 16697 2112
rect 517 2072 555 2106
rect 589 2072 3701 2106
rect 3735 2072 3773 2106
rect 3807 2072 6943 2106
rect 6977 2072 7015 2106
rect 7049 2072 10185 2106
rect 10219 2072 10257 2106
rect 10291 2072 13451 2106
rect 13485 2072 13523 2106
rect 13557 2072 16697 2106
rect 19925 2073 19977 2079
rect 459 2066 16697 2072
tri 579 1984 626 2031 se
rect 626 2021 3632 2031
rect 626 1984 959 2021
rect 579 1950 679 1984
rect 713 1950 752 1984
rect 786 1950 825 1984
rect 859 1950 898 1984
rect 932 1969 959 1984
rect 1011 1969 1043 2021
rect 1095 1984 1127 2021
rect 1179 1984 1210 2021
rect 1262 1984 3632 2021
tri 3632 1984 3679 2031 sw
tri 3821 1984 3868 2031 se
rect 3868 2021 6874 2031
tri 6874 2021 6884 2031 sw
tri 7100 2021 7110 2031 se
rect 7110 2021 10116 2031
tri 10116 2021 10126 2031 sw
tri 10342 2021 10352 2031 se
rect 10352 2021 13358 2031
tri 13358 2021 13368 2031 sw
tri 13584 2021 13594 2031 se
rect 13594 2021 16600 2031
rect 3868 1984 6333 2021
rect 1095 1969 1117 1984
rect 1179 1969 1190 1984
rect 1262 1969 1263 1984
rect 932 1957 971 1969
rect 1005 1957 1044 1969
rect 1078 1957 1117 1969
rect 1151 1957 1190 1969
rect 1224 1957 1263 1969
rect 932 1950 959 1957
rect 579 1912 959 1950
rect 579 1878 679 1912
rect 713 1878 752 1912
rect 786 1878 825 1912
rect 859 1878 898 1912
rect 932 1905 959 1912
rect 1011 1905 1043 1957
rect 1095 1950 1117 1957
rect 1179 1950 1190 1957
rect 1262 1950 1263 1957
rect 1297 1950 1336 1984
rect 1370 1950 1409 1984
rect 1443 1950 1482 1984
rect 1516 1950 1555 1984
rect 1589 1950 1628 1984
rect 1662 1950 1701 1984
rect 1735 1950 1774 1984
rect 1808 1950 1847 1984
rect 1881 1950 1920 1984
rect 1954 1950 1993 1984
rect 2027 1950 2066 1984
rect 2100 1950 2139 1984
rect 2173 1950 2213 1984
rect 2247 1950 2287 1984
rect 2321 1950 2361 1984
rect 2395 1950 2435 1984
rect 2469 1950 2509 1984
rect 2543 1950 2583 1984
rect 2617 1950 2657 1984
rect 2691 1950 2731 1984
rect 2765 1950 2805 1984
rect 2839 1950 2879 1984
rect 2913 1950 2953 1984
rect 2987 1950 3027 1984
rect 3061 1950 3101 1984
rect 3135 1950 3175 1984
rect 3209 1950 3249 1984
rect 3283 1950 3323 1984
rect 3357 1950 3397 1984
rect 3431 1950 3471 1984
rect 3505 1950 3545 1984
rect 3579 1950 3921 1984
rect 3955 1950 3995 1984
rect 4029 1950 4069 1984
rect 4103 1950 4143 1984
rect 4177 1950 4217 1984
rect 4251 1950 4291 1984
rect 4325 1950 4365 1984
rect 4399 1950 4439 1984
rect 4473 1950 4513 1984
rect 4547 1950 4587 1984
rect 4621 1950 4661 1984
rect 4695 1950 4735 1984
rect 4769 1950 4809 1984
rect 4843 1950 4883 1984
rect 4917 1950 4957 1984
rect 4991 1950 5031 1984
rect 5065 1950 5105 1984
rect 5139 1950 5179 1984
rect 5213 1950 5253 1984
rect 5287 1950 5327 1984
rect 5361 1950 5400 1984
rect 5434 1950 5473 1984
rect 5507 1950 5546 1984
rect 5580 1950 5619 1984
rect 5653 1950 5692 1984
rect 5726 1950 5765 1984
rect 5799 1950 5838 1984
rect 5872 1950 5911 1984
rect 5945 1950 5984 1984
rect 6018 1950 6057 1984
rect 6091 1950 6130 1984
rect 6164 1950 6203 1984
rect 6237 1950 6276 1984
rect 6310 1969 6333 1984
rect 6385 1969 6400 2021
rect 6452 1984 6467 2021
rect 6519 1984 6534 2021
rect 6586 1984 6601 2021
rect 6653 1984 6668 2021
rect 6720 1984 6884 2021
tri 6884 1984 6921 2021 sw
tri 7063 1984 7100 2021 se
rect 7100 1984 7264 2021
rect 7316 1984 7331 2021
rect 7383 1984 7398 2021
rect 7450 1984 7465 2021
rect 7517 1984 7532 2021
rect 6456 1969 6467 1984
rect 6529 1969 6534 1984
rect 6310 1957 6349 1969
rect 6383 1957 6422 1969
rect 6456 1957 6495 1969
rect 6529 1957 6568 1969
rect 6602 1957 6641 1969
rect 6675 1957 6714 1969
rect 6310 1950 6333 1957
rect 1095 1912 1127 1950
rect 1179 1912 1210 1950
rect 1262 1912 6333 1950
rect 1095 1905 1117 1912
rect 1179 1905 1190 1912
rect 1262 1905 1263 1912
rect 932 1893 971 1905
rect 1005 1893 1044 1905
rect 1078 1893 1117 1905
rect 1151 1893 1190 1905
rect 1224 1893 1263 1905
rect 932 1878 959 1893
tri 579 1831 626 1878 ne
rect 626 1841 959 1878
rect 1011 1841 1043 1893
rect 1095 1878 1117 1893
rect 1179 1878 1190 1893
rect 1262 1878 1263 1893
rect 1297 1878 1336 1912
rect 1370 1878 1409 1912
rect 1443 1878 1482 1912
rect 1516 1878 1555 1912
rect 1589 1878 1628 1912
rect 1662 1878 1701 1912
rect 1735 1878 1774 1912
rect 1808 1878 1847 1912
rect 1881 1878 1920 1912
rect 1954 1878 1993 1912
rect 2027 1878 2066 1912
rect 2100 1878 2139 1912
rect 2173 1878 2213 1912
rect 2247 1878 2287 1912
rect 2321 1878 2361 1912
rect 2395 1878 2435 1912
rect 2469 1878 2509 1912
rect 2543 1878 2583 1912
rect 2617 1878 2657 1912
rect 2691 1878 2731 1912
rect 2765 1878 2805 1912
rect 2839 1878 2879 1912
rect 2913 1878 2953 1912
rect 2987 1878 3027 1912
rect 3061 1878 3101 1912
rect 3135 1878 3175 1912
rect 3209 1878 3249 1912
rect 3283 1878 3323 1912
rect 3357 1878 3397 1912
rect 3431 1878 3471 1912
rect 3505 1878 3545 1912
rect 3579 1878 3921 1912
rect 3955 1878 3995 1912
rect 4029 1878 4069 1912
rect 4103 1878 4143 1912
rect 4177 1878 4217 1912
rect 4251 1878 4291 1912
rect 4325 1878 4365 1912
rect 4399 1878 4439 1912
rect 4473 1878 4513 1912
rect 4547 1878 4587 1912
rect 4621 1878 4661 1912
rect 4695 1878 4735 1912
rect 4769 1878 4809 1912
rect 4843 1878 4883 1912
rect 4917 1878 4957 1912
rect 4991 1878 5031 1912
rect 5065 1878 5105 1912
rect 5139 1878 5179 1912
rect 5213 1878 5253 1912
rect 5287 1878 5327 1912
rect 5361 1878 5400 1912
rect 5434 1878 5473 1912
rect 5507 1878 5546 1912
rect 5580 1878 5619 1912
rect 5653 1878 5692 1912
rect 5726 1878 5765 1912
rect 5799 1878 5838 1912
rect 5872 1878 5911 1912
rect 5945 1878 5984 1912
rect 6018 1878 6057 1912
rect 6091 1878 6130 1912
rect 6164 1878 6203 1912
rect 6237 1878 6276 1912
rect 6310 1905 6333 1912
rect 6385 1905 6400 1957
rect 6456 1950 6467 1957
rect 6529 1950 6534 1957
rect 6748 1950 6787 1984
rect 6821 1950 7163 1984
rect 7197 1950 7236 1984
rect 7450 1969 7455 1984
rect 7517 1969 7528 1984
rect 7584 1969 7599 2021
rect 7651 1984 10126 2021
tri 10126 1984 10163 2021 sw
tri 10305 1984 10342 2021 se
rect 10342 1984 12817 2021
rect 7651 1969 7674 1984
rect 7270 1957 7309 1969
rect 7343 1957 7382 1969
rect 7416 1957 7455 1969
rect 7489 1957 7528 1969
rect 7562 1957 7601 1969
rect 7635 1957 7674 1969
rect 7450 1950 7455 1957
rect 7517 1950 7528 1957
rect 6452 1912 6467 1950
rect 6519 1912 6534 1950
rect 6586 1912 6601 1950
rect 6653 1912 6668 1950
rect 6720 1912 7264 1950
rect 7316 1912 7331 1950
rect 7383 1912 7398 1950
rect 7450 1912 7465 1950
rect 7517 1912 7532 1950
rect 6456 1905 6467 1912
rect 6529 1905 6534 1912
rect 6310 1893 6349 1905
rect 6383 1893 6422 1905
rect 6456 1893 6495 1905
rect 6529 1893 6568 1905
rect 6602 1893 6641 1905
rect 6675 1893 6714 1905
rect 6310 1878 6333 1893
rect 1095 1841 1127 1878
rect 1179 1841 1210 1878
rect 1262 1841 3632 1878
rect 626 1831 3632 1841
tri 3632 1831 3679 1878 nw
tri 3821 1831 3868 1878 ne
rect 3868 1841 6333 1878
rect 6385 1841 6400 1893
rect 6456 1878 6467 1893
rect 6529 1878 6534 1893
rect 6748 1878 6787 1912
rect 6821 1878 7163 1912
rect 7197 1878 7236 1912
rect 7450 1905 7455 1912
rect 7517 1905 7528 1912
rect 7584 1905 7599 1957
rect 7651 1950 7674 1957
rect 7708 1950 7747 1984
rect 7781 1950 7820 1984
rect 7854 1950 7893 1984
rect 7927 1950 7966 1984
rect 8000 1950 8039 1984
rect 8073 1950 8112 1984
rect 8146 1950 8185 1984
rect 8219 1950 8258 1984
rect 8292 1950 8331 1984
rect 8365 1950 8404 1984
rect 8438 1950 8477 1984
rect 8511 1950 8550 1984
rect 8584 1950 8623 1984
rect 8657 1950 8697 1984
rect 8731 1950 8771 1984
rect 8805 1950 8845 1984
rect 8879 1950 8919 1984
rect 8953 1950 8993 1984
rect 9027 1950 9067 1984
rect 9101 1950 9141 1984
rect 9175 1950 9215 1984
rect 9249 1950 9289 1984
rect 9323 1950 9363 1984
rect 9397 1950 9437 1984
rect 9471 1950 9511 1984
rect 9545 1950 9585 1984
rect 9619 1950 9659 1984
rect 9693 1950 9733 1984
rect 9767 1950 9807 1984
rect 9841 1950 9881 1984
rect 9915 1950 9955 1984
rect 9989 1950 10029 1984
rect 10063 1950 10405 1984
rect 10439 1950 10479 1984
rect 10513 1950 10553 1984
rect 10587 1950 10627 1984
rect 10661 1950 10701 1984
rect 10735 1950 10775 1984
rect 10809 1950 10849 1984
rect 10883 1950 10923 1984
rect 10957 1950 10997 1984
rect 11031 1950 11071 1984
rect 11105 1950 11145 1984
rect 11179 1950 11219 1984
rect 11253 1950 11293 1984
rect 11327 1950 11367 1984
rect 11401 1950 11441 1984
rect 11475 1950 11515 1984
rect 11549 1950 11589 1984
rect 11623 1950 11663 1984
rect 11697 1950 11737 1984
rect 11771 1950 11811 1984
rect 11845 1950 11884 1984
rect 11918 1950 11957 1984
rect 11991 1950 12030 1984
rect 12064 1950 12103 1984
rect 12137 1950 12176 1984
rect 12210 1950 12249 1984
rect 12283 1950 12322 1984
rect 12356 1950 12395 1984
rect 12429 1950 12468 1984
rect 12502 1950 12541 1984
rect 12575 1950 12614 1984
rect 12648 1950 12687 1984
rect 12721 1950 12760 1984
rect 12794 1969 12817 1984
rect 12869 1969 12884 2021
rect 12936 1984 12951 2021
rect 13003 1984 13018 2021
rect 13070 1984 13085 2021
rect 13137 1984 13152 2021
rect 13204 1984 13368 2021
tri 13368 1984 13405 2021 sw
tri 13547 1984 13584 2021 se
rect 13584 1984 13748 2021
rect 13800 1984 13815 2021
rect 13867 1984 13882 2021
rect 13934 1984 13949 2021
rect 14001 1984 14016 2021
rect 12940 1969 12951 1984
rect 13013 1969 13018 1984
rect 12794 1957 12833 1969
rect 12867 1957 12906 1969
rect 12940 1957 12979 1969
rect 13013 1957 13052 1969
rect 13086 1957 13125 1969
rect 13159 1957 13198 1969
rect 12794 1950 12817 1957
rect 7651 1912 12817 1950
rect 7651 1905 7674 1912
rect 7270 1893 7309 1905
rect 7343 1893 7382 1905
rect 7416 1893 7455 1905
rect 7489 1893 7528 1905
rect 7562 1893 7601 1905
rect 7635 1893 7674 1905
rect 7450 1878 7455 1893
rect 7517 1878 7528 1893
rect 6452 1841 6467 1878
rect 6519 1841 6534 1878
rect 6586 1841 6601 1878
rect 6653 1841 6668 1878
rect 6720 1841 6884 1878
tri 6884 1841 6921 1878 nw
tri 7063 1841 7100 1878 ne
rect 7100 1841 7264 1878
rect 7316 1841 7331 1878
rect 7383 1841 7398 1878
rect 7450 1841 7465 1878
rect 7517 1841 7532 1878
rect 7584 1841 7599 1893
rect 7651 1878 7674 1893
rect 7708 1878 7747 1912
rect 7781 1878 7820 1912
rect 7854 1878 7893 1912
rect 7927 1878 7966 1912
rect 8000 1878 8039 1912
rect 8073 1878 8112 1912
rect 8146 1878 8185 1912
rect 8219 1878 8258 1912
rect 8292 1878 8331 1912
rect 8365 1878 8404 1912
rect 8438 1878 8477 1912
rect 8511 1878 8550 1912
rect 8584 1878 8623 1912
rect 8657 1878 8697 1912
rect 8731 1878 8771 1912
rect 8805 1878 8845 1912
rect 8879 1878 8919 1912
rect 8953 1878 8993 1912
rect 9027 1878 9067 1912
rect 9101 1878 9141 1912
rect 9175 1878 9215 1912
rect 9249 1878 9289 1912
rect 9323 1878 9363 1912
rect 9397 1878 9437 1912
rect 9471 1878 9511 1912
rect 9545 1878 9585 1912
rect 9619 1878 9659 1912
rect 9693 1878 9733 1912
rect 9767 1878 9807 1912
rect 9841 1878 9881 1912
rect 9915 1878 9955 1912
rect 9989 1878 10029 1912
rect 10063 1878 10405 1912
rect 10439 1878 10479 1912
rect 10513 1878 10553 1912
rect 10587 1878 10627 1912
rect 10661 1878 10701 1912
rect 10735 1878 10775 1912
rect 10809 1878 10849 1912
rect 10883 1878 10923 1912
rect 10957 1878 10997 1912
rect 11031 1878 11071 1912
rect 11105 1878 11145 1912
rect 11179 1878 11219 1912
rect 11253 1878 11293 1912
rect 11327 1878 11367 1912
rect 11401 1878 11441 1912
rect 11475 1878 11515 1912
rect 11549 1878 11589 1912
rect 11623 1878 11663 1912
rect 11697 1878 11737 1912
rect 11771 1878 11811 1912
rect 11845 1878 11884 1912
rect 11918 1878 11957 1912
rect 11991 1878 12030 1912
rect 12064 1878 12103 1912
rect 12137 1878 12176 1912
rect 12210 1878 12249 1912
rect 12283 1878 12322 1912
rect 12356 1878 12395 1912
rect 12429 1878 12468 1912
rect 12502 1878 12541 1912
rect 12575 1878 12614 1912
rect 12648 1878 12687 1912
rect 12721 1878 12760 1912
rect 12794 1905 12817 1912
rect 12869 1905 12884 1957
rect 12940 1950 12951 1957
rect 13013 1950 13018 1957
rect 13232 1950 13271 1984
rect 13305 1950 13647 1984
rect 13681 1950 13720 1984
rect 13934 1969 13939 1984
rect 14001 1969 14012 1984
rect 14068 1969 14083 2021
rect 14135 1984 16600 2021
tri 16600 1984 16647 2031 sw
tri 16826 2021 16836 2031 se
rect 16836 2021 19842 2031
tri 19842 2021 19852 2031 sw
tri 16789 1984 16826 2021 se
rect 16826 1984 19386 2021
rect 19438 1984 19469 2021
rect 19521 1984 19552 2021
rect 19604 1984 19636 2021
rect 19688 1984 19852 2021
tri 19852 1984 19889 2021 sw
rect 14135 1969 14158 1984
rect 13754 1957 13793 1969
rect 13827 1957 13866 1969
rect 13900 1957 13939 1969
rect 13973 1957 14012 1969
rect 14046 1957 14085 1969
rect 14119 1957 14158 1969
rect 13934 1950 13939 1957
rect 14001 1950 14012 1957
rect 12936 1912 12951 1950
rect 13003 1912 13018 1950
rect 13070 1912 13085 1950
rect 13137 1912 13152 1950
rect 13204 1912 13748 1950
rect 13800 1912 13815 1950
rect 13867 1912 13882 1950
rect 13934 1912 13949 1950
rect 14001 1912 14016 1950
rect 12940 1905 12951 1912
rect 13013 1905 13018 1912
rect 12794 1893 12833 1905
rect 12867 1893 12906 1905
rect 12940 1893 12979 1905
rect 13013 1893 13052 1905
rect 13086 1893 13125 1905
rect 13159 1893 13198 1905
rect 12794 1878 12817 1893
rect 7651 1841 10126 1878
tri 10126 1841 10163 1878 nw
tri 10305 1841 10342 1878 ne
rect 10342 1841 12817 1878
rect 12869 1841 12884 1893
rect 12940 1878 12951 1893
rect 13013 1878 13018 1893
rect 13232 1878 13271 1912
rect 13305 1878 13647 1912
rect 13681 1878 13720 1912
rect 13934 1905 13939 1912
rect 14001 1905 14012 1912
rect 14068 1905 14083 1957
rect 14135 1950 14158 1957
rect 14192 1950 14231 1984
rect 14265 1950 14304 1984
rect 14338 1950 14377 1984
rect 14411 1950 14450 1984
rect 14484 1950 14523 1984
rect 14557 1950 14596 1984
rect 14630 1950 14669 1984
rect 14703 1950 14742 1984
rect 14776 1950 14815 1984
rect 14849 1950 14888 1984
rect 14922 1950 14961 1984
rect 14995 1950 15034 1984
rect 15068 1950 15107 1984
rect 15141 1950 15181 1984
rect 15215 1950 15255 1984
rect 15289 1950 15329 1984
rect 15363 1950 15403 1984
rect 15437 1950 15477 1984
rect 15511 1950 15551 1984
rect 15585 1950 15625 1984
rect 15659 1950 15699 1984
rect 15733 1950 15773 1984
rect 15807 1950 15847 1984
rect 15881 1950 15921 1984
rect 15955 1950 15995 1984
rect 16029 1950 16069 1984
rect 16103 1950 16143 1984
rect 16177 1950 16217 1984
rect 16251 1950 16291 1984
rect 16325 1950 16365 1984
rect 16399 1950 16439 1984
rect 16473 1950 16513 1984
rect 16547 1950 16889 1984
rect 16923 1950 16963 1984
rect 16997 1950 17037 1984
rect 17071 1950 17111 1984
rect 17145 1950 17185 1984
rect 17219 1950 17259 1984
rect 17293 1950 17333 1984
rect 17367 1950 17407 1984
rect 17441 1950 17481 1984
rect 17515 1950 17555 1984
rect 17589 1950 17629 1984
rect 17663 1950 17703 1984
rect 17737 1950 17777 1984
rect 17811 1950 17851 1984
rect 17885 1950 17925 1984
rect 17959 1950 17999 1984
rect 18033 1950 18073 1984
rect 18107 1950 18147 1984
rect 18181 1950 18221 1984
rect 18255 1950 18295 1984
rect 18329 1950 18368 1984
rect 18402 1950 18441 1984
rect 18475 1950 18514 1984
rect 18548 1950 18587 1984
rect 18621 1950 18660 1984
rect 18694 1950 18733 1984
rect 18767 1950 18806 1984
rect 18840 1950 18879 1984
rect 18913 1950 18952 1984
rect 18986 1950 19025 1984
rect 19059 1950 19098 1984
rect 19132 1950 19171 1984
rect 19205 1950 19244 1984
rect 19278 1950 19317 1984
rect 19351 1969 19386 1984
rect 19438 1969 19463 1984
rect 19521 1969 19536 1984
rect 19604 1969 19609 1984
rect 19351 1957 19390 1969
rect 19424 1957 19463 1969
rect 19497 1957 19536 1969
rect 19570 1957 19609 1969
rect 19643 1957 19682 1969
rect 19351 1950 19386 1957
rect 19438 1950 19463 1957
rect 19521 1950 19536 1957
rect 19604 1950 19609 1957
rect 19716 1950 19755 1984
rect 19789 1950 19889 1984
rect 14135 1912 19386 1950
rect 19438 1912 19469 1950
rect 19521 1912 19552 1950
rect 19604 1912 19636 1950
rect 19688 1912 19889 1950
rect 14135 1905 14158 1912
rect 13754 1893 13793 1905
rect 13827 1893 13866 1905
rect 13900 1893 13939 1905
rect 13973 1893 14012 1905
rect 14046 1893 14085 1905
rect 14119 1893 14158 1905
rect 13934 1878 13939 1893
rect 14001 1878 14012 1893
rect 12936 1841 12951 1878
rect 13003 1841 13018 1878
rect 13070 1841 13085 1878
rect 13137 1841 13152 1878
rect 13204 1841 13368 1878
tri 13368 1841 13405 1878 nw
tri 13547 1841 13584 1878 ne
rect 13584 1841 13748 1878
rect 13800 1841 13815 1878
rect 13867 1841 13882 1878
rect 13934 1841 13949 1878
rect 14001 1841 14016 1878
rect 14068 1841 14083 1893
rect 14135 1878 14158 1893
rect 14192 1878 14231 1912
rect 14265 1878 14304 1912
rect 14338 1878 14377 1912
rect 14411 1878 14450 1912
rect 14484 1878 14523 1912
rect 14557 1878 14596 1912
rect 14630 1878 14669 1912
rect 14703 1878 14742 1912
rect 14776 1878 14815 1912
rect 14849 1878 14888 1912
rect 14922 1878 14961 1912
rect 14995 1878 15034 1912
rect 15068 1878 15107 1912
rect 15141 1878 15181 1912
rect 15215 1878 15255 1912
rect 15289 1878 15329 1912
rect 15363 1878 15403 1912
rect 15437 1878 15477 1912
rect 15511 1878 15551 1912
rect 15585 1878 15625 1912
rect 15659 1878 15699 1912
rect 15733 1878 15773 1912
rect 15807 1878 15847 1912
rect 15881 1878 15921 1912
rect 15955 1878 15995 1912
rect 16029 1878 16069 1912
rect 16103 1878 16143 1912
rect 16177 1878 16217 1912
rect 16251 1878 16291 1912
rect 16325 1878 16365 1912
rect 16399 1878 16439 1912
rect 16473 1878 16513 1912
rect 16547 1878 16889 1912
rect 16923 1878 16963 1912
rect 16997 1878 17037 1912
rect 17071 1878 17111 1912
rect 17145 1878 17185 1912
rect 17219 1878 17259 1912
rect 17293 1878 17333 1912
rect 17367 1878 17407 1912
rect 17441 1878 17481 1912
rect 17515 1878 17555 1912
rect 17589 1878 17629 1912
rect 17663 1878 17703 1912
rect 17737 1878 17777 1912
rect 17811 1878 17851 1912
rect 17885 1878 17925 1912
rect 17959 1878 17999 1912
rect 18033 1878 18073 1912
rect 18107 1878 18147 1912
rect 18181 1878 18221 1912
rect 18255 1878 18295 1912
rect 18329 1878 18368 1912
rect 18402 1878 18441 1912
rect 18475 1878 18514 1912
rect 18548 1878 18587 1912
rect 18621 1878 18660 1912
rect 18694 1878 18733 1912
rect 18767 1878 18806 1912
rect 18840 1878 18879 1912
rect 18913 1878 18952 1912
rect 18986 1878 19025 1912
rect 19059 1878 19098 1912
rect 19132 1878 19171 1912
rect 19205 1878 19244 1912
rect 19278 1878 19317 1912
rect 19351 1905 19386 1912
rect 19438 1905 19463 1912
rect 19521 1905 19536 1912
rect 19604 1905 19609 1912
rect 19351 1893 19390 1905
rect 19424 1893 19463 1905
rect 19497 1893 19536 1905
rect 19570 1893 19609 1905
rect 19643 1893 19682 1905
rect 19351 1878 19386 1893
rect 19438 1878 19463 1893
rect 19521 1878 19536 1893
rect 19604 1878 19609 1893
rect 19716 1878 19755 1912
rect 19789 1878 19889 1912
rect 14135 1841 16600 1878
rect 3868 1831 6874 1841
tri 6874 1831 6884 1841 nw
tri 7100 1831 7110 1841 ne
rect 7110 1831 10116 1841
tri 10116 1831 10126 1841 nw
tri 10342 1831 10352 1841 ne
rect 10352 1831 13358 1841
tri 13358 1831 13368 1841 nw
tri 13584 1831 13594 1841 ne
rect 13594 1831 16600 1841
tri 16600 1831 16647 1878 nw
tri 16789 1841 16826 1878 ne
rect 16826 1841 19386 1878
rect 19438 1841 19469 1878
rect 19521 1841 19552 1878
rect 19604 1841 19636 1878
rect 19688 1841 19852 1878
tri 19852 1841 19889 1878 nw
tri 16826 1831 16836 1841 ne
rect 16836 1831 19842 1841
tri 19842 1831 19852 1841 nw
rect 6327 -179 6333 -127
rect 6385 -179 6400 -127
rect 6452 -179 6467 -127
rect 6519 -179 6534 -127
rect 6586 -179 6601 -127
rect 6653 -179 6668 -127
rect 6720 -179 6726 -127
rect 7258 -179 7264 -127
rect 7316 -179 7331 -127
rect 7383 -179 7398 -127
rect 7450 -179 7465 -127
rect 7517 -179 7532 -127
rect 7584 -179 7599 -127
rect 7651 -179 7657 -127
rect 12811 -178 12817 -126
rect 12869 -178 12884 -126
rect 12936 -178 12951 -126
rect 13003 -178 13018 -126
rect 13070 -178 13085 -126
rect 13137 -178 13152 -126
rect 13204 -178 13210 -126
rect 13742 -179 13748 -127
rect 13800 -179 13815 -127
rect 13867 -179 13882 -127
rect 13934 -179 13949 -127
rect 14001 -179 14016 -127
rect 14068 -179 14083 -127
rect 14135 -179 14141 -127
rect 19380 -179 19386 -127
rect 19438 -179 19470 -127
rect 19522 -179 19553 -127
rect 19605 -179 19636 -127
rect 19688 -179 19694 -127
rect 872 -1595 878 -1543
rect 930 -1595 944 -1543
rect 996 -1595 1010 -1543
rect 1062 -1595 1076 -1543
rect 1128 -1595 1141 -1543
rect 1193 -1595 1206 -1543
rect 1258 -1595 6334 -1543
rect 6386 -1595 6400 -1543
rect 6452 -1595 6466 -1543
rect 6518 -1595 6532 -1543
rect 6584 -1595 6597 -1543
rect 6649 -1595 6662 -1543
rect 6714 -1595 7266 -1543
rect 7318 -1595 7332 -1543
rect 7384 -1595 7398 -1543
rect 7450 -1595 7464 -1543
rect 7516 -1595 7529 -1543
rect 7581 -1595 7594 -1543
rect 7646 -1595 12819 -1543
rect 12871 -1595 12885 -1543
rect 12937 -1595 12951 -1543
rect 13003 -1595 13017 -1543
rect 13069 -1595 13082 -1543
rect 13134 -1595 13147 -1543
rect 13199 -1595 13750 -1543
rect 13802 -1595 13816 -1543
rect 13868 -1595 13882 -1543
rect 13934 -1595 13948 -1543
rect 14000 -1595 14013 -1543
rect 14065 -1595 14078 -1543
rect 14130 -1595 19303 -1543
rect 19355 -1595 19369 -1543
rect 19421 -1595 19435 -1543
rect 19487 -1595 19501 -1543
rect 19553 -1595 19566 -1543
rect 19618 -1595 19631 -1543
rect 19683 -1595 19689 -1543
rect 872 -1607 19689 -1595
rect 872 -1659 878 -1607
rect 930 -1659 944 -1607
rect 996 -1659 1010 -1607
rect 1062 -1659 1076 -1607
rect 1128 -1659 1141 -1607
rect 1193 -1659 1206 -1607
rect 1258 -1659 6334 -1607
rect 6386 -1659 6400 -1607
rect 6452 -1659 6466 -1607
rect 6518 -1659 6532 -1607
rect 6584 -1659 6597 -1607
rect 6649 -1659 6662 -1607
rect 6714 -1659 7266 -1607
rect 7318 -1659 7332 -1607
rect 7384 -1659 7398 -1607
rect 7450 -1659 7464 -1607
rect 7516 -1659 7529 -1607
rect 7581 -1659 7594 -1607
rect 7646 -1659 12819 -1607
rect 12871 -1659 12885 -1607
rect 12937 -1659 12951 -1607
rect 13003 -1659 13017 -1607
rect 13069 -1659 13082 -1607
rect 13134 -1659 13147 -1607
rect 13199 -1659 13750 -1607
rect 13802 -1659 13816 -1607
rect 13868 -1659 13882 -1607
rect 13934 -1659 13948 -1607
rect 14000 -1659 14013 -1607
rect 14065 -1659 14078 -1607
rect 14130 -1659 19303 -1607
rect 19355 -1659 19369 -1607
rect 19421 -1659 19435 -1607
rect 19487 -1659 19501 -1607
rect 19553 -1659 19566 -1607
rect 19618 -1659 19631 -1607
rect 19683 -1659 19689 -1607
rect 872 -1671 19689 -1659
rect 872 -1723 878 -1671
rect 930 -1723 944 -1671
rect 996 -1723 1010 -1671
rect 1062 -1723 1076 -1671
rect 1128 -1723 1141 -1671
rect 1193 -1723 1206 -1671
rect 1258 -1723 6334 -1671
rect 6386 -1723 6400 -1671
rect 6452 -1723 6466 -1671
rect 6518 -1723 6532 -1671
rect 6584 -1723 6597 -1671
rect 6649 -1723 6662 -1671
rect 6714 -1723 7266 -1671
rect 7318 -1723 7332 -1671
rect 7384 -1723 7398 -1671
rect 7450 -1723 7464 -1671
rect 7516 -1723 7529 -1671
rect 7581 -1723 7594 -1671
rect 7646 -1723 12819 -1671
rect 12871 -1723 12885 -1671
rect 12937 -1723 12951 -1671
rect 13003 -1723 13017 -1671
rect 13069 -1723 13082 -1671
rect 13134 -1723 13147 -1671
rect 13199 -1723 13750 -1671
rect 13802 -1723 13816 -1671
rect 13868 -1723 13882 -1671
rect 13934 -1723 13948 -1671
rect 14000 -1723 14013 -1671
rect 14065 -1723 14078 -1671
rect 14130 -1723 19303 -1671
rect 19355 -1723 19369 -1671
rect 19421 -1723 19435 -1671
rect 19487 -1723 19501 -1671
rect 19553 -1723 19566 -1671
rect 19618 -1723 19631 -1671
rect 19683 -1723 19689 -1671
<< via1 >>
rect 1115 4397 1167 4449
rect 6333 4397 6385 4449
rect 6400 4397 6452 4449
rect 6467 4397 6519 4449
rect 6534 4397 6586 4449
rect 6601 4397 6653 4449
rect 6668 4397 6720 4449
rect 7264 4397 7316 4449
rect 7331 4397 7383 4449
rect 7398 4397 7450 4449
rect 7465 4397 7517 4449
rect 7532 4397 7584 4449
rect 7599 4397 7651 4449
rect 12817 4397 12869 4449
rect 12884 4397 12936 4449
rect 12951 4397 13003 4449
rect 13018 4397 13070 4449
rect 13085 4397 13137 4449
rect 13152 4397 13204 4449
rect 13748 4397 13800 4449
rect 13815 4397 13867 4449
rect 13882 4397 13934 4449
rect 13949 4397 14001 4449
rect 14016 4397 14068 4449
rect 14083 4397 14135 4449
rect 19382 4397 19434 4449
rect 19467 4397 19519 4449
rect 19552 4397 19604 4449
rect 19636 4397 19688 4449
rect 1115 4317 1167 4369
rect 6333 4317 6385 4369
rect 6400 4317 6452 4369
rect 6467 4317 6519 4369
rect 6534 4317 6586 4369
rect 6601 4317 6653 4369
rect 6668 4317 6720 4369
rect 7264 4317 7316 4369
rect 7331 4317 7383 4369
rect 7398 4317 7450 4369
rect 7465 4317 7517 4369
rect 7532 4317 7584 4369
rect 7599 4317 7651 4369
rect 12817 4317 12869 4369
rect 12884 4317 12936 4369
rect 12951 4317 13003 4369
rect 13018 4317 13070 4369
rect 13085 4317 13137 4369
rect 13152 4317 13204 4369
rect 13748 4317 13800 4369
rect 13815 4317 13867 4369
rect 13882 4317 13934 4369
rect 13949 4317 14001 4369
rect 14016 4317 14068 4369
rect 14083 4317 14135 4369
rect 19382 4317 19434 4369
rect 19467 4317 19519 4369
rect 19552 4317 19604 4369
rect 19636 4317 19688 4369
rect 6333 3009 6385 3061
rect 6400 3009 6452 3061
rect 6467 3009 6519 3061
rect 6534 3009 6586 3061
rect 6601 3009 6653 3061
rect 6668 3009 6720 3061
rect 6333 2929 6385 2981
rect 6400 2929 6452 2981
rect 6467 2929 6519 2981
rect 6534 2929 6586 2981
rect 6601 2929 6653 2981
rect 6668 2929 6720 2981
rect 7264 3009 7316 3061
rect 7331 3009 7383 3061
rect 7398 3009 7450 3061
rect 7465 3009 7517 3061
rect 7532 3009 7584 3061
rect 7599 3009 7651 3061
rect 7264 2929 7316 2981
rect 7331 2929 7383 2981
rect 7398 2929 7450 2981
rect 7465 2929 7517 2981
rect 7532 2929 7584 2981
rect 7599 2929 7651 2981
rect 12817 3009 12869 3061
rect 12884 3009 12936 3061
rect 12951 3009 13003 3061
rect 13018 3009 13070 3061
rect 13085 3009 13137 3061
rect 13152 3009 13204 3061
rect 12817 2929 12869 2981
rect 12884 2929 12936 2981
rect 12951 2929 13003 2981
rect 13018 2929 13070 2981
rect 13085 2929 13137 2981
rect 13152 2929 13204 2981
rect 13748 3009 13800 3061
rect 13815 3009 13867 3061
rect 13882 3009 13934 3061
rect 13949 3009 14001 3061
rect 14016 3009 14068 3061
rect 14083 3009 14135 3061
rect 13748 2929 13800 2981
rect 13815 2929 13867 2981
rect 13882 2929 13934 2981
rect 13949 2929 14001 2981
rect 14016 2929 14068 2981
rect 14083 2929 14135 2981
rect 19386 3009 19438 3061
rect 19470 3009 19522 3061
rect 19553 3009 19605 3061
rect 19636 3009 19688 3061
rect 19386 2929 19438 2981
rect 19470 2929 19522 2981
rect 19553 2929 19605 2981
rect 19636 2929 19688 2981
rect 959 2808 1011 2840
rect 959 2788 971 2808
rect 971 2788 1005 2808
rect 1005 2788 1011 2808
rect 1043 2808 1095 2840
rect 1127 2808 1179 2840
rect 1210 2808 1262 2840
rect 6333 2808 6385 2840
rect 1043 2788 1044 2808
rect 1044 2788 1078 2808
rect 1078 2788 1095 2808
rect 1127 2788 1151 2808
rect 1151 2788 1179 2808
rect 1210 2788 1224 2808
rect 1224 2788 1262 2808
rect 959 2774 971 2776
rect 971 2774 1005 2776
rect 1005 2774 1011 2776
rect 959 2736 1011 2774
rect 959 2724 971 2736
rect 971 2724 1005 2736
rect 1005 2724 1011 2736
rect 1043 2774 1044 2776
rect 1044 2774 1078 2776
rect 1078 2774 1095 2776
rect 1127 2774 1151 2776
rect 1151 2774 1179 2776
rect 1210 2774 1224 2776
rect 1224 2774 1262 2776
rect 6333 2788 6349 2808
rect 6349 2788 6383 2808
rect 6383 2788 6385 2808
rect 6400 2808 6452 2840
rect 6467 2808 6519 2840
rect 6534 2808 6586 2840
rect 6601 2808 6653 2840
rect 6668 2808 6720 2840
rect 7264 2808 7316 2840
rect 7331 2808 7383 2840
rect 7398 2808 7450 2840
rect 7465 2808 7517 2840
rect 7532 2808 7584 2840
rect 6400 2788 6422 2808
rect 6422 2788 6452 2808
rect 6467 2788 6495 2808
rect 6495 2788 6519 2808
rect 6534 2788 6568 2808
rect 6568 2788 6586 2808
rect 6601 2788 6602 2808
rect 6602 2788 6641 2808
rect 6641 2788 6653 2808
rect 6668 2788 6675 2808
rect 6675 2788 6714 2808
rect 6714 2788 6720 2808
rect 6333 2774 6349 2776
rect 6349 2774 6383 2776
rect 6383 2774 6385 2776
rect 1043 2736 1095 2774
rect 1127 2736 1179 2774
rect 1210 2736 1262 2774
rect 6333 2736 6385 2774
rect 1043 2724 1044 2736
rect 1044 2724 1078 2736
rect 1078 2724 1095 2736
rect 1127 2724 1151 2736
rect 1151 2724 1179 2736
rect 1210 2724 1224 2736
rect 1224 2724 1262 2736
rect 959 2702 971 2712
rect 971 2702 1005 2712
rect 1005 2702 1011 2712
rect 959 2660 1011 2702
rect 1043 2702 1044 2712
rect 1044 2702 1078 2712
rect 1078 2702 1095 2712
rect 1127 2702 1151 2712
rect 1151 2702 1179 2712
rect 1210 2702 1224 2712
rect 1224 2702 1262 2712
rect 6333 2724 6349 2736
rect 6349 2724 6383 2736
rect 6383 2724 6385 2736
rect 6400 2774 6422 2776
rect 6422 2774 6452 2776
rect 6467 2774 6495 2776
rect 6495 2774 6519 2776
rect 6534 2774 6568 2776
rect 6568 2774 6586 2776
rect 6601 2774 6602 2776
rect 6602 2774 6641 2776
rect 6641 2774 6653 2776
rect 6668 2774 6675 2776
rect 6675 2774 6714 2776
rect 6714 2774 6720 2776
rect 7264 2788 7270 2808
rect 7270 2788 7309 2808
rect 7309 2788 7316 2808
rect 7331 2788 7343 2808
rect 7343 2788 7382 2808
rect 7382 2788 7383 2808
rect 7398 2788 7416 2808
rect 7416 2788 7450 2808
rect 7465 2788 7489 2808
rect 7489 2788 7517 2808
rect 7532 2788 7562 2808
rect 7562 2788 7584 2808
rect 7599 2808 7651 2840
rect 12817 2808 12869 2840
rect 7599 2788 7601 2808
rect 7601 2788 7635 2808
rect 7635 2788 7651 2808
rect 7264 2774 7270 2776
rect 7270 2774 7309 2776
rect 7309 2774 7316 2776
rect 7331 2774 7343 2776
rect 7343 2774 7382 2776
rect 7382 2774 7383 2776
rect 7398 2774 7416 2776
rect 7416 2774 7450 2776
rect 7465 2774 7489 2776
rect 7489 2774 7517 2776
rect 7532 2774 7562 2776
rect 7562 2774 7584 2776
rect 6400 2736 6452 2774
rect 6467 2736 6519 2774
rect 6534 2736 6586 2774
rect 6601 2736 6653 2774
rect 6668 2736 6720 2774
rect 7264 2736 7316 2774
rect 7331 2736 7383 2774
rect 7398 2736 7450 2774
rect 7465 2736 7517 2774
rect 7532 2736 7584 2774
rect 6400 2724 6422 2736
rect 6422 2724 6452 2736
rect 6467 2724 6495 2736
rect 6495 2724 6519 2736
rect 6534 2724 6568 2736
rect 6568 2724 6586 2736
rect 6601 2724 6602 2736
rect 6602 2724 6641 2736
rect 6641 2724 6653 2736
rect 6668 2724 6675 2736
rect 6675 2724 6714 2736
rect 6714 2724 6720 2736
rect 6333 2702 6349 2712
rect 6349 2702 6383 2712
rect 6383 2702 6385 2712
rect 1043 2660 1095 2702
rect 1127 2660 1179 2702
rect 1210 2660 1262 2702
rect 6333 2660 6385 2702
rect 6400 2702 6422 2712
rect 6422 2702 6452 2712
rect 6467 2702 6495 2712
rect 6495 2702 6519 2712
rect 6534 2702 6568 2712
rect 6568 2702 6586 2712
rect 6601 2702 6602 2712
rect 6602 2702 6641 2712
rect 6641 2702 6653 2712
rect 6668 2702 6675 2712
rect 6675 2702 6714 2712
rect 6714 2702 6720 2712
rect 7264 2724 7270 2736
rect 7270 2724 7309 2736
rect 7309 2724 7316 2736
rect 7331 2724 7343 2736
rect 7343 2724 7382 2736
rect 7382 2724 7383 2736
rect 7398 2724 7416 2736
rect 7416 2724 7450 2736
rect 7465 2724 7489 2736
rect 7489 2724 7517 2736
rect 7532 2724 7562 2736
rect 7562 2724 7584 2736
rect 7599 2774 7601 2776
rect 7601 2774 7635 2776
rect 7635 2774 7651 2776
rect 12817 2788 12833 2808
rect 12833 2788 12867 2808
rect 12867 2788 12869 2808
rect 12884 2808 12936 2840
rect 12951 2808 13003 2840
rect 13018 2808 13070 2840
rect 13085 2808 13137 2840
rect 13152 2808 13204 2840
rect 13748 2808 13800 2840
rect 13815 2808 13867 2840
rect 13882 2808 13934 2840
rect 13949 2808 14001 2840
rect 14016 2808 14068 2840
rect 12884 2788 12906 2808
rect 12906 2788 12936 2808
rect 12951 2788 12979 2808
rect 12979 2788 13003 2808
rect 13018 2788 13052 2808
rect 13052 2788 13070 2808
rect 13085 2788 13086 2808
rect 13086 2788 13125 2808
rect 13125 2788 13137 2808
rect 13152 2788 13159 2808
rect 13159 2788 13198 2808
rect 13198 2788 13204 2808
rect 12817 2774 12833 2776
rect 12833 2774 12867 2776
rect 12867 2774 12869 2776
rect 7599 2736 7651 2774
rect 12817 2736 12869 2774
rect 7599 2724 7601 2736
rect 7601 2724 7635 2736
rect 7635 2724 7651 2736
rect 7264 2702 7270 2712
rect 7270 2702 7309 2712
rect 7309 2702 7316 2712
rect 7331 2702 7343 2712
rect 7343 2702 7382 2712
rect 7382 2702 7383 2712
rect 7398 2702 7416 2712
rect 7416 2702 7450 2712
rect 7465 2702 7489 2712
rect 7489 2702 7517 2712
rect 7532 2702 7562 2712
rect 7562 2702 7584 2712
rect 6400 2660 6452 2702
rect 6467 2660 6519 2702
rect 6534 2660 6586 2702
rect 6601 2660 6653 2702
rect 6668 2660 6720 2702
rect 7264 2660 7316 2702
rect 7331 2660 7383 2702
rect 7398 2660 7450 2702
rect 7465 2660 7517 2702
rect 7532 2660 7584 2702
rect 7599 2702 7601 2712
rect 7601 2702 7635 2712
rect 7635 2702 7651 2712
rect 12817 2724 12833 2736
rect 12833 2724 12867 2736
rect 12867 2724 12869 2736
rect 12884 2774 12906 2776
rect 12906 2774 12936 2776
rect 12951 2774 12979 2776
rect 12979 2774 13003 2776
rect 13018 2774 13052 2776
rect 13052 2774 13070 2776
rect 13085 2774 13086 2776
rect 13086 2774 13125 2776
rect 13125 2774 13137 2776
rect 13152 2774 13159 2776
rect 13159 2774 13198 2776
rect 13198 2774 13204 2776
rect 13748 2788 13754 2808
rect 13754 2788 13793 2808
rect 13793 2788 13800 2808
rect 13815 2788 13827 2808
rect 13827 2788 13866 2808
rect 13866 2788 13867 2808
rect 13882 2788 13900 2808
rect 13900 2788 13934 2808
rect 13949 2788 13973 2808
rect 13973 2788 14001 2808
rect 14016 2788 14046 2808
rect 14046 2788 14068 2808
rect 14083 2808 14135 2840
rect 19386 2808 19438 2840
rect 19469 2808 19521 2840
rect 19552 2808 19604 2840
rect 19636 2808 19688 2840
rect 14083 2788 14085 2808
rect 14085 2788 14119 2808
rect 14119 2788 14135 2808
rect 13748 2774 13754 2776
rect 13754 2774 13793 2776
rect 13793 2774 13800 2776
rect 13815 2774 13827 2776
rect 13827 2774 13866 2776
rect 13866 2774 13867 2776
rect 13882 2774 13900 2776
rect 13900 2774 13934 2776
rect 13949 2774 13973 2776
rect 13973 2774 14001 2776
rect 14016 2774 14046 2776
rect 14046 2774 14068 2776
rect 12884 2736 12936 2774
rect 12951 2736 13003 2774
rect 13018 2736 13070 2774
rect 13085 2736 13137 2774
rect 13152 2736 13204 2774
rect 13748 2736 13800 2774
rect 13815 2736 13867 2774
rect 13882 2736 13934 2774
rect 13949 2736 14001 2774
rect 14016 2736 14068 2774
rect 12884 2724 12906 2736
rect 12906 2724 12936 2736
rect 12951 2724 12979 2736
rect 12979 2724 13003 2736
rect 13018 2724 13052 2736
rect 13052 2724 13070 2736
rect 13085 2724 13086 2736
rect 13086 2724 13125 2736
rect 13125 2724 13137 2736
rect 13152 2724 13159 2736
rect 13159 2724 13198 2736
rect 13198 2724 13204 2736
rect 12817 2702 12833 2712
rect 12833 2702 12867 2712
rect 12867 2702 12869 2712
rect 7599 2660 7651 2702
rect 12817 2660 12869 2702
rect 12884 2702 12906 2712
rect 12906 2702 12936 2712
rect 12951 2702 12979 2712
rect 12979 2702 13003 2712
rect 13018 2702 13052 2712
rect 13052 2702 13070 2712
rect 13085 2702 13086 2712
rect 13086 2702 13125 2712
rect 13125 2702 13137 2712
rect 13152 2702 13159 2712
rect 13159 2702 13198 2712
rect 13198 2702 13204 2712
rect 13748 2724 13754 2736
rect 13754 2724 13793 2736
rect 13793 2724 13800 2736
rect 13815 2724 13827 2736
rect 13827 2724 13866 2736
rect 13866 2724 13867 2736
rect 13882 2724 13900 2736
rect 13900 2724 13934 2736
rect 13949 2724 13973 2736
rect 13973 2724 14001 2736
rect 14016 2724 14046 2736
rect 14046 2724 14068 2736
rect 14083 2774 14085 2776
rect 14085 2774 14119 2776
rect 14119 2774 14135 2776
rect 19386 2788 19390 2808
rect 19390 2788 19424 2808
rect 19424 2788 19438 2808
rect 19469 2788 19497 2808
rect 19497 2788 19521 2808
rect 19552 2788 19570 2808
rect 19570 2788 19604 2808
rect 19636 2788 19643 2808
rect 19643 2788 19682 2808
rect 19682 2788 19688 2808
rect 19386 2774 19390 2776
rect 19390 2774 19424 2776
rect 19424 2774 19438 2776
rect 19469 2774 19497 2776
rect 19497 2774 19521 2776
rect 19552 2774 19570 2776
rect 19570 2774 19604 2776
rect 19636 2774 19643 2776
rect 19643 2774 19682 2776
rect 19682 2774 19688 2776
rect 14083 2736 14135 2774
rect 19386 2736 19438 2774
rect 19469 2736 19521 2774
rect 19552 2736 19604 2774
rect 19636 2736 19688 2774
rect 14083 2724 14085 2736
rect 14085 2724 14119 2736
rect 14119 2724 14135 2736
rect 13748 2702 13754 2712
rect 13754 2702 13793 2712
rect 13793 2702 13800 2712
rect 13815 2702 13827 2712
rect 13827 2702 13866 2712
rect 13866 2702 13867 2712
rect 13882 2702 13900 2712
rect 13900 2702 13934 2712
rect 13949 2702 13973 2712
rect 13973 2702 14001 2712
rect 14016 2702 14046 2712
rect 14046 2702 14068 2712
rect 12884 2660 12936 2702
rect 12951 2660 13003 2702
rect 13018 2660 13070 2702
rect 13085 2660 13137 2702
rect 13152 2660 13204 2702
rect 13748 2660 13800 2702
rect 13815 2660 13867 2702
rect 13882 2660 13934 2702
rect 13949 2660 14001 2702
rect 14016 2660 14068 2702
rect 14083 2702 14085 2712
rect 14085 2702 14119 2712
rect 14119 2702 14135 2712
rect 19386 2724 19390 2736
rect 19390 2724 19424 2736
rect 19424 2724 19438 2736
rect 19469 2724 19497 2736
rect 19497 2724 19521 2736
rect 19552 2724 19570 2736
rect 19570 2724 19604 2736
rect 19636 2724 19643 2736
rect 19643 2724 19682 2736
rect 19682 2724 19688 2736
rect 19386 2702 19390 2712
rect 19390 2702 19424 2712
rect 19424 2702 19438 2712
rect 19469 2702 19497 2712
rect 19497 2702 19521 2712
rect 19552 2702 19570 2712
rect 19570 2702 19604 2712
rect 19636 2702 19643 2712
rect 19643 2702 19682 2712
rect 19682 2702 19688 2712
rect 14083 2660 14135 2702
rect 19386 2660 19438 2702
rect 19469 2660 19521 2702
rect 19552 2660 19604 2702
rect 19636 2660 19688 2702
rect 19925 2603 19977 2607
rect 19925 2569 19937 2603
rect 19937 2569 19971 2603
rect 19971 2569 19977 2603
rect 19925 2555 19977 2569
rect 0 2136 52 2188
rect 178 2136 230 2188
rect 0 2072 52 2124
rect 178 2072 230 2124
rect 459 2136 511 2188
rect 1342 2487 1394 2539
rect 1407 2487 1459 2539
rect 1472 2487 1524 2539
rect 1537 2487 1589 2539
rect 1601 2487 1653 2539
rect 1665 2487 1717 2539
rect 1729 2487 1781 2539
rect 1793 2487 1845 2539
rect 1857 2487 1909 2539
rect 1921 2487 1973 2539
rect 1985 2487 2037 2539
rect 2049 2487 2101 2539
rect 2113 2487 2165 2539
rect 2177 2487 2229 2539
rect 5271 2487 5323 2539
rect 5335 2487 5387 2539
rect 5399 2487 5451 2539
rect 5463 2487 5515 2539
rect 5527 2487 5579 2539
rect 5591 2487 5643 2539
rect 5655 2487 5707 2539
rect 5719 2487 5771 2539
rect 5783 2487 5835 2539
rect 5847 2487 5899 2539
rect 5911 2487 5963 2539
rect 5976 2487 6028 2539
rect 6041 2487 6093 2539
rect 6106 2487 6158 2539
rect 7826 2487 7878 2539
rect 7891 2487 7943 2539
rect 7956 2487 8008 2539
rect 8021 2487 8073 2539
rect 8085 2487 8137 2539
rect 8149 2487 8201 2539
rect 8213 2487 8265 2539
rect 8277 2487 8329 2539
rect 8341 2487 8393 2539
rect 8405 2487 8457 2539
rect 8469 2487 8521 2539
rect 8533 2487 8585 2539
rect 8597 2487 8649 2539
rect 8661 2487 8713 2539
rect 11755 2487 11807 2539
rect 11819 2487 11871 2539
rect 11883 2487 11935 2539
rect 11947 2487 11999 2539
rect 12011 2487 12063 2539
rect 12075 2487 12127 2539
rect 12139 2487 12191 2539
rect 12203 2487 12255 2539
rect 12267 2487 12319 2539
rect 12331 2487 12383 2539
rect 12395 2487 12447 2539
rect 12460 2487 12512 2539
rect 12525 2487 12577 2539
rect 12590 2487 12642 2539
rect 14310 2487 14362 2539
rect 14375 2487 14427 2539
rect 14440 2487 14492 2539
rect 14505 2487 14557 2539
rect 14569 2487 14621 2539
rect 14633 2487 14685 2539
rect 14697 2487 14749 2539
rect 14761 2487 14813 2539
rect 14825 2487 14877 2539
rect 14889 2487 14941 2539
rect 14953 2487 15005 2539
rect 15017 2487 15069 2539
rect 15081 2487 15133 2539
rect 15145 2487 15197 2539
rect 18239 2487 18291 2539
rect 18303 2487 18355 2539
rect 18367 2487 18419 2539
rect 18431 2487 18483 2539
rect 18495 2487 18547 2539
rect 18559 2487 18611 2539
rect 18623 2487 18675 2539
rect 18687 2487 18739 2539
rect 18751 2487 18803 2539
rect 18815 2487 18867 2539
rect 18879 2487 18931 2539
rect 18944 2487 18996 2539
rect 19009 2487 19061 2539
rect 19074 2487 19126 2539
rect 19925 2531 19977 2543
rect 19925 2497 19937 2531
rect 19937 2497 19971 2531
rect 19971 2497 19977 2531
rect 1342 2419 1394 2471
rect 1407 2419 1459 2471
rect 1472 2419 1524 2471
rect 1537 2419 1589 2471
rect 1601 2419 1653 2471
rect 1665 2419 1717 2471
rect 1729 2419 1781 2471
rect 1793 2419 1845 2471
rect 1857 2419 1909 2471
rect 1921 2419 1973 2471
rect 1985 2419 2037 2471
rect 2049 2419 2101 2471
rect 2113 2419 2165 2471
rect 2177 2419 2229 2471
rect 5271 2419 5323 2471
rect 5335 2419 5387 2471
rect 5399 2419 5451 2471
rect 5463 2419 5515 2471
rect 5527 2419 5579 2471
rect 5591 2419 5643 2471
rect 5655 2419 5707 2471
rect 5719 2419 5771 2471
rect 5783 2419 5835 2471
rect 5847 2419 5899 2471
rect 5911 2419 5963 2471
rect 5976 2419 6028 2471
rect 6041 2419 6093 2471
rect 6106 2419 6158 2471
rect 7826 2419 7878 2471
rect 7891 2419 7943 2471
rect 7956 2419 8008 2471
rect 8021 2419 8073 2471
rect 8085 2419 8137 2471
rect 8149 2419 8201 2471
rect 8213 2419 8265 2471
rect 8277 2419 8329 2471
rect 8341 2419 8393 2471
rect 8405 2419 8457 2471
rect 8469 2419 8521 2471
rect 8533 2419 8585 2471
rect 8597 2419 8649 2471
rect 8661 2419 8713 2471
rect 11755 2419 11807 2471
rect 11819 2419 11871 2471
rect 11883 2419 11935 2471
rect 11947 2419 11999 2471
rect 12011 2419 12063 2471
rect 12075 2419 12127 2471
rect 12139 2419 12191 2471
rect 12203 2419 12255 2471
rect 12267 2419 12319 2471
rect 12331 2419 12383 2471
rect 12395 2419 12447 2471
rect 12460 2419 12512 2471
rect 12525 2419 12577 2471
rect 12590 2419 12642 2471
rect 14310 2419 14362 2471
rect 14375 2419 14427 2471
rect 14440 2419 14492 2471
rect 14505 2419 14557 2471
rect 14569 2419 14621 2471
rect 14633 2419 14685 2471
rect 14697 2419 14749 2471
rect 14761 2419 14813 2471
rect 14825 2419 14877 2471
rect 14889 2419 14941 2471
rect 14953 2419 15005 2471
rect 15017 2419 15069 2471
rect 15081 2419 15133 2471
rect 15145 2419 15197 2471
rect 18239 2419 18291 2471
rect 18303 2419 18355 2471
rect 18367 2419 18419 2471
rect 18431 2419 18483 2471
rect 18495 2419 18547 2471
rect 18559 2419 18611 2471
rect 18623 2419 18675 2471
rect 18687 2419 18739 2471
rect 18751 2419 18803 2471
rect 18815 2419 18867 2471
rect 18879 2419 18931 2471
rect 18944 2419 18996 2471
rect 19009 2419 19061 2471
rect 19074 2419 19126 2471
rect 1342 2396 1394 2403
rect 1342 2362 1370 2396
rect 1370 2362 1394 2396
rect 1342 2351 1394 2362
rect 1407 2396 1459 2403
rect 1407 2362 1409 2396
rect 1409 2362 1443 2396
rect 1443 2362 1459 2396
rect 1407 2351 1459 2362
rect 1472 2396 1524 2403
rect 1472 2362 1482 2396
rect 1482 2362 1516 2396
rect 1516 2362 1524 2396
rect 1472 2351 1524 2362
rect 1537 2396 1589 2403
rect 1537 2362 1555 2396
rect 1555 2362 1589 2396
rect 1537 2351 1589 2362
rect 1601 2396 1653 2403
rect 1665 2396 1717 2403
rect 1729 2396 1781 2403
rect 1793 2396 1845 2403
rect 1857 2396 1909 2403
rect 1921 2396 1973 2403
rect 1601 2362 1628 2396
rect 1628 2362 1653 2396
rect 1665 2362 1701 2396
rect 1701 2362 1717 2396
rect 1729 2362 1735 2396
rect 1735 2362 1774 2396
rect 1774 2362 1781 2396
rect 1793 2362 1808 2396
rect 1808 2362 1845 2396
rect 1857 2362 1881 2396
rect 1881 2362 1909 2396
rect 1921 2362 1954 2396
rect 1954 2362 1973 2396
rect 1601 2351 1653 2362
rect 1665 2351 1717 2362
rect 1729 2351 1781 2362
rect 1793 2351 1845 2362
rect 1857 2351 1909 2362
rect 1921 2351 1973 2362
rect 1985 2396 2037 2403
rect 1985 2362 1993 2396
rect 1993 2362 2027 2396
rect 2027 2362 2037 2396
rect 1985 2351 2037 2362
rect 2049 2396 2101 2403
rect 2049 2362 2066 2396
rect 2066 2362 2100 2396
rect 2100 2362 2101 2396
rect 2049 2351 2101 2362
rect 2113 2396 2165 2403
rect 2177 2396 2229 2403
rect 5271 2396 5323 2403
rect 5335 2396 5387 2403
rect 2113 2362 2139 2396
rect 2139 2362 2165 2396
rect 2177 2362 2213 2396
rect 2213 2362 2229 2396
rect 5271 2362 5287 2396
rect 5287 2362 5323 2396
rect 5335 2362 5361 2396
rect 5361 2362 5387 2396
rect 2113 2351 2165 2362
rect 2177 2351 2229 2362
rect 5271 2351 5323 2362
rect 5335 2351 5387 2362
rect 5399 2396 5451 2403
rect 5399 2362 5400 2396
rect 5400 2362 5434 2396
rect 5434 2362 5451 2396
rect 5399 2351 5451 2362
rect 5463 2396 5515 2403
rect 5463 2362 5473 2396
rect 5473 2362 5507 2396
rect 5507 2362 5515 2396
rect 5463 2351 5515 2362
rect 5527 2396 5579 2403
rect 5591 2396 5643 2403
rect 5655 2396 5707 2403
rect 5719 2396 5771 2403
rect 5783 2396 5835 2403
rect 5847 2396 5899 2403
rect 5527 2362 5546 2396
rect 5546 2362 5579 2396
rect 5591 2362 5619 2396
rect 5619 2362 5643 2396
rect 5655 2362 5692 2396
rect 5692 2362 5707 2396
rect 5719 2362 5726 2396
rect 5726 2362 5765 2396
rect 5765 2362 5771 2396
rect 5783 2362 5799 2396
rect 5799 2362 5835 2396
rect 5847 2362 5872 2396
rect 5872 2362 5899 2396
rect 5527 2351 5579 2362
rect 5591 2351 5643 2362
rect 5655 2351 5707 2362
rect 5719 2351 5771 2362
rect 5783 2351 5835 2362
rect 5847 2351 5899 2362
rect 5911 2396 5963 2403
rect 5911 2362 5945 2396
rect 5945 2362 5963 2396
rect 5911 2351 5963 2362
rect 5976 2396 6028 2403
rect 5976 2362 5984 2396
rect 5984 2362 6018 2396
rect 6018 2362 6028 2396
rect 5976 2351 6028 2362
rect 6041 2396 6093 2403
rect 6041 2362 6057 2396
rect 6057 2362 6091 2396
rect 6091 2362 6093 2396
rect 6041 2351 6093 2362
rect 6106 2396 6158 2403
rect 7826 2396 7878 2403
rect 6106 2362 6130 2396
rect 6130 2362 6158 2396
rect 7826 2362 7854 2396
rect 7854 2362 7878 2396
rect 6106 2351 6158 2362
rect 7826 2351 7878 2362
rect 7891 2396 7943 2403
rect 7891 2362 7893 2396
rect 7893 2362 7927 2396
rect 7927 2362 7943 2396
rect 7891 2351 7943 2362
rect 7956 2396 8008 2403
rect 7956 2362 7966 2396
rect 7966 2362 8000 2396
rect 8000 2362 8008 2396
rect 7956 2351 8008 2362
rect 8021 2396 8073 2403
rect 8021 2362 8039 2396
rect 8039 2362 8073 2396
rect 8021 2351 8073 2362
rect 8085 2396 8137 2403
rect 8149 2396 8201 2403
rect 8213 2396 8265 2403
rect 8277 2396 8329 2403
rect 8341 2396 8393 2403
rect 8405 2396 8457 2403
rect 8085 2362 8112 2396
rect 8112 2362 8137 2396
rect 8149 2362 8185 2396
rect 8185 2362 8201 2396
rect 8213 2362 8219 2396
rect 8219 2362 8258 2396
rect 8258 2362 8265 2396
rect 8277 2362 8292 2396
rect 8292 2362 8329 2396
rect 8341 2362 8365 2396
rect 8365 2362 8393 2396
rect 8405 2362 8438 2396
rect 8438 2362 8457 2396
rect 8085 2351 8137 2362
rect 8149 2351 8201 2362
rect 8213 2351 8265 2362
rect 8277 2351 8329 2362
rect 8341 2351 8393 2362
rect 8405 2351 8457 2362
rect 8469 2396 8521 2403
rect 8469 2362 8477 2396
rect 8477 2362 8511 2396
rect 8511 2362 8521 2396
rect 8469 2351 8521 2362
rect 8533 2396 8585 2403
rect 8533 2362 8550 2396
rect 8550 2362 8584 2396
rect 8584 2362 8585 2396
rect 8533 2351 8585 2362
rect 8597 2396 8649 2403
rect 8661 2396 8713 2403
rect 11755 2396 11807 2403
rect 11819 2396 11871 2403
rect 8597 2362 8623 2396
rect 8623 2362 8649 2396
rect 8661 2362 8697 2396
rect 8697 2362 8713 2396
rect 11755 2362 11771 2396
rect 11771 2362 11807 2396
rect 11819 2362 11845 2396
rect 11845 2362 11871 2396
rect 8597 2351 8649 2362
rect 8661 2351 8713 2362
rect 11755 2351 11807 2362
rect 11819 2351 11871 2362
rect 11883 2396 11935 2403
rect 11883 2362 11884 2396
rect 11884 2362 11918 2396
rect 11918 2362 11935 2396
rect 11883 2351 11935 2362
rect 11947 2396 11999 2403
rect 11947 2362 11957 2396
rect 11957 2362 11991 2396
rect 11991 2362 11999 2396
rect 11947 2351 11999 2362
rect 12011 2396 12063 2403
rect 12075 2396 12127 2403
rect 12139 2396 12191 2403
rect 12203 2396 12255 2403
rect 12267 2396 12319 2403
rect 12331 2396 12383 2403
rect 12011 2362 12030 2396
rect 12030 2362 12063 2396
rect 12075 2362 12103 2396
rect 12103 2362 12127 2396
rect 12139 2362 12176 2396
rect 12176 2362 12191 2396
rect 12203 2362 12210 2396
rect 12210 2362 12249 2396
rect 12249 2362 12255 2396
rect 12267 2362 12283 2396
rect 12283 2362 12319 2396
rect 12331 2362 12356 2396
rect 12356 2362 12383 2396
rect 12011 2351 12063 2362
rect 12075 2351 12127 2362
rect 12139 2351 12191 2362
rect 12203 2351 12255 2362
rect 12267 2351 12319 2362
rect 12331 2351 12383 2362
rect 12395 2396 12447 2403
rect 12395 2362 12429 2396
rect 12429 2362 12447 2396
rect 12395 2351 12447 2362
rect 12460 2396 12512 2403
rect 12460 2362 12468 2396
rect 12468 2362 12502 2396
rect 12502 2362 12512 2396
rect 12460 2351 12512 2362
rect 12525 2396 12577 2403
rect 12525 2362 12541 2396
rect 12541 2362 12575 2396
rect 12575 2362 12577 2396
rect 12525 2351 12577 2362
rect 12590 2396 12642 2403
rect 14310 2396 14362 2403
rect 12590 2362 12614 2396
rect 12614 2362 12642 2396
rect 14310 2362 14338 2396
rect 14338 2362 14362 2396
rect 12590 2351 12642 2362
rect 14310 2351 14362 2362
rect 14375 2396 14427 2403
rect 14375 2362 14377 2396
rect 14377 2362 14411 2396
rect 14411 2362 14427 2396
rect 14375 2351 14427 2362
rect 14440 2396 14492 2403
rect 14440 2362 14450 2396
rect 14450 2362 14484 2396
rect 14484 2362 14492 2396
rect 14440 2351 14492 2362
rect 14505 2396 14557 2403
rect 14505 2362 14523 2396
rect 14523 2362 14557 2396
rect 14505 2351 14557 2362
rect 14569 2396 14621 2403
rect 14633 2396 14685 2403
rect 14697 2396 14749 2403
rect 14761 2396 14813 2403
rect 14825 2396 14877 2403
rect 14889 2396 14941 2403
rect 14569 2362 14596 2396
rect 14596 2362 14621 2396
rect 14633 2362 14669 2396
rect 14669 2362 14685 2396
rect 14697 2362 14703 2396
rect 14703 2362 14742 2396
rect 14742 2362 14749 2396
rect 14761 2362 14776 2396
rect 14776 2362 14813 2396
rect 14825 2362 14849 2396
rect 14849 2362 14877 2396
rect 14889 2362 14922 2396
rect 14922 2362 14941 2396
rect 14569 2351 14621 2362
rect 14633 2351 14685 2362
rect 14697 2351 14749 2362
rect 14761 2351 14813 2362
rect 14825 2351 14877 2362
rect 14889 2351 14941 2362
rect 14953 2396 15005 2403
rect 14953 2362 14961 2396
rect 14961 2362 14995 2396
rect 14995 2362 15005 2396
rect 14953 2351 15005 2362
rect 15017 2396 15069 2403
rect 15017 2362 15034 2396
rect 15034 2362 15068 2396
rect 15068 2362 15069 2396
rect 15017 2351 15069 2362
rect 15081 2396 15133 2403
rect 15145 2396 15197 2403
rect 18239 2396 18291 2403
rect 18303 2396 18355 2403
rect 15081 2362 15107 2396
rect 15107 2362 15133 2396
rect 15145 2362 15181 2396
rect 15181 2362 15197 2396
rect 18239 2362 18255 2396
rect 18255 2362 18291 2396
rect 18303 2362 18329 2396
rect 18329 2362 18355 2396
rect 15081 2351 15133 2362
rect 15145 2351 15197 2362
rect 18239 2351 18291 2362
rect 18303 2351 18355 2362
rect 18367 2396 18419 2403
rect 18367 2362 18368 2396
rect 18368 2362 18402 2396
rect 18402 2362 18419 2396
rect 18367 2351 18419 2362
rect 18431 2396 18483 2403
rect 18431 2362 18441 2396
rect 18441 2362 18475 2396
rect 18475 2362 18483 2396
rect 18431 2351 18483 2362
rect 18495 2396 18547 2403
rect 18559 2396 18611 2403
rect 18623 2396 18675 2403
rect 18687 2396 18739 2403
rect 18751 2396 18803 2403
rect 18815 2396 18867 2403
rect 18495 2362 18514 2396
rect 18514 2362 18547 2396
rect 18559 2362 18587 2396
rect 18587 2362 18611 2396
rect 18623 2362 18660 2396
rect 18660 2362 18675 2396
rect 18687 2362 18694 2396
rect 18694 2362 18733 2396
rect 18733 2362 18739 2396
rect 18751 2362 18767 2396
rect 18767 2362 18803 2396
rect 18815 2362 18840 2396
rect 18840 2362 18867 2396
rect 18495 2351 18547 2362
rect 18559 2351 18611 2362
rect 18623 2351 18675 2362
rect 18687 2351 18739 2362
rect 18751 2351 18803 2362
rect 18815 2351 18867 2362
rect 18879 2396 18931 2403
rect 18879 2362 18913 2396
rect 18913 2362 18931 2396
rect 18879 2351 18931 2362
rect 18944 2396 18996 2403
rect 18944 2362 18952 2396
rect 18952 2362 18986 2396
rect 18986 2362 18996 2396
rect 18944 2351 18996 2362
rect 19009 2396 19061 2403
rect 19009 2362 19025 2396
rect 19025 2362 19059 2396
rect 19059 2362 19061 2396
rect 19009 2351 19061 2362
rect 19074 2396 19126 2403
rect 19074 2362 19098 2396
rect 19098 2362 19126 2396
rect 19074 2351 19126 2362
rect 1342 2324 1394 2335
rect 1342 2290 1370 2324
rect 1370 2290 1394 2324
rect 1342 2283 1394 2290
rect 1407 2324 1459 2335
rect 1407 2290 1409 2324
rect 1409 2290 1443 2324
rect 1443 2290 1459 2324
rect 1407 2283 1459 2290
rect 1472 2324 1524 2335
rect 1472 2290 1482 2324
rect 1482 2290 1516 2324
rect 1516 2290 1524 2324
rect 1472 2283 1524 2290
rect 1537 2324 1589 2335
rect 1537 2290 1555 2324
rect 1555 2290 1589 2324
rect 1537 2283 1589 2290
rect 1601 2324 1653 2335
rect 1665 2324 1717 2335
rect 1729 2324 1781 2335
rect 1793 2324 1845 2335
rect 1857 2324 1909 2335
rect 1921 2324 1973 2335
rect 1601 2290 1628 2324
rect 1628 2290 1653 2324
rect 1665 2290 1701 2324
rect 1701 2290 1717 2324
rect 1729 2290 1735 2324
rect 1735 2290 1774 2324
rect 1774 2290 1781 2324
rect 1793 2290 1808 2324
rect 1808 2290 1845 2324
rect 1857 2290 1881 2324
rect 1881 2290 1909 2324
rect 1921 2290 1954 2324
rect 1954 2290 1973 2324
rect 1601 2283 1653 2290
rect 1665 2283 1717 2290
rect 1729 2283 1781 2290
rect 1793 2283 1845 2290
rect 1857 2283 1909 2290
rect 1921 2283 1973 2290
rect 1985 2324 2037 2335
rect 1985 2290 1993 2324
rect 1993 2290 2027 2324
rect 2027 2290 2037 2324
rect 1985 2283 2037 2290
rect 2049 2324 2101 2335
rect 2049 2290 2066 2324
rect 2066 2290 2100 2324
rect 2100 2290 2101 2324
rect 2049 2283 2101 2290
rect 2113 2324 2165 2335
rect 2177 2324 2229 2335
rect 5271 2324 5323 2335
rect 5335 2324 5387 2335
rect 2113 2290 2139 2324
rect 2139 2290 2165 2324
rect 2177 2290 2213 2324
rect 2213 2290 2229 2324
rect 5271 2290 5287 2324
rect 5287 2290 5323 2324
rect 5335 2290 5361 2324
rect 5361 2290 5387 2324
rect 2113 2283 2165 2290
rect 2177 2283 2229 2290
rect 5271 2283 5323 2290
rect 5335 2283 5387 2290
rect 5399 2324 5451 2335
rect 5399 2290 5400 2324
rect 5400 2290 5434 2324
rect 5434 2290 5451 2324
rect 5399 2283 5451 2290
rect 5463 2324 5515 2335
rect 5463 2290 5473 2324
rect 5473 2290 5507 2324
rect 5507 2290 5515 2324
rect 5463 2283 5515 2290
rect 5527 2324 5579 2335
rect 5591 2324 5643 2335
rect 5655 2324 5707 2335
rect 5719 2324 5771 2335
rect 5783 2324 5835 2335
rect 5847 2324 5899 2335
rect 5527 2290 5546 2324
rect 5546 2290 5579 2324
rect 5591 2290 5619 2324
rect 5619 2290 5643 2324
rect 5655 2290 5692 2324
rect 5692 2290 5707 2324
rect 5719 2290 5726 2324
rect 5726 2290 5765 2324
rect 5765 2290 5771 2324
rect 5783 2290 5799 2324
rect 5799 2290 5835 2324
rect 5847 2290 5872 2324
rect 5872 2290 5899 2324
rect 5527 2283 5579 2290
rect 5591 2283 5643 2290
rect 5655 2283 5707 2290
rect 5719 2283 5771 2290
rect 5783 2283 5835 2290
rect 5847 2283 5899 2290
rect 5911 2324 5963 2335
rect 5911 2290 5945 2324
rect 5945 2290 5963 2324
rect 5911 2283 5963 2290
rect 5976 2324 6028 2335
rect 5976 2290 5984 2324
rect 5984 2290 6018 2324
rect 6018 2290 6028 2324
rect 5976 2283 6028 2290
rect 6041 2324 6093 2335
rect 6041 2290 6057 2324
rect 6057 2290 6091 2324
rect 6091 2290 6093 2324
rect 6041 2283 6093 2290
rect 6106 2324 6158 2335
rect 7826 2324 7878 2335
rect 6106 2290 6130 2324
rect 6130 2290 6158 2324
rect 7826 2290 7854 2324
rect 7854 2290 7878 2324
rect 6106 2283 6158 2290
rect 7826 2283 7878 2290
rect 7891 2324 7943 2335
rect 7891 2290 7893 2324
rect 7893 2290 7927 2324
rect 7927 2290 7943 2324
rect 7891 2283 7943 2290
rect 7956 2324 8008 2335
rect 7956 2290 7966 2324
rect 7966 2290 8000 2324
rect 8000 2290 8008 2324
rect 7956 2283 8008 2290
rect 8021 2324 8073 2335
rect 8021 2290 8039 2324
rect 8039 2290 8073 2324
rect 8021 2283 8073 2290
rect 8085 2324 8137 2335
rect 8149 2324 8201 2335
rect 8213 2324 8265 2335
rect 8277 2324 8329 2335
rect 8341 2324 8393 2335
rect 8405 2324 8457 2335
rect 8085 2290 8112 2324
rect 8112 2290 8137 2324
rect 8149 2290 8185 2324
rect 8185 2290 8201 2324
rect 8213 2290 8219 2324
rect 8219 2290 8258 2324
rect 8258 2290 8265 2324
rect 8277 2290 8292 2324
rect 8292 2290 8329 2324
rect 8341 2290 8365 2324
rect 8365 2290 8393 2324
rect 8405 2290 8438 2324
rect 8438 2290 8457 2324
rect 8085 2283 8137 2290
rect 8149 2283 8201 2290
rect 8213 2283 8265 2290
rect 8277 2283 8329 2290
rect 8341 2283 8393 2290
rect 8405 2283 8457 2290
rect 8469 2324 8521 2335
rect 8469 2290 8477 2324
rect 8477 2290 8511 2324
rect 8511 2290 8521 2324
rect 8469 2283 8521 2290
rect 8533 2324 8585 2335
rect 8533 2290 8550 2324
rect 8550 2290 8584 2324
rect 8584 2290 8585 2324
rect 8533 2283 8585 2290
rect 8597 2324 8649 2335
rect 8661 2324 8713 2335
rect 11755 2324 11807 2335
rect 11819 2324 11871 2335
rect 8597 2290 8623 2324
rect 8623 2290 8649 2324
rect 8661 2290 8697 2324
rect 8697 2290 8713 2324
rect 11755 2290 11771 2324
rect 11771 2290 11807 2324
rect 11819 2290 11845 2324
rect 11845 2290 11871 2324
rect 8597 2283 8649 2290
rect 8661 2283 8713 2290
rect 11755 2283 11807 2290
rect 11819 2283 11871 2290
rect 11883 2324 11935 2335
rect 11883 2290 11884 2324
rect 11884 2290 11918 2324
rect 11918 2290 11935 2324
rect 11883 2283 11935 2290
rect 11947 2324 11999 2335
rect 11947 2290 11957 2324
rect 11957 2290 11991 2324
rect 11991 2290 11999 2324
rect 11947 2283 11999 2290
rect 12011 2324 12063 2335
rect 12075 2324 12127 2335
rect 12139 2324 12191 2335
rect 12203 2324 12255 2335
rect 12267 2324 12319 2335
rect 12331 2324 12383 2335
rect 12011 2290 12030 2324
rect 12030 2290 12063 2324
rect 12075 2290 12103 2324
rect 12103 2290 12127 2324
rect 12139 2290 12176 2324
rect 12176 2290 12191 2324
rect 12203 2290 12210 2324
rect 12210 2290 12249 2324
rect 12249 2290 12255 2324
rect 12267 2290 12283 2324
rect 12283 2290 12319 2324
rect 12331 2290 12356 2324
rect 12356 2290 12383 2324
rect 12011 2283 12063 2290
rect 12075 2283 12127 2290
rect 12139 2283 12191 2290
rect 12203 2283 12255 2290
rect 12267 2283 12319 2290
rect 12331 2283 12383 2290
rect 12395 2324 12447 2335
rect 12395 2290 12429 2324
rect 12429 2290 12447 2324
rect 12395 2283 12447 2290
rect 12460 2324 12512 2335
rect 12460 2290 12468 2324
rect 12468 2290 12502 2324
rect 12502 2290 12512 2324
rect 12460 2283 12512 2290
rect 12525 2324 12577 2335
rect 12525 2290 12541 2324
rect 12541 2290 12575 2324
rect 12575 2290 12577 2324
rect 12525 2283 12577 2290
rect 12590 2324 12642 2335
rect 14310 2324 14362 2335
rect 12590 2290 12614 2324
rect 12614 2290 12642 2324
rect 14310 2290 14338 2324
rect 14338 2290 14362 2324
rect 12590 2283 12642 2290
rect 14310 2283 14362 2290
rect 14375 2324 14427 2335
rect 14375 2290 14377 2324
rect 14377 2290 14411 2324
rect 14411 2290 14427 2324
rect 14375 2283 14427 2290
rect 14440 2324 14492 2335
rect 14440 2290 14450 2324
rect 14450 2290 14484 2324
rect 14484 2290 14492 2324
rect 14440 2283 14492 2290
rect 14505 2324 14557 2335
rect 14505 2290 14523 2324
rect 14523 2290 14557 2324
rect 14505 2283 14557 2290
rect 14569 2324 14621 2335
rect 14633 2324 14685 2335
rect 14697 2324 14749 2335
rect 14761 2324 14813 2335
rect 14825 2324 14877 2335
rect 14889 2324 14941 2335
rect 14569 2290 14596 2324
rect 14596 2290 14621 2324
rect 14633 2290 14669 2324
rect 14669 2290 14685 2324
rect 14697 2290 14703 2324
rect 14703 2290 14742 2324
rect 14742 2290 14749 2324
rect 14761 2290 14776 2324
rect 14776 2290 14813 2324
rect 14825 2290 14849 2324
rect 14849 2290 14877 2324
rect 14889 2290 14922 2324
rect 14922 2290 14941 2324
rect 14569 2283 14621 2290
rect 14633 2283 14685 2290
rect 14697 2283 14749 2290
rect 14761 2283 14813 2290
rect 14825 2283 14877 2290
rect 14889 2283 14941 2290
rect 14953 2324 15005 2335
rect 14953 2290 14961 2324
rect 14961 2290 14995 2324
rect 14995 2290 15005 2324
rect 14953 2283 15005 2290
rect 15017 2324 15069 2335
rect 15017 2290 15034 2324
rect 15034 2290 15068 2324
rect 15068 2290 15069 2324
rect 15017 2283 15069 2290
rect 15081 2324 15133 2335
rect 15145 2324 15197 2335
rect 18239 2324 18291 2335
rect 18303 2324 18355 2335
rect 15081 2290 15107 2324
rect 15107 2290 15133 2324
rect 15145 2290 15181 2324
rect 15181 2290 15197 2324
rect 18239 2290 18255 2324
rect 18255 2290 18291 2324
rect 18303 2290 18329 2324
rect 18329 2290 18355 2324
rect 15081 2283 15133 2290
rect 15145 2283 15197 2290
rect 18239 2283 18291 2290
rect 18303 2283 18355 2290
rect 18367 2324 18419 2335
rect 18367 2290 18368 2324
rect 18368 2290 18402 2324
rect 18402 2290 18419 2324
rect 18367 2283 18419 2290
rect 18431 2324 18483 2335
rect 18431 2290 18441 2324
rect 18441 2290 18475 2324
rect 18475 2290 18483 2324
rect 18431 2283 18483 2290
rect 18495 2324 18547 2335
rect 18559 2324 18611 2335
rect 18623 2324 18675 2335
rect 18687 2324 18739 2335
rect 18751 2324 18803 2335
rect 18815 2324 18867 2335
rect 18495 2290 18514 2324
rect 18514 2290 18547 2324
rect 18559 2290 18587 2324
rect 18587 2290 18611 2324
rect 18623 2290 18660 2324
rect 18660 2290 18675 2324
rect 18687 2290 18694 2324
rect 18694 2290 18733 2324
rect 18733 2290 18739 2324
rect 18751 2290 18767 2324
rect 18767 2290 18803 2324
rect 18815 2290 18840 2324
rect 18840 2290 18867 2324
rect 18495 2283 18547 2290
rect 18559 2283 18611 2290
rect 18623 2283 18675 2290
rect 18687 2283 18739 2290
rect 18751 2283 18803 2290
rect 18815 2283 18867 2290
rect 18879 2324 18931 2335
rect 18879 2290 18913 2324
rect 18913 2290 18931 2324
rect 18879 2283 18931 2290
rect 18944 2324 18996 2335
rect 18944 2290 18952 2324
rect 18952 2290 18986 2324
rect 18986 2290 18996 2324
rect 18944 2283 18996 2290
rect 19009 2324 19061 2335
rect 19009 2290 19025 2324
rect 19025 2290 19059 2324
rect 19059 2290 19061 2324
rect 19009 2283 19061 2290
rect 19074 2324 19126 2335
rect 19074 2290 19098 2324
rect 19098 2290 19126 2324
rect 19074 2283 19126 2290
rect 1342 2215 1394 2267
rect 1407 2215 1459 2267
rect 1472 2215 1524 2267
rect 1537 2215 1589 2267
rect 1601 2215 1653 2267
rect 1665 2215 1717 2267
rect 1729 2215 1781 2267
rect 1793 2215 1845 2267
rect 1857 2215 1909 2267
rect 1921 2215 1973 2267
rect 1985 2215 2037 2267
rect 2049 2215 2101 2267
rect 2113 2215 2165 2267
rect 2177 2215 2229 2267
rect 5271 2215 5323 2267
rect 5335 2215 5387 2267
rect 5399 2215 5451 2267
rect 5463 2215 5515 2267
rect 5527 2215 5579 2267
rect 5591 2215 5643 2267
rect 5655 2215 5707 2267
rect 5719 2215 5771 2267
rect 5783 2215 5835 2267
rect 5847 2215 5899 2267
rect 5911 2215 5963 2267
rect 5976 2215 6028 2267
rect 6041 2215 6093 2267
rect 6106 2215 6158 2267
rect 7826 2215 7878 2267
rect 7891 2215 7943 2267
rect 7956 2215 8008 2267
rect 8021 2215 8073 2267
rect 8085 2215 8137 2267
rect 8149 2215 8201 2267
rect 8213 2215 8265 2267
rect 8277 2215 8329 2267
rect 8341 2215 8393 2267
rect 8405 2215 8457 2267
rect 8469 2215 8521 2267
rect 8533 2215 8585 2267
rect 8597 2215 8649 2267
rect 8661 2215 8713 2267
rect 11755 2215 11807 2267
rect 11819 2215 11871 2267
rect 11883 2215 11935 2267
rect 11947 2215 11999 2267
rect 12011 2215 12063 2267
rect 12075 2215 12127 2267
rect 12139 2215 12191 2267
rect 12203 2215 12255 2267
rect 12267 2215 12319 2267
rect 12331 2215 12383 2267
rect 12395 2215 12447 2267
rect 12460 2215 12512 2267
rect 12525 2215 12577 2267
rect 12590 2215 12642 2267
rect 14310 2215 14362 2267
rect 14375 2215 14427 2267
rect 14440 2215 14492 2267
rect 14505 2215 14557 2267
rect 14569 2215 14621 2267
rect 14633 2215 14685 2267
rect 14697 2215 14749 2267
rect 14761 2215 14813 2267
rect 14825 2215 14877 2267
rect 14889 2215 14941 2267
rect 14953 2215 15005 2267
rect 15017 2215 15069 2267
rect 15081 2215 15133 2267
rect 15145 2215 15197 2267
rect 18239 2215 18291 2267
rect 18303 2215 18355 2267
rect 18367 2215 18419 2267
rect 18431 2215 18483 2267
rect 18495 2215 18547 2267
rect 18559 2215 18611 2267
rect 18623 2215 18675 2267
rect 18687 2215 18739 2267
rect 18751 2215 18803 2267
rect 18815 2215 18867 2267
rect 18879 2215 18931 2267
rect 18944 2215 18996 2267
rect 19009 2215 19061 2267
rect 19074 2215 19126 2267
rect 1342 2147 1394 2199
rect 1407 2147 1459 2199
rect 1472 2147 1524 2199
rect 1537 2147 1589 2199
rect 1601 2147 1653 2199
rect 1665 2147 1717 2199
rect 1729 2147 1781 2199
rect 1793 2147 1845 2199
rect 1857 2147 1909 2199
rect 1921 2147 1973 2199
rect 1985 2147 2037 2199
rect 2049 2147 2101 2199
rect 2113 2147 2165 2199
rect 2177 2147 2229 2199
rect 5271 2147 5323 2199
rect 5335 2147 5387 2199
rect 5399 2147 5451 2199
rect 5463 2147 5515 2199
rect 5527 2147 5579 2199
rect 5591 2147 5643 2199
rect 5655 2147 5707 2199
rect 5719 2147 5771 2199
rect 5783 2147 5835 2199
rect 5847 2147 5899 2199
rect 5911 2147 5963 2199
rect 5976 2147 6028 2199
rect 6041 2147 6093 2199
rect 6106 2147 6158 2199
rect 7826 2147 7878 2199
rect 7891 2147 7943 2199
rect 7956 2147 8008 2199
rect 8021 2147 8073 2199
rect 8085 2147 8137 2199
rect 8149 2147 8201 2199
rect 8213 2147 8265 2199
rect 8277 2147 8329 2199
rect 8341 2147 8393 2199
rect 8405 2147 8457 2199
rect 8469 2147 8521 2199
rect 8533 2147 8585 2199
rect 8597 2147 8649 2199
rect 8661 2147 8713 2199
rect 11755 2147 11807 2199
rect 11819 2147 11871 2199
rect 11883 2147 11935 2199
rect 11947 2147 11999 2199
rect 12011 2147 12063 2199
rect 12075 2147 12127 2199
rect 12139 2147 12191 2199
rect 12203 2147 12255 2199
rect 12267 2147 12319 2199
rect 12331 2147 12383 2199
rect 12395 2147 12447 2199
rect 12460 2147 12512 2199
rect 12525 2147 12577 2199
rect 12590 2147 12642 2199
rect 14310 2147 14362 2199
rect 14375 2147 14427 2199
rect 14440 2147 14492 2199
rect 14505 2147 14557 2199
rect 14569 2147 14621 2199
rect 14633 2147 14685 2199
rect 14697 2147 14749 2199
rect 14761 2147 14813 2199
rect 14825 2147 14877 2199
rect 14889 2147 14941 2199
rect 14953 2147 15005 2199
rect 15017 2147 15069 2199
rect 15081 2147 15133 2199
rect 15145 2147 15197 2199
rect 18239 2147 18291 2199
rect 18303 2147 18355 2199
rect 18367 2147 18419 2199
rect 18431 2147 18483 2199
rect 18495 2147 18547 2199
rect 18559 2147 18611 2199
rect 18623 2147 18675 2199
rect 18687 2147 18739 2199
rect 18751 2147 18803 2199
rect 18815 2147 18867 2199
rect 18879 2147 18931 2199
rect 18944 2147 18996 2199
rect 19009 2147 19061 2199
rect 19074 2147 19126 2199
rect 19925 2491 19977 2497
rect 19925 2191 19977 2195
rect 19925 2157 19937 2191
rect 19937 2157 19971 2191
rect 19971 2157 19977 2191
rect 19925 2143 19977 2157
rect 459 2106 511 2124
rect 19925 2119 19977 2131
rect 459 2072 483 2106
rect 483 2072 511 2106
rect 19925 2085 19937 2119
rect 19937 2085 19971 2119
rect 19971 2085 19977 2119
rect 19925 2079 19977 2085
rect 959 1984 1011 2021
rect 959 1969 971 1984
rect 971 1969 1005 1984
rect 1005 1969 1011 1984
rect 1043 1984 1095 2021
rect 1127 1984 1179 2021
rect 1210 1984 1262 2021
rect 6333 1984 6385 2021
rect 1043 1969 1044 1984
rect 1044 1969 1078 1984
rect 1078 1969 1095 1984
rect 1127 1969 1151 1984
rect 1151 1969 1179 1984
rect 1210 1969 1224 1984
rect 1224 1969 1262 1984
rect 959 1950 971 1957
rect 971 1950 1005 1957
rect 1005 1950 1011 1957
rect 959 1912 1011 1950
rect 959 1905 971 1912
rect 971 1905 1005 1912
rect 1005 1905 1011 1912
rect 1043 1950 1044 1957
rect 1044 1950 1078 1957
rect 1078 1950 1095 1957
rect 1127 1950 1151 1957
rect 1151 1950 1179 1957
rect 1210 1950 1224 1957
rect 1224 1950 1262 1957
rect 6333 1969 6349 1984
rect 6349 1969 6383 1984
rect 6383 1969 6385 1984
rect 6400 1984 6452 2021
rect 6467 1984 6519 2021
rect 6534 1984 6586 2021
rect 6601 1984 6653 2021
rect 6668 1984 6720 2021
rect 7264 1984 7316 2021
rect 7331 1984 7383 2021
rect 7398 1984 7450 2021
rect 7465 1984 7517 2021
rect 7532 1984 7584 2021
rect 6400 1969 6422 1984
rect 6422 1969 6452 1984
rect 6467 1969 6495 1984
rect 6495 1969 6519 1984
rect 6534 1969 6568 1984
rect 6568 1969 6586 1984
rect 6601 1969 6602 1984
rect 6602 1969 6641 1984
rect 6641 1969 6653 1984
rect 6668 1969 6675 1984
rect 6675 1969 6714 1984
rect 6714 1969 6720 1984
rect 6333 1950 6349 1957
rect 6349 1950 6383 1957
rect 6383 1950 6385 1957
rect 1043 1912 1095 1950
rect 1127 1912 1179 1950
rect 1210 1912 1262 1950
rect 6333 1912 6385 1950
rect 1043 1905 1044 1912
rect 1044 1905 1078 1912
rect 1078 1905 1095 1912
rect 1127 1905 1151 1912
rect 1151 1905 1179 1912
rect 1210 1905 1224 1912
rect 1224 1905 1262 1912
rect 959 1878 971 1893
rect 971 1878 1005 1893
rect 1005 1878 1011 1893
rect 959 1841 1011 1878
rect 1043 1878 1044 1893
rect 1044 1878 1078 1893
rect 1078 1878 1095 1893
rect 1127 1878 1151 1893
rect 1151 1878 1179 1893
rect 1210 1878 1224 1893
rect 1224 1878 1262 1893
rect 6333 1905 6349 1912
rect 6349 1905 6383 1912
rect 6383 1905 6385 1912
rect 6400 1950 6422 1957
rect 6422 1950 6452 1957
rect 6467 1950 6495 1957
rect 6495 1950 6519 1957
rect 6534 1950 6568 1957
rect 6568 1950 6586 1957
rect 6601 1950 6602 1957
rect 6602 1950 6641 1957
rect 6641 1950 6653 1957
rect 6668 1950 6675 1957
rect 6675 1950 6714 1957
rect 6714 1950 6720 1957
rect 7264 1969 7270 1984
rect 7270 1969 7309 1984
rect 7309 1969 7316 1984
rect 7331 1969 7343 1984
rect 7343 1969 7382 1984
rect 7382 1969 7383 1984
rect 7398 1969 7416 1984
rect 7416 1969 7450 1984
rect 7465 1969 7489 1984
rect 7489 1969 7517 1984
rect 7532 1969 7562 1984
rect 7562 1969 7584 1984
rect 7599 1984 7651 2021
rect 12817 1984 12869 2021
rect 7599 1969 7601 1984
rect 7601 1969 7635 1984
rect 7635 1969 7651 1984
rect 7264 1950 7270 1957
rect 7270 1950 7309 1957
rect 7309 1950 7316 1957
rect 7331 1950 7343 1957
rect 7343 1950 7382 1957
rect 7382 1950 7383 1957
rect 7398 1950 7416 1957
rect 7416 1950 7450 1957
rect 7465 1950 7489 1957
rect 7489 1950 7517 1957
rect 7532 1950 7562 1957
rect 7562 1950 7584 1957
rect 6400 1912 6452 1950
rect 6467 1912 6519 1950
rect 6534 1912 6586 1950
rect 6601 1912 6653 1950
rect 6668 1912 6720 1950
rect 7264 1912 7316 1950
rect 7331 1912 7383 1950
rect 7398 1912 7450 1950
rect 7465 1912 7517 1950
rect 7532 1912 7584 1950
rect 6400 1905 6422 1912
rect 6422 1905 6452 1912
rect 6467 1905 6495 1912
rect 6495 1905 6519 1912
rect 6534 1905 6568 1912
rect 6568 1905 6586 1912
rect 6601 1905 6602 1912
rect 6602 1905 6641 1912
rect 6641 1905 6653 1912
rect 6668 1905 6675 1912
rect 6675 1905 6714 1912
rect 6714 1905 6720 1912
rect 6333 1878 6349 1893
rect 6349 1878 6383 1893
rect 6383 1878 6385 1893
rect 1043 1841 1095 1878
rect 1127 1841 1179 1878
rect 1210 1841 1262 1878
rect 6333 1841 6385 1878
rect 6400 1878 6422 1893
rect 6422 1878 6452 1893
rect 6467 1878 6495 1893
rect 6495 1878 6519 1893
rect 6534 1878 6568 1893
rect 6568 1878 6586 1893
rect 6601 1878 6602 1893
rect 6602 1878 6641 1893
rect 6641 1878 6653 1893
rect 6668 1878 6675 1893
rect 6675 1878 6714 1893
rect 6714 1878 6720 1893
rect 7264 1905 7270 1912
rect 7270 1905 7309 1912
rect 7309 1905 7316 1912
rect 7331 1905 7343 1912
rect 7343 1905 7382 1912
rect 7382 1905 7383 1912
rect 7398 1905 7416 1912
rect 7416 1905 7450 1912
rect 7465 1905 7489 1912
rect 7489 1905 7517 1912
rect 7532 1905 7562 1912
rect 7562 1905 7584 1912
rect 7599 1950 7601 1957
rect 7601 1950 7635 1957
rect 7635 1950 7651 1957
rect 12817 1969 12833 1984
rect 12833 1969 12867 1984
rect 12867 1969 12869 1984
rect 12884 1984 12936 2021
rect 12951 1984 13003 2021
rect 13018 1984 13070 2021
rect 13085 1984 13137 2021
rect 13152 1984 13204 2021
rect 13748 1984 13800 2021
rect 13815 1984 13867 2021
rect 13882 1984 13934 2021
rect 13949 1984 14001 2021
rect 14016 1984 14068 2021
rect 12884 1969 12906 1984
rect 12906 1969 12936 1984
rect 12951 1969 12979 1984
rect 12979 1969 13003 1984
rect 13018 1969 13052 1984
rect 13052 1969 13070 1984
rect 13085 1969 13086 1984
rect 13086 1969 13125 1984
rect 13125 1969 13137 1984
rect 13152 1969 13159 1984
rect 13159 1969 13198 1984
rect 13198 1969 13204 1984
rect 12817 1950 12833 1957
rect 12833 1950 12867 1957
rect 12867 1950 12869 1957
rect 7599 1912 7651 1950
rect 12817 1912 12869 1950
rect 7599 1905 7601 1912
rect 7601 1905 7635 1912
rect 7635 1905 7651 1912
rect 7264 1878 7270 1893
rect 7270 1878 7309 1893
rect 7309 1878 7316 1893
rect 7331 1878 7343 1893
rect 7343 1878 7382 1893
rect 7382 1878 7383 1893
rect 7398 1878 7416 1893
rect 7416 1878 7450 1893
rect 7465 1878 7489 1893
rect 7489 1878 7517 1893
rect 7532 1878 7562 1893
rect 7562 1878 7584 1893
rect 6400 1841 6452 1878
rect 6467 1841 6519 1878
rect 6534 1841 6586 1878
rect 6601 1841 6653 1878
rect 6668 1841 6720 1878
rect 7264 1841 7316 1878
rect 7331 1841 7383 1878
rect 7398 1841 7450 1878
rect 7465 1841 7517 1878
rect 7532 1841 7584 1878
rect 7599 1878 7601 1893
rect 7601 1878 7635 1893
rect 7635 1878 7651 1893
rect 12817 1905 12833 1912
rect 12833 1905 12867 1912
rect 12867 1905 12869 1912
rect 12884 1950 12906 1957
rect 12906 1950 12936 1957
rect 12951 1950 12979 1957
rect 12979 1950 13003 1957
rect 13018 1950 13052 1957
rect 13052 1950 13070 1957
rect 13085 1950 13086 1957
rect 13086 1950 13125 1957
rect 13125 1950 13137 1957
rect 13152 1950 13159 1957
rect 13159 1950 13198 1957
rect 13198 1950 13204 1957
rect 13748 1969 13754 1984
rect 13754 1969 13793 1984
rect 13793 1969 13800 1984
rect 13815 1969 13827 1984
rect 13827 1969 13866 1984
rect 13866 1969 13867 1984
rect 13882 1969 13900 1984
rect 13900 1969 13934 1984
rect 13949 1969 13973 1984
rect 13973 1969 14001 1984
rect 14016 1969 14046 1984
rect 14046 1969 14068 1984
rect 14083 1984 14135 2021
rect 19386 1984 19438 2021
rect 19469 1984 19521 2021
rect 19552 1984 19604 2021
rect 19636 1984 19688 2021
rect 14083 1969 14085 1984
rect 14085 1969 14119 1984
rect 14119 1969 14135 1984
rect 13748 1950 13754 1957
rect 13754 1950 13793 1957
rect 13793 1950 13800 1957
rect 13815 1950 13827 1957
rect 13827 1950 13866 1957
rect 13866 1950 13867 1957
rect 13882 1950 13900 1957
rect 13900 1950 13934 1957
rect 13949 1950 13973 1957
rect 13973 1950 14001 1957
rect 14016 1950 14046 1957
rect 14046 1950 14068 1957
rect 12884 1912 12936 1950
rect 12951 1912 13003 1950
rect 13018 1912 13070 1950
rect 13085 1912 13137 1950
rect 13152 1912 13204 1950
rect 13748 1912 13800 1950
rect 13815 1912 13867 1950
rect 13882 1912 13934 1950
rect 13949 1912 14001 1950
rect 14016 1912 14068 1950
rect 12884 1905 12906 1912
rect 12906 1905 12936 1912
rect 12951 1905 12979 1912
rect 12979 1905 13003 1912
rect 13018 1905 13052 1912
rect 13052 1905 13070 1912
rect 13085 1905 13086 1912
rect 13086 1905 13125 1912
rect 13125 1905 13137 1912
rect 13152 1905 13159 1912
rect 13159 1905 13198 1912
rect 13198 1905 13204 1912
rect 12817 1878 12833 1893
rect 12833 1878 12867 1893
rect 12867 1878 12869 1893
rect 7599 1841 7651 1878
rect 12817 1841 12869 1878
rect 12884 1878 12906 1893
rect 12906 1878 12936 1893
rect 12951 1878 12979 1893
rect 12979 1878 13003 1893
rect 13018 1878 13052 1893
rect 13052 1878 13070 1893
rect 13085 1878 13086 1893
rect 13086 1878 13125 1893
rect 13125 1878 13137 1893
rect 13152 1878 13159 1893
rect 13159 1878 13198 1893
rect 13198 1878 13204 1893
rect 13748 1905 13754 1912
rect 13754 1905 13793 1912
rect 13793 1905 13800 1912
rect 13815 1905 13827 1912
rect 13827 1905 13866 1912
rect 13866 1905 13867 1912
rect 13882 1905 13900 1912
rect 13900 1905 13934 1912
rect 13949 1905 13973 1912
rect 13973 1905 14001 1912
rect 14016 1905 14046 1912
rect 14046 1905 14068 1912
rect 14083 1950 14085 1957
rect 14085 1950 14119 1957
rect 14119 1950 14135 1957
rect 19386 1969 19390 1984
rect 19390 1969 19424 1984
rect 19424 1969 19438 1984
rect 19469 1969 19497 1984
rect 19497 1969 19521 1984
rect 19552 1969 19570 1984
rect 19570 1969 19604 1984
rect 19636 1969 19643 1984
rect 19643 1969 19682 1984
rect 19682 1969 19688 1984
rect 19386 1950 19390 1957
rect 19390 1950 19424 1957
rect 19424 1950 19438 1957
rect 19469 1950 19497 1957
rect 19497 1950 19521 1957
rect 19552 1950 19570 1957
rect 19570 1950 19604 1957
rect 19636 1950 19643 1957
rect 19643 1950 19682 1957
rect 19682 1950 19688 1957
rect 14083 1912 14135 1950
rect 19386 1912 19438 1950
rect 19469 1912 19521 1950
rect 19552 1912 19604 1950
rect 19636 1912 19688 1950
rect 14083 1905 14085 1912
rect 14085 1905 14119 1912
rect 14119 1905 14135 1912
rect 13748 1878 13754 1893
rect 13754 1878 13793 1893
rect 13793 1878 13800 1893
rect 13815 1878 13827 1893
rect 13827 1878 13866 1893
rect 13866 1878 13867 1893
rect 13882 1878 13900 1893
rect 13900 1878 13934 1893
rect 13949 1878 13973 1893
rect 13973 1878 14001 1893
rect 14016 1878 14046 1893
rect 14046 1878 14068 1893
rect 12884 1841 12936 1878
rect 12951 1841 13003 1878
rect 13018 1841 13070 1878
rect 13085 1841 13137 1878
rect 13152 1841 13204 1878
rect 13748 1841 13800 1878
rect 13815 1841 13867 1878
rect 13882 1841 13934 1878
rect 13949 1841 14001 1878
rect 14016 1841 14068 1878
rect 14083 1878 14085 1893
rect 14085 1878 14119 1893
rect 14119 1878 14135 1893
rect 19386 1905 19390 1912
rect 19390 1905 19424 1912
rect 19424 1905 19438 1912
rect 19469 1905 19497 1912
rect 19497 1905 19521 1912
rect 19552 1905 19570 1912
rect 19570 1905 19604 1912
rect 19636 1905 19643 1912
rect 19643 1905 19682 1912
rect 19682 1905 19688 1912
rect 19386 1878 19390 1893
rect 19390 1878 19424 1893
rect 19424 1878 19438 1893
rect 19469 1878 19497 1893
rect 19497 1878 19521 1893
rect 19552 1878 19570 1893
rect 19570 1878 19604 1893
rect 19636 1878 19643 1893
rect 19643 1878 19682 1893
rect 19682 1878 19688 1893
rect 14083 1841 14135 1878
rect 19386 1841 19438 1878
rect 19469 1841 19521 1878
rect 19552 1841 19604 1878
rect 19636 1841 19688 1878
rect 6333 -179 6385 -127
rect 6400 -179 6452 -127
rect 6467 -179 6519 -127
rect 6534 -179 6586 -127
rect 6601 -179 6653 -127
rect 6668 -179 6720 -127
rect 7264 -179 7316 -127
rect 7331 -179 7383 -127
rect 7398 -179 7450 -127
rect 7465 -179 7517 -127
rect 7532 -179 7584 -127
rect 7599 -179 7651 -127
rect 12817 -178 12869 -126
rect 12884 -178 12936 -126
rect 12951 -178 13003 -126
rect 13018 -178 13070 -126
rect 13085 -178 13137 -126
rect 13152 -178 13204 -126
rect 13748 -179 13800 -127
rect 13815 -179 13867 -127
rect 13882 -179 13934 -127
rect 13949 -179 14001 -127
rect 14016 -179 14068 -127
rect 14083 -179 14135 -127
rect 19386 -179 19438 -127
rect 19470 -179 19522 -127
rect 19553 -179 19605 -127
rect 19636 -179 19688 -127
rect 878 -1595 930 -1543
rect 944 -1595 996 -1543
rect 1010 -1595 1062 -1543
rect 1076 -1595 1128 -1543
rect 1141 -1595 1193 -1543
rect 1206 -1595 1258 -1543
rect 6334 -1595 6386 -1543
rect 6400 -1595 6452 -1543
rect 6466 -1595 6518 -1543
rect 6532 -1595 6584 -1543
rect 6597 -1595 6649 -1543
rect 6662 -1595 6714 -1543
rect 7266 -1595 7318 -1543
rect 7332 -1595 7384 -1543
rect 7398 -1595 7450 -1543
rect 7464 -1595 7516 -1543
rect 7529 -1595 7581 -1543
rect 7594 -1595 7646 -1543
rect 12819 -1595 12871 -1543
rect 12885 -1595 12937 -1543
rect 12951 -1595 13003 -1543
rect 13017 -1595 13069 -1543
rect 13082 -1595 13134 -1543
rect 13147 -1595 13199 -1543
rect 13750 -1595 13802 -1543
rect 13816 -1595 13868 -1543
rect 13882 -1595 13934 -1543
rect 13948 -1595 14000 -1543
rect 14013 -1595 14065 -1543
rect 14078 -1595 14130 -1543
rect 19303 -1595 19355 -1543
rect 19369 -1595 19421 -1543
rect 19435 -1595 19487 -1543
rect 19501 -1595 19553 -1543
rect 19566 -1595 19618 -1543
rect 19631 -1595 19683 -1543
rect 878 -1659 930 -1607
rect 944 -1659 996 -1607
rect 1010 -1659 1062 -1607
rect 1076 -1659 1128 -1607
rect 1141 -1659 1193 -1607
rect 1206 -1659 1258 -1607
rect 6334 -1659 6386 -1607
rect 6400 -1659 6452 -1607
rect 6466 -1659 6518 -1607
rect 6532 -1659 6584 -1607
rect 6597 -1659 6649 -1607
rect 6662 -1659 6714 -1607
rect 7266 -1659 7318 -1607
rect 7332 -1659 7384 -1607
rect 7398 -1659 7450 -1607
rect 7464 -1659 7516 -1607
rect 7529 -1659 7581 -1607
rect 7594 -1659 7646 -1607
rect 12819 -1659 12871 -1607
rect 12885 -1659 12937 -1607
rect 12951 -1659 13003 -1607
rect 13017 -1659 13069 -1607
rect 13082 -1659 13134 -1607
rect 13147 -1659 13199 -1607
rect 13750 -1659 13802 -1607
rect 13816 -1659 13868 -1607
rect 13882 -1659 13934 -1607
rect 13948 -1659 14000 -1607
rect 14013 -1659 14065 -1607
rect 14078 -1659 14130 -1607
rect 19303 -1659 19355 -1607
rect 19369 -1659 19421 -1607
rect 19435 -1659 19487 -1607
rect 19501 -1659 19553 -1607
rect 19566 -1659 19618 -1607
rect 19631 -1659 19683 -1607
rect 878 -1723 930 -1671
rect 944 -1723 996 -1671
rect 1010 -1723 1062 -1671
rect 1076 -1723 1128 -1671
rect 1141 -1723 1193 -1671
rect 1206 -1723 1258 -1671
rect 6334 -1723 6386 -1671
rect 6400 -1723 6452 -1671
rect 6466 -1723 6518 -1671
rect 6532 -1723 6584 -1671
rect 6597 -1723 6649 -1671
rect 6662 -1723 6714 -1671
rect 7266 -1723 7318 -1671
rect 7332 -1723 7384 -1671
rect 7398 -1723 7450 -1671
rect 7464 -1723 7516 -1671
rect 7529 -1723 7581 -1671
rect 7594 -1723 7646 -1671
rect 12819 -1723 12871 -1671
rect 12885 -1723 12937 -1671
rect 12951 -1723 13003 -1671
rect 13017 -1723 13069 -1671
rect 13082 -1723 13134 -1671
rect 13147 -1723 13199 -1671
rect 13750 -1723 13802 -1671
rect 13816 -1723 13868 -1671
rect 13882 -1723 13934 -1671
rect 13948 -1723 14000 -1671
rect 14013 -1723 14065 -1671
rect 14078 -1723 14130 -1671
rect 19303 -1723 19355 -1671
rect 19369 -1723 19421 -1671
rect 19435 -1723 19487 -1671
rect 19501 -1723 19553 -1671
rect 19566 -1723 19618 -1671
rect 19631 -1723 19683 -1671
<< metal2 >>
rect 953 4397 962 4453
rect 1018 4397 1044 4453
rect 1100 4449 1126 4453
rect 1100 4397 1115 4449
rect 1182 4397 1207 4453
rect 1263 4397 1272 4453
rect 953 4369 1272 4397
rect 953 4313 962 4369
rect 1018 4313 1044 4369
rect 1100 4317 1115 4369
rect 1100 4313 1126 4317
rect 1182 4313 1207 4369
rect 1263 4313 1272 4369
rect 6327 4449 6336 4453
rect 6392 4449 6418 4453
rect 6474 4449 6499 4453
rect 6555 4449 6580 4453
rect 6636 4449 6661 4453
rect 6717 4449 6726 4453
rect 6327 4397 6333 4449
rect 6392 4397 6400 4449
rect 6653 4397 6661 4449
rect 6720 4397 6726 4449
rect 6327 4369 6726 4397
rect 6327 4317 6333 4369
rect 6392 4317 6400 4369
rect 6653 4317 6661 4369
rect 6720 4317 6726 4369
rect 6327 4313 6336 4317
rect 6392 4313 6418 4317
rect 6474 4313 6499 4317
rect 6555 4313 6580 4317
rect 6636 4313 6661 4317
rect 6717 4313 6726 4317
rect 7258 4449 7267 4453
rect 7323 4449 7349 4453
rect 7405 4449 7430 4453
rect 7486 4449 7511 4453
rect 7567 4449 7592 4453
rect 7648 4449 7657 4453
rect 7258 4397 7264 4449
rect 7323 4397 7331 4449
rect 7584 4397 7592 4449
rect 7651 4397 7657 4449
rect 7258 4369 7657 4397
rect 7258 4317 7264 4369
rect 7323 4317 7331 4369
rect 7584 4317 7592 4369
rect 7651 4317 7657 4369
rect 7258 4313 7267 4317
rect 7323 4313 7349 4317
rect 7405 4313 7430 4317
rect 7486 4313 7511 4317
rect 7567 4313 7592 4317
rect 7648 4313 7657 4317
rect 12811 4449 12820 4453
rect 12876 4449 12902 4453
rect 12958 4449 12983 4453
rect 13039 4449 13064 4453
rect 13120 4449 13145 4453
rect 13201 4449 13210 4453
rect 12811 4397 12817 4449
rect 12876 4397 12884 4449
rect 13137 4397 13145 4449
rect 13204 4397 13210 4449
rect 12811 4369 13210 4397
rect 12811 4317 12817 4369
rect 12876 4317 12884 4369
rect 13137 4317 13145 4369
rect 13204 4317 13210 4369
rect 12811 4313 12820 4317
rect 12876 4313 12902 4317
rect 12958 4313 12983 4317
rect 13039 4313 13064 4317
rect 13120 4313 13145 4317
rect 13201 4313 13210 4317
rect 13742 4449 13751 4453
rect 13807 4449 13833 4453
rect 13889 4449 13914 4453
rect 13970 4449 13995 4453
rect 14051 4449 14076 4453
rect 14132 4449 14141 4453
rect 13742 4397 13748 4449
rect 13807 4397 13815 4449
rect 14068 4397 14076 4449
rect 14135 4397 14141 4449
rect 13742 4369 14141 4397
rect 13742 4317 13748 4369
rect 13807 4317 13815 4369
rect 14068 4317 14076 4369
rect 14135 4317 14141 4369
rect 13742 4313 13751 4317
rect 13807 4313 13833 4317
rect 13889 4313 13914 4317
rect 13970 4313 13995 4317
rect 14051 4313 14076 4317
rect 14132 4313 14141 4317
rect 19376 4449 19385 4453
rect 19376 4397 19382 4449
rect 19441 4397 19467 4453
rect 19523 4397 19548 4453
rect 19604 4397 19629 4453
rect 19685 4449 19694 4453
rect 19688 4397 19694 4449
rect 19376 4369 19694 4397
rect 19376 4317 19382 4369
rect 19376 4313 19385 4317
rect 19441 4313 19467 4369
rect 19523 4313 19548 4369
rect 19604 4313 19629 4369
rect 19688 4317 19694 4369
rect 19685 4313 19694 4317
rect 953 3009 962 3065
rect 1018 3009 1043 3065
rect 1099 3009 1123 3065
rect 1179 3009 1203 3065
rect 1259 3009 1268 3065
rect 953 2981 1268 3009
rect 953 2925 962 2981
rect 1018 2925 1043 2981
rect 1099 2925 1123 2981
rect 1179 2925 1203 2981
rect 1259 2925 1268 2981
rect 6327 3061 6336 3065
rect 6392 3061 6418 3065
rect 6474 3061 6499 3065
rect 6555 3061 6580 3065
rect 6636 3061 6661 3065
rect 6717 3061 6726 3065
rect 6327 3009 6333 3061
rect 6392 3009 6400 3061
rect 6653 3009 6661 3061
rect 6720 3009 6726 3061
rect 6327 2981 6726 3009
rect 6327 2929 6333 2981
rect 6392 2929 6400 2981
rect 6653 2929 6661 2981
rect 6720 2929 6726 2981
rect 6327 2925 6336 2929
rect 6392 2925 6418 2929
rect 6474 2925 6499 2929
rect 6555 2925 6580 2929
rect 6636 2925 6661 2929
rect 6717 2925 6726 2929
rect 7258 3061 7267 3065
rect 7323 3061 7349 3065
rect 7405 3061 7430 3065
rect 7486 3061 7511 3065
rect 7567 3061 7592 3065
rect 7648 3061 7657 3065
rect 7258 3009 7264 3061
rect 7323 3009 7331 3061
rect 7584 3009 7592 3061
rect 7651 3009 7657 3061
rect 7258 2981 7657 3009
rect 7258 2929 7264 2981
rect 7323 2929 7331 2981
rect 7584 2929 7592 2981
rect 7651 2929 7657 2981
rect 7258 2925 7267 2929
rect 7323 2925 7349 2929
rect 7405 2925 7430 2929
rect 7486 2925 7511 2929
rect 7567 2925 7592 2929
rect 7648 2925 7657 2929
rect 12811 3061 12820 3065
rect 12876 3061 12902 3065
rect 12958 3061 12983 3065
rect 13039 3061 13064 3065
rect 13120 3061 13145 3065
rect 13201 3061 13210 3065
rect 12811 3009 12817 3061
rect 12876 3009 12884 3061
rect 13137 3009 13145 3061
rect 13204 3009 13210 3061
rect 12811 2981 13210 3009
rect 12811 2929 12817 2981
rect 12876 2929 12884 2981
rect 13137 2929 13145 2981
rect 13204 2929 13210 2981
rect 12811 2925 12820 2929
rect 12876 2925 12902 2929
rect 12958 2925 12983 2929
rect 13039 2925 13064 2929
rect 13120 2925 13145 2929
rect 13201 2925 13210 2929
rect 13742 3061 13751 3065
rect 13807 3061 13833 3065
rect 13889 3061 13914 3065
rect 13970 3061 13995 3065
rect 14051 3061 14076 3065
rect 14132 3061 14141 3065
rect 13742 3009 13748 3061
rect 13807 3009 13815 3061
rect 14068 3009 14076 3061
rect 14135 3009 14141 3061
rect 13742 2981 14141 3009
rect 13742 2929 13748 2981
rect 13807 2929 13815 2981
rect 14068 2929 14076 2981
rect 14135 2929 14141 2981
rect 13742 2925 13751 2929
rect 13807 2925 13833 2929
rect 13889 2925 13914 2929
rect 13970 2925 13995 2929
rect 14051 2925 14076 2929
rect 14132 2925 14141 2929
rect 19380 3061 19389 3065
rect 19380 3009 19386 3061
rect 19445 3009 19469 3065
rect 19525 3009 19549 3065
rect 19605 3009 19629 3065
rect 19685 3061 19694 3065
rect 19688 3009 19694 3061
rect 19380 2981 19694 3009
rect 19380 2929 19386 2981
rect 19380 2925 19389 2929
rect 19445 2925 19469 2981
rect 19525 2925 19549 2981
rect 19605 2925 19629 2981
rect 19688 2929 19694 2981
rect 19685 2925 19694 2929
tri 20647 2840 20662 2855 se
rect 20662 2840 20790 3201
rect 953 2788 959 2840
rect 953 2784 962 2788
rect 1018 2784 1043 2840
rect 1099 2784 1123 2840
rect 1179 2784 1203 2840
rect 1262 2788 1268 2840
rect 1259 2784 1268 2788
rect 953 2776 1268 2784
rect 953 2724 959 2776
rect 1011 2724 1043 2776
rect 1095 2724 1127 2776
rect 1179 2724 1210 2776
rect 1262 2724 1268 2776
rect 953 2716 1268 2724
rect 953 2712 962 2716
rect 953 2660 959 2712
rect 1018 2660 1043 2716
rect 1099 2660 1123 2716
rect 1179 2660 1203 2716
rect 1259 2712 1268 2716
rect 1262 2660 1268 2712
rect 6327 2788 6333 2840
rect 6392 2788 6400 2840
rect 6653 2788 6661 2840
rect 6720 2788 6726 2840
rect 6327 2784 6336 2788
rect 6392 2784 6417 2788
rect 6473 2784 6498 2788
rect 6554 2784 6579 2788
rect 6635 2784 6661 2788
rect 6717 2784 6726 2788
rect 6327 2776 6726 2784
rect 6327 2724 6333 2776
rect 6385 2724 6400 2776
rect 6452 2724 6467 2776
rect 6519 2724 6534 2776
rect 6586 2724 6601 2776
rect 6653 2724 6668 2776
rect 6720 2724 6726 2776
rect 6327 2716 6726 2724
rect 6327 2712 6336 2716
rect 6392 2712 6417 2716
rect 6473 2712 6498 2716
rect 6554 2712 6579 2716
rect 6635 2712 6661 2716
rect 6717 2712 6726 2716
rect 6327 2660 6333 2712
rect 6392 2660 6400 2712
rect 6653 2660 6661 2712
rect 6720 2660 6726 2712
rect 7258 2788 7264 2840
rect 7323 2788 7331 2840
rect 7584 2788 7592 2840
rect 7651 2788 7657 2840
rect 7258 2784 7267 2788
rect 7323 2784 7349 2788
rect 7405 2784 7430 2788
rect 7486 2784 7511 2788
rect 7567 2784 7592 2788
rect 7648 2784 7657 2788
rect 7258 2776 7657 2784
rect 7258 2724 7264 2776
rect 7316 2724 7331 2776
rect 7383 2724 7398 2776
rect 7450 2724 7465 2776
rect 7517 2724 7532 2776
rect 7584 2724 7599 2776
rect 7651 2724 7657 2776
rect 7258 2716 7657 2724
rect 7258 2712 7267 2716
rect 7323 2712 7349 2716
rect 7405 2712 7430 2716
rect 7486 2712 7511 2716
rect 7567 2712 7592 2716
rect 7648 2712 7657 2716
rect 7258 2660 7264 2712
rect 7323 2660 7331 2712
rect 7584 2660 7592 2712
rect 7651 2660 7657 2712
rect 12811 2788 12817 2840
rect 12876 2788 12884 2840
rect 13137 2788 13145 2840
rect 13204 2788 13210 2840
rect 12811 2784 12820 2788
rect 12876 2784 12901 2788
rect 12957 2784 12982 2788
rect 13038 2784 13063 2788
rect 13119 2784 13145 2788
rect 13201 2784 13210 2788
rect 12811 2776 13210 2784
rect 12811 2724 12817 2776
rect 12869 2724 12884 2776
rect 12936 2724 12951 2776
rect 13003 2724 13018 2776
rect 13070 2724 13085 2776
rect 13137 2724 13152 2776
rect 13204 2724 13210 2776
rect 12811 2716 13210 2724
rect 12811 2712 12820 2716
rect 12876 2712 12901 2716
rect 12957 2712 12982 2716
rect 13038 2712 13063 2716
rect 13119 2712 13145 2716
rect 13201 2712 13210 2716
rect 12811 2660 12817 2712
rect 12876 2660 12884 2712
rect 13137 2660 13145 2712
rect 13204 2660 13210 2712
rect 13742 2788 13748 2840
rect 13807 2788 13815 2840
rect 14068 2788 14076 2840
rect 14135 2788 14141 2840
rect 13742 2784 13751 2788
rect 13807 2784 13833 2788
rect 13889 2784 13914 2788
rect 13970 2784 13995 2788
rect 14051 2784 14076 2788
rect 14132 2784 14141 2788
rect 13742 2776 14141 2784
rect 13742 2724 13748 2776
rect 13800 2724 13815 2776
rect 13867 2724 13882 2776
rect 13934 2724 13949 2776
rect 14001 2724 14016 2776
rect 14068 2724 14083 2776
rect 14135 2724 14141 2776
rect 13742 2716 14141 2724
rect 13742 2712 13751 2716
rect 13807 2712 13833 2716
rect 13889 2712 13914 2716
rect 13970 2712 13995 2716
rect 14051 2712 14076 2716
rect 14132 2712 14141 2716
rect 13742 2660 13748 2712
rect 13807 2660 13815 2712
rect 14068 2660 14076 2712
rect 14135 2660 14141 2712
rect 19380 2788 19386 2840
rect 19380 2784 19389 2788
rect 19445 2784 19469 2840
rect 19525 2784 19549 2840
rect 19605 2784 19629 2840
rect 19688 2788 19694 2840
tri 20628 2821 20647 2840 se
rect 20647 2821 20790 2840
rect 19685 2784 19694 2788
rect 19380 2776 19694 2784
rect 19380 2724 19386 2776
rect 19438 2724 19469 2776
rect 19521 2724 19552 2776
rect 19604 2724 19636 2776
rect 19688 2724 19694 2776
rect 19925 2783 20501 2821
rect 20563 2783 20790 2821
rect 19925 2781 20003 2783
tri 20003 2781 20005 2783 nw
tri 20628 2781 20630 2783 ne
rect 20630 2781 20790 2783
rect 19925 2729 19977 2781
tri 19977 2755 20003 2781 nw
tri 20630 2755 20656 2781 ne
rect 20656 2755 20790 2781
tri 20656 2749 20662 2755 ne
rect 19926 2727 19976 2728
rect 19380 2716 19694 2724
rect 19380 2712 19389 2716
rect 19380 2660 19386 2712
rect 19445 2660 19469 2716
rect 19525 2660 19549 2716
rect 19605 2660 19629 2716
rect 19685 2712 19694 2716
rect 19688 2660 19694 2712
rect 19380 2655 19694 2660
rect 19380 2640 19679 2655
tri 19679 2640 19694 2655 nw
rect 19926 2666 19976 2667
rect 19925 2640 19977 2665
tri 20656 2642 20662 2648 se
rect 20662 2642 20790 2755
tri 19977 2640 19979 2642 sw
tri 20654 2640 20656 2642 se
rect 20656 2640 20790 2642
rect 19925 2614 19979 2640
tri 19979 2614 20005 2640 sw
tri 20628 2614 20654 2640 se
rect 20654 2614 20790 2640
rect 19925 2607 20790 2614
rect 19977 2576 20790 2607
rect 19925 2543 19977 2555
tri 19977 2549 20004 2576 nw
rect 1336 2539 2235 2543
rect 1336 2487 1342 2539
rect 1589 2487 1599 2539
rect 1655 2487 1665 2539
rect 1909 2487 1921 2539
rect 1982 2487 1985 2539
rect 2165 2487 2169 2539
rect 2229 2487 2235 2539
rect 1336 2483 1353 2487
rect 1409 2483 1435 2487
rect 1491 2483 1517 2487
rect 1573 2483 1599 2487
rect 1655 2483 1681 2487
rect 1737 2483 1763 2487
rect 1819 2483 1845 2487
rect 1901 2483 1926 2487
rect 1982 2483 2007 2487
rect 2063 2483 2088 2487
rect 2144 2483 2169 2487
rect 2225 2483 2235 2487
rect 1336 2471 2235 2483
rect 1336 2419 1342 2471
rect 1394 2455 1407 2471
rect 1459 2455 1472 2471
rect 1524 2455 1537 2471
rect 1589 2455 1601 2471
rect 1653 2455 1665 2471
rect 1717 2455 1729 2471
rect 1781 2455 1793 2471
rect 1845 2455 1857 2471
rect 1589 2419 1599 2455
rect 1655 2419 1665 2455
rect 1909 2419 1921 2471
rect 1973 2455 1985 2471
rect 2037 2455 2049 2471
rect 2101 2455 2113 2471
rect 2165 2455 2177 2471
rect 1982 2419 1985 2455
rect 2165 2419 2169 2455
rect 2229 2419 2235 2471
rect 1336 2403 1353 2419
rect 1409 2403 1435 2419
rect 1491 2403 1517 2419
rect 1573 2403 1599 2419
rect 1655 2403 1681 2419
rect 1737 2403 1763 2419
rect 1819 2403 1845 2419
rect 1901 2403 1926 2419
rect 1982 2403 2007 2419
rect 2063 2403 2088 2419
rect 2144 2403 2169 2419
rect 2225 2403 2235 2419
rect 1336 2351 1342 2403
rect 1589 2399 1599 2403
rect 1655 2399 1665 2403
rect 1394 2371 1407 2399
rect 1459 2371 1472 2399
rect 1524 2371 1537 2399
rect 1589 2371 1601 2399
rect 1653 2371 1665 2399
rect 1717 2371 1729 2399
rect 1781 2371 1793 2399
rect 1845 2371 1857 2399
rect 1589 2351 1599 2371
rect 1655 2351 1665 2371
rect 1909 2351 1921 2403
rect 1982 2399 1985 2403
rect 2165 2399 2169 2403
rect 1973 2371 1985 2399
rect 2037 2371 2049 2399
rect 2101 2371 2113 2399
rect 2165 2371 2177 2399
rect 1982 2351 1985 2371
rect 2165 2351 2169 2371
rect 2229 2351 2235 2403
rect 1336 2335 1353 2351
rect 1409 2335 1435 2351
rect 1491 2335 1517 2351
rect 1573 2335 1599 2351
rect 1655 2335 1681 2351
rect 1737 2335 1763 2351
rect 1819 2335 1845 2351
rect 1901 2335 1926 2351
rect 1982 2335 2007 2351
rect 2063 2335 2088 2351
rect 2144 2335 2169 2351
rect 2225 2335 2235 2351
rect 1336 2283 1342 2335
rect 1589 2315 1599 2335
rect 1655 2315 1665 2335
rect 1394 2287 1407 2315
rect 1459 2287 1472 2315
rect 1524 2287 1537 2315
rect 1589 2287 1601 2315
rect 1653 2287 1665 2315
rect 1717 2287 1729 2315
rect 1781 2287 1793 2315
rect 1845 2287 1857 2315
rect 1589 2283 1599 2287
rect 1655 2283 1665 2287
rect 1909 2283 1921 2335
rect 1982 2315 1985 2335
rect 2165 2315 2169 2335
rect 1973 2287 1985 2315
rect 2037 2287 2049 2315
rect 2101 2287 2113 2315
rect 2165 2287 2177 2315
rect 1982 2283 1985 2287
rect 2165 2283 2169 2287
rect 2229 2283 2235 2335
rect 1336 2267 1353 2283
rect 1409 2267 1435 2283
rect 1491 2267 1517 2283
rect 1573 2267 1599 2283
rect 1655 2267 1681 2283
rect 1737 2267 1763 2283
rect 1819 2267 1845 2283
rect 1901 2267 1926 2283
rect 1982 2267 2007 2283
rect 2063 2267 2088 2283
rect 2144 2267 2169 2283
rect 2225 2267 2235 2283
rect 1336 2215 1342 2267
rect 1589 2231 1599 2267
rect 1655 2231 1665 2267
rect 1394 2215 1407 2231
rect 1459 2215 1472 2231
rect 1524 2215 1537 2231
rect 1589 2215 1601 2231
rect 1653 2215 1665 2231
rect 1717 2215 1729 2231
rect 1781 2215 1793 2231
rect 1845 2215 1857 2231
rect 1909 2215 1921 2267
rect 1982 2231 1985 2267
rect 2165 2231 2169 2267
rect 1973 2215 1985 2231
rect 2037 2215 2049 2231
rect 2101 2215 2113 2231
rect 2165 2215 2177 2231
rect 2229 2215 2235 2267
rect 1336 2203 2235 2215
rect 1336 2199 1353 2203
rect 1409 2199 1435 2203
rect 1491 2199 1517 2203
rect 1573 2199 1599 2203
rect 1655 2199 1681 2203
rect 1737 2199 1763 2203
rect 1819 2199 1845 2203
rect 1901 2199 1926 2203
rect 1982 2199 2007 2203
rect 2063 2199 2088 2203
rect 2144 2199 2169 2203
rect 2225 2199 2235 2203
rect 0 2188 52 2194
rect 0 2124 52 2136
rect 0 2066 52 2072
rect 178 2188 511 2194
rect 230 2136 459 2188
rect 1336 2147 1342 2199
rect 1589 2147 1599 2199
rect 1655 2147 1665 2199
rect 1909 2147 1921 2199
rect 1982 2147 1985 2199
rect 2165 2147 2169 2199
rect 2229 2147 2235 2199
rect 1336 2143 2235 2147
rect 5265 2539 6164 2543
rect 5265 2487 5271 2539
rect 5331 2487 5335 2539
rect 5515 2487 5518 2539
rect 5579 2487 5591 2539
rect 5835 2487 5845 2539
rect 5901 2487 5911 2539
rect 6158 2487 6164 2539
rect 5265 2483 5275 2487
rect 5331 2483 5356 2487
rect 5412 2483 5437 2487
rect 5493 2483 5518 2487
rect 5574 2483 5599 2487
rect 5655 2483 5681 2487
rect 5737 2483 5763 2487
rect 5819 2483 5845 2487
rect 5901 2483 5927 2487
rect 5983 2483 6009 2487
rect 6065 2483 6091 2487
rect 6147 2483 6164 2487
rect 5265 2471 6164 2483
rect 5265 2419 5271 2471
rect 5323 2455 5335 2471
rect 5387 2455 5399 2471
rect 5451 2455 5463 2471
rect 5515 2455 5527 2471
rect 5331 2419 5335 2455
rect 5515 2419 5518 2455
rect 5579 2419 5591 2471
rect 5643 2455 5655 2471
rect 5707 2455 5719 2471
rect 5771 2455 5783 2471
rect 5835 2455 5847 2471
rect 5899 2455 5911 2471
rect 5963 2455 5976 2471
rect 6028 2455 6041 2471
rect 6093 2455 6106 2471
rect 5835 2419 5845 2455
rect 5901 2419 5911 2455
rect 6158 2419 6164 2471
rect 5265 2403 5275 2419
rect 5331 2403 5356 2419
rect 5412 2403 5437 2419
rect 5493 2403 5518 2419
rect 5574 2403 5599 2419
rect 5655 2403 5681 2419
rect 5737 2403 5763 2419
rect 5819 2403 5845 2419
rect 5901 2403 5927 2419
rect 5983 2403 6009 2419
rect 6065 2403 6091 2419
rect 6147 2403 6164 2419
rect 5265 2351 5271 2403
rect 5331 2399 5335 2403
rect 5515 2399 5518 2403
rect 5323 2371 5335 2399
rect 5387 2371 5399 2399
rect 5451 2371 5463 2399
rect 5515 2371 5527 2399
rect 5331 2351 5335 2371
rect 5515 2351 5518 2371
rect 5579 2351 5591 2403
rect 5835 2399 5845 2403
rect 5901 2399 5911 2403
rect 5643 2371 5655 2399
rect 5707 2371 5719 2399
rect 5771 2371 5783 2399
rect 5835 2371 5847 2399
rect 5899 2371 5911 2399
rect 5963 2371 5976 2399
rect 6028 2371 6041 2399
rect 6093 2371 6106 2399
rect 5835 2351 5845 2371
rect 5901 2351 5911 2371
rect 6158 2351 6164 2403
rect 5265 2335 5275 2351
rect 5331 2335 5356 2351
rect 5412 2335 5437 2351
rect 5493 2335 5518 2351
rect 5574 2335 5599 2351
rect 5655 2335 5681 2351
rect 5737 2335 5763 2351
rect 5819 2335 5845 2351
rect 5901 2335 5927 2351
rect 5983 2335 6009 2351
rect 6065 2335 6091 2351
rect 6147 2335 6164 2351
rect 5265 2283 5271 2335
rect 5331 2315 5335 2335
rect 5515 2315 5518 2335
rect 5323 2287 5335 2315
rect 5387 2287 5399 2315
rect 5451 2287 5463 2315
rect 5515 2287 5527 2315
rect 5331 2283 5335 2287
rect 5515 2283 5518 2287
rect 5579 2283 5591 2335
rect 5835 2315 5845 2335
rect 5901 2315 5911 2335
rect 5643 2287 5655 2315
rect 5707 2287 5719 2315
rect 5771 2287 5783 2315
rect 5835 2287 5847 2315
rect 5899 2287 5911 2315
rect 5963 2287 5976 2315
rect 6028 2287 6041 2315
rect 6093 2287 6106 2315
rect 5835 2283 5845 2287
rect 5901 2283 5911 2287
rect 6158 2283 6164 2335
rect 5265 2267 5275 2283
rect 5331 2267 5356 2283
rect 5412 2267 5437 2283
rect 5493 2267 5518 2283
rect 5574 2267 5599 2283
rect 5655 2267 5681 2283
rect 5737 2267 5763 2283
rect 5819 2267 5845 2283
rect 5901 2267 5927 2283
rect 5983 2267 6009 2283
rect 6065 2267 6091 2283
rect 6147 2267 6164 2283
rect 5265 2215 5271 2267
rect 5331 2231 5335 2267
rect 5515 2231 5518 2267
rect 5323 2215 5335 2231
rect 5387 2215 5399 2231
rect 5451 2215 5463 2231
rect 5515 2215 5527 2231
rect 5579 2215 5591 2267
rect 5835 2231 5845 2267
rect 5901 2231 5911 2267
rect 5643 2215 5655 2231
rect 5707 2215 5719 2231
rect 5771 2215 5783 2231
rect 5835 2215 5847 2231
rect 5899 2215 5911 2231
rect 5963 2215 5976 2231
rect 6028 2215 6041 2231
rect 6093 2215 6106 2231
rect 6158 2215 6164 2267
rect 5265 2203 6164 2215
rect 5265 2199 5275 2203
rect 5331 2199 5356 2203
rect 5412 2199 5437 2203
rect 5493 2199 5518 2203
rect 5574 2199 5599 2203
rect 5655 2199 5681 2203
rect 5737 2199 5763 2203
rect 5819 2199 5845 2203
rect 5901 2199 5927 2203
rect 5983 2199 6009 2203
rect 6065 2199 6091 2203
rect 6147 2199 6164 2203
rect 5265 2147 5271 2199
rect 5331 2147 5335 2199
rect 5515 2147 5518 2199
rect 5579 2147 5591 2199
rect 5835 2147 5845 2199
rect 5901 2147 5911 2199
rect 6158 2147 6164 2199
rect 5265 2143 6164 2147
rect 7820 2539 8719 2543
rect 7820 2487 7826 2539
rect 8073 2487 8083 2539
rect 8139 2487 8149 2539
rect 8393 2487 8405 2539
rect 8466 2487 8469 2539
rect 8649 2487 8653 2539
rect 8713 2487 8719 2539
rect 7820 2483 7837 2487
rect 7893 2483 7919 2487
rect 7975 2483 8001 2487
rect 8057 2483 8083 2487
rect 8139 2483 8165 2487
rect 8221 2483 8247 2487
rect 8303 2483 8329 2487
rect 8385 2483 8410 2487
rect 8466 2483 8491 2487
rect 8547 2483 8572 2487
rect 8628 2483 8653 2487
rect 8709 2483 8719 2487
rect 7820 2471 8719 2483
rect 7820 2419 7826 2471
rect 7878 2455 7891 2471
rect 7943 2455 7956 2471
rect 8008 2455 8021 2471
rect 8073 2455 8085 2471
rect 8137 2455 8149 2471
rect 8201 2455 8213 2471
rect 8265 2455 8277 2471
rect 8329 2455 8341 2471
rect 8073 2419 8083 2455
rect 8139 2419 8149 2455
rect 8393 2419 8405 2471
rect 8457 2455 8469 2471
rect 8521 2455 8533 2471
rect 8585 2455 8597 2471
rect 8649 2455 8661 2471
rect 8466 2419 8469 2455
rect 8649 2419 8653 2455
rect 8713 2419 8719 2471
rect 7820 2403 7837 2419
rect 7893 2403 7919 2419
rect 7975 2403 8001 2419
rect 8057 2403 8083 2419
rect 8139 2403 8165 2419
rect 8221 2403 8247 2419
rect 8303 2403 8329 2419
rect 8385 2403 8410 2419
rect 8466 2403 8491 2419
rect 8547 2403 8572 2419
rect 8628 2403 8653 2419
rect 8709 2403 8719 2419
rect 7820 2351 7826 2403
rect 8073 2399 8083 2403
rect 8139 2399 8149 2403
rect 7878 2371 7891 2399
rect 7943 2371 7956 2399
rect 8008 2371 8021 2399
rect 8073 2371 8085 2399
rect 8137 2371 8149 2399
rect 8201 2371 8213 2399
rect 8265 2371 8277 2399
rect 8329 2371 8341 2399
rect 8073 2351 8083 2371
rect 8139 2351 8149 2371
rect 8393 2351 8405 2403
rect 8466 2399 8469 2403
rect 8649 2399 8653 2403
rect 8457 2371 8469 2399
rect 8521 2371 8533 2399
rect 8585 2371 8597 2399
rect 8649 2371 8661 2399
rect 8466 2351 8469 2371
rect 8649 2351 8653 2371
rect 8713 2351 8719 2403
rect 7820 2335 7837 2351
rect 7893 2335 7919 2351
rect 7975 2335 8001 2351
rect 8057 2335 8083 2351
rect 8139 2335 8165 2351
rect 8221 2335 8247 2351
rect 8303 2335 8329 2351
rect 8385 2335 8410 2351
rect 8466 2335 8491 2351
rect 8547 2335 8572 2351
rect 8628 2335 8653 2351
rect 8709 2335 8719 2351
rect 7820 2283 7826 2335
rect 8073 2315 8083 2335
rect 8139 2315 8149 2335
rect 7878 2287 7891 2315
rect 7943 2287 7956 2315
rect 8008 2287 8021 2315
rect 8073 2287 8085 2315
rect 8137 2287 8149 2315
rect 8201 2287 8213 2315
rect 8265 2287 8277 2315
rect 8329 2287 8341 2315
rect 8073 2283 8083 2287
rect 8139 2283 8149 2287
rect 8393 2283 8405 2335
rect 8466 2315 8469 2335
rect 8649 2315 8653 2335
rect 8457 2287 8469 2315
rect 8521 2287 8533 2315
rect 8585 2287 8597 2315
rect 8649 2287 8661 2315
rect 8466 2283 8469 2287
rect 8649 2283 8653 2287
rect 8713 2283 8719 2335
rect 7820 2267 7837 2283
rect 7893 2267 7919 2283
rect 7975 2267 8001 2283
rect 8057 2267 8083 2283
rect 8139 2267 8165 2283
rect 8221 2267 8247 2283
rect 8303 2267 8329 2283
rect 8385 2267 8410 2283
rect 8466 2267 8491 2283
rect 8547 2267 8572 2283
rect 8628 2267 8653 2283
rect 8709 2267 8719 2283
rect 7820 2215 7826 2267
rect 8073 2231 8083 2267
rect 8139 2231 8149 2267
rect 7878 2215 7891 2231
rect 7943 2215 7956 2231
rect 8008 2215 8021 2231
rect 8073 2215 8085 2231
rect 8137 2215 8149 2231
rect 8201 2215 8213 2231
rect 8265 2215 8277 2231
rect 8329 2215 8341 2231
rect 8393 2215 8405 2267
rect 8466 2231 8469 2267
rect 8649 2231 8653 2267
rect 8457 2215 8469 2231
rect 8521 2215 8533 2231
rect 8585 2215 8597 2231
rect 8649 2215 8661 2231
rect 8713 2215 8719 2267
rect 7820 2203 8719 2215
rect 7820 2199 7837 2203
rect 7893 2199 7919 2203
rect 7975 2199 8001 2203
rect 8057 2199 8083 2203
rect 8139 2199 8165 2203
rect 8221 2199 8247 2203
rect 8303 2199 8329 2203
rect 8385 2199 8410 2203
rect 8466 2199 8491 2203
rect 8547 2199 8572 2203
rect 8628 2199 8653 2203
rect 8709 2199 8719 2203
rect 7820 2147 7826 2199
rect 8073 2147 8083 2199
rect 8139 2147 8149 2199
rect 8393 2147 8405 2199
rect 8466 2147 8469 2199
rect 8649 2147 8653 2199
rect 8713 2147 8719 2199
rect 7820 2143 8719 2147
rect 11749 2539 12648 2543
rect 11749 2487 11755 2539
rect 11815 2487 11819 2539
rect 11999 2487 12002 2539
rect 12063 2487 12075 2539
rect 12319 2487 12329 2539
rect 12385 2487 12395 2539
rect 12642 2487 12648 2539
rect 11749 2483 11759 2487
rect 11815 2483 11840 2487
rect 11896 2483 11921 2487
rect 11977 2483 12002 2487
rect 12058 2483 12083 2487
rect 12139 2483 12165 2487
rect 12221 2483 12247 2487
rect 12303 2483 12329 2487
rect 12385 2483 12411 2487
rect 12467 2483 12493 2487
rect 12549 2483 12575 2487
rect 12631 2483 12648 2487
rect 11749 2471 12648 2483
rect 11749 2419 11755 2471
rect 11807 2455 11819 2471
rect 11871 2455 11883 2471
rect 11935 2455 11947 2471
rect 11999 2455 12011 2471
rect 11815 2419 11819 2455
rect 11999 2419 12002 2455
rect 12063 2419 12075 2471
rect 12127 2455 12139 2471
rect 12191 2455 12203 2471
rect 12255 2455 12267 2471
rect 12319 2455 12331 2471
rect 12383 2455 12395 2471
rect 12447 2455 12460 2471
rect 12512 2455 12525 2471
rect 12577 2455 12590 2471
rect 12319 2419 12329 2455
rect 12385 2419 12395 2455
rect 12642 2419 12648 2471
rect 11749 2403 11759 2419
rect 11815 2403 11840 2419
rect 11896 2403 11921 2419
rect 11977 2403 12002 2419
rect 12058 2403 12083 2419
rect 12139 2403 12165 2419
rect 12221 2403 12247 2419
rect 12303 2403 12329 2419
rect 12385 2403 12411 2419
rect 12467 2403 12493 2419
rect 12549 2403 12575 2419
rect 12631 2403 12648 2419
rect 11749 2351 11755 2403
rect 11815 2399 11819 2403
rect 11999 2399 12002 2403
rect 11807 2371 11819 2399
rect 11871 2371 11883 2399
rect 11935 2371 11947 2399
rect 11999 2371 12011 2399
rect 11815 2351 11819 2371
rect 11999 2351 12002 2371
rect 12063 2351 12075 2403
rect 12319 2399 12329 2403
rect 12385 2399 12395 2403
rect 12127 2371 12139 2399
rect 12191 2371 12203 2399
rect 12255 2371 12267 2399
rect 12319 2371 12331 2399
rect 12383 2371 12395 2399
rect 12447 2371 12460 2399
rect 12512 2371 12525 2399
rect 12577 2371 12590 2399
rect 12319 2351 12329 2371
rect 12385 2351 12395 2371
rect 12642 2351 12648 2403
rect 11749 2335 11759 2351
rect 11815 2335 11840 2351
rect 11896 2335 11921 2351
rect 11977 2335 12002 2351
rect 12058 2335 12083 2351
rect 12139 2335 12165 2351
rect 12221 2335 12247 2351
rect 12303 2335 12329 2351
rect 12385 2335 12411 2351
rect 12467 2335 12493 2351
rect 12549 2335 12575 2351
rect 12631 2335 12648 2351
rect 11749 2283 11755 2335
rect 11815 2315 11819 2335
rect 11999 2315 12002 2335
rect 11807 2287 11819 2315
rect 11871 2287 11883 2315
rect 11935 2287 11947 2315
rect 11999 2287 12011 2315
rect 11815 2283 11819 2287
rect 11999 2283 12002 2287
rect 12063 2283 12075 2335
rect 12319 2315 12329 2335
rect 12385 2315 12395 2335
rect 12127 2287 12139 2315
rect 12191 2287 12203 2315
rect 12255 2287 12267 2315
rect 12319 2287 12331 2315
rect 12383 2287 12395 2315
rect 12447 2287 12460 2315
rect 12512 2287 12525 2315
rect 12577 2287 12590 2315
rect 12319 2283 12329 2287
rect 12385 2283 12395 2287
rect 12642 2283 12648 2335
rect 11749 2267 11759 2283
rect 11815 2267 11840 2283
rect 11896 2267 11921 2283
rect 11977 2267 12002 2283
rect 12058 2267 12083 2283
rect 12139 2267 12165 2283
rect 12221 2267 12247 2283
rect 12303 2267 12329 2283
rect 12385 2267 12411 2283
rect 12467 2267 12493 2283
rect 12549 2267 12575 2283
rect 12631 2267 12648 2283
rect 11749 2215 11755 2267
rect 11815 2231 11819 2267
rect 11999 2231 12002 2267
rect 11807 2215 11819 2231
rect 11871 2215 11883 2231
rect 11935 2215 11947 2231
rect 11999 2215 12011 2231
rect 12063 2215 12075 2267
rect 12319 2231 12329 2267
rect 12385 2231 12395 2267
rect 12127 2215 12139 2231
rect 12191 2215 12203 2231
rect 12255 2215 12267 2231
rect 12319 2215 12331 2231
rect 12383 2215 12395 2231
rect 12447 2215 12460 2231
rect 12512 2215 12525 2231
rect 12577 2215 12590 2231
rect 12642 2215 12648 2267
rect 11749 2203 12648 2215
rect 11749 2199 11759 2203
rect 11815 2199 11840 2203
rect 11896 2199 11921 2203
rect 11977 2199 12002 2203
rect 12058 2199 12083 2203
rect 12139 2199 12165 2203
rect 12221 2199 12247 2203
rect 12303 2199 12329 2203
rect 12385 2199 12411 2203
rect 12467 2199 12493 2203
rect 12549 2199 12575 2203
rect 12631 2199 12648 2203
rect 11749 2147 11755 2199
rect 11815 2147 11819 2199
rect 11999 2147 12002 2199
rect 12063 2147 12075 2199
rect 12319 2147 12329 2199
rect 12385 2147 12395 2199
rect 12642 2147 12648 2199
rect 11749 2143 12648 2147
rect 14304 2539 15203 2543
rect 14304 2487 14310 2539
rect 14557 2487 14567 2539
rect 14623 2487 14633 2539
rect 14877 2487 14889 2539
rect 14950 2487 14953 2539
rect 15133 2487 15137 2539
rect 15197 2487 15203 2539
rect 14304 2483 14321 2487
rect 14377 2483 14403 2487
rect 14459 2483 14485 2487
rect 14541 2483 14567 2487
rect 14623 2483 14649 2487
rect 14705 2483 14731 2487
rect 14787 2483 14813 2487
rect 14869 2483 14894 2487
rect 14950 2483 14975 2487
rect 15031 2483 15056 2487
rect 15112 2483 15137 2487
rect 15193 2483 15203 2487
rect 14304 2471 15203 2483
rect 14304 2419 14310 2471
rect 14362 2455 14375 2471
rect 14427 2455 14440 2471
rect 14492 2455 14505 2471
rect 14557 2455 14569 2471
rect 14621 2455 14633 2471
rect 14685 2455 14697 2471
rect 14749 2455 14761 2471
rect 14813 2455 14825 2471
rect 14557 2419 14567 2455
rect 14623 2419 14633 2455
rect 14877 2419 14889 2471
rect 14941 2455 14953 2471
rect 15005 2455 15017 2471
rect 15069 2455 15081 2471
rect 15133 2455 15145 2471
rect 14950 2419 14953 2455
rect 15133 2419 15137 2455
rect 15197 2419 15203 2471
rect 14304 2403 14321 2419
rect 14377 2403 14403 2419
rect 14459 2403 14485 2419
rect 14541 2403 14567 2419
rect 14623 2403 14649 2419
rect 14705 2403 14731 2419
rect 14787 2403 14813 2419
rect 14869 2403 14894 2419
rect 14950 2403 14975 2419
rect 15031 2403 15056 2419
rect 15112 2403 15137 2419
rect 15193 2403 15203 2419
rect 14304 2351 14310 2403
rect 14557 2399 14567 2403
rect 14623 2399 14633 2403
rect 14362 2371 14375 2399
rect 14427 2371 14440 2399
rect 14492 2371 14505 2399
rect 14557 2371 14569 2399
rect 14621 2371 14633 2399
rect 14685 2371 14697 2399
rect 14749 2371 14761 2399
rect 14813 2371 14825 2399
rect 14557 2351 14567 2371
rect 14623 2351 14633 2371
rect 14877 2351 14889 2403
rect 14950 2399 14953 2403
rect 15133 2399 15137 2403
rect 14941 2371 14953 2399
rect 15005 2371 15017 2399
rect 15069 2371 15081 2399
rect 15133 2371 15145 2399
rect 14950 2351 14953 2371
rect 15133 2351 15137 2371
rect 15197 2351 15203 2403
rect 14304 2335 14321 2351
rect 14377 2335 14403 2351
rect 14459 2335 14485 2351
rect 14541 2335 14567 2351
rect 14623 2335 14649 2351
rect 14705 2335 14731 2351
rect 14787 2335 14813 2351
rect 14869 2335 14894 2351
rect 14950 2335 14975 2351
rect 15031 2335 15056 2351
rect 15112 2335 15137 2351
rect 15193 2335 15203 2351
rect 14304 2283 14310 2335
rect 14557 2315 14567 2335
rect 14623 2315 14633 2335
rect 14362 2287 14375 2315
rect 14427 2287 14440 2315
rect 14492 2287 14505 2315
rect 14557 2287 14569 2315
rect 14621 2287 14633 2315
rect 14685 2287 14697 2315
rect 14749 2287 14761 2315
rect 14813 2287 14825 2315
rect 14557 2283 14567 2287
rect 14623 2283 14633 2287
rect 14877 2283 14889 2335
rect 14950 2315 14953 2335
rect 15133 2315 15137 2335
rect 14941 2287 14953 2315
rect 15005 2287 15017 2315
rect 15069 2287 15081 2315
rect 15133 2287 15145 2315
rect 14950 2283 14953 2287
rect 15133 2283 15137 2287
rect 15197 2283 15203 2335
rect 14304 2267 14321 2283
rect 14377 2267 14403 2283
rect 14459 2267 14485 2283
rect 14541 2267 14567 2283
rect 14623 2267 14649 2283
rect 14705 2267 14731 2283
rect 14787 2267 14813 2283
rect 14869 2267 14894 2283
rect 14950 2267 14975 2283
rect 15031 2267 15056 2283
rect 15112 2267 15137 2283
rect 15193 2267 15203 2283
rect 14304 2215 14310 2267
rect 14557 2231 14567 2267
rect 14623 2231 14633 2267
rect 14362 2215 14375 2231
rect 14427 2215 14440 2231
rect 14492 2215 14505 2231
rect 14557 2215 14569 2231
rect 14621 2215 14633 2231
rect 14685 2215 14697 2231
rect 14749 2215 14761 2231
rect 14813 2215 14825 2231
rect 14877 2215 14889 2267
rect 14950 2231 14953 2267
rect 15133 2231 15137 2267
rect 14941 2215 14953 2231
rect 15005 2215 15017 2231
rect 15069 2215 15081 2231
rect 15133 2215 15145 2231
rect 15197 2215 15203 2267
rect 14304 2203 15203 2215
rect 14304 2199 14321 2203
rect 14377 2199 14403 2203
rect 14459 2199 14485 2203
rect 14541 2199 14567 2203
rect 14623 2199 14649 2203
rect 14705 2199 14731 2203
rect 14787 2199 14813 2203
rect 14869 2199 14894 2203
rect 14950 2199 14975 2203
rect 15031 2199 15056 2203
rect 15112 2199 15137 2203
rect 15193 2199 15203 2203
rect 14304 2147 14310 2199
rect 14557 2147 14567 2199
rect 14623 2147 14633 2199
rect 14877 2147 14889 2199
rect 14950 2147 14953 2199
rect 15133 2147 15137 2199
rect 15197 2147 15203 2199
rect 14304 2143 15203 2147
rect 18233 2539 19132 2543
rect 18233 2487 18239 2539
rect 18299 2487 18303 2539
rect 18483 2487 18486 2539
rect 18547 2487 18559 2539
rect 18803 2487 18813 2539
rect 18869 2487 18879 2539
rect 19126 2487 19132 2539
rect 18233 2483 18243 2487
rect 18299 2483 18324 2487
rect 18380 2483 18405 2487
rect 18461 2483 18486 2487
rect 18542 2483 18567 2487
rect 18623 2483 18649 2487
rect 18705 2483 18731 2487
rect 18787 2483 18813 2487
rect 18869 2483 18895 2487
rect 18951 2483 18977 2487
rect 19033 2483 19059 2487
rect 19115 2483 19132 2487
rect 19925 2485 19977 2491
rect 18233 2471 19132 2483
rect 18233 2419 18239 2471
rect 18291 2455 18303 2471
rect 18355 2455 18367 2471
rect 18419 2455 18431 2471
rect 18483 2455 18495 2471
rect 18299 2419 18303 2455
rect 18483 2419 18486 2455
rect 18547 2419 18559 2471
rect 18611 2455 18623 2471
rect 18675 2455 18687 2471
rect 18739 2455 18751 2471
rect 18803 2455 18815 2471
rect 18867 2455 18879 2471
rect 18931 2455 18944 2471
rect 18996 2455 19009 2471
rect 19061 2455 19074 2471
rect 18803 2419 18813 2455
rect 18869 2419 18879 2455
rect 19126 2419 19132 2471
rect 18233 2403 18243 2419
rect 18299 2403 18324 2419
rect 18380 2403 18405 2419
rect 18461 2403 18486 2419
rect 18542 2403 18567 2419
rect 18623 2403 18649 2419
rect 18705 2403 18731 2419
rect 18787 2403 18813 2419
rect 18869 2403 18895 2419
rect 18951 2403 18977 2419
rect 19033 2403 19059 2419
rect 19115 2403 19132 2419
rect 18233 2351 18239 2403
rect 18299 2399 18303 2403
rect 18483 2399 18486 2403
rect 18291 2371 18303 2399
rect 18355 2371 18367 2399
rect 18419 2371 18431 2399
rect 18483 2371 18495 2399
rect 18299 2351 18303 2371
rect 18483 2351 18486 2371
rect 18547 2351 18559 2403
rect 18803 2399 18813 2403
rect 18869 2399 18879 2403
rect 18611 2371 18623 2399
rect 18675 2371 18687 2399
rect 18739 2371 18751 2399
rect 18803 2371 18815 2399
rect 18867 2371 18879 2399
rect 18931 2371 18944 2399
rect 18996 2371 19009 2399
rect 19061 2371 19074 2399
rect 18803 2351 18813 2371
rect 18869 2351 18879 2371
rect 19126 2351 19132 2403
rect 18233 2335 18243 2351
rect 18299 2335 18324 2351
rect 18380 2335 18405 2351
rect 18461 2335 18486 2351
rect 18542 2335 18567 2351
rect 18623 2335 18649 2351
rect 18705 2335 18731 2351
rect 18787 2335 18813 2351
rect 18869 2335 18895 2351
rect 18951 2335 18977 2351
rect 19033 2335 19059 2351
rect 19115 2335 19132 2351
rect 18233 2283 18239 2335
rect 18299 2315 18303 2335
rect 18483 2315 18486 2335
rect 18291 2287 18303 2315
rect 18355 2287 18367 2315
rect 18419 2287 18431 2315
rect 18483 2287 18495 2315
rect 18299 2283 18303 2287
rect 18483 2283 18486 2287
rect 18547 2283 18559 2335
rect 18803 2315 18813 2335
rect 18869 2315 18879 2335
rect 18611 2287 18623 2315
rect 18675 2287 18687 2315
rect 18739 2287 18751 2315
rect 18803 2287 18815 2315
rect 18867 2287 18879 2315
rect 18931 2287 18944 2315
rect 18996 2287 19009 2315
rect 19061 2287 19074 2315
rect 18803 2283 18813 2287
rect 18869 2283 18879 2287
rect 19126 2283 19132 2335
rect 18233 2267 18243 2283
rect 18299 2267 18324 2283
rect 18380 2267 18405 2283
rect 18461 2267 18486 2283
rect 18542 2267 18567 2283
rect 18623 2267 18649 2283
rect 18705 2267 18731 2283
rect 18787 2267 18813 2283
rect 18869 2267 18895 2283
rect 18951 2267 18977 2283
rect 19033 2267 19059 2283
rect 19115 2267 19132 2283
rect 18233 2215 18239 2267
rect 18299 2231 18303 2267
rect 18483 2231 18486 2267
rect 18291 2215 18303 2231
rect 18355 2215 18367 2231
rect 18419 2215 18431 2231
rect 18483 2215 18495 2231
rect 18547 2215 18559 2267
rect 18803 2231 18813 2267
rect 18869 2231 18879 2267
rect 18611 2215 18623 2231
rect 18675 2215 18687 2231
rect 18739 2215 18751 2231
rect 18803 2215 18815 2231
rect 18867 2215 18879 2231
rect 18931 2215 18944 2231
rect 18996 2215 19009 2231
rect 19061 2215 19074 2231
rect 19126 2215 19132 2267
rect 18233 2203 19132 2215
rect 18233 2199 18243 2203
rect 18299 2199 18324 2203
rect 18380 2199 18405 2203
rect 18461 2199 18486 2203
rect 18542 2199 18567 2203
rect 18623 2199 18649 2203
rect 18705 2199 18731 2203
rect 18787 2199 18813 2203
rect 18869 2199 18895 2203
rect 18951 2199 18977 2203
rect 19033 2199 19059 2203
rect 19115 2199 19132 2203
rect 18233 2147 18239 2199
rect 18299 2147 18303 2199
rect 18483 2147 18486 2199
rect 18547 2147 18559 2199
rect 18803 2147 18813 2199
rect 18869 2147 18879 2199
rect 19126 2147 19132 2199
rect 18233 2143 19132 2147
rect 19925 2195 19977 2201
rect 178 2124 511 2136
rect 230 2072 459 2124
rect 19925 2131 19977 2143
rect 19925 2073 19977 2079
rect 178 2066 511 2072
rect 953 1969 959 2021
rect 953 1965 962 1969
rect 1018 1965 1043 2021
rect 1099 1965 1123 2021
rect 1179 1965 1203 2021
rect 1262 1969 1268 2021
rect 1259 1965 1268 1969
rect 953 1957 1268 1965
rect 953 1905 959 1957
rect 1011 1905 1043 1957
rect 1095 1905 1127 1957
rect 1179 1905 1210 1957
rect 1262 1905 1268 1957
rect 953 1897 1268 1905
rect 953 1893 962 1897
rect 953 1841 959 1893
rect 1018 1841 1043 1897
rect 1099 1841 1123 1897
rect 1179 1841 1203 1897
rect 1259 1893 1268 1897
rect 1262 1841 1268 1893
rect 6327 1969 6333 2021
rect 6392 1969 6400 2021
rect 6653 1969 6661 2021
rect 6720 1969 6726 2021
rect 6327 1965 6336 1969
rect 6392 1965 6417 1969
rect 6473 1965 6498 1969
rect 6554 1965 6579 1969
rect 6635 1965 6661 1969
rect 6717 1965 6726 1969
rect 6327 1957 6726 1965
rect 6327 1905 6333 1957
rect 6385 1905 6400 1957
rect 6452 1905 6467 1957
rect 6519 1905 6534 1957
rect 6586 1905 6601 1957
rect 6653 1905 6668 1957
rect 6720 1905 6726 1957
rect 6327 1897 6726 1905
rect 6327 1893 6336 1897
rect 6392 1893 6417 1897
rect 6473 1893 6498 1897
rect 6554 1893 6579 1897
rect 6635 1893 6661 1897
rect 6717 1893 6726 1897
rect 6327 1841 6333 1893
rect 6392 1841 6400 1893
rect 6653 1841 6661 1893
rect 6720 1841 6726 1893
rect 7258 1969 7264 2021
rect 7323 1969 7331 2021
rect 7584 1969 7592 2021
rect 7651 1969 7657 2021
rect 7258 1965 7267 1969
rect 7323 1965 7349 1969
rect 7405 1965 7430 1969
rect 7486 1965 7511 1969
rect 7567 1965 7592 1969
rect 7648 1965 7657 1969
rect 7258 1957 7657 1965
rect 7258 1905 7264 1957
rect 7316 1905 7331 1957
rect 7383 1905 7398 1957
rect 7450 1905 7465 1957
rect 7517 1905 7532 1957
rect 7584 1905 7599 1957
rect 7651 1905 7657 1957
rect 7258 1897 7657 1905
rect 7258 1893 7267 1897
rect 7323 1893 7349 1897
rect 7405 1893 7430 1897
rect 7486 1893 7511 1897
rect 7567 1893 7592 1897
rect 7648 1893 7657 1897
rect 7258 1841 7264 1893
rect 7323 1841 7331 1893
rect 7584 1841 7592 1893
rect 7651 1841 7657 1893
rect 12811 1969 12817 2021
rect 12876 1969 12884 2021
rect 13137 1969 13145 2021
rect 13204 1969 13210 2021
rect 12811 1965 12820 1969
rect 12876 1965 12901 1969
rect 12957 1965 12982 1969
rect 13038 1965 13063 1969
rect 13119 1965 13145 1969
rect 13201 1965 13210 1969
rect 12811 1957 13210 1965
rect 12811 1905 12817 1957
rect 12869 1905 12884 1957
rect 12936 1905 12951 1957
rect 13003 1905 13018 1957
rect 13070 1905 13085 1957
rect 13137 1905 13152 1957
rect 13204 1905 13210 1957
rect 12811 1897 13210 1905
rect 12811 1893 12820 1897
rect 12876 1893 12901 1897
rect 12957 1893 12982 1897
rect 13038 1893 13063 1897
rect 13119 1893 13145 1897
rect 13201 1893 13210 1897
rect 12811 1841 12817 1893
rect 12876 1841 12884 1893
rect 13137 1841 13145 1893
rect 13204 1841 13210 1893
rect 13742 1969 13748 2021
rect 13807 1969 13815 2021
rect 14068 1969 14076 2021
rect 14135 1969 14141 2021
rect 13742 1965 13751 1969
rect 13807 1965 13833 1969
rect 13889 1965 13914 1969
rect 13970 1965 13995 1969
rect 14051 1965 14076 1969
rect 14132 1965 14141 1969
rect 13742 1957 14141 1965
rect 13742 1905 13748 1957
rect 13800 1905 13815 1957
rect 13867 1905 13882 1957
rect 13934 1905 13949 1957
rect 14001 1905 14016 1957
rect 14068 1905 14083 1957
rect 14135 1905 14141 1957
rect 13742 1897 14141 1905
rect 13742 1893 13751 1897
rect 13807 1893 13833 1897
rect 13889 1893 13914 1897
rect 13970 1893 13995 1897
rect 14051 1893 14076 1897
rect 14132 1893 14141 1897
rect 13742 1841 13748 1893
rect 13807 1841 13815 1893
rect 14068 1841 14076 1893
rect 14135 1841 14141 1893
rect 19380 1969 19386 2021
rect 19380 1965 19389 1969
rect 19445 1965 19469 2021
rect 19525 1965 19549 2021
rect 19605 1965 19629 2021
rect 19688 1969 19694 2021
rect 19685 1965 19694 1969
rect 19380 1957 19694 1965
rect 19380 1905 19386 1957
rect 19438 1905 19469 1957
rect 19521 1905 19552 1957
rect 19604 1905 19636 1957
rect 19688 1905 19694 1957
rect 19380 1897 19694 1905
rect 19380 1893 19389 1897
rect 19380 1841 19386 1893
rect 19445 1841 19469 1897
rect 19525 1841 19549 1897
rect 19605 1841 19629 1897
rect 19685 1893 19694 1897
rect 19688 1841 19694 1893
rect 957 -109 966 -53
rect 1022 -109 1085 -53
rect 1141 -109 1203 -53
rect 1259 -109 1268 -53
rect 957 -137 1268 -109
rect 957 -193 966 -137
rect 1022 -193 1085 -137
rect 1141 -193 1203 -137
rect 1259 -193 1268 -137
rect 6327 -109 6336 -53
rect 6392 -109 6418 -53
rect 6474 -109 6499 -53
rect 6555 -109 6580 -53
rect 6636 -109 6661 -53
rect 6717 -109 6726 -53
rect 6327 -127 6726 -109
rect 6327 -179 6333 -127
rect 6385 -137 6400 -127
rect 6452 -137 6467 -127
rect 6519 -137 6534 -127
rect 6586 -137 6601 -127
rect 6653 -137 6668 -127
rect 6392 -179 6400 -137
rect 6653 -179 6661 -137
rect 6720 -179 6726 -127
rect 6327 -193 6336 -179
rect 6392 -193 6418 -179
rect 6474 -193 6499 -179
rect 6555 -193 6580 -179
rect 6636 -193 6661 -179
rect 6717 -193 6726 -179
rect 7258 -109 7267 -53
rect 7323 -109 7349 -53
rect 7405 -109 7430 -53
rect 7486 -109 7511 -53
rect 7567 -109 7592 -53
rect 7648 -109 7657 -53
rect 7258 -127 7657 -109
rect 7258 -179 7264 -127
rect 7316 -137 7331 -127
rect 7383 -137 7398 -127
rect 7450 -137 7465 -127
rect 7517 -137 7532 -127
rect 7584 -137 7599 -127
rect 7323 -179 7331 -137
rect 7584 -179 7592 -137
rect 7651 -179 7657 -127
rect 7258 -193 7267 -179
rect 7323 -193 7349 -179
rect 7405 -193 7430 -179
rect 7486 -193 7511 -179
rect 7567 -193 7592 -179
rect 7648 -193 7657 -179
rect 12811 -109 12820 -53
rect 12876 -109 12902 -53
rect 12958 -109 12983 -53
rect 13039 -109 13064 -53
rect 13120 -109 13145 -53
rect 13201 -109 13210 -53
rect 12811 -126 13210 -109
rect 12811 -178 12817 -126
rect 12869 -137 12884 -126
rect 12936 -137 12951 -126
rect 13003 -137 13018 -126
rect 13070 -137 13085 -126
rect 13137 -137 13152 -126
rect 12876 -178 12884 -137
rect 13137 -178 13145 -137
rect 13204 -178 13210 -126
rect 12811 -193 12820 -178
rect 12876 -193 12902 -178
rect 12958 -193 12983 -178
rect 13039 -193 13064 -178
rect 13120 -193 13145 -178
rect 13201 -193 13210 -178
rect 13742 -109 13751 -53
rect 13807 -109 13833 -53
rect 13889 -109 13914 -53
rect 13970 -109 13995 -53
rect 14051 -109 14076 -53
rect 14132 -109 14141 -53
rect 13742 -127 14141 -109
rect 13742 -179 13748 -127
rect 13800 -137 13815 -127
rect 13867 -137 13882 -127
rect 13934 -137 13949 -127
rect 14001 -137 14016 -127
rect 14068 -137 14083 -127
rect 13807 -179 13815 -137
rect 14068 -179 14076 -137
rect 14135 -179 14141 -127
rect 13742 -193 13751 -179
rect 13807 -193 13833 -179
rect 13889 -193 13914 -179
rect 13970 -193 13995 -179
rect 14051 -193 14076 -179
rect 14132 -193 14141 -179
rect 19380 -109 19389 -53
rect 19445 -109 19469 -53
rect 19525 -109 19549 -53
rect 19605 -109 19629 -53
rect 19685 -109 19694 -53
rect 19380 -127 19694 -109
rect 19380 -179 19386 -127
rect 19438 -137 19470 -127
rect 19522 -137 19553 -127
rect 19605 -137 19636 -127
rect 19380 -193 19389 -179
rect 19445 -193 19469 -137
rect 19525 -193 19549 -137
rect 19605 -193 19629 -137
rect 19688 -179 19694 -127
rect 19685 -193 19694 -179
rect 12811 -1543 13210 -1538
rect 872 -1595 878 -1543
rect 930 -1595 944 -1543
rect 996 -1595 1010 -1543
rect 1062 -1595 1076 -1543
rect 1128 -1595 1141 -1543
rect 1193 -1595 1206 -1543
rect 1258 -1595 1264 -1543
rect 872 -1607 1264 -1595
rect 872 -1659 878 -1607
rect 930 -1659 944 -1607
rect 996 -1659 1010 -1607
rect 1062 -1659 1076 -1607
rect 1128 -1659 1141 -1607
rect 1193 -1659 1206 -1607
rect 1258 -1659 1264 -1607
rect 872 -1671 1264 -1659
rect 872 -1723 878 -1671
rect 930 -1723 944 -1671
rect 996 -1723 1010 -1671
rect 1062 -1723 1076 -1671
rect 1128 -1723 1141 -1671
rect 1193 -1723 1206 -1671
rect 1258 -1723 1264 -1671
rect 6328 -1595 6334 -1543
rect 6386 -1565 6400 -1543
rect 6452 -1565 6466 -1543
rect 6393 -1595 6400 -1565
rect 6518 -1595 6532 -1543
rect 6584 -1565 6597 -1543
rect 6649 -1565 6662 -1543
rect 6649 -1595 6655 -1565
rect 6714 -1595 6720 -1543
rect 6328 -1607 6337 -1595
rect 6393 -1607 6443 -1595
rect 6499 -1607 6549 -1595
rect 6605 -1607 6655 -1595
rect 6711 -1607 6720 -1595
rect 6328 -1659 6334 -1607
rect 6393 -1621 6400 -1607
rect 6386 -1645 6400 -1621
rect 6452 -1645 6466 -1621
rect 6393 -1659 6400 -1645
rect 6518 -1659 6532 -1607
rect 6649 -1621 6655 -1607
rect 6584 -1645 6597 -1621
rect 6649 -1645 6662 -1621
rect 6649 -1659 6655 -1645
rect 6714 -1659 6720 -1607
rect 6328 -1671 6337 -1659
rect 6393 -1671 6443 -1659
rect 6499 -1671 6549 -1659
rect 6605 -1671 6655 -1659
rect 6711 -1671 6720 -1659
rect 6328 -1723 6334 -1671
rect 6393 -1701 6400 -1671
rect 6386 -1723 6400 -1701
rect 6452 -1723 6466 -1701
rect 6518 -1723 6532 -1671
rect 6649 -1701 6655 -1671
rect 6584 -1723 6597 -1701
rect 6649 -1723 6662 -1701
rect 6714 -1723 6720 -1671
rect 7260 -1595 7266 -1543
rect 7318 -1565 7332 -1543
rect 7384 -1565 7398 -1543
rect 7325 -1595 7332 -1565
rect 7450 -1595 7464 -1543
rect 7516 -1565 7529 -1543
rect 7581 -1565 7594 -1543
rect 7581 -1595 7587 -1565
rect 7646 -1595 7652 -1543
rect 7260 -1607 7269 -1595
rect 7325 -1607 7375 -1595
rect 7431 -1607 7481 -1595
rect 7537 -1607 7587 -1595
rect 7643 -1607 7652 -1595
rect 7260 -1659 7266 -1607
rect 7325 -1621 7332 -1607
rect 7318 -1645 7332 -1621
rect 7384 -1645 7398 -1621
rect 7325 -1659 7332 -1645
rect 7450 -1659 7464 -1607
rect 7581 -1621 7587 -1607
rect 7516 -1645 7529 -1621
rect 7581 -1645 7594 -1621
rect 7581 -1659 7587 -1645
rect 7646 -1659 7652 -1607
rect 7260 -1671 7269 -1659
rect 7325 -1671 7375 -1659
rect 7431 -1671 7481 -1659
rect 7537 -1671 7587 -1659
rect 7643 -1671 7652 -1659
rect 7260 -1723 7266 -1671
rect 7325 -1701 7332 -1671
rect 7318 -1723 7332 -1701
rect 7384 -1723 7398 -1701
rect 7450 -1723 7464 -1671
rect 7581 -1701 7587 -1671
rect 7516 -1723 7529 -1701
rect 7581 -1723 7594 -1701
rect 7646 -1723 7652 -1671
rect 12811 -1595 12819 -1543
rect 12871 -1565 12885 -1543
rect 12937 -1565 12951 -1543
rect 13003 -1565 13017 -1543
rect 13069 -1565 13082 -1543
rect 13134 -1565 13147 -1543
rect 13199 -1565 13210 -1543
rect 12878 -1595 12885 -1565
rect 12811 -1607 12822 -1595
rect 12878 -1607 12903 -1595
rect 12959 -1607 12984 -1595
rect 12811 -1659 12819 -1607
rect 12878 -1621 12885 -1607
rect 12871 -1645 12885 -1621
rect 12937 -1645 12951 -1621
rect 12878 -1659 12885 -1645
rect 12811 -1671 12822 -1659
rect 12878 -1671 12903 -1659
rect 12959 -1671 12984 -1659
rect 12811 -1723 12819 -1671
rect 12878 -1701 12885 -1671
rect 13200 -1701 13210 -1565
rect 12871 -1723 12885 -1701
rect 12937 -1723 12951 -1701
rect 13003 -1723 13017 -1701
rect 13069 -1723 13082 -1701
rect 13134 -1723 13147 -1701
rect 13199 -1723 13210 -1701
rect 12811 -1728 13210 -1723
rect 13742 -1543 14141 -1538
rect 13742 -1595 13750 -1543
rect 13802 -1565 13816 -1543
rect 13868 -1565 13882 -1543
rect 13934 -1565 13948 -1543
rect 14000 -1565 14013 -1543
rect 14065 -1565 14078 -1543
rect 14130 -1565 14141 -1543
rect 13809 -1595 13816 -1565
rect 13742 -1607 13753 -1595
rect 13809 -1607 13834 -1595
rect 13890 -1607 13915 -1595
rect 13742 -1659 13750 -1607
rect 13809 -1621 13816 -1607
rect 13802 -1645 13816 -1621
rect 13868 -1645 13882 -1621
rect 13809 -1659 13816 -1645
rect 13742 -1671 13753 -1659
rect 13809 -1671 13834 -1659
rect 13890 -1671 13915 -1659
rect 13742 -1723 13750 -1671
rect 13809 -1701 13816 -1671
rect 14131 -1701 14141 -1565
rect 13802 -1723 13816 -1701
rect 13868 -1723 13882 -1701
rect 13934 -1723 13948 -1701
rect 14000 -1723 14013 -1701
rect 14065 -1723 14078 -1701
rect 14130 -1723 14141 -1701
rect 13742 -1728 14141 -1723
rect 19295 -1543 19694 -1538
rect 19295 -1595 19303 -1543
rect 19355 -1595 19369 -1543
rect 19421 -1565 19435 -1543
rect 19487 -1565 19501 -1543
rect 19553 -1565 19566 -1543
rect 19618 -1565 19631 -1543
rect 19683 -1565 19694 -1543
rect 19618 -1595 19628 -1565
rect 19295 -1607 19385 -1595
rect 19441 -1607 19466 -1595
rect 19522 -1607 19547 -1595
rect 19603 -1607 19628 -1595
rect 19295 -1659 19303 -1607
rect 19355 -1659 19369 -1607
rect 19618 -1621 19628 -1607
rect 19684 -1621 19694 -1565
rect 19421 -1645 19435 -1621
rect 19487 -1645 19501 -1621
rect 19553 -1645 19566 -1621
rect 19618 -1645 19631 -1621
rect 19683 -1645 19694 -1621
rect 19618 -1659 19628 -1645
rect 19295 -1671 19385 -1659
rect 19441 -1671 19466 -1659
rect 19522 -1671 19547 -1659
rect 19603 -1671 19628 -1659
rect 19295 -1723 19303 -1671
rect 19355 -1723 19369 -1671
rect 19618 -1701 19628 -1671
rect 19684 -1701 19694 -1645
rect 19421 -1723 19435 -1701
rect 19487 -1723 19501 -1701
rect 19553 -1723 19566 -1701
rect 19618 -1723 19631 -1701
rect 19683 -1723 19694 -1701
rect 19295 -1728 19694 -1723
<< rmetal2 >>
rect 19925 2728 19977 2729
rect 19925 2727 19926 2728
rect 19976 2727 19977 2728
rect 19925 2666 19926 2667
rect 19976 2666 19977 2667
rect 19925 2665 19977 2666
<< via2 >>
rect 962 4397 1018 4453
rect 1044 4397 1100 4453
rect 1126 4449 1182 4453
rect 1126 4397 1167 4449
rect 1167 4397 1182 4449
rect 1207 4397 1263 4453
rect 962 4313 1018 4369
rect 1044 4313 1100 4369
rect 1126 4317 1167 4369
rect 1167 4317 1182 4369
rect 1126 4313 1182 4317
rect 1207 4313 1263 4369
rect 6336 4449 6392 4453
rect 6418 4449 6474 4453
rect 6499 4449 6555 4453
rect 6580 4449 6636 4453
rect 6661 4449 6717 4453
rect 6336 4397 6385 4449
rect 6385 4397 6392 4449
rect 6418 4397 6452 4449
rect 6452 4397 6467 4449
rect 6467 4397 6474 4449
rect 6499 4397 6519 4449
rect 6519 4397 6534 4449
rect 6534 4397 6555 4449
rect 6580 4397 6586 4449
rect 6586 4397 6601 4449
rect 6601 4397 6636 4449
rect 6661 4397 6668 4449
rect 6668 4397 6717 4449
rect 6336 4317 6385 4369
rect 6385 4317 6392 4369
rect 6418 4317 6452 4369
rect 6452 4317 6467 4369
rect 6467 4317 6474 4369
rect 6499 4317 6519 4369
rect 6519 4317 6534 4369
rect 6534 4317 6555 4369
rect 6580 4317 6586 4369
rect 6586 4317 6601 4369
rect 6601 4317 6636 4369
rect 6661 4317 6668 4369
rect 6668 4317 6717 4369
rect 6336 4313 6392 4317
rect 6418 4313 6474 4317
rect 6499 4313 6555 4317
rect 6580 4313 6636 4317
rect 6661 4313 6717 4317
rect 7267 4449 7323 4453
rect 7349 4449 7405 4453
rect 7430 4449 7486 4453
rect 7511 4449 7567 4453
rect 7592 4449 7648 4453
rect 7267 4397 7316 4449
rect 7316 4397 7323 4449
rect 7349 4397 7383 4449
rect 7383 4397 7398 4449
rect 7398 4397 7405 4449
rect 7430 4397 7450 4449
rect 7450 4397 7465 4449
rect 7465 4397 7486 4449
rect 7511 4397 7517 4449
rect 7517 4397 7532 4449
rect 7532 4397 7567 4449
rect 7592 4397 7599 4449
rect 7599 4397 7648 4449
rect 7267 4317 7316 4369
rect 7316 4317 7323 4369
rect 7349 4317 7383 4369
rect 7383 4317 7398 4369
rect 7398 4317 7405 4369
rect 7430 4317 7450 4369
rect 7450 4317 7465 4369
rect 7465 4317 7486 4369
rect 7511 4317 7517 4369
rect 7517 4317 7532 4369
rect 7532 4317 7567 4369
rect 7592 4317 7599 4369
rect 7599 4317 7648 4369
rect 7267 4313 7323 4317
rect 7349 4313 7405 4317
rect 7430 4313 7486 4317
rect 7511 4313 7567 4317
rect 7592 4313 7648 4317
rect 12820 4449 12876 4453
rect 12902 4449 12958 4453
rect 12983 4449 13039 4453
rect 13064 4449 13120 4453
rect 13145 4449 13201 4453
rect 12820 4397 12869 4449
rect 12869 4397 12876 4449
rect 12902 4397 12936 4449
rect 12936 4397 12951 4449
rect 12951 4397 12958 4449
rect 12983 4397 13003 4449
rect 13003 4397 13018 4449
rect 13018 4397 13039 4449
rect 13064 4397 13070 4449
rect 13070 4397 13085 4449
rect 13085 4397 13120 4449
rect 13145 4397 13152 4449
rect 13152 4397 13201 4449
rect 12820 4317 12869 4369
rect 12869 4317 12876 4369
rect 12902 4317 12936 4369
rect 12936 4317 12951 4369
rect 12951 4317 12958 4369
rect 12983 4317 13003 4369
rect 13003 4317 13018 4369
rect 13018 4317 13039 4369
rect 13064 4317 13070 4369
rect 13070 4317 13085 4369
rect 13085 4317 13120 4369
rect 13145 4317 13152 4369
rect 13152 4317 13201 4369
rect 12820 4313 12876 4317
rect 12902 4313 12958 4317
rect 12983 4313 13039 4317
rect 13064 4313 13120 4317
rect 13145 4313 13201 4317
rect 13751 4449 13807 4453
rect 13833 4449 13889 4453
rect 13914 4449 13970 4453
rect 13995 4449 14051 4453
rect 14076 4449 14132 4453
rect 13751 4397 13800 4449
rect 13800 4397 13807 4449
rect 13833 4397 13867 4449
rect 13867 4397 13882 4449
rect 13882 4397 13889 4449
rect 13914 4397 13934 4449
rect 13934 4397 13949 4449
rect 13949 4397 13970 4449
rect 13995 4397 14001 4449
rect 14001 4397 14016 4449
rect 14016 4397 14051 4449
rect 14076 4397 14083 4449
rect 14083 4397 14132 4449
rect 13751 4317 13800 4369
rect 13800 4317 13807 4369
rect 13833 4317 13867 4369
rect 13867 4317 13882 4369
rect 13882 4317 13889 4369
rect 13914 4317 13934 4369
rect 13934 4317 13949 4369
rect 13949 4317 13970 4369
rect 13995 4317 14001 4369
rect 14001 4317 14016 4369
rect 14016 4317 14051 4369
rect 14076 4317 14083 4369
rect 14083 4317 14132 4369
rect 13751 4313 13807 4317
rect 13833 4313 13889 4317
rect 13914 4313 13970 4317
rect 13995 4313 14051 4317
rect 14076 4313 14132 4317
rect 19385 4449 19441 4453
rect 19385 4397 19434 4449
rect 19434 4397 19441 4449
rect 19467 4449 19523 4453
rect 19467 4397 19519 4449
rect 19519 4397 19523 4449
rect 19548 4449 19604 4453
rect 19548 4397 19552 4449
rect 19552 4397 19604 4449
rect 19629 4449 19685 4453
rect 19629 4397 19636 4449
rect 19636 4397 19685 4449
rect 19385 4317 19434 4369
rect 19434 4317 19441 4369
rect 19385 4313 19441 4317
rect 19467 4317 19519 4369
rect 19519 4317 19523 4369
rect 19467 4313 19523 4317
rect 19548 4317 19552 4369
rect 19552 4317 19604 4369
rect 19548 4313 19604 4317
rect 19629 4317 19636 4369
rect 19636 4317 19685 4369
rect 19629 4313 19685 4317
rect 962 3009 1018 3065
rect 1043 3009 1099 3065
rect 1123 3009 1179 3065
rect 1203 3009 1259 3065
rect 962 2925 1018 2981
rect 1043 2925 1099 2981
rect 1123 2925 1179 2981
rect 1203 2925 1259 2981
rect 6336 3061 6392 3065
rect 6418 3061 6474 3065
rect 6499 3061 6555 3065
rect 6580 3061 6636 3065
rect 6661 3061 6717 3065
rect 6336 3009 6385 3061
rect 6385 3009 6392 3061
rect 6418 3009 6452 3061
rect 6452 3009 6467 3061
rect 6467 3009 6474 3061
rect 6499 3009 6519 3061
rect 6519 3009 6534 3061
rect 6534 3009 6555 3061
rect 6580 3009 6586 3061
rect 6586 3009 6601 3061
rect 6601 3009 6636 3061
rect 6661 3009 6668 3061
rect 6668 3009 6717 3061
rect 6336 2929 6385 2981
rect 6385 2929 6392 2981
rect 6418 2929 6452 2981
rect 6452 2929 6467 2981
rect 6467 2929 6474 2981
rect 6499 2929 6519 2981
rect 6519 2929 6534 2981
rect 6534 2929 6555 2981
rect 6580 2929 6586 2981
rect 6586 2929 6601 2981
rect 6601 2929 6636 2981
rect 6661 2929 6668 2981
rect 6668 2929 6717 2981
rect 6336 2925 6392 2929
rect 6418 2925 6474 2929
rect 6499 2925 6555 2929
rect 6580 2925 6636 2929
rect 6661 2925 6717 2929
rect 7267 3061 7323 3065
rect 7349 3061 7405 3065
rect 7430 3061 7486 3065
rect 7511 3061 7567 3065
rect 7592 3061 7648 3065
rect 7267 3009 7316 3061
rect 7316 3009 7323 3061
rect 7349 3009 7383 3061
rect 7383 3009 7398 3061
rect 7398 3009 7405 3061
rect 7430 3009 7450 3061
rect 7450 3009 7465 3061
rect 7465 3009 7486 3061
rect 7511 3009 7517 3061
rect 7517 3009 7532 3061
rect 7532 3009 7567 3061
rect 7592 3009 7599 3061
rect 7599 3009 7648 3061
rect 7267 2929 7316 2981
rect 7316 2929 7323 2981
rect 7349 2929 7383 2981
rect 7383 2929 7398 2981
rect 7398 2929 7405 2981
rect 7430 2929 7450 2981
rect 7450 2929 7465 2981
rect 7465 2929 7486 2981
rect 7511 2929 7517 2981
rect 7517 2929 7532 2981
rect 7532 2929 7567 2981
rect 7592 2929 7599 2981
rect 7599 2929 7648 2981
rect 7267 2925 7323 2929
rect 7349 2925 7405 2929
rect 7430 2925 7486 2929
rect 7511 2925 7567 2929
rect 7592 2925 7648 2929
rect 12820 3061 12876 3065
rect 12902 3061 12958 3065
rect 12983 3061 13039 3065
rect 13064 3061 13120 3065
rect 13145 3061 13201 3065
rect 12820 3009 12869 3061
rect 12869 3009 12876 3061
rect 12902 3009 12936 3061
rect 12936 3009 12951 3061
rect 12951 3009 12958 3061
rect 12983 3009 13003 3061
rect 13003 3009 13018 3061
rect 13018 3009 13039 3061
rect 13064 3009 13070 3061
rect 13070 3009 13085 3061
rect 13085 3009 13120 3061
rect 13145 3009 13152 3061
rect 13152 3009 13201 3061
rect 12820 2929 12869 2981
rect 12869 2929 12876 2981
rect 12902 2929 12936 2981
rect 12936 2929 12951 2981
rect 12951 2929 12958 2981
rect 12983 2929 13003 2981
rect 13003 2929 13018 2981
rect 13018 2929 13039 2981
rect 13064 2929 13070 2981
rect 13070 2929 13085 2981
rect 13085 2929 13120 2981
rect 13145 2929 13152 2981
rect 13152 2929 13201 2981
rect 12820 2925 12876 2929
rect 12902 2925 12958 2929
rect 12983 2925 13039 2929
rect 13064 2925 13120 2929
rect 13145 2925 13201 2929
rect 13751 3061 13807 3065
rect 13833 3061 13889 3065
rect 13914 3061 13970 3065
rect 13995 3061 14051 3065
rect 14076 3061 14132 3065
rect 13751 3009 13800 3061
rect 13800 3009 13807 3061
rect 13833 3009 13867 3061
rect 13867 3009 13882 3061
rect 13882 3009 13889 3061
rect 13914 3009 13934 3061
rect 13934 3009 13949 3061
rect 13949 3009 13970 3061
rect 13995 3009 14001 3061
rect 14001 3009 14016 3061
rect 14016 3009 14051 3061
rect 14076 3009 14083 3061
rect 14083 3009 14132 3061
rect 13751 2929 13800 2981
rect 13800 2929 13807 2981
rect 13833 2929 13867 2981
rect 13867 2929 13882 2981
rect 13882 2929 13889 2981
rect 13914 2929 13934 2981
rect 13934 2929 13949 2981
rect 13949 2929 13970 2981
rect 13995 2929 14001 2981
rect 14001 2929 14016 2981
rect 14016 2929 14051 2981
rect 14076 2929 14083 2981
rect 14083 2929 14132 2981
rect 13751 2925 13807 2929
rect 13833 2925 13889 2929
rect 13914 2925 13970 2929
rect 13995 2925 14051 2929
rect 14076 2925 14132 2929
rect 19389 3061 19445 3065
rect 19389 3009 19438 3061
rect 19438 3009 19445 3061
rect 19469 3061 19525 3065
rect 19469 3009 19470 3061
rect 19470 3009 19522 3061
rect 19522 3009 19525 3061
rect 19549 3061 19605 3065
rect 19549 3009 19553 3061
rect 19553 3009 19605 3061
rect 19629 3061 19685 3065
rect 19629 3009 19636 3061
rect 19636 3009 19685 3061
rect 19389 2929 19438 2981
rect 19438 2929 19445 2981
rect 19389 2925 19445 2929
rect 19469 2929 19470 2981
rect 19470 2929 19522 2981
rect 19522 2929 19525 2981
rect 19469 2925 19525 2929
rect 19549 2929 19553 2981
rect 19553 2929 19605 2981
rect 19549 2925 19605 2929
rect 19629 2929 19636 2981
rect 19636 2929 19685 2981
rect 19629 2925 19685 2929
rect 962 2788 1011 2840
rect 1011 2788 1018 2840
rect 962 2784 1018 2788
rect 1043 2788 1095 2840
rect 1095 2788 1099 2840
rect 1043 2784 1099 2788
rect 1123 2788 1127 2840
rect 1127 2788 1179 2840
rect 1123 2784 1179 2788
rect 1203 2788 1210 2840
rect 1210 2788 1259 2840
rect 1203 2784 1259 2788
rect 962 2712 1018 2716
rect 962 2660 1011 2712
rect 1011 2660 1018 2712
rect 1043 2712 1099 2716
rect 1043 2660 1095 2712
rect 1095 2660 1099 2712
rect 1123 2712 1179 2716
rect 1123 2660 1127 2712
rect 1127 2660 1179 2712
rect 1203 2712 1259 2716
rect 1203 2660 1210 2712
rect 1210 2660 1259 2712
rect 6336 2788 6385 2840
rect 6385 2788 6392 2840
rect 6417 2788 6452 2840
rect 6452 2788 6467 2840
rect 6467 2788 6473 2840
rect 6498 2788 6519 2840
rect 6519 2788 6534 2840
rect 6534 2788 6554 2840
rect 6579 2788 6586 2840
rect 6586 2788 6601 2840
rect 6601 2788 6635 2840
rect 6661 2788 6668 2840
rect 6668 2788 6717 2840
rect 6336 2784 6392 2788
rect 6417 2784 6473 2788
rect 6498 2784 6554 2788
rect 6579 2784 6635 2788
rect 6661 2784 6717 2788
rect 6336 2712 6392 2716
rect 6417 2712 6473 2716
rect 6498 2712 6554 2716
rect 6579 2712 6635 2716
rect 6661 2712 6717 2716
rect 6336 2660 6385 2712
rect 6385 2660 6392 2712
rect 6417 2660 6452 2712
rect 6452 2660 6467 2712
rect 6467 2660 6473 2712
rect 6498 2660 6519 2712
rect 6519 2660 6534 2712
rect 6534 2660 6554 2712
rect 6579 2660 6586 2712
rect 6586 2660 6601 2712
rect 6601 2660 6635 2712
rect 6661 2660 6668 2712
rect 6668 2660 6717 2712
rect 7267 2788 7316 2840
rect 7316 2788 7323 2840
rect 7349 2788 7383 2840
rect 7383 2788 7398 2840
rect 7398 2788 7405 2840
rect 7430 2788 7450 2840
rect 7450 2788 7465 2840
rect 7465 2788 7486 2840
rect 7511 2788 7517 2840
rect 7517 2788 7532 2840
rect 7532 2788 7567 2840
rect 7592 2788 7599 2840
rect 7599 2788 7648 2840
rect 7267 2784 7323 2788
rect 7349 2784 7405 2788
rect 7430 2784 7486 2788
rect 7511 2784 7567 2788
rect 7592 2784 7648 2788
rect 7267 2712 7323 2716
rect 7349 2712 7405 2716
rect 7430 2712 7486 2716
rect 7511 2712 7567 2716
rect 7592 2712 7648 2716
rect 7267 2660 7316 2712
rect 7316 2660 7323 2712
rect 7349 2660 7383 2712
rect 7383 2660 7398 2712
rect 7398 2660 7405 2712
rect 7430 2660 7450 2712
rect 7450 2660 7465 2712
rect 7465 2660 7486 2712
rect 7511 2660 7517 2712
rect 7517 2660 7532 2712
rect 7532 2660 7567 2712
rect 7592 2660 7599 2712
rect 7599 2660 7648 2712
rect 12820 2788 12869 2840
rect 12869 2788 12876 2840
rect 12901 2788 12936 2840
rect 12936 2788 12951 2840
rect 12951 2788 12957 2840
rect 12982 2788 13003 2840
rect 13003 2788 13018 2840
rect 13018 2788 13038 2840
rect 13063 2788 13070 2840
rect 13070 2788 13085 2840
rect 13085 2788 13119 2840
rect 13145 2788 13152 2840
rect 13152 2788 13201 2840
rect 12820 2784 12876 2788
rect 12901 2784 12957 2788
rect 12982 2784 13038 2788
rect 13063 2784 13119 2788
rect 13145 2784 13201 2788
rect 12820 2712 12876 2716
rect 12901 2712 12957 2716
rect 12982 2712 13038 2716
rect 13063 2712 13119 2716
rect 13145 2712 13201 2716
rect 12820 2660 12869 2712
rect 12869 2660 12876 2712
rect 12901 2660 12936 2712
rect 12936 2660 12951 2712
rect 12951 2660 12957 2712
rect 12982 2660 13003 2712
rect 13003 2660 13018 2712
rect 13018 2660 13038 2712
rect 13063 2660 13070 2712
rect 13070 2660 13085 2712
rect 13085 2660 13119 2712
rect 13145 2660 13152 2712
rect 13152 2660 13201 2712
rect 13751 2788 13800 2840
rect 13800 2788 13807 2840
rect 13833 2788 13867 2840
rect 13867 2788 13882 2840
rect 13882 2788 13889 2840
rect 13914 2788 13934 2840
rect 13934 2788 13949 2840
rect 13949 2788 13970 2840
rect 13995 2788 14001 2840
rect 14001 2788 14016 2840
rect 14016 2788 14051 2840
rect 14076 2788 14083 2840
rect 14083 2788 14132 2840
rect 13751 2784 13807 2788
rect 13833 2784 13889 2788
rect 13914 2784 13970 2788
rect 13995 2784 14051 2788
rect 14076 2784 14132 2788
rect 13751 2712 13807 2716
rect 13833 2712 13889 2716
rect 13914 2712 13970 2716
rect 13995 2712 14051 2716
rect 14076 2712 14132 2716
rect 13751 2660 13800 2712
rect 13800 2660 13807 2712
rect 13833 2660 13867 2712
rect 13867 2660 13882 2712
rect 13882 2660 13889 2712
rect 13914 2660 13934 2712
rect 13934 2660 13949 2712
rect 13949 2660 13970 2712
rect 13995 2660 14001 2712
rect 14001 2660 14016 2712
rect 14016 2660 14051 2712
rect 14076 2660 14083 2712
rect 14083 2660 14132 2712
rect 19389 2788 19438 2840
rect 19438 2788 19445 2840
rect 19389 2784 19445 2788
rect 19469 2788 19521 2840
rect 19521 2788 19525 2840
rect 19469 2784 19525 2788
rect 19549 2788 19552 2840
rect 19552 2788 19604 2840
rect 19604 2788 19605 2840
rect 19549 2784 19605 2788
rect 19629 2788 19636 2840
rect 19636 2788 19685 2840
rect 19629 2784 19685 2788
rect 19389 2712 19445 2716
rect 19389 2660 19438 2712
rect 19438 2660 19445 2712
rect 19469 2712 19525 2716
rect 19469 2660 19521 2712
rect 19521 2660 19525 2712
rect 19549 2712 19605 2716
rect 19549 2660 19552 2712
rect 19552 2660 19604 2712
rect 19604 2660 19605 2712
rect 19629 2712 19685 2716
rect 19629 2660 19636 2712
rect 19636 2660 19685 2712
rect 1353 2487 1394 2539
rect 1394 2487 1407 2539
rect 1407 2487 1409 2539
rect 1435 2487 1459 2539
rect 1459 2487 1472 2539
rect 1472 2487 1491 2539
rect 1517 2487 1524 2539
rect 1524 2487 1537 2539
rect 1537 2487 1573 2539
rect 1599 2487 1601 2539
rect 1601 2487 1653 2539
rect 1653 2487 1655 2539
rect 1681 2487 1717 2539
rect 1717 2487 1729 2539
rect 1729 2487 1737 2539
rect 1763 2487 1781 2539
rect 1781 2487 1793 2539
rect 1793 2487 1819 2539
rect 1845 2487 1857 2539
rect 1857 2487 1901 2539
rect 1926 2487 1973 2539
rect 1973 2487 1982 2539
rect 2007 2487 2037 2539
rect 2037 2487 2049 2539
rect 2049 2487 2063 2539
rect 2088 2487 2101 2539
rect 2101 2487 2113 2539
rect 2113 2487 2144 2539
rect 2169 2487 2177 2539
rect 2177 2487 2225 2539
rect 1353 2483 1409 2487
rect 1435 2483 1491 2487
rect 1517 2483 1573 2487
rect 1599 2483 1655 2487
rect 1681 2483 1737 2487
rect 1763 2483 1819 2487
rect 1845 2483 1901 2487
rect 1926 2483 1982 2487
rect 2007 2483 2063 2487
rect 2088 2483 2144 2487
rect 2169 2483 2225 2487
rect 1353 2419 1394 2455
rect 1394 2419 1407 2455
rect 1407 2419 1409 2455
rect 1435 2419 1459 2455
rect 1459 2419 1472 2455
rect 1472 2419 1491 2455
rect 1517 2419 1524 2455
rect 1524 2419 1537 2455
rect 1537 2419 1573 2455
rect 1599 2419 1601 2455
rect 1601 2419 1653 2455
rect 1653 2419 1655 2455
rect 1681 2419 1717 2455
rect 1717 2419 1729 2455
rect 1729 2419 1737 2455
rect 1763 2419 1781 2455
rect 1781 2419 1793 2455
rect 1793 2419 1819 2455
rect 1845 2419 1857 2455
rect 1857 2419 1901 2455
rect 1926 2419 1973 2455
rect 1973 2419 1982 2455
rect 2007 2419 2037 2455
rect 2037 2419 2049 2455
rect 2049 2419 2063 2455
rect 2088 2419 2101 2455
rect 2101 2419 2113 2455
rect 2113 2419 2144 2455
rect 2169 2419 2177 2455
rect 2177 2419 2225 2455
rect 1353 2403 1409 2419
rect 1435 2403 1491 2419
rect 1517 2403 1573 2419
rect 1599 2403 1655 2419
rect 1681 2403 1737 2419
rect 1763 2403 1819 2419
rect 1845 2403 1901 2419
rect 1926 2403 1982 2419
rect 2007 2403 2063 2419
rect 2088 2403 2144 2419
rect 2169 2403 2225 2419
rect 1353 2399 1394 2403
rect 1394 2399 1407 2403
rect 1407 2399 1409 2403
rect 1435 2399 1459 2403
rect 1459 2399 1472 2403
rect 1472 2399 1491 2403
rect 1517 2399 1524 2403
rect 1524 2399 1537 2403
rect 1537 2399 1573 2403
rect 1599 2399 1601 2403
rect 1601 2399 1653 2403
rect 1653 2399 1655 2403
rect 1681 2399 1717 2403
rect 1717 2399 1729 2403
rect 1729 2399 1737 2403
rect 1763 2399 1781 2403
rect 1781 2399 1793 2403
rect 1793 2399 1819 2403
rect 1845 2399 1857 2403
rect 1857 2399 1901 2403
rect 1353 2351 1394 2371
rect 1394 2351 1407 2371
rect 1407 2351 1409 2371
rect 1435 2351 1459 2371
rect 1459 2351 1472 2371
rect 1472 2351 1491 2371
rect 1517 2351 1524 2371
rect 1524 2351 1537 2371
rect 1537 2351 1573 2371
rect 1599 2351 1601 2371
rect 1601 2351 1653 2371
rect 1653 2351 1655 2371
rect 1681 2351 1717 2371
rect 1717 2351 1729 2371
rect 1729 2351 1737 2371
rect 1763 2351 1781 2371
rect 1781 2351 1793 2371
rect 1793 2351 1819 2371
rect 1845 2351 1857 2371
rect 1857 2351 1901 2371
rect 1926 2399 1973 2403
rect 1973 2399 1982 2403
rect 2007 2399 2037 2403
rect 2037 2399 2049 2403
rect 2049 2399 2063 2403
rect 2088 2399 2101 2403
rect 2101 2399 2113 2403
rect 2113 2399 2144 2403
rect 2169 2399 2177 2403
rect 2177 2399 2225 2403
rect 1926 2351 1973 2371
rect 1973 2351 1982 2371
rect 2007 2351 2037 2371
rect 2037 2351 2049 2371
rect 2049 2351 2063 2371
rect 2088 2351 2101 2371
rect 2101 2351 2113 2371
rect 2113 2351 2144 2371
rect 2169 2351 2177 2371
rect 2177 2351 2225 2371
rect 1353 2335 1409 2351
rect 1435 2335 1491 2351
rect 1517 2335 1573 2351
rect 1599 2335 1655 2351
rect 1681 2335 1737 2351
rect 1763 2335 1819 2351
rect 1845 2335 1901 2351
rect 1926 2335 1982 2351
rect 2007 2335 2063 2351
rect 2088 2335 2144 2351
rect 2169 2335 2225 2351
rect 1353 2315 1394 2335
rect 1394 2315 1407 2335
rect 1407 2315 1409 2335
rect 1435 2315 1459 2335
rect 1459 2315 1472 2335
rect 1472 2315 1491 2335
rect 1517 2315 1524 2335
rect 1524 2315 1537 2335
rect 1537 2315 1573 2335
rect 1599 2315 1601 2335
rect 1601 2315 1653 2335
rect 1653 2315 1655 2335
rect 1681 2315 1717 2335
rect 1717 2315 1729 2335
rect 1729 2315 1737 2335
rect 1763 2315 1781 2335
rect 1781 2315 1793 2335
rect 1793 2315 1819 2335
rect 1845 2315 1857 2335
rect 1857 2315 1901 2335
rect 1353 2283 1394 2287
rect 1394 2283 1407 2287
rect 1407 2283 1409 2287
rect 1435 2283 1459 2287
rect 1459 2283 1472 2287
rect 1472 2283 1491 2287
rect 1517 2283 1524 2287
rect 1524 2283 1537 2287
rect 1537 2283 1573 2287
rect 1599 2283 1601 2287
rect 1601 2283 1653 2287
rect 1653 2283 1655 2287
rect 1681 2283 1717 2287
rect 1717 2283 1729 2287
rect 1729 2283 1737 2287
rect 1763 2283 1781 2287
rect 1781 2283 1793 2287
rect 1793 2283 1819 2287
rect 1845 2283 1857 2287
rect 1857 2283 1901 2287
rect 1926 2315 1973 2335
rect 1973 2315 1982 2335
rect 2007 2315 2037 2335
rect 2037 2315 2049 2335
rect 2049 2315 2063 2335
rect 2088 2315 2101 2335
rect 2101 2315 2113 2335
rect 2113 2315 2144 2335
rect 2169 2315 2177 2335
rect 2177 2315 2225 2335
rect 1926 2283 1973 2287
rect 1973 2283 1982 2287
rect 2007 2283 2037 2287
rect 2037 2283 2049 2287
rect 2049 2283 2063 2287
rect 2088 2283 2101 2287
rect 2101 2283 2113 2287
rect 2113 2283 2144 2287
rect 2169 2283 2177 2287
rect 2177 2283 2225 2287
rect 1353 2267 1409 2283
rect 1435 2267 1491 2283
rect 1517 2267 1573 2283
rect 1599 2267 1655 2283
rect 1681 2267 1737 2283
rect 1763 2267 1819 2283
rect 1845 2267 1901 2283
rect 1926 2267 1982 2283
rect 2007 2267 2063 2283
rect 2088 2267 2144 2283
rect 2169 2267 2225 2283
rect 1353 2231 1394 2267
rect 1394 2231 1407 2267
rect 1407 2231 1409 2267
rect 1435 2231 1459 2267
rect 1459 2231 1472 2267
rect 1472 2231 1491 2267
rect 1517 2231 1524 2267
rect 1524 2231 1537 2267
rect 1537 2231 1573 2267
rect 1599 2231 1601 2267
rect 1601 2231 1653 2267
rect 1653 2231 1655 2267
rect 1681 2231 1717 2267
rect 1717 2231 1729 2267
rect 1729 2231 1737 2267
rect 1763 2231 1781 2267
rect 1781 2231 1793 2267
rect 1793 2231 1819 2267
rect 1845 2231 1857 2267
rect 1857 2231 1901 2267
rect 1926 2231 1973 2267
rect 1973 2231 1982 2267
rect 2007 2231 2037 2267
rect 2037 2231 2049 2267
rect 2049 2231 2063 2267
rect 2088 2231 2101 2267
rect 2101 2231 2113 2267
rect 2113 2231 2144 2267
rect 2169 2231 2177 2267
rect 2177 2231 2225 2267
rect 1353 2199 1409 2203
rect 1435 2199 1491 2203
rect 1517 2199 1573 2203
rect 1599 2199 1655 2203
rect 1681 2199 1737 2203
rect 1763 2199 1819 2203
rect 1845 2199 1901 2203
rect 1926 2199 1982 2203
rect 2007 2199 2063 2203
rect 2088 2199 2144 2203
rect 2169 2199 2225 2203
rect 1353 2147 1394 2199
rect 1394 2147 1407 2199
rect 1407 2147 1409 2199
rect 1435 2147 1459 2199
rect 1459 2147 1472 2199
rect 1472 2147 1491 2199
rect 1517 2147 1524 2199
rect 1524 2147 1537 2199
rect 1537 2147 1573 2199
rect 1599 2147 1601 2199
rect 1601 2147 1653 2199
rect 1653 2147 1655 2199
rect 1681 2147 1717 2199
rect 1717 2147 1729 2199
rect 1729 2147 1737 2199
rect 1763 2147 1781 2199
rect 1781 2147 1793 2199
rect 1793 2147 1819 2199
rect 1845 2147 1857 2199
rect 1857 2147 1901 2199
rect 1926 2147 1973 2199
rect 1973 2147 1982 2199
rect 2007 2147 2037 2199
rect 2037 2147 2049 2199
rect 2049 2147 2063 2199
rect 2088 2147 2101 2199
rect 2101 2147 2113 2199
rect 2113 2147 2144 2199
rect 2169 2147 2177 2199
rect 2177 2147 2225 2199
rect 5275 2487 5323 2539
rect 5323 2487 5331 2539
rect 5356 2487 5387 2539
rect 5387 2487 5399 2539
rect 5399 2487 5412 2539
rect 5437 2487 5451 2539
rect 5451 2487 5463 2539
rect 5463 2487 5493 2539
rect 5518 2487 5527 2539
rect 5527 2487 5574 2539
rect 5599 2487 5643 2539
rect 5643 2487 5655 2539
rect 5681 2487 5707 2539
rect 5707 2487 5719 2539
rect 5719 2487 5737 2539
rect 5763 2487 5771 2539
rect 5771 2487 5783 2539
rect 5783 2487 5819 2539
rect 5845 2487 5847 2539
rect 5847 2487 5899 2539
rect 5899 2487 5901 2539
rect 5927 2487 5963 2539
rect 5963 2487 5976 2539
rect 5976 2487 5983 2539
rect 6009 2487 6028 2539
rect 6028 2487 6041 2539
rect 6041 2487 6065 2539
rect 6091 2487 6093 2539
rect 6093 2487 6106 2539
rect 6106 2487 6147 2539
rect 5275 2483 5331 2487
rect 5356 2483 5412 2487
rect 5437 2483 5493 2487
rect 5518 2483 5574 2487
rect 5599 2483 5655 2487
rect 5681 2483 5737 2487
rect 5763 2483 5819 2487
rect 5845 2483 5901 2487
rect 5927 2483 5983 2487
rect 6009 2483 6065 2487
rect 6091 2483 6147 2487
rect 5275 2419 5323 2455
rect 5323 2419 5331 2455
rect 5356 2419 5387 2455
rect 5387 2419 5399 2455
rect 5399 2419 5412 2455
rect 5437 2419 5451 2455
rect 5451 2419 5463 2455
rect 5463 2419 5493 2455
rect 5518 2419 5527 2455
rect 5527 2419 5574 2455
rect 5599 2419 5643 2455
rect 5643 2419 5655 2455
rect 5681 2419 5707 2455
rect 5707 2419 5719 2455
rect 5719 2419 5737 2455
rect 5763 2419 5771 2455
rect 5771 2419 5783 2455
rect 5783 2419 5819 2455
rect 5845 2419 5847 2455
rect 5847 2419 5899 2455
rect 5899 2419 5901 2455
rect 5927 2419 5963 2455
rect 5963 2419 5976 2455
rect 5976 2419 5983 2455
rect 6009 2419 6028 2455
rect 6028 2419 6041 2455
rect 6041 2419 6065 2455
rect 6091 2419 6093 2455
rect 6093 2419 6106 2455
rect 6106 2419 6147 2455
rect 5275 2403 5331 2419
rect 5356 2403 5412 2419
rect 5437 2403 5493 2419
rect 5518 2403 5574 2419
rect 5599 2403 5655 2419
rect 5681 2403 5737 2419
rect 5763 2403 5819 2419
rect 5845 2403 5901 2419
rect 5927 2403 5983 2419
rect 6009 2403 6065 2419
rect 6091 2403 6147 2419
rect 5275 2399 5323 2403
rect 5323 2399 5331 2403
rect 5356 2399 5387 2403
rect 5387 2399 5399 2403
rect 5399 2399 5412 2403
rect 5437 2399 5451 2403
rect 5451 2399 5463 2403
rect 5463 2399 5493 2403
rect 5518 2399 5527 2403
rect 5527 2399 5574 2403
rect 5275 2351 5323 2371
rect 5323 2351 5331 2371
rect 5356 2351 5387 2371
rect 5387 2351 5399 2371
rect 5399 2351 5412 2371
rect 5437 2351 5451 2371
rect 5451 2351 5463 2371
rect 5463 2351 5493 2371
rect 5518 2351 5527 2371
rect 5527 2351 5574 2371
rect 5599 2399 5643 2403
rect 5643 2399 5655 2403
rect 5681 2399 5707 2403
rect 5707 2399 5719 2403
rect 5719 2399 5737 2403
rect 5763 2399 5771 2403
rect 5771 2399 5783 2403
rect 5783 2399 5819 2403
rect 5845 2399 5847 2403
rect 5847 2399 5899 2403
rect 5899 2399 5901 2403
rect 5927 2399 5963 2403
rect 5963 2399 5976 2403
rect 5976 2399 5983 2403
rect 6009 2399 6028 2403
rect 6028 2399 6041 2403
rect 6041 2399 6065 2403
rect 6091 2399 6093 2403
rect 6093 2399 6106 2403
rect 6106 2399 6147 2403
rect 5599 2351 5643 2371
rect 5643 2351 5655 2371
rect 5681 2351 5707 2371
rect 5707 2351 5719 2371
rect 5719 2351 5737 2371
rect 5763 2351 5771 2371
rect 5771 2351 5783 2371
rect 5783 2351 5819 2371
rect 5845 2351 5847 2371
rect 5847 2351 5899 2371
rect 5899 2351 5901 2371
rect 5927 2351 5963 2371
rect 5963 2351 5976 2371
rect 5976 2351 5983 2371
rect 6009 2351 6028 2371
rect 6028 2351 6041 2371
rect 6041 2351 6065 2371
rect 6091 2351 6093 2371
rect 6093 2351 6106 2371
rect 6106 2351 6147 2371
rect 5275 2335 5331 2351
rect 5356 2335 5412 2351
rect 5437 2335 5493 2351
rect 5518 2335 5574 2351
rect 5599 2335 5655 2351
rect 5681 2335 5737 2351
rect 5763 2335 5819 2351
rect 5845 2335 5901 2351
rect 5927 2335 5983 2351
rect 6009 2335 6065 2351
rect 6091 2335 6147 2351
rect 5275 2315 5323 2335
rect 5323 2315 5331 2335
rect 5356 2315 5387 2335
rect 5387 2315 5399 2335
rect 5399 2315 5412 2335
rect 5437 2315 5451 2335
rect 5451 2315 5463 2335
rect 5463 2315 5493 2335
rect 5518 2315 5527 2335
rect 5527 2315 5574 2335
rect 5275 2283 5323 2287
rect 5323 2283 5331 2287
rect 5356 2283 5387 2287
rect 5387 2283 5399 2287
rect 5399 2283 5412 2287
rect 5437 2283 5451 2287
rect 5451 2283 5463 2287
rect 5463 2283 5493 2287
rect 5518 2283 5527 2287
rect 5527 2283 5574 2287
rect 5599 2315 5643 2335
rect 5643 2315 5655 2335
rect 5681 2315 5707 2335
rect 5707 2315 5719 2335
rect 5719 2315 5737 2335
rect 5763 2315 5771 2335
rect 5771 2315 5783 2335
rect 5783 2315 5819 2335
rect 5845 2315 5847 2335
rect 5847 2315 5899 2335
rect 5899 2315 5901 2335
rect 5927 2315 5963 2335
rect 5963 2315 5976 2335
rect 5976 2315 5983 2335
rect 6009 2315 6028 2335
rect 6028 2315 6041 2335
rect 6041 2315 6065 2335
rect 6091 2315 6093 2335
rect 6093 2315 6106 2335
rect 6106 2315 6147 2335
rect 5599 2283 5643 2287
rect 5643 2283 5655 2287
rect 5681 2283 5707 2287
rect 5707 2283 5719 2287
rect 5719 2283 5737 2287
rect 5763 2283 5771 2287
rect 5771 2283 5783 2287
rect 5783 2283 5819 2287
rect 5845 2283 5847 2287
rect 5847 2283 5899 2287
rect 5899 2283 5901 2287
rect 5927 2283 5963 2287
rect 5963 2283 5976 2287
rect 5976 2283 5983 2287
rect 6009 2283 6028 2287
rect 6028 2283 6041 2287
rect 6041 2283 6065 2287
rect 6091 2283 6093 2287
rect 6093 2283 6106 2287
rect 6106 2283 6147 2287
rect 5275 2267 5331 2283
rect 5356 2267 5412 2283
rect 5437 2267 5493 2283
rect 5518 2267 5574 2283
rect 5599 2267 5655 2283
rect 5681 2267 5737 2283
rect 5763 2267 5819 2283
rect 5845 2267 5901 2283
rect 5927 2267 5983 2283
rect 6009 2267 6065 2283
rect 6091 2267 6147 2283
rect 5275 2231 5323 2267
rect 5323 2231 5331 2267
rect 5356 2231 5387 2267
rect 5387 2231 5399 2267
rect 5399 2231 5412 2267
rect 5437 2231 5451 2267
rect 5451 2231 5463 2267
rect 5463 2231 5493 2267
rect 5518 2231 5527 2267
rect 5527 2231 5574 2267
rect 5599 2231 5643 2267
rect 5643 2231 5655 2267
rect 5681 2231 5707 2267
rect 5707 2231 5719 2267
rect 5719 2231 5737 2267
rect 5763 2231 5771 2267
rect 5771 2231 5783 2267
rect 5783 2231 5819 2267
rect 5845 2231 5847 2267
rect 5847 2231 5899 2267
rect 5899 2231 5901 2267
rect 5927 2231 5963 2267
rect 5963 2231 5976 2267
rect 5976 2231 5983 2267
rect 6009 2231 6028 2267
rect 6028 2231 6041 2267
rect 6041 2231 6065 2267
rect 6091 2231 6093 2267
rect 6093 2231 6106 2267
rect 6106 2231 6147 2267
rect 5275 2199 5331 2203
rect 5356 2199 5412 2203
rect 5437 2199 5493 2203
rect 5518 2199 5574 2203
rect 5599 2199 5655 2203
rect 5681 2199 5737 2203
rect 5763 2199 5819 2203
rect 5845 2199 5901 2203
rect 5927 2199 5983 2203
rect 6009 2199 6065 2203
rect 6091 2199 6147 2203
rect 5275 2147 5323 2199
rect 5323 2147 5331 2199
rect 5356 2147 5387 2199
rect 5387 2147 5399 2199
rect 5399 2147 5412 2199
rect 5437 2147 5451 2199
rect 5451 2147 5463 2199
rect 5463 2147 5493 2199
rect 5518 2147 5527 2199
rect 5527 2147 5574 2199
rect 5599 2147 5643 2199
rect 5643 2147 5655 2199
rect 5681 2147 5707 2199
rect 5707 2147 5719 2199
rect 5719 2147 5737 2199
rect 5763 2147 5771 2199
rect 5771 2147 5783 2199
rect 5783 2147 5819 2199
rect 5845 2147 5847 2199
rect 5847 2147 5899 2199
rect 5899 2147 5901 2199
rect 5927 2147 5963 2199
rect 5963 2147 5976 2199
rect 5976 2147 5983 2199
rect 6009 2147 6028 2199
rect 6028 2147 6041 2199
rect 6041 2147 6065 2199
rect 6091 2147 6093 2199
rect 6093 2147 6106 2199
rect 6106 2147 6147 2199
rect 7837 2487 7878 2539
rect 7878 2487 7891 2539
rect 7891 2487 7893 2539
rect 7919 2487 7943 2539
rect 7943 2487 7956 2539
rect 7956 2487 7975 2539
rect 8001 2487 8008 2539
rect 8008 2487 8021 2539
rect 8021 2487 8057 2539
rect 8083 2487 8085 2539
rect 8085 2487 8137 2539
rect 8137 2487 8139 2539
rect 8165 2487 8201 2539
rect 8201 2487 8213 2539
rect 8213 2487 8221 2539
rect 8247 2487 8265 2539
rect 8265 2487 8277 2539
rect 8277 2487 8303 2539
rect 8329 2487 8341 2539
rect 8341 2487 8385 2539
rect 8410 2487 8457 2539
rect 8457 2487 8466 2539
rect 8491 2487 8521 2539
rect 8521 2487 8533 2539
rect 8533 2487 8547 2539
rect 8572 2487 8585 2539
rect 8585 2487 8597 2539
rect 8597 2487 8628 2539
rect 8653 2487 8661 2539
rect 8661 2487 8709 2539
rect 7837 2483 7893 2487
rect 7919 2483 7975 2487
rect 8001 2483 8057 2487
rect 8083 2483 8139 2487
rect 8165 2483 8221 2487
rect 8247 2483 8303 2487
rect 8329 2483 8385 2487
rect 8410 2483 8466 2487
rect 8491 2483 8547 2487
rect 8572 2483 8628 2487
rect 8653 2483 8709 2487
rect 7837 2419 7878 2455
rect 7878 2419 7891 2455
rect 7891 2419 7893 2455
rect 7919 2419 7943 2455
rect 7943 2419 7956 2455
rect 7956 2419 7975 2455
rect 8001 2419 8008 2455
rect 8008 2419 8021 2455
rect 8021 2419 8057 2455
rect 8083 2419 8085 2455
rect 8085 2419 8137 2455
rect 8137 2419 8139 2455
rect 8165 2419 8201 2455
rect 8201 2419 8213 2455
rect 8213 2419 8221 2455
rect 8247 2419 8265 2455
rect 8265 2419 8277 2455
rect 8277 2419 8303 2455
rect 8329 2419 8341 2455
rect 8341 2419 8385 2455
rect 8410 2419 8457 2455
rect 8457 2419 8466 2455
rect 8491 2419 8521 2455
rect 8521 2419 8533 2455
rect 8533 2419 8547 2455
rect 8572 2419 8585 2455
rect 8585 2419 8597 2455
rect 8597 2419 8628 2455
rect 8653 2419 8661 2455
rect 8661 2419 8709 2455
rect 7837 2403 7893 2419
rect 7919 2403 7975 2419
rect 8001 2403 8057 2419
rect 8083 2403 8139 2419
rect 8165 2403 8221 2419
rect 8247 2403 8303 2419
rect 8329 2403 8385 2419
rect 8410 2403 8466 2419
rect 8491 2403 8547 2419
rect 8572 2403 8628 2419
rect 8653 2403 8709 2419
rect 7837 2399 7878 2403
rect 7878 2399 7891 2403
rect 7891 2399 7893 2403
rect 7919 2399 7943 2403
rect 7943 2399 7956 2403
rect 7956 2399 7975 2403
rect 8001 2399 8008 2403
rect 8008 2399 8021 2403
rect 8021 2399 8057 2403
rect 8083 2399 8085 2403
rect 8085 2399 8137 2403
rect 8137 2399 8139 2403
rect 8165 2399 8201 2403
rect 8201 2399 8213 2403
rect 8213 2399 8221 2403
rect 8247 2399 8265 2403
rect 8265 2399 8277 2403
rect 8277 2399 8303 2403
rect 8329 2399 8341 2403
rect 8341 2399 8385 2403
rect 7837 2351 7878 2371
rect 7878 2351 7891 2371
rect 7891 2351 7893 2371
rect 7919 2351 7943 2371
rect 7943 2351 7956 2371
rect 7956 2351 7975 2371
rect 8001 2351 8008 2371
rect 8008 2351 8021 2371
rect 8021 2351 8057 2371
rect 8083 2351 8085 2371
rect 8085 2351 8137 2371
rect 8137 2351 8139 2371
rect 8165 2351 8201 2371
rect 8201 2351 8213 2371
rect 8213 2351 8221 2371
rect 8247 2351 8265 2371
rect 8265 2351 8277 2371
rect 8277 2351 8303 2371
rect 8329 2351 8341 2371
rect 8341 2351 8385 2371
rect 8410 2399 8457 2403
rect 8457 2399 8466 2403
rect 8491 2399 8521 2403
rect 8521 2399 8533 2403
rect 8533 2399 8547 2403
rect 8572 2399 8585 2403
rect 8585 2399 8597 2403
rect 8597 2399 8628 2403
rect 8653 2399 8661 2403
rect 8661 2399 8709 2403
rect 8410 2351 8457 2371
rect 8457 2351 8466 2371
rect 8491 2351 8521 2371
rect 8521 2351 8533 2371
rect 8533 2351 8547 2371
rect 8572 2351 8585 2371
rect 8585 2351 8597 2371
rect 8597 2351 8628 2371
rect 8653 2351 8661 2371
rect 8661 2351 8709 2371
rect 7837 2335 7893 2351
rect 7919 2335 7975 2351
rect 8001 2335 8057 2351
rect 8083 2335 8139 2351
rect 8165 2335 8221 2351
rect 8247 2335 8303 2351
rect 8329 2335 8385 2351
rect 8410 2335 8466 2351
rect 8491 2335 8547 2351
rect 8572 2335 8628 2351
rect 8653 2335 8709 2351
rect 7837 2315 7878 2335
rect 7878 2315 7891 2335
rect 7891 2315 7893 2335
rect 7919 2315 7943 2335
rect 7943 2315 7956 2335
rect 7956 2315 7975 2335
rect 8001 2315 8008 2335
rect 8008 2315 8021 2335
rect 8021 2315 8057 2335
rect 8083 2315 8085 2335
rect 8085 2315 8137 2335
rect 8137 2315 8139 2335
rect 8165 2315 8201 2335
rect 8201 2315 8213 2335
rect 8213 2315 8221 2335
rect 8247 2315 8265 2335
rect 8265 2315 8277 2335
rect 8277 2315 8303 2335
rect 8329 2315 8341 2335
rect 8341 2315 8385 2335
rect 7837 2283 7878 2287
rect 7878 2283 7891 2287
rect 7891 2283 7893 2287
rect 7919 2283 7943 2287
rect 7943 2283 7956 2287
rect 7956 2283 7975 2287
rect 8001 2283 8008 2287
rect 8008 2283 8021 2287
rect 8021 2283 8057 2287
rect 8083 2283 8085 2287
rect 8085 2283 8137 2287
rect 8137 2283 8139 2287
rect 8165 2283 8201 2287
rect 8201 2283 8213 2287
rect 8213 2283 8221 2287
rect 8247 2283 8265 2287
rect 8265 2283 8277 2287
rect 8277 2283 8303 2287
rect 8329 2283 8341 2287
rect 8341 2283 8385 2287
rect 8410 2315 8457 2335
rect 8457 2315 8466 2335
rect 8491 2315 8521 2335
rect 8521 2315 8533 2335
rect 8533 2315 8547 2335
rect 8572 2315 8585 2335
rect 8585 2315 8597 2335
rect 8597 2315 8628 2335
rect 8653 2315 8661 2335
rect 8661 2315 8709 2335
rect 8410 2283 8457 2287
rect 8457 2283 8466 2287
rect 8491 2283 8521 2287
rect 8521 2283 8533 2287
rect 8533 2283 8547 2287
rect 8572 2283 8585 2287
rect 8585 2283 8597 2287
rect 8597 2283 8628 2287
rect 8653 2283 8661 2287
rect 8661 2283 8709 2287
rect 7837 2267 7893 2283
rect 7919 2267 7975 2283
rect 8001 2267 8057 2283
rect 8083 2267 8139 2283
rect 8165 2267 8221 2283
rect 8247 2267 8303 2283
rect 8329 2267 8385 2283
rect 8410 2267 8466 2283
rect 8491 2267 8547 2283
rect 8572 2267 8628 2283
rect 8653 2267 8709 2283
rect 7837 2231 7878 2267
rect 7878 2231 7891 2267
rect 7891 2231 7893 2267
rect 7919 2231 7943 2267
rect 7943 2231 7956 2267
rect 7956 2231 7975 2267
rect 8001 2231 8008 2267
rect 8008 2231 8021 2267
rect 8021 2231 8057 2267
rect 8083 2231 8085 2267
rect 8085 2231 8137 2267
rect 8137 2231 8139 2267
rect 8165 2231 8201 2267
rect 8201 2231 8213 2267
rect 8213 2231 8221 2267
rect 8247 2231 8265 2267
rect 8265 2231 8277 2267
rect 8277 2231 8303 2267
rect 8329 2231 8341 2267
rect 8341 2231 8385 2267
rect 8410 2231 8457 2267
rect 8457 2231 8466 2267
rect 8491 2231 8521 2267
rect 8521 2231 8533 2267
rect 8533 2231 8547 2267
rect 8572 2231 8585 2267
rect 8585 2231 8597 2267
rect 8597 2231 8628 2267
rect 8653 2231 8661 2267
rect 8661 2231 8709 2267
rect 7837 2199 7893 2203
rect 7919 2199 7975 2203
rect 8001 2199 8057 2203
rect 8083 2199 8139 2203
rect 8165 2199 8221 2203
rect 8247 2199 8303 2203
rect 8329 2199 8385 2203
rect 8410 2199 8466 2203
rect 8491 2199 8547 2203
rect 8572 2199 8628 2203
rect 8653 2199 8709 2203
rect 7837 2147 7878 2199
rect 7878 2147 7891 2199
rect 7891 2147 7893 2199
rect 7919 2147 7943 2199
rect 7943 2147 7956 2199
rect 7956 2147 7975 2199
rect 8001 2147 8008 2199
rect 8008 2147 8021 2199
rect 8021 2147 8057 2199
rect 8083 2147 8085 2199
rect 8085 2147 8137 2199
rect 8137 2147 8139 2199
rect 8165 2147 8201 2199
rect 8201 2147 8213 2199
rect 8213 2147 8221 2199
rect 8247 2147 8265 2199
rect 8265 2147 8277 2199
rect 8277 2147 8303 2199
rect 8329 2147 8341 2199
rect 8341 2147 8385 2199
rect 8410 2147 8457 2199
rect 8457 2147 8466 2199
rect 8491 2147 8521 2199
rect 8521 2147 8533 2199
rect 8533 2147 8547 2199
rect 8572 2147 8585 2199
rect 8585 2147 8597 2199
rect 8597 2147 8628 2199
rect 8653 2147 8661 2199
rect 8661 2147 8709 2199
rect 11759 2487 11807 2539
rect 11807 2487 11815 2539
rect 11840 2487 11871 2539
rect 11871 2487 11883 2539
rect 11883 2487 11896 2539
rect 11921 2487 11935 2539
rect 11935 2487 11947 2539
rect 11947 2487 11977 2539
rect 12002 2487 12011 2539
rect 12011 2487 12058 2539
rect 12083 2487 12127 2539
rect 12127 2487 12139 2539
rect 12165 2487 12191 2539
rect 12191 2487 12203 2539
rect 12203 2487 12221 2539
rect 12247 2487 12255 2539
rect 12255 2487 12267 2539
rect 12267 2487 12303 2539
rect 12329 2487 12331 2539
rect 12331 2487 12383 2539
rect 12383 2487 12385 2539
rect 12411 2487 12447 2539
rect 12447 2487 12460 2539
rect 12460 2487 12467 2539
rect 12493 2487 12512 2539
rect 12512 2487 12525 2539
rect 12525 2487 12549 2539
rect 12575 2487 12577 2539
rect 12577 2487 12590 2539
rect 12590 2487 12631 2539
rect 11759 2483 11815 2487
rect 11840 2483 11896 2487
rect 11921 2483 11977 2487
rect 12002 2483 12058 2487
rect 12083 2483 12139 2487
rect 12165 2483 12221 2487
rect 12247 2483 12303 2487
rect 12329 2483 12385 2487
rect 12411 2483 12467 2487
rect 12493 2483 12549 2487
rect 12575 2483 12631 2487
rect 11759 2419 11807 2455
rect 11807 2419 11815 2455
rect 11840 2419 11871 2455
rect 11871 2419 11883 2455
rect 11883 2419 11896 2455
rect 11921 2419 11935 2455
rect 11935 2419 11947 2455
rect 11947 2419 11977 2455
rect 12002 2419 12011 2455
rect 12011 2419 12058 2455
rect 12083 2419 12127 2455
rect 12127 2419 12139 2455
rect 12165 2419 12191 2455
rect 12191 2419 12203 2455
rect 12203 2419 12221 2455
rect 12247 2419 12255 2455
rect 12255 2419 12267 2455
rect 12267 2419 12303 2455
rect 12329 2419 12331 2455
rect 12331 2419 12383 2455
rect 12383 2419 12385 2455
rect 12411 2419 12447 2455
rect 12447 2419 12460 2455
rect 12460 2419 12467 2455
rect 12493 2419 12512 2455
rect 12512 2419 12525 2455
rect 12525 2419 12549 2455
rect 12575 2419 12577 2455
rect 12577 2419 12590 2455
rect 12590 2419 12631 2455
rect 11759 2403 11815 2419
rect 11840 2403 11896 2419
rect 11921 2403 11977 2419
rect 12002 2403 12058 2419
rect 12083 2403 12139 2419
rect 12165 2403 12221 2419
rect 12247 2403 12303 2419
rect 12329 2403 12385 2419
rect 12411 2403 12467 2419
rect 12493 2403 12549 2419
rect 12575 2403 12631 2419
rect 11759 2399 11807 2403
rect 11807 2399 11815 2403
rect 11840 2399 11871 2403
rect 11871 2399 11883 2403
rect 11883 2399 11896 2403
rect 11921 2399 11935 2403
rect 11935 2399 11947 2403
rect 11947 2399 11977 2403
rect 12002 2399 12011 2403
rect 12011 2399 12058 2403
rect 11759 2351 11807 2371
rect 11807 2351 11815 2371
rect 11840 2351 11871 2371
rect 11871 2351 11883 2371
rect 11883 2351 11896 2371
rect 11921 2351 11935 2371
rect 11935 2351 11947 2371
rect 11947 2351 11977 2371
rect 12002 2351 12011 2371
rect 12011 2351 12058 2371
rect 12083 2399 12127 2403
rect 12127 2399 12139 2403
rect 12165 2399 12191 2403
rect 12191 2399 12203 2403
rect 12203 2399 12221 2403
rect 12247 2399 12255 2403
rect 12255 2399 12267 2403
rect 12267 2399 12303 2403
rect 12329 2399 12331 2403
rect 12331 2399 12383 2403
rect 12383 2399 12385 2403
rect 12411 2399 12447 2403
rect 12447 2399 12460 2403
rect 12460 2399 12467 2403
rect 12493 2399 12512 2403
rect 12512 2399 12525 2403
rect 12525 2399 12549 2403
rect 12575 2399 12577 2403
rect 12577 2399 12590 2403
rect 12590 2399 12631 2403
rect 12083 2351 12127 2371
rect 12127 2351 12139 2371
rect 12165 2351 12191 2371
rect 12191 2351 12203 2371
rect 12203 2351 12221 2371
rect 12247 2351 12255 2371
rect 12255 2351 12267 2371
rect 12267 2351 12303 2371
rect 12329 2351 12331 2371
rect 12331 2351 12383 2371
rect 12383 2351 12385 2371
rect 12411 2351 12447 2371
rect 12447 2351 12460 2371
rect 12460 2351 12467 2371
rect 12493 2351 12512 2371
rect 12512 2351 12525 2371
rect 12525 2351 12549 2371
rect 12575 2351 12577 2371
rect 12577 2351 12590 2371
rect 12590 2351 12631 2371
rect 11759 2335 11815 2351
rect 11840 2335 11896 2351
rect 11921 2335 11977 2351
rect 12002 2335 12058 2351
rect 12083 2335 12139 2351
rect 12165 2335 12221 2351
rect 12247 2335 12303 2351
rect 12329 2335 12385 2351
rect 12411 2335 12467 2351
rect 12493 2335 12549 2351
rect 12575 2335 12631 2351
rect 11759 2315 11807 2335
rect 11807 2315 11815 2335
rect 11840 2315 11871 2335
rect 11871 2315 11883 2335
rect 11883 2315 11896 2335
rect 11921 2315 11935 2335
rect 11935 2315 11947 2335
rect 11947 2315 11977 2335
rect 12002 2315 12011 2335
rect 12011 2315 12058 2335
rect 11759 2283 11807 2287
rect 11807 2283 11815 2287
rect 11840 2283 11871 2287
rect 11871 2283 11883 2287
rect 11883 2283 11896 2287
rect 11921 2283 11935 2287
rect 11935 2283 11947 2287
rect 11947 2283 11977 2287
rect 12002 2283 12011 2287
rect 12011 2283 12058 2287
rect 12083 2315 12127 2335
rect 12127 2315 12139 2335
rect 12165 2315 12191 2335
rect 12191 2315 12203 2335
rect 12203 2315 12221 2335
rect 12247 2315 12255 2335
rect 12255 2315 12267 2335
rect 12267 2315 12303 2335
rect 12329 2315 12331 2335
rect 12331 2315 12383 2335
rect 12383 2315 12385 2335
rect 12411 2315 12447 2335
rect 12447 2315 12460 2335
rect 12460 2315 12467 2335
rect 12493 2315 12512 2335
rect 12512 2315 12525 2335
rect 12525 2315 12549 2335
rect 12575 2315 12577 2335
rect 12577 2315 12590 2335
rect 12590 2315 12631 2335
rect 12083 2283 12127 2287
rect 12127 2283 12139 2287
rect 12165 2283 12191 2287
rect 12191 2283 12203 2287
rect 12203 2283 12221 2287
rect 12247 2283 12255 2287
rect 12255 2283 12267 2287
rect 12267 2283 12303 2287
rect 12329 2283 12331 2287
rect 12331 2283 12383 2287
rect 12383 2283 12385 2287
rect 12411 2283 12447 2287
rect 12447 2283 12460 2287
rect 12460 2283 12467 2287
rect 12493 2283 12512 2287
rect 12512 2283 12525 2287
rect 12525 2283 12549 2287
rect 12575 2283 12577 2287
rect 12577 2283 12590 2287
rect 12590 2283 12631 2287
rect 11759 2267 11815 2283
rect 11840 2267 11896 2283
rect 11921 2267 11977 2283
rect 12002 2267 12058 2283
rect 12083 2267 12139 2283
rect 12165 2267 12221 2283
rect 12247 2267 12303 2283
rect 12329 2267 12385 2283
rect 12411 2267 12467 2283
rect 12493 2267 12549 2283
rect 12575 2267 12631 2283
rect 11759 2231 11807 2267
rect 11807 2231 11815 2267
rect 11840 2231 11871 2267
rect 11871 2231 11883 2267
rect 11883 2231 11896 2267
rect 11921 2231 11935 2267
rect 11935 2231 11947 2267
rect 11947 2231 11977 2267
rect 12002 2231 12011 2267
rect 12011 2231 12058 2267
rect 12083 2231 12127 2267
rect 12127 2231 12139 2267
rect 12165 2231 12191 2267
rect 12191 2231 12203 2267
rect 12203 2231 12221 2267
rect 12247 2231 12255 2267
rect 12255 2231 12267 2267
rect 12267 2231 12303 2267
rect 12329 2231 12331 2267
rect 12331 2231 12383 2267
rect 12383 2231 12385 2267
rect 12411 2231 12447 2267
rect 12447 2231 12460 2267
rect 12460 2231 12467 2267
rect 12493 2231 12512 2267
rect 12512 2231 12525 2267
rect 12525 2231 12549 2267
rect 12575 2231 12577 2267
rect 12577 2231 12590 2267
rect 12590 2231 12631 2267
rect 11759 2199 11815 2203
rect 11840 2199 11896 2203
rect 11921 2199 11977 2203
rect 12002 2199 12058 2203
rect 12083 2199 12139 2203
rect 12165 2199 12221 2203
rect 12247 2199 12303 2203
rect 12329 2199 12385 2203
rect 12411 2199 12467 2203
rect 12493 2199 12549 2203
rect 12575 2199 12631 2203
rect 11759 2147 11807 2199
rect 11807 2147 11815 2199
rect 11840 2147 11871 2199
rect 11871 2147 11883 2199
rect 11883 2147 11896 2199
rect 11921 2147 11935 2199
rect 11935 2147 11947 2199
rect 11947 2147 11977 2199
rect 12002 2147 12011 2199
rect 12011 2147 12058 2199
rect 12083 2147 12127 2199
rect 12127 2147 12139 2199
rect 12165 2147 12191 2199
rect 12191 2147 12203 2199
rect 12203 2147 12221 2199
rect 12247 2147 12255 2199
rect 12255 2147 12267 2199
rect 12267 2147 12303 2199
rect 12329 2147 12331 2199
rect 12331 2147 12383 2199
rect 12383 2147 12385 2199
rect 12411 2147 12447 2199
rect 12447 2147 12460 2199
rect 12460 2147 12467 2199
rect 12493 2147 12512 2199
rect 12512 2147 12525 2199
rect 12525 2147 12549 2199
rect 12575 2147 12577 2199
rect 12577 2147 12590 2199
rect 12590 2147 12631 2199
rect 14321 2487 14362 2539
rect 14362 2487 14375 2539
rect 14375 2487 14377 2539
rect 14403 2487 14427 2539
rect 14427 2487 14440 2539
rect 14440 2487 14459 2539
rect 14485 2487 14492 2539
rect 14492 2487 14505 2539
rect 14505 2487 14541 2539
rect 14567 2487 14569 2539
rect 14569 2487 14621 2539
rect 14621 2487 14623 2539
rect 14649 2487 14685 2539
rect 14685 2487 14697 2539
rect 14697 2487 14705 2539
rect 14731 2487 14749 2539
rect 14749 2487 14761 2539
rect 14761 2487 14787 2539
rect 14813 2487 14825 2539
rect 14825 2487 14869 2539
rect 14894 2487 14941 2539
rect 14941 2487 14950 2539
rect 14975 2487 15005 2539
rect 15005 2487 15017 2539
rect 15017 2487 15031 2539
rect 15056 2487 15069 2539
rect 15069 2487 15081 2539
rect 15081 2487 15112 2539
rect 15137 2487 15145 2539
rect 15145 2487 15193 2539
rect 14321 2483 14377 2487
rect 14403 2483 14459 2487
rect 14485 2483 14541 2487
rect 14567 2483 14623 2487
rect 14649 2483 14705 2487
rect 14731 2483 14787 2487
rect 14813 2483 14869 2487
rect 14894 2483 14950 2487
rect 14975 2483 15031 2487
rect 15056 2483 15112 2487
rect 15137 2483 15193 2487
rect 14321 2419 14362 2455
rect 14362 2419 14375 2455
rect 14375 2419 14377 2455
rect 14403 2419 14427 2455
rect 14427 2419 14440 2455
rect 14440 2419 14459 2455
rect 14485 2419 14492 2455
rect 14492 2419 14505 2455
rect 14505 2419 14541 2455
rect 14567 2419 14569 2455
rect 14569 2419 14621 2455
rect 14621 2419 14623 2455
rect 14649 2419 14685 2455
rect 14685 2419 14697 2455
rect 14697 2419 14705 2455
rect 14731 2419 14749 2455
rect 14749 2419 14761 2455
rect 14761 2419 14787 2455
rect 14813 2419 14825 2455
rect 14825 2419 14869 2455
rect 14894 2419 14941 2455
rect 14941 2419 14950 2455
rect 14975 2419 15005 2455
rect 15005 2419 15017 2455
rect 15017 2419 15031 2455
rect 15056 2419 15069 2455
rect 15069 2419 15081 2455
rect 15081 2419 15112 2455
rect 15137 2419 15145 2455
rect 15145 2419 15193 2455
rect 14321 2403 14377 2419
rect 14403 2403 14459 2419
rect 14485 2403 14541 2419
rect 14567 2403 14623 2419
rect 14649 2403 14705 2419
rect 14731 2403 14787 2419
rect 14813 2403 14869 2419
rect 14894 2403 14950 2419
rect 14975 2403 15031 2419
rect 15056 2403 15112 2419
rect 15137 2403 15193 2419
rect 14321 2399 14362 2403
rect 14362 2399 14375 2403
rect 14375 2399 14377 2403
rect 14403 2399 14427 2403
rect 14427 2399 14440 2403
rect 14440 2399 14459 2403
rect 14485 2399 14492 2403
rect 14492 2399 14505 2403
rect 14505 2399 14541 2403
rect 14567 2399 14569 2403
rect 14569 2399 14621 2403
rect 14621 2399 14623 2403
rect 14649 2399 14685 2403
rect 14685 2399 14697 2403
rect 14697 2399 14705 2403
rect 14731 2399 14749 2403
rect 14749 2399 14761 2403
rect 14761 2399 14787 2403
rect 14813 2399 14825 2403
rect 14825 2399 14869 2403
rect 14321 2351 14362 2371
rect 14362 2351 14375 2371
rect 14375 2351 14377 2371
rect 14403 2351 14427 2371
rect 14427 2351 14440 2371
rect 14440 2351 14459 2371
rect 14485 2351 14492 2371
rect 14492 2351 14505 2371
rect 14505 2351 14541 2371
rect 14567 2351 14569 2371
rect 14569 2351 14621 2371
rect 14621 2351 14623 2371
rect 14649 2351 14685 2371
rect 14685 2351 14697 2371
rect 14697 2351 14705 2371
rect 14731 2351 14749 2371
rect 14749 2351 14761 2371
rect 14761 2351 14787 2371
rect 14813 2351 14825 2371
rect 14825 2351 14869 2371
rect 14894 2399 14941 2403
rect 14941 2399 14950 2403
rect 14975 2399 15005 2403
rect 15005 2399 15017 2403
rect 15017 2399 15031 2403
rect 15056 2399 15069 2403
rect 15069 2399 15081 2403
rect 15081 2399 15112 2403
rect 15137 2399 15145 2403
rect 15145 2399 15193 2403
rect 14894 2351 14941 2371
rect 14941 2351 14950 2371
rect 14975 2351 15005 2371
rect 15005 2351 15017 2371
rect 15017 2351 15031 2371
rect 15056 2351 15069 2371
rect 15069 2351 15081 2371
rect 15081 2351 15112 2371
rect 15137 2351 15145 2371
rect 15145 2351 15193 2371
rect 14321 2335 14377 2351
rect 14403 2335 14459 2351
rect 14485 2335 14541 2351
rect 14567 2335 14623 2351
rect 14649 2335 14705 2351
rect 14731 2335 14787 2351
rect 14813 2335 14869 2351
rect 14894 2335 14950 2351
rect 14975 2335 15031 2351
rect 15056 2335 15112 2351
rect 15137 2335 15193 2351
rect 14321 2315 14362 2335
rect 14362 2315 14375 2335
rect 14375 2315 14377 2335
rect 14403 2315 14427 2335
rect 14427 2315 14440 2335
rect 14440 2315 14459 2335
rect 14485 2315 14492 2335
rect 14492 2315 14505 2335
rect 14505 2315 14541 2335
rect 14567 2315 14569 2335
rect 14569 2315 14621 2335
rect 14621 2315 14623 2335
rect 14649 2315 14685 2335
rect 14685 2315 14697 2335
rect 14697 2315 14705 2335
rect 14731 2315 14749 2335
rect 14749 2315 14761 2335
rect 14761 2315 14787 2335
rect 14813 2315 14825 2335
rect 14825 2315 14869 2335
rect 14321 2283 14362 2287
rect 14362 2283 14375 2287
rect 14375 2283 14377 2287
rect 14403 2283 14427 2287
rect 14427 2283 14440 2287
rect 14440 2283 14459 2287
rect 14485 2283 14492 2287
rect 14492 2283 14505 2287
rect 14505 2283 14541 2287
rect 14567 2283 14569 2287
rect 14569 2283 14621 2287
rect 14621 2283 14623 2287
rect 14649 2283 14685 2287
rect 14685 2283 14697 2287
rect 14697 2283 14705 2287
rect 14731 2283 14749 2287
rect 14749 2283 14761 2287
rect 14761 2283 14787 2287
rect 14813 2283 14825 2287
rect 14825 2283 14869 2287
rect 14894 2315 14941 2335
rect 14941 2315 14950 2335
rect 14975 2315 15005 2335
rect 15005 2315 15017 2335
rect 15017 2315 15031 2335
rect 15056 2315 15069 2335
rect 15069 2315 15081 2335
rect 15081 2315 15112 2335
rect 15137 2315 15145 2335
rect 15145 2315 15193 2335
rect 14894 2283 14941 2287
rect 14941 2283 14950 2287
rect 14975 2283 15005 2287
rect 15005 2283 15017 2287
rect 15017 2283 15031 2287
rect 15056 2283 15069 2287
rect 15069 2283 15081 2287
rect 15081 2283 15112 2287
rect 15137 2283 15145 2287
rect 15145 2283 15193 2287
rect 14321 2267 14377 2283
rect 14403 2267 14459 2283
rect 14485 2267 14541 2283
rect 14567 2267 14623 2283
rect 14649 2267 14705 2283
rect 14731 2267 14787 2283
rect 14813 2267 14869 2283
rect 14894 2267 14950 2283
rect 14975 2267 15031 2283
rect 15056 2267 15112 2283
rect 15137 2267 15193 2283
rect 14321 2231 14362 2267
rect 14362 2231 14375 2267
rect 14375 2231 14377 2267
rect 14403 2231 14427 2267
rect 14427 2231 14440 2267
rect 14440 2231 14459 2267
rect 14485 2231 14492 2267
rect 14492 2231 14505 2267
rect 14505 2231 14541 2267
rect 14567 2231 14569 2267
rect 14569 2231 14621 2267
rect 14621 2231 14623 2267
rect 14649 2231 14685 2267
rect 14685 2231 14697 2267
rect 14697 2231 14705 2267
rect 14731 2231 14749 2267
rect 14749 2231 14761 2267
rect 14761 2231 14787 2267
rect 14813 2231 14825 2267
rect 14825 2231 14869 2267
rect 14894 2231 14941 2267
rect 14941 2231 14950 2267
rect 14975 2231 15005 2267
rect 15005 2231 15017 2267
rect 15017 2231 15031 2267
rect 15056 2231 15069 2267
rect 15069 2231 15081 2267
rect 15081 2231 15112 2267
rect 15137 2231 15145 2267
rect 15145 2231 15193 2267
rect 14321 2199 14377 2203
rect 14403 2199 14459 2203
rect 14485 2199 14541 2203
rect 14567 2199 14623 2203
rect 14649 2199 14705 2203
rect 14731 2199 14787 2203
rect 14813 2199 14869 2203
rect 14894 2199 14950 2203
rect 14975 2199 15031 2203
rect 15056 2199 15112 2203
rect 15137 2199 15193 2203
rect 14321 2147 14362 2199
rect 14362 2147 14375 2199
rect 14375 2147 14377 2199
rect 14403 2147 14427 2199
rect 14427 2147 14440 2199
rect 14440 2147 14459 2199
rect 14485 2147 14492 2199
rect 14492 2147 14505 2199
rect 14505 2147 14541 2199
rect 14567 2147 14569 2199
rect 14569 2147 14621 2199
rect 14621 2147 14623 2199
rect 14649 2147 14685 2199
rect 14685 2147 14697 2199
rect 14697 2147 14705 2199
rect 14731 2147 14749 2199
rect 14749 2147 14761 2199
rect 14761 2147 14787 2199
rect 14813 2147 14825 2199
rect 14825 2147 14869 2199
rect 14894 2147 14941 2199
rect 14941 2147 14950 2199
rect 14975 2147 15005 2199
rect 15005 2147 15017 2199
rect 15017 2147 15031 2199
rect 15056 2147 15069 2199
rect 15069 2147 15081 2199
rect 15081 2147 15112 2199
rect 15137 2147 15145 2199
rect 15145 2147 15193 2199
rect 18243 2487 18291 2539
rect 18291 2487 18299 2539
rect 18324 2487 18355 2539
rect 18355 2487 18367 2539
rect 18367 2487 18380 2539
rect 18405 2487 18419 2539
rect 18419 2487 18431 2539
rect 18431 2487 18461 2539
rect 18486 2487 18495 2539
rect 18495 2487 18542 2539
rect 18567 2487 18611 2539
rect 18611 2487 18623 2539
rect 18649 2487 18675 2539
rect 18675 2487 18687 2539
rect 18687 2487 18705 2539
rect 18731 2487 18739 2539
rect 18739 2487 18751 2539
rect 18751 2487 18787 2539
rect 18813 2487 18815 2539
rect 18815 2487 18867 2539
rect 18867 2487 18869 2539
rect 18895 2487 18931 2539
rect 18931 2487 18944 2539
rect 18944 2487 18951 2539
rect 18977 2487 18996 2539
rect 18996 2487 19009 2539
rect 19009 2487 19033 2539
rect 19059 2487 19061 2539
rect 19061 2487 19074 2539
rect 19074 2487 19115 2539
rect 18243 2483 18299 2487
rect 18324 2483 18380 2487
rect 18405 2483 18461 2487
rect 18486 2483 18542 2487
rect 18567 2483 18623 2487
rect 18649 2483 18705 2487
rect 18731 2483 18787 2487
rect 18813 2483 18869 2487
rect 18895 2483 18951 2487
rect 18977 2483 19033 2487
rect 19059 2483 19115 2487
rect 18243 2419 18291 2455
rect 18291 2419 18299 2455
rect 18324 2419 18355 2455
rect 18355 2419 18367 2455
rect 18367 2419 18380 2455
rect 18405 2419 18419 2455
rect 18419 2419 18431 2455
rect 18431 2419 18461 2455
rect 18486 2419 18495 2455
rect 18495 2419 18542 2455
rect 18567 2419 18611 2455
rect 18611 2419 18623 2455
rect 18649 2419 18675 2455
rect 18675 2419 18687 2455
rect 18687 2419 18705 2455
rect 18731 2419 18739 2455
rect 18739 2419 18751 2455
rect 18751 2419 18787 2455
rect 18813 2419 18815 2455
rect 18815 2419 18867 2455
rect 18867 2419 18869 2455
rect 18895 2419 18931 2455
rect 18931 2419 18944 2455
rect 18944 2419 18951 2455
rect 18977 2419 18996 2455
rect 18996 2419 19009 2455
rect 19009 2419 19033 2455
rect 19059 2419 19061 2455
rect 19061 2419 19074 2455
rect 19074 2419 19115 2455
rect 18243 2403 18299 2419
rect 18324 2403 18380 2419
rect 18405 2403 18461 2419
rect 18486 2403 18542 2419
rect 18567 2403 18623 2419
rect 18649 2403 18705 2419
rect 18731 2403 18787 2419
rect 18813 2403 18869 2419
rect 18895 2403 18951 2419
rect 18977 2403 19033 2419
rect 19059 2403 19115 2419
rect 18243 2399 18291 2403
rect 18291 2399 18299 2403
rect 18324 2399 18355 2403
rect 18355 2399 18367 2403
rect 18367 2399 18380 2403
rect 18405 2399 18419 2403
rect 18419 2399 18431 2403
rect 18431 2399 18461 2403
rect 18486 2399 18495 2403
rect 18495 2399 18542 2403
rect 18243 2351 18291 2371
rect 18291 2351 18299 2371
rect 18324 2351 18355 2371
rect 18355 2351 18367 2371
rect 18367 2351 18380 2371
rect 18405 2351 18419 2371
rect 18419 2351 18431 2371
rect 18431 2351 18461 2371
rect 18486 2351 18495 2371
rect 18495 2351 18542 2371
rect 18567 2399 18611 2403
rect 18611 2399 18623 2403
rect 18649 2399 18675 2403
rect 18675 2399 18687 2403
rect 18687 2399 18705 2403
rect 18731 2399 18739 2403
rect 18739 2399 18751 2403
rect 18751 2399 18787 2403
rect 18813 2399 18815 2403
rect 18815 2399 18867 2403
rect 18867 2399 18869 2403
rect 18895 2399 18931 2403
rect 18931 2399 18944 2403
rect 18944 2399 18951 2403
rect 18977 2399 18996 2403
rect 18996 2399 19009 2403
rect 19009 2399 19033 2403
rect 19059 2399 19061 2403
rect 19061 2399 19074 2403
rect 19074 2399 19115 2403
rect 18567 2351 18611 2371
rect 18611 2351 18623 2371
rect 18649 2351 18675 2371
rect 18675 2351 18687 2371
rect 18687 2351 18705 2371
rect 18731 2351 18739 2371
rect 18739 2351 18751 2371
rect 18751 2351 18787 2371
rect 18813 2351 18815 2371
rect 18815 2351 18867 2371
rect 18867 2351 18869 2371
rect 18895 2351 18931 2371
rect 18931 2351 18944 2371
rect 18944 2351 18951 2371
rect 18977 2351 18996 2371
rect 18996 2351 19009 2371
rect 19009 2351 19033 2371
rect 19059 2351 19061 2371
rect 19061 2351 19074 2371
rect 19074 2351 19115 2371
rect 18243 2335 18299 2351
rect 18324 2335 18380 2351
rect 18405 2335 18461 2351
rect 18486 2335 18542 2351
rect 18567 2335 18623 2351
rect 18649 2335 18705 2351
rect 18731 2335 18787 2351
rect 18813 2335 18869 2351
rect 18895 2335 18951 2351
rect 18977 2335 19033 2351
rect 19059 2335 19115 2351
rect 18243 2315 18291 2335
rect 18291 2315 18299 2335
rect 18324 2315 18355 2335
rect 18355 2315 18367 2335
rect 18367 2315 18380 2335
rect 18405 2315 18419 2335
rect 18419 2315 18431 2335
rect 18431 2315 18461 2335
rect 18486 2315 18495 2335
rect 18495 2315 18542 2335
rect 18243 2283 18291 2287
rect 18291 2283 18299 2287
rect 18324 2283 18355 2287
rect 18355 2283 18367 2287
rect 18367 2283 18380 2287
rect 18405 2283 18419 2287
rect 18419 2283 18431 2287
rect 18431 2283 18461 2287
rect 18486 2283 18495 2287
rect 18495 2283 18542 2287
rect 18567 2315 18611 2335
rect 18611 2315 18623 2335
rect 18649 2315 18675 2335
rect 18675 2315 18687 2335
rect 18687 2315 18705 2335
rect 18731 2315 18739 2335
rect 18739 2315 18751 2335
rect 18751 2315 18787 2335
rect 18813 2315 18815 2335
rect 18815 2315 18867 2335
rect 18867 2315 18869 2335
rect 18895 2315 18931 2335
rect 18931 2315 18944 2335
rect 18944 2315 18951 2335
rect 18977 2315 18996 2335
rect 18996 2315 19009 2335
rect 19009 2315 19033 2335
rect 19059 2315 19061 2335
rect 19061 2315 19074 2335
rect 19074 2315 19115 2335
rect 18567 2283 18611 2287
rect 18611 2283 18623 2287
rect 18649 2283 18675 2287
rect 18675 2283 18687 2287
rect 18687 2283 18705 2287
rect 18731 2283 18739 2287
rect 18739 2283 18751 2287
rect 18751 2283 18787 2287
rect 18813 2283 18815 2287
rect 18815 2283 18867 2287
rect 18867 2283 18869 2287
rect 18895 2283 18931 2287
rect 18931 2283 18944 2287
rect 18944 2283 18951 2287
rect 18977 2283 18996 2287
rect 18996 2283 19009 2287
rect 19009 2283 19033 2287
rect 19059 2283 19061 2287
rect 19061 2283 19074 2287
rect 19074 2283 19115 2287
rect 18243 2267 18299 2283
rect 18324 2267 18380 2283
rect 18405 2267 18461 2283
rect 18486 2267 18542 2283
rect 18567 2267 18623 2283
rect 18649 2267 18705 2283
rect 18731 2267 18787 2283
rect 18813 2267 18869 2283
rect 18895 2267 18951 2283
rect 18977 2267 19033 2283
rect 19059 2267 19115 2283
rect 18243 2231 18291 2267
rect 18291 2231 18299 2267
rect 18324 2231 18355 2267
rect 18355 2231 18367 2267
rect 18367 2231 18380 2267
rect 18405 2231 18419 2267
rect 18419 2231 18431 2267
rect 18431 2231 18461 2267
rect 18486 2231 18495 2267
rect 18495 2231 18542 2267
rect 18567 2231 18611 2267
rect 18611 2231 18623 2267
rect 18649 2231 18675 2267
rect 18675 2231 18687 2267
rect 18687 2231 18705 2267
rect 18731 2231 18739 2267
rect 18739 2231 18751 2267
rect 18751 2231 18787 2267
rect 18813 2231 18815 2267
rect 18815 2231 18867 2267
rect 18867 2231 18869 2267
rect 18895 2231 18931 2267
rect 18931 2231 18944 2267
rect 18944 2231 18951 2267
rect 18977 2231 18996 2267
rect 18996 2231 19009 2267
rect 19009 2231 19033 2267
rect 19059 2231 19061 2267
rect 19061 2231 19074 2267
rect 19074 2231 19115 2267
rect 18243 2199 18299 2203
rect 18324 2199 18380 2203
rect 18405 2199 18461 2203
rect 18486 2199 18542 2203
rect 18567 2199 18623 2203
rect 18649 2199 18705 2203
rect 18731 2199 18787 2203
rect 18813 2199 18869 2203
rect 18895 2199 18951 2203
rect 18977 2199 19033 2203
rect 19059 2199 19115 2203
rect 18243 2147 18291 2199
rect 18291 2147 18299 2199
rect 18324 2147 18355 2199
rect 18355 2147 18367 2199
rect 18367 2147 18380 2199
rect 18405 2147 18419 2199
rect 18419 2147 18431 2199
rect 18431 2147 18461 2199
rect 18486 2147 18495 2199
rect 18495 2147 18542 2199
rect 18567 2147 18611 2199
rect 18611 2147 18623 2199
rect 18649 2147 18675 2199
rect 18675 2147 18687 2199
rect 18687 2147 18705 2199
rect 18731 2147 18739 2199
rect 18739 2147 18751 2199
rect 18751 2147 18787 2199
rect 18813 2147 18815 2199
rect 18815 2147 18867 2199
rect 18867 2147 18869 2199
rect 18895 2147 18931 2199
rect 18931 2147 18944 2199
rect 18944 2147 18951 2199
rect 18977 2147 18996 2199
rect 18996 2147 19009 2199
rect 19009 2147 19033 2199
rect 19059 2147 19061 2199
rect 19061 2147 19074 2199
rect 19074 2147 19115 2199
rect 962 1969 1011 2021
rect 1011 1969 1018 2021
rect 962 1965 1018 1969
rect 1043 1969 1095 2021
rect 1095 1969 1099 2021
rect 1043 1965 1099 1969
rect 1123 1969 1127 2021
rect 1127 1969 1179 2021
rect 1123 1965 1179 1969
rect 1203 1969 1210 2021
rect 1210 1969 1259 2021
rect 1203 1965 1259 1969
rect 962 1893 1018 1897
rect 962 1841 1011 1893
rect 1011 1841 1018 1893
rect 1043 1893 1099 1897
rect 1043 1841 1095 1893
rect 1095 1841 1099 1893
rect 1123 1893 1179 1897
rect 1123 1841 1127 1893
rect 1127 1841 1179 1893
rect 1203 1893 1259 1897
rect 1203 1841 1210 1893
rect 1210 1841 1259 1893
rect 6336 1969 6385 2021
rect 6385 1969 6392 2021
rect 6417 1969 6452 2021
rect 6452 1969 6467 2021
rect 6467 1969 6473 2021
rect 6498 1969 6519 2021
rect 6519 1969 6534 2021
rect 6534 1969 6554 2021
rect 6579 1969 6586 2021
rect 6586 1969 6601 2021
rect 6601 1969 6635 2021
rect 6661 1969 6668 2021
rect 6668 1969 6717 2021
rect 6336 1965 6392 1969
rect 6417 1965 6473 1969
rect 6498 1965 6554 1969
rect 6579 1965 6635 1969
rect 6661 1965 6717 1969
rect 6336 1893 6392 1897
rect 6417 1893 6473 1897
rect 6498 1893 6554 1897
rect 6579 1893 6635 1897
rect 6661 1893 6717 1897
rect 6336 1841 6385 1893
rect 6385 1841 6392 1893
rect 6417 1841 6452 1893
rect 6452 1841 6467 1893
rect 6467 1841 6473 1893
rect 6498 1841 6519 1893
rect 6519 1841 6534 1893
rect 6534 1841 6554 1893
rect 6579 1841 6586 1893
rect 6586 1841 6601 1893
rect 6601 1841 6635 1893
rect 6661 1841 6668 1893
rect 6668 1841 6717 1893
rect 7267 1969 7316 2021
rect 7316 1969 7323 2021
rect 7349 1969 7383 2021
rect 7383 1969 7398 2021
rect 7398 1969 7405 2021
rect 7430 1969 7450 2021
rect 7450 1969 7465 2021
rect 7465 1969 7486 2021
rect 7511 1969 7517 2021
rect 7517 1969 7532 2021
rect 7532 1969 7567 2021
rect 7592 1969 7599 2021
rect 7599 1969 7648 2021
rect 7267 1965 7323 1969
rect 7349 1965 7405 1969
rect 7430 1965 7486 1969
rect 7511 1965 7567 1969
rect 7592 1965 7648 1969
rect 7267 1893 7323 1897
rect 7349 1893 7405 1897
rect 7430 1893 7486 1897
rect 7511 1893 7567 1897
rect 7592 1893 7648 1897
rect 7267 1841 7316 1893
rect 7316 1841 7323 1893
rect 7349 1841 7383 1893
rect 7383 1841 7398 1893
rect 7398 1841 7405 1893
rect 7430 1841 7450 1893
rect 7450 1841 7465 1893
rect 7465 1841 7486 1893
rect 7511 1841 7517 1893
rect 7517 1841 7532 1893
rect 7532 1841 7567 1893
rect 7592 1841 7599 1893
rect 7599 1841 7648 1893
rect 12820 1969 12869 2021
rect 12869 1969 12876 2021
rect 12901 1969 12936 2021
rect 12936 1969 12951 2021
rect 12951 1969 12957 2021
rect 12982 1969 13003 2021
rect 13003 1969 13018 2021
rect 13018 1969 13038 2021
rect 13063 1969 13070 2021
rect 13070 1969 13085 2021
rect 13085 1969 13119 2021
rect 13145 1969 13152 2021
rect 13152 1969 13201 2021
rect 12820 1965 12876 1969
rect 12901 1965 12957 1969
rect 12982 1965 13038 1969
rect 13063 1965 13119 1969
rect 13145 1965 13201 1969
rect 12820 1893 12876 1897
rect 12901 1893 12957 1897
rect 12982 1893 13038 1897
rect 13063 1893 13119 1897
rect 13145 1893 13201 1897
rect 12820 1841 12869 1893
rect 12869 1841 12876 1893
rect 12901 1841 12936 1893
rect 12936 1841 12951 1893
rect 12951 1841 12957 1893
rect 12982 1841 13003 1893
rect 13003 1841 13018 1893
rect 13018 1841 13038 1893
rect 13063 1841 13070 1893
rect 13070 1841 13085 1893
rect 13085 1841 13119 1893
rect 13145 1841 13152 1893
rect 13152 1841 13201 1893
rect 13751 1969 13800 2021
rect 13800 1969 13807 2021
rect 13833 1969 13867 2021
rect 13867 1969 13882 2021
rect 13882 1969 13889 2021
rect 13914 1969 13934 2021
rect 13934 1969 13949 2021
rect 13949 1969 13970 2021
rect 13995 1969 14001 2021
rect 14001 1969 14016 2021
rect 14016 1969 14051 2021
rect 14076 1969 14083 2021
rect 14083 1969 14132 2021
rect 13751 1965 13807 1969
rect 13833 1965 13889 1969
rect 13914 1965 13970 1969
rect 13995 1965 14051 1969
rect 14076 1965 14132 1969
rect 13751 1893 13807 1897
rect 13833 1893 13889 1897
rect 13914 1893 13970 1897
rect 13995 1893 14051 1897
rect 14076 1893 14132 1897
rect 13751 1841 13800 1893
rect 13800 1841 13807 1893
rect 13833 1841 13867 1893
rect 13867 1841 13882 1893
rect 13882 1841 13889 1893
rect 13914 1841 13934 1893
rect 13934 1841 13949 1893
rect 13949 1841 13970 1893
rect 13995 1841 14001 1893
rect 14001 1841 14016 1893
rect 14016 1841 14051 1893
rect 14076 1841 14083 1893
rect 14083 1841 14132 1893
rect 19389 1969 19438 2021
rect 19438 1969 19445 2021
rect 19389 1965 19445 1969
rect 19469 1969 19521 2021
rect 19521 1969 19525 2021
rect 19469 1965 19525 1969
rect 19549 1969 19552 2021
rect 19552 1969 19604 2021
rect 19604 1969 19605 2021
rect 19549 1965 19605 1969
rect 19629 1969 19636 2021
rect 19636 1969 19685 2021
rect 19629 1965 19685 1969
rect 19389 1893 19445 1897
rect 19389 1841 19438 1893
rect 19438 1841 19445 1893
rect 19469 1893 19525 1897
rect 19469 1841 19521 1893
rect 19521 1841 19525 1893
rect 19549 1893 19605 1897
rect 19549 1841 19552 1893
rect 19552 1841 19604 1893
rect 19604 1841 19605 1893
rect 19629 1893 19685 1897
rect 19629 1841 19636 1893
rect 19636 1841 19685 1893
rect 966 -109 1022 -53
rect 1085 -109 1141 -53
rect 1203 -109 1259 -53
rect 966 -193 1022 -137
rect 1085 -193 1141 -137
rect 1203 -193 1259 -137
rect 6336 -109 6392 -53
rect 6418 -109 6474 -53
rect 6499 -109 6555 -53
rect 6580 -109 6636 -53
rect 6661 -109 6717 -53
rect 6336 -179 6385 -137
rect 6385 -179 6392 -137
rect 6418 -179 6452 -137
rect 6452 -179 6467 -137
rect 6467 -179 6474 -137
rect 6499 -179 6519 -137
rect 6519 -179 6534 -137
rect 6534 -179 6555 -137
rect 6580 -179 6586 -137
rect 6586 -179 6601 -137
rect 6601 -179 6636 -137
rect 6661 -179 6668 -137
rect 6668 -179 6717 -137
rect 6336 -193 6392 -179
rect 6418 -193 6474 -179
rect 6499 -193 6555 -179
rect 6580 -193 6636 -179
rect 6661 -193 6717 -179
rect 7267 -109 7323 -53
rect 7349 -109 7405 -53
rect 7430 -109 7486 -53
rect 7511 -109 7567 -53
rect 7592 -109 7648 -53
rect 7267 -179 7316 -137
rect 7316 -179 7323 -137
rect 7349 -179 7383 -137
rect 7383 -179 7398 -137
rect 7398 -179 7405 -137
rect 7430 -179 7450 -137
rect 7450 -179 7465 -137
rect 7465 -179 7486 -137
rect 7511 -179 7517 -137
rect 7517 -179 7532 -137
rect 7532 -179 7567 -137
rect 7592 -179 7599 -137
rect 7599 -179 7648 -137
rect 7267 -193 7323 -179
rect 7349 -193 7405 -179
rect 7430 -193 7486 -179
rect 7511 -193 7567 -179
rect 7592 -193 7648 -179
rect 12820 -109 12876 -53
rect 12902 -109 12958 -53
rect 12983 -109 13039 -53
rect 13064 -109 13120 -53
rect 13145 -109 13201 -53
rect 12820 -178 12869 -137
rect 12869 -178 12876 -137
rect 12902 -178 12936 -137
rect 12936 -178 12951 -137
rect 12951 -178 12958 -137
rect 12983 -178 13003 -137
rect 13003 -178 13018 -137
rect 13018 -178 13039 -137
rect 13064 -178 13070 -137
rect 13070 -178 13085 -137
rect 13085 -178 13120 -137
rect 13145 -178 13152 -137
rect 13152 -178 13201 -137
rect 12820 -193 12876 -178
rect 12902 -193 12958 -178
rect 12983 -193 13039 -178
rect 13064 -193 13120 -178
rect 13145 -193 13201 -178
rect 13751 -109 13807 -53
rect 13833 -109 13889 -53
rect 13914 -109 13970 -53
rect 13995 -109 14051 -53
rect 14076 -109 14132 -53
rect 13751 -179 13800 -137
rect 13800 -179 13807 -137
rect 13833 -179 13867 -137
rect 13867 -179 13882 -137
rect 13882 -179 13889 -137
rect 13914 -179 13934 -137
rect 13934 -179 13949 -137
rect 13949 -179 13970 -137
rect 13995 -179 14001 -137
rect 14001 -179 14016 -137
rect 14016 -179 14051 -137
rect 14076 -179 14083 -137
rect 14083 -179 14132 -137
rect 13751 -193 13807 -179
rect 13833 -193 13889 -179
rect 13914 -193 13970 -179
rect 13995 -193 14051 -179
rect 14076 -193 14132 -179
rect 19389 -109 19445 -53
rect 19469 -109 19525 -53
rect 19549 -109 19605 -53
rect 19629 -109 19685 -53
rect 19389 -179 19438 -137
rect 19438 -179 19445 -137
rect 19389 -193 19445 -179
rect 19469 -179 19470 -137
rect 19470 -179 19522 -137
rect 19522 -179 19525 -137
rect 19469 -193 19525 -179
rect 19549 -179 19553 -137
rect 19553 -179 19605 -137
rect 19549 -193 19605 -179
rect 19629 -179 19636 -137
rect 19636 -179 19685 -137
rect 19629 -193 19685 -179
rect 6337 -1595 6386 -1565
rect 6386 -1595 6393 -1565
rect 6443 -1595 6452 -1565
rect 6452 -1595 6466 -1565
rect 6466 -1595 6499 -1565
rect 6549 -1595 6584 -1565
rect 6584 -1595 6597 -1565
rect 6597 -1595 6605 -1565
rect 6655 -1595 6662 -1565
rect 6662 -1595 6711 -1565
rect 6337 -1607 6393 -1595
rect 6443 -1607 6499 -1595
rect 6549 -1607 6605 -1595
rect 6655 -1607 6711 -1595
rect 6337 -1621 6386 -1607
rect 6386 -1621 6393 -1607
rect 6443 -1621 6452 -1607
rect 6452 -1621 6466 -1607
rect 6466 -1621 6499 -1607
rect 6337 -1659 6386 -1645
rect 6386 -1659 6393 -1645
rect 6443 -1659 6452 -1645
rect 6452 -1659 6466 -1645
rect 6466 -1659 6499 -1645
rect 6549 -1621 6584 -1607
rect 6584 -1621 6597 -1607
rect 6597 -1621 6605 -1607
rect 6655 -1621 6662 -1607
rect 6662 -1621 6711 -1607
rect 6549 -1659 6584 -1645
rect 6584 -1659 6597 -1645
rect 6597 -1659 6605 -1645
rect 6655 -1659 6662 -1645
rect 6662 -1659 6711 -1645
rect 6337 -1671 6393 -1659
rect 6443 -1671 6499 -1659
rect 6549 -1671 6605 -1659
rect 6655 -1671 6711 -1659
rect 6337 -1701 6386 -1671
rect 6386 -1701 6393 -1671
rect 6443 -1701 6452 -1671
rect 6452 -1701 6466 -1671
rect 6466 -1701 6499 -1671
rect 6549 -1701 6584 -1671
rect 6584 -1701 6597 -1671
rect 6597 -1701 6605 -1671
rect 6655 -1701 6662 -1671
rect 6662 -1701 6711 -1671
rect 7269 -1595 7318 -1565
rect 7318 -1595 7325 -1565
rect 7375 -1595 7384 -1565
rect 7384 -1595 7398 -1565
rect 7398 -1595 7431 -1565
rect 7481 -1595 7516 -1565
rect 7516 -1595 7529 -1565
rect 7529 -1595 7537 -1565
rect 7587 -1595 7594 -1565
rect 7594 -1595 7643 -1565
rect 7269 -1607 7325 -1595
rect 7375 -1607 7431 -1595
rect 7481 -1607 7537 -1595
rect 7587 -1607 7643 -1595
rect 7269 -1621 7318 -1607
rect 7318 -1621 7325 -1607
rect 7375 -1621 7384 -1607
rect 7384 -1621 7398 -1607
rect 7398 -1621 7431 -1607
rect 7269 -1659 7318 -1645
rect 7318 -1659 7325 -1645
rect 7375 -1659 7384 -1645
rect 7384 -1659 7398 -1645
rect 7398 -1659 7431 -1645
rect 7481 -1621 7516 -1607
rect 7516 -1621 7529 -1607
rect 7529 -1621 7537 -1607
rect 7587 -1621 7594 -1607
rect 7594 -1621 7643 -1607
rect 7481 -1659 7516 -1645
rect 7516 -1659 7529 -1645
rect 7529 -1659 7537 -1645
rect 7587 -1659 7594 -1645
rect 7594 -1659 7643 -1645
rect 7269 -1671 7325 -1659
rect 7375 -1671 7431 -1659
rect 7481 -1671 7537 -1659
rect 7587 -1671 7643 -1659
rect 7269 -1701 7318 -1671
rect 7318 -1701 7325 -1671
rect 7375 -1701 7384 -1671
rect 7384 -1701 7398 -1671
rect 7398 -1701 7431 -1671
rect 7481 -1701 7516 -1671
rect 7516 -1701 7529 -1671
rect 7529 -1701 7537 -1671
rect 7587 -1701 7594 -1671
rect 7594 -1701 7643 -1671
rect 12822 -1595 12871 -1565
rect 12871 -1595 12878 -1565
rect 12903 -1595 12937 -1565
rect 12937 -1595 12951 -1565
rect 12951 -1595 12959 -1565
rect 12984 -1595 13003 -1565
rect 13003 -1595 13017 -1565
rect 13017 -1595 13069 -1565
rect 13069 -1595 13082 -1565
rect 13082 -1595 13134 -1565
rect 13134 -1595 13147 -1565
rect 13147 -1595 13199 -1565
rect 13199 -1595 13200 -1565
rect 12822 -1607 12878 -1595
rect 12903 -1607 12959 -1595
rect 12984 -1607 13200 -1595
rect 12822 -1621 12871 -1607
rect 12871 -1621 12878 -1607
rect 12903 -1621 12937 -1607
rect 12937 -1621 12951 -1607
rect 12951 -1621 12959 -1607
rect 12822 -1659 12871 -1645
rect 12871 -1659 12878 -1645
rect 12903 -1659 12937 -1645
rect 12937 -1659 12951 -1645
rect 12951 -1659 12959 -1645
rect 12984 -1659 13003 -1607
rect 13003 -1659 13017 -1607
rect 13017 -1659 13069 -1607
rect 13069 -1659 13082 -1607
rect 13082 -1659 13134 -1607
rect 13134 -1659 13147 -1607
rect 13147 -1659 13199 -1607
rect 13199 -1659 13200 -1607
rect 12822 -1671 12878 -1659
rect 12903 -1671 12959 -1659
rect 12984 -1671 13200 -1659
rect 12822 -1701 12871 -1671
rect 12871 -1701 12878 -1671
rect 12903 -1701 12937 -1671
rect 12937 -1701 12951 -1671
rect 12951 -1701 12959 -1671
rect 12984 -1701 13003 -1671
rect 13003 -1701 13017 -1671
rect 13017 -1701 13069 -1671
rect 13069 -1701 13082 -1671
rect 13082 -1701 13134 -1671
rect 13134 -1701 13147 -1671
rect 13147 -1701 13199 -1671
rect 13199 -1701 13200 -1671
rect 13753 -1595 13802 -1565
rect 13802 -1595 13809 -1565
rect 13834 -1595 13868 -1565
rect 13868 -1595 13882 -1565
rect 13882 -1595 13890 -1565
rect 13915 -1595 13934 -1565
rect 13934 -1595 13948 -1565
rect 13948 -1595 14000 -1565
rect 14000 -1595 14013 -1565
rect 14013 -1595 14065 -1565
rect 14065 -1595 14078 -1565
rect 14078 -1595 14130 -1565
rect 14130 -1595 14131 -1565
rect 13753 -1607 13809 -1595
rect 13834 -1607 13890 -1595
rect 13915 -1607 14131 -1595
rect 13753 -1621 13802 -1607
rect 13802 -1621 13809 -1607
rect 13834 -1621 13868 -1607
rect 13868 -1621 13882 -1607
rect 13882 -1621 13890 -1607
rect 13753 -1659 13802 -1645
rect 13802 -1659 13809 -1645
rect 13834 -1659 13868 -1645
rect 13868 -1659 13882 -1645
rect 13882 -1659 13890 -1645
rect 13915 -1659 13934 -1607
rect 13934 -1659 13948 -1607
rect 13948 -1659 14000 -1607
rect 14000 -1659 14013 -1607
rect 14013 -1659 14065 -1607
rect 14065 -1659 14078 -1607
rect 14078 -1659 14130 -1607
rect 14130 -1659 14131 -1607
rect 13753 -1671 13809 -1659
rect 13834 -1671 13890 -1659
rect 13915 -1671 14131 -1659
rect 13753 -1701 13802 -1671
rect 13802 -1701 13809 -1671
rect 13834 -1701 13868 -1671
rect 13868 -1701 13882 -1671
rect 13882 -1701 13890 -1671
rect 13915 -1701 13934 -1671
rect 13934 -1701 13948 -1671
rect 13948 -1701 14000 -1671
rect 14000 -1701 14013 -1671
rect 14013 -1701 14065 -1671
rect 14065 -1701 14078 -1671
rect 14078 -1701 14130 -1671
rect 14130 -1701 14131 -1671
rect 19385 -1595 19421 -1565
rect 19421 -1595 19435 -1565
rect 19435 -1595 19441 -1565
rect 19466 -1595 19487 -1565
rect 19487 -1595 19501 -1565
rect 19501 -1595 19522 -1565
rect 19547 -1595 19553 -1565
rect 19553 -1595 19566 -1565
rect 19566 -1595 19603 -1565
rect 19628 -1595 19631 -1565
rect 19631 -1595 19683 -1565
rect 19683 -1595 19684 -1565
rect 19385 -1607 19441 -1595
rect 19466 -1607 19522 -1595
rect 19547 -1607 19603 -1595
rect 19628 -1607 19684 -1595
rect 19385 -1621 19421 -1607
rect 19421 -1621 19435 -1607
rect 19435 -1621 19441 -1607
rect 19466 -1621 19487 -1607
rect 19487 -1621 19501 -1607
rect 19501 -1621 19522 -1607
rect 19547 -1621 19553 -1607
rect 19553 -1621 19566 -1607
rect 19566 -1621 19603 -1607
rect 19628 -1621 19631 -1607
rect 19631 -1621 19683 -1607
rect 19683 -1621 19684 -1607
rect 19385 -1659 19421 -1645
rect 19421 -1659 19435 -1645
rect 19435 -1659 19441 -1645
rect 19466 -1659 19487 -1645
rect 19487 -1659 19501 -1645
rect 19501 -1659 19522 -1645
rect 19547 -1659 19553 -1645
rect 19553 -1659 19566 -1645
rect 19566 -1659 19603 -1645
rect 19628 -1659 19631 -1645
rect 19631 -1659 19683 -1645
rect 19683 -1659 19684 -1645
rect 19385 -1671 19441 -1659
rect 19466 -1671 19522 -1659
rect 19547 -1671 19603 -1659
rect 19628 -1671 19684 -1659
rect 19385 -1701 19421 -1671
rect 19421 -1701 19435 -1671
rect 19435 -1701 19441 -1671
rect 19466 -1701 19487 -1671
rect 19487 -1701 19501 -1671
rect 19501 -1701 19522 -1671
rect 19547 -1701 19553 -1671
rect 19553 -1701 19566 -1671
rect 19566 -1701 19603 -1671
rect 19628 -1701 19631 -1671
rect 19631 -1701 19683 -1671
rect 19683 -1701 19684 -1671
<< metal3 >>
rect 957 4453 1268 4478
rect 957 4397 962 4453
rect 1018 4397 1044 4453
rect 1100 4397 1126 4453
rect 1182 4397 1207 4453
rect 1263 4397 1268 4453
rect 957 4369 1268 4397
rect 957 4313 962 4369
rect 1018 4313 1044 4369
rect 1100 4313 1126 4369
rect 1182 4313 1207 4369
rect 1263 4313 1268 4369
rect 957 3065 1268 4313
rect 957 3009 962 3065
rect 1018 3009 1043 3065
rect 1099 3009 1123 3065
rect 1179 3009 1203 3065
rect 1259 3009 1268 3065
rect 957 2981 1268 3009
rect 957 2925 962 2981
rect 1018 2925 1043 2981
rect 1099 2925 1123 2981
rect 1179 2925 1203 2981
rect 1259 2925 1268 2981
rect 957 2840 1268 2925
rect 957 2784 962 2840
rect 1018 2784 1043 2840
rect 1099 2784 1123 2840
rect 1179 2784 1203 2840
rect 1259 2784 1268 2840
rect 957 2716 1268 2784
rect 957 2660 962 2716
rect 1018 2660 1043 2716
rect 1099 2660 1123 2716
rect 1179 2660 1203 2716
rect 1259 2660 1268 2716
rect 957 2021 1268 2660
rect 6327 4453 6726 4469
rect 6327 4397 6336 4453
rect 6392 4397 6418 4453
rect 6474 4397 6499 4453
rect 6555 4397 6580 4453
rect 6636 4397 6661 4453
rect 6717 4397 6726 4453
rect 6327 4369 6726 4397
rect 6327 4313 6336 4369
rect 6392 4313 6418 4369
rect 6474 4313 6499 4369
rect 6555 4313 6580 4369
rect 6636 4313 6661 4369
rect 6717 4313 6726 4369
rect 6327 3065 6726 4313
rect 6327 3009 6336 3065
rect 6392 3009 6418 3065
rect 6474 3009 6499 3065
rect 6555 3009 6580 3065
rect 6636 3009 6661 3065
rect 6717 3009 6726 3065
rect 6327 2981 6726 3009
rect 6327 2925 6336 2981
rect 6392 2925 6418 2981
rect 6474 2925 6499 2981
rect 6555 2925 6580 2981
rect 6636 2925 6661 2981
rect 6717 2925 6726 2981
rect 6327 2840 6726 2925
rect 6327 2784 6336 2840
rect 6392 2784 6417 2840
rect 6473 2784 6498 2840
rect 6554 2784 6579 2840
rect 6635 2784 6661 2840
rect 6717 2784 6726 2840
rect 6327 2716 6726 2784
rect 6327 2660 6336 2716
rect 6392 2660 6417 2716
rect 6473 2660 6498 2716
rect 6554 2660 6579 2716
rect 6635 2660 6661 2716
rect 6717 2660 6726 2716
rect 1348 2539 2230 2546
rect 1348 2483 1353 2539
rect 1409 2483 1435 2539
rect 1491 2483 1517 2539
rect 1573 2483 1599 2539
rect 1655 2483 1681 2539
rect 1737 2483 1763 2539
rect 1819 2483 1845 2539
rect 1901 2483 1926 2539
rect 1982 2483 2007 2539
rect 2063 2483 2088 2539
rect 2144 2483 2169 2539
rect 2225 2483 2230 2539
rect 1348 2455 2230 2483
rect 1348 2399 1353 2455
rect 1409 2399 1435 2455
rect 1491 2399 1517 2455
rect 1573 2399 1599 2455
rect 1655 2399 1681 2455
rect 1737 2399 1763 2455
rect 1819 2399 1845 2455
rect 1901 2399 1926 2455
rect 1982 2399 2007 2455
rect 2063 2399 2088 2455
rect 2144 2399 2169 2455
rect 2225 2399 2230 2455
rect 1348 2371 2230 2399
rect 1348 2315 1353 2371
rect 1409 2315 1435 2371
rect 1491 2315 1517 2371
rect 1573 2315 1599 2371
rect 1655 2315 1681 2371
rect 1737 2315 1763 2371
rect 1819 2315 1845 2371
rect 1901 2315 1926 2371
rect 1982 2315 2007 2371
rect 2063 2315 2088 2371
rect 2144 2315 2169 2371
rect 2225 2315 2230 2371
rect 1348 2287 2230 2315
rect 1348 2231 1353 2287
rect 1409 2231 1435 2287
rect 1491 2231 1517 2287
rect 1573 2231 1599 2287
rect 1655 2231 1681 2287
rect 1737 2231 1763 2287
rect 1819 2231 1845 2287
rect 1901 2231 1926 2287
rect 1982 2231 2007 2287
rect 2063 2231 2088 2287
rect 2144 2231 2169 2287
rect 2225 2231 2230 2287
rect 1348 2203 2230 2231
rect 1348 2147 1353 2203
rect 1409 2147 1435 2203
rect 1491 2147 1517 2203
rect 1573 2147 1599 2203
rect 1655 2147 1681 2203
rect 1737 2147 1763 2203
rect 1819 2147 1845 2203
rect 1901 2147 1926 2203
rect 1982 2147 2007 2203
rect 2063 2147 2088 2203
rect 2144 2147 2169 2203
rect 2225 2147 2230 2203
rect 1348 2140 2230 2147
rect 5270 2539 6152 2546
rect 5270 2483 5275 2539
rect 5331 2483 5356 2539
rect 5412 2483 5437 2539
rect 5493 2483 5518 2539
rect 5574 2483 5599 2539
rect 5655 2483 5681 2539
rect 5737 2483 5763 2539
rect 5819 2483 5845 2539
rect 5901 2483 5927 2539
rect 5983 2483 6009 2539
rect 6065 2483 6091 2539
rect 6147 2483 6152 2539
rect 5270 2455 6152 2483
rect 5270 2399 5275 2455
rect 5331 2399 5356 2455
rect 5412 2399 5437 2455
rect 5493 2399 5518 2455
rect 5574 2399 5599 2455
rect 5655 2399 5681 2455
rect 5737 2399 5763 2455
rect 5819 2399 5845 2455
rect 5901 2399 5927 2455
rect 5983 2399 6009 2455
rect 6065 2399 6091 2455
rect 6147 2399 6152 2455
rect 5270 2371 6152 2399
rect 5270 2315 5275 2371
rect 5331 2315 5356 2371
rect 5412 2315 5437 2371
rect 5493 2315 5518 2371
rect 5574 2315 5599 2371
rect 5655 2315 5681 2371
rect 5737 2315 5763 2371
rect 5819 2315 5845 2371
rect 5901 2315 5927 2371
rect 5983 2315 6009 2371
rect 6065 2315 6091 2371
rect 6147 2315 6152 2371
rect 5270 2287 6152 2315
rect 5270 2231 5275 2287
rect 5331 2231 5356 2287
rect 5412 2231 5437 2287
rect 5493 2231 5518 2287
rect 5574 2231 5599 2287
rect 5655 2231 5681 2287
rect 5737 2231 5763 2287
rect 5819 2231 5845 2287
rect 5901 2231 5927 2287
rect 5983 2231 6009 2287
rect 6065 2231 6091 2287
rect 6147 2231 6152 2287
rect 5270 2203 6152 2231
rect 5270 2147 5275 2203
rect 5331 2147 5356 2203
rect 5412 2147 5437 2203
rect 5493 2147 5518 2203
rect 5574 2147 5599 2203
rect 5655 2147 5681 2203
rect 5737 2147 5763 2203
rect 5819 2147 5845 2203
rect 5901 2147 5927 2203
rect 5983 2147 6009 2203
rect 6065 2147 6091 2203
rect 6147 2147 6152 2203
rect 5270 2140 6152 2147
rect 957 1965 962 2021
rect 1018 1965 1043 2021
rect 1099 1965 1123 2021
rect 1179 1965 1203 2021
rect 1259 1965 1268 2021
rect 957 1897 1268 1965
rect 957 1841 962 1897
rect 1018 1841 1043 1897
rect 1099 1841 1123 1897
rect 1179 1841 1203 1897
rect 1259 1841 1268 1897
rect 957 -53 1268 1841
rect 957 -109 966 -53
rect 1022 -109 1085 -53
rect 1141 -109 1203 -53
rect 1259 -109 1268 -53
rect 957 -137 1268 -109
rect 957 -193 966 -137
rect 1022 -193 1085 -137
rect 1141 -193 1203 -137
rect 1259 -193 1268 -137
rect 957 -1683 1268 -193
rect 6327 2021 6726 2660
rect 6327 1965 6336 2021
rect 6392 1965 6417 2021
rect 6473 1965 6498 2021
rect 6554 1965 6579 2021
rect 6635 1965 6661 2021
rect 6717 1965 6726 2021
rect 6327 1897 6726 1965
rect 6327 1841 6336 1897
rect 6392 1841 6417 1897
rect 6473 1841 6498 1897
rect 6554 1841 6579 1897
rect 6635 1841 6661 1897
rect 6717 1841 6726 1897
rect 6327 -53 6726 1841
rect 6327 -109 6336 -53
rect 6392 -109 6418 -53
rect 6474 -109 6499 -53
rect 6555 -109 6580 -53
rect 6636 -109 6661 -53
rect 6717 -109 6726 -53
rect 6327 -137 6726 -109
rect 6327 -193 6336 -137
rect 6392 -193 6418 -137
rect 6474 -193 6499 -137
rect 6555 -193 6580 -137
rect 6636 -193 6661 -137
rect 6717 -193 6726 -137
rect 6327 -1565 6726 -193
rect 6327 -1621 6337 -1565
rect 6393 -1621 6443 -1565
rect 6499 -1621 6549 -1565
rect 6605 -1621 6655 -1565
rect 6711 -1621 6726 -1565
rect 6327 -1645 6726 -1621
rect 6327 -1701 6337 -1645
rect 6393 -1701 6443 -1645
rect 6499 -1701 6549 -1645
rect 6605 -1701 6655 -1645
rect 6711 -1701 6726 -1645
rect 6327 -1723 6726 -1701
rect 7258 4453 7657 4469
rect 7258 4397 7267 4453
rect 7323 4397 7349 4453
rect 7405 4397 7430 4453
rect 7486 4397 7511 4453
rect 7567 4397 7592 4453
rect 7648 4397 7657 4453
rect 7258 4369 7657 4397
rect 7258 4313 7267 4369
rect 7323 4313 7349 4369
rect 7405 4313 7430 4369
rect 7486 4313 7511 4369
rect 7567 4313 7592 4369
rect 7648 4313 7657 4369
rect 7258 3065 7657 4313
rect 7258 3009 7267 3065
rect 7323 3009 7349 3065
rect 7405 3009 7430 3065
rect 7486 3009 7511 3065
rect 7567 3009 7592 3065
rect 7648 3009 7657 3065
rect 7258 2981 7657 3009
rect 7258 2925 7267 2981
rect 7323 2925 7349 2981
rect 7405 2925 7430 2981
rect 7486 2925 7511 2981
rect 7567 2925 7592 2981
rect 7648 2925 7657 2981
rect 7258 2840 7657 2925
rect 7258 2784 7267 2840
rect 7323 2784 7349 2840
rect 7405 2784 7430 2840
rect 7486 2784 7511 2840
rect 7567 2784 7592 2840
rect 7648 2784 7657 2840
rect 7258 2716 7657 2784
rect 7258 2660 7267 2716
rect 7323 2660 7349 2716
rect 7405 2660 7430 2716
rect 7486 2660 7511 2716
rect 7567 2660 7592 2716
rect 7648 2660 7657 2716
rect 7258 2021 7657 2660
rect 12811 4453 13210 4469
rect 12811 4397 12820 4453
rect 12876 4397 12902 4453
rect 12958 4397 12983 4453
rect 13039 4397 13064 4453
rect 13120 4397 13145 4453
rect 13201 4397 13210 4453
rect 12811 4369 13210 4397
rect 12811 4313 12820 4369
rect 12876 4313 12902 4369
rect 12958 4313 12983 4369
rect 13039 4313 13064 4369
rect 13120 4313 13145 4369
rect 13201 4313 13210 4369
rect 12811 3065 13210 4313
rect 12811 3009 12820 3065
rect 12876 3009 12902 3065
rect 12958 3009 12983 3065
rect 13039 3009 13064 3065
rect 13120 3009 13145 3065
rect 13201 3009 13210 3065
rect 12811 2981 13210 3009
rect 12811 2925 12820 2981
rect 12876 2925 12902 2981
rect 12958 2925 12983 2981
rect 13039 2925 13064 2981
rect 13120 2925 13145 2981
rect 13201 2925 13210 2981
rect 12811 2840 13210 2925
rect 12811 2784 12820 2840
rect 12876 2784 12901 2840
rect 12957 2784 12982 2840
rect 13038 2784 13063 2840
rect 13119 2784 13145 2840
rect 13201 2784 13210 2840
rect 12811 2716 13210 2784
rect 12811 2660 12820 2716
rect 12876 2660 12901 2716
rect 12957 2660 12982 2716
rect 13038 2660 13063 2716
rect 13119 2660 13145 2716
rect 13201 2660 13210 2716
rect 7832 2539 8714 2546
rect 7832 2483 7837 2539
rect 7893 2483 7919 2539
rect 7975 2483 8001 2539
rect 8057 2483 8083 2539
rect 8139 2483 8165 2539
rect 8221 2483 8247 2539
rect 8303 2483 8329 2539
rect 8385 2483 8410 2539
rect 8466 2483 8491 2539
rect 8547 2483 8572 2539
rect 8628 2483 8653 2539
rect 8709 2483 8714 2539
rect 7832 2455 8714 2483
rect 7832 2399 7837 2455
rect 7893 2399 7919 2455
rect 7975 2399 8001 2455
rect 8057 2399 8083 2455
rect 8139 2399 8165 2455
rect 8221 2399 8247 2455
rect 8303 2399 8329 2455
rect 8385 2399 8410 2455
rect 8466 2399 8491 2455
rect 8547 2399 8572 2455
rect 8628 2399 8653 2455
rect 8709 2399 8714 2455
rect 7832 2371 8714 2399
rect 7832 2315 7837 2371
rect 7893 2315 7919 2371
rect 7975 2315 8001 2371
rect 8057 2315 8083 2371
rect 8139 2315 8165 2371
rect 8221 2315 8247 2371
rect 8303 2315 8329 2371
rect 8385 2315 8410 2371
rect 8466 2315 8491 2371
rect 8547 2315 8572 2371
rect 8628 2315 8653 2371
rect 8709 2315 8714 2371
rect 7832 2287 8714 2315
rect 7832 2231 7837 2287
rect 7893 2231 7919 2287
rect 7975 2231 8001 2287
rect 8057 2231 8083 2287
rect 8139 2231 8165 2287
rect 8221 2231 8247 2287
rect 8303 2231 8329 2287
rect 8385 2231 8410 2287
rect 8466 2231 8491 2287
rect 8547 2231 8572 2287
rect 8628 2231 8653 2287
rect 8709 2231 8714 2287
rect 7832 2203 8714 2231
rect 7832 2147 7837 2203
rect 7893 2147 7919 2203
rect 7975 2147 8001 2203
rect 8057 2147 8083 2203
rect 8139 2147 8165 2203
rect 8221 2147 8247 2203
rect 8303 2147 8329 2203
rect 8385 2147 8410 2203
rect 8466 2147 8491 2203
rect 8547 2147 8572 2203
rect 8628 2147 8653 2203
rect 8709 2147 8714 2203
rect 7832 2140 8714 2147
rect 11754 2539 12636 2546
rect 11754 2483 11759 2539
rect 11815 2483 11840 2539
rect 11896 2483 11921 2539
rect 11977 2483 12002 2539
rect 12058 2483 12083 2539
rect 12139 2483 12165 2539
rect 12221 2483 12247 2539
rect 12303 2483 12329 2539
rect 12385 2483 12411 2539
rect 12467 2483 12493 2539
rect 12549 2483 12575 2539
rect 12631 2483 12636 2539
rect 11754 2455 12636 2483
rect 11754 2399 11759 2455
rect 11815 2399 11840 2455
rect 11896 2399 11921 2455
rect 11977 2399 12002 2455
rect 12058 2399 12083 2455
rect 12139 2399 12165 2455
rect 12221 2399 12247 2455
rect 12303 2399 12329 2455
rect 12385 2399 12411 2455
rect 12467 2399 12493 2455
rect 12549 2399 12575 2455
rect 12631 2399 12636 2455
rect 11754 2371 12636 2399
rect 11754 2315 11759 2371
rect 11815 2315 11840 2371
rect 11896 2315 11921 2371
rect 11977 2315 12002 2371
rect 12058 2315 12083 2371
rect 12139 2315 12165 2371
rect 12221 2315 12247 2371
rect 12303 2315 12329 2371
rect 12385 2315 12411 2371
rect 12467 2315 12493 2371
rect 12549 2315 12575 2371
rect 12631 2315 12636 2371
rect 11754 2287 12636 2315
rect 11754 2231 11759 2287
rect 11815 2231 11840 2287
rect 11896 2231 11921 2287
rect 11977 2231 12002 2287
rect 12058 2231 12083 2287
rect 12139 2231 12165 2287
rect 12221 2231 12247 2287
rect 12303 2231 12329 2287
rect 12385 2231 12411 2287
rect 12467 2231 12493 2287
rect 12549 2231 12575 2287
rect 12631 2231 12636 2287
rect 11754 2203 12636 2231
rect 11754 2147 11759 2203
rect 11815 2147 11840 2203
rect 11896 2147 11921 2203
rect 11977 2147 12002 2203
rect 12058 2147 12083 2203
rect 12139 2147 12165 2203
rect 12221 2147 12247 2203
rect 12303 2147 12329 2203
rect 12385 2147 12411 2203
rect 12467 2147 12493 2203
rect 12549 2147 12575 2203
rect 12631 2147 12636 2203
rect 11754 2140 12636 2147
rect 7258 1965 7267 2021
rect 7323 1965 7349 2021
rect 7405 1965 7430 2021
rect 7486 1965 7511 2021
rect 7567 1965 7592 2021
rect 7648 1965 7657 2021
rect 7258 1897 7657 1965
rect 7258 1841 7267 1897
rect 7323 1841 7349 1897
rect 7405 1841 7430 1897
rect 7486 1841 7511 1897
rect 7567 1841 7592 1897
rect 7648 1841 7657 1897
rect 7258 -53 7657 1841
rect 7258 -109 7267 -53
rect 7323 -109 7349 -53
rect 7405 -109 7430 -53
rect 7486 -109 7511 -53
rect 7567 -109 7592 -53
rect 7648 -109 7657 -53
rect 7258 -137 7657 -109
rect 7258 -193 7267 -137
rect 7323 -193 7349 -137
rect 7405 -193 7430 -137
rect 7486 -193 7511 -137
rect 7567 -193 7592 -137
rect 7648 -193 7657 -137
rect 7258 -1565 7657 -193
rect 7258 -1621 7269 -1565
rect 7325 -1621 7375 -1565
rect 7431 -1621 7481 -1565
rect 7537 -1621 7587 -1565
rect 7643 -1621 7657 -1565
rect 7258 -1645 7657 -1621
rect 7258 -1701 7269 -1645
rect 7325 -1701 7375 -1645
rect 7431 -1701 7481 -1645
rect 7537 -1701 7587 -1645
rect 7643 -1701 7657 -1645
rect 7258 -1723 7657 -1701
rect 12811 2021 13210 2660
rect 12811 1965 12820 2021
rect 12876 1965 12901 2021
rect 12957 1965 12982 2021
rect 13038 1965 13063 2021
rect 13119 1965 13145 2021
rect 13201 1965 13210 2021
rect 12811 1897 13210 1965
rect 12811 1841 12820 1897
rect 12876 1841 12901 1897
rect 12957 1841 12982 1897
rect 13038 1841 13063 1897
rect 13119 1841 13145 1897
rect 13201 1841 13210 1897
rect 12811 -53 13210 1841
rect 12811 -109 12820 -53
rect 12876 -109 12902 -53
rect 12958 -109 12983 -53
rect 13039 -109 13064 -53
rect 13120 -109 13145 -53
rect 13201 -109 13210 -53
rect 12811 -137 13210 -109
rect 12811 -193 12820 -137
rect 12876 -193 12902 -137
rect 12958 -193 12983 -137
rect 13039 -193 13064 -137
rect 13120 -193 13145 -137
rect 13201 -193 13210 -137
rect 12811 -1565 13210 -193
rect 12811 -1621 12822 -1565
rect 12878 -1621 12903 -1565
rect 12959 -1621 12984 -1565
rect 12811 -1645 12984 -1621
rect 12811 -1701 12822 -1645
rect 12878 -1701 12903 -1645
rect 12959 -1701 12984 -1645
rect 13200 -1701 13210 -1565
rect 12811 -1728 13210 -1701
rect 13742 4453 14141 4469
rect 13742 4397 13751 4453
rect 13807 4397 13833 4453
rect 13889 4397 13914 4453
rect 13970 4397 13995 4453
rect 14051 4397 14076 4453
rect 14132 4397 14141 4453
rect 13742 4369 14141 4397
rect 13742 4313 13751 4369
rect 13807 4313 13833 4369
rect 13889 4313 13914 4369
rect 13970 4313 13995 4369
rect 14051 4313 14076 4369
rect 14132 4313 14141 4369
rect 13742 3065 14141 4313
rect 13742 3009 13751 3065
rect 13807 3009 13833 3065
rect 13889 3009 13914 3065
rect 13970 3009 13995 3065
rect 14051 3009 14076 3065
rect 14132 3009 14141 3065
rect 13742 2981 14141 3009
rect 13742 2925 13751 2981
rect 13807 2925 13833 2981
rect 13889 2925 13914 2981
rect 13970 2925 13995 2981
rect 14051 2925 14076 2981
rect 14132 2925 14141 2981
rect 13742 2840 14141 2925
rect 13742 2784 13751 2840
rect 13807 2784 13833 2840
rect 13889 2784 13914 2840
rect 13970 2784 13995 2840
rect 14051 2784 14076 2840
rect 14132 2784 14141 2840
rect 13742 2716 14141 2784
rect 13742 2660 13751 2716
rect 13807 2660 13833 2716
rect 13889 2660 13914 2716
rect 13970 2660 13995 2716
rect 14051 2660 14076 2716
rect 14132 2660 14141 2716
rect 13742 2021 14141 2660
rect 19380 4453 19694 4469
rect 19380 4397 19385 4453
rect 19441 4397 19467 4453
rect 19523 4397 19548 4453
rect 19604 4397 19629 4453
rect 19685 4397 19694 4453
rect 19380 4369 19694 4397
rect 19380 4313 19385 4369
rect 19441 4313 19467 4369
rect 19523 4313 19548 4369
rect 19604 4313 19629 4369
rect 19685 4313 19694 4369
rect 19380 3065 19694 4313
rect 19380 3009 19389 3065
rect 19445 3009 19469 3065
rect 19525 3009 19549 3065
rect 19605 3009 19629 3065
rect 19685 3009 19694 3065
rect 19380 2981 19694 3009
rect 19380 2925 19389 2981
rect 19445 2925 19469 2981
rect 19525 2925 19549 2981
rect 19605 2925 19629 2981
rect 19685 2925 19694 2981
rect 19380 2840 19694 2925
rect 19380 2784 19389 2840
rect 19445 2784 19469 2840
rect 19525 2784 19549 2840
rect 19605 2784 19629 2840
rect 19685 2784 19694 2840
rect 19380 2716 19694 2784
rect 19380 2660 19389 2716
rect 19445 2660 19469 2716
rect 19525 2660 19549 2716
rect 19605 2660 19629 2716
rect 19685 2660 19694 2716
rect 14316 2539 15198 2546
rect 14316 2483 14321 2539
rect 14377 2483 14403 2539
rect 14459 2483 14485 2539
rect 14541 2483 14567 2539
rect 14623 2483 14649 2539
rect 14705 2483 14731 2539
rect 14787 2483 14813 2539
rect 14869 2483 14894 2539
rect 14950 2483 14975 2539
rect 15031 2483 15056 2539
rect 15112 2483 15137 2539
rect 15193 2483 15198 2539
rect 14316 2455 15198 2483
rect 14316 2399 14321 2455
rect 14377 2399 14403 2455
rect 14459 2399 14485 2455
rect 14541 2399 14567 2455
rect 14623 2399 14649 2455
rect 14705 2399 14731 2455
rect 14787 2399 14813 2455
rect 14869 2399 14894 2455
rect 14950 2399 14975 2455
rect 15031 2399 15056 2455
rect 15112 2399 15137 2455
rect 15193 2399 15198 2455
rect 14316 2371 15198 2399
rect 14316 2315 14321 2371
rect 14377 2315 14403 2371
rect 14459 2315 14485 2371
rect 14541 2315 14567 2371
rect 14623 2315 14649 2371
rect 14705 2315 14731 2371
rect 14787 2315 14813 2371
rect 14869 2315 14894 2371
rect 14950 2315 14975 2371
rect 15031 2315 15056 2371
rect 15112 2315 15137 2371
rect 15193 2315 15198 2371
rect 14316 2287 15198 2315
rect 14316 2231 14321 2287
rect 14377 2231 14403 2287
rect 14459 2231 14485 2287
rect 14541 2231 14567 2287
rect 14623 2231 14649 2287
rect 14705 2231 14731 2287
rect 14787 2231 14813 2287
rect 14869 2231 14894 2287
rect 14950 2231 14975 2287
rect 15031 2231 15056 2287
rect 15112 2231 15137 2287
rect 15193 2231 15198 2287
rect 14316 2203 15198 2231
rect 14316 2147 14321 2203
rect 14377 2147 14403 2203
rect 14459 2147 14485 2203
rect 14541 2147 14567 2203
rect 14623 2147 14649 2203
rect 14705 2147 14731 2203
rect 14787 2147 14813 2203
rect 14869 2147 14894 2203
rect 14950 2147 14975 2203
rect 15031 2147 15056 2203
rect 15112 2147 15137 2203
rect 15193 2147 15198 2203
rect 14316 2140 15198 2147
rect 18238 2539 19120 2546
rect 18238 2483 18243 2539
rect 18299 2483 18324 2539
rect 18380 2483 18405 2539
rect 18461 2483 18486 2539
rect 18542 2483 18567 2539
rect 18623 2483 18649 2539
rect 18705 2483 18731 2539
rect 18787 2483 18813 2539
rect 18869 2483 18895 2539
rect 18951 2483 18977 2539
rect 19033 2483 19059 2539
rect 19115 2483 19120 2539
rect 18238 2455 19120 2483
rect 18238 2399 18243 2455
rect 18299 2399 18324 2455
rect 18380 2399 18405 2455
rect 18461 2399 18486 2455
rect 18542 2399 18567 2455
rect 18623 2399 18649 2455
rect 18705 2399 18731 2455
rect 18787 2399 18813 2455
rect 18869 2399 18895 2455
rect 18951 2399 18977 2455
rect 19033 2399 19059 2455
rect 19115 2399 19120 2455
rect 18238 2371 19120 2399
rect 18238 2315 18243 2371
rect 18299 2315 18324 2371
rect 18380 2315 18405 2371
rect 18461 2315 18486 2371
rect 18542 2315 18567 2371
rect 18623 2315 18649 2371
rect 18705 2315 18731 2371
rect 18787 2315 18813 2371
rect 18869 2315 18895 2371
rect 18951 2315 18977 2371
rect 19033 2315 19059 2371
rect 19115 2315 19120 2371
rect 18238 2287 19120 2315
rect 18238 2231 18243 2287
rect 18299 2231 18324 2287
rect 18380 2231 18405 2287
rect 18461 2231 18486 2287
rect 18542 2231 18567 2287
rect 18623 2231 18649 2287
rect 18705 2231 18731 2287
rect 18787 2231 18813 2287
rect 18869 2231 18895 2287
rect 18951 2231 18977 2287
rect 19033 2231 19059 2287
rect 19115 2231 19120 2287
rect 18238 2203 19120 2231
rect 18238 2147 18243 2203
rect 18299 2147 18324 2203
rect 18380 2147 18405 2203
rect 18461 2147 18486 2203
rect 18542 2147 18567 2203
rect 18623 2147 18649 2203
rect 18705 2147 18731 2203
rect 18787 2147 18813 2203
rect 18869 2147 18895 2203
rect 18951 2147 18977 2203
rect 19033 2147 19059 2203
rect 19115 2147 19120 2203
rect 18238 2140 19120 2147
rect 13742 1965 13751 2021
rect 13807 1965 13833 2021
rect 13889 1965 13914 2021
rect 13970 1965 13995 2021
rect 14051 1965 14076 2021
rect 14132 1965 14141 2021
rect 13742 1897 14141 1965
rect 13742 1841 13751 1897
rect 13807 1841 13833 1897
rect 13889 1841 13914 1897
rect 13970 1841 13995 1897
rect 14051 1841 14076 1897
rect 14132 1841 14141 1897
rect 13742 -53 14141 1841
rect 13742 -109 13751 -53
rect 13807 -109 13833 -53
rect 13889 -109 13914 -53
rect 13970 -109 13995 -53
rect 14051 -109 14076 -53
rect 14132 -109 14141 -53
rect 13742 -137 14141 -109
rect 13742 -193 13751 -137
rect 13807 -193 13833 -137
rect 13889 -193 13914 -137
rect 13970 -193 13995 -137
rect 14051 -193 14076 -137
rect 14132 -193 14141 -137
rect 13742 -1565 14141 -193
rect 13742 -1621 13753 -1565
rect 13809 -1621 13834 -1565
rect 13890 -1621 13915 -1565
rect 13742 -1645 13915 -1621
rect 13742 -1701 13753 -1645
rect 13809 -1701 13834 -1645
rect 13890 -1701 13915 -1645
rect 14131 -1701 14141 -1565
rect 13742 -1728 14141 -1701
rect 19380 2021 19694 2660
rect 19380 1965 19389 2021
rect 19445 1965 19469 2021
rect 19525 1965 19549 2021
rect 19605 1965 19629 2021
rect 19685 1965 19694 2021
rect 19380 1897 19694 1965
rect 19380 1841 19389 1897
rect 19445 1841 19469 1897
rect 19525 1841 19549 1897
rect 19605 1841 19629 1897
rect 19685 1841 19694 1897
rect 19380 -53 19694 1841
rect 19380 -109 19389 -53
rect 19445 -109 19469 -53
rect 19525 -109 19549 -53
rect 19605 -109 19629 -53
rect 19685 -109 19694 -53
rect 19380 -137 19694 -109
rect 19380 -193 19389 -137
rect 19445 -193 19469 -137
rect 19525 -193 19549 -137
rect 19605 -193 19629 -137
rect 19685 -193 19694 -137
rect 19380 -1565 19694 -193
rect 19380 -1621 19385 -1565
rect 19441 -1621 19466 -1565
rect 19522 -1621 19547 -1565
rect 19603 -1621 19628 -1565
rect 19684 -1621 19694 -1565
rect 19380 -1645 19694 -1621
rect 19380 -1701 19385 -1645
rect 19441 -1701 19466 -1645
rect 19522 -1701 19547 -1645
rect 19603 -1701 19628 -1645
rect 19684 -1701 19694 -1645
rect 19380 -1706 19694 -1701
use sky130_fd_io__gpio_ovtv2_hotswap_guardrings  sky130_fd_io__gpio_ovtv2_hotswap_guardrings_0
timestamp 1701704242
transform 1 0 -2627 0 1 -3247
box 0 0 26980 8664
use sky130_fd_io__tk_em2o_cdns_55959141808167  sky130_fd_io__tk_em2o_cdns_55959141808167_0
timestamp 1701704242
transform 0 1 19925 -1 0 2781
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_0
timestamp 1701704242
transform -1 0 7030 0 1 2482
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_1
timestamp 1701704242
transform -1 0 547 0 -1 2614
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_2
timestamp 1701704242
transform -1 0 547 0 1 2070
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_3
timestamp 1701704242
transform -1 0 3788 0 1 2070
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_4
timestamp 1701704242
transform -1 0 3788 0 1 2482
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_5
timestamp 1701704242
transform -1 0 7030 0 1 2070
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_6
timestamp 1701704242
transform -1 0 10272 0 -1 2614
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_7
timestamp 1701704242
transform -1 0 10272 0 1 2072
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_8
timestamp 1701704242
transform -1 0 13515 0 1 2070
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_9
timestamp 1701704242
transform -1 0 13515 0 -1 2614
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_10
timestamp 1701704242
transform 1 0 19921 0 1 2070
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_11
timestamp 1701704242
transform 1 0 19921 0 1 2482
box 0 0 1 1
<< labels >>
flabel metal2 s 20255 2576 20342 2614 3 FreeSans 200 0 0 0 SOFT_VCC_IO
port 4 nsew
flabel metal2 s 20280 2783 20355 2821 3 FreeSans 200 0 0 0 TIE_HI
port 5 nsew
flabel metal1 s 471 2345 532 2407 3 FreeSans 200 0 0 0 P2G
port 1 nsew
flabel metal1 s 10621 2255 10944 2490 3 FreeSans 200 0 0 0 PAD
port 2 nsew
flabel metal3 s 19380 3237 19694 3316 3 FreeSans 200 0 0 0 VPB_DRVR
port 3 nsew
<< properties >>
string GDS_END 70783934
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 70461792
<< end >>
