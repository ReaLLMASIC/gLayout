magic
tech sky130A
timestamp 1701704242
<< properties >>
string GDS_END 21561458
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 21561070
<< end >>
