magic
tech sky130B
timestamp 1701704242
<< viali >>
rect 0 0 449 89
<< metal1 >>
rect -6 89 455 92
rect -6 0 0 89
rect 449 0 455 89
rect -6 -3 455 0
<< properties >>
string GDS_END 86378038
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86375410
<< end >>
