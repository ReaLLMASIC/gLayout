magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< pwell >>
rect -76 -26 876 626
<< mvnmos >>
rect 0 0 800 600
<< mvndiff >>
rect -50 0 0 600
rect 800 0 850 600
<< poly >>
rect 0 600 800 626
rect 0 -26 800 0
<< metal1 >>
rect -51 -16 -5 546
rect 805 -16 851 546
use hvDFM1sd_CDNS_52468879185149  hvDFM1sd_CDNS_52468879185149_0
timestamp 1701704242
transform -1 0 0 0 1 0
box -26 -26 79 626
use hvDFM1sd_CDNS_52468879185149  hvDFM1sd_CDNS_52468879185149_1
timestamp 1701704242
transform 1 0 800 0 1 0
box -26 -26 79 626
<< labels >>
flabel comment s -28 265 -28 265 0 FreeSans 300 0 0 0 S
flabel comment s 828 265 828 265 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 86879154
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86878264
<< end >>
