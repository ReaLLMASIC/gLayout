magic
tech sky130A
timestamp 1701704242
<< properties >>
string GDS_END 20472658
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 20471758
<< end >>
