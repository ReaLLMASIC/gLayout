magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< pwell >>
rect -76 -26 10322 1426
<< nmos >>
rect 0 0 36 1400
rect 238 0 274 1400
rect 554 0 590 1400
rect 792 0 828 1400
rect 1108 0 1144 1400
rect 1346 0 1382 1400
rect 1662 0 1698 1400
rect 1900 0 1936 1400
rect 2216 0 2252 1400
rect 2454 0 2490 1400
rect 2770 0 2806 1400
rect 3008 0 3044 1400
rect 3324 0 3360 1400
rect 3562 0 3598 1400
rect 3878 0 3914 1400
rect 4116 0 4152 1400
rect 4432 0 4468 1400
rect 4670 0 4706 1400
rect 4986 0 5022 1400
rect 5224 0 5260 1400
rect 5540 0 5576 1400
rect 5778 0 5814 1400
rect 6094 0 6130 1400
rect 6332 0 6368 1400
rect 6648 0 6684 1400
rect 6886 0 6922 1400
rect 7202 0 7238 1400
rect 7440 0 7476 1400
rect 7756 0 7792 1400
rect 7994 0 8030 1400
rect 8310 0 8346 1400
rect 8548 0 8584 1400
rect 8864 0 8900 1400
rect 9102 0 9138 1400
rect 9418 0 9454 1400
rect 9656 0 9692 1400
rect 9972 0 10008 1400
rect 10210 0 10246 1400
<< ndiff >>
rect -50 0 0 1400
rect 36 0 238 1400
rect 274 0 314 1400
rect 514 0 554 1400
rect 590 0 792 1400
rect 828 0 868 1400
rect 1068 0 1108 1400
rect 1144 0 1346 1400
rect 1382 0 1422 1400
rect 1622 0 1662 1400
rect 1698 0 1900 1400
rect 1936 0 1976 1400
rect 2176 0 2216 1400
rect 2252 0 2454 1400
rect 2490 0 2530 1400
rect 2730 0 2770 1400
rect 2806 0 3008 1400
rect 3044 0 3084 1400
rect 3284 0 3324 1400
rect 3360 0 3562 1400
rect 3598 0 3638 1400
rect 3838 0 3878 1400
rect 3914 0 4116 1400
rect 4152 0 4192 1400
rect 4392 0 4432 1400
rect 4468 0 4670 1400
rect 4706 0 4746 1400
rect 4946 0 4986 1400
rect 5022 0 5224 1400
rect 5260 0 5300 1400
rect 5500 0 5540 1400
rect 5576 0 5778 1400
rect 5814 0 5854 1400
rect 6054 0 6094 1400
rect 6130 0 6332 1400
rect 6368 0 6408 1400
rect 6608 0 6648 1400
rect 6684 0 6886 1400
rect 6922 0 6962 1400
rect 7162 0 7202 1400
rect 7238 0 7440 1400
rect 7476 0 7516 1400
rect 7716 0 7756 1400
rect 7792 0 7994 1400
rect 8030 0 8070 1400
rect 8270 0 8310 1400
rect 8346 0 8548 1400
rect 8584 0 8624 1400
rect 8824 0 8864 1400
rect 8900 0 9102 1400
rect 9138 0 9178 1400
rect 9378 0 9418 1400
rect 9454 0 9656 1400
rect 9692 0 9732 1400
rect 9932 0 9972 1400
rect 10008 0 10210 1400
rect 10246 0 10296 1400
<< poly >>
rect 0 1400 36 1432
rect 238 1400 274 1432
rect 554 1400 590 1432
rect 792 1400 828 1432
rect 1108 1400 1144 1432
rect 1346 1400 1382 1432
rect 1662 1400 1698 1432
rect 1900 1400 1936 1432
rect 2216 1400 2252 1432
rect 2454 1400 2490 1432
rect 2770 1400 2806 1432
rect 3008 1400 3044 1432
rect 3324 1400 3360 1432
rect 3562 1400 3598 1432
rect 3878 1400 3914 1432
rect 4116 1400 4152 1432
rect 4432 1400 4468 1432
rect 4670 1400 4706 1432
rect 4986 1400 5022 1432
rect 5224 1400 5260 1432
rect 5540 1400 5576 1432
rect 5778 1400 5814 1432
rect 6094 1400 6130 1432
rect 6332 1400 6368 1432
rect 6648 1400 6684 1432
rect 6886 1400 6922 1432
rect 7202 1400 7238 1432
rect 7440 1400 7476 1432
rect 7756 1400 7792 1432
rect 7994 1400 8030 1432
rect 8310 1400 8346 1432
rect 8548 1400 8584 1432
rect 8864 1400 8900 1432
rect 9102 1400 9138 1432
rect 9418 1400 9454 1432
rect 9656 1400 9692 1432
rect 9972 1400 10008 1432
rect 10210 1400 10246 1432
rect 0 -32 36 0
rect 238 -32 274 0
rect 554 -32 590 0
rect 792 -32 828 0
rect 1108 -32 1144 0
rect 1346 -32 1382 0
rect 1662 -32 1698 0
rect 1900 -32 1936 0
rect 2216 -32 2252 0
rect 2454 -32 2490 0
rect 2770 -32 2806 0
rect 3008 -32 3044 0
rect 3324 -32 3360 0
rect 3562 -32 3598 0
rect 3878 -32 3914 0
rect 4116 -32 4152 0
rect 4432 -32 4468 0
rect 4670 -32 4706 0
rect 4986 -32 5022 0
rect 5224 -32 5260 0
rect 5540 -32 5576 0
rect 5778 -32 5814 0
rect 6094 -32 6130 0
rect 6332 -32 6368 0
rect 6648 -32 6684 0
rect 6886 -32 6922 0
rect 7202 -32 7238 0
rect 7440 -32 7476 0
rect 7756 -32 7792 0
rect 7994 -32 8030 0
rect 8310 -32 8346 0
rect 8548 -32 8584 0
rect 8864 -32 8900 0
rect 9102 -32 9138 0
rect 9418 -32 9454 0
rect 9656 -32 9692 0
rect 9972 -32 10008 0
rect 10210 -32 10246 0
<< locali >>
rect -229 -4 -51 1354
rect 325 -4 503 1354
rect 879 -4 1057 1354
rect 1433 -4 1611 1354
rect 1987 -4 2165 1354
rect 2541 -4 2719 1354
rect 3095 -4 3273 1354
rect 3649 -4 3827 1354
rect 4203 -4 4381 1354
rect 4757 -4 4935 1354
rect 5311 -4 5489 1354
rect 5865 -4 6043 1354
rect 6419 -4 6597 1354
rect 6973 -4 7151 1354
rect 7527 -4 7705 1354
rect 8081 -4 8259 1354
rect 8635 -4 8813 1354
rect 9189 -4 9367 1354
rect 9743 -4 9921 1354
rect 10297 -4 10475 1354
use DFTPL1s2_CDNS_55959141808702  DFTPL1s2_CDNS_55959141808702_0
timestamp 1701704242
transform -1 0 -40 0 1 0
box -26 -26 226 1426
use DFTPL1s2_CDNS_55959141808702  DFTPL1s2_CDNS_55959141808702_1
timestamp 1701704242
transform 1 0 314 0 1 0
box -26 -26 226 1426
use DFTPL1s2_CDNS_55959141808702  DFTPL1s2_CDNS_55959141808702_2
timestamp 1701704242
transform 1 0 868 0 1 0
box -26 -26 226 1426
use DFTPL1s2_CDNS_55959141808702  DFTPL1s2_CDNS_55959141808702_3
timestamp 1701704242
transform 1 0 1422 0 1 0
box -26 -26 226 1426
use DFTPL1s2_CDNS_55959141808702  DFTPL1s2_CDNS_55959141808702_4
timestamp 1701704242
transform 1 0 1976 0 1 0
box -26 -26 226 1426
use DFTPL1s2_CDNS_55959141808702  DFTPL1s2_CDNS_55959141808702_5
timestamp 1701704242
transform 1 0 2530 0 1 0
box -26 -26 226 1426
use DFTPL1s2_CDNS_55959141808702  DFTPL1s2_CDNS_55959141808702_6
timestamp 1701704242
transform 1 0 3084 0 1 0
box -26 -26 226 1426
use DFTPL1s2_CDNS_55959141808702  DFTPL1s2_CDNS_55959141808702_7
timestamp 1701704242
transform 1 0 3638 0 1 0
box -26 -26 226 1426
use DFTPL1s2_CDNS_55959141808702  DFTPL1s2_CDNS_55959141808702_8
timestamp 1701704242
transform 1 0 4192 0 1 0
box -26 -26 226 1426
use DFTPL1s2_CDNS_55959141808702  DFTPL1s2_CDNS_55959141808702_9
timestamp 1701704242
transform 1 0 4746 0 1 0
box -26 -26 226 1426
use DFTPL1s2_CDNS_55959141808702  DFTPL1s2_CDNS_55959141808702_10
timestamp 1701704242
transform 1 0 5300 0 1 0
box -26 -26 226 1426
use DFTPL1s2_CDNS_55959141808702  DFTPL1s2_CDNS_55959141808702_11
timestamp 1701704242
transform 1 0 5854 0 1 0
box -26 -26 226 1426
use DFTPL1s2_CDNS_55959141808702  DFTPL1s2_CDNS_55959141808702_12
timestamp 1701704242
transform 1 0 6408 0 1 0
box -26 -26 226 1426
use DFTPL1s2_CDNS_55959141808702  DFTPL1s2_CDNS_55959141808702_13
timestamp 1701704242
transform 1 0 6962 0 1 0
box -26 -26 226 1426
use DFTPL1s2_CDNS_55959141808702  DFTPL1s2_CDNS_55959141808702_14
timestamp 1701704242
transform 1 0 7516 0 1 0
box -26 -26 226 1426
use DFTPL1s2_CDNS_55959141808702  DFTPL1s2_CDNS_55959141808702_15
timestamp 1701704242
transform 1 0 8070 0 1 0
box -26 -26 226 1426
use DFTPL1s2_CDNS_55959141808702  DFTPL1s2_CDNS_55959141808702_16
timestamp 1701704242
transform 1 0 8624 0 1 0
box -26 -26 226 1426
use DFTPL1s2_CDNS_55959141808702  DFTPL1s2_CDNS_55959141808702_17
timestamp 1701704242
transform 1 0 9178 0 1 0
box -26 -26 226 1426
use DFTPL1s2_CDNS_55959141808702  DFTPL1s2_CDNS_55959141808702_18
timestamp 1701704242
transform 1 0 9732 0 1 0
box -26 -26 226 1426
use DFTPL1s2_CDNS_55959141808702  DFTPL1s2_CDNS_55959141808702_19
timestamp 1701704242
transform 1 0 10286 0 1 0
box -26 -26 226 1426
<< labels >>
flabel comment s 10386 675 10386 675 0 FreeSans 300 0 0 0 S
flabel comment s 10109 700 10109 700 0 FreeSans 300 0 0 0 D
flabel comment s 9832 675 9832 675 0 FreeSans 300 0 0 0 S
flabel comment s 9555 700 9555 700 0 FreeSans 300 0 0 0 D
flabel comment s 9278 675 9278 675 0 FreeSans 300 0 0 0 S
flabel comment s 9001 700 9001 700 0 FreeSans 300 0 0 0 D
flabel comment s 8724 675 8724 675 0 FreeSans 300 0 0 0 S
flabel comment s 8447 700 8447 700 0 FreeSans 300 0 0 0 D
flabel comment s 8170 675 8170 675 0 FreeSans 300 0 0 0 S
flabel comment s 7893 700 7893 700 0 FreeSans 300 0 0 0 D
flabel comment s 7616 675 7616 675 0 FreeSans 300 0 0 0 S
flabel comment s 7339 700 7339 700 0 FreeSans 300 0 0 0 D
flabel comment s 7062 675 7062 675 0 FreeSans 300 0 0 0 S
flabel comment s 6785 700 6785 700 0 FreeSans 300 0 0 0 D
flabel comment s 6508 675 6508 675 0 FreeSans 300 0 0 0 S
flabel comment s 6231 700 6231 700 0 FreeSans 300 0 0 0 D
flabel comment s 5954 675 5954 675 0 FreeSans 300 0 0 0 S
flabel comment s 5677 700 5677 700 0 FreeSans 300 0 0 0 D
flabel comment s 5400 675 5400 675 0 FreeSans 300 0 0 0 S
flabel comment s 5123 700 5123 700 0 FreeSans 300 0 0 0 D
flabel comment s 4846 675 4846 675 0 FreeSans 300 0 0 0 S
flabel comment s 4569 700 4569 700 0 FreeSans 300 0 0 0 D
flabel comment s 4292 675 4292 675 0 FreeSans 300 0 0 0 S
flabel comment s 4015 700 4015 700 0 FreeSans 300 0 0 0 D
flabel comment s 3738 675 3738 675 0 FreeSans 300 0 0 0 S
flabel comment s 3461 700 3461 700 0 FreeSans 300 0 0 0 D
flabel comment s 3184 675 3184 675 0 FreeSans 300 0 0 0 S
flabel comment s 2907 700 2907 700 0 FreeSans 300 0 0 0 D
flabel comment s 2630 675 2630 675 0 FreeSans 300 0 0 0 S
flabel comment s 2353 700 2353 700 0 FreeSans 300 0 0 0 D
flabel comment s 2076 675 2076 675 0 FreeSans 300 0 0 0 S
flabel comment s 1799 700 1799 700 0 FreeSans 300 0 0 0 D
flabel comment s 1522 675 1522 675 0 FreeSans 300 0 0 0 S
flabel comment s 1245 700 1245 700 0 FreeSans 300 0 0 0 D
flabel comment s 968 675 968 675 0 FreeSans 300 0 0 0 S
flabel comment s 691 700 691 700 0 FreeSans 300 0 0 0 D
flabel comment s 414 675 414 675 0 FreeSans 300 0 0 0 S
flabel comment s 137 700 137 700 0 FreeSans 300 0 0 0 D
flabel comment s -140 675 -140 675 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 43080326
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 43060846
<< end >>
