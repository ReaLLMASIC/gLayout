magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -38 261 1142 582
<< pwell >>
rect 1 21 1103 203
rect 29 -17 63 21
<< scnmos >>
rect 96 47 126 177
rect 182 47 212 177
rect 268 47 298 177
rect 354 47 384 177
rect 551 47 581 177
rect 637 47 667 177
rect 723 47 753 177
rect 809 47 839 177
rect 895 47 925 177
rect 981 47 1011 177
<< scpmoshvt >>
rect 96 297 126 497
rect 182 297 212 497
rect 268 297 298 497
rect 354 297 384 497
rect 440 297 470 497
rect 526 297 556 497
rect 723 297 753 497
rect 809 297 839 497
rect 895 297 925 497
rect 981 297 1011 497
<< ndiff >>
rect 27 157 96 177
rect 27 123 51 157
rect 85 123 96 157
rect 27 89 96 123
rect 27 55 51 89
rect 85 55 96 89
rect 27 47 96 55
rect 126 157 182 177
rect 126 123 137 157
rect 171 123 182 157
rect 126 47 182 123
rect 212 141 268 177
rect 212 107 224 141
rect 258 107 268 141
rect 212 47 268 107
rect 298 89 354 177
rect 298 55 310 89
rect 344 55 354 89
rect 298 47 354 55
rect 384 158 443 177
rect 384 124 401 158
rect 435 124 443 158
rect 384 47 443 124
rect 497 165 551 177
rect 497 131 506 165
rect 540 131 551 165
rect 497 47 551 131
rect 581 89 637 177
rect 581 55 592 89
rect 626 55 637 89
rect 581 47 637 55
rect 667 132 723 177
rect 667 98 677 132
rect 711 98 723 132
rect 667 47 723 98
rect 753 94 809 177
rect 753 60 764 94
rect 798 60 809 94
rect 753 47 809 60
rect 839 132 895 177
rect 839 98 850 132
rect 884 98 895 132
rect 839 47 895 98
rect 925 94 981 177
rect 925 60 936 94
rect 970 60 981 94
rect 925 47 981 60
rect 1011 133 1077 177
rect 1011 99 1034 133
rect 1068 99 1077 133
rect 1011 47 1077 99
<< pdiff >>
rect 43 477 96 497
rect 43 443 51 477
rect 85 443 96 477
rect 43 386 96 443
rect 43 352 51 386
rect 85 352 96 386
rect 43 297 96 352
rect 126 477 182 497
rect 126 443 137 477
rect 171 443 182 477
rect 126 384 182 443
rect 126 350 137 384
rect 171 350 182 384
rect 126 297 182 350
rect 212 485 268 497
rect 212 451 223 485
rect 257 451 268 485
rect 212 417 268 451
rect 212 383 223 417
rect 257 383 268 417
rect 212 297 268 383
rect 298 477 354 497
rect 298 443 309 477
rect 343 443 354 477
rect 298 386 354 443
rect 298 352 309 386
rect 343 352 354 386
rect 298 297 354 352
rect 384 485 440 497
rect 384 451 395 485
rect 429 451 440 485
rect 384 417 440 451
rect 384 383 395 417
rect 429 383 440 417
rect 384 297 440 383
rect 470 477 526 497
rect 470 443 481 477
rect 515 443 526 477
rect 470 386 526 443
rect 470 352 481 386
rect 515 352 526 386
rect 470 297 526 352
rect 556 485 609 497
rect 556 451 567 485
rect 601 451 609 485
rect 556 417 609 451
rect 556 383 567 417
rect 601 383 609 417
rect 556 297 609 383
rect 664 489 723 497
rect 664 455 678 489
rect 712 455 723 489
rect 664 417 723 455
rect 664 383 678 417
rect 712 383 723 417
rect 664 297 723 383
rect 753 397 809 497
rect 753 363 764 397
rect 798 363 809 397
rect 753 297 809 363
rect 839 489 895 497
rect 839 455 850 489
rect 884 455 895 489
rect 839 421 895 455
rect 839 387 850 421
rect 884 387 895 421
rect 839 353 895 387
rect 839 319 850 353
rect 884 319 895 353
rect 839 297 895 319
rect 925 489 981 497
rect 925 455 936 489
rect 970 455 981 489
rect 925 421 981 455
rect 925 387 936 421
rect 970 387 981 421
rect 925 297 981 387
rect 1011 477 1077 497
rect 1011 443 1022 477
rect 1056 443 1077 477
rect 1011 380 1077 443
rect 1011 346 1022 380
rect 1056 346 1077 380
rect 1011 297 1077 346
<< ndiffc >>
rect 51 123 85 157
rect 51 55 85 89
rect 137 123 171 157
rect 224 107 258 141
rect 310 55 344 89
rect 401 124 435 158
rect 506 131 540 165
rect 592 55 626 89
rect 677 98 711 132
rect 764 60 798 94
rect 850 98 884 132
rect 936 60 970 94
rect 1034 99 1068 133
<< pdiffc >>
rect 51 443 85 477
rect 51 352 85 386
rect 137 443 171 477
rect 137 350 171 384
rect 223 451 257 485
rect 223 383 257 417
rect 309 443 343 477
rect 309 352 343 386
rect 395 451 429 485
rect 395 383 429 417
rect 481 443 515 477
rect 481 352 515 386
rect 567 451 601 485
rect 567 383 601 417
rect 678 455 712 489
rect 678 383 712 417
rect 764 363 798 397
rect 850 455 884 489
rect 850 387 884 421
rect 850 319 884 353
rect 936 455 970 489
rect 936 387 970 421
rect 1022 443 1056 477
rect 1022 346 1056 380
<< poly >>
rect 96 497 126 523
rect 182 497 212 523
rect 268 497 298 523
rect 354 497 384 523
rect 440 497 470 523
rect 526 497 556 523
rect 723 497 753 523
rect 809 497 839 523
rect 895 497 925 523
rect 981 497 1011 523
rect 96 265 126 297
rect 182 265 212 297
rect 25 249 212 265
rect 25 215 35 249
rect 69 215 212 249
rect 25 199 212 215
rect 96 177 126 199
rect 182 177 212 199
rect 268 259 298 297
rect 354 259 384 297
rect 268 249 384 259
rect 268 215 308 249
rect 342 215 384 249
rect 268 205 384 215
rect 440 259 470 297
rect 526 259 556 297
rect 723 259 753 297
rect 809 259 839 297
rect 440 249 667 259
rect 440 215 456 249
rect 490 215 587 249
rect 621 215 667 249
rect 440 205 667 215
rect 268 177 298 205
rect 354 177 384 205
rect 551 177 581 205
rect 637 177 667 205
rect 723 249 839 259
rect 723 215 766 249
rect 800 215 839 249
rect 723 205 839 215
rect 723 177 753 205
rect 809 177 839 205
rect 895 259 925 297
rect 981 259 1011 297
rect 895 249 1011 259
rect 895 215 943 249
rect 977 215 1011 249
rect 895 205 1011 215
rect 895 177 925 205
rect 981 177 1011 205
rect 96 21 126 47
rect 182 21 212 47
rect 268 21 298 47
rect 354 21 384 47
rect 551 21 581 47
rect 637 21 667 47
rect 723 21 753 47
rect 809 21 839 47
rect 895 21 925 47
rect 981 21 1011 47
<< polycont >>
rect 35 215 69 249
rect 308 215 342 249
rect 456 215 490 249
rect 587 215 621 249
rect 766 215 800 249
rect 943 215 977 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 35 477 85 527
rect 35 443 51 477
rect 35 386 85 443
rect 35 352 51 386
rect 35 305 85 352
rect 121 477 173 493
rect 121 443 137 477
rect 171 443 173 477
rect 121 384 173 443
rect 121 350 137 384
rect 171 350 173 384
rect 207 485 273 527
rect 207 451 223 485
rect 257 451 273 485
rect 207 417 273 451
rect 207 383 223 417
rect 257 383 273 417
rect 207 367 273 383
rect 307 477 345 493
rect 307 443 309 477
rect 343 443 345 477
rect 307 386 345 443
rect 121 333 173 350
rect 307 352 309 386
rect 343 352 345 386
rect 379 485 445 527
rect 379 451 395 485
rect 429 451 445 485
rect 379 417 445 451
rect 379 383 395 417
rect 429 383 445 417
rect 379 368 445 383
rect 479 477 515 493
rect 479 443 481 477
rect 479 386 515 443
rect 307 333 345 352
rect 479 352 481 386
rect 551 485 617 527
rect 551 451 567 485
rect 601 451 617 485
rect 551 417 617 451
rect 551 383 567 417
rect 601 383 617 417
rect 551 367 617 383
rect 662 489 900 493
rect 662 455 678 489
rect 712 455 850 489
rect 884 455 900 489
rect 662 417 714 455
rect 848 421 900 455
rect 662 383 678 417
rect 712 383 714 417
rect 662 367 714 383
rect 763 397 801 421
rect 479 333 515 352
rect 763 363 764 397
rect 798 363 801 397
rect 763 333 801 363
rect 121 299 801 333
rect 848 387 850 421
rect 884 387 900 421
rect 848 353 900 387
rect 934 489 986 527
rect 934 455 936 489
rect 970 455 986 489
rect 934 421 986 455
rect 934 387 936 421
rect 970 387 986 421
rect 934 371 986 387
rect 1020 477 1072 493
rect 1020 443 1022 477
rect 1056 443 1072 477
rect 1020 380 1072 443
rect 848 319 850 353
rect 884 337 900 353
rect 1020 346 1022 380
rect 1056 346 1072 380
rect 1020 337 1072 346
rect 884 319 1072 337
rect 848 303 1072 319
rect 17 249 85 271
rect 17 215 35 249
rect 69 215 85 249
rect 121 181 173 299
rect 209 249 358 265
rect 209 215 308 249
rect 342 215 358 249
rect 440 249 637 265
rect 440 215 456 249
rect 490 215 587 249
rect 621 215 637 249
rect 673 249 891 265
rect 673 215 766 249
rect 800 215 891 249
rect 927 249 1087 265
rect 927 215 943 249
rect 977 215 1087 249
rect 35 157 87 173
rect 35 123 51 157
rect 85 123 87 157
rect 121 157 187 181
rect 121 123 137 157
rect 171 123 187 157
rect 223 158 455 181
rect 223 147 401 158
rect 223 141 260 147
rect 35 89 87 123
rect 223 107 224 141
rect 258 107 260 141
rect 385 124 401 147
rect 435 124 455 158
rect 490 165 1087 168
rect 490 131 506 165
rect 540 133 1087 165
rect 540 132 1034 133
rect 540 131 677 132
rect 223 89 260 107
rect 35 55 51 89
rect 85 55 260 89
rect 35 52 260 55
rect 294 106 352 113
rect 294 89 355 106
rect 676 98 677 131
rect 711 131 850 132
rect 711 98 714 131
rect 576 89 642 97
rect 294 55 310 89
rect 344 55 592 89
rect 626 55 642 89
rect 676 73 714 98
rect 848 98 850 131
rect 884 130 1034 132
rect 884 98 886 130
rect 748 94 814 97
rect 294 51 642 55
rect 748 60 764 94
rect 798 60 814 94
rect 848 73 886 98
rect 1020 99 1034 130
rect 1068 99 1087 133
rect 920 94 986 96
rect 748 17 814 60
rect 920 60 936 94
rect 970 60 986 94
rect 1020 73 1087 99
rect 920 17 986 60
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
<< metal1 >>
rect 0 561 1104 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 0 496 1104 527
rect 0 17 1104 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
rect 0 -48 1104 -17
<< labels >>
flabel locali s 1041 221 1075 255 0 FreeSans 400 0 0 0 A1
port 1 nsew signal input
flabel locali s 949 221 983 255 0 FreeSans 400 0 0 0 A1
port 1 nsew signal input
flabel locali s 765 221 799 255 0 FreeSans 400 0 0 0 A2
port 2 nsew signal input
flabel locali s 581 221 615 255 0 FreeSans 400 0 0 0 B1
port 3 nsew signal input
flabel locali s 489 221 523 255 0 FreeSans 400 0 0 0 B1
port 3 nsew signal input
flabel locali s 305 221 339 255 0 FreeSans 400 0 0 0 C1
port 4 nsew signal input
flabel locali s 29 221 63 255 0 FreeSans 400 0 0 0 D1
port 5 nsew signal input
flabel locali s 121 289 155 323 0 FreeSans 400 0 0 0 Y
port 10 nsew signal output
flabel locali s 121 221 155 255 0 FreeSans 400 0 0 0 Y
port 10 nsew signal output
flabel locali s 121 153 155 187 0 FreeSans 400 0 0 0 Y
port 10 nsew signal output
flabel locali s 121 425 155 459 0 FreeSans 400 0 0 0 Y
port 10 nsew signal output
flabel locali s 121 357 155 391 0 FreeSans 400 0 0 0 Y
port 10 nsew signal output
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional abutment
rlabel comment s 0 0 0 0 4 o2111ai_2
rlabel metal1 s 0 -48 1104 48 1 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1104 592 1 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1104 544
string GDS_END 960620
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 951156
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 5.520 0.000 
<< end >>
