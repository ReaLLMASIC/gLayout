magic
tech sky130B
magscale 1 2
timestamp 1701704242
use sky130_fd_pr__hvdftpm1s2__example_55959141808649  sky130_fd_pr__hvdftpm1s2__example_55959141808649_0
timestamp 1701704242
transform -1 0 -91 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 17339324
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 17338466
<< end >>
