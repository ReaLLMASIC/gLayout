magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< pwell >>
rect -76 -26 1732 326
<< mvnmos >>
rect 0 0 800 300
rect 856 0 1656 300
<< mvndiff >>
rect -50 0 0 300
rect 1656 0 1706 300
<< poly >>
rect 0 300 800 332
rect 0 -32 800 0
rect 856 300 1656 332
rect 856 -32 1656 0
<< metal1 >>
rect -51 -16 -5 258
rect 805 -16 851 258
rect 1661 -16 1707 258
use hvDFM1sd2_CDNS_52468879185892  hvDFM1sd2_CDNS_52468879185892_0
timestamp 1701704242
transform -1 0 0 0 1 0
box -26 -26 82 326
use hvDFM1sd2_CDNS_52468879185892  hvDFM1sd2_CDNS_52468879185892_1
timestamp 1701704242
transform 1 0 1656 0 1 0
box -26 -26 82 326
use hvDFM1sd2_CDNS_52468879185892  hvDFM1sd2_CDNS_52468879185892_2
timestamp 1701704242
transform 1 0 800 0 1 0
box -26 -26 82 326
<< labels >>
flabel comment s -28 121 -28 121 0 FreeSans 300 0 0 0 S
flabel comment s 828 121 828 121 0 FreeSans 300 0 0 0 D
flabel comment s 1684 121 1684 121 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 6104066
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 6102672
<< end >>
