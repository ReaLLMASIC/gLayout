magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -119 -66 4623 666
<< mvpmos >>
rect 0 0 400 600
rect 456 0 856 600
rect 912 0 1312 600
rect 1368 0 1768 600
rect 1824 0 2224 600
rect 2280 0 2680 600
rect 2736 0 3136 600
rect 3192 0 3592 600
rect 3648 0 4048 600
rect 4104 0 4504 600
<< mvpdiff >>
rect -50 0 0 600
rect 4504 0 4554 600
<< poly >>
rect 0 600 400 626
rect 0 -26 400 0
rect 456 600 856 626
rect 456 -26 856 0
rect 912 600 1312 626
rect 912 -26 1312 0
rect 1368 600 1768 626
rect 1368 -26 1768 0
rect 1824 600 2224 626
rect 1824 -26 2224 0
rect 2280 600 2680 626
rect 2280 -26 2680 0
rect 2736 600 3136 626
rect 2736 -26 3136 0
rect 3192 600 3592 626
rect 3192 -26 3592 0
rect 3648 600 4048 626
rect 3648 -26 4048 0
rect 4104 600 4504 626
rect 4104 -26 4504 0
<< metal1 >>
rect -51 -16 -5 546
rect 405 -16 451 546
rect 861 -16 907 546
rect 1317 -16 1363 546
rect 1773 -16 1819 546
rect 2229 -16 2275 546
rect 2685 -16 2731 546
rect 3141 -16 3187 546
rect 3597 -16 3643 546
rect 4053 -16 4099 546
rect 4509 -16 4555 546
use hvDFM1sd2_CDNS_5246887918599  hvDFM1sd2_CDNS_5246887918599_0
timestamp 1701704242
transform 1 0 4048 0 1 0
box -36 -36 92 636
use hvDFM1sd2_CDNS_5246887918599  hvDFM1sd2_CDNS_5246887918599_1
timestamp 1701704242
transform 1 0 3592 0 1 0
box -36 -36 92 636
use hvDFM1sd2_CDNS_5246887918599  hvDFM1sd2_CDNS_5246887918599_2
timestamp 1701704242
transform 1 0 3136 0 1 0
box -36 -36 92 636
use hvDFM1sd2_CDNS_5246887918599  hvDFM1sd2_CDNS_5246887918599_3
timestamp 1701704242
transform 1 0 2680 0 1 0
box -36 -36 92 636
use hvDFM1sd2_CDNS_5246887918599  hvDFM1sd2_CDNS_5246887918599_4
timestamp 1701704242
transform 1 0 2224 0 1 0
box -36 -36 92 636
use hvDFM1sd2_CDNS_5246887918599  hvDFM1sd2_CDNS_5246887918599_5
timestamp 1701704242
transform 1 0 1768 0 1 0
box -36 -36 92 636
use hvDFM1sd2_CDNS_5246887918599  hvDFM1sd2_CDNS_5246887918599_6
timestamp 1701704242
transform 1 0 1312 0 1 0
box -36 -36 92 636
use hvDFM1sd2_CDNS_5246887918599  hvDFM1sd2_CDNS_5246887918599_7
timestamp 1701704242
transform 1 0 856 0 1 0
box -36 -36 92 636
use hvDFM1sd2_CDNS_5246887918599  hvDFM1sd2_CDNS_5246887918599_8
timestamp 1701704242
transform 1 0 400 0 1 0
box -36 -36 92 636
use hvDFM1sd_CDNS_52468879185167  hvDFM1sd_CDNS_52468879185167_0
timestamp 1701704242
transform -1 0 0 0 1 0
box -36 -36 89 636
use hvDFM1sd_CDNS_52468879185167  hvDFM1sd_CDNS_52468879185167_1
timestamp 1701704242
transform 1 0 4504 0 1 0
box -36 -36 89 636
<< labels >>
flabel comment s -28 265 -28 265 0 FreeSans 300 0 0 0 S
flabel comment s 428 265 428 265 0 FreeSans 300 0 0 0 D
flabel comment s 884 265 884 265 0 FreeSans 300 0 0 0 S
flabel comment s 1340 265 1340 265 0 FreeSans 300 0 0 0 D
flabel comment s 1796 265 1796 265 0 FreeSans 300 0 0 0 S
flabel comment s 2252 265 2252 265 0 FreeSans 300 0 0 0 D
flabel comment s 2708 265 2708 265 0 FreeSans 300 0 0 0 S
flabel comment s 3164 265 3164 265 0 FreeSans 300 0 0 0 D
flabel comment s 3620 265 3620 265 0 FreeSans 300 0 0 0 S
flabel comment s 4076 265 4076 265 0 FreeSans 300 0 0 0 D
flabel comment s 4532 265 4532 265 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 86846762
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86841262
<< end >>
