magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< pwell >>
rect 4478 858 5187 1328
rect 4965 -7 5187 858
<< psubdiff >>
rect 4504 1278 5161 1302
rect 4504 1244 4565 1278
rect 4599 1244 4633 1278
rect 4667 1244 4701 1278
rect 4735 1244 4769 1278
rect 4803 1244 4837 1278
rect 4871 1244 4905 1278
rect 4939 1244 4991 1278
rect 5025 1244 5059 1278
rect 5093 1244 5127 1278
rect 4504 1207 5161 1244
rect 4504 1194 4991 1207
rect 4504 1160 4565 1194
rect 4599 1160 4633 1194
rect 4667 1160 4701 1194
rect 4735 1160 4769 1194
rect 4803 1160 4837 1194
rect 4871 1160 4905 1194
rect 4939 1173 4991 1194
rect 5025 1173 5059 1207
rect 5093 1173 5127 1207
rect 4939 1160 5161 1173
rect 4504 1136 5161 1160
rect 4504 1111 4991 1136
rect 4504 1077 4565 1111
rect 4599 1077 4633 1111
rect 4667 1077 4701 1111
rect 4735 1077 4769 1111
rect 4803 1077 4837 1111
rect 4871 1077 4905 1111
rect 4939 1102 4991 1111
rect 5025 1102 5059 1136
rect 5093 1102 5127 1136
rect 4939 1077 5161 1102
rect 4504 1065 5161 1077
rect 4504 1031 4991 1065
rect 5025 1031 5059 1065
rect 5093 1031 5127 1065
rect 4504 1028 5161 1031
rect 4504 994 4565 1028
rect 4599 994 4633 1028
rect 4667 994 4701 1028
rect 4735 994 4769 1028
rect 4803 994 4837 1028
rect 4871 994 4905 1028
rect 4939 994 5161 1028
rect 4504 960 4991 994
rect 5025 960 5059 994
rect 5093 960 5127 994
rect 4504 923 5161 960
rect 4504 889 4991 923
rect 5025 889 5059 923
rect 5093 889 5127 923
rect 4504 884 5161 889
rect 4991 852 5161 884
rect 5025 818 5059 852
rect 5093 818 5127 852
rect 4991 781 5161 818
rect 5025 747 5059 781
rect 5093 747 5127 781
rect 4991 710 5161 747
rect 5025 676 5059 710
rect 5093 676 5127 710
rect 4991 639 5161 676
rect 5025 605 5059 639
rect 5093 605 5127 639
rect 4991 568 5161 605
rect 5025 534 5059 568
rect 5093 534 5127 568
rect 4991 497 5161 534
rect 5025 463 5059 497
rect 5093 463 5127 497
rect 4991 427 5161 463
rect 5025 393 5059 427
rect 5093 393 5127 427
rect 4991 357 5161 393
rect 5025 323 5059 357
rect 5093 323 5127 357
rect 4991 287 5161 323
rect 5025 253 5059 287
rect 5093 253 5127 287
rect 4991 217 5161 253
rect 5025 183 5059 217
rect 5093 183 5127 217
rect 4991 147 5161 183
rect 5025 113 5059 147
rect 5093 113 5127 147
rect 4991 77 5161 113
rect 5025 43 5059 77
rect 5093 43 5127 77
rect 4991 19 5161 43
<< psubdiffcont >>
rect 4565 1244 4599 1278
rect 4633 1244 4667 1278
rect 4701 1244 4735 1278
rect 4769 1244 4803 1278
rect 4837 1244 4871 1278
rect 4905 1244 4939 1278
rect 4991 1244 5025 1278
rect 5059 1244 5093 1278
rect 5127 1244 5161 1278
rect 4565 1160 4599 1194
rect 4633 1160 4667 1194
rect 4701 1160 4735 1194
rect 4769 1160 4803 1194
rect 4837 1160 4871 1194
rect 4905 1160 4939 1194
rect 4991 1173 5025 1207
rect 5059 1173 5093 1207
rect 5127 1173 5161 1207
rect 4565 1077 4599 1111
rect 4633 1077 4667 1111
rect 4701 1077 4735 1111
rect 4769 1077 4803 1111
rect 4837 1077 4871 1111
rect 4905 1077 4939 1111
rect 4991 1102 5025 1136
rect 5059 1102 5093 1136
rect 5127 1102 5161 1136
rect 4991 1031 5025 1065
rect 5059 1031 5093 1065
rect 5127 1031 5161 1065
rect 4565 994 4599 1028
rect 4633 994 4667 1028
rect 4701 994 4735 1028
rect 4769 994 4803 1028
rect 4837 994 4871 1028
rect 4905 994 4939 1028
rect 4991 960 5025 994
rect 5059 960 5093 994
rect 5127 960 5161 994
rect 4991 889 5025 923
rect 5059 889 5093 923
rect 5127 889 5161 923
rect 4991 818 5025 852
rect 5059 818 5093 852
rect 5127 818 5161 852
rect 4991 747 5025 781
rect 5059 747 5093 781
rect 5127 747 5161 781
rect 4991 676 5025 710
rect 5059 676 5093 710
rect 5127 676 5161 710
rect 4991 605 5025 639
rect 5059 605 5093 639
rect 5127 605 5161 639
rect 4991 534 5025 568
rect 5059 534 5093 568
rect 5127 534 5161 568
rect 4991 463 5025 497
rect 5059 463 5093 497
rect 5127 463 5161 497
rect 4991 393 5025 427
rect 5059 393 5093 427
rect 5127 393 5161 427
rect 4991 323 5025 357
rect 5059 323 5093 357
rect 5127 323 5161 357
rect 4991 253 5025 287
rect 5059 253 5093 287
rect 5127 253 5161 287
rect 4991 183 5025 217
rect 5059 183 5093 217
rect 5127 183 5161 217
rect 4991 113 5025 147
rect 5059 113 5093 147
rect 5127 113 5161 147
rect 4991 43 5025 77
rect 5059 43 5093 77
rect 5127 43 5161 77
<< locali >>
rect 126 2634 160 2668
rect 302 2634 336 2668
rect 1578 2634 1612 2668
rect 1822 2634 1856 2668
rect 2394 2634 2428 2668
rect 2678 2634 2712 2668
rect 3316 2634 3350 2668
rect 3492 2634 3526 2668
rect 3954 2634 3988 2668
rect 4768 2634 4802 2668
rect 5122 2634 5156 2668
rect 5474 2634 5508 2668
rect 5528 2474 5562 2508
rect 4164 2332 4198 2370
rect 5262 2388 5296 2426
rect 4362 1802 4396 1840
rect 4504 1278 5161 1302
rect 4504 1244 4565 1278
rect 4599 1244 4633 1278
rect 4667 1244 4701 1278
rect 4735 1244 4769 1278
rect 4803 1244 4837 1278
rect 4871 1244 4905 1278
rect 4939 1244 4991 1278
rect 5025 1244 5059 1278
rect 5093 1244 5127 1278
rect 498 1194 536 1228
rect 870 1194 908 1228
rect 2162 1194 2200 1228
rect 2516 1194 2554 1228
rect 3776 1148 3882 1234
rect 4162 1194 4200 1228
rect 4504 1207 5161 1244
rect 4504 1194 4991 1207
rect 3810 1114 3848 1148
rect 4504 1160 4565 1194
rect 4599 1160 4633 1194
rect 4667 1160 4701 1194
rect 4735 1160 4769 1194
rect 4803 1160 4837 1194
rect 4871 1160 4905 1194
rect 4939 1173 4991 1194
rect 5025 1173 5059 1207
rect 5093 1173 5127 1207
rect 4939 1160 5161 1173
rect 4504 1136 5161 1160
rect 4504 1111 4991 1136
rect 4504 1077 4565 1111
rect 4599 1077 4633 1111
rect 4667 1077 4701 1111
rect 4735 1077 4769 1111
rect 4803 1077 4837 1111
rect 4871 1077 4905 1111
rect 4939 1102 4991 1111
rect 5025 1102 5059 1136
rect 5093 1102 5127 1136
rect 4939 1077 5161 1102
rect 4504 1065 5161 1077
rect 4504 1031 4991 1065
rect 5025 1031 5059 1065
rect 5093 1031 5127 1065
rect 4504 1028 5161 1031
rect 4504 994 4565 1028
rect 4599 994 4633 1028
rect 4667 994 4701 1028
rect 4735 994 4769 1028
rect 4803 994 4837 1028
rect 4871 994 4905 1028
rect 4939 994 5161 1028
rect 4504 960 4991 994
rect 5025 960 5059 994
rect 5093 960 5127 994
rect 4504 923 5161 960
rect 1359 884 1393 918
rect 4504 889 4991 923
rect 5025 889 5059 923
rect 5093 889 5127 923
rect 4504 884 5161 889
rect 4991 852 5161 884
rect 5025 818 5059 852
rect 5093 818 5127 852
rect 4991 781 5161 818
rect 5025 747 5059 781
rect 5093 747 5127 781
rect 4991 710 5161 747
rect 5025 676 5059 710
rect 5093 676 5127 710
rect 129 622 163 656
rect 1263 622 1296 656
rect 1775 622 1809 656
rect 2909 622 2943 656
rect 3421 622 3455 656
rect 4555 622 4589 656
rect 4991 639 5161 676
rect 5025 605 5059 639
rect 5093 605 5127 639
rect 4991 568 5161 605
rect 5025 534 5059 568
rect 5093 534 5127 568
rect 4991 497 5161 534
rect 5025 463 5059 497
rect 5093 463 5127 497
rect 4991 427 5161 463
rect 5025 393 5059 427
rect 5093 393 5127 427
rect 4991 357 5161 393
rect 5025 323 5059 357
rect 5093 323 5127 357
rect 4991 287 5161 323
rect 5025 253 5059 287
rect 5093 253 5127 287
rect 4991 217 5161 253
rect 5025 183 5059 217
rect 5093 183 5127 217
rect 4991 147 5161 183
rect 5025 113 5059 147
rect 5093 113 5127 147
rect 4991 77 5161 113
rect 1611 36 1646 70
rect 5025 43 5059 77
rect 5093 43 5127 77
rect 4991 19 5161 43
<< viali >>
rect 5262 2426 5296 2460
rect 4164 2370 4198 2404
rect 5262 2354 5296 2388
rect 4164 2298 4198 2332
rect 4362 1840 4396 1874
rect 4362 1768 4396 1802
rect 464 1194 498 1228
rect 536 1194 570 1228
rect 836 1194 870 1228
rect 908 1194 942 1228
rect 2128 1194 2162 1228
rect 2200 1194 2234 1228
rect 2482 1194 2516 1228
rect 2554 1194 2588 1228
rect 4128 1194 4162 1228
rect 4200 1194 4234 1228
rect 3776 1114 3810 1148
rect 3848 1114 3882 1148
<< metal1 >>
tri 4122 2460 4128 2466 se
rect 4128 2460 5308 2466
tri 4104 2442 4122 2460 se
rect 4122 2442 5262 2460
rect -210 2414 1269 2442
tri 1239 2404 1249 2414 ne
rect 1249 2404 1269 2414
tri 1249 2390 1263 2404 ne
rect 1263 2390 1269 2404
rect 1321 2390 1333 2442
rect 1385 2426 2256 2442
tri 2256 2426 2272 2442 sw
tri 3716 2426 3732 2442 se
rect 3732 2438 5262 2442
rect 3732 2426 4128 2438
tri 4128 2426 4140 2438 nw
tri 5075 2426 5087 2438 ne
rect 5087 2426 5262 2438
rect 5296 2426 5308 2460
rect 1385 2414 2272 2426
rect 1385 2410 1411 2414
tri 1411 2410 1415 2414 nw
tri 2244 2410 2248 2414 ne
rect 2248 2410 2272 2414
tri 2272 2410 2288 2426 sw
tri 3700 2410 3716 2426 se
rect 3716 2414 4116 2426
tri 4116 2414 4128 2426 nw
tri 5087 2414 5099 2426 ne
rect 5099 2414 5308 2426
rect 3716 2410 3740 2414
tri 3740 2410 3744 2414 nw
tri 5099 2410 5103 2414 ne
rect 5103 2410 5308 2414
rect 1385 2404 1405 2410
tri 1405 2404 1411 2410 nw
tri 2248 2404 2254 2410 ne
rect 2254 2404 2288 2410
tri 2288 2404 2294 2410 sw
tri 3694 2404 3700 2410 se
rect 3700 2404 3734 2410
tri 3734 2404 3740 2410 nw
tri 4146 2404 4152 2410 se
rect 4152 2404 4210 2410
rect 1385 2402 1403 2404
tri 1403 2402 1405 2404 nw
tri 2254 2402 2256 2404 ne
rect 2256 2402 2294 2404
tri 2294 2402 2296 2404 sw
tri 3692 2402 3694 2404 se
rect 3694 2402 3732 2404
tri 3732 2402 3734 2404 nw
tri 4144 2402 4146 2404 se
rect 4146 2402 4164 2404
rect 1385 2390 1391 2402
tri 1391 2390 1403 2402 nw
tri 2256 2390 2268 2402 ne
rect 2268 2390 2296 2402
tri 2296 2390 2308 2402 sw
tri 3680 2390 3692 2402 se
rect 3692 2390 3700 2402
tri 2268 2386 2272 2390 ne
rect 2272 2386 2308 2390
tri 2308 2386 2312 2390 sw
tri 3676 2386 3680 2390 se
rect 3680 2386 3700 2390
rect -210 2358 204 2386
tri 174 2354 178 2358 ne
rect 178 2354 204 2358
tri 178 2334 198 2354 ne
rect 198 2334 204 2354
rect 256 2334 268 2386
rect 320 2370 781 2386
tri 781 2370 797 2386 sw
tri 2001 2370 2017 2386 se
rect 2017 2370 2232 2386
tri 2232 2370 2248 2386 sw
tri 2272 2370 2288 2386 ne
rect 2288 2370 2312 2386
tri 2312 2370 2328 2386 sw
tri 3660 2370 3676 2386 se
rect 3676 2370 3700 2386
tri 3700 2370 3732 2402 nw
tri 4128 2386 4144 2402 se
rect 4144 2386 4164 2402
tri 3759 2370 3775 2386 se
rect 3775 2370 4164 2386
rect 4198 2370 4210 2404
tri 5103 2388 5125 2410 ne
rect 5125 2388 5308 2410
rect 320 2361 797 2370
tri 797 2361 806 2370 sw
tri 1992 2361 2001 2370 se
rect 2001 2361 2248 2370
rect 320 2358 806 2361
rect 320 2354 346 2358
tri 346 2354 350 2358 nw
tri 768 2354 772 2358 ne
rect 772 2354 806 2358
tri 806 2354 813 2361 sw
tri 1985 2354 1992 2361 se
rect 1992 2358 2248 2361
rect 1992 2354 2025 2358
tri 2025 2354 2029 2358 nw
tri 2220 2354 2224 2358 ne
rect 2224 2354 2248 2358
tri 2248 2354 2264 2370 sw
tri 2288 2354 2304 2370 ne
rect 2304 2354 3684 2370
tri 3684 2354 3700 2370 nw
tri 3743 2354 3759 2370 se
rect 3759 2358 4210 2370
rect 3759 2354 3783 2358
tri 3783 2354 3787 2358 nw
tri 4127 2354 4131 2358 ne
rect 4131 2354 4210 2358
tri 5125 2354 5159 2388 ne
rect 5159 2354 5262 2388
rect 5296 2354 5308 2388
rect 320 2334 326 2354
tri 326 2334 346 2354 nw
tri 772 2334 792 2354 ne
rect 792 2346 813 2354
tri 813 2346 821 2354 sw
tri 1977 2346 1985 2354 se
rect 1985 2346 2017 2354
tri 2017 2346 2025 2354 nw
tri 2224 2346 2232 2354 ne
rect 2232 2346 2264 2354
rect 792 2334 821 2346
tri 821 2334 833 2346 sw
tri 1965 2334 1977 2346 se
rect 1977 2334 2003 2346
tri 792 2332 794 2334 ne
rect 794 2332 833 2334
tri 833 2332 835 2334 sw
tri 1963 2332 1965 2334 se
rect 1965 2332 2003 2334
tri 2003 2332 2017 2346 nw
tri 2232 2332 2246 2346 ne
rect 2246 2342 2264 2346
tri 2264 2342 2276 2354 sw
tri 2304 2342 2316 2354 ne
rect 2316 2342 3672 2354
tri 3672 2342 3684 2354 nw
tri 3735 2346 3743 2354 se
rect 3743 2346 3775 2354
tri 3775 2346 3783 2354 nw
tri 4131 2346 4139 2354 ne
rect 4139 2346 4210 2354
tri 5159 2348 5165 2354 ne
rect 5165 2348 5308 2354
tri 3731 2342 3735 2346 se
rect 3735 2342 3761 2346
rect 2246 2334 2276 2342
tri 2276 2334 2284 2342 sw
tri 3723 2334 3731 2342 se
rect 3731 2334 3761 2342
rect 2246 2332 2284 2334
tri 2284 2332 2286 2334 sw
tri 3721 2332 3723 2334 se
rect 3723 2332 3761 2334
tri 3761 2332 3775 2346 nw
tri 4139 2333 4152 2346 ne
rect 4152 2332 4210 2346
tri 794 2320 806 2332 ne
rect 806 2320 835 2332
tri 835 2320 847 2332 sw
tri 1951 2320 1963 2332 se
rect 1963 2320 1991 2332
tri 1991 2320 2003 2332 nw
tri 2246 2320 2258 2332 ne
rect 2258 2320 2286 2332
tri 806 2314 812 2320 ne
rect 812 2314 1985 2320
tri 1985 2314 1991 2320 nw
tri 2258 2314 2264 2320 ne
rect 2264 2314 2286 2320
tri 2286 2314 2304 2332 sw
tri 3703 2314 3721 2332 se
rect 3721 2314 3743 2332
tri 3743 2314 3761 2332 nw
tri 812 2298 828 2314 ne
rect 828 2298 1969 2314
tri 1969 2298 1985 2314 nw
tri 2264 2298 2280 2314 ne
rect 2280 2298 3727 2314
tri 3727 2298 3743 2314 nw
rect 4152 2298 4164 2332
rect 4198 2298 4210 2332
tri 828 2292 834 2298 ne
rect 834 2292 1963 2298
tri 1963 2292 1969 2298 nw
tri 2280 2292 2286 2298 ne
rect 2286 2292 3721 2298
tri 3721 2292 3727 2298 nw
rect 4152 2292 4210 2298
tri 2286 2286 2292 2292 ne
rect 2292 2286 3715 2292
tri 3715 2286 3721 2292 nw
rect 1823 2212 1829 2264
rect 1881 2212 1893 2264
rect 1945 2212 1951 2264
rect -210 1982 60 2184
rect 72 2059 105 2092
tri -14 1908 60 1982 ne
rect 4344 1828 4350 1880
rect 4402 1828 4408 1880
rect 4344 1816 4408 1828
rect 4344 1764 4350 1816
rect 4402 1764 4408 1816
rect 4344 1762 4408 1764
rect 4452 1826 4458 1878
rect 4510 1826 4516 1878
rect 4452 1814 4516 1826
rect 4452 1760 4458 1814
rect 4510 1762 4516 1814
tri -14 1658 60 1732 se
rect 66 1692 100 1726
rect -210 1456 60 1658
rect 69 1593 106 1628
rect 2023 1356 2029 1408
rect 2081 1356 2093 1408
rect 2145 1356 2151 1408
rect -210 1262 5801 1328
rect 198 1182 204 1234
rect 256 1182 268 1234
rect 320 1228 582 1234
rect 320 1194 464 1228
rect 498 1194 536 1228
rect 570 1194 582 1228
rect 320 1182 582 1194
rect 720 1228 1315 1234
rect 720 1194 836 1228
rect 870 1194 908 1228
rect 942 1194 1263 1228
rect 720 1182 1263 1194
tri 1238 1157 1263 1182 ne
rect 2023 1182 2029 1234
rect 2081 1182 2093 1234
rect 2145 1228 2246 1234
rect 2162 1194 2200 1228
rect 2234 1194 2246 1228
rect 2145 1182 2246 1194
rect 2470 1228 2600 1234
rect 2470 1194 2482 1228
rect 2516 1194 2554 1228
rect 2588 1194 2600 1228
rect 1263 1164 1315 1176
tri 2445 1154 2470 1179 se
rect 2470 1154 2600 1194
rect 4116 1228 4286 1234
rect 4116 1194 4128 1228
rect 4162 1194 4200 1228
rect 4234 1194 4286 1228
rect 4116 1182 4286 1194
rect 4338 1182 4350 1234
rect 4402 1182 4408 1234
rect 1263 1106 1315 1112
rect 1823 1102 1829 1154
rect 1881 1102 1893 1154
rect 1945 1102 2600 1154
rect 3764 1148 4394 1154
rect 3764 1114 3776 1148
rect 3810 1114 3848 1148
rect 3882 1114 4394 1148
rect 3764 1102 4394 1114
rect 4446 1102 4458 1154
rect 4510 1102 4516 1154
rect 1519 816 1553 850
rect 1519 338 1553 372
<< via1 >>
rect 1269 2390 1321 2442
rect 1333 2390 1385 2442
rect 204 2334 256 2386
rect 268 2334 320 2386
rect 1829 2212 1881 2264
rect 1893 2212 1945 2264
rect 4350 1874 4402 1880
rect 4350 1840 4362 1874
rect 4362 1840 4396 1874
rect 4396 1840 4402 1874
rect 4350 1828 4402 1840
rect 4350 1802 4402 1816
rect 4350 1768 4362 1802
rect 4362 1768 4396 1802
rect 4396 1768 4402 1802
rect 4350 1764 4402 1768
rect 4458 1826 4510 1878
rect 4458 1762 4510 1814
rect 2029 1356 2081 1408
rect 2093 1356 2145 1408
rect 204 1182 256 1234
rect 268 1182 320 1234
rect 1263 1176 1315 1228
rect 2029 1182 2081 1234
rect 2093 1228 2145 1234
rect 2093 1194 2128 1228
rect 2128 1194 2145 1228
rect 2093 1182 2145 1194
rect 1263 1112 1315 1164
rect 4286 1182 4338 1234
rect 4350 1182 4402 1234
rect 1829 1102 1881 1154
rect 1893 1102 1945 1154
rect 4394 1102 4446 1154
rect 4458 1102 4510 1154
<< metal2 >>
rect 1263 2390 1269 2442
rect 1321 2390 1333 2442
rect 1385 2390 1391 2442
rect 1263 2386 1336 2390
tri 1336 2386 1340 2390 nw
rect 198 2334 204 2386
rect 256 2334 268 2386
rect 320 2334 326 2386
rect 198 1234 326 2334
rect 198 1182 204 1234
rect 256 1182 268 1234
rect 320 1182 326 1234
rect 1263 1228 1315 2386
tri 1315 2365 1336 2386 nw
rect 1263 1164 1315 1176
rect 1263 1106 1315 1112
rect 1823 2212 1829 2264
rect 1881 2212 1893 2264
rect 1945 2212 1951 2264
rect 1823 1154 1951 2212
rect 4344 1828 4350 1880
rect 4402 1828 4408 1880
rect 4344 1816 4408 1828
rect 4344 1764 4350 1816
rect 4402 1764 4408 1816
rect 2023 1356 2029 1408
rect 2081 1356 2093 1408
rect 2145 1356 2151 1408
rect 2023 1234 2151 1356
tri 4319 1234 4344 1259 se
rect 4344 1234 4408 1764
rect 2023 1182 2029 1234
rect 2081 1182 2093 1234
rect 2145 1182 2151 1234
rect 4280 1182 4286 1234
rect 4338 1182 4350 1234
rect 4402 1182 4408 1234
rect 4452 1826 4458 1878
rect 4510 1826 4516 1878
rect 4452 1814 4516 1826
rect 4452 1762 4458 1814
rect 4510 1762 4516 1814
tri 4427 1154 4452 1179 se
rect 4452 1154 4516 1762
rect 1823 1102 1829 1154
rect 1881 1102 1893 1154
rect 1945 1102 1951 1154
rect 4388 1102 4394 1154
rect 4446 1102 4458 1154
rect 4510 1102 4516 1154
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_0
timestamp 1701704242
transform -1 0 4198 0 1 2298
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_1
timestamp 1701704242
transform 1 0 5262 0 -1 2460
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_2
timestamp 1701704242
transform 1 0 4362 0 -1 1874
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1701704242
transform 1 0 464 0 1 1194
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1701704242
transform 1 0 836 0 1 1194
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1701704242
transform 1 0 2128 0 1 1194
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_3
timestamp 1701704242
transform 1 0 2482 0 1 1194
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_4
timestamp 1701704242
transform 1 0 3776 0 1 1114
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_5
timestamp 1701704242
transform 1 0 4128 0 1 1194
box 0 0 1 1
use L1M1_CDNS_52468879185316  L1M1_CDNS_52468879185316_0
timestamp 1701704242
transform 1 0 4551 0 1 1268
box -12 -6 622 40
use L1M1_CDNS_52468879185955  L1M1_CDNS_52468879185955_0
timestamp 1701704242
transform -1 0 2835 0 1 1268
box -12 -6 982 40
use L1M1_CDNS_52468879185955  L1M1_CDNS_52468879185955_1
timestamp 1701704242
transform -1 0 1186 0 1 1268
box -12 -6 982 40
use L1M1_CDNS_52468879185955  L1M1_CDNS_52468879185955_2
timestamp 1701704242
transform -1 0 4480 0 1 1268
box -12 -6 982 40
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_0
timestamp 1701704242
transform 0 1 1263 -1 0 1234
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_1
timestamp 1701704242
transform -1 0 1391 0 -1 2442
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_2
timestamp 1701704242
transform 1 0 198 0 1 1182
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_3
timestamp 1701704242
transform 1 0 2023 0 1 1182
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_4
timestamp 1701704242
transform 1 0 4280 0 1 1182
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_5
timestamp 1701704242
transform 1 0 198 0 1 2334
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_6
timestamp 1701704242
transform 1 0 2023 0 1 1356
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_7
timestamp 1701704242
transform 1 0 1823 0 1 2212
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_8
timestamp 1701704242
transform 1 0 1823 0 1 1102
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_9
timestamp 1701704242
transform 1 0 4388 0 1 1102
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_0
timestamp 1701704242
transform 1 0 4344 0 -1 1880
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_1
timestamp 1701704242
transform 1 0 4452 0 -1 1878
box 0 0 1 1
use sky130_fd_io__sio_com_ictl_logic  sky130_fd_io__sio_com_ictl_logic_0
timestamp 1701704242
transform 1 0 -50 0 1 1315
box 32 0 5818 1369
use sky130_fd_io__sio_com_ictl_outls_bank  sky130_fd_io__sio_com_ictl_outls_bank_0
timestamp 1701704242
transform 1 0 -110 0 1 53
box -94 -53 5015 1275
<< labels >>
flabel comment s 4232 1209 4232 1209 0 FreeSans 200 0 0 0 ie_diff_sel__h
flabel comment s 4232 1131 4232 1131 0 FreeSans 200 0 0 0 ie_diff_sel__h_n
flabel comment s 1966 1136 1966 1136 0 FreeSans 200 0 0 0 inp_dis_i_h
flabel comment s 2282 1384 2282 1384 0 FreeSans 200 0 0 0 inp_dis_i_h_n
flabel comment s -102 2376 -102 2376 0 FreeSans 200 0 0 0 ie_se_sel_h_n
flabel comment s -102 2429 -102 2429 0 FreeSans 200 0 0 0 ie_se_sel_h
flabel metal1 s 66 1692 100 1726 0 FreeSans 200 0 0 0 vgnd
port 3 nsew
flabel metal1 s 69 1593 106 1628 0 FreeSans 200 0 0 0 vgnd
port 3 nsew
flabel metal1 s 1519 338 1553 372 0 FreeSans 200 0 0 0 vpwr_ka
port 2 nsew
flabel metal1 s 1519 816 1553 850 0 FreeSans 200 0 0 0 vgnd
port 3 nsew
flabel metal1 s 72 2059 105 2092 0 FreeSans 200 0 0 0 vcc_io
port 4 nsew
flabel metal1 s 2554 1194 2589 1228 0 FreeSans 200 0 0 0 inp_dis_i_h
port 5 nsew
flabel locali s 1359 884 1393 918 0 FreeSans 200 0 0 0 vgnd
port 3 nsew
flabel locali s 5122 2634 5156 2668 0 FreeSans 200 0 0 0 vtrip_sel_h
port 6 nsew
flabel locali s 1611 36 1646 70 0 FreeSans 200 0 0 0 vpb_ka
port 7 nsew
flabel locali s 5474 2634 5508 2668 0 FreeSans 200 0 0 0 tripsel_i_h_n
port 8 nsew
flabel locali s 5528 2474 5562 2508 0 FreeSans 200 0 0 0 tripsel_i_h
port 9 nsew
flabel locali s 2909 622 2943 656 0 FreeSans 200 0 0 0 inp_dis_i_n
port 10 nsew
flabel locali s 1775 622 1809 656 0 FreeSans 200 0 0 0 inp_dis_i
port 11 nsew
flabel locali s 1822 2634 1856 2668 0 FreeSans 200 0 0 0 inp_dis_h
port 12 nsew
flabel locali s 1263 622 1296 656 0 FreeSans 200 0 0 0 ie_se_sel_n
port 13 nsew
flabel locali s 129 622 163 656 0 FreeSans 200 0 0 0 ie_se_sel
port 14 nsew
flabel locali s 4555 622 4589 656 0 FreeSans 200 0 0 0 ie_diff_sel_n
port 15 nsew
flabel locali s 3421 622 3455 656 0 FreeSans 200 0 0 0 ie_diff_sel
port 16 nsew
flabel locali s 3954 2634 3988 2668 0 FreeSans 200 0 0 0 ibuf_sel_h_n
port 17 nsew
flabel locali s 4768 2634 4802 2668 0 FreeSans 200 0 0 0 ibuf_sel_h
port 18 nsew
flabel locali s 2678 2634 2712 2668 0 FreeSans 200 0 0 0 dm_h_n<2>
port 19 nsew
flabel locali s 3316 2634 3350 2668 0 FreeSans 200 0 0 0 dm_h_n<1>
port 20 nsew
flabel locali s 3492 2634 3526 2668 0 FreeSans 200 0 0 0 dm_h_n<0>
port 21 nsew
flabel locali s 302 2634 336 2668 0 FreeSans 200 0 0 0 dm_h<2>
port 22 nsew
flabel locali s 126 2634 160 2668 0 FreeSans 200 0 0 0 dm_h<1>
port 23 nsew
flabel locali s 1578 2634 1612 2668 0 FreeSans 200 0 0 0 dm_h<0>
port 24 nsew
flabel locali s 2394 2634 2428 2668 0 FreeSans 200 0 0 0 inp_dis_h_n
port 25 nsew
flabel metal2 s 2072 1193 2102 1223 0 FreeSans 200 0 0 0 inp_dis_i_h_n
port 26 nsew
flabel metal2 s 215 1193 245 1223 0 FreeSans 200 0 0 0 ie_se_sel_h_n
port 27 nsew
flabel metal2 s 1273 1187 1304 1217 0 FreeSans 200 0 0 0 ie_se_sel_h
port 28 nsew
flabel metal2 s 4405 1113 4435 1143 0 FreeSans 200 0 0 0 ie_diff_sel_h_n
port 29 nsew
flabel metal2 s 4298 1193 4327 1223 0 FreeSans 200 0 0 0 ie_diff_sel_h
port 30 nsew
<< properties >>
string GDS_END 85555696
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85541568
string path 126.900 32.550 126.900 0.475 
<< end >>
