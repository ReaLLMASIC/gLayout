magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< via4 >>
rect 1247 14758 1483 14994
rect 1567 14758 1803 14994
rect 1887 14758 2123 14994
rect 2207 14758 2443 14994
rect 2527 14758 2763 14994
rect 2847 14758 3083 14994
rect 3167 14758 3403 14994
rect 3487 14758 3723 14994
rect 3807 14758 4043 14994
rect 4127 14758 4363 14994
rect 4447 14758 4683 14994
rect 4767 14758 5003 14994
rect 5087 14758 5323 14994
rect 5407 14758 5643 14994
rect 5727 14758 5963 14994
rect 6047 14758 6283 14994
rect 6367 14758 6603 14994
rect 6687 14758 6923 14994
rect 7007 14758 7243 14994
rect 7327 14758 7563 14994
rect 7647 14758 7883 14994
rect 7967 14758 8203 14994
rect 8287 14758 8523 14994
rect 8607 14758 8843 14994
rect 8927 14758 9163 14994
rect 9247 14758 9483 14994
rect 9567 14758 9803 14994
rect 9887 14758 10123 14994
rect 10207 14758 10443 14994
rect 10527 14758 10763 14994
rect 10847 14758 11083 14994
rect 11167 14758 11403 14994
rect 11487 14758 11723 14994
rect 925 14450 1161 14686
rect 11849 14396 12085 14632
rect 605 14130 841 14366
rect 12169 14076 12405 14312
rect 285 13810 521 14046
rect 12489 13756 12725 13992
rect -38 13487 198 13723
rect -38 13167 198 13403
rect 12758 13393 12994 13629
rect -38 12847 198 13083
rect 12758 13073 12994 13309
rect -38 12527 198 12763
rect 12758 12753 12994 12989
rect -38 12207 198 12443
rect 12758 12433 12994 12669
rect -38 11887 198 12123
rect 12758 12113 12994 12349
rect -38 11567 198 11803
rect 12758 11793 12994 12029
rect -38 11247 198 11483
rect 12758 11473 12994 11709
rect -38 10927 198 11163
rect 12758 11153 12994 11389
rect -38 10607 198 10843
rect 12758 10833 12994 11069
rect -38 10287 198 10523
rect 12758 10513 12994 10749
rect -38 9967 198 10203
rect 12758 10193 12994 10429
rect -38 9647 198 9883
rect 12758 9873 12994 10109
rect -38 9327 198 9563
rect 12758 9553 12994 9789
rect -38 9007 198 9243
rect 12758 9233 12994 9469
rect -38 8687 198 8923
rect 12758 8913 12994 9149
rect -38 8367 198 8603
rect 12758 8593 12994 8829
rect -38 8047 198 8283
rect 12758 8273 12994 8509
rect -38 7727 198 7963
rect 12758 7953 12994 8189
rect -38 7407 198 7643
rect 12758 7633 12994 7869
rect -38 7087 198 7323
rect 12758 7313 12994 7549
rect -38 6767 198 7003
rect 12758 6993 12994 7229
rect -38 6447 198 6683
rect 12758 6673 12994 6909
rect -38 6127 198 6363
rect 12758 6353 12994 6589
rect -38 5807 198 6043
rect 12758 6033 12994 6269
rect -38 5487 198 5723
rect 12758 5713 12994 5949
rect -38 5167 198 5403
rect 12758 5393 12994 5629
rect -38 4847 198 5083
rect 12758 5073 12994 5309
rect -38 4527 198 4763
rect 12758 4753 12994 4989
rect -38 4207 198 4443
rect 12758 4433 12994 4669
rect -38 3887 198 4123
rect 12758 4113 12994 4349
rect -38 3567 198 3803
rect 12758 3793 12994 4029
rect -38 3247 198 3483
rect 12758 3473 12994 3709
rect -38 2927 198 3163
rect 12758 3153 12994 3389
rect -38 2607 198 2843
rect 12758 2833 12994 3069
rect -38 2287 198 2523
rect 12758 2513 12994 2749
rect -38 1967 198 2203
rect 12758 2193 12994 2429
rect -38 1647 198 1883
rect 12758 1873 12994 2109
rect -38 1327 198 1563
rect 12758 1553 12994 1789
rect 12758 1233 12994 1469
rect 231 964 467 1200
rect 12435 910 12671 1146
rect 551 644 787 880
rect 12115 590 12351 826
rect 871 324 1107 560
rect 11795 270 12031 506
rect 1233 -38 1469 198
rect 1553 -38 1789 198
rect 1873 -38 2109 198
rect 2193 -38 2429 198
rect 2513 -38 2749 198
rect 2833 -38 3069 198
rect 3153 -38 3389 198
rect 3473 -38 3709 198
rect 3793 -38 4029 198
rect 4113 -38 4349 198
rect 4433 -38 4669 198
rect 4753 -38 4989 198
rect 5073 -38 5309 198
rect 5393 -38 5629 198
rect 5713 -38 5949 198
rect 6033 -38 6269 198
rect 6353 -38 6589 198
rect 6673 -38 6909 198
rect 6993 -38 7229 198
rect 7313 -38 7549 198
rect 7633 -38 7869 198
rect 7953 -38 8189 198
rect 8273 -38 8509 198
rect 8593 -38 8829 198
rect 8913 -38 9149 198
rect 9233 -38 9469 198
rect 9553 -38 9789 198
rect 9873 -38 10109 198
rect 10193 -38 10429 198
rect 10513 -38 10749 198
rect 10833 -38 11069 198
rect 11153 -38 11389 198
rect 11473 -38 11709 198
<< properties >>
string GDS_END 85508626
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85498638
<< end >>
