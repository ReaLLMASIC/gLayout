magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -119 -66 999 1066
<< mvpmos >>
rect 0 0 100 1000
rect 156 0 256 1000
rect 312 0 412 1000
rect 468 0 568 1000
rect 624 0 724 1000
rect 780 0 880 1000
<< mvpdiff >>
rect -50 0 0 1000
rect 880 0 930 1000
<< poly >>
rect 0 1000 100 1026
rect 0 -26 100 0
rect 156 1000 256 1026
rect 156 -26 256 0
rect 312 1000 412 1026
rect 312 -26 412 0
rect 468 1000 568 1026
rect 468 -26 568 0
rect 624 1000 724 1026
rect 624 -26 724 0
rect 780 1000 880 1026
rect 780 -26 880 0
<< locali >>
rect -45 -4 -11 946
rect 111 -4 145 946
rect 267 -4 301 946
rect 423 -4 457 946
rect 579 -4 613 946
rect 735 -4 769 946
rect 891 -4 925 946
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_0
timestamp 1701704242
transform 1 0 724 0 1 0
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_1
timestamp 1701704242
transform 1 0 568 0 1 0
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_2
timestamp 1701704242
transform 1 0 412 0 1 0
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_3
timestamp 1701704242
transform 1 0 256 0 1 0
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_4
timestamp 1701704242
transform 1 0 100 0 1 0
box -36 -36 92 1036
use hvDFL1sd_CDNS_52468879185112  hvDFL1sd_CDNS_52468879185112_0
timestamp 1701704242
transform -1 0 0 0 1 0
box -36 -36 89 1036
use hvDFL1sd_CDNS_52468879185112  hvDFL1sd_CDNS_52468879185112_1
timestamp 1701704242
transform 1 0 880 0 1 0
box -36 -36 89 1036
<< labels >>
flabel comment s -28 471 -28 471 0 FreeSans 300 0 0 0 S
flabel comment s 128 471 128 471 0 FreeSans 300 0 0 0 D
flabel comment s 284 471 284 471 0 FreeSans 300 0 0 0 S
flabel comment s 440 471 440 471 0 FreeSans 300 0 0 0 D
flabel comment s 596 471 596 471 0 FreeSans 300 0 0 0 S
flabel comment s 752 471 752 471 0 FreeSans 300 0 0 0 D
flabel comment s 908 471 908 471 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 87563398
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 87559890
<< end >>
