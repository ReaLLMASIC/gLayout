magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< dnwell >>
tri -500 6514 -414 6600 se
rect -414 6514 564 6600
tri 564 6514 650 6600 sw
rect -500 -514 650 6514
tri -500 -600 -414 -514 ne
rect -414 -600 564 -514
tri 564 -600 650 -514 nw
<< nwell >>
rect -10 0 160 6000
<< pwell >>
rect -1866 6874 2016 7008
rect -1866 6026 -1732 6874
rect 1882 6026 2016 6874
rect -1866 -26 -374 6026
rect 524 -26 2016 6026
rect -1866 -874 -1732 -26
rect 1882 -874 2016 -26
rect -1866 -1008 2016 -874
<< mvnnmos >>
rect -1600 0 -400 6000
rect 550 0 1750 6000
<< mvndiff >>
rect -1658 5975 -1600 6000
rect -1658 5941 -1646 5975
rect -1612 5941 -1600 5975
rect -1658 5907 -1600 5941
rect -1658 5873 -1646 5907
rect -1612 5873 -1600 5907
rect -1658 5839 -1600 5873
rect -1658 5805 -1646 5839
rect -1612 5805 -1600 5839
rect -1658 5771 -1600 5805
rect -1658 5737 -1646 5771
rect -1612 5737 -1600 5771
rect -1658 5703 -1600 5737
rect -1658 5669 -1646 5703
rect -1612 5669 -1600 5703
rect -1658 5635 -1600 5669
rect -1658 5601 -1646 5635
rect -1612 5601 -1600 5635
rect -1658 5567 -1600 5601
rect -1658 5533 -1646 5567
rect -1612 5533 -1600 5567
rect -1658 5499 -1600 5533
rect -1658 5465 -1646 5499
rect -1612 5465 -1600 5499
rect -1658 5431 -1600 5465
rect -1658 5397 -1646 5431
rect -1612 5397 -1600 5431
rect -1658 5363 -1600 5397
rect -1658 5329 -1646 5363
rect -1612 5329 -1600 5363
rect -1658 5295 -1600 5329
rect -1658 5261 -1646 5295
rect -1612 5261 -1600 5295
rect -1658 5227 -1600 5261
rect -1658 5193 -1646 5227
rect -1612 5193 -1600 5227
rect -1658 5159 -1600 5193
rect -1658 5125 -1646 5159
rect -1612 5125 -1600 5159
rect -1658 5091 -1600 5125
rect -1658 5057 -1646 5091
rect -1612 5057 -1600 5091
rect -1658 5023 -1600 5057
rect -1658 4989 -1646 5023
rect -1612 4989 -1600 5023
rect -1658 4955 -1600 4989
rect -1658 4921 -1646 4955
rect -1612 4921 -1600 4955
rect -1658 4887 -1600 4921
rect -1658 4853 -1646 4887
rect -1612 4853 -1600 4887
rect -1658 4819 -1600 4853
rect -1658 4785 -1646 4819
rect -1612 4785 -1600 4819
rect -1658 4751 -1600 4785
rect -1658 4717 -1646 4751
rect -1612 4717 -1600 4751
rect -1658 4683 -1600 4717
rect -1658 4649 -1646 4683
rect -1612 4649 -1600 4683
rect -1658 4615 -1600 4649
rect -1658 4581 -1646 4615
rect -1612 4581 -1600 4615
rect -1658 4547 -1600 4581
rect -1658 4513 -1646 4547
rect -1612 4513 -1600 4547
rect -1658 4479 -1600 4513
rect -1658 4445 -1646 4479
rect -1612 4445 -1600 4479
rect -1658 4411 -1600 4445
rect -1658 4377 -1646 4411
rect -1612 4377 -1600 4411
rect -1658 4343 -1600 4377
rect -1658 4309 -1646 4343
rect -1612 4309 -1600 4343
rect -1658 4275 -1600 4309
rect -1658 4241 -1646 4275
rect -1612 4241 -1600 4275
rect -1658 4207 -1600 4241
rect -1658 4173 -1646 4207
rect -1612 4173 -1600 4207
rect -1658 4139 -1600 4173
rect -1658 4105 -1646 4139
rect -1612 4105 -1600 4139
rect -1658 4071 -1600 4105
rect -1658 4037 -1646 4071
rect -1612 4037 -1600 4071
rect -1658 4003 -1600 4037
rect -1658 3969 -1646 4003
rect -1612 3969 -1600 4003
rect -1658 3935 -1600 3969
rect -1658 3901 -1646 3935
rect -1612 3901 -1600 3935
rect -1658 3867 -1600 3901
rect -1658 3833 -1646 3867
rect -1612 3833 -1600 3867
rect -1658 3799 -1600 3833
rect -1658 3765 -1646 3799
rect -1612 3765 -1600 3799
rect -1658 3731 -1600 3765
rect -1658 3697 -1646 3731
rect -1612 3697 -1600 3731
rect -1658 3663 -1600 3697
rect -1658 3629 -1646 3663
rect -1612 3629 -1600 3663
rect -1658 3595 -1600 3629
rect -1658 3561 -1646 3595
rect -1612 3561 -1600 3595
rect -1658 3527 -1600 3561
rect -1658 3493 -1646 3527
rect -1612 3493 -1600 3527
rect -1658 3459 -1600 3493
rect -1658 3425 -1646 3459
rect -1612 3425 -1600 3459
rect -1658 3391 -1600 3425
rect -1658 3357 -1646 3391
rect -1612 3357 -1600 3391
rect -1658 3323 -1600 3357
rect -1658 3289 -1646 3323
rect -1612 3289 -1600 3323
rect -1658 3255 -1600 3289
rect -1658 3221 -1646 3255
rect -1612 3221 -1600 3255
rect -1658 3187 -1600 3221
rect -1658 3153 -1646 3187
rect -1612 3153 -1600 3187
rect -1658 3119 -1600 3153
rect -1658 3085 -1646 3119
rect -1612 3085 -1600 3119
rect -1658 3051 -1600 3085
rect -1658 3017 -1646 3051
rect -1612 3017 -1600 3051
rect -1658 2983 -1600 3017
rect -1658 2949 -1646 2983
rect -1612 2949 -1600 2983
rect -1658 2915 -1600 2949
rect -1658 2881 -1646 2915
rect -1612 2881 -1600 2915
rect -1658 2847 -1600 2881
rect -1658 2813 -1646 2847
rect -1612 2813 -1600 2847
rect -1658 2779 -1600 2813
rect -1658 2745 -1646 2779
rect -1612 2745 -1600 2779
rect -1658 2711 -1600 2745
rect -1658 2677 -1646 2711
rect -1612 2677 -1600 2711
rect -1658 2643 -1600 2677
rect -1658 2609 -1646 2643
rect -1612 2609 -1600 2643
rect -1658 2575 -1600 2609
rect -1658 2541 -1646 2575
rect -1612 2541 -1600 2575
rect -1658 2507 -1600 2541
rect -1658 2473 -1646 2507
rect -1612 2473 -1600 2507
rect -1658 2439 -1600 2473
rect -1658 2405 -1646 2439
rect -1612 2405 -1600 2439
rect -1658 2371 -1600 2405
rect -1658 2337 -1646 2371
rect -1612 2337 -1600 2371
rect -1658 2303 -1600 2337
rect -1658 2269 -1646 2303
rect -1612 2269 -1600 2303
rect -1658 2235 -1600 2269
rect -1658 2201 -1646 2235
rect -1612 2201 -1600 2235
rect -1658 2167 -1600 2201
rect -1658 2133 -1646 2167
rect -1612 2133 -1600 2167
rect -1658 2099 -1600 2133
rect -1658 2065 -1646 2099
rect -1612 2065 -1600 2099
rect -1658 2031 -1600 2065
rect -1658 1997 -1646 2031
rect -1612 1997 -1600 2031
rect -1658 1963 -1600 1997
rect -1658 1929 -1646 1963
rect -1612 1929 -1600 1963
rect -1658 1895 -1600 1929
rect -1658 1861 -1646 1895
rect -1612 1861 -1600 1895
rect -1658 1827 -1600 1861
rect -1658 1793 -1646 1827
rect -1612 1793 -1600 1827
rect -1658 1759 -1600 1793
rect -1658 1725 -1646 1759
rect -1612 1725 -1600 1759
rect -1658 1691 -1600 1725
rect -1658 1657 -1646 1691
rect -1612 1657 -1600 1691
rect -1658 1623 -1600 1657
rect -1658 1589 -1646 1623
rect -1612 1589 -1600 1623
rect -1658 1555 -1600 1589
rect -1658 1521 -1646 1555
rect -1612 1521 -1600 1555
rect -1658 1487 -1600 1521
rect -1658 1453 -1646 1487
rect -1612 1453 -1600 1487
rect -1658 1419 -1600 1453
rect -1658 1385 -1646 1419
rect -1612 1385 -1600 1419
rect -1658 1351 -1600 1385
rect -1658 1317 -1646 1351
rect -1612 1317 -1600 1351
rect -1658 1283 -1600 1317
rect -1658 1249 -1646 1283
rect -1612 1249 -1600 1283
rect -1658 1215 -1600 1249
rect -1658 1181 -1646 1215
rect -1612 1181 -1600 1215
rect -1658 1147 -1600 1181
rect -1658 1113 -1646 1147
rect -1612 1113 -1600 1147
rect -1658 1079 -1600 1113
rect -1658 1045 -1646 1079
rect -1612 1045 -1600 1079
rect -1658 1011 -1600 1045
rect -1658 977 -1646 1011
rect -1612 977 -1600 1011
rect -1658 943 -1600 977
rect -1658 909 -1646 943
rect -1612 909 -1600 943
rect -1658 875 -1600 909
rect -1658 841 -1646 875
rect -1612 841 -1600 875
rect -1658 807 -1600 841
rect -1658 773 -1646 807
rect -1612 773 -1600 807
rect -1658 739 -1600 773
rect -1658 705 -1646 739
rect -1612 705 -1600 739
rect -1658 671 -1600 705
rect -1658 637 -1646 671
rect -1612 637 -1600 671
rect -1658 603 -1600 637
rect -1658 569 -1646 603
rect -1612 569 -1600 603
rect -1658 535 -1600 569
rect -1658 501 -1646 535
rect -1612 501 -1600 535
rect -1658 467 -1600 501
rect -1658 433 -1646 467
rect -1612 433 -1600 467
rect -1658 399 -1600 433
rect -1658 365 -1646 399
rect -1612 365 -1600 399
rect -1658 331 -1600 365
rect -1658 297 -1646 331
rect -1612 297 -1600 331
rect -1658 263 -1600 297
rect -1658 229 -1646 263
rect -1612 229 -1600 263
rect -1658 195 -1600 229
rect -1658 161 -1646 195
rect -1612 161 -1600 195
rect -1658 127 -1600 161
rect -1658 93 -1646 127
rect -1612 93 -1600 127
rect -1658 59 -1600 93
rect -1658 25 -1646 59
rect -1612 25 -1600 59
rect -1658 0 -1600 25
rect 1750 5975 1808 6000
rect 1750 5941 1762 5975
rect 1796 5941 1808 5975
rect 1750 5907 1808 5941
rect 1750 5873 1762 5907
rect 1796 5873 1808 5907
rect 1750 5839 1808 5873
rect 1750 5805 1762 5839
rect 1796 5805 1808 5839
rect 1750 5771 1808 5805
rect 1750 5737 1762 5771
rect 1796 5737 1808 5771
rect 1750 5703 1808 5737
rect 1750 5669 1762 5703
rect 1796 5669 1808 5703
rect 1750 5635 1808 5669
rect 1750 5601 1762 5635
rect 1796 5601 1808 5635
rect 1750 5567 1808 5601
rect 1750 5533 1762 5567
rect 1796 5533 1808 5567
rect 1750 5499 1808 5533
rect 1750 5465 1762 5499
rect 1796 5465 1808 5499
rect 1750 5431 1808 5465
rect 1750 5397 1762 5431
rect 1796 5397 1808 5431
rect 1750 5363 1808 5397
rect 1750 5329 1762 5363
rect 1796 5329 1808 5363
rect 1750 5295 1808 5329
rect 1750 5261 1762 5295
rect 1796 5261 1808 5295
rect 1750 5227 1808 5261
rect 1750 5193 1762 5227
rect 1796 5193 1808 5227
rect 1750 5159 1808 5193
rect 1750 5125 1762 5159
rect 1796 5125 1808 5159
rect 1750 5091 1808 5125
rect 1750 5057 1762 5091
rect 1796 5057 1808 5091
rect 1750 5023 1808 5057
rect 1750 4989 1762 5023
rect 1796 4989 1808 5023
rect 1750 4955 1808 4989
rect 1750 4921 1762 4955
rect 1796 4921 1808 4955
rect 1750 4887 1808 4921
rect 1750 4853 1762 4887
rect 1796 4853 1808 4887
rect 1750 4819 1808 4853
rect 1750 4785 1762 4819
rect 1796 4785 1808 4819
rect 1750 4751 1808 4785
rect 1750 4717 1762 4751
rect 1796 4717 1808 4751
rect 1750 4683 1808 4717
rect 1750 4649 1762 4683
rect 1796 4649 1808 4683
rect 1750 4615 1808 4649
rect 1750 4581 1762 4615
rect 1796 4581 1808 4615
rect 1750 4547 1808 4581
rect 1750 4513 1762 4547
rect 1796 4513 1808 4547
rect 1750 4479 1808 4513
rect 1750 4445 1762 4479
rect 1796 4445 1808 4479
rect 1750 4411 1808 4445
rect 1750 4377 1762 4411
rect 1796 4377 1808 4411
rect 1750 4343 1808 4377
rect 1750 4309 1762 4343
rect 1796 4309 1808 4343
rect 1750 4275 1808 4309
rect 1750 4241 1762 4275
rect 1796 4241 1808 4275
rect 1750 4207 1808 4241
rect 1750 4173 1762 4207
rect 1796 4173 1808 4207
rect 1750 4139 1808 4173
rect 1750 4105 1762 4139
rect 1796 4105 1808 4139
rect 1750 4071 1808 4105
rect 1750 4037 1762 4071
rect 1796 4037 1808 4071
rect 1750 4003 1808 4037
rect 1750 3969 1762 4003
rect 1796 3969 1808 4003
rect 1750 3935 1808 3969
rect 1750 3901 1762 3935
rect 1796 3901 1808 3935
rect 1750 3867 1808 3901
rect 1750 3833 1762 3867
rect 1796 3833 1808 3867
rect 1750 3799 1808 3833
rect 1750 3765 1762 3799
rect 1796 3765 1808 3799
rect 1750 3731 1808 3765
rect 1750 3697 1762 3731
rect 1796 3697 1808 3731
rect 1750 3663 1808 3697
rect 1750 3629 1762 3663
rect 1796 3629 1808 3663
rect 1750 3595 1808 3629
rect 1750 3561 1762 3595
rect 1796 3561 1808 3595
rect 1750 3527 1808 3561
rect 1750 3493 1762 3527
rect 1796 3493 1808 3527
rect 1750 3459 1808 3493
rect 1750 3425 1762 3459
rect 1796 3425 1808 3459
rect 1750 3391 1808 3425
rect 1750 3357 1762 3391
rect 1796 3357 1808 3391
rect 1750 3323 1808 3357
rect 1750 3289 1762 3323
rect 1796 3289 1808 3323
rect 1750 3255 1808 3289
rect 1750 3221 1762 3255
rect 1796 3221 1808 3255
rect 1750 3187 1808 3221
rect 1750 3153 1762 3187
rect 1796 3153 1808 3187
rect 1750 3119 1808 3153
rect 1750 3085 1762 3119
rect 1796 3085 1808 3119
rect 1750 3051 1808 3085
rect 1750 3017 1762 3051
rect 1796 3017 1808 3051
rect 1750 2983 1808 3017
rect 1750 2949 1762 2983
rect 1796 2949 1808 2983
rect 1750 2915 1808 2949
rect 1750 2881 1762 2915
rect 1796 2881 1808 2915
rect 1750 2847 1808 2881
rect 1750 2813 1762 2847
rect 1796 2813 1808 2847
rect 1750 2779 1808 2813
rect 1750 2745 1762 2779
rect 1796 2745 1808 2779
rect 1750 2711 1808 2745
rect 1750 2677 1762 2711
rect 1796 2677 1808 2711
rect 1750 2643 1808 2677
rect 1750 2609 1762 2643
rect 1796 2609 1808 2643
rect 1750 2575 1808 2609
rect 1750 2541 1762 2575
rect 1796 2541 1808 2575
rect 1750 2507 1808 2541
rect 1750 2473 1762 2507
rect 1796 2473 1808 2507
rect 1750 2439 1808 2473
rect 1750 2405 1762 2439
rect 1796 2405 1808 2439
rect 1750 2371 1808 2405
rect 1750 2337 1762 2371
rect 1796 2337 1808 2371
rect 1750 2303 1808 2337
rect 1750 2269 1762 2303
rect 1796 2269 1808 2303
rect 1750 2235 1808 2269
rect 1750 2201 1762 2235
rect 1796 2201 1808 2235
rect 1750 2167 1808 2201
rect 1750 2133 1762 2167
rect 1796 2133 1808 2167
rect 1750 2099 1808 2133
rect 1750 2065 1762 2099
rect 1796 2065 1808 2099
rect 1750 2031 1808 2065
rect 1750 1997 1762 2031
rect 1796 1997 1808 2031
rect 1750 1963 1808 1997
rect 1750 1929 1762 1963
rect 1796 1929 1808 1963
rect 1750 1895 1808 1929
rect 1750 1861 1762 1895
rect 1796 1861 1808 1895
rect 1750 1827 1808 1861
rect 1750 1793 1762 1827
rect 1796 1793 1808 1827
rect 1750 1759 1808 1793
rect 1750 1725 1762 1759
rect 1796 1725 1808 1759
rect 1750 1691 1808 1725
rect 1750 1657 1762 1691
rect 1796 1657 1808 1691
rect 1750 1623 1808 1657
rect 1750 1589 1762 1623
rect 1796 1589 1808 1623
rect 1750 1555 1808 1589
rect 1750 1521 1762 1555
rect 1796 1521 1808 1555
rect 1750 1487 1808 1521
rect 1750 1453 1762 1487
rect 1796 1453 1808 1487
rect 1750 1419 1808 1453
rect 1750 1385 1762 1419
rect 1796 1385 1808 1419
rect 1750 1351 1808 1385
rect 1750 1317 1762 1351
rect 1796 1317 1808 1351
rect 1750 1283 1808 1317
rect 1750 1249 1762 1283
rect 1796 1249 1808 1283
rect 1750 1215 1808 1249
rect 1750 1181 1762 1215
rect 1796 1181 1808 1215
rect 1750 1147 1808 1181
rect 1750 1113 1762 1147
rect 1796 1113 1808 1147
rect 1750 1079 1808 1113
rect 1750 1045 1762 1079
rect 1796 1045 1808 1079
rect 1750 1011 1808 1045
rect 1750 977 1762 1011
rect 1796 977 1808 1011
rect 1750 943 1808 977
rect 1750 909 1762 943
rect 1796 909 1808 943
rect 1750 875 1808 909
rect 1750 841 1762 875
rect 1796 841 1808 875
rect 1750 807 1808 841
rect 1750 773 1762 807
rect 1796 773 1808 807
rect 1750 739 1808 773
rect 1750 705 1762 739
rect 1796 705 1808 739
rect 1750 671 1808 705
rect 1750 637 1762 671
rect 1796 637 1808 671
rect 1750 603 1808 637
rect 1750 569 1762 603
rect 1796 569 1808 603
rect 1750 535 1808 569
rect 1750 501 1762 535
rect 1796 501 1808 535
rect 1750 467 1808 501
rect 1750 433 1762 467
rect 1796 433 1808 467
rect 1750 399 1808 433
rect 1750 365 1762 399
rect 1796 365 1808 399
rect 1750 331 1808 365
rect 1750 297 1762 331
rect 1796 297 1808 331
rect 1750 263 1808 297
rect 1750 229 1762 263
rect 1796 229 1808 263
rect 1750 195 1808 229
rect 1750 161 1762 195
rect 1796 161 1808 195
rect 1750 127 1808 161
rect 1750 93 1762 127
rect 1796 93 1808 127
rect 1750 59 1808 93
rect 1750 25 1762 59
rect 1796 25 1808 59
rect 1750 0 1808 25
<< mvndiffc >>
rect -1646 5941 -1612 5975
rect -1646 5873 -1612 5907
rect -1646 5805 -1612 5839
rect -1646 5737 -1612 5771
rect -1646 5669 -1612 5703
rect -1646 5601 -1612 5635
rect -1646 5533 -1612 5567
rect -1646 5465 -1612 5499
rect -1646 5397 -1612 5431
rect -1646 5329 -1612 5363
rect -1646 5261 -1612 5295
rect -1646 5193 -1612 5227
rect -1646 5125 -1612 5159
rect -1646 5057 -1612 5091
rect -1646 4989 -1612 5023
rect -1646 4921 -1612 4955
rect -1646 4853 -1612 4887
rect -1646 4785 -1612 4819
rect -1646 4717 -1612 4751
rect -1646 4649 -1612 4683
rect -1646 4581 -1612 4615
rect -1646 4513 -1612 4547
rect -1646 4445 -1612 4479
rect -1646 4377 -1612 4411
rect -1646 4309 -1612 4343
rect -1646 4241 -1612 4275
rect -1646 4173 -1612 4207
rect -1646 4105 -1612 4139
rect -1646 4037 -1612 4071
rect -1646 3969 -1612 4003
rect -1646 3901 -1612 3935
rect -1646 3833 -1612 3867
rect -1646 3765 -1612 3799
rect -1646 3697 -1612 3731
rect -1646 3629 -1612 3663
rect -1646 3561 -1612 3595
rect -1646 3493 -1612 3527
rect -1646 3425 -1612 3459
rect -1646 3357 -1612 3391
rect -1646 3289 -1612 3323
rect -1646 3221 -1612 3255
rect -1646 3153 -1612 3187
rect -1646 3085 -1612 3119
rect -1646 3017 -1612 3051
rect -1646 2949 -1612 2983
rect -1646 2881 -1612 2915
rect -1646 2813 -1612 2847
rect -1646 2745 -1612 2779
rect -1646 2677 -1612 2711
rect -1646 2609 -1612 2643
rect -1646 2541 -1612 2575
rect -1646 2473 -1612 2507
rect -1646 2405 -1612 2439
rect -1646 2337 -1612 2371
rect -1646 2269 -1612 2303
rect -1646 2201 -1612 2235
rect -1646 2133 -1612 2167
rect -1646 2065 -1612 2099
rect -1646 1997 -1612 2031
rect -1646 1929 -1612 1963
rect -1646 1861 -1612 1895
rect -1646 1793 -1612 1827
rect -1646 1725 -1612 1759
rect -1646 1657 -1612 1691
rect -1646 1589 -1612 1623
rect -1646 1521 -1612 1555
rect -1646 1453 -1612 1487
rect -1646 1385 -1612 1419
rect -1646 1317 -1612 1351
rect -1646 1249 -1612 1283
rect -1646 1181 -1612 1215
rect -1646 1113 -1612 1147
rect -1646 1045 -1612 1079
rect -1646 977 -1612 1011
rect -1646 909 -1612 943
rect -1646 841 -1612 875
rect -1646 773 -1612 807
rect -1646 705 -1612 739
rect -1646 637 -1612 671
rect -1646 569 -1612 603
rect -1646 501 -1612 535
rect -1646 433 -1612 467
rect -1646 365 -1612 399
rect -1646 297 -1612 331
rect -1646 229 -1612 263
rect -1646 161 -1612 195
rect -1646 93 -1612 127
rect -1646 25 -1612 59
rect 1762 5941 1796 5975
rect 1762 5873 1796 5907
rect 1762 5805 1796 5839
rect 1762 5737 1796 5771
rect 1762 5669 1796 5703
rect 1762 5601 1796 5635
rect 1762 5533 1796 5567
rect 1762 5465 1796 5499
rect 1762 5397 1796 5431
rect 1762 5329 1796 5363
rect 1762 5261 1796 5295
rect 1762 5193 1796 5227
rect 1762 5125 1796 5159
rect 1762 5057 1796 5091
rect 1762 4989 1796 5023
rect 1762 4921 1796 4955
rect 1762 4853 1796 4887
rect 1762 4785 1796 4819
rect 1762 4717 1796 4751
rect 1762 4649 1796 4683
rect 1762 4581 1796 4615
rect 1762 4513 1796 4547
rect 1762 4445 1796 4479
rect 1762 4377 1796 4411
rect 1762 4309 1796 4343
rect 1762 4241 1796 4275
rect 1762 4173 1796 4207
rect 1762 4105 1796 4139
rect 1762 4037 1796 4071
rect 1762 3969 1796 4003
rect 1762 3901 1796 3935
rect 1762 3833 1796 3867
rect 1762 3765 1796 3799
rect 1762 3697 1796 3731
rect 1762 3629 1796 3663
rect 1762 3561 1796 3595
rect 1762 3493 1796 3527
rect 1762 3425 1796 3459
rect 1762 3357 1796 3391
rect 1762 3289 1796 3323
rect 1762 3221 1796 3255
rect 1762 3153 1796 3187
rect 1762 3085 1796 3119
rect 1762 3017 1796 3051
rect 1762 2949 1796 2983
rect 1762 2881 1796 2915
rect 1762 2813 1796 2847
rect 1762 2745 1796 2779
rect 1762 2677 1796 2711
rect 1762 2609 1796 2643
rect 1762 2541 1796 2575
rect 1762 2473 1796 2507
rect 1762 2405 1796 2439
rect 1762 2337 1796 2371
rect 1762 2269 1796 2303
rect 1762 2201 1796 2235
rect 1762 2133 1796 2167
rect 1762 2065 1796 2099
rect 1762 1997 1796 2031
rect 1762 1929 1796 1963
rect 1762 1861 1796 1895
rect 1762 1793 1796 1827
rect 1762 1725 1796 1759
rect 1762 1657 1796 1691
rect 1762 1589 1796 1623
rect 1762 1521 1796 1555
rect 1762 1453 1796 1487
rect 1762 1385 1796 1419
rect 1762 1317 1796 1351
rect 1762 1249 1796 1283
rect 1762 1181 1796 1215
rect 1762 1113 1796 1147
rect 1762 1045 1796 1079
rect 1762 977 1796 1011
rect 1762 909 1796 943
rect 1762 841 1796 875
rect 1762 773 1796 807
rect 1762 705 1796 739
rect 1762 637 1796 671
rect 1762 569 1796 603
rect 1762 501 1796 535
rect 1762 433 1796 467
rect 1762 365 1796 399
rect 1762 297 1796 331
rect 1762 229 1796 263
rect 1762 161 1796 195
rect 1762 93 1796 127
rect 1762 25 1796 59
<< mvpsubdiff >>
rect -1840 6958 1990 6982
rect -1840 6924 -1608 6958
rect -1574 6924 -1540 6958
rect -1506 6924 -1472 6958
rect -1438 6924 -1404 6958
rect -1370 6924 -1336 6958
rect -1302 6924 -1268 6958
rect -1234 6924 -1200 6958
rect -1166 6924 -1132 6958
rect -1098 6924 -1064 6958
rect -1030 6924 -996 6958
rect -962 6924 -928 6958
rect -894 6924 -860 6958
rect -826 6924 -792 6958
rect -758 6924 -724 6958
rect -690 6924 -656 6958
rect -622 6924 -588 6958
rect -554 6924 -520 6958
rect -486 6924 -452 6958
rect -418 6924 -384 6958
rect -350 6924 -316 6958
rect -282 6924 -248 6958
rect -214 6924 -180 6958
rect -146 6924 -112 6958
rect -78 6924 -44 6958
rect -10 6924 24 6958
rect 58 6924 92 6958
rect 126 6924 160 6958
rect 194 6924 228 6958
rect 262 6924 296 6958
rect 330 6924 364 6958
rect 398 6924 432 6958
rect 466 6924 500 6958
rect 534 6924 568 6958
rect 602 6924 636 6958
rect 670 6924 704 6958
rect 738 6924 772 6958
rect 806 6924 840 6958
rect 874 6924 908 6958
rect 942 6924 976 6958
rect 1010 6924 1044 6958
rect 1078 6924 1112 6958
rect 1146 6924 1180 6958
rect 1214 6924 1248 6958
rect 1282 6924 1316 6958
rect 1350 6924 1384 6958
rect 1418 6924 1452 6958
rect 1486 6924 1520 6958
rect 1554 6924 1588 6958
rect 1622 6924 1656 6958
rect 1690 6924 1724 6958
rect 1758 6924 1990 6958
rect -1840 6900 1990 6924
rect -1840 6825 -1758 6900
rect -1840 6791 -1816 6825
rect -1782 6791 -1758 6825
rect 1908 6825 1990 6900
rect -1840 6757 -1758 6791
rect -1840 6723 -1816 6757
rect -1782 6723 -1758 6757
rect -1840 6689 -1758 6723
rect -1840 6655 -1816 6689
rect -1782 6655 -1758 6689
rect -1840 6621 -1758 6655
rect -1840 6587 -1816 6621
rect -1782 6587 -1758 6621
rect -1840 6553 -1758 6587
rect -1840 6519 -1816 6553
rect -1782 6519 -1758 6553
rect -1840 6485 -1758 6519
rect -1840 6451 -1816 6485
rect -1782 6451 -1758 6485
rect -1840 6417 -1758 6451
rect -1840 6383 -1816 6417
rect -1782 6383 -1758 6417
rect -1840 6349 -1758 6383
rect -1840 6315 -1816 6349
rect -1782 6315 -1758 6349
rect -1840 6281 -1758 6315
rect -1840 6247 -1816 6281
rect -1782 6247 -1758 6281
rect -1840 6213 -1758 6247
rect -1840 6179 -1816 6213
rect -1782 6179 -1758 6213
rect -1840 6145 -1758 6179
rect -1840 6111 -1816 6145
rect -1782 6111 -1758 6145
rect -1840 6077 -1758 6111
rect -1840 6043 -1816 6077
rect -1782 6043 -1758 6077
rect -1840 6009 -1758 6043
rect -1840 5975 -1816 6009
rect -1782 5975 -1758 6009
rect 1908 6791 1932 6825
rect 1966 6791 1990 6825
rect 1908 6757 1990 6791
rect 1908 6723 1932 6757
rect 1966 6723 1990 6757
rect 1908 6689 1990 6723
rect 1908 6655 1932 6689
rect 1966 6655 1990 6689
rect 1908 6621 1990 6655
rect 1908 6587 1932 6621
rect 1966 6587 1990 6621
rect 1908 6553 1990 6587
rect 1908 6519 1932 6553
rect 1966 6519 1990 6553
rect 1908 6485 1990 6519
rect 1908 6451 1932 6485
rect 1966 6451 1990 6485
rect 1908 6417 1990 6451
rect 1908 6383 1932 6417
rect 1966 6383 1990 6417
rect 1908 6349 1990 6383
rect 1908 6315 1932 6349
rect 1966 6315 1990 6349
rect 1908 6281 1990 6315
rect 1908 6247 1932 6281
rect 1966 6247 1990 6281
rect 1908 6213 1990 6247
rect 1908 6179 1932 6213
rect 1966 6179 1990 6213
rect 1908 6145 1990 6179
rect 1908 6111 1932 6145
rect 1966 6111 1990 6145
rect 1908 6077 1990 6111
rect 1908 6043 1932 6077
rect 1966 6043 1990 6077
rect 1908 6009 1990 6043
rect -1840 5941 -1758 5975
rect -1840 5907 -1816 5941
rect -1782 5907 -1758 5941
rect -1840 5873 -1758 5907
rect -1840 5839 -1816 5873
rect -1782 5839 -1758 5873
rect -1840 5805 -1758 5839
rect -1840 5771 -1816 5805
rect -1782 5771 -1758 5805
rect -1840 5737 -1758 5771
rect -1840 5703 -1816 5737
rect -1782 5703 -1758 5737
rect -1840 5669 -1758 5703
rect -1840 5635 -1816 5669
rect -1782 5635 -1758 5669
rect -1840 5601 -1758 5635
rect -1840 5567 -1816 5601
rect -1782 5567 -1758 5601
rect -1840 5533 -1758 5567
rect -1840 5499 -1816 5533
rect -1782 5499 -1758 5533
rect -1840 5465 -1758 5499
rect -1840 5431 -1816 5465
rect -1782 5431 -1758 5465
rect -1840 5397 -1758 5431
rect -1840 5363 -1816 5397
rect -1782 5363 -1758 5397
rect -1840 5329 -1758 5363
rect -1840 5295 -1816 5329
rect -1782 5295 -1758 5329
rect -1840 5261 -1758 5295
rect -1840 5227 -1816 5261
rect -1782 5227 -1758 5261
rect -1840 5193 -1758 5227
rect -1840 5159 -1816 5193
rect -1782 5159 -1758 5193
rect -1840 5125 -1758 5159
rect -1840 5091 -1816 5125
rect -1782 5091 -1758 5125
rect -1840 5057 -1758 5091
rect -1840 5023 -1816 5057
rect -1782 5023 -1758 5057
rect -1840 4989 -1758 5023
rect -1840 4955 -1816 4989
rect -1782 4955 -1758 4989
rect -1840 4921 -1758 4955
rect -1840 4887 -1816 4921
rect -1782 4887 -1758 4921
rect -1840 4853 -1758 4887
rect -1840 4819 -1816 4853
rect -1782 4819 -1758 4853
rect -1840 4785 -1758 4819
rect -1840 4751 -1816 4785
rect -1782 4751 -1758 4785
rect -1840 4717 -1758 4751
rect -1840 4683 -1816 4717
rect -1782 4683 -1758 4717
rect -1840 4649 -1758 4683
rect -1840 4615 -1816 4649
rect -1782 4615 -1758 4649
rect -1840 4581 -1758 4615
rect -1840 4547 -1816 4581
rect -1782 4547 -1758 4581
rect -1840 4513 -1758 4547
rect -1840 4479 -1816 4513
rect -1782 4479 -1758 4513
rect -1840 4445 -1758 4479
rect -1840 4411 -1816 4445
rect -1782 4411 -1758 4445
rect -1840 4377 -1758 4411
rect -1840 4343 -1816 4377
rect -1782 4343 -1758 4377
rect -1840 4309 -1758 4343
rect -1840 4275 -1816 4309
rect -1782 4275 -1758 4309
rect -1840 4241 -1758 4275
rect -1840 4207 -1816 4241
rect -1782 4207 -1758 4241
rect -1840 4173 -1758 4207
rect -1840 4139 -1816 4173
rect -1782 4139 -1758 4173
rect -1840 4105 -1758 4139
rect -1840 4071 -1816 4105
rect -1782 4071 -1758 4105
rect -1840 4037 -1758 4071
rect -1840 4003 -1816 4037
rect -1782 4003 -1758 4037
rect -1840 3969 -1758 4003
rect -1840 3935 -1816 3969
rect -1782 3935 -1758 3969
rect -1840 3901 -1758 3935
rect -1840 3867 -1816 3901
rect -1782 3867 -1758 3901
rect -1840 3833 -1758 3867
rect -1840 3799 -1816 3833
rect -1782 3799 -1758 3833
rect -1840 3765 -1758 3799
rect -1840 3731 -1816 3765
rect -1782 3731 -1758 3765
rect -1840 3697 -1758 3731
rect -1840 3663 -1816 3697
rect -1782 3663 -1758 3697
rect -1840 3629 -1758 3663
rect -1840 3595 -1816 3629
rect -1782 3595 -1758 3629
rect -1840 3561 -1758 3595
rect -1840 3527 -1816 3561
rect -1782 3527 -1758 3561
rect -1840 3493 -1758 3527
rect -1840 3459 -1816 3493
rect -1782 3459 -1758 3493
rect -1840 3425 -1758 3459
rect -1840 3391 -1816 3425
rect -1782 3391 -1758 3425
rect -1840 3357 -1758 3391
rect -1840 3323 -1816 3357
rect -1782 3323 -1758 3357
rect -1840 3289 -1758 3323
rect -1840 3255 -1816 3289
rect -1782 3255 -1758 3289
rect -1840 3221 -1758 3255
rect -1840 3187 -1816 3221
rect -1782 3187 -1758 3221
rect -1840 3153 -1758 3187
rect -1840 3119 -1816 3153
rect -1782 3119 -1758 3153
rect -1840 3085 -1758 3119
rect -1840 3051 -1816 3085
rect -1782 3051 -1758 3085
rect -1840 3017 -1758 3051
rect -1840 2983 -1816 3017
rect -1782 2983 -1758 3017
rect -1840 2949 -1758 2983
rect -1840 2915 -1816 2949
rect -1782 2915 -1758 2949
rect -1840 2881 -1758 2915
rect -1840 2847 -1816 2881
rect -1782 2847 -1758 2881
rect -1840 2813 -1758 2847
rect -1840 2779 -1816 2813
rect -1782 2779 -1758 2813
rect -1840 2745 -1758 2779
rect -1840 2711 -1816 2745
rect -1782 2711 -1758 2745
rect -1840 2677 -1758 2711
rect -1840 2643 -1816 2677
rect -1782 2643 -1758 2677
rect -1840 2609 -1758 2643
rect -1840 2575 -1816 2609
rect -1782 2575 -1758 2609
rect -1840 2541 -1758 2575
rect -1840 2507 -1816 2541
rect -1782 2507 -1758 2541
rect -1840 2473 -1758 2507
rect -1840 2439 -1816 2473
rect -1782 2439 -1758 2473
rect -1840 2405 -1758 2439
rect -1840 2371 -1816 2405
rect -1782 2371 -1758 2405
rect -1840 2337 -1758 2371
rect -1840 2303 -1816 2337
rect -1782 2303 -1758 2337
rect -1840 2269 -1758 2303
rect -1840 2235 -1816 2269
rect -1782 2235 -1758 2269
rect -1840 2201 -1758 2235
rect -1840 2167 -1816 2201
rect -1782 2167 -1758 2201
rect -1840 2133 -1758 2167
rect -1840 2099 -1816 2133
rect -1782 2099 -1758 2133
rect -1840 2065 -1758 2099
rect -1840 2031 -1816 2065
rect -1782 2031 -1758 2065
rect -1840 1997 -1758 2031
rect -1840 1963 -1816 1997
rect -1782 1963 -1758 1997
rect -1840 1929 -1758 1963
rect -1840 1895 -1816 1929
rect -1782 1895 -1758 1929
rect -1840 1861 -1758 1895
rect -1840 1827 -1816 1861
rect -1782 1827 -1758 1861
rect -1840 1793 -1758 1827
rect -1840 1759 -1816 1793
rect -1782 1759 -1758 1793
rect -1840 1725 -1758 1759
rect -1840 1691 -1816 1725
rect -1782 1691 -1758 1725
rect -1840 1657 -1758 1691
rect -1840 1623 -1816 1657
rect -1782 1623 -1758 1657
rect -1840 1589 -1758 1623
rect -1840 1555 -1816 1589
rect -1782 1555 -1758 1589
rect -1840 1521 -1758 1555
rect -1840 1487 -1816 1521
rect -1782 1487 -1758 1521
rect -1840 1453 -1758 1487
rect -1840 1419 -1816 1453
rect -1782 1419 -1758 1453
rect -1840 1385 -1758 1419
rect -1840 1351 -1816 1385
rect -1782 1351 -1758 1385
rect -1840 1317 -1758 1351
rect -1840 1283 -1816 1317
rect -1782 1283 -1758 1317
rect -1840 1249 -1758 1283
rect -1840 1215 -1816 1249
rect -1782 1215 -1758 1249
rect -1840 1181 -1758 1215
rect -1840 1147 -1816 1181
rect -1782 1147 -1758 1181
rect -1840 1113 -1758 1147
rect -1840 1079 -1816 1113
rect -1782 1079 -1758 1113
rect -1840 1045 -1758 1079
rect -1840 1011 -1816 1045
rect -1782 1011 -1758 1045
rect -1840 977 -1758 1011
rect -1840 943 -1816 977
rect -1782 943 -1758 977
rect -1840 909 -1758 943
rect -1840 875 -1816 909
rect -1782 875 -1758 909
rect -1840 841 -1758 875
rect -1840 807 -1816 841
rect -1782 807 -1758 841
rect -1840 773 -1758 807
rect -1840 739 -1816 773
rect -1782 739 -1758 773
rect -1840 705 -1758 739
rect -1840 671 -1816 705
rect -1782 671 -1758 705
rect -1840 637 -1758 671
rect -1840 603 -1816 637
rect -1782 603 -1758 637
rect -1840 569 -1758 603
rect -1840 535 -1816 569
rect -1782 535 -1758 569
rect -1840 501 -1758 535
rect -1840 467 -1816 501
rect -1782 467 -1758 501
rect -1840 433 -1758 467
rect -1840 399 -1816 433
rect -1782 399 -1758 433
rect -1840 365 -1758 399
rect -1840 331 -1816 365
rect -1782 331 -1758 365
rect -1840 297 -1758 331
rect -1840 263 -1816 297
rect -1782 263 -1758 297
rect -1840 229 -1758 263
rect -1840 195 -1816 229
rect -1782 195 -1758 229
rect -1840 161 -1758 195
rect -1840 127 -1816 161
rect -1782 127 -1758 161
rect -1840 93 -1758 127
rect -1840 59 -1816 93
rect -1782 59 -1758 93
rect -1840 25 -1758 59
rect -1840 -9 -1816 25
rect -1782 -9 -1758 25
rect 1908 5975 1932 6009
rect 1966 5975 1990 6009
rect 1908 5941 1990 5975
rect 1908 5907 1932 5941
rect 1966 5907 1990 5941
rect 1908 5873 1990 5907
rect 1908 5839 1932 5873
rect 1966 5839 1990 5873
rect 1908 5805 1990 5839
rect 1908 5771 1932 5805
rect 1966 5771 1990 5805
rect 1908 5737 1990 5771
rect 1908 5703 1932 5737
rect 1966 5703 1990 5737
rect 1908 5669 1990 5703
rect 1908 5635 1932 5669
rect 1966 5635 1990 5669
rect 1908 5601 1990 5635
rect 1908 5567 1932 5601
rect 1966 5567 1990 5601
rect 1908 5533 1990 5567
rect 1908 5499 1932 5533
rect 1966 5499 1990 5533
rect 1908 5465 1990 5499
rect 1908 5431 1932 5465
rect 1966 5431 1990 5465
rect 1908 5397 1990 5431
rect 1908 5363 1932 5397
rect 1966 5363 1990 5397
rect 1908 5329 1990 5363
rect 1908 5295 1932 5329
rect 1966 5295 1990 5329
rect 1908 5261 1990 5295
rect 1908 5227 1932 5261
rect 1966 5227 1990 5261
rect 1908 5193 1990 5227
rect 1908 5159 1932 5193
rect 1966 5159 1990 5193
rect 1908 5125 1990 5159
rect 1908 5091 1932 5125
rect 1966 5091 1990 5125
rect 1908 5057 1990 5091
rect 1908 5023 1932 5057
rect 1966 5023 1990 5057
rect 1908 4989 1990 5023
rect 1908 4955 1932 4989
rect 1966 4955 1990 4989
rect 1908 4921 1990 4955
rect 1908 4887 1932 4921
rect 1966 4887 1990 4921
rect 1908 4853 1990 4887
rect 1908 4819 1932 4853
rect 1966 4819 1990 4853
rect 1908 4785 1990 4819
rect 1908 4751 1932 4785
rect 1966 4751 1990 4785
rect 1908 4717 1990 4751
rect 1908 4683 1932 4717
rect 1966 4683 1990 4717
rect 1908 4649 1990 4683
rect 1908 4615 1932 4649
rect 1966 4615 1990 4649
rect 1908 4581 1990 4615
rect 1908 4547 1932 4581
rect 1966 4547 1990 4581
rect 1908 4513 1990 4547
rect 1908 4479 1932 4513
rect 1966 4479 1990 4513
rect 1908 4445 1990 4479
rect 1908 4411 1932 4445
rect 1966 4411 1990 4445
rect 1908 4377 1990 4411
rect 1908 4343 1932 4377
rect 1966 4343 1990 4377
rect 1908 4309 1990 4343
rect 1908 4275 1932 4309
rect 1966 4275 1990 4309
rect 1908 4241 1990 4275
rect 1908 4207 1932 4241
rect 1966 4207 1990 4241
rect 1908 4173 1990 4207
rect 1908 4139 1932 4173
rect 1966 4139 1990 4173
rect 1908 4105 1990 4139
rect 1908 4071 1932 4105
rect 1966 4071 1990 4105
rect 1908 4037 1990 4071
rect 1908 4003 1932 4037
rect 1966 4003 1990 4037
rect 1908 3969 1990 4003
rect 1908 3935 1932 3969
rect 1966 3935 1990 3969
rect 1908 3901 1990 3935
rect 1908 3867 1932 3901
rect 1966 3867 1990 3901
rect 1908 3833 1990 3867
rect 1908 3799 1932 3833
rect 1966 3799 1990 3833
rect 1908 3765 1990 3799
rect 1908 3731 1932 3765
rect 1966 3731 1990 3765
rect 1908 3697 1990 3731
rect 1908 3663 1932 3697
rect 1966 3663 1990 3697
rect 1908 3629 1990 3663
rect 1908 3595 1932 3629
rect 1966 3595 1990 3629
rect 1908 3561 1990 3595
rect 1908 3527 1932 3561
rect 1966 3527 1990 3561
rect 1908 3493 1990 3527
rect 1908 3459 1932 3493
rect 1966 3459 1990 3493
rect 1908 3425 1990 3459
rect 1908 3391 1932 3425
rect 1966 3391 1990 3425
rect 1908 3357 1990 3391
rect 1908 3323 1932 3357
rect 1966 3323 1990 3357
rect 1908 3289 1990 3323
rect 1908 3255 1932 3289
rect 1966 3255 1990 3289
rect 1908 3221 1990 3255
rect 1908 3187 1932 3221
rect 1966 3187 1990 3221
rect 1908 3153 1990 3187
rect 1908 3119 1932 3153
rect 1966 3119 1990 3153
rect 1908 3085 1990 3119
rect 1908 3051 1932 3085
rect 1966 3051 1990 3085
rect 1908 3017 1990 3051
rect 1908 2983 1932 3017
rect 1966 2983 1990 3017
rect 1908 2949 1990 2983
rect 1908 2915 1932 2949
rect 1966 2915 1990 2949
rect 1908 2881 1990 2915
rect 1908 2847 1932 2881
rect 1966 2847 1990 2881
rect 1908 2813 1990 2847
rect 1908 2779 1932 2813
rect 1966 2779 1990 2813
rect 1908 2745 1990 2779
rect 1908 2711 1932 2745
rect 1966 2711 1990 2745
rect 1908 2677 1990 2711
rect 1908 2643 1932 2677
rect 1966 2643 1990 2677
rect 1908 2609 1990 2643
rect 1908 2575 1932 2609
rect 1966 2575 1990 2609
rect 1908 2541 1990 2575
rect 1908 2507 1932 2541
rect 1966 2507 1990 2541
rect 1908 2473 1990 2507
rect 1908 2439 1932 2473
rect 1966 2439 1990 2473
rect 1908 2405 1990 2439
rect 1908 2371 1932 2405
rect 1966 2371 1990 2405
rect 1908 2337 1990 2371
rect 1908 2303 1932 2337
rect 1966 2303 1990 2337
rect 1908 2269 1990 2303
rect 1908 2235 1932 2269
rect 1966 2235 1990 2269
rect 1908 2201 1990 2235
rect 1908 2167 1932 2201
rect 1966 2167 1990 2201
rect 1908 2133 1990 2167
rect 1908 2099 1932 2133
rect 1966 2099 1990 2133
rect 1908 2065 1990 2099
rect 1908 2031 1932 2065
rect 1966 2031 1990 2065
rect 1908 1997 1990 2031
rect 1908 1963 1932 1997
rect 1966 1963 1990 1997
rect 1908 1929 1990 1963
rect 1908 1895 1932 1929
rect 1966 1895 1990 1929
rect 1908 1861 1990 1895
rect 1908 1827 1932 1861
rect 1966 1827 1990 1861
rect 1908 1793 1990 1827
rect 1908 1759 1932 1793
rect 1966 1759 1990 1793
rect 1908 1725 1990 1759
rect 1908 1691 1932 1725
rect 1966 1691 1990 1725
rect 1908 1657 1990 1691
rect 1908 1623 1932 1657
rect 1966 1623 1990 1657
rect 1908 1589 1990 1623
rect 1908 1555 1932 1589
rect 1966 1555 1990 1589
rect 1908 1521 1990 1555
rect 1908 1487 1932 1521
rect 1966 1487 1990 1521
rect 1908 1453 1990 1487
rect 1908 1419 1932 1453
rect 1966 1419 1990 1453
rect 1908 1385 1990 1419
rect 1908 1351 1932 1385
rect 1966 1351 1990 1385
rect 1908 1317 1990 1351
rect 1908 1283 1932 1317
rect 1966 1283 1990 1317
rect 1908 1249 1990 1283
rect 1908 1215 1932 1249
rect 1966 1215 1990 1249
rect 1908 1181 1990 1215
rect 1908 1147 1932 1181
rect 1966 1147 1990 1181
rect 1908 1113 1990 1147
rect 1908 1079 1932 1113
rect 1966 1079 1990 1113
rect 1908 1045 1990 1079
rect 1908 1011 1932 1045
rect 1966 1011 1990 1045
rect 1908 977 1990 1011
rect 1908 943 1932 977
rect 1966 943 1990 977
rect 1908 909 1990 943
rect 1908 875 1932 909
rect 1966 875 1990 909
rect 1908 841 1990 875
rect 1908 807 1932 841
rect 1966 807 1990 841
rect 1908 773 1990 807
rect 1908 739 1932 773
rect 1966 739 1990 773
rect 1908 705 1990 739
rect 1908 671 1932 705
rect 1966 671 1990 705
rect 1908 637 1990 671
rect 1908 603 1932 637
rect 1966 603 1990 637
rect 1908 569 1990 603
rect 1908 535 1932 569
rect 1966 535 1990 569
rect 1908 501 1990 535
rect 1908 467 1932 501
rect 1966 467 1990 501
rect 1908 433 1990 467
rect 1908 399 1932 433
rect 1966 399 1990 433
rect 1908 365 1990 399
rect 1908 331 1932 365
rect 1966 331 1990 365
rect 1908 297 1990 331
rect 1908 263 1932 297
rect 1966 263 1990 297
rect 1908 229 1990 263
rect 1908 195 1932 229
rect 1966 195 1990 229
rect 1908 161 1990 195
rect 1908 127 1932 161
rect 1966 127 1990 161
rect 1908 93 1990 127
rect 1908 59 1932 93
rect 1966 59 1990 93
rect 1908 25 1990 59
rect -1840 -43 -1758 -9
rect -1840 -77 -1816 -43
rect -1782 -77 -1758 -43
rect -1840 -111 -1758 -77
rect -1840 -145 -1816 -111
rect -1782 -145 -1758 -111
rect -1840 -179 -1758 -145
rect -1840 -213 -1816 -179
rect -1782 -213 -1758 -179
rect -1840 -247 -1758 -213
rect -1840 -281 -1816 -247
rect -1782 -281 -1758 -247
rect -1840 -315 -1758 -281
rect -1840 -349 -1816 -315
rect -1782 -349 -1758 -315
rect -1840 -383 -1758 -349
rect -1840 -417 -1816 -383
rect -1782 -417 -1758 -383
rect -1840 -451 -1758 -417
rect -1840 -485 -1816 -451
rect -1782 -485 -1758 -451
rect -1840 -519 -1758 -485
rect -1840 -553 -1816 -519
rect -1782 -553 -1758 -519
rect -1840 -587 -1758 -553
rect -1840 -621 -1816 -587
rect -1782 -621 -1758 -587
rect -1840 -655 -1758 -621
rect -1840 -689 -1816 -655
rect -1782 -689 -1758 -655
rect -1840 -723 -1758 -689
rect -1840 -757 -1816 -723
rect -1782 -757 -1758 -723
rect -1840 -791 -1758 -757
rect -1840 -825 -1816 -791
rect -1782 -825 -1758 -791
rect 1908 -9 1932 25
rect 1966 -9 1990 25
rect 1908 -43 1990 -9
rect 1908 -77 1932 -43
rect 1966 -77 1990 -43
rect 1908 -111 1990 -77
rect 1908 -145 1932 -111
rect 1966 -145 1990 -111
rect 1908 -179 1990 -145
rect 1908 -213 1932 -179
rect 1966 -213 1990 -179
rect 1908 -247 1990 -213
rect 1908 -281 1932 -247
rect 1966 -281 1990 -247
rect 1908 -315 1990 -281
rect 1908 -349 1932 -315
rect 1966 -349 1990 -315
rect 1908 -383 1990 -349
rect 1908 -417 1932 -383
rect 1966 -417 1990 -383
rect 1908 -451 1990 -417
rect 1908 -485 1932 -451
rect 1966 -485 1990 -451
rect 1908 -519 1990 -485
rect 1908 -553 1932 -519
rect 1966 -553 1990 -519
rect 1908 -587 1990 -553
rect 1908 -621 1932 -587
rect 1966 -621 1990 -587
rect 1908 -655 1990 -621
rect 1908 -689 1932 -655
rect 1966 -689 1990 -655
rect 1908 -723 1990 -689
rect 1908 -757 1932 -723
rect 1966 -757 1990 -723
rect 1908 -791 1990 -757
rect -1840 -900 -1758 -825
rect 1908 -825 1932 -791
rect 1966 -825 1990 -791
rect 1908 -900 1990 -825
rect -1840 -924 1990 -900
rect -1840 -958 -1608 -924
rect -1574 -958 -1540 -924
rect -1506 -958 -1472 -924
rect -1438 -958 -1404 -924
rect -1370 -958 -1336 -924
rect -1302 -958 -1268 -924
rect -1234 -958 -1200 -924
rect -1166 -958 -1132 -924
rect -1098 -958 -1064 -924
rect -1030 -958 -996 -924
rect -962 -958 -928 -924
rect -894 -958 -860 -924
rect -826 -958 -792 -924
rect -758 -958 -724 -924
rect -690 -958 -656 -924
rect -622 -958 -588 -924
rect -554 -958 -520 -924
rect -486 -958 -452 -924
rect -418 -958 -384 -924
rect -350 -958 -316 -924
rect -282 -958 -248 -924
rect -214 -958 -180 -924
rect -146 -958 -112 -924
rect -78 -958 -44 -924
rect -10 -958 24 -924
rect 58 -958 92 -924
rect 126 -958 160 -924
rect 194 -958 228 -924
rect 262 -958 296 -924
rect 330 -958 364 -924
rect 398 -958 432 -924
rect 466 -958 500 -924
rect 534 -958 568 -924
rect 602 -958 636 -924
rect 670 -958 704 -924
rect 738 -958 772 -924
rect 806 -958 840 -924
rect 874 -958 908 -924
rect 942 -958 976 -924
rect 1010 -958 1044 -924
rect 1078 -958 1112 -924
rect 1146 -958 1180 -924
rect 1214 -958 1248 -924
rect 1282 -958 1316 -924
rect 1350 -958 1384 -924
rect 1418 -958 1452 -924
rect 1486 -958 1520 -924
rect 1554 -958 1588 -924
rect 1622 -958 1656 -924
rect 1690 -958 1724 -924
rect 1758 -958 1990 -924
rect -1840 -982 1990 -958
<< mvnsubdiff >>
tri 0 5970 30 6000 se
rect 30 5970 120 6000
tri 120 5970 150 6000 sw
rect 0 5941 150 5970
rect 0 59 24 5941
rect 126 59 150 5941
rect 0 30 150 59
tri 0 0 30 30 ne
rect 30 0 120 30
tri 120 0 150 30 nw
<< mvpsubdiffcont >>
rect -1608 6924 -1574 6958
rect -1540 6924 -1506 6958
rect -1472 6924 -1438 6958
rect -1404 6924 -1370 6958
rect -1336 6924 -1302 6958
rect -1268 6924 -1234 6958
rect -1200 6924 -1166 6958
rect -1132 6924 -1098 6958
rect -1064 6924 -1030 6958
rect -996 6924 -962 6958
rect -928 6924 -894 6958
rect -860 6924 -826 6958
rect -792 6924 -758 6958
rect -724 6924 -690 6958
rect -656 6924 -622 6958
rect -588 6924 -554 6958
rect -520 6924 -486 6958
rect -452 6924 -418 6958
rect -384 6924 -350 6958
rect -316 6924 -282 6958
rect -248 6924 -214 6958
rect -180 6924 -146 6958
rect -112 6924 -78 6958
rect -44 6924 -10 6958
rect 24 6924 58 6958
rect 92 6924 126 6958
rect 160 6924 194 6958
rect 228 6924 262 6958
rect 296 6924 330 6958
rect 364 6924 398 6958
rect 432 6924 466 6958
rect 500 6924 534 6958
rect 568 6924 602 6958
rect 636 6924 670 6958
rect 704 6924 738 6958
rect 772 6924 806 6958
rect 840 6924 874 6958
rect 908 6924 942 6958
rect 976 6924 1010 6958
rect 1044 6924 1078 6958
rect 1112 6924 1146 6958
rect 1180 6924 1214 6958
rect 1248 6924 1282 6958
rect 1316 6924 1350 6958
rect 1384 6924 1418 6958
rect 1452 6924 1486 6958
rect 1520 6924 1554 6958
rect 1588 6924 1622 6958
rect 1656 6924 1690 6958
rect 1724 6924 1758 6958
rect -1816 6791 -1782 6825
rect -1816 6723 -1782 6757
rect -1816 6655 -1782 6689
rect -1816 6587 -1782 6621
rect -1816 6519 -1782 6553
rect -1816 6451 -1782 6485
rect -1816 6383 -1782 6417
rect -1816 6315 -1782 6349
rect -1816 6247 -1782 6281
rect -1816 6179 -1782 6213
rect -1816 6111 -1782 6145
rect -1816 6043 -1782 6077
rect -1816 5975 -1782 6009
rect 1932 6791 1966 6825
rect 1932 6723 1966 6757
rect 1932 6655 1966 6689
rect 1932 6587 1966 6621
rect 1932 6519 1966 6553
rect 1932 6451 1966 6485
rect 1932 6383 1966 6417
rect 1932 6315 1966 6349
rect 1932 6247 1966 6281
rect 1932 6179 1966 6213
rect 1932 6111 1966 6145
rect 1932 6043 1966 6077
rect -1816 5907 -1782 5941
rect -1816 5839 -1782 5873
rect -1816 5771 -1782 5805
rect -1816 5703 -1782 5737
rect -1816 5635 -1782 5669
rect -1816 5567 -1782 5601
rect -1816 5499 -1782 5533
rect -1816 5431 -1782 5465
rect -1816 5363 -1782 5397
rect -1816 5295 -1782 5329
rect -1816 5227 -1782 5261
rect -1816 5159 -1782 5193
rect -1816 5091 -1782 5125
rect -1816 5023 -1782 5057
rect -1816 4955 -1782 4989
rect -1816 4887 -1782 4921
rect -1816 4819 -1782 4853
rect -1816 4751 -1782 4785
rect -1816 4683 -1782 4717
rect -1816 4615 -1782 4649
rect -1816 4547 -1782 4581
rect -1816 4479 -1782 4513
rect -1816 4411 -1782 4445
rect -1816 4343 -1782 4377
rect -1816 4275 -1782 4309
rect -1816 4207 -1782 4241
rect -1816 4139 -1782 4173
rect -1816 4071 -1782 4105
rect -1816 4003 -1782 4037
rect -1816 3935 -1782 3969
rect -1816 3867 -1782 3901
rect -1816 3799 -1782 3833
rect -1816 3731 -1782 3765
rect -1816 3663 -1782 3697
rect -1816 3595 -1782 3629
rect -1816 3527 -1782 3561
rect -1816 3459 -1782 3493
rect -1816 3391 -1782 3425
rect -1816 3323 -1782 3357
rect -1816 3255 -1782 3289
rect -1816 3187 -1782 3221
rect -1816 3119 -1782 3153
rect -1816 3051 -1782 3085
rect -1816 2983 -1782 3017
rect -1816 2915 -1782 2949
rect -1816 2847 -1782 2881
rect -1816 2779 -1782 2813
rect -1816 2711 -1782 2745
rect -1816 2643 -1782 2677
rect -1816 2575 -1782 2609
rect -1816 2507 -1782 2541
rect -1816 2439 -1782 2473
rect -1816 2371 -1782 2405
rect -1816 2303 -1782 2337
rect -1816 2235 -1782 2269
rect -1816 2167 -1782 2201
rect -1816 2099 -1782 2133
rect -1816 2031 -1782 2065
rect -1816 1963 -1782 1997
rect -1816 1895 -1782 1929
rect -1816 1827 -1782 1861
rect -1816 1759 -1782 1793
rect -1816 1691 -1782 1725
rect -1816 1623 -1782 1657
rect -1816 1555 -1782 1589
rect -1816 1487 -1782 1521
rect -1816 1419 -1782 1453
rect -1816 1351 -1782 1385
rect -1816 1283 -1782 1317
rect -1816 1215 -1782 1249
rect -1816 1147 -1782 1181
rect -1816 1079 -1782 1113
rect -1816 1011 -1782 1045
rect -1816 943 -1782 977
rect -1816 875 -1782 909
rect -1816 807 -1782 841
rect -1816 739 -1782 773
rect -1816 671 -1782 705
rect -1816 603 -1782 637
rect -1816 535 -1782 569
rect -1816 467 -1782 501
rect -1816 399 -1782 433
rect -1816 331 -1782 365
rect -1816 263 -1782 297
rect -1816 195 -1782 229
rect -1816 127 -1782 161
rect -1816 59 -1782 93
rect -1816 -9 -1782 25
rect 1932 5975 1966 6009
rect 1932 5907 1966 5941
rect 1932 5839 1966 5873
rect 1932 5771 1966 5805
rect 1932 5703 1966 5737
rect 1932 5635 1966 5669
rect 1932 5567 1966 5601
rect 1932 5499 1966 5533
rect 1932 5431 1966 5465
rect 1932 5363 1966 5397
rect 1932 5295 1966 5329
rect 1932 5227 1966 5261
rect 1932 5159 1966 5193
rect 1932 5091 1966 5125
rect 1932 5023 1966 5057
rect 1932 4955 1966 4989
rect 1932 4887 1966 4921
rect 1932 4819 1966 4853
rect 1932 4751 1966 4785
rect 1932 4683 1966 4717
rect 1932 4615 1966 4649
rect 1932 4547 1966 4581
rect 1932 4479 1966 4513
rect 1932 4411 1966 4445
rect 1932 4343 1966 4377
rect 1932 4275 1966 4309
rect 1932 4207 1966 4241
rect 1932 4139 1966 4173
rect 1932 4071 1966 4105
rect 1932 4003 1966 4037
rect 1932 3935 1966 3969
rect 1932 3867 1966 3901
rect 1932 3799 1966 3833
rect 1932 3731 1966 3765
rect 1932 3663 1966 3697
rect 1932 3595 1966 3629
rect 1932 3527 1966 3561
rect 1932 3459 1966 3493
rect 1932 3391 1966 3425
rect 1932 3323 1966 3357
rect 1932 3255 1966 3289
rect 1932 3187 1966 3221
rect 1932 3119 1966 3153
rect 1932 3051 1966 3085
rect 1932 2983 1966 3017
rect 1932 2915 1966 2949
rect 1932 2847 1966 2881
rect 1932 2779 1966 2813
rect 1932 2711 1966 2745
rect 1932 2643 1966 2677
rect 1932 2575 1966 2609
rect 1932 2507 1966 2541
rect 1932 2439 1966 2473
rect 1932 2371 1966 2405
rect 1932 2303 1966 2337
rect 1932 2235 1966 2269
rect 1932 2167 1966 2201
rect 1932 2099 1966 2133
rect 1932 2031 1966 2065
rect 1932 1963 1966 1997
rect 1932 1895 1966 1929
rect 1932 1827 1966 1861
rect 1932 1759 1966 1793
rect 1932 1691 1966 1725
rect 1932 1623 1966 1657
rect 1932 1555 1966 1589
rect 1932 1487 1966 1521
rect 1932 1419 1966 1453
rect 1932 1351 1966 1385
rect 1932 1283 1966 1317
rect 1932 1215 1966 1249
rect 1932 1147 1966 1181
rect 1932 1079 1966 1113
rect 1932 1011 1966 1045
rect 1932 943 1966 977
rect 1932 875 1966 909
rect 1932 807 1966 841
rect 1932 739 1966 773
rect 1932 671 1966 705
rect 1932 603 1966 637
rect 1932 535 1966 569
rect 1932 467 1966 501
rect 1932 399 1966 433
rect 1932 331 1966 365
rect 1932 263 1966 297
rect 1932 195 1966 229
rect 1932 127 1966 161
rect 1932 59 1966 93
rect -1816 -77 -1782 -43
rect -1816 -145 -1782 -111
rect -1816 -213 -1782 -179
rect -1816 -281 -1782 -247
rect -1816 -349 -1782 -315
rect -1816 -417 -1782 -383
rect -1816 -485 -1782 -451
rect -1816 -553 -1782 -519
rect -1816 -621 -1782 -587
rect -1816 -689 -1782 -655
rect -1816 -757 -1782 -723
rect -1816 -825 -1782 -791
rect 1932 -9 1966 25
rect 1932 -77 1966 -43
rect 1932 -145 1966 -111
rect 1932 -213 1966 -179
rect 1932 -281 1966 -247
rect 1932 -349 1966 -315
rect 1932 -417 1966 -383
rect 1932 -485 1966 -451
rect 1932 -553 1966 -519
rect 1932 -621 1966 -587
rect 1932 -689 1966 -655
rect 1932 -757 1966 -723
rect 1932 -825 1966 -791
rect -1608 -958 -1574 -924
rect -1540 -958 -1506 -924
rect -1472 -958 -1438 -924
rect -1404 -958 -1370 -924
rect -1336 -958 -1302 -924
rect -1268 -958 -1234 -924
rect -1200 -958 -1166 -924
rect -1132 -958 -1098 -924
rect -1064 -958 -1030 -924
rect -996 -958 -962 -924
rect -928 -958 -894 -924
rect -860 -958 -826 -924
rect -792 -958 -758 -924
rect -724 -958 -690 -924
rect -656 -958 -622 -924
rect -588 -958 -554 -924
rect -520 -958 -486 -924
rect -452 -958 -418 -924
rect -384 -958 -350 -924
rect -316 -958 -282 -924
rect -248 -958 -214 -924
rect -180 -958 -146 -924
rect -112 -958 -78 -924
rect -44 -958 -10 -924
rect 24 -958 58 -924
rect 92 -958 126 -924
rect 160 -958 194 -924
rect 228 -958 262 -924
rect 296 -958 330 -924
rect 364 -958 398 -924
rect 432 -958 466 -924
rect 500 -958 534 -924
rect 568 -958 602 -924
rect 636 -958 670 -924
rect 704 -958 738 -924
rect 772 -958 806 -924
rect 840 -958 874 -924
rect 908 -958 942 -924
rect 976 -958 1010 -924
rect 1044 -958 1078 -924
rect 1112 -958 1146 -924
rect 1180 -958 1214 -924
rect 1248 -958 1282 -924
rect 1316 -958 1350 -924
rect 1384 -958 1418 -924
rect 1452 -958 1486 -924
rect 1520 -958 1554 -924
rect 1588 -958 1622 -924
rect 1656 -958 1690 -924
rect 1724 -958 1758 -924
<< mvnsubdiffcont >>
rect 24 59 126 5941
<< poly >>
rect -1600 6300 1750 6800
rect -1600 6000 -200 6300
rect 350 6000 1750 6300
rect -400 0 -200 6000
rect 350 0 550 6000
rect -1600 -300 -200 0
rect 350 -300 1750 0
rect -1600 -459 1750 -300
rect -1600 -493 -280 -459
rect -246 -493 -206 -459
rect -172 -493 -132 -459
rect -98 -493 -58 -459
rect -24 -493 16 -459
rect 50 -493 90 -459
rect 124 -493 164 -459
rect 198 -493 238 -459
rect 272 -493 312 -459
rect 346 -493 386 -459
rect 420 -493 1750 -459
rect -1600 -533 1750 -493
rect -1600 -567 -280 -533
rect -246 -567 -206 -533
rect -172 -567 -132 -533
rect -98 -567 -58 -533
rect -24 -567 16 -533
rect 50 -567 90 -533
rect 124 -567 164 -533
rect 198 -567 238 -533
rect 272 -567 312 -533
rect 346 -567 386 -533
rect 420 -567 1750 -533
rect -1600 -607 1750 -567
rect -1600 -641 -280 -607
rect -246 -641 -206 -607
rect -172 -641 -132 -607
rect -98 -641 -58 -607
rect -24 -641 16 -607
rect 50 -641 90 -607
rect 124 -641 164 -607
rect 198 -641 238 -607
rect 272 -641 312 -607
rect 346 -641 386 -607
rect 420 -641 1750 -607
rect -1600 -800 1750 -641
<< polycont >>
rect -280 -493 -246 -459
rect -206 -493 -172 -459
rect -132 -493 -98 -459
rect -58 -493 -24 -459
rect 16 -493 50 -459
rect 90 -493 124 -459
rect 164 -493 198 -459
rect 238 -493 272 -459
rect 312 -493 346 -459
rect 386 -493 420 -459
rect -280 -567 -246 -533
rect -206 -567 -172 -533
rect -132 -567 -98 -533
rect -58 -567 -24 -533
rect 16 -567 50 -533
rect 90 -567 124 -533
rect 164 -567 198 -533
rect 238 -567 272 -533
rect 312 -567 346 -533
rect 386 -567 420 -533
rect -280 -641 -246 -607
rect -206 -641 -172 -607
rect -132 -641 -98 -607
rect -58 -641 -24 -607
rect 16 -641 50 -607
rect 90 -641 124 -607
rect 164 -641 198 -607
rect 238 -641 272 -607
rect 312 -641 346 -607
rect 386 -641 420 -607
<< locali >>
rect -1840 6958 1990 6982
rect -1840 6924 -1608 6958
rect -1574 6924 -1540 6958
rect -1506 6924 -1472 6958
rect -1438 6924 -1404 6958
rect -1370 6924 -1336 6958
rect -1302 6924 -1268 6958
rect -1234 6924 -1200 6958
rect -1166 6924 -1132 6958
rect -1098 6924 -1064 6958
rect -1030 6924 -996 6958
rect -962 6924 -928 6958
rect -894 6924 -860 6958
rect -826 6924 -792 6958
rect -758 6924 -724 6958
rect -690 6924 -656 6958
rect -622 6924 -588 6958
rect -554 6924 -520 6958
rect -486 6924 -452 6958
rect -418 6924 -384 6958
rect -350 6924 -316 6958
rect -282 6924 -248 6958
rect -214 6924 -180 6958
rect -146 6924 -112 6958
rect -78 6924 -44 6958
rect -10 6924 24 6958
rect 58 6924 92 6958
rect 126 6924 160 6958
rect 194 6924 228 6958
rect 262 6924 296 6958
rect 330 6924 364 6958
rect 398 6924 432 6958
rect 466 6924 500 6958
rect 534 6924 568 6958
rect 602 6924 636 6958
rect 670 6924 704 6958
rect 738 6924 772 6958
rect 806 6924 840 6958
rect 874 6924 908 6958
rect 942 6924 976 6958
rect 1010 6924 1044 6958
rect 1078 6924 1112 6958
rect 1146 6924 1180 6958
rect 1214 6924 1248 6958
rect 1282 6924 1316 6958
rect 1350 6924 1384 6958
rect 1418 6924 1452 6958
rect 1486 6924 1520 6958
rect 1554 6924 1588 6958
rect 1622 6924 1656 6958
rect 1690 6924 1724 6958
rect 1758 6924 1990 6958
rect -1840 6900 1990 6924
rect -1840 6825 -1758 6900
rect -1840 6791 -1816 6825
rect -1782 6791 -1758 6825
rect -1840 6757 -1758 6791
rect -1840 6723 -1816 6757
rect -1782 6723 -1758 6757
rect -1840 6689 -1758 6723
rect -1840 6655 -1816 6689
rect -1782 6655 -1758 6689
rect -1840 6621 -1758 6655
rect -1840 6587 -1816 6621
rect -1782 6587 -1758 6621
rect -1840 6553 -1758 6587
rect -1840 6519 -1816 6553
rect -1782 6519 -1758 6553
rect -1840 6485 -1758 6519
rect -1840 6451 -1816 6485
rect -1782 6451 -1758 6485
rect -1840 6417 -1758 6451
rect -1840 6383 -1816 6417
rect -1782 6383 -1758 6417
rect -1840 6349 -1758 6383
rect -1840 6315 -1816 6349
rect -1782 6315 -1758 6349
rect -1840 6281 -1758 6315
rect -1840 6247 -1816 6281
rect -1782 6247 -1758 6281
rect -1840 6213 -1758 6247
rect -1840 6179 -1816 6213
rect -1782 6179 -1758 6213
rect -1840 6145 -1758 6179
rect -1840 6111 -1816 6145
rect -1782 6111 -1758 6145
rect -1840 6077 -1758 6111
rect -1840 6043 -1816 6077
rect -1782 6043 -1758 6077
rect 1908 6825 1990 6900
rect 1908 6791 1932 6825
rect 1966 6791 1990 6825
rect 1908 6757 1990 6791
rect 1908 6723 1932 6757
rect 1966 6723 1990 6757
rect 1908 6689 1990 6723
rect 1908 6655 1932 6689
rect 1966 6655 1990 6689
rect 1908 6621 1990 6655
rect 1908 6587 1932 6621
rect 1966 6587 1990 6621
rect 1908 6553 1990 6587
rect 1908 6519 1932 6553
rect 1966 6519 1990 6553
rect 1908 6485 1990 6519
rect 1908 6451 1932 6485
rect 1966 6451 1990 6485
rect 1908 6417 1990 6451
rect 1908 6383 1932 6417
rect 1966 6383 1990 6417
rect 1908 6349 1990 6383
rect 1908 6315 1932 6349
rect 1966 6315 1990 6349
rect 1908 6281 1990 6315
rect 1908 6247 1932 6281
rect 1966 6247 1990 6281
rect 1908 6213 1990 6247
rect 1908 6179 1932 6213
rect 1966 6179 1990 6213
rect 1908 6145 1990 6179
rect 1908 6111 1932 6145
rect 1966 6111 1990 6145
rect 1908 6077 1990 6111
rect -1840 6009 -1758 6043
rect -1840 5975 -1816 6009
rect -1782 5975 -1758 6009
rect -1840 5941 -1758 5975
rect -1840 5907 -1816 5941
rect -1782 5907 -1758 5941
rect -1840 5873 -1758 5907
rect -1840 5839 -1816 5873
rect -1782 5839 -1758 5873
rect -1840 5805 -1758 5839
rect -1840 5771 -1816 5805
rect -1782 5771 -1758 5805
rect -1840 5737 -1758 5771
rect -1840 5703 -1816 5737
rect -1782 5703 -1758 5737
rect -1840 5669 -1758 5703
rect -1840 5635 -1816 5669
rect -1782 5635 -1758 5669
rect -1840 5601 -1758 5635
rect -1840 5567 -1816 5601
rect -1782 5567 -1758 5601
rect -1840 5533 -1758 5567
rect -1840 5499 -1816 5533
rect -1782 5499 -1758 5533
rect -1840 5465 -1758 5499
rect -1840 5431 -1816 5465
rect -1782 5431 -1758 5465
rect -1840 5397 -1758 5431
rect -1840 5363 -1816 5397
rect -1782 5363 -1758 5397
rect -1840 5329 -1758 5363
rect -1840 5295 -1816 5329
rect -1782 5295 -1758 5329
rect -1840 5261 -1758 5295
rect -1840 5227 -1816 5261
rect -1782 5227 -1758 5261
rect -1840 5193 -1758 5227
rect -1840 5159 -1816 5193
rect -1782 5159 -1758 5193
rect -1840 5125 -1758 5159
rect -1840 5091 -1816 5125
rect -1782 5091 -1758 5125
rect -1840 5057 -1758 5091
rect -1840 5023 -1816 5057
rect -1782 5023 -1758 5057
rect -1840 4989 -1758 5023
rect -1840 4955 -1816 4989
rect -1782 4955 -1758 4989
rect -1840 4921 -1758 4955
rect -1840 4887 -1816 4921
rect -1782 4887 -1758 4921
rect -1840 4853 -1758 4887
rect -1840 4819 -1816 4853
rect -1782 4819 -1758 4853
rect -1840 4785 -1758 4819
rect -1840 4751 -1816 4785
rect -1782 4751 -1758 4785
rect -1840 4717 -1758 4751
rect -1840 4683 -1816 4717
rect -1782 4683 -1758 4717
rect -1840 4649 -1758 4683
rect -1840 4615 -1816 4649
rect -1782 4615 -1758 4649
rect -1840 4581 -1758 4615
rect -1840 4547 -1816 4581
rect -1782 4547 -1758 4581
rect -1840 4513 -1758 4547
rect -1840 4479 -1816 4513
rect -1782 4479 -1758 4513
rect -1840 4445 -1758 4479
rect -1840 4411 -1816 4445
rect -1782 4411 -1758 4445
rect -1840 4377 -1758 4411
rect -1840 4343 -1816 4377
rect -1782 4343 -1758 4377
rect -1840 4309 -1758 4343
rect -1840 4275 -1816 4309
rect -1782 4275 -1758 4309
rect -1840 4241 -1758 4275
rect -1840 4207 -1816 4241
rect -1782 4207 -1758 4241
rect -1840 4173 -1758 4207
rect -1840 4139 -1816 4173
rect -1782 4139 -1758 4173
rect -1840 4105 -1758 4139
rect -1840 4071 -1816 4105
rect -1782 4071 -1758 4105
rect -1840 4037 -1758 4071
rect -1840 4003 -1816 4037
rect -1782 4003 -1758 4037
rect -1840 3969 -1758 4003
rect -1840 3935 -1816 3969
rect -1782 3935 -1758 3969
rect -1840 3901 -1758 3935
rect -1840 3867 -1816 3901
rect -1782 3867 -1758 3901
rect -1840 3833 -1758 3867
rect -1840 3799 -1816 3833
rect -1782 3799 -1758 3833
rect -1840 3765 -1758 3799
rect -1840 3731 -1816 3765
rect -1782 3731 -1758 3765
rect -1840 3697 -1758 3731
rect -1840 3663 -1816 3697
rect -1782 3663 -1758 3697
rect -1840 3629 -1758 3663
rect -1840 3595 -1816 3629
rect -1782 3595 -1758 3629
rect -1840 3561 -1758 3595
rect -1840 3527 -1816 3561
rect -1782 3527 -1758 3561
rect -1840 3493 -1758 3527
rect -1840 3459 -1816 3493
rect -1782 3459 -1758 3493
rect -1840 3425 -1758 3459
rect -1840 3391 -1816 3425
rect -1782 3391 -1758 3425
rect -1840 3357 -1758 3391
rect -1840 3323 -1816 3357
rect -1782 3323 -1758 3357
rect -1840 3289 -1758 3323
rect -1840 3255 -1816 3289
rect -1782 3255 -1758 3289
rect -1840 3221 -1758 3255
rect -1840 3187 -1816 3221
rect -1782 3187 -1758 3221
rect -1840 3153 -1758 3187
rect -1840 3119 -1816 3153
rect -1782 3119 -1758 3153
rect -1840 3085 -1758 3119
rect -1840 3051 -1816 3085
rect -1782 3051 -1758 3085
rect -1840 3017 -1758 3051
rect -1840 2983 -1816 3017
rect -1782 2983 -1758 3017
rect -1840 2949 -1758 2983
rect -1840 2915 -1816 2949
rect -1782 2915 -1758 2949
rect -1840 2881 -1758 2915
rect -1840 2847 -1816 2881
rect -1782 2847 -1758 2881
rect -1840 2813 -1758 2847
rect -1840 2779 -1816 2813
rect -1782 2779 -1758 2813
rect -1840 2745 -1758 2779
rect -1840 2711 -1816 2745
rect -1782 2711 -1758 2745
rect -1840 2677 -1758 2711
rect -1840 2643 -1816 2677
rect -1782 2643 -1758 2677
rect -1840 2609 -1758 2643
rect -1840 2575 -1816 2609
rect -1782 2575 -1758 2609
rect -1840 2541 -1758 2575
rect -1840 2507 -1816 2541
rect -1782 2507 -1758 2541
rect -1840 2473 -1758 2507
rect -1840 2439 -1816 2473
rect -1782 2439 -1758 2473
rect -1840 2405 -1758 2439
rect -1840 2371 -1816 2405
rect -1782 2371 -1758 2405
rect -1840 2337 -1758 2371
rect -1840 2303 -1816 2337
rect -1782 2303 -1758 2337
rect -1840 2269 -1758 2303
rect -1840 2235 -1816 2269
rect -1782 2235 -1758 2269
rect -1840 2201 -1758 2235
rect -1840 2167 -1816 2201
rect -1782 2167 -1758 2201
rect -1840 2133 -1758 2167
rect -1840 2099 -1816 2133
rect -1782 2099 -1758 2133
rect -1840 2065 -1758 2099
rect -1840 2031 -1816 2065
rect -1782 2031 -1758 2065
rect -1840 1997 -1758 2031
rect -1840 1963 -1816 1997
rect -1782 1963 -1758 1997
rect -1840 1929 -1758 1963
rect -1840 1895 -1816 1929
rect -1782 1895 -1758 1929
rect -1840 1861 -1758 1895
rect -1840 1827 -1816 1861
rect -1782 1827 -1758 1861
rect -1840 1793 -1758 1827
rect -1840 1759 -1816 1793
rect -1782 1759 -1758 1793
rect -1840 1725 -1758 1759
rect -1840 1691 -1816 1725
rect -1782 1691 -1758 1725
rect -1840 1657 -1758 1691
rect -1840 1623 -1816 1657
rect -1782 1623 -1758 1657
rect -1840 1589 -1758 1623
rect -1840 1555 -1816 1589
rect -1782 1555 -1758 1589
rect -1840 1521 -1758 1555
rect -1840 1487 -1816 1521
rect -1782 1487 -1758 1521
rect -1840 1453 -1758 1487
rect -1840 1419 -1816 1453
rect -1782 1419 -1758 1453
rect -1840 1385 -1758 1419
rect -1840 1351 -1816 1385
rect -1782 1351 -1758 1385
rect -1840 1317 -1758 1351
rect -1840 1283 -1816 1317
rect -1782 1283 -1758 1317
rect -1840 1249 -1758 1283
rect -1840 1215 -1816 1249
rect -1782 1215 -1758 1249
rect -1840 1181 -1758 1215
rect -1840 1147 -1816 1181
rect -1782 1147 -1758 1181
rect -1840 1113 -1758 1147
rect -1840 1079 -1816 1113
rect -1782 1079 -1758 1113
rect -1840 1045 -1758 1079
rect -1840 1011 -1816 1045
rect -1782 1011 -1758 1045
rect -1840 977 -1758 1011
rect -1840 943 -1816 977
rect -1782 943 -1758 977
rect -1840 909 -1758 943
rect -1840 875 -1816 909
rect -1782 875 -1758 909
rect -1840 841 -1758 875
rect -1840 807 -1816 841
rect -1782 807 -1758 841
rect -1840 773 -1758 807
rect -1840 739 -1816 773
rect -1782 739 -1758 773
rect -1840 705 -1758 739
rect -1840 671 -1816 705
rect -1782 671 -1758 705
rect -1840 637 -1758 671
rect -1840 603 -1816 637
rect -1782 603 -1758 637
rect -1840 569 -1758 603
rect -1840 535 -1816 569
rect -1782 535 -1758 569
rect -1840 501 -1758 535
rect -1840 467 -1816 501
rect -1782 467 -1758 501
rect -1840 433 -1758 467
rect -1840 399 -1816 433
rect -1782 399 -1758 433
rect -1840 365 -1758 399
rect -1840 331 -1816 365
rect -1782 331 -1758 365
rect -1840 297 -1758 331
rect -1840 263 -1816 297
rect -1782 263 -1758 297
rect -1840 229 -1758 263
rect -1840 195 -1816 229
rect -1782 195 -1758 229
rect -1840 161 -1758 195
rect -1840 127 -1816 161
rect -1782 127 -1758 161
rect -1840 93 -1758 127
rect -1840 59 -1816 93
rect -1782 59 -1758 93
rect -1840 25 -1758 59
rect -1840 -9 -1816 25
rect -1782 -9 -1758 25
rect -1662 5975 -1596 5991
rect -1662 5935 -1646 5975
rect -1612 5935 -1596 5975
rect -1662 5907 -1596 5935
rect -1662 5863 -1646 5907
rect -1612 5863 -1596 5907
rect -1662 5839 -1596 5863
rect -1662 5791 -1646 5839
rect -1612 5791 -1596 5839
rect -1662 5771 -1596 5791
rect -1662 5719 -1646 5771
rect -1612 5719 -1596 5771
rect -1662 5703 -1596 5719
rect -1662 5647 -1646 5703
rect -1612 5647 -1596 5703
rect -1662 5635 -1596 5647
rect -1662 5575 -1646 5635
rect -1612 5575 -1596 5635
rect -1662 5567 -1596 5575
rect -1662 5503 -1646 5567
rect -1612 5503 -1596 5567
rect -1662 5499 -1596 5503
rect -1662 5397 -1646 5499
rect -1612 5397 -1596 5499
rect -1662 5393 -1596 5397
rect -1662 5329 -1646 5393
rect -1612 5329 -1596 5393
rect -1662 5321 -1596 5329
rect -1662 5261 -1646 5321
rect -1612 5261 -1596 5321
rect -1662 5249 -1596 5261
rect -1662 5193 -1646 5249
rect -1612 5193 -1596 5249
rect -1662 5177 -1596 5193
rect -1662 5125 -1646 5177
rect -1612 5125 -1596 5177
rect -1662 5105 -1596 5125
rect -1662 5057 -1646 5105
rect -1612 5057 -1596 5105
rect -1662 5033 -1596 5057
rect -1662 4989 -1646 5033
rect -1612 4989 -1596 5033
rect -1662 4961 -1596 4989
rect -1662 4921 -1646 4961
rect -1612 4921 -1596 4961
rect -1662 4889 -1596 4921
rect -1662 4853 -1646 4889
rect -1612 4853 -1596 4889
rect -1662 4819 -1596 4853
rect -1662 4783 -1646 4819
rect -1612 4783 -1596 4819
rect -1662 4751 -1596 4783
rect -1662 4711 -1646 4751
rect -1612 4711 -1596 4751
rect -1662 4683 -1596 4711
rect -1662 4639 -1646 4683
rect -1612 4639 -1596 4683
rect -1662 4615 -1596 4639
rect -1662 4567 -1646 4615
rect -1612 4567 -1596 4615
rect -1662 4547 -1596 4567
rect -1662 4495 -1646 4547
rect -1612 4495 -1596 4547
rect -1662 4479 -1596 4495
rect -1662 4423 -1646 4479
rect -1612 4423 -1596 4479
rect -1662 4411 -1596 4423
rect -1662 4351 -1646 4411
rect -1612 4351 -1596 4411
rect -1662 4343 -1596 4351
rect -1662 4279 -1646 4343
rect -1612 4279 -1596 4343
rect -1662 4275 -1596 4279
rect -1662 4173 -1646 4275
rect -1612 4173 -1596 4275
rect -1662 4169 -1596 4173
rect -1662 4105 -1646 4169
rect -1612 4105 -1596 4169
rect -1662 4097 -1596 4105
rect -1662 4037 -1646 4097
rect -1612 4037 -1596 4097
rect -1662 4025 -1596 4037
rect -1662 3969 -1646 4025
rect -1612 3969 -1596 4025
rect -1662 3953 -1596 3969
rect -1662 3901 -1646 3953
rect -1612 3901 -1596 3953
rect -1662 3881 -1596 3901
rect -1662 3833 -1646 3881
rect -1612 3833 -1596 3881
rect -1662 3809 -1596 3833
rect -1662 3765 -1646 3809
rect -1612 3765 -1596 3809
rect -1662 3737 -1596 3765
rect -1662 3697 -1646 3737
rect -1612 3697 -1596 3737
rect -1662 3665 -1596 3697
rect -1662 3629 -1646 3665
rect -1612 3629 -1596 3665
rect -1662 3595 -1596 3629
rect -1662 3559 -1646 3595
rect -1612 3559 -1596 3595
rect -1662 3527 -1596 3559
rect -1662 3487 -1646 3527
rect -1612 3487 -1596 3527
rect -1662 3459 -1596 3487
rect -1662 3415 -1646 3459
rect -1612 3415 -1596 3459
rect -1662 3391 -1596 3415
rect -1662 3343 -1646 3391
rect -1612 3343 -1596 3391
rect -1662 3323 -1596 3343
rect -1662 3271 -1646 3323
rect -1612 3271 -1596 3323
rect -1662 3255 -1596 3271
rect -1662 3199 -1646 3255
rect -1612 3199 -1596 3255
rect -1662 3187 -1596 3199
rect -1662 3127 -1646 3187
rect -1612 3127 -1596 3187
rect -1662 3119 -1596 3127
rect -1662 3055 -1646 3119
rect -1612 3055 -1596 3119
rect -1662 3051 -1596 3055
rect -1662 2949 -1646 3051
rect -1612 2949 -1596 3051
rect -1662 2945 -1596 2949
rect -1662 2881 -1646 2945
rect -1612 2881 -1596 2945
rect -1662 2873 -1596 2881
rect -1662 2813 -1646 2873
rect -1612 2813 -1596 2873
rect -1662 2801 -1596 2813
rect -1662 2745 -1646 2801
rect -1612 2745 -1596 2801
rect -1662 2729 -1596 2745
rect -1662 2677 -1646 2729
rect -1612 2677 -1596 2729
rect -1662 2657 -1596 2677
rect -1662 2609 -1646 2657
rect -1612 2609 -1596 2657
rect -1662 2585 -1596 2609
rect -1662 2541 -1646 2585
rect -1612 2541 -1596 2585
rect -1662 2513 -1596 2541
rect -1662 2473 -1646 2513
rect -1612 2473 -1596 2513
rect -1662 2441 -1596 2473
rect -1662 2405 -1646 2441
rect -1612 2405 -1596 2441
rect -1662 2371 -1596 2405
rect -1662 2335 -1646 2371
rect -1612 2335 -1596 2371
rect -1662 2303 -1596 2335
rect -1662 2263 -1646 2303
rect -1612 2263 -1596 2303
rect -1662 2235 -1596 2263
rect -1662 2191 -1646 2235
rect -1612 2191 -1596 2235
rect -1662 2167 -1596 2191
rect -1662 2119 -1646 2167
rect -1612 2119 -1596 2167
rect -1662 2099 -1596 2119
rect -1662 2047 -1646 2099
rect -1612 2047 -1596 2099
rect -1662 2031 -1596 2047
rect -1662 1975 -1646 2031
rect -1612 1975 -1596 2031
rect -1662 1963 -1596 1975
rect -1662 1903 -1646 1963
rect -1612 1903 -1596 1963
rect -1662 1895 -1596 1903
rect -1662 1831 -1646 1895
rect -1612 1831 -1596 1895
rect -1662 1827 -1596 1831
rect -1662 1725 -1646 1827
rect -1612 1725 -1596 1827
rect -1662 1721 -1596 1725
rect -1662 1657 -1646 1721
rect -1612 1657 -1596 1721
rect -1662 1649 -1596 1657
rect -1662 1589 -1646 1649
rect -1612 1589 -1596 1649
rect -1662 1577 -1596 1589
rect -1662 1521 -1646 1577
rect -1612 1521 -1596 1577
rect -1662 1505 -1596 1521
rect -1662 1453 -1646 1505
rect -1612 1453 -1596 1505
rect -1662 1433 -1596 1453
rect -1662 1385 -1646 1433
rect -1612 1385 -1596 1433
rect -1662 1361 -1596 1385
rect -1662 1317 -1646 1361
rect -1612 1317 -1596 1361
rect -1662 1289 -1596 1317
rect -1662 1249 -1646 1289
rect -1612 1249 -1596 1289
rect -1662 1217 -1596 1249
rect -1662 1181 -1646 1217
rect -1612 1181 -1596 1217
rect -1662 1147 -1596 1181
rect -1662 1111 -1646 1147
rect -1612 1111 -1596 1147
rect -1662 1079 -1596 1111
rect -1662 1039 -1646 1079
rect -1612 1039 -1596 1079
rect -1662 1011 -1596 1039
rect -1662 967 -1646 1011
rect -1612 967 -1596 1011
rect -1662 943 -1596 967
rect -1662 895 -1646 943
rect -1612 895 -1596 943
rect -1662 875 -1596 895
rect -1662 823 -1646 875
rect -1612 823 -1596 875
rect -1662 807 -1596 823
rect -1662 751 -1646 807
rect -1612 751 -1596 807
rect -1662 739 -1596 751
rect -1662 679 -1646 739
rect -1612 679 -1596 739
rect -1662 671 -1596 679
rect -1662 607 -1646 671
rect -1612 607 -1596 671
rect -1662 603 -1596 607
rect -1662 501 -1646 603
rect -1612 501 -1596 603
rect -1662 497 -1596 501
rect -1662 433 -1646 497
rect -1612 433 -1596 497
rect -1662 425 -1596 433
rect -1662 365 -1646 425
rect -1612 365 -1596 425
rect -1662 353 -1596 365
rect -1662 297 -1646 353
rect -1612 297 -1596 353
rect -1662 281 -1596 297
rect -1662 229 -1646 281
rect -1612 229 -1596 281
rect -1662 209 -1596 229
rect -1662 161 -1646 209
rect -1612 161 -1596 209
rect -1662 137 -1596 161
rect -1662 93 -1646 137
rect -1612 93 -1596 137
rect -1662 65 -1596 93
rect -1662 25 -1646 65
rect -1612 25 -1596 65
rect -1662 9 -1596 25
rect -25 5969 175 6050
rect 1908 6043 1932 6077
rect 1966 6043 1990 6077
rect 1908 6009 1990 6043
rect -25 31 22 5969
rect 128 31 175 5969
rect -1840 -43 -1758 -9
rect -1840 -77 -1816 -43
rect -1782 -77 -1758 -43
rect -25 -50 175 31
rect 1746 5975 1812 5991
rect 1746 5935 1762 5975
rect 1796 5935 1812 5975
rect 1746 5907 1812 5935
rect 1746 5863 1762 5907
rect 1796 5863 1812 5907
rect 1746 5839 1812 5863
rect 1746 5791 1762 5839
rect 1796 5791 1812 5839
rect 1746 5771 1812 5791
rect 1746 5719 1762 5771
rect 1796 5719 1812 5771
rect 1746 5703 1812 5719
rect 1746 5647 1762 5703
rect 1796 5647 1812 5703
rect 1746 5635 1812 5647
rect 1746 5575 1762 5635
rect 1796 5575 1812 5635
rect 1746 5567 1812 5575
rect 1746 5503 1762 5567
rect 1796 5503 1812 5567
rect 1746 5499 1812 5503
rect 1746 5397 1762 5499
rect 1796 5397 1812 5499
rect 1746 5393 1812 5397
rect 1746 5329 1762 5393
rect 1796 5329 1812 5393
rect 1746 5321 1812 5329
rect 1746 5261 1762 5321
rect 1796 5261 1812 5321
rect 1746 5249 1812 5261
rect 1746 5193 1762 5249
rect 1796 5193 1812 5249
rect 1746 5177 1812 5193
rect 1746 5125 1762 5177
rect 1796 5125 1812 5177
rect 1746 5105 1812 5125
rect 1746 5057 1762 5105
rect 1796 5057 1812 5105
rect 1746 5033 1812 5057
rect 1746 4989 1762 5033
rect 1796 4989 1812 5033
rect 1746 4961 1812 4989
rect 1746 4921 1762 4961
rect 1796 4921 1812 4961
rect 1746 4889 1812 4921
rect 1746 4853 1762 4889
rect 1796 4853 1812 4889
rect 1746 4819 1812 4853
rect 1746 4783 1762 4819
rect 1796 4783 1812 4819
rect 1746 4751 1812 4783
rect 1746 4711 1762 4751
rect 1796 4711 1812 4751
rect 1746 4683 1812 4711
rect 1746 4639 1762 4683
rect 1796 4639 1812 4683
rect 1746 4615 1812 4639
rect 1746 4567 1762 4615
rect 1796 4567 1812 4615
rect 1746 4547 1812 4567
rect 1746 4495 1762 4547
rect 1796 4495 1812 4547
rect 1746 4479 1812 4495
rect 1746 4423 1762 4479
rect 1796 4423 1812 4479
rect 1746 4411 1812 4423
rect 1746 4351 1762 4411
rect 1796 4351 1812 4411
rect 1746 4343 1812 4351
rect 1746 4279 1762 4343
rect 1796 4279 1812 4343
rect 1746 4275 1812 4279
rect 1746 4173 1762 4275
rect 1796 4173 1812 4275
rect 1746 4169 1812 4173
rect 1746 4105 1762 4169
rect 1796 4105 1812 4169
rect 1746 4097 1812 4105
rect 1746 4037 1762 4097
rect 1796 4037 1812 4097
rect 1746 4025 1812 4037
rect 1746 3969 1762 4025
rect 1796 3969 1812 4025
rect 1746 3953 1812 3969
rect 1746 3901 1762 3953
rect 1796 3901 1812 3953
rect 1746 3881 1812 3901
rect 1746 3833 1762 3881
rect 1796 3833 1812 3881
rect 1746 3809 1812 3833
rect 1746 3765 1762 3809
rect 1796 3765 1812 3809
rect 1746 3737 1812 3765
rect 1746 3697 1762 3737
rect 1796 3697 1812 3737
rect 1746 3665 1812 3697
rect 1746 3629 1762 3665
rect 1796 3629 1812 3665
rect 1746 3595 1812 3629
rect 1746 3559 1762 3595
rect 1796 3559 1812 3595
rect 1746 3527 1812 3559
rect 1746 3487 1762 3527
rect 1796 3487 1812 3527
rect 1746 3459 1812 3487
rect 1746 3415 1762 3459
rect 1796 3415 1812 3459
rect 1746 3391 1812 3415
rect 1746 3343 1762 3391
rect 1796 3343 1812 3391
rect 1746 3323 1812 3343
rect 1746 3271 1762 3323
rect 1796 3271 1812 3323
rect 1746 3255 1812 3271
rect 1746 3199 1762 3255
rect 1796 3199 1812 3255
rect 1746 3187 1812 3199
rect 1746 3127 1762 3187
rect 1796 3127 1812 3187
rect 1746 3119 1812 3127
rect 1746 3055 1762 3119
rect 1796 3055 1812 3119
rect 1746 3051 1812 3055
rect 1746 2949 1762 3051
rect 1796 2949 1812 3051
rect 1746 2945 1812 2949
rect 1746 2881 1762 2945
rect 1796 2881 1812 2945
rect 1746 2873 1812 2881
rect 1746 2813 1762 2873
rect 1796 2813 1812 2873
rect 1746 2801 1812 2813
rect 1746 2745 1762 2801
rect 1796 2745 1812 2801
rect 1746 2729 1812 2745
rect 1746 2677 1762 2729
rect 1796 2677 1812 2729
rect 1746 2657 1812 2677
rect 1746 2609 1762 2657
rect 1796 2609 1812 2657
rect 1746 2585 1812 2609
rect 1746 2541 1762 2585
rect 1796 2541 1812 2585
rect 1746 2513 1812 2541
rect 1746 2473 1762 2513
rect 1796 2473 1812 2513
rect 1746 2441 1812 2473
rect 1746 2405 1762 2441
rect 1796 2405 1812 2441
rect 1746 2371 1812 2405
rect 1746 2335 1762 2371
rect 1796 2335 1812 2371
rect 1746 2303 1812 2335
rect 1746 2263 1762 2303
rect 1796 2263 1812 2303
rect 1746 2235 1812 2263
rect 1746 2191 1762 2235
rect 1796 2191 1812 2235
rect 1746 2167 1812 2191
rect 1746 2119 1762 2167
rect 1796 2119 1812 2167
rect 1746 2099 1812 2119
rect 1746 2047 1762 2099
rect 1796 2047 1812 2099
rect 1746 2031 1812 2047
rect 1746 1975 1762 2031
rect 1796 1975 1812 2031
rect 1746 1963 1812 1975
rect 1746 1903 1762 1963
rect 1796 1903 1812 1963
rect 1746 1895 1812 1903
rect 1746 1831 1762 1895
rect 1796 1831 1812 1895
rect 1746 1827 1812 1831
rect 1746 1725 1762 1827
rect 1796 1725 1812 1827
rect 1746 1721 1812 1725
rect 1746 1657 1762 1721
rect 1796 1657 1812 1721
rect 1746 1649 1812 1657
rect 1746 1589 1762 1649
rect 1796 1589 1812 1649
rect 1746 1577 1812 1589
rect 1746 1521 1762 1577
rect 1796 1521 1812 1577
rect 1746 1505 1812 1521
rect 1746 1453 1762 1505
rect 1796 1453 1812 1505
rect 1746 1433 1812 1453
rect 1746 1385 1762 1433
rect 1796 1385 1812 1433
rect 1746 1361 1812 1385
rect 1746 1317 1762 1361
rect 1796 1317 1812 1361
rect 1746 1289 1812 1317
rect 1746 1249 1762 1289
rect 1796 1249 1812 1289
rect 1746 1217 1812 1249
rect 1746 1181 1762 1217
rect 1796 1181 1812 1217
rect 1746 1147 1812 1181
rect 1746 1111 1762 1147
rect 1796 1111 1812 1147
rect 1746 1079 1812 1111
rect 1746 1039 1762 1079
rect 1796 1039 1812 1079
rect 1746 1011 1812 1039
rect 1746 967 1762 1011
rect 1796 967 1812 1011
rect 1746 943 1812 967
rect 1746 895 1762 943
rect 1796 895 1812 943
rect 1746 875 1812 895
rect 1746 823 1762 875
rect 1796 823 1812 875
rect 1746 807 1812 823
rect 1746 751 1762 807
rect 1796 751 1812 807
rect 1746 739 1812 751
rect 1746 679 1762 739
rect 1796 679 1812 739
rect 1746 671 1812 679
rect 1746 607 1762 671
rect 1796 607 1812 671
rect 1746 603 1812 607
rect 1746 501 1762 603
rect 1796 501 1812 603
rect 1746 497 1812 501
rect 1746 433 1762 497
rect 1796 433 1812 497
rect 1746 425 1812 433
rect 1746 365 1762 425
rect 1796 365 1812 425
rect 1746 353 1812 365
rect 1746 297 1762 353
rect 1796 297 1812 353
rect 1746 281 1812 297
rect 1746 229 1762 281
rect 1796 229 1812 281
rect 1746 209 1812 229
rect 1746 161 1762 209
rect 1796 161 1812 209
rect 1746 137 1812 161
rect 1746 93 1762 137
rect 1796 93 1812 137
rect 1746 65 1812 93
rect 1746 25 1762 65
rect 1796 25 1812 65
rect 1746 9 1812 25
rect 1908 5975 1932 6009
rect 1966 5975 1990 6009
rect 1908 5941 1990 5975
rect 1908 5907 1932 5941
rect 1966 5907 1990 5941
rect 1908 5873 1990 5907
rect 1908 5839 1932 5873
rect 1966 5839 1990 5873
rect 1908 5805 1990 5839
rect 1908 5771 1932 5805
rect 1966 5771 1990 5805
rect 1908 5737 1990 5771
rect 1908 5703 1932 5737
rect 1966 5703 1990 5737
rect 1908 5669 1990 5703
rect 1908 5635 1932 5669
rect 1966 5635 1990 5669
rect 1908 5601 1990 5635
rect 1908 5567 1932 5601
rect 1966 5567 1990 5601
rect 1908 5533 1990 5567
rect 1908 5499 1932 5533
rect 1966 5499 1990 5533
rect 1908 5465 1990 5499
rect 1908 5431 1932 5465
rect 1966 5431 1990 5465
rect 1908 5397 1990 5431
rect 1908 5363 1932 5397
rect 1966 5363 1990 5397
rect 1908 5329 1990 5363
rect 1908 5295 1932 5329
rect 1966 5295 1990 5329
rect 1908 5261 1990 5295
rect 1908 5227 1932 5261
rect 1966 5227 1990 5261
rect 1908 5193 1990 5227
rect 1908 5159 1932 5193
rect 1966 5159 1990 5193
rect 1908 5125 1990 5159
rect 1908 5091 1932 5125
rect 1966 5091 1990 5125
rect 1908 5057 1990 5091
rect 1908 5023 1932 5057
rect 1966 5023 1990 5057
rect 1908 4989 1990 5023
rect 1908 4955 1932 4989
rect 1966 4955 1990 4989
rect 1908 4921 1990 4955
rect 1908 4887 1932 4921
rect 1966 4887 1990 4921
rect 1908 4853 1990 4887
rect 1908 4819 1932 4853
rect 1966 4819 1990 4853
rect 1908 4785 1990 4819
rect 1908 4751 1932 4785
rect 1966 4751 1990 4785
rect 1908 4717 1990 4751
rect 1908 4683 1932 4717
rect 1966 4683 1990 4717
rect 1908 4649 1990 4683
rect 1908 4615 1932 4649
rect 1966 4615 1990 4649
rect 1908 4581 1990 4615
rect 1908 4547 1932 4581
rect 1966 4547 1990 4581
rect 1908 4513 1990 4547
rect 1908 4479 1932 4513
rect 1966 4479 1990 4513
rect 1908 4445 1990 4479
rect 1908 4411 1932 4445
rect 1966 4411 1990 4445
rect 1908 4377 1990 4411
rect 1908 4343 1932 4377
rect 1966 4343 1990 4377
rect 1908 4309 1990 4343
rect 1908 4275 1932 4309
rect 1966 4275 1990 4309
rect 1908 4241 1990 4275
rect 1908 4207 1932 4241
rect 1966 4207 1990 4241
rect 1908 4173 1990 4207
rect 1908 4139 1932 4173
rect 1966 4139 1990 4173
rect 1908 4105 1990 4139
rect 1908 4071 1932 4105
rect 1966 4071 1990 4105
rect 1908 4037 1990 4071
rect 1908 4003 1932 4037
rect 1966 4003 1990 4037
rect 1908 3969 1990 4003
rect 1908 3935 1932 3969
rect 1966 3935 1990 3969
rect 1908 3901 1990 3935
rect 1908 3867 1932 3901
rect 1966 3867 1990 3901
rect 1908 3833 1990 3867
rect 1908 3799 1932 3833
rect 1966 3799 1990 3833
rect 1908 3765 1990 3799
rect 1908 3731 1932 3765
rect 1966 3731 1990 3765
rect 1908 3697 1990 3731
rect 1908 3663 1932 3697
rect 1966 3663 1990 3697
rect 1908 3629 1990 3663
rect 1908 3595 1932 3629
rect 1966 3595 1990 3629
rect 1908 3561 1990 3595
rect 1908 3527 1932 3561
rect 1966 3527 1990 3561
rect 1908 3493 1990 3527
rect 1908 3459 1932 3493
rect 1966 3459 1990 3493
rect 1908 3425 1990 3459
rect 1908 3391 1932 3425
rect 1966 3391 1990 3425
rect 1908 3357 1990 3391
rect 1908 3323 1932 3357
rect 1966 3323 1990 3357
rect 1908 3289 1990 3323
rect 1908 3255 1932 3289
rect 1966 3255 1990 3289
rect 1908 3221 1990 3255
rect 1908 3187 1932 3221
rect 1966 3187 1990 3221
rect 1908 3153 1990 3187
rect 1908 3119 1932 3153
rect 1966 3119 1990 3153
rect 1908 3085 1990 3119
rect 1908 3051 1932 3085
rect 1966 3051 1990 3085
rect 1908 3017 1990 3051
rect 1908 2983 1932 3017
rect 1966 2983 1990 3017
rect 1908 2949 1990 2983
rect 1908 2915 1932 2949
rect 1966 2915 1990 2949
rect 1908 2881 1990 2915
rect 1908 2847 1932 2881
rect 1966 2847 1990 2881
rect 1908 2813 1990 2847
rect 1908 2779 1932 2813
rect 1966 2779 1990 2813
rect 1908 2745 1990 2779
rect 1908 2711 1932 2745
rect 1966 2711 1990 2745
rect 1908 2677 1990 2711
rect 1908 2643 1932 2677
rect 1966 2643 1990 2677
rect 1908 2609 1990 2643
rect 1908 2575 1932 2609
rect 1966 2575 1990 2609
rect 1908 2541 1990 2575
rect 1908 2507 1932 2541
rect 1966 2507 1990 2541
rect 1908 2473 1990 2507
rect 1908 2439 1932 2473
rect 1966 2439 1990 2473
rect 1908 2405 1990 2439
rect 1908 2371 1932 2405
rect 1966 2371 1990 2405
rect 1908 2337 1990 2371
rect 1908 2303 1932 2337
rect 1966 2303 1990 2337
rect 1908 2269 1990 2303
rect 1908 2235 1932 2269
rect 1966 2235 1990 2269
rect 1908 2201 1990 2235
rect 1908 2167 1932 2201
rect 1966 2167 1990 2201
rect 1908 2133 1990 2167
rect 1908 2099 1932 2133
rect 1966 2099 1990 2133
rect 1908 2065 1990 2099
rect 1908 2031 1932 2065
rect 1966 2031 1990 2065
rect 1908 1997 1990 2031
rect 1908 1963 1932 1997
rect 1966 1963 1990 1997
rect 1908 1929 1990 1963
rect 1908 1895 1932 1929
rect 1966 1895 1990 1929
rect 1908 1861 1990 1895
rect 1908 1827 1932 1861
rect 1966 1827 1990 1861
rect 1908 1793 1990 1827
rect 1908 1759 1932 1793
rect 1966 1759 1990 1793
rect 1908 1725 1990 1759
rect 1908 1691 1932 1725
rect 1966 1691 1990 1725
rect 1908 1657 1990 1691
rect 1908 1623 1932 1657
rect 1966 1623 1990 1657
rect 1908 1589 1990 1623
rect 1908 1555 1932 1589
rect 1966 1555 1990 1589
rect 1908 1521 1990 1555
rect 1908 1487 1932 1521
rect 1966 1487 1990 1521
rect 1908 1453 1990 1487
rect 1908 1419 1932 1453
rect 1966 1419 1990 1453
rect 1908 1385 1990 1419
rect 1908 1351 1932 1385
rect 1966 1351 1990 1385
rect 1908 1317 1990 1351
rect 1908 1283 1932 1317
rect 1966 1283 1990 1317
rect 1908 1249 1990 1283
rect 1908 1215 1932 1249
rect 1966 1215 1990 1249
rect 1908 1181 1990 1215
rect 1908 1147 1932 1181
rect 1966 1147 1990 1181
rect 1908 1113 1990 1147
rect 1908 1079 1932 1113
rect 1966 1079 1990 1113
rect 1908 1045 1990 1079
rect 1908 1011 1932 1045
rect 1966 1011 1990 1045
rect 1908 977 1990 1011
rect 1908 943 1932 977
rect 1966 943 1990 977
rect 1908 909 1990 943
rect 1908 875 1932 909
rect 1966 875 1990 909
rect 1908 841 1990 875
rect 1908 807 1932 841
rect 1966 807 1990 841
rect 1908 773 1990 807
rect 1908 739 1932 773
rect 1966 739 1990 773
rect 1908 705 1990 739
rect 1908 671 1932 705
rect 1966 671 1990 705
rect 1908 637 1990 671
rect 1908 603 1932 637
rect 1966 603 1990 637
rect 1908 569 1990 603
rect 1908 535 1932 569
rect 1966 535 1990 569
rect 1908 501 1990 535
rect 1908 467 1932 501
rect 1966 467 1990 501
rect 1908 433 1990 467
rect 1908 399 1932 433
rect 1966 399 1990 433
rect 1908 365 1990 399
rect 1908 331 1932 365
rect 1966 331 1990 365
rect 1908 297 1990 331
rect 1908 263 1932 297
rect 1966 263 1990 297
rect 1908 229 1990 263
rect 1908 195 1932 229
rect 1966 195 1990 229
rect 1908 161 1990 195
rect 1908 127 1932 161
rect 1966 127 1990 161
rect 1908 93 1990 127
rect 1908 59 1932 93
rect 1966 59 1990 93
rect 1908 25 1990 59
rect 1908 -9 1932 25
rect 1966 -9 1990 25
rect 1908 -43 1990 -9
rect -1840 -111 -1758 -77
rect -1840 -145 -1816 -111
rect -1782 -145 -1758 -111
rect -1840 -179 -1758 -145
rect -1840 -213 -1816 -179
rect -1782 -213 -1758 -179
rect -1840 -247 -1758 -213
rect -1840 -281 -1816 -247
rect -1782 -281 -1758 -247
rect -1840 -315 -1758 -281
rect -1840 -349 -1816 -315
rect -1782 -349 -1758 -315
rect -1840 -383 -1758 -349
rect -1840 -417 -1816 -383
rect -1782 -417 -1758 -383
rect -1840 -451 -1758 -417
rect 1908 -77 1932 -43
rect 1966 -77 1990 -43
rect 1908 -111 1990 -77
rect 1908 -145 1932 -111
rect 1966 -145 1990 -111
rect 1908 -179 1990 -145
rect 1908 -213 1932 -179
rect 1966 -213 1990 -179
rect 1908 -247 1990 -213
rect 1908 -281 1932 -247
rect 1966 -281 1990 -247
rect 1908 -315 1990 -281
rect 1908 -349 1932 -315
rect 1966 -349 1990 -315
rect 1908 -383 1990 -349
rect 1908 -417 1932 -383
rect 1966 -417 1990 -383
rect -1840 -485 -1816 -451
rect -1782 -485 -1758 -451
rect -1840 -519 -1758 -485
rect -1840 -553 -1816 -519
rect -1782 -553 -1758 -519
rect -1840 -587 -1758 -553
rect -1840 -621 -1816 -587
rect -1782 -621 -1758 -587
rect -1840 -655 -1758 -621
rect -1840 -689 -1816 -655
rect -1782 -689 -1758 -655
rect -296 -459 460 -443
rect -296 -493 -280 -459
rect -246 -493 -206 -459
rect -172 -493 -132 -459
rect -98 -493 -58 -459
rect -24 -493 16 -459
rect 50 -493 90 -459
rect 124 -493 164 -459
rect 198 -493 238 -459
rect 272 -493 312 -459
rect 346 -493 386 -459
rect 420 -493 460 -459
rect -296 -533 460 -493
rect -296 -567 -280 -533
rect -246 -567 -206 -533
rect -172 -567 -132 -533
rect -98 -567 -58 -533
rect -24 -567 16 -533
rect 50 -567 90 -533
rect 124 -567 164 -533
rect 198 -567 238 -533
rect 272 -567 312 -533
rect 346 -567 386 -533
rect 420 -567 460 -533
rect -296 -607 460 -567
rect -296 -641 -280 -607
rect -246 -641 -206 -607
rect -172 -641 -132 -607
rect -98 -641 -58 -607
rect -24 -641 16 -607
rect 50 -641 90 -607
rect 124 -641 164 -607
rect 198 -641 238 -607
rect 272 -641 312 -607
rect 346 -641 386 -607
rect 420 -641 460 -607
rect -296 -657 460 -641
rect 1908 -451 1990 -417
rect 1908 -485 1932 -451
rect 1966 -485 1990 -451
rect 1908 -519 1990 -485
rect 1908 -553 1932 -519
rect 1966 -553 1990 -519
rect 1908 -587 1990 -553
rect 1908 -621 1932 -587
rect 1966 -621 1990 -587
rect 1908 -655 1990 -621
rect -1840 -723 -1758 -689
rect -1840 -757 -1816 -723
rect -1782 -757 -1758 -723
rect -1840 -791 -1758 -757
rect -1840 -825 -1816 -791
rect -1782 -825 -1758 -791
rect -1840 -900 -1758 -825
rect 1908 -689 1932 -655
rect 1966 -689 1990 -655
rect 1908 -723 1990 -689
rect 1908 -757 1932 -723
rect 1966 -757 1990 -723
rect 1908 -791 1990 -757
rect 1908 -825 1932 -791
rect 1966 -825 1990 -791
rect 1908 -900 1990 -825
rect -1840 -924 1990 -900
rect -1840 -958 -1608 -924
rect -1574 -958 -1540 -924
rect -1506 -958 -1472 -924
rect -1438 -958 -1404 -924
rect -1370 -958 -1336 -924
rect -1302 -958 -1268 -924
rect -1234 -958 -1200 -924
rect -1166 -958 -1132 -924
rect -1098 -958 -1064 -924
rect -1030 -958 -996 -924
rect -962 -958 -928 -924
rect -894 -958 -860 -924
rect -826 -958 -792 -924
rect -758 -958 -724 -924
rect -690 -958 -656 -924
rect -622 -958 -588 -924
rect -554 -958 -520 -924
rect -486 -958 -452 -924
rect -418 -958 -384 -924
rect -350 -958 -316 -924
rect -282 -958 -248 -924
rect -214 -958 -180 -924
rect -146 -958 -112 -924
rect -78 -958 -44 -924
rect -10 -958 24 -924
rect 58 -958 92 -924
rect 126 -958 160 -924
rect 194 -958 228 -924
rect 262 -958 296 -924
rect 330 -958 364 -924
rect 398 -958 432 -924
rect 466 -958 500 -924
rect 534 -958 568 -924
rect 602 -958 636 -924
rect 670 -958 704 -924
rect 738 -958 772 -924
rect 806 -958 840 -924
rect 874 -958 908 -924
rect 942 -958 976 -924
rect 1010 -958 1044 -924
rect 1078 -958 1112 -924
rect 1146 -958 1180 -924
rect 1214 -958 1248 -924
rect 1282 -958 1316 -924
rect 1350 -958 1384 -924
rect 1418 -958 1452 -924
rect 1486 -958 1520 -924
rect 1554 -958 1588 -924
rect 1622 -958 1656 -924
rect 1690 -958 1724 -924
rect 1758 -958 1990 -924
rect -1840 -982 1990 -958
<< viali >>
rect -1646 5941 -1612 5969
rect -1646 5935 -1612 5941
rect -1646 5873 -1612 5897
rect -1646 5863 -1612 5873
rect -1646 5805 -1612 5825
rect -1646 5791 -1612 5805
rect -1646 5737 -1612 5753
rect -1646 5719 -1612 5737
rect -1646 5669 -1612 5681
rect -1646 5647 -1612 5669
rect -1646 5601 -1612 5609
rect -1646 5575 -1612 5601
rect -1646 5533 -1612 5537
rect -1646 5503 -1612 5533
rect -1646 5431 -1612 5465
rect -1646 5363 -1612 5393
rect -1646 5359 -1612 5363
rect -1646 5295 -1612 5321
rect -1646 5287 -1612 5295
rect -1646 5227 -1612 5249
rect -1646 5215 -1612 5227
rect -1646 5159 -1612 5177
rect -1646 5143 -1612 5159
rect -1646 5091 -1612 5105
rect -1646 5071 -1612 5091
rect -1646 5023 -1612 5033
rect -1646 4999 -1612 5023
rect -1646 4955 -1612 4961
rect -1646 4927 -1612 4955
rect -1646 4887 -1612 4889
rect -1646 4855 -1612 4887
rect -1646 4785 -1612 4817
rect -1646 4783 -1612 4785
rect -1646 4717 -1612 4745
rect -1646 4711 -1612 4717
rect -1646 4649 -1612 4673
rect -1646 4639 -1612 4649
rect -1646 4581 -1612 4601
rect -1646 4567 -1612 4581
rect -1646 4513 -1612 4529
rect -1646 4495 -1612 4513
rect -1646 4445 -1612 4457
rect -1646 4423 -1612 4445
rect -1646 4377 -1612 4385
rect -1646 4351 -1612 4377
rect -1646 4309 -1612 4313
rect -1646 4279 -1612 4309
rect -1646 4207 -1612 4241
rect -1646 4139 -1612 4169
rect -1646 4135 -1612 4139
rect -1646 4071 -1612 4097
rect -1646 4063 -1612 4071
rect -1646 4003 -1612 4025
rect -1646 3991 -1612 4003
rect -1646 3935 -1612 3953
rect -1646 3919 -1612 3935
rect -1646 3867 -1612 3881
rect -1646 3847 -1612 3867
rect -1646 3799 -1612 3809
rect -1646 3775 -1612 3799
rect -1646 3731 -1612 3737
rect -1646 3703 -1612 3731
rect -1646 3663 -1612 3665
rect -1646 3631 -1612 3663
rect -1646 3561 -1612 3593
rect -1646 3559 -1612 3561
rect -1646 3493 -1612 3521
rect -1646 3487 -1612 3493
rect -1646 3425 -1612 3449
rect -1646 3415 -1612 3425
rect -1646 3357 -1612 3377
rect -1646 3343 -1612 3357
rect -1646 3289 -1612 3305
rect -1646 3271 -1612 3289
rect -1646 3221 -1612 3233
rect -1646 3199 -1612 3221
rect -1646 3153 -1612 3161
rect -1646 3127 -1612 3153
rect -1646 3085 -1612 3089
rect -1646 3055 -1612 3085
rect -1646 2983 -1612 3017
rect -1646 2915 -1612 2945
rect -1646 2911 -1612 2915
rect -1646 2847 -1612 2873
rect -1646 2839 -1612 2847
rect -1646 2779 -1612 2801
rect -1646 2767 -1612 2779
rect -1646 2711 -1612 2729
rect -1646 2695 -1612 2711
rect -1646 2643 -1612 2657
rect -1646 2623 -1612 2643
rect -1646 2575 -1612 2585
rect -1646 2551 -1612 2575
rect -1646 2507 -1612 2513
rect -1646 2479 -1612 2507
rect -1646 2439 -1612 2441
rect -1646 2407 -1612 2439
rect -1646 2337 -1612 2369
rect -1646 2335 -1612 2337
rect -1646 2269 -1612 2297
rect -1646 2263 -1612 2269
rect -1646 2201 -1612 2225
rect -1646 2191 -1612 2201
rect -1646 2133 -1612 2153
rect -1646 2119 -1612 2133
rect -1646 2065 -1612 2081
rect -1646 2047 -1612 2065
rect -1646 1997 -1612 2009
rect -1646 1975 -1612 1997
rect -1646 1929 -1612 1937
rect -1646 1903 -1612 1929
rect -1646 1861 -1612 1865
rect -1646 1831 -1612 1861
rect -1646 1759 -1612 1793
rect -1646 1691 -1612 1721
rect -1646 1687 -1612 1691
rect -1646 1623 -1612 1649
rect -1646 1615 -1612 1623
rect -1646 1555 -1612 1577
rect -1646 1543 -1612 1555
rect -1646 1487 -1612 1505
rect -1646 1471 -1612 1487
rect -1646 1419 -1612 1433
rect -1646 1399 -1612 1419
rect -1646 1351 -1612 1361
rect -1646 1327 -1612 1351
rect -1646 1283 -1612 1289
rect -1646 1255 -1612 1283
rect -1646 1215 -1612 1217
rect -1646 1183 -1612 1215
rect -1646 1113 -1612 1145
rect -1646 1111 -1612 1113
rect -1646 1045 -1612 1073
rect -1646 1039 -1612 1045
rect -1646 977 -1612 1001
rect -1646 967 -1612 977
rect -1646 909 -1612 929
rect -1646 895 -1612 909
rect -1646 841 -1612 857
rect -1646 823 -1612 841
rect -1646 773 -1612 785
rect -1646 751 -1612 773
rect -1646 705 -1612 713
rect -1646 679 -1612 705
rect -1646 637 -1612 641
rect -1646 607 -1612 637
rect -1646 535 -1612 569
rect -1646 467 -1612 497
rect -1646 463 -1612 467
rect -1646 399 -1612 425
rect -1646 391 -1612 399
rect -1646 331 -1612 353
rect -1646 319 -1612 331
rect -1646 263 -1612 281
rect -1646 247 -1612 263
rect -1646 195 -1612 209
rect -1646 175 -1612 195
rect -1646 127 -1612 137
rect -1646 103 -1612 127
rect -1646 59 -1612 65
rect -1646 31 -1612 59
rect 22 5941 128 5969
rect 22 59 24 5941
rect 24 59 126 5941
rect 126 59 128 5941
rect 22 31 128 59
rect 1762 5941 1796 5969
rect 1762 5935 1796 5941
rect 1762 5873 1796 5897
rect 1762 5863 1796 5873
rect 1762 5805 1796 5825
rect 1762 5791 1796 5805
rect 1762 5737 1796 5753
rect 1762 5719 1796 5737
rect 1762 5669 1796 5681
rect 1762 5647 1796 5669
rect 1762 5601 1796 5609
rect 1762 5575 1796 5601
rect 1762 5533 1796 5537
rect 1762 5503 1796 5533
rect 1762 5431 1796 5465
rect 1762 5363 1796 5393
rect 1762 5359 1796 5363
rect 1762 5295 1796 5321
rect 1762 5287 1796 5295
rect 1762 5227 1796 5249
rect 1762 5215 1796 5227
rect 1762 5159 1796 5177
rect 1762 5143 1796 5159
rect 1762 5091 1796 5105
rect 1762 5071 1796 5091
rect 1762 5023 1796 5033
rect 1762 4999 1796 5023
rect 1762 4955 1796 4961
rect 1762 4927 1796 4955
rect 1762 4887 1796 4889
rect 1762 4855 1796 4887
rect 1762 4785 1796 4817
rect 1762 4783 1796 4785
rect 1762 4717 1796 4745
rect 1762 4711 1796 4717
rect 1762 4649 1796 4673
rect 1762 4639 1796 4649
rect 1762 4581 1796 4601
rect 1762 4567 1796 4581
rect 1762 4513 1796 4529
rect 1762 4495 1796 4513
rect 1762 4445 1796 4457
rect 1762 4423 1796 4445
rect 1762 4377 1796 4385
rect 1762 4351 1796 4377
rect 1762 4309 1796 4313
rect 1762 4279 1796 4309
rect 1762 4207 1796 4241
rect 1762 4139 1796 4169
rect 1762 4135 1796 4139
rect 1762 4071 1796 4097
rect 1762 4063 1796 4071
rect 1762 4003 1796 4025
rect 1762 3991 1796 4003
rect 1762 3935 1796 3953
rect 1762 3919 1796 3935
rect 1762 3867 1796 3881
rect 1762 3847 1796 3867
rect 1762 3799 1796 3809
rect 1762 3775 1796 3799
rect 1762 3731 1796 3737
rect 1762 3703 1796 3731
rect 1762 3663 1796 3665
rect 1762 3631 1796 3663
rect 1762 3561 1796 3593
rect 1762 3559 1796 3561
rect 1762 3493 1796 3521
rect 1762 3487 1796 3493
rect 1762 3425 1796 3449
rect 1762 3415 1796 3425
rect 1762 3357 1796 3377
rect 1762 3343 1796 3357
rect 1762 3289 1796 3305
rect 1762 3271 1796 3289
rect 1762 3221 1796 3233
rect 1762 3199 1796 3221
rect 1762 3153 1796 3161
rect 1762 3127 1796 3153
rect 1762 3085 1796 3089
rect 1762 3055 1796 3085
rect 1762 2983 1796 3017
rect 1762 2915 1796 2945
rect 1762 2911 1796 2915
rect 1762 2847 1796 2873
rect 1762 2839 1796 2847
rect 1762 2779 1796 2801
rect 1762 2767 1796 2779
rect 1762 2711 1796 2729
rect 1762 2695 1796 2711
rect 1762 2643 1796 2657
rect 1762 2623 1796 2643
rect 1762 2575 1796 2585
rect 1762 2551 1796 2575
rect 1762 2507 1796 2513
rect 1762 2479 1796 2507
rect 1762 2439 1796 2441
rect 1762 2407 1796 2439
rect 1762 2337 1796 2369
rect 1762 2335 1796 2337
rect 1762 2269 1796 2297
rect 1762 2263 1796 2269
rect 1762 2201 1796 2225
rect 1762 2191 1796 2201
rect 1762 2133 1796 2153
rect 1762 2119 1796 2133
rect 1762 2065 1796 2081
rect 1762 2047 1796 2065
rect 1762 1997 1796 2009
rect 1762 1975 1796 1997
rect 1762 1929 1796 1937
rect 1762 1903 1796 1929
rect 1762 1861 1796 1865
rect 1762 1831 1796 1861
rect 1762 1759 1796 1793
rect 1762 1691 1796 1721
rect 1762 1687 1796 1691
rect 1762 1623 1796 1649
rect 1762 1615 1796 1623
rect 1762 1555 1796 1577
rect 1762 1543 1796 1555
rect 1762 1487 1796 1505
rect 1762 1471 1796 1487
rect 1762 1419 1796 1433
rect 1762 1399 1796 1419
rect 1762 1351 1796 1361
rect 1762 1327 1796 1351
rect 1762 1283 1796 1289
rect 1762 1255 1796 1283
rect 1762 1215 1796 1217
rect 1762 1183 1796 1215
rect 1762 1113 1796 1145
rect 1762 1111 1796 1113
rect 1762 1045 1796 1073
rect 1762 1039 1796 1045
rect 1762 977 1796 1001
rect 1762 967 1796 977
rect 1762 909 1796 929
rect 1762 895 1796 909
rect 1762 841 1796 857
rect 1762 823 1796 841
rect 1762 773 1796 785
rect 1762 751 1796 773
rect 1762 705 1796 713
rect 1762 679 1796 705
rect 1762 637 1796 641
rect 1762 607 1796 637
rect 1762 535 1796 569
rect 1762 467 1796 497
rect 1762 463 1796 467
rect 1762 399 1796 425
rect 1762 391 1796 399
rect 1762 331 1796 353
rect 1762 319 1796 331
rect 1762 263 1796 281
rect 1762 247 1796 263
rect 1762 195 1796 209
rect 1762 175 1796 195
rect 1762 127 1796 137
rect 1762 103 1796 127
rect 1762 59 1796 65
rect 1762 31 1796 59
rect -280 -493 -246 -459
rect -206 -493 -172 -459
rect -132 -493 -98 -459
rect -58 -493 -24 -459
rect 16 -493 50 -459
rect 90 -493 124 -459
rect 164 -493 198 -459
rect 238 -493 272 -459
rect 312 -493 346 -459
rect 386 -493 420 -459
rect -280 -567 -246 -533
rect -206 -567 -172 -533
rect -132 -567 -98 -533
rect -58 -567 -24 -533
rect 16 -567 50 -533
rect 90 -567 124 -533
rect 164 -567 198 -533
rect 238 -567 272 -533
rect 312 -567 346 -533
rect 386 -567 420 -533
rect -280 -641 -246 -607
rect -206 -641 -172 -607
rect -132 -641 -98 -607
rect -58 -641 -24 -607
rect 16 -641 50 -607
rect 90 -641 124 -607
rect 164 -641 198 -607
rect 238 -641 272 -607
rect 312 -641 346 -607
rect 386 -641 420 -607
<< metal1 >>
rect -1712 5969 -1112 6200
rect -1712 5935 -1646 5969
rect -1612 5935 -1112 5969
rect -1712 5897 -1112 5935
rect -1712 5863 -1646 5897
rect -1612 5863 -1112 5897
rect -1712 5825 -1112 5863
rect -1712 5791 -1646 5825
rect -1612 5791 -1112 5825
rect -1712 5753 -1112 5791
rect -1712 5719 -1646 5753
rect -1612 5719 -1112 5753
rect -1712 5681 -1112 5719
rect -1712 5647 -1646 5681
rect -1612 5647 -1112 5681
rect -1712 5609 -1112 5647
rect -1712 5575 -1646 5609
rect -1612 5575 -1112 5609
rect -1712 5537 -1112 5575
rect -1712 5503 -1646 5537
rect -1612 5503 -1112 5537
rect -1712 5465 -1112 5503
rect -1712 5431 -1646 5465
rect -1612 5431 -1112 5465
rect -1712 5393 -1112 5431
rect -1712 5359 -1646 5393
rect -1612 5359 -1112 5393
rect -1712 5321 -1112 5359
rect -1712 5287 -1646 5321
rect -1612 5287 -1112 5321
rect -1712 5249 -1112 5287
rect -1712 5215 -1646 5249
rect -1612 5215 -1112 5249
rect -1712 5177 -1112 5215
rect -1712 5143 -1646 5177
rect -1612 5143 -1112 5177
rect -1712 5105 -1112 5143
rect -1712 5071 -1646 5105
rect -1612 5071 -1112 5105
rect -1712 5033 -1112 5071
rect -1712 4999 -1646 5033
rect -1612 4999 -1112 5033
rect -1712 4961 -1112 4999
rect -1712 4927 -1646 4961
rect -1612 4927 -1112 4961
rect -1712 4889 -1112 4927
rect -1712 4855 -1646 4889
rect -1612 4855 -1112 4889
rect -1712 4817 -1112 4855
rect -1712 4783 -1646 4817
rect -1612 4783 -1112 4817
rect -1712 4745 -1112 4783
rect -1712 4711 -1646 4745
rect -1612 4711 -1112 4745
rect -1712 4673 -1112 4711
rect -1712 4639 -1646 4673
rect -1612 4639 -1112 4673
rect -1712 4601 -1112 4639
rect -1712 4567 -1646 4601
rect -1612 4567 -1112 4601
rect -1712 4529 -1112 4567
rect -1712 4495 -1646 4529
rect -1612 4495 -1112 4529
rect -1712 4457 -1112 4495
rect -1712 4423 -1646 4457
rect -1612 4423 -1112 4457
rect -1712 4385 -1112 4423
rect -1712 4351 -1646 4385
rect -1612 4351 -1112 4385
rect -1712 4313 -1112 4351
rect -1712 4279 -1646 4313
rect -1612 4279 -1112 4313
rect -1712 4241 -1112 4279
rect -1712 4207 -1646 4241
rect -1612 4207 -1112 4241
rect -1712 4169 -1112 4207
rect -1712 4135 -1646 4169
rect -1612 4135 -1112 4169
rect -1712 4097 -1112 4135
rect -1712 4063 -1646 4097
rect -1612 4063 -1112 4097
rect -1712 4025 -1112 4063
rect -1712 3991 -1646 4025
rect -1612 3991 -1112 4025
rect -1712 3953 -1112 3991
rect -1712 3919 -1646 3953
rect -1612 3919 -1112 3953
rect -1712 3881 -1112 3919
rect -1712 3847 -1646 3881
rect -1612 3847 -1112 3881
rect -1712 3809 -1112 3847
rect -1712 3775 -1646 3809
rect -1612 3775 -1112 3809
rect -1712 3737 -1112 3775
rect -1712 3703 -1646 3737
rect -1612 3703 -1112 3737
rect -1712 3665 -1112 3703
rect -1712 3631 -1646 3665
rect -1612 3631 -1112 3665
rect -1712 3593 -1112 3631
rect -1712 3559 -1646 3593
rect -1612 3559 -1112 3593
rect -1712 3521 -1112 3559
rect -1712 3487 -1646 3521
rect -1612 3487 -1112 3521
rect -1712 3449 -1112 3487
rect -1712 3415 -1646 3449
rect -1612 3415 -1112 3449
rect -1712 3377 -1112 3415
rect -1712 3343 -1646 3377
rect -1612 3343 -1112 3377
rect -1712 3305 -1112 3343
rect -1712 3271 -1646 3305
rect -1612 3271 -1112 3305
rect -1712 3233 -1112 3271
rect -1712 3199 -1646 3233
rect -1612 3199 -1112 3233
rect -1712 3161 -1112 3199
rect -1712 3127 -1646 3161
rect -1612 3127 -1112 3161
rect -1712 3089 -1112 3127
rect -1712 3055 -1646 3089
rect -1612 3055 -1112 3089
rect -1712 3017 -1112 3055
rect -1712 2983 -1646 3017
rect -1612 2983 -1112 3017
rect -1712 2945 -1112 2983
rect -1712 2911 -1646 2945
rect -1612 2911 -1112 2945
rect -1712 2873 -1112 2911
rect -1712 2839 -1646 2873
rect -1612 2839 -1112 2873
rect -1712 2801 -1112 2839
rect -1712 2767 -1646 2801
rect -1612 2767 -1112 2801
rect -1712 2729 -1112 2767
rect -1712 2695 -1646 2729
rect -1612 2695 -1112 2729
rect -1712 2657 -1112 2695
rect -1712 2623 -1646 2657
rect -1612 2623 -1112 2657
rect -1712 2585 -1112 2623
rect -1712 2551 -1646 2585
rect -1612 2551 -1112 2585
rect -1712 2513 -1112 2551
rect -1712 2479 -1646 2513
rect -1612 2479 -1112 2513
rect -1712 2441 -1112 2479
rect -1712 2407 -1646 2441
rect -1612 2407 -1112 2441
rect -1712 2369 -1112 2407
rect -1712 2335 -1646 2369
rect -1612 2335 -1112 2369
rect -1712 2297 -1112 2335
rect -1712 2263 -1646 2297
rect -1612 2263 -1112 2297
rect -1712 2225 -1112 2263
rect -1712 2191 -1646 2225
rect -1612 2191 -1112 2225
rect -1712 2153 -1112 2191
rect -1712 2119 -1646 2153
rect -1612 2119 -1112 2153
rect -1712 2081 -1112 2119
rect -1712 2047 -1646 2081
rect -1612 2047 -1112 2081
rect -1712 2009 -1112 2047
rect -1712 1975 -1646 2009
rect -1612 1975 -1112 2009
rect -1712 1937 -1112 1975
rect -1712 1903 -1646 1937
rect -1612 1903 -1112 1937
rect -1712 1865 -1112 1903
rect -1712 1831 -1646 1865
rect -1612 1831 -1112 1865
rect -1712 1793 -1112 1831
rect -1712 1759 -1646 1793
rect -1612 1759 -1112 1793
rect -1712 1721 -1112 1759
rect -1712 1687 -1646 1721
rect -1612 1687 -1112 1721
rect -1712 1649 -1112 1687
rect -1712 1615 -1646 1649
rect -1612 1615 -1112 1649
rect -1712 1577 -1112 1615
rect -1712 1543 -1646 1577
rect -1612 1543 -1112 1577
rect -1712 1505 -1112 1543
rect -1712 1471 -1646 1505
rect -1612 1471 -1112 1505
rect -1712 1433 -1112 1471
rect -1712 1399 -1646 1433
rect -1612 1399 -1112 1433
rect -1712 1361 -1112 1399
rect -1712 1327 -1646 1361
rect -1612 1327 -1112 1361
rect -1712 1289 -1112 1327
rect -1712 1255 -1646 1289
rect -1612 1255 -1112 1289
rect -1712 1217 -1112 1255
rect -1712 1183 -1646 1217
rect -1612 1183 -1112 1217
rect -1712 1145 -1112 1183
rect -1712 1111 -1646 1145
rect -1612 1111 -1112 1145
rect -1712 1073 -1112 1111
rect -1712 1039 -1646 1073
rect -1612 1039 -1112 1073
rect -1712 1001 -1112 1039
rect -1712 967 -1646 1001
rect -1612 967 -1112 1001
rect -1712 929 -1112 967
rect -1712 895 -1646 929
rect -1612 895 -1112 929
rect -1712 857 -1112 895
rect -1712 823 -1646 857
rect -1612 823 -1112 857
rect -1712 785 -1112 823
rect -1712 751 -1646 785
rect -1612 751 -1112 785
rect -1712 713 -1112 751
rect -1712 679 -1646 713
rect -1612 679 -1112 713
rect -1712 641 -1112 679
rect -1712 607 -1646 641
rect -1612 607 -1112 641
rect -1712 569 -1112 607
rect -1712 535 -1646 569
rect -1612 535 -1112 569
rect -1712 497 -1112 535
rect -1712 463 -1646 497
rect -1612 463 -1112 497
rect -1712 425 -1112 463
rect -1712 391 -1646 425
rect -1612 391 -1112 425
rect -1712 353 -1112 391
rect -1712 319 -1646 353
rect -1612 319 -1112 353
rect -1712 281 -1112 319
rect -1712 247 -1646 281
rect -1612 247 -1112 281
rect -1712 209 -1112 247
rect -1712 175 -1646 209
rect -1612 175 -1112 209
rect -1712 137 -1112 175
rect -1712 103 -1646 137
rect -1612 103 -1112 137
rect -1712 65 -1112 103
rect -1712 31 -1646 65
rect -1612 31 -1112 65
rect -1712 -200 -1112 31
rect -275 5969 425 6200
rect -275 31 22 5969
rect 128 31 425 5969
rect -275 -200 425 31
rect 1262 5969 1862 6200
rect 1262 5935 1762 5969
rect 1796 5935 1862 5969
rect 1262 5897 1862 5935
rect 1262 5863 1762 5897
rect 1796 5863 1862 5897
rect 1262 5825 1862 5863
rect 1262 5791 1762 5825
rect 1796 5791 1862 5825
rect 1262 5753 1862 5791
rect 1262 5719 1762 5753
rect 1796 5719 1862 5753
rect 1262 5681 1862 5719
rect 1262 5647 1762 5681
rect 1796 5647 1862 5681
rect 1262 5609 1862 5647
rect 1262 5575 1762 5609
rect 1796 5575 1862 5609
rect 1262 5537 1862 5575
rect 1262 5503 1762 5537
rect 1796 5503 1862 5537
rect 1262 5465 1862 5503
rect 1262 5431 1762 5465
rect 1796 5431 1862 5465
rect 1262 5393 1862 5431
rect 1262 5359 1762 5393
rect 1796 5359 1862 5393
rect 1262 5321 1862 5359
rect 1262 5287 1762 5321
rect 1796 5287 1862 5321
rect 1262 5249 1862 5287
rect 1262 5215 1762 5249
rect 1796 5215 1862 5249
rect 1262 5177 1862 5215
rect 1262 5143 1762 5177
rect 1796 5143 1862 5177
rect 1262 5105 1862 5143
rect 1262 5071 1762 5105
rect 1796 5071 1862 5105
rect 1262 5033 1862 5071
rect 1262 4999 1762 5033
rect 1796 4999 1862 5033
rect 1262 4961 1862 4999
rect 1262 4927 1762 4961
rect 1796 4927 1862 4961
rect 1262 4889 1862 4927
rect 1262 4855 1762 4889
rect 1796 4855 1862 4889
rect 1262 4817 1862 4855
rect 1262 4783 1762 4817
rect 1796 4783 1862 4817
rect 1262 4745 1862 4783
rect 1262 4711 1762 4745
rect 1796 4711 1862 4745
rect 1262 4673 1862 4711
rect 1262 4639 1762 4673
rect 1796 4639 1862 4673
rect 1262 4601 1862 4639
rect 1262 4567 1762 4601
rect 1796 4567 1862 4601
rect 1262 4529 1862 4567
rect 1262 4495 1762 4529
rect 1796 4495 1862 4529
rect 1262 4457 1862 4495
rect 1262 4423 1762 4457
rect 1796 4423 1862 4457
rect 1262 4385 1862 4423
rect 1262 4351 1762 4385
rect 1796 4351 1862 4385
rect 1262 4313 1862 4351
rect 1262 4279 1762 4313
rect 1796 4279 1862 4313
rect 1262 4241 1862 4279
rect 1262 4207 1762 4241
rect 1796 4207 1862 4241
rect 1262 4169 1862 4207
rect 1262 4135 1762 4169
rect 1796 4135 1862 4169
rect 1262 4097 1862 4135
rect 1262 4063 1762 4097
rect 1796 4063 1862 4097
rect 1262 4025 1862 4063
rect 1262 3991 1762 4025
rect 1796 3991 1862 4025
rect 1262 3953 1862 3991
rect 1262 3919 1762 3953
rect 1796 3919 1862 3953
rect 1262 3881 1862 3919
rect 1262 3847 1762 3881
rect 1796 3847 1862 3881
rect 1262 3809 1862 3847
rect 1262 3775 1762 3809
rect 1796 3775 1862 3809
rect 1262 3737 1862 3775
rect 1262 3703 1762 3737
rect 1796 3703 1862 3737
rect 1262 3665 1862 3703
rect 1262 3631 1762 3665
rect 1796 3631 1862 3665
rect 1262 3593 1862 3631
rect 1262 3559 1762 3593
rect 1796 3559 1862 3593
rect 1262 3521 1862 3559
rect 1262 3487 1762 3521
rect 1796 3487 1862 3521
rect 1262 3449 1862 3487
rect 1262 3415 1762 3449
rect 1796 3415 1862 3449
rect 1262 3377 1862 3415
rect 1262 3343 1762 3377
rect 1796 3343 1862 3377
rect 1262 3305 1862 3343
rect 1262 3271 1762 3305
rect 1796 3271 1862 3305
rect 1262 3233 1862 3271
rect 1262 3199 1762 3233
rect 1796 3199 1862 3233
rect 1262 3161 1862 3199
rect 1262 3127 1762 3161
rect 1796 3127 1862 3161
rect 1262 3089 1862 3127
rect 1262 3055 1762 3089
rect 1796 3055 1862 3089
rect 1262 3017 1862 3055
rect 1262 2983 1762 3017
rect 1796 2983 1862 3017
rect 1262 2945 1862 2983
rect 1262 2911 1762 2945
rect 1796 2911 1862 2945
rect 1262 2873 1862 2911
rect 1262 2839 1762 2873
rect 1796 2839 1862 2873
rect 1262 2801 1862 2839
rect 1262 2767 1762 2801
rect 1796 2767 1862 2801
rect 1262 2729 1862 2767
rect 1262 2695 1762 2729
rect 1796 2695 1862 2729
rect 1262 2657 1862 2695
rect 1262 2623 1762 2657
rect 1796 2623 1862 2657
rect 1262 2585 1862 2623
rect 1262 2551 1762 2585
rect 1796 2551 1862 2585
rect 1262 2513 1862 2551
rect 1262 2479 1762 2513
rect 1796 2479 1862 2513
rect 1262 2441 1862 2479
rect 1262 2407 1762 2441
rect 1796 2407 1862 2441
rect 1262 2369 1862 2407
rect 1262 2335 1762 2369
rect 1796 2335 1862 2369
rect 1262 2297 1862 2335
rect 1262 2263 1762 2297
rect 1796 2263 1862 2297
rect 1262 2225 1862 2263
rect 1262 2191 1762 2225
rect 1796 2191 1862 2225
rect 1262 2153 1862 2191
rect 1262 2119 1762 2153
rect 1796 2119 1862 2153
rect 1262 2081 1862 2119
rect 1262 2047 1762 2081
rect 1796 2047 1862 2081
rect 1262 2009 1862 2047
rect 1262 1975 1762 2009
rect 1796 1975 1862 2009
rect 1262 1937 1862 1975
rect 1262 1903 1762 1937
rect 1796 1903 1862 1937
rect 1262 1865 1862 1903
rect 1262 1831 1762 1865
rect 1796 1831 1862 1865
rect 1262 1793 1862 1831
rect 1262 1759 1762 1793
rect 1796 1759 1862 1793
rect 1262 1721 1862 1759
rect 1262 1687 1762 1721
rect 1796 1687 1862 1721
rect 1262 1649 1862 1687
rect 1262 1615 1762 1649
rect 1796 1615 1862 1649
rect 1262 1577 1862 1615
rect 1262 1543 1762 1577
rect 1796 1543 1862 1577
rect 1262 1505 1862 1543
rect 1262 1471 1762 1505
rect 1796 1471 1862 1505
rect 1262 1433 1862 1471
rect 1262 1399 1762 1433
rect 1796 1399 1862 1433
rect 1262 1361 1862 1399
rect 1262 1327 1762 1361
rect 1796 1327 1862 1361
rect 1262 1289 1862 1327
rect 1262 1255 1762 1289
rect 1796 1255 1862 1289
rect 1262 1217 1862 1255
rect 1262 1183 1762 1217
rect 1796 1183 1862 1217
rect 1262 1145 1862 1183
rect 1262 1111 1762 1145
rect 1796 1111 1862 1145
rect 1262 1073 1862 1111
rect 1262 1039 1762 1073
rect 1796 1039 1862 1073
rect 1262 1001 1862 1039
rect 1262 967 1762 1001
rect 1796 967 1862 1001
rect 1262 929 1862 967
rect 1262 895 1762 929
rect 1796 895 1862 929
rect 1262 857 1862 895
rect 1262 823 1762 857
rect 1796 823 1862 857
rect 1262 785 1862 823
rect 1262 751 1762 785
rect 1796 751 1862 785
rect 1262 713 1862 751
rect 1262 679 1762 713
rect 1796 679 1862 713
rect 1262 641 1862 679
rect 1262 607 1762 641
rect 1796 607 1862 641
rect 1262 569 1862 607
rect 1262 535 1762 569
rect 1796 535 1862 569
rect 1262 497 1862 535
rect 1262 463 1762 497
rect 1796 463 1862 497
rect 1262 425 1862 463
rect 1262 391 1762 425
rect 1796 391 1862 425
rect 1262 353 1862 391
rect 1262 319 1762 353
rect 1796 319 1862 353
rect 1262 281 1862 319
rect 1262 247 1762 281
rect 1796 247 1862 281
rect 1262 209 1862 247
rect 1262 175 1762 209
rect 1796 175 1862 209
rect 1262 137 1862 175
rect 1262 103 1762 137
rect 1796 103 1862 137
rect 1262 65 1862 103
rect 1262 31 1762 65
rect 1796 31 1862 65
rect 1262 -200 1862 31
rect -296 -450 460 -443
rect -296 -502 -289 -450
rect -237 -502 -215 -450
rect -163 -502 -141 -450
rect -89 -502 -67 -450
rect -15 -502 7 -450
rect 59 -502 81 -450
rect 133 -502 155 -450
rect 207 -502 229 -450
rect 281 -502 303 -450
rect 355 -502 377 -450
rect 429 -502 460 -450
rect -296 -524 460 -502
rect -296 -576 -289 -524
rect -237 -576 -215 -524
rect -163 -576 -141 -524
rect -89 -576 -67 -524
rect -15 -576 7 -524
rect 59 -576 81 -524
rect 133 -576 155 -524
rect 207 -576 229 -524
rect 281 -576 303 -524
rect 355 -576 377 -524
rect 429 -576 460 -524
rect -296 -598 460 -576
rect -296 -650 -289 -598
rect -237 -650 -215 -598
rect -163 -650 -141 -598
rect -89 -650 -67 -598
rect -15 -650 7 -598
rect 59 -650 81 -598
rect 133 -650 155 -598
rect 207 -650 229 -598
rect 281 -650 303 -598
rect 355 -650 377 -598
rect 429 -650 460 -598
rect -296 -657 460 -650
<< via1 >>
rect -289 -459 -237 -450
rect -289 -493 -280 -459
rect -280 -493 -246 -459
rect -246 -493 -237 -459
rect -289 -502 -237 -493
rect -215 -459 -163 -450
rect -215 -493 -206 -459
rect -206 -493 -172 -459
rect -172 -493 -163 -459
rect -215 -502 -163 -493
rect -141 -459 -89 -450
rect -141 -493 -132 -459
rect -132 -493 -98 -459
rect -98 -493 -89 -459
rect -141 -502 -89 -493
rect -67 -459 -15 -450
rect -67 -493 -58 -459
rect -58 -493 -24 -459
rect -24 -493 -15 -459
rect -67 -502 -15 -493
rect 7 -459 59 -450
rect 7 -493 16 -459
rect 16 -493 50 -459
rect 50 -493 59 -459
rect 7 -502 59 -493
rect 81 -459 133 -450
rect 81 -493 90 -459
rect 90 -493 124 -459
rect 124 -493 133 -459
rect 81 -502 133 -493
rect 155 -459 207 -450
rect 155 -493 164 -459
rect 164 -493 198 -459
rect 198 -493 207 -459
rect 155 -502 207 -493
rect 229 -459 281 -450
rect 229 -493 238 -459
rect 238 -493 272 -459
rect 272 -493 281 -459
rect 229 -502 281 -493
rect 303 -459 355 -450
rect 303 -493 312 -459
rect 312 -493 346 -459
rect 346 -493 355 -459
rect 303 -502 355 -493
rect 377 -459 429 -450
rect 377 -493 386 -459
rect 386 -493 420 -459
rect 420 -493 429 -459
rect 377 -502 429 -493
rect -289 -533 -237 -524
rect -289 -567 -280 -533
rect -280 -567 -246 -533
rect -246 -567 -237 -533
rect -289 -576 -237 -567
rect -215 -533 -163 -524
rect -215 -567 -206 -533
rect -206 -567 -172 -533
rect -172 -567 -163 -533
rect -215 -576 -163 -567
rect -141 -533 -89 -524
rect -141 -567 -132 -533
rect -132 -567 -98 -533
rect -98 -567 -89 -533
rect -141 -576 -89 -567
rect -67 -533 -15 -524
rect -67 -567 -58 -533
rect -58 -567 -24 -533
rect -24 -567 -15 -533
rect -67 -576 -15 -567
rect 7 -533 59 -524
rect 7 -567 16 -533
rect 16 -567 50 -533
rect 50 -567 59 -533
rect 7 -576 59 -567
rect 81 -533 133 -524
rect 81 -567 90 -533
rect 90 -567 124 -533
rect 124 -567 133 -533
rect 81 -576 133 -567
rect 155 -533 207 -524
rect 155 -567 164 -533
rect 164 -567 198 -533
rect 198 -567 207 -533
rect 155 -576 207 -567
rect 229 -533 281 -524
rect 229 -567 238 -533
rect 238 -567 272 -533
rect 272 -567 281 -533
rect 229 -576 281 -567
rect 303 -533 355 -524
rect 303 -567 312 -533
rect 312 -567 346 -533
rect 346 -567 355 -533
rect 303 -576 355 -567
rect 377 -533 429 -524
rect 377 -567 386 -533
rect 386 -567 420 -533
rect 420 -567 429 -533
rect 377 -576 429 -567
rect -289 -607 -237 -598
rect -289 -641 -280 -607
rect -280 -641 -246 -607
rect -246 -641 -237 -607
rect -289 -650 -237 -641
rect -215 -607 -163 -598
rect -215 -641 -206 -607
rect -206 -641 -172 -607
rect -172 -641 -163 -607
rect -215 -650 -163 -641
rect -141 -607 -89 -598
rect -141 -641 -132 -607
rect -132 -641 -98 -607
rect -98 -641 -89 -607
rect -141 -650 -89 -641
rect -67 -607 -15 -598
rect -67 -641 -58 -607
rect -58 -641 -24 -607
rect -24 -641 -15 -607
rect -67 -650 -15 -641
rect 7 -607 59 -598
rect 7 -641 16 -607
rect 16 -641 50 -607
rect 50 -641 59 -607
rect 7 -650 59 -641
rect 81 -607 133 -598
rect 81 -641 90 -607
rect 90 -641 124 -607
rect 124 -641 133 -607
rect 81 -650 133 -641
rect 155 -607 207 -598
rect 155 -641 164 -607
rect 164 -641 198 -607
rect 198 -641 207 -607
rect 155 -650 207 -641
rect 229 -607 281 -598
rect 229 -641 238 -607
rect 238 -641 272 -607
rect 272 -641 281 -607
rect 229 -650 281 -641
rect 303 -607 355 -598
rect 303 -641 312 -607
rect 312 -641 346 -607
rect 346 -641 355 -607
rect 303 -650 355 -641
rect 377 -607 429 -598
rect 377 -641 386 -607
rect 386 -641 420 -607
rect 420 -641 429 -607
rect 377 -650 429 -641
<< metal2 >>
rect -296 -450 460 -443
rect -296 -502 -289 -450
rect -237 -502 -215 -450
rect -163 -502 -141 -450
rect -89 -502 -67 -450
rect -15 -502 7 -450
rect 59 -502 81 -450
rect 133 -502 155 -450
rect 207 -502 229 -450
rect 281 -502 303 -450
rect 355 -502 377 -450
rect 429 -502 460 -450
rect -296 -524 460 -502
rect -296 -576 -289 -524
rect -237 -576 -215 -524
rect -163 -576 -141 -524
rect -89 -576 -67 -524
rect -15 -576 7 -524
rect 59 -576 81 -524
rect 133 -576 155 -524
rect 207 -576 229 -524
rect 281 -576 303 -524
rect 355 -576 377 -524
rect 429 -576 460 -524
rect -296 -598 460 -576
rect -296 -650 -289 -598
rect -237 -650 -215 -598
rect -163 -650 -141 -598
rect -89 -650 -67 -598
rect -15 -650 7 -598
rect 59 -650 81 -598
rect 133 -650 155 -598
rect 207 -650 229 -598
rect 281 -650 303 -598
rect 355 -650 377 -598
rect 429 -650 460 -598
rect -296 -657 460 -650
<< labels >>
flabel locali s 1835 6920 1990 6982 0 FreeSans 400 0 0 0 PSUB
port 1 nsew
flabel locali s 1779 28 1779 28 0 FreeSans 400 0 0 0 S
flabel locali s -1630 31 -1630 31 0 FreeSans 400 0 0 0 S
flabel locali s 8 43 142 47 0 FreeSans 400 0 0 0 D
port 2 nsew
flabel comment s 885 159 885 159 0 FreeSans 1600 0 0 0 S
flabel comment s -725 159 -725 159 0 FreeSans 1600 0 0 0 S
flabel comment s 67 159 67 159 0 FreeSans 1600 0 0 0 D
<< properties >>
string GDS_END 7852598
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 7760932
<< end >>
