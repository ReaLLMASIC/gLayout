magic
tech sky130B
timestamp 1701704242
<< metal1 >>
rect 0 0 3 218
rect 93 0 96 218
<< via1 >>
rect 3 0 93 218
<< metal2 >>
rect 0 0 3 218
rect 93 0 96 218
<< properties >>
string GDS_END 78488558
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 78487082
<< end >>
