magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< pwell >>
rect -26 -26 286 1026
<< psubdiff >>
rect 0 930 60 1000
rect 0 896 11 930
rect 45 896 60 930
rect 0 862 60 896
rect 0 828 11 862
rect 45 828 60 862
rect 0 794 60 828
rect 0 760 11 794
rect 45 760 60 794
rect 0 726 60 760
rect 0 692 11 726
rect 45 692 60 726
rect 0 658 60 692
rect 0 624 11 658
rect 45 624 60 658
rect 0 590 60 624
rect 0 556 11 590
rect 45 556 60 590
rect 0 522 60 556
rect 0 488 11 522
rect 45 488 60 522
rect 0 454 60 488
rect 0 420 11 454
rect 45 420 60 454
rect 0 386 60 420
rect 0 352 11 386
rect 45 352 60 386
rect 0 318 60 352
rect 0 284 11 318
rect 45 284 60 318
rect 0 250 60 284
rect 0 216 11 250
rect 45 216 60 250
rect 0 182 60 216
rect 0 148 11 182
rect 45 148 60 182
rect 0 114 60 148
rect 0 80 11 114
rect 45 80 60 114
rect 0 46 60 80
rect 0 12 11 46
rect 45 12 60 46
rect 0 0 60 12
rect 200 930 260 1000
rect 200 896 215 930
rect 249 896 260 930
rect 200 862 260 896
rect 200 828 215 862
rect 249 828 260 862
rect 200 794 260 828
rect 200 760 215 794
rect 249 760 260 794
rect 200 726 260 760
rect 200 692 215 726
rect 249 692 260 726
rect 200 658 260 692
rect 200 624 215 658
rect 249 624 260 658
rect 200 590 260 624
rect 200 556 215 590
rect 249 556 260 590
rect 200 522 260 556
rect 200 488 215 522
rect 249 488 260 522
rect 200 454 260 488
rect 200 420 215 454
rect 249 420 260 454
rect 200 386 260 420
rect 200 352 215 386
rect 249 352 260 386
rect 200 318 260 352
rect 200 284 215 318
rect 249 284 260 318
rect 200 250 260 284
rect 200 216 215 250
rect 249 216 260 250
rect 200 182 260 216
rect 200 148 215 182
rect 249 148 260 182
rect 200 114 260 148
rect 200 80 215 114
rect 249 80 260 114
rect 200 46 260 80
rect 200 12 215 46
rect 249 12 260 46
rect 200 0 260 12
<< nsubdiff >>
rect 60 0 200 1000
<< psubdiffcont >>
rect 11 896 45 930
rect 11 828 45 862
rect 11 760 45 794
rect 11 692 45 726
rect 11 624 45 658
rect 11 556 45 590
rect 11 488 45 522
rect 11 420 45 454
rect 11 352 45 386
rect 11 284 45 318
rect 11 216 45 250
rect 11 148 45 182
rect 11 80 45 114
rect 11 12 45 46
rect 215 896 249 930
rect 215 828 249 862
rect 215 760 249 794
rect 215 692 249 726
rect 215 624 249 658
rect 215 556 249 590
rect 215 488 249 522
rect 215 420 249 454
rect 215 352 249 386
rect 215 284 249 318
rect 215 216 249 250
rect 215 148 249 182
rect 215 80 249 114
rect 215 12 249 46
<< locali >>
rect 11 932 113 966
rect 147 932 249 966
rect 11 930 249 932
rect 45 896 215 930
rect 11 894 249 896
rect 11 862 113 894
rect 45 860 113 862
rect 147 862 249 894
rect 147 860 215 862
rect 45 828 215 860
rect 11 822 249 828
rect 11 794 113 822
rect 45 788 113 794
rect 147 794 249 822
rect 147 788 215 794
rect 45 760 215 788
rect 11 750 249 760
rect 11 726 113 750
rect 45 716 113 726
rect 147 726 249 750
rect 147 716 215 726
rect 45 692 215 716
rect 11 678 249 692
rect 11 658 113 678
rect 45 644 113 658
rect 147 658 249 678
rect 147 644 215 658
rect 45 624 215 644
rect 11 606 249 624
rect 11 590 113 606
rect 45 572 113 590
rect 147 590 249 606
rect 147 572 215 590
rect 45 556 215 572
rect 11 534 249 556
rect 11 522 113 534
rect 45 500 113 522
rect 147 522 249 534
rect 147 500 215 522
rect 45 488 215 500
rect 11 462 249 488
rect 11 454 113 462
rect 45 428 113 454
rect 147 454 249 462
rect 147 428 215 454
rect 45 420 215 428
rect 11 390 249 420
rect 11 386 113 390
rect 45 356 113 386
rect 147 386 249 390
rect 147 356 215 386
rect 45 352 215 356
rect 11 318 249 352
rect 45 284 113 318
rect 147 284 215 318
rect 11 250 249 284
rect 45 246 215 250
rect 45 216 113 246
rect 11 212 113 216
rect 147 216 215 246
rect 147 212 249 216
rect 11 182 249 212
rect 45 174 215 182
rect 45 148 113 174
rect 11 140 113 148
rect 147 148 215 174
rect 147 140 249 148
rect 11 114 249 140
rect 45 102 215 114
rect 45 80 113 102
rect 11 68 113 80
rect 147 80 215 102
rect 147 68 249 80
rect 11 46 249 68
rect 45 30 215 46
rect 45 12 113 30
rect 11 -4 113 12
rect 147 12 215 30
rect 147 -4 249 12
<< viali >>
rect 113 932 147 966
rect 113 860 147 894
rect 113 788 147 822
rect 113 716 147 750
rect 113 644 147 678
rect 113 572 147 606
rect 113 500 147 534
rect 113 428 147 462
rect 113 356 147 390
rect 113 284 147 318
rect 113 212 147 246
rect 113 140 147 174
rect 113 68 147 102
rect 113 -4 147 30
<< metal1 >>
rect 107 966 153 978
rect 107 932 113 966
rect 147 932 153 966
rect 107 894 153 932
rect 107 860 113 894
rect 147 860 153 894
rect 107 822 153 860
rect 107 788 113 822
rect 147 788 153 822
rect 107 750 153 788
rect 107 716 113 750
rect 147 716 153 750
rect 107 678 153 716
rect 107 644 113 678
rect 147 644 153 678
rect 107 606 153 644
rect 107 572 113 606
rect 147 572 153 606
rect 107 534 153 572
rect 107 500 113 534
rect 147 500 153 534
rect 107 462 153 500
rect 107 428 113 462
rect 147 428 153 462
rect 107 390 153 428
rect 107 356 113 390
rect 147 356 153 390
rect 107 318 153 356
rect 107 284 113 318
rect 147 284 153 318
rect 107 246 153 284
rect 107 212 113 246
rect 147 212 153 246
rect 107 174 153 212
rect 107 140 113 174
rect 147 140 153 174
rect 107 102 153 140
rect 107 68 113 102
rect 147 68 153 102
rect 107 30 153 68
rect 107 -4 113 30
rect 147 -4 153 30
rect 107 -16 153 -4
<< properties >>
string GDS_END 12827908
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 12823680
<< end >>
