magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< pwell >>
rect 0 0 952 7015
<< ndiff >>
rect 26 6981 86 6989
rect 26 6947 39 6981
rect 73 6947 86 6981
rect 26 6913 86 6947
rect 26 6879 39 6913
rect 73 6879 86 6913
rect 866 6975 926 6989
rect 866 6941 879 6975
rect 913 6941 926 6975
rect 866 6907 926 6941
rect 866 6873 879 6907
rect 913 6873 926 6907
<< ndiffc >>
rect 39 6947 73 6981
rect 39 6879 73 6913
rect 879 6941 913 6975
rect 879 6873 913 6907
<< ndiffres >>
rect 26 86 86 6879
rect 146 6929 326 6989
rect 146 86 206 6929
rect 26 26 206 86
rect 266 86 326 6929
rect 386 6929 566 6989
rect 386 86 446 6929
rect 266 26 446 86
rect 506 86 566 6929
rect 626 6929 806 6989
rect 626 86 686 6929
rect 506 26 686 86
rect 746 86 806 6929
rect 866 86 926 6873
rect 746 26 926 86
<< locali >>
rect 23 6947 39 6981
rect 73 6947 89 6981
rect 23 6913 89 6947
rect 23 6879 39 6913
rect 73 6879 89 6913
rect 863 6975 929 6981
rect 863 6941 879 6975
rect 913 6941 929 6975
rect 863 6907 929 6941
rect 863 6873 879 6907
rect 913 6873 929 6907
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_0
timestamp 1701704242
transform 0 -1 85 -1 0 6921
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_1
timestamp 1701704242
transform 0 -1 925 -1 0 6983
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_2
timestamp 1701704242
transform 0 -1 85 -1 0 6989
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_3
timestamp 1701704242
transform 0 -1 925 -1 0 6915
box 0 0 1 1
<< properties >>
string GDS_END 6069612
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 6066976
<< end >>
