magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< nwell >>
rect 16 900 1362 2140
<< pwell >>
rect 1290 86 1376 760
rect 42 0 1376 86
<< mvpsubdiff >>
rect 1316 710 1350 734
rect 1316 641 1350 676
rect 1316 572 1350 607
rect 1316 503 1350 538
rect 1316 434 1350 469
rect 1316 364 1350 400
rect 1316 294 1350 330
rect 1316 224 1350 260
rect 1316 154 1350 190
rect 1316 84 1350 120
rect 68 26 92 60
rect 126 26 163 60
rect 197 26 234 60
rect 268 26 305 60
rect 339 26 376 60
rect 410 26 447 60
rect 481 26 518 60
rect 552 26 589 60
rect 623 26 660 60
rect 694 26 730 60
rect 764 26 800 60
rect 834 26 870 60
rect 904 26 940 60
rect 974 26 1010 60
rect 1044 26 1080 60
rect 1114 26 1150 60
rect 1184 26 1220 60
rect 1254 50 1316 60
rect 1254 26 1350 50
<< mvnsubdiff >>
rect 82 2040 106 2074
rect 140 2040 177 2074
rect 211 2040 248 2074
rect 282 2040 319 2074
rect 353 2040 390 2074
rect 424 2040 461 2074
rect 495 2040 532 2074
rect 566 2040 603 2074
rect 637 2040 674 2074
rect 708 2040 745 2074
rect 779 2040 816 2074
rect 850 2040 886 2074
rect 920 2040 956 2074
rect 990 2040 1026 2074
rect 1060 2040 1096 2074
rect 1130 2040 1166 2074
rect 1200 2050 1296 2074
rect 1200 2040 1262 2050
rect 1262 1981 1296 2016
rect 1262 1912 1296 1947
rect 1262 1843 1296 1878
rect 1262 1774 1296 1809
rect 1262 1705 1296 1740
rect 1262 1636 1296 1671
rect 1262 1568 1296 1602
rect 1262 1500 1296 1534
rect 1262 1432 1296 1466
rect 1262 1364 1296 1398
rect 1262 1296 1296 1330
rect 1262 1228 1296 1262
rect 1262 1160 1296 1194
rect 1262 1092 1296 1126
rect 1262 1024 1296 1058
rect 1262 966 1296 990
<< mvpsubdiffcont >>
rect 1316 676 1350 710
rect 1316 607 1350 641
rect 1316 538 1350 572
rect 1316 469 1350 503
rect 1316 400 1350 434
rect 1316 330 1350 364
rect 1316 260 1350 294
rect 1316 190 1350 224
rect 1316 120 1350 154
rect 92 26 126 60
rect 163 26 197 60
rect 234 26 268 60
rect 305 26 339 60
rect 376 26 410 60
rect 447 26 481 60
rect 518 26 552 60
rect 589 26 623 60
rect 660 26 694 60
rect 730 26 764 60
rect 800 26 834 60
rect 870 26 904 60
rect 940 26 974 60
rect 1010 26 1044 60
rect 1080 26 1114 60
rect 1150 26 1184 60
rect 1220 26 1254 60
rect 1316 50 1350 84
<< mvnsubdiffcont >>
rect 106 2040 140 2074
rect 177 2040 211 2074
rect 248 2040 282 2074
rect 319 2040 353 2074
rect 390 2040 424 2074
rect 461 2040 495 2074
rect 532 2040 566 2074
rect 603 2040 637 2074
rect 674 2040 708 2074
rect 745 2040 779 2074
rect 816 2040 850 2074
rect 886 2040 920 2074
rect 956 2040 990 2074
rect 1026 2040 1060 2074
rect 1096 2040 1130 2074
rect 1166 2040 1200 2074
rect 1262 2016 1296 2050
rect 1262 1947 1296 1981
rect 1262 1878 1296 1912
rect 1262 1809 1296 1843
rect 1262 1740 1296 1774
rect 1262 1671 1296 1705
rect 1262 1602 1296 1636
rect 1262 1534 1296 1568
rect 1262 1466 1296 1500
rect 1262 1398 1296 1432
rect 1262 1330 1296 1364
rect 1262 1262 1296 1296
rect 1262 1194 1296 1228
rect 1262 1126 1296 1160
rect 1262 1058 1296 1092
rect 1262 990 1296 1024
<< poly >>
rect 135 826 255 940
rect 311 918 959 940
rect 311 884 705 918
rect 739 884 773 918
rect 807 884 841 918
rect 875 884 909 918
rect 943 884 959 918
rect 311 868 959 884
rect 1015 933 1135 940
rect 79 810 375 826
rect 79 776 155 810
rect 189 776 223 810
rect 257 776 291 810
rect 325 776 375 810
rect 79 760 375 776
rect 541 760 837 868
rect 1015 826 1189 933
rect 893 810 1189 826
rect 893 776 935 810
rect 969 776 1003 810
rect 1037 776 1071 810
rect 1105 776 1139 810
rect 1173 776 1189 810
rect 893 760 1189 776
<< polycont >>
rect 705 884 739 918
rect 773 884 807 918
rect 841 884 875 918
rect 909 884 943 918
rect 155 776 189 810
rect 223 776 257 810
rect 291 776 325 810
rect 935 776 969 810
rect 1003 776 1037 810
rect 1071 776 1105 810
rect 1139 776 1173 810
<< locali >>
rect 82 2040 106 2074
rect 140 2040 177 2074
rect 211 2040 248 2074
rect 282 2040 319 2074
rect 353 2040 390 2074
rect 424 2040 461 2074
rect 495 2040 532 2074
rect 566 2040 603 2074
rect 637 2040 674 2074
rect 708 2040 745 2074
rect 779 2040 816 2074
rect 850 2040 886 2074
rect 920 2040 956 2074
rect 990 2040 1026 2074
rect 1060 2040 1096 2074
rect 1130 2040 1166 2074
rect 1200 2050 1296 2074
rect 1200 2040 1262 2050
rect 90 1912 124 2040
rect 442 1912 476 2040
rect 794 1912 828 2040
rect 1146 1912 1180 2040
rect 1262 1981 1296 2016
rect 1262 1912 1296 1947
rect 1262 1843 1296 1878
rect 1262 1774 1296 1809
rect 300 1676 338 1710
rect 616 1676 654 1710
rect 931 1676 969 1710
rect 1262 1705 1296 1740
rect 1262 1636 1296 1671
rect 1262 1568 1296 1602
rect 1262 1500 1296 1534
rect 1262 1432 1296 1466
rect 90 1336 124 1374
rect 90 1264 124 1302
rect 442 1336 476 1374
rect 442 1264 476 1302
rect 794 1336 828 1374
rect 794 1264 828 1302
rect 1146 1336 1180 1374
rect 1146 1264 1180 1302
rect 1262 1364 1296 1374
rect 1262 1296 1296 1302
rect 1262 1228 1296 1230
rect 1262 1160 1296 1194
rect 1262 1092 1296 1126
rect 34 739 68 777
rect 139 776 155 810
rect 189 776 223 810
rect 257 776 291 810
rect 325 776 341 810
rect 386 739 420 777
rect 618 738 652 1044
rect 1262 1024 1296 1058
rect 1262 966 1296 990
rect 689 884 705 918
rect 739 884 773 918
rect 807 884 841 918
rect 875 884 909 918
rect 943 884 959 918
rect 919 776 935 810
rect 969 776 1003 810
rect 1037 776 1071 810
rect 1105 776 1139 810
rect 1173 776 1189 810
rect 1316 739 1350 777
rect 618 704 689 738
rect 1316 641 1350 676
rect 1316 572 1350 607
rect 1316 503 1350 538
rect 1316 434 1350 469
rect 1316 364 1350 400
rect 1316 294 1350 330
rect 232 241 270 275
rect 986 241 1024 275
rect 1316 224 1350 260
rect 34 195 68 196
rect 34 123 68 161
rect 34 60 68 89
rect 386 195 420 196
rect 386 123 420 161
rect 496 162 530 198
rect 848 162 882 198
rect 1200 162 1234 199
rect 496 128 1234 162
rect 1316 154 1350 161
rect 386 60 420 89
rect 1316 84 1350 89
rect 34 26 92 60
rect 134 26 163 60
rect 206 26 234 60
rect 278 26 305 60
rect 350 26 376 60
rect 410 26 447 60
rect 481 26 518 60
rect 552 26 589 60
rect 623 26 660 60
rect 694 26 730 60
rect 764 26 800 60
rect 834 26 870 60
rect 904 26 940 60
rect 974 26 1010 60
rect 1044 26 1080 60
rect 1114 26 1150 60
rect 1184 26 1220 60
rect 1254 50 1316 60
rect 1254 26 1350 50
<< viali >>
rect 266 1676 300 1710
rect 338 1676 372 1710
rect 582 1676 616 1710
rect 654 1676 688 1710
rect 897 1676 931 1710
rect 969 1676 1003 1710
rect 90 1374 124 1408
rect 90 1302 124 1336
rect 90 1230 124 1264
rect 442 1374 476 1408
rect 442 1302 476 1336
rect 442 1230 476 1264
rect 794 1374 828 1408
rect 794 1302 828 1336
rect 794 1230 828 1264
rect 1146 1374 1180 1408
rect 1146 1302 1180 1336
rect 1146 1230 1180 1264
rect 1262 1398 1296 1408
rect 1262 1374 1296 1398
rect 1262 1330 1296 1336
rect 1262 1302 1296 1330
rect 1262 1262 1296 1264
rect 1262 1230 1296 1262
rect 34 777 68 811
rect 386 777 420 811
rect 34 705 68 739
rect 386 705 420 739
rect 1316 777 1350 811
rect 1316 710 1350 739
rect 1316 705 1350 710
rect 198 241 232 275
rect 270 241 304 275
rect 952 241 986 275
rect 1024 241 1058 275
rect 34 161 68 195
rect 34 89 68 123
rect 386 161 420 195
rect 1316 190 1350 195
rect 1316 161 1350 190
rect 386 89 420 123
rect 1316 120 1350 123
rect 1316 89 1350 120
rect 100 26 126 60
rect 126 26 134 60
rect 172 26 197 60
rect 197 26 206 60
rect 244 26 268 60
rect 268 26 278 60
rect 316 26 339 60
rect 339 26 350 60
<< metal1 >>
rect 254 1710 1015 1716
rect 254 1676 266 1710
rect 300 1676 338 1710
rect 372 1676 582 1710
rect 616 1676 654 1710
rect 688 1676 897 1710
rect 931 1676 969 1710
rect 1003 1676 1015 1710
rect 254 1670 1015 1676
rect -8 1408 1378 1420
rect -8 1374 90 1408
rect 124 1374 442 1408
rect 476 1374 794 1408
rect 828 1374 1146 1408
rect 1180 1374 1262 1408
rect 1296 1374 1378 1408
rect -8 1336 1378 1374
rect -8 1302 90 1336
rect 124 1302 442 1336
rect 476 1302 794 1336
rect 828 1302 1146 1336
rect 1180 1302 1262 1336
rect 1296 1302 1378 1336
rect -8 1264 1378 1302
rect -8 1230 90 1264
rect 124 1230 442 1264
rect 476 1230 794 1264
rect 828 1230 1146 1264
rect 1180 1230 1262 1264
rect 1296 1230 1378 1264
rect -8 1218 1378 1230
rect 28 811 1371 823
rect 28 777 34 811
rect 68 777 386 811
rect 420 777 1316 811
rect 1350 777 1371 811
rect 28 739 1371 777
rect 28 705 34 739
rect 68 705 386 739
rect 420 705 1316 739
rect 1350 705 1371 739
rect 28 693 1371 705
rect 186 275 1070 281
rect 186 241 198 275
rect 232 241 270 275
rect 304 241 952 275
rect 986 241 1024 275
rect 1058 241 1070 275
rect 186 235 1070 241
rect -8 195 1376 207
rect -8 161 34 195
rect 68 161 386 195
rect 420 161 1316 195
rect 1350 161 1376 195
rect -8 123 1376 161
rect -8 89 34 123
rect 68 89 386 123
rect 420 89 1316 123
rect 1350 89 1376 123
rect -8 77 1376 89
rect -8 66 1338 77
tri 1338 66 1349 77 nw
rect -8 60 1292 66
rect -8 26 100 60
rect 134 26 172 60
rect 206 26 244 60
rect 278 26 316 60
rect 350 26 1292 60
rect -8 20 1292 26
tri 1292 20 1338 66 nw
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1701704242
transform 0 1 34 -1 0 195
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1701704242
transform 0 1 386 -1 0 195
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1701704242
transform 0 1 1316 -1 0 195
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_3
timestamp 1701704242
transform 0 1 34 -1 0 811
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_4
timestamp 1701704242
transform 0 1 1316 -1 0 811
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_5
timestamp 1701704242
transform 0 1 386 -1 0 811
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_6
timestamp 1701704242
transform -1 0 1058 0 1 241
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_7
timestamp 1701704242
transform 1 0 266 0 1 1676
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_8
timestamp 1701704242
transform 1 0 198 0 1 241
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_9
timestamp 1701704242
transform 1 0 582 0 1 1676
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_10
timestamp 1701704242
transform 1 0 897 0 1 1676
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_0
timestamp 1701704242
transform 0 -1 1180 -1 0 1408
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_1
timestamp 1701704242
transform 0 -1 828 -1 0 1408
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_2
timestamp 1701704242
transform 0 -1 476 -1 0 1408
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_3
timestamp 1701704242
transform 0 -1 124 -1 0 1408
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_4
timestamp 1701704242
transform 0 -1 1296 -1 0 1408
box 0 0 1 1
use L1M1_CDNS_52468879185191  L1M1_CDNS_52468879185191_0
timestamp 1701704242
transform -1 0 1280 0 1 26
box -12 -6 838 40
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_0
timestamp 1701704242
transform 1 0 100 0 1 26
box 0 0 1 1
use nfet_CDNS_52468879185365  nfet_CDNS_52468879185365_0
timestamp 1701704242
transform -1 0 1189 0 -1 734
box -79 -26 375 626
use nfet_CDNS_52468879185365  nfet_CDNS_52468879185365_1
timestamp 1701704242
transform -1 0 837 0 -1 734
box -79 -26 375 626
use nfet_CDNS_52468879185365  nfet_CDNS_52468879185365_2
timestamp 1701704242
transform -1 0 375 0 -1 734
box -79 -26 375 626
use pfet_CDNS_52468879185313  pfet_CDNS_52468879185313_0
timestamp 1701704242
transform -1 0 431 0 -1 1966
box -119 -66 239 1066
use pfet_CDNS_524688791851428  pfet_CDNS_524688791851428_0
timestamp 1701704242
transform 1 0 487 0 -1 1966
box -119 -66 767 1066
use pfet_CDNS_524688791851429  pfet_CDNS_524688791851429_0
timestamp 1701704242
transform 1 0 135 0 -1 1966
box -119 -66 239 1066
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_0
timestamp 1701704242
transform 0 1 139 1 0 760
box 0 0 1 1
use PYL1_CDNS_52468879185309  PYL1_CDNS_52468879185309_0
timestamp 1701704242
transform 0 1 689 1 0 868
box 0 0 1 1
use PYL1_CDNS_52468879185309  PYL1_CDNS_52468879185309_1
timestamp 1701704242
transform 0 -1 1189 1 0 760
box 0 0 1 1
<< labels >>
flabel metal1 s 53 20 74 207 3 FreeSans 200 0 0 0 vgnd_io
port 1 nsew
flabel metal1 s 711 1670 768 1716 0 FreeSans 200 0 0 0 pu_h_n
port 3 nsew
flabel metal1 s 1366 1218 1378 1420 7 FreeSans 200 0 0 0 vcc_io
port 2 nsew
flabel locali s 223 776 257 810 0 FreeSans 200 180 0 0 slow_h_n
port 5 nsew
flabel locali s 1037 776 1071 810 0 FreeSans 200 180 0 0 puen_h
port 6 nsew
flabel locali s 807 884 841 918 0 FreeSans 200 180 0 0 drvhi_h
port 7 nsew
<< properties >>
string GDS_END 88128816
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 88120364
string path 1.400 51.425 31.975 51.425 31.975 23.500 
<< end >>
