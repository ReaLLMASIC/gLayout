magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< dnwell >>
rect -68 68 10427 5860
<< nwell >>
rect -148 5586 10507 5940
rect -148 342 206 5586
rect 460 596 3152 5332
rect 3406 342 3710 5586
rect 4529 342 4833 5586
rect 10153 342 10507 5586
rect -148 -12 10507 342
<< pwell >>
rect 300 5414 3312 5500
rect 300 514 386 5414
rect 3226 514 3312 5414
rect 300 428 3312 514
rect 3784 1446 3870 2518
rect 4343 1446 4429 2518
rect 4907 5320 10053 5474
rect 4907 3038 5061 5320
rect 9899 3038 10053 5320
rect 4907 2884 10053 3038
rect 4907 608 5061 2884
rect 9899 608 10053 2884
rect 4907 454 10053 608
<< mvpsubdiff >>
rect 326 5440 396 5474
rect 430 5440 464 5474
rect 498 5440 532 5474
rect 566 5440 600 5474
rect 634 5440 668 5474
rect 702 5440 736 5474
rect 770 5440 804 5474
rect 838 5440 872 5474
rect 906 5440 940 5474
rect 974 5440 1008 5474
rect 1042 5440 1076 5474
rect 1110 5440 1144 5474
rect 1178 5440 1212 5474
rect 1246 5440 1280 5474
rect 1314 5440 1348 5474
rect 1382 5440 1416 5474
rect 1450 5440 1484 5474
rect 1518 5440 1552 5474
rect 1586 5440 1620 5474
rect 1654 5440 1688 5474
rect 1722 5440 1756 5474
rect 1790 5440 1824 5474
rect 1858 5440 1892 5474
rect 1926 5440 1960 5474
rect 1994 5440 2028 5474
rect 2062 5440 2096 5474
rect 2130 5440 2164 5474
rect 2198 5440 2232 5474
rect 2266 5440 2300 5474
rect 2334 5440 2368 5474
rect 2402 5440 2436 5474
rect 2470 5440 2504 5474
rect 2538 5440 2572 5474
rect 2606 5440 2640 5474
rect 2674 5440 2708 5474
rect 2742 5440 2776 5474
rect 2810 5440 2844 5474
rect 2878 5440 2912 5474
rect 2946 5440 2980 5474
rect 3014 5440 3048 5474
rect 3082 5440 3116 5474
rect 3150 5440 3184 5474
rect 3218 5440 3286 5474
rect 326 5406 360 5440
rect 326 5338 360 5372
rect 326 5270 360 5304
rect 3252 5384 3286 5440
rect 3252 5316 3286 5350
rect 326 5202 360 5236
rect 326 5134 360 5168
rect 326 5066 360 5100
rect 326 4998 360 5032
rect 326 4930 360 4964
rect 326 4862 360 4896
rect 326 4794 360 4828
rect 326 4726 360 4760
rect 326 4658 360 4692
rect 326 4590 360 4624
rect 326 4522 360 4556
rect 326 4454 360 4488
rect 326 4386 360 4420
rect 326 4318 360 4352
rect 326 4250 360 4284
rect 326 4182 360 4216
rect 326 4114 360 4148
rect 326 4046 360 4080
rect 326 3978 360 4012
rect 326 3910 360 3944
rect 326 3842 360 3876
rect 326 3774 360 3808
rect 326 3706 360 3740
rect 326 3638 360 3672
rect 326 3570 360 3604
rect 326 3502 360 3536
rect 326 3434 360 3468
rect 326 3366 360 3400
rect 326 3298 360 3332
rect 326 3230 360 3264
rect 326 3162 360 3196
rect 326 3094 360 3128
rect 326 3026 360 3060
rect 326 2958 360 2992
rect 326 2890 360 2924
rect 326 2822 360 2856
rect 326 2754 360 2788
rect 326 2686 360 2720
rect 326 2618 360 2652
rect 326 2550 360 2584
rect 326 2482 360 2516
rect 326 2414 360 2448
rect 326 2346 360 2380
rect 326 2278 360 2312
rect 326 2210 360 2244
rect 326 2142 360 2176
rect 326 2074 360 2108
rect 326 2006 360 2040
rect 326 1938 360 1972
rect 326 1870 360 1904
rect 326 1802 360 1836
rect 326 1734 360 1768
rect 326 1666 360 1700
rect 326 1598 360 1632
rect 326 1530 360 1564
rect 326 1462 360 1496
rect 326 1394 360 1428
rect 326 1326 360 1360
rect 326 1258 360 1292
rect 326 1190 360 1224
rect 326 1122 360 1156
rect 326 1054 360 1088
rect 326 986 360 1020
rect 326 918 360 952
rect 326 850 360 884
rect 326 782 360 816
rect 326 714 360 748
rect 326 646 360 680
rect 3252 5248 3286 5282
rect 3252 5180 3286 5214
rect 3252 5112 3286 5146
rect 3252 5044 3286 5078
rect 3252 4976 3286 5010
rect 3252 4908 3286 4942
rect 3252 4840 3286 4874
rect 3252 4772 3286 4806
rect 3252 4704 3286 4738
rect 3252 4636 3286 4670
rect 3252 4568 3286 4602
rect 3252 4500 3286 4534
rect 3252 4432 3286 4466
rect 3252 4364 3286 4398
rect 3252 4296 3286 4330
rect 3252 4228 3286 4262
rect 3252 4160 3286 4194
rect 3252 4092 3286 4126
rect 3252 4024 3286 4058
rect 3252 3956 3286 3990
rect 3252 3888 3286 3922
rect 3252 3820 3286 3854
rect 3252 3752 3286 3786
rect 3252 3684 3286 3718
rect 3252 3616 3286 3650
rect 3252 3548 3286 3582
rect 3252 3480 3286 3514
rect 3252 3412 3286 3446
rect 3252 3344 3286 3378
rect 3252 3276 3286 3310
rect 3252 3208 3286 3242
rect 3252 3140 3286 3174
rect 3252 3072 3286 3106
rect 3252 3004 3286 3038
rect 3252 2936 3286 2970
rect 3252 2868 3286 2902
rect 3252 2800 3286 2834
rect 3252 2732 3286 2766
rect 3252 2664 3286 2698
rect 3252 2596 3286 2630
rect 3252 2528 3286 2562
rect 3252 2460 3286 2494
rect 3252 2392 3286 2426
rect 3252 2324 3286 2358
rect 3252 2256 3286 2290
rect 3252 2188 3286 2222
rect 3252 2120 3286 2154
rect 3252 2052 3286 2086
rect 3252 1984 3286 2018
rect 3252 1916 3286 1950
rect 3252 1848 3286 1882
rect 3252 1780 3286 1814
rect 3252 1712 3286 1746
rect 3252 1644 3286 1678
rect 3252 1576 3286 1610
rect 3252 1508 3286 1542
rect 3252 1440 3286 1474
rect 3252 1372 3286 1406
rect 3252 1304 3286 1338
rect 3252 1236 3286 1270
rect 3252 1168 3286 1202
rect 3252 1100 3286 1134
rect 3252 1032 3286 1066
rect 3252 964 3286 998
rect 3252 896 3286 930
rect 3252 828 3286 862
rect 3252 760 3286 794
rect 3252 692 3286 726
rect 326 488 360 612
rect 3252 624 3286 658
rect 3252 556 3286 590
rect 3252 488 3286 522
rect 326 454 394 488
rect 428 454 462 488
rect 496 454 530 488
rect 564 454 598 488
rect 632 454 666 488
rect 700 454 734 488
rect 768 454 802 488
rect 836 454 870 488
rect 904 454 938 488
rect 972 454 1006 488
rect 1040 454 1074 488
rect 1108 454 1142 488
rect 1176 454 1210 488
rect 1244 454 1278 488
rect 1312 454 1346 488
rect 1380 454 1414 488
rect 1448 454 1482 488
rect 1516 454 1550 488
rect 1584 454 1618 488
rect 1652 454 1686 488
rect 1720 454 1754 488
rect 1788 454 1822 488
rect 1856 454 1890 488
rect 1924 454 1958 488
rect 1992 454 2026 488
rect 2060 454 2094 488
rect 2128 454 2162 488
rect 2196 454 2230 488
rect 2264 454 2298 488
rect 2332 454 2366 488
rect 2400 454 2434 488
rect 2468 454 2502 488
rect 2536 454 2570 488
rect 2604 454 2638 488
rect 2672 454 2706 488
rect 2740 454 2774 488
rect 2808 454 2842 488
rect 2876 454 2910 488
rect 2944 454 2978 488
rect 3012 454 3046 488
rect 3080 454 3114 488
rect 3148 454 3182 488
rect 3216 454 3286 488
rect 3810 2468 3844 2492
rect 3810 2395 3844 2434
rect 3810 2322 3844 2361
rect 3810 2250 3844 2288
rect 3810 2178 3844 2216
rect 3810 2106 3844 2144
rect 3810 2034 3844 2072
rect 3810 1962 3844 2000
rect 3810 1890 3844 1928
rect 3810 1818 3844 1856
rect 3810 1746 3844 1784
rect 3810 1674 3844 1712
rect 3810 1602 3844 1640
rect 3810 1530 3844 1568
rect 3810 1472 3844 1496
rect 4369 2468 4403 2492
rect 4369 2395 4403 2434
rect 4369 2322 4403 2361
rect 4369 2250 4403 2288
rect 4369 2178 4403 2216
rect 4369 2106 4403 2144
rect 4369 2034 4403 2072
rect 4369 1962 4403 2000
rect 4369 1890 4403 1928
rect 4369 1818 4403 1856
rect 4369 1746 4403 1784
rect 4369 1674 4403 1712
rect 4369 1602 4403 1640
rect 4369 1530 4403 1568
rect 4369 1472 4403 1496
rect 4933 5346 5001 5448
rect 9863 5414 9897 5448
rect 9931 5414 10027 5448
rect 9863 5380 10027 5414
rect 9863 5346 9925 5380
rect 4933 5342 5035 5346
rect 4967 5308 5035 5342
rect 4933 5274 5035 5308
rect 5035 2910 5097 3012
rect 9891 2910 10027 2966
rect 9925 2838 10027 2910
rect 9925 594 10027 628
rect 9925 582 9993 594
rect 5035 548 5097 582
rect 4933 514 5097 548
rect 4933 480 5029 514
rect 5063 480 5097 514
rect 9959 560 9993 582
rect 9959 480 10027 560
<< mvnsubdiff >>
rect -22 5724 46 5814
rect 12 5712 46 5724
rect 10212 5780 10246 5814
rect 10280 5780 10381 5814
rect 10212 5746 10381 5780
rect 10212 5712 10279 5746
rect 12 5690 80 5712
rect -22 5656 80 5690
rect 3473 5656 3643 5712
rect 527 5231 603 5265
rect 637 5231 671 5265
rect 527 5197 671 5231
rect 629 5163 671 5197
rect 3017 5185 3085 5265
rect 3017 5163 3051 5185
rect 2983 5151 3051 5163
rect 2983 5117 3085 5151
rect 527 765 629 879
rect 527 663 595 765
rect 2941 731 2983 765
rect 2941 697 3085 731
rect 2941 663 2975 697
rect 3009 663 3085 697
rect 4596 5656 4766 5712
rect 10279 1376 10381 1496
rect 10279 220 10381 254
rect 10279 216 10347 220
rect 80 182 147 216
rect -22 148 147 182
rect -22 114 79 148
rect 113 114 147 148
rect 10313 186 10347 216
rect 10313 114 10381 186
<< mvpsubdiffcont >>
rect 396 5440 430 5474
rect 464 5440 498 5474
rect 532 5440 566 5474
rect 600 5440 634 5474
rect 668 5440 702 5474
rect 736 5440 770 5474
rect 804 5440 838 5474
rect 872 5440 906 5474
rect 940 5440 974 5474
rect 1008 5440 1042 5474
rect 1076 5440 1110 5474
rect 1144 5440 1178 5474
rect 1212 5440 1246 5474
rect 1280 5440 1314 5474
rect 1348 5440 1382 5474
rect 1416 5440 1450 5474
rect 1484 5440 1518 5474
rect 1552 5440 1586 5474
rect 1620 5440 1654 5474
rect 1688 5440 1722 5474
rect 1756 5440 1790 5474
rect 1824 5440 1858 5474
rect 1892 5440 1926 5474
rect 1960 5440 1994 5474
rect 2028 5440 2062 5474
rect 2096 5440 2130 5474
rect 2164 5440 2198 5474
rect 2232 5440 2266 5474
rect 2300 5440 2334 5474
rect 2368 5440 2402 5474
rect 2436 5440 2470 5474
rect 2504 5440 2538 5474
rect 2572 5440 2606 5474
rect 2640 5440 2674 5474
rect 2708 5440 2742 5474
rect 2776 5440 2810 5474
rect 2844 5440 2878 5474
rect 2912 5440 2946 5474
rect 2980 5440 3014 5474
rect 3048 5440 3082 5474
rect 3116 5440 3150 5474
rect 3184 5440 3218 5474
rect 326 5372 360 5406
rect 326 5304 360 5338
rect 326 5236 360 5270
rect 3252 5350 3286 5384
rect 3252 5282 3286 5316
rect 326 5168 360 5202
rect 326 5100 360 5134
rect 326 5032 360 5066
rect 326 4964 360 4998
rect 326 4896 360 4930
rect 326 4828 360 4862
rect 326 4760 360 4794
rect 326 4692 360 4726
rect 326 4624 360 4658
rect 326 4556 360 4590
rect 326 4488 360 4522
rect 326 4420 360 4454
rect 326 4352 360 4386
rect 326 4284 360 4318
rect 326 4216 360 4250
rect 326 4148 360 4182
rect 326 4080 360 4114
rect 326 4012 360 4046
rect 326 3944 360 3978
rect 326 3876 360 3910
rect 326 3808 360 3842
rect 326 3740 360 3774
rect 326 3672 360 3706
rect 326 3604 360 3638
rect 326 3536 360 3570
rect 326 3468 360 3502
rect 326 3400 360 3434
rect 326 3332 360 3366
rect 326 3264 360 3298
rect 326 3196 360 3230
rect 326 3128 360 3162
rect 326 3060 360 3094
rect 326 2992 360 3026
rect 326 2924 360 2958
rect 326 2856 360 2890
rect 326 2788 360 2822
rect 326 2720 360 2754
rect 326 2652 360 2686
rect 326 2584 360 2618
rect 326 2516 360 2550
rect 326 2448 360 2482
rect 326 2380 360 2414
rect 326 2312 360 2346
rect 326 2244 360 2278
rect 326 2176 360 2210
rect 326 2108 360 2142
rect 326 2040 360 2074
rect 326 1972 360 2006
rect 326 1904 360 1938
rect 326 1836 360 1870
rect 326 1768 360 1802
rect 326 1700 360 1734
rect 326 1632 360 1666
rect 326 1564 360 1598
rect 326 1496 360 1530
rect 326 1428 360 1462
rect 326 1360 360 1394
rect 326 1292 360 1326
rect 326 1224 360 1258
rect 326 1156 360 1190
rect 326 1088 360 1122
rect 326 1020 360 1054
rect 326 952 360 986
rect 326 884 360 918
rect 326 816 360 850
rect 326 748 360 782
rect 326 680 360 714
rect 3252 5214 3286 5248
rect 3252 5146 3286 5180
rect 3252 5078 3286 5112
rect 3252 5010 3286 5044
rect 3252 4942 3286 4976
rect 3252 4874 3286 4908
rect 3252 4806 3286 4840
rect 3252 4738 3286 4772
rect 3252 4670 3286 4704
rect 3252 4602 3286 4636
rect 3252 4534 3286 4568
rect 3252 4466 3286 4500
rect 3252 4398 3286 4432
rect 3252 4330 3286 4364
rect 3252 4262 3286 4296
rect 3252 4194 3286 4228
rect 3252 4126 3286 4160
rect 3252 4058 3286 4092
rect 3252 3990 3286 4024
rect 3252 3922 3286 3956
rect 3252 3854 3286 3888
rect 3252 3786 3286 3820
rect 3252 3718 3286 3752
rect 3252 3650 3286 3684
rect 3252 3582 3286 3616
rect 3252 3514 3286 3548
rect 3252 3446 3286 3480
rect 3252 3378 3286 3412
rect 3252 3310 3286 3344
rect 3252 3242 3286 3276
rect 3252 3174 3286 3208
rect 3252 3106 3286 3140
rect 3252 3038 3286 3072
rect 3252 2970 3286 3004
rect 3252 2902 3286 2936
rect 3252 2834 3286 2868
rect 3252 2766 3286 2800
rect 3252 2698 3286 2732
rect 3252 2630 3286 2664
rect 3252 2562 3286 2596
rect 3252 2494 3286 2528
rect 3252 2426 3286 2460
rect 3252 2358 3286 2392
rect 3252 2290 3286 2324
rect 3252 2222 3286 2256
rect 3252 2154 3286 2188
rect 3252 2086 3286 2120
rect 3252 2018 3286 2052
rect 3252 1950 3286 1984
rect 3252 1882 3286 1916
rect 3252 1814 3286 1848
rect 3252 1746 3286 1780
rect 3252 1678 3286 1712
rect 3252 1610 3286 1644
rect 3252 1542 3286 1576
rect 3252 1474 3286 1508
rect 3252 1406 3286 1440
rect 3252 1338 3286 1372
rect 3252 1270 3286 1304
rect 3252 1202 3286 1236
rect 3252 1134 3286 1168
rect 3252 1066 3286 1100
rect 3252 998 3286 1032
rect 3252 930 3286 964
rect 3252 862 3286 896
rect 3252 794 3286 828
rect 3252 726 3286 760
rect 326 612 360 646
rect 3252 658 3286 692
rect 3252 590 3286 624
rect 3252 522 3286 556
rect 394 454 428 488
rect 462 454 496 488
rect 530 454 564 488
rect 598 454 632 488
rect 666 454 700 488
rect 734 454 768 488
rect 802 454 836 488
rect 870 454 904 488
rect 938 454 972 488
rect 1006 454 1040 488
rect 1074 454 1108 488
rect 1142 454 1176 488
rect 1210 454 1244 488
rect 1278 454 1312 488
rect 1346 454 1380 488
rect 1414 454 1448 488
rect 1482 454 1516 488
rect 1550 454 1584 488
rect 1618 454 1652 488
rect 1686 454 1720 488
rect 1754 454 1788 488
rect 1822 454 1856 488
rect 1890 454 1924 488
rect 1958 454 1992 488
rect 2026 454 2060 488
rect 2094 454 2128 488
rect 2162 454 2196 488
rect 2230 454 2264 488
rect 2298 454 2332 488
rect 2366 454 2400 488
rect 2434 454 2468 488
rect 2502 454 2536 488
rect 2570 454 2604 488
rect 2638 454 2672 488
rect 2706 454 2740 488
rect 2774 454 2808 488
rect 2842 454 2876 488
rect 2910 454 2944 488
rect 2978 454 3012 488
rect 3046 454 3080 488
rect 3114 454 3148 488
rect 3182 454 3216 488
rect 3810 2434 3844 2468
rect 3810 2361 3844 2395
rect 3810 2288 3844 2322
rect 3810 2216 3844 2250
rect 3810 2144 3844 2178
rect 3810 2072 3844 2106
rect 3810 2000 3844 2034
rect 3810 1928 3844 1962
rect 3810 1856 3844 1890
rect 3810 1784 3844 1818
rect 3810 1712 3844 1746
rect 3810 1640 3844 1674
rect 3810 1568 3844 1602
rect 3810 1496 3844 1530
rect 4369 2434 4403 2468
rect 4369 2361 4403 2395
rect 4369 2288 4403 2322
rect 4369 2216 4403 2250
rect 4369 2144 4403 2178
rect 4369 2072 4403 2106
rect 4369 2000 4403 2034
rect 4369 1928 4403 1962
rect 4369 1856 4403 1890
rect 4369 1784 4403 1818
rect 4369 1712 4403 1746
rect 4369 1640 4403 1674
rect 4369 1568 4403 1602
rect 4369 1496 4403 1530
rect 5001 5346 9863 5448
rect 9897 5414 9931 5448
rect 4933 5308 4967 5342
rect 4933 548 5035 5274
rect 9925 3012 10027 5380
rect 5097 2966 10027 3012
rect 5097 2910 9891 2966
rect 9925 628 10027 2838
rect 5029 480 5063 514
rect 5097 480 9959 582
rect 9993 560 10027 594
<< mvnsubdiffcont >>
rect -22 5690 12 5724
rect 46 5712 10212 5814
rect 10246 5780 10280 5814
rect -22 182 80 5656
rect 603 5231 637 5265
rect 527 879 629 5197
rect 671 5163 3017 5265
rect 3051 5151 3085 5185
rect 595 663 2941 765
rect 2983 731 3085 5117
rect 2975 663 3009 697
rect 3473 216 3643 5656
rect 4596 216 4766 5656
rect 10279 1496 10381 5746
rect 10279 254 10381 1376
rect 79 114 113 148
rect 147 114 10313 216
rect 10347 186 10381 220
<< poly >>
rect 742 3041 2870 3057
rect 742 3007 758 3041
rect 792 3007 827 3041
rect 861 3007 896 3041
rect 930 3007 965 3041
rect 999 3007 1034 3041
rect 1068 3007 1103 3041
rect 1137 3007 1172 3041
rect 1206 3007 1241 3041
rect 1275 3007 1310 3041
rect 1344 3007 1379 3041
rect 1413 3007 1448 3041
rect 1482 3007 1517 3041
rect 1551 3007 1586 3041
rect 1620 3007 1655 3041
rect 1689 3007 1724 3041
rect 1758 3007 1793 3041
rect 1827 3007 1862 3041
rect 1896 3007 1931 3041
rect 1965 3007 2000 3041
rect 2034 3007 2069 3041
rect 2103 3007 2138 3041
rect 2172 3007 2207 3041
rect 2241 3007 2276 3041
rect 2310 3007 2344 3041
rect 2378 3007 2412 3041
rect 2446 3007 2480 3041
rect 2514 3007 2548 3041
rect 2582 3007 2616 3041
rect 2650 3007 2684 3041
rect 2718 3007 2752 3041
rect 2786 3007 2820 3041
rect 2854 3007 2870 3041
rect 742 2991 2870 3007
rect 742 2921 2870 2937
rect 742 2887 758 2921
rect 792 2887 827 2921
rect 861 2887 896 2921
rect 930 2887 965 2921
rect 999 2887 1034 2921
rect 1068 2887 1103 2921
rect 1137 2887 1172 2921
rect 1206 2887 1241 2921
rect 1275 2887 1310 2921
rect 1344 2887 1379 2921
rect 1413 2887 1448 2921
rect 1482 2887 1517 2921
rect 1551 2887 1586 2921
rect 1620 2887 1655 2921
rect 1689 2887 1724 2921
rect 1758 2887 1793 2921
rect 1827 2887 1862 2921
rect 1896 2887 1931 2921
rect 1965 2887 2000 2921
rect 2034 2887 2069 2921
rect 2103 2887 2138 2921
rect 2172 2887 2207 2921
rect 2241 2887 2276 2921
rect 2310 2887 2344 2921
rect 2378 2887 2412 2921
rect 2446 2887 2480 2921
rect 2514 2887 2548 2921
rect 2582 2887 2616 2921
rect 2650 2887 2684 2921
rect 2718 2887 2752 2921
rect 2786 2887 2820 2921
rect 2854 2887 2870 2921
rect 742 2871 2870 2887
rect 3977 2564 4233 2580
rect 3977 2530 3993 2564
rect 4027 2530 4088 2564
rect 4122 2530 4183 2564
rect 4217 2530 4233 2564
rect 3977 2514 4233 2530
rect 5168 3216 9792 3232
rect 5168 3182 5184 3216
rect 5218 3182 5252 3216
rect 5286 3182 5320 3216
rect 5354 3182 5388 3216
rect 5422 3182 5456 3216
rect 5490 3182 5524 3216
rect 5558 3182 5592 3216
rect 5626 3182 5660 3216
rect 5694 3182 5728 3216
rect 5762 3182 5796 3216
rect 5830 3182 5864 3216
rect 5898 3182 5932 3216
rect 5966 3182 6000 3216
rect 6034 3182 6068 3216
rect 6102 3182 6136 3216
rect 6170 3182 6204 3216
rect 6238 3182 6272 3216
rect 6306 3182 6340 3216
rect 6374 3182 6408 3216
rect 6442 3182 6476 3216
rect 6510 3182 6544 3216
rect 6578 3182 6612 3216
rect 6646 3182 6680 3216
rect 6714 3182 6748 3216
rect 6782 3182 6816 3216
rect 6850 3182 6884 3216
rect 6918 3182 6952 3216
rect 6986 3182 7020 3216
rect 7054 3182 7088 3216
rect 7122 3182 7156 3216
rect 7190 3182 7224 3216
rect 7258 3182 7292 3216
rect 7326 3182 7360 3216
rect 7394 3182 7428 3216
rect 7462 3182 7496 3216
rect 7530 3182 7564 3216
rect 7598 3182 7632 3216
rect 7666 3182 7700 3216
rect 7734 3182 7768 3216
rect 7802 3182 7836 3216
rect 7870 3182 7904 3216
rect 7938 3182 7972 3216
rect 8006 3182 8040 3216
rect 8074 3182 8108 3216
rect 8142 3182 8176 3216
rect 8210 3182 8244 3216
rect 8278 3182 8312 3216
rect 8346 3182 8380 3216
rect 8414 3182 8448 3216
rect 8482 3182 8516 3216
rect 8550 3182 8584 3216
rect 8618 3182 8652 3216
rect 8686 3182 8720 3216
rect 8754 3182 8788 3216
rect 8822 3182 8856 3216
rect 8890 3182 8924 3216
rect 8958 3182 8992 3216
rect 9026 3182 9060 3216
rect 9094 3182 9128 3216
rect 9162 3182 9196 3216
rect 9230 3182 9264 3216
rect 9298 3182 9332 3216
rect 9366 3182 9400 3216
rect 9434 3182 9468 3216
rect 9502 3182 9536 3216
rect 9570 3182 9604 3216
rect 9638 3182 9673 3216
rect 9707 3182 9742 3216
rect 9776 3182 9792 3216
rect 5168 3166 9792 3182
rect 5168 2746 9792 2762
rect 5168 2712 5184 2746
rect 5218 2712 5252 2746
rect 5286 2712 5320 2746
rect 5354 2712 5388 2746
rect 5422 2712 5456 2746
rect 5490 2712 5524 2746
rect 5558 2712 5592 2746
rect 5626 2712 5660 2746
rect 5694 2712 5728 2746
rect 5762 2712 5796 2746
rect 5830 2712 5864 2746
rect 5898 2712 5932 2746
rect 5966 2712 6000 2746
rect 6034 2712 6068 2746
rect 6102 2712 6136 2746
rect 6170 2712 6204 2746
rect 6238 2712 6272 2746
rect 6306 2712 6340 2746
rect 6374 2712 6408 2746
rect 6442 2712 6476 2746
rect 6510 2712 6544 2746
rect 6578 2712 6612 2746
rect 6646 2712 6680 2746
rect 6714 2712 6748 2746
rect 6782 2712 6816 2746
rect 6850 2712 6884 2746
rect 6918 2712 6952 2746
rect 6986 2712 7020 2746
rect 7054 2712 7088 2746
rect 7122 2712 7156 2746
rect 7190 2712 7224 2746
rect 7258 2712 7292 2746
rect 7326 2712 7360 2746
rect 7394 2712 7428 2746
rect 7462 2712 7496 2746
rect 7530 2712 7564 2746
rect 7598 2712 7632 2746
rect 7666 2712 7700 2746
rect 7734 2712 7768 2746
rect 7802 2712 7836 2746
rect 7870 2712 7904 2746
rect 7938 2712 7972 2746
rect 8006 2712 8040 2746
rect 8074 2712 8108 2746
rect 8142 2712 8176 2746
rect 8210 2712 8244 2746
rect 8278 2712 8312 2746
rect 8346 2712 8380 2746
rect 8414 2712 8448 2746
rect 8482 2712 8516 2746
rect 8550 2712 8584 2746
rect 8618 2712 8652 2746
rect 8686 2712 8720 2746
rect 8754 2712 8788 2746
rect 8822 2712 8856 2746
rect 8890 2712 8924 2746
rect 8958 2712 8992 2746
rect 9026 2712 9060 2746
rect 9094 2712 9128 2746
rect 9162 2712 9196 2746
rect 9230 2712 9264 2746
rect 9298 2712 9332 2746
rect 9366 2712 9400 2746
rect 9434 2712 9468 2746
rect 9502 2712 9536 2746
rect 9570 2712 9604 2746
rect 9638 2712 9673 2746
rect 9707 2712 9742 2746
rect 9776 2712 9792 2746
rect 5168 2696 9792 2712
<< polycont >>
rect 758 3007 792 3041
rect 827 3007 861 3041
rect 896 3007 930 3041
rect 965 3007 999 3041
rect 1034 3007 1068 3041
rect 1103 3007 1137 3041
rect 1172 3007 1206 3041
rect 1241 3007 1275 3041
rect 1310 3007 1344 3041
rect 1379 3007 1413 3041
rect 1448 3007 1482 3041
rect 1517 3007 1551 3041
rect 1586 3007 1620 3041
rect 1655 3007 1689 3041
rect 1724 3007 1758 3041
rect 1793 3007 1827 3041
rect 1862 3007 1896 3041
rect 1931 3007 1965 3041
rect 2000 3007 2034 3041
rect 2069 3007 2103 3041
rect 2138 3007 2172 3041
rect 2207 3007 2241 3041
rect 2276 3007 2310 3041
rect 2344 3007 2378 3041
rect 2412 3007 2446 3041
rect 2480 3007 2514 3041
rect 2548 3007 2582 3041
rect 2616 3007 2650 3041
rect 2684 3007 2718 3041
rect 2752 3007 2786 3041
rect 2820 3007 2854 3041
rect 758 2887 792 2921
rect 827 2887 861 2921
rect 896 2887 930 2921
rect 965 2887 999 2921
rect 1034 2887 1068 2921
rect 1103 2887 1137 2921
rect 1172 2887 1206 2921
rect 1241 2887 1275 2921
rect 1310 2887 1344 2921
rect 1379 2887 1413 2921
rect 1448 2887 1482 2921
rect 1517 2887 1551 2921
rect 1586 2887 1620 2921
rect 1655 2887 1689 2921
rect 1724 2887 1758 2921
rect 1793 2887 1827 2921
rect 1862 2887 1896 2921
rect 1931 2887 1965 2921
rect 2000 2887 2034 2921
rect 2069 2887 2103 2921
rect 2138 2887 2172 2921
rect 2207 2887 2241 2921
rect 2276 2887 2310 2921
rect 2344 2887 2378 2921
rect 2412 2887 2446 2921
rect 2480 2887 2514 2921
rect 2548 2887 2582 2921
rect 2616 2887 2650 2921
rect 2684 2887 2718 2921
rect 2752 2887 2786 2921
rect 2820 2887 2854 2921
rect 3993 2530 4027 2564
rect 4088 2530 4122 2564
rect 4183 2530 4217 2564
rect 5184 3182 5218 3216
rect 5252 3182 5286 3216
rect 5320 3182 5354 3216
rect 5388 3182 5422 3216
rect 5456 3182 5490 3216
rect 5524 3182 5558 3216
rect 5592 3182 5626 3216
rect 5660 3182 5694 3216
rect 5728 3182 5762 3216
rect 5796 3182 5830 3216
rect 5864 3182 5898 3216
rect 5932 3182 5966 3216
rect 6000 3182 6034 3216
rect 6068 3182 6102 3216
rect 6136 3182 6170 3216
rect 6204 3182 6238 3216
rect 6272 3182 6306 3216
rect 6340 3182 6374 3216
rect 6408 3182 6442 3216
rect 6476 3182 6510 3216
rect 6544 3182 6578 3216
rect 6612 3182 6646 3216
rect 6680 3182 6714 3216
rect 6748 3182 6782 3216
rect 6816 3182 6850 3216
rect 6884 3182 6918 3216
rect 6952 3182 6986 3216
rect 7020 3182 7054 3216
rect 7088 3182 7122 3216
rect 7156 3182 7190 3216
rect 7224 3182 7258 3216
rect 7292 3182 7326 3216
rect 7360 3182 7394 3216
rect 7428 3182 7462 3216
rect 7496 3182 7530 3216
rect 7564 3182 7598 3216
rect 7632 3182 7666 3216
rect 7700 3182 7734 3216
rect 7768 3182 7802 3216
rect 7836 3182 7870 3216
rect 7904 3182 7938 3216
rect 7972 3182 8006 3216
rect 8040 3182 8074 3216
rect 8108 3182 8142 3216
rect 8176 3182 8210 3216
rect 8244 3182 8278 3216
rect 8312 3182 8346 3216
rect 8380 3182 8414 3216
rect 8448 3182 8482 3216
rect 8516 3182 8550 3216
rect 8584 3182 8618 3216
rect 8652 3182 8686 3216
rect 8720 3182 8754 3216
rect 8788 3182 8822 3216
rect 8856 3182 8890 3216
rect 8924 3182 8958 3216
rect 8992 3182 9026 3216
rect 9060 3182 9094 3216
rect 9128 3182 9162 3216
rect 9196 3182 9230 3216
rect 9264 3182 9298 3216
rect 9332 3182 9366 3216
rect 9400 3182 9434 3216
rect 9468 3182 9502 3216
rect 9536 3182 9570 3216
rect 9604 3182 9638 3216
rect 9673 3182 9707 3216
rect 9742 3182 9776 3216
rect 5184 2712 5218 2746
rect 5252 2712 5286 2746
rect 5320 2712 5354 2746
rect 5388 2712 5422 2746
rect 5456 2712 5490 2746
rect 5524 2712 5558 2746
rect 5592 2712 5626 2746
rect 5660 2712 5694 2746
rect 5728 2712 5762 2746
rect 5796 2712 5830 2746
rect 5864 2712 5898 2746
rect 5932 2712 5966 2746
rect 6000 2712 6034 2746
rect 6068 2712 6102 2746
rect 6136 2712 6170 2746
rect 6204 2712 6238 2746
rect 6272 2712 6306 2746
rect 6340 2712 6374 2746
rect 6408 2712 6442 2746
rect 6476 2712 6510 2746
rect 6544 2712 6578 2746
rect 6612 2712 6646 2746
rect 6680 2712 6714 2746
rect 6748 2712 6782 2746
rect 6816 2712 6850 2746
rect 6884 2712 6918 2746
rect 6952 2712 6986 2746
rect 7020 2712 7054 2746
rect 7088 2712 7122 2746
rect 7156 2712 7190 2746
rect 7224 2712 7258 2746
rect 7292 2712 7326 2746
rect 7360 2712 7394 2746
rect 7428 2712 7462 2746
rect 7496 2712 7530 2746
rect 7564 2712 7598 2746
rect 7632 2712 7666 2746
rect 7700 2712 7734 2746
rect 7768 2712 7802 2746
rect 7836 2712 7870 2746
rect 7904 2712 7938 2746
rect 7972 2712 8006 2746
rect 8040 2712 8074 2746
rect 8108 2712 8142 2746
rect 8176 2712 8210 2746
rect 8244 2712 8278 2746
rect 8312 2712 8346 2746
rect 8380 2712 8414 2746
rect 8448 2712 8482 2746
rect 8516 2712 8550 2746
rect 8584 2712 8618 2746
rect 8652 2712 8686 2746
rect 8720 2712 8754 2746
rect 8788 2712 8822 2746
rect 8856 2712 8890 2746
rect 8924 2712 8958 2746
rect 8992 2712 9026 2746
rect 9060 2712 9094 2746
rect 9128 2712 9162 2746
rect 9196 2712 9230 2746
rect 9264 2712 9298 2746
rect 9332 2712 9366 2746
rect 9400 2712 9434 2746
rect 9468 2712 9502 2746
rect 9536 2712 9570 2746
rect 9604 2712 9638 2746
rect 9673 2712 9707 2746
rect 9742 2712 9776 2746
<< locali >>
rect -30 5816 10389 5822
rect -30 5814 48 5816
rect 82 5814 121 5816
rect 155 5814 194 5816
rect 228 5814 267 5816
rect 301 5814 340 5816
rect 374 5814 413 5816
rect 447 5814 486 5816
rect 520 5814 559 5816
rect 593 5814 632 5816
rect 666 5814 705 5816
rect 739 5814 778 5816
rect 812 5814 851 5816
rect 885 5814 924 5816
rect 958 5814 997 5816
rect 1031 5814 1070 5816
rect 1104 5814 1143 5816
rect 1177 5814 1216 5816
rect 9458 5814 9534 5816
rect 9568 5814 9609 5816
rect 9643 5814 9683 5816
rect 9717 5814 9757 5816
rect 9791 5814 9831 5816
rect 9865 5814 9905 5816
rect 9939 5814 9979 5816
rect 10013 5814 10053 5816
rect 10087 5814 10127 5816
rect 10161 5814 10201 5816
rect 10235 5814 10275 5816
rect -30 5744 46 5814
rect -30 4126 -24 5744
rect 10235 5782 10246 5814
rect 10309 5782 10389 5816
rect 10212 5780 10246 5782
rect 10280 5780 10389 5782
rect 10212 5746 10389 5780
rect 10212 5744 10279 5746
rect 10381 5744 10389 5746
rect 82 5710 121 5712
rect 155 5710 194 5712
rect 228 5710 267 5712
rect 301 5710 340 5712
rect 374 5710 413 5712
rect 447 5710 486 5712
rect 520 5710 559 5712
rect 593 5710 632 5712
rect 666 5710 705 5712
rect 739 5710 778 5712
rect 812 5710 851 5712
rect 885 5710 924 5712
rect 958 5710 997 5712
rect 1031 5710 1070 5712
rect 1104 5710 1143 5712
rect 1177 5710 1216 5712
rect 9458 5710 9534 5712
rect 9568 5710 9609 5712
rect 9643 5710 9683 5712
rect 9717 5710 9757 5712
rect 9791 5710 9831 5712
rect 9865 5710 9905 5712
rect 9939 5710 9979 5712
rect 10013 5710 10053 5712
rect 10087 5710 10127 5712
rect 10161 5710 10201 5712
rect 10235 5710 10277 5744
rect 10383 5710 10389 5744
rect 82 5704 3469 5710
rect 82 4126 88 5704
rect 3463 5638 3469 5704
rect 3647 5704 4592 5710
rect 3647 5638 3653 5704
rect 3463 5599 3473 5638
rect 3643 5599 3653 5638
rect 3463 5565 3469 5599
rect 3647 5565 3653 5599
rect 3463 5526 3473 5565
rect 3643 5526 3653 5565
rect 3463 5492 3469 5526
rect 3647 5492 3653 5526
rect -30 4087 -22 4126
rect 80 4087 88 4126
rect -30 4053 -24 4087
rect 82 4053 88 4087
rect -30 4014 -22 4053
rect 80 4014 88 4053
rect -30 3980 -24 4014
rect 82 3980 88 4014
rect -30 3941 -22 3980
rect 80 3941 88 3980
rect -30 3907 -24 3941
rect 82 3907 88 3941
rect -30 3868 -22 3907
rect 80 3868 88 3907
rect -30 3834 -24 3868
rect 82 3834 88 3868
rect -30 3795 -22 3834
rect 80 3795 88 3834
rect -30 3761 -24 3795
rect 82 3761 88 3795
rect -30 3722 -22 3761
rect 80 3722 88 3761
rect -30 3688 -24 3722
rect 82 3688 88 3722
rect -30 3649 -22 3688
rect 80 3649 88 3688
rect -30 3615 -24 3649
rect 82 3615 88 3649
rect -30 3576 -22 3615
rect 80 3576 88 3615
rect -30 3542 -24 3576
rect 82 3542 88 3576
rect -30 3503 -22 3542
rect 80 3503 88 3542
rect -30 3469 -24 3503
rect 82 3469 88 3503
rect -30 3430 -22 3469
rect 80 3430 88 3469
rect -30 3396 -24 3430
rect 82 3396 88 3430
rect -30 3357 -22 3396
rect 80 3357 88 3396
rect -30 3323 -24 3357
rect 82 3323 88 3357
rect -30 3284 -22 3323
rect 80 3284 88 3323
rect -30 3250 -24 3284
rect 82 3250 88 3284
rect -30 3211 -22 3250
rect 80 3211 88 3250
rect -30 3177 -24 3211
rect 82 3177 88 3211
rect -30 3138 -22 3177
rect 80 3138 88 3177
rect -30 3104 -24 3138
rect 82 3104 88 3138
rect -30 3065 -22 3104
rect 80 3065 88 3104
rect -30 3031 -24 3065
rect 82 3031 88 3065
rect -30 2992 -22 3031
rect 80 2992 88 3031
rect -30 2958 -24 2992
rect 82 2958 88 2992
rect -30 2919 -22 2958
rect 80 2919 88 2958
rect -30 2885 -24 2919
rect 82 2885 88 2919
rect -30 2846 -22 2885
rect 80 2846 88 2885
rect -30 2812 -24 2846
rect 82 2812 88 2846
rect -30 2773 -22 2812
rect 80 2773 88 2812
rect -30 2739 -24 2773
rect 82 2739 88 2773
rect -30 2700 -22 2739
rect 80 2700 88 2739
rect -30 2666 -24 2700
rect 82 2666 88 2700
rect -30 2627 -22 2666
rect 80 2627 88 2666
rect -30 2593 -24 2627
rect 82 2593 88 2627
rect -30 2554 -22 2593
rect 80 2554 88 2593
rect -30 2520 -24 2554
rect 82 2520 88 2554
rect -30 2481 -22 2520
rect 80 2481 88 2520
rect -30 2447 -24 2481
rect 82 2447 88 2481
rect -30 2408 -22 2447
rect 80 2408 88 2447
rect -30 2374 -24 2408
rect 82 2374 88 2408
rect -30 2335 -22 2374
rect 80 2335 88 2374
rect -30 2301 -24 2335
rect 82 2301 88 2335
rect -30 2262 -22 2301
rect 80 2262 88 2301
rect -30 2228 -24 2262
rect 82 2228 88 2262
rect -30 2189 -22 2228
rect 80 2189 88 2228
rect -30 2155 -24 2189
rect 82 2155 88 2189
rect -30 2116 -22 2155
rect 80 2116 88 2155
rect -30 2082 -24 2116
rect 82 2082 88 2116
rect -30 2043 -22 2082
rect 80 2043 88 2082
rect -30 2009 -24 2043
rect 82 2009 88 2043
rect -30 1970 -22 2009
rect 80 1970 88 2009
rect -30 1936 -24 1970
rect 82 1936 88 1970
rect -30 1897 -22 1936
rect 80 1897 88 1936
rect -30 1863 -24 1897
rect 82 1863 88 1897
rect -30 1824 -22 1863
rect 80 1824 88 1863
rect -30 1790 -24 1824
rect 82 1790 88 1824
rect -30 1751 -22 1790
rect 80 1751 88 1790
rect -30 1717 -24 1751
rect 82 1717 88 1751
rect -30 1678 -22 1717
rect 80 1678 88 1717
rect -30 1644 -24 1678
rect 82 1644 88 1678
rect -30 1605 -22 1644
rect 80 1605 88 1644
rect -30 1571 -24 1605
rect 82 1571 88 1605
rect -30 1532 -22 1571
rect 80 1532 88 1571
rect -30 1498 -24 1532
rect 82 1498 88 1532
rect -30 1459 -22 1498
rect 80 1459 88 1498
rect -30 1425 -24 1459
rect 82 1425 88 1459
rect -30 1386 -22 1425
rect 80 1386 88 1425
rect -30 1352 -24 1386
rect 82 1352 88 1386
rect -30 1313 -22 1352
rect 80 1313 88 1352
rect -30 1279 -24 1313
rect 82 1279 88 1313
rect -30 1240 -22 1279
rect 80 1240 88 1279
rect -30 1206 -24 1240
rect 82 1206 88 1240
rect -30 1167 -22 1206
rect 80 1167 88 1206
rect -30 1133 -24 1167
rect 82 1133 88 1167
rect -30 1094 -22 1133
rect 80 1094 88 1133
rect -30 1060 -24 1094
rect 82 1060 88 1094
rect -30 1021 -22 1060
rect 80 1021 88 1060
rect -30 987 -24 1021
rect 82 987 88 1021
rect -30 948 -22 987
rect 80 948 88 987
rect -30 914 -24 948
rect 82 914 88 948
rect -30 875 -22 914
rect 80 875 88 914
rect -30 841 -24 875
rect 82 841 88 875
rect -30 802 -22 841
rect 80 802 88 841
rect -30 768 -24 802
rect 82 768 88 802
rect -30 729 -22 768
rect 80 729 88 768
rect -30 695 -24 729
rect 82 695 88 729
rect -30 656 -22 695
rect 80 656 88 695
rect -30 622 -24 656
rect 82 622 88 656
rect -30 583 -22 622
rect 80 583 88 622
rect -30 549 -24 583
rect 82 549 88 583
rect -30 510 -22 549
rect 80 510 88 549
rect -30 476 -24 510
rect 82 476 88 510
rect -30 437 -22 476
rect 80 437 88 476
rect 320 5474 3293 5480
rect 320 5440 396 5474
rect 442 5440 464 5474
rect 524 5440 532 5474
rect 566 5440 572 5474
rect 634 5440 654 5474
rect 702 5440 736 5474
rect 770 5440 804 5474
rect 853 5440 872 5474
rect 906 5440 929 5474
rect 974 5440 1001 5474
rect 1042 5440 1073 5474
rect 1110 5440 1144 5474
rect 1179 5440 1212 5474
rect 1251 5440 1280 5474
rect 1323 5440 1348 5474
rect 1395 5440 1416 5474
rect 1467 5440 1484 5474
rect 1539 5440 1552 5474
rect 1611 5440 1620 5474
rect 1683 5440 1688 5474
rect 1755 5440 1756 5474
rect 1790 5440 1794 5474
rect 1858 5440 1867 5474
rect 1926 5440 1940 5474
rect 1994 5440 2013 5474
rect 2062 5440 2086 5474
rect 2130 5440 2159 5474
rect 2198 5440 2232 5474
rect 2266 5440 2300 5474
rect 2339 5440 2368 5474
rect 2412 5440 2436 5474
rect 2485 5440 2504 5474
rect 2558 5440 2572 5474
rect 2631 5440 2640 5474
rect 2704 5440 2708 5474
rect 2742 5440 2743 5474
rect 2810 5440 2816 5474
rect 2878 5440 2889 5474
rect 2946 5440 2962 5474
rect 3014 5440 3035 5474
rect 3082 5440 3108 5474
rect 3150 5440 3181 5474
rect 3218 5440 3293 5474
rect 320 5434 3293 5440
rect 320 5406 366 5434
rect 320 5368 326 5406
rect 360 5368 366 5406
rect 320 5338 366 5368
rect 320 5295 326 5338
rect 360 5295 366 5338
rect 320 5270 366 5295
rect 3247 5402 3293 5434
rect 3247 5384 3253 5402
rect 3247 5350 3252 5384
rect 3287 5368 3293 5402
rect 3286 5350 3293 5368
rect 3247 5330 3293 5350
rect 3247 5316 3253 5330
rect 3247 5282 3252 5316
rect 3287 5296 3293 5330
rect 3286 5282 3293 5296
rect 320 5222 326 5270
rect 360 5222 366 5270
rect 320 5202 366 5222
rect 320 5149 326 5202
rect 360 5149 366 5202
rect 320 5134 366 5149
rect 320 5076 326 5134
rect 360 5076 366 5134
rect 320 5066 366 5076
rect 320 5003 326 5066
rect 360 5003 366 5066
rect 320 4998 366 5003
rect 320 4896 326 4998
rect 360 4896 366 4998
rect 320 4891 366 4896
rect 320 4828 326 4891
rect 360 4828 366 4891
rect 320 4818 366 4828
rect 320 4760 326 4818
rect 360 4760 366 4818
rect 320 4745 366 4760
rect 320 4692 326 4745
rect 360 4692 366 4745
rect 320 4672 366 4692
rect 320 4624 326 4672
rect 360 4624 366 4672
rect 320 4599 366 4624
rect 320 4556 326 4599
rect 360 4556 366 4599
rect 320 4526 366 4556
rect 320 4488 326 4526
rect 360 4488 366 4526
rect 320 4454 366 4488
rect 320 4419 326 4454
rect 360 4419 366 4454
rect 320 4386 366 4419
rect 320 4346 326 4386
rect 360 4346 366 4386
rect 320 4318 366 4346
rect 320 4273 326 4318
rect 360 4273 366 4318
rect 320 4250 366 4273
rect 320 4200 326 4250
rect 360 4200 366 4250
rect 320 4182 366 4200
rect 320 4127 326 4182
rect 360 4127 366 4182
rect 320 4114 366 4127
rect 320 4054 326 4114
rect 360 4054 366 4114
rect 320 4046 366 4054
rect 320 3982 326 4046
rect 360 3982 366 4046
rect 320 3978 366 3982
rect 320 3876 326 3978
rect 360 3876 366 3978
rect 320 3872 366 3876
rect 320 3808 326 3872
rect 360 3808 366 3872
rect 320 3800 366 3808
rect 320 3740 326 3800
rect 360 3740 366 3800
rect 320 3728 366 3740
rect 320 3672 326 3728
rect 360 3672 366 3728
rect 320 3656 366 3672
rect 320 3604 326 3656
rect 360 3604 366 3656
rect 320 3584 366 3604
rect 320 3536 326 3584
rect 360 3536 366 3584
rect 320 3512 366 3536
rect 320 3468 326 3512
rect 360 3468 366 3512
rect 320 3440 366 3468
rect 320 3400 326 3440
rect 360 3400 366 3440
rect 320 3368 366 3400
rect 320 3332 326 3368
rect 360 3332 366 3368
rect 320 3298 366 3332
rect 320 3262 326 3298
rect 360 3262 366 3298
rect 320 3230 366 3262
rect 320 3190 326 3230
rect 360 3190 366 3230
rect 320 3162 366 3190
rect 320 3118 326 3162
rect 360 3118 366 3162
rect 320 3094 366 3118
rect 320 3046 326 3094
rect 360 3046 366 3094
rect 320 3026 366 3046
rect 320 2974 326 3026
rect 360 2974 366 3026
rect 320 2958 366 2974
rect 320 2902 326 2958
rect 360 2902 366 2958
rect 320 2890 366 2902
rect 320 2830 326 2890
rect 360 2830 366 2890
rect 320 2822 366 2830
rect 320 2758 326 2822
rect 360 2758 366 2822
rect 320 2754 366 2758
rect 320 2652 326 2754
rect 360 2652 366 2754
rect 320 2648 366 2652
rect 320 2584 326 2648
rect 360 2584 366 2648
rect 320 2576 366 2584
rect 320 2516 326 2576
rect 360 2516 366 2576
rect 320 2504 366 2516
rect 320 2448 326 2504
rect 360 2448 366 2504
rect 320 2432 366 2448
rect 320 2380 326 2432
rect 360 2380 366 2432
rect 320 2360 366 2380
rect 320 2312 326 2360
rect 360 2312 366 2360
rect 320 2288 366 2312
rect 320 2244 326 2288
rect 360 2244 366 2288
rect 320 2216 366 2244
rect 320 2176 326 2216
rect 360 2176 366 2216
rect 320 2144 366 2176
rect 320 2108 326 2144
rect 360 2108 366 2144
rect 320 2074 366 2108
rect 320 2038 326 2074
rect 360 2038 366 2074
rect 320 2006 366 2038
rect 320 1966 326 2006
rect 360 1966 366 2006
rect 320 1938 366 1966
rect 320 1894 326 1938
rect 360 1894 366 1938
rect 320 1870 366 1894
rect 320 1822 326 1870
rect 360 1822 366 1870
rect 320 1802 366 1822
rect 320 1750 326 1802
rect 360 1750 366 1802
rect 320 1734 366 1750
rect 320 1678 326 1734
rect 360 1678 366 1734
rect 320 1666 366 1678
rect 320 1606 326 1666
rect 360 1606 366 1666
rect 320 1598 366 1606
rect 320 1534 326 1598
rect 360 1534 366 1598
rect 320 1530 366 1534
rect 320 1428 326 1530
rect 360 1428 366 1530
rect 320 1424 366 1428
rect 320 1360 326 1424
rect 360 1360 366 1424
rect 320 1352 366 1360
rect 320 1292 326 1352
rect 360 1292 366 1352
rect 320 1280 366 1292
rect 320 1224 326 1280
rect 360 1224 366 1280
rect 320 1208 366 1224
rect 320 1156 326 1208
rect 360 1156 366 1208
rect 320 1136 366 1156
rect 320 1088 326 1136
rect 360 1088 366 1136
rect 320 1064 366 1088
rect 320 1020 326 1064
rect 360 1020 366 1064
rect 320 992 366 1020
rect 320 952 326 992
rect 360 952 366 992
rect 320 920 366 952
rect 320 884 326 920
rect 360 884 366 920
rect 320 850 366 884
rect 320 814 326 850
rect 360 814 366 850
rect 320 782 366 814
rect 320 742 326 782
rect 360 742 366 782
rect 320 714 366 742
rect 320 670 326 714
rect 360 670 366 714
rect 320 646 366 670
rect 519 5274 3093 5280
rect 519 5240 600 5274
rect 634 5265 675 5274
rect 709 5265 750 5274
rect 784 5265 825 5274
rect 859 5265 900 5274
rect 934 5265 976 5274
rect 1010 5265 1052 5274
rect 1086 5265 1128 5274
rect 1162 5265 1204 5274
rect 1238 5265 1280 5274
rect 1314 5265 1356 5274
rect 1390 5265 1432 5274
rect 1466 5265 1508 5274
rect 1542 5265 1584 5274
rect 1618 5265 1660 5274
rect 1694 5265 1736 5274
rect 1770 5265 1846 5274
rect 1880 5265 1921 5274
rect 1955 5265 1996 5274
rect 2030 5265 2071 5274
rect 2105 5265 2146 5274
rect 2180 5265 2221 5274
rect 2255 5265 2297 5274
rect 2331 5265 2373 5274
rect 2407 5265 2449 5274
rect 2483 5265 2525 5274
rect 2559 5265 2601 5274
rect 2635 5265 2677 5274
rect 2711 5265 2753 5274
rect 2787 5265 2829 5274
rect 2863 5265 2905 5274
rect 2939 5265 2981 5274
rect 3015 5265 3093 5274
rect 519 5231 603 5240
rect 637 5231 671 5265
rect 519 5202 671 5231
rect 3017 5202 3093 5265
rect 519 5168 525 5202
rect 559 5197 597 5202
rect 631 5168 671 5202
rect 519 5129 527 5168
rect 629 5163 671 5168
rect 629 5162 2981 5163
rect 629 5129 637 5162
rect 519 5095 525 5129
rect 631 5095 637 5129
rect 519 5056 527 5095
rect 629 5056 637 5095
rect 519 5022 525 5056
rect 631 5022 637 5056
rect 519 4983 527 5022
rect 629 4983 637 5022
rect 519 4949 525 4983
rect 631 4949 637 4983
rect 519 4910 527 4949
rect 629 4910 637 4949
rect 519 4876 525 4910
rect 631 4876 637 4910
rect 519 4837 527 4876
rect 629 4837 637 4876
rect 519 4803 525 4837
rect 631 4803 637 4837
rect 519 4764 527 4803
rect 629 4764 637 4803
rect 519 4730 525 4764
rect 631 4730 637 4764
rect 519 4691 527 4730
rect 629 4691 637 4730
rect 519 4657 525 4691
rect 631 4657 637 4691
rect 519 4618 527 4657
rect 629 4618 637 4657
rect 519 4584 525 4618
rect 631 4584 637 4618
rect 519 4545 527 4584
rect 629 4545 637 4584
rect 519 4511 525 4545
rect 631 4511 637 4545
rect 519 4472 527 4511
rect 629 4472 637 4511
rect 519 4438 525 4472
rect 631 4438 637 4472
rect 519 4399 527 4438
rect 629 4399 637 4438
rect 519 4365 525 4399
rect 631 4365 637 4399
rect 519 4326 527 4365
rect 629 4326 637 4365
rect 519 4292 525 4326
rect 631 4292 637 4326
rect 519 4253 527 4292
rect 629 4253 637 4292
rect 519 4219 525 4253
rect 631 4219 637 4253
rect 519 4180 527 4219
rect 629 4180 637 4219
rect 519 4146 525 4180
rect 631 4146 637 4180
rect 519 4107 527 4146
rect 629 4107 637 4146
rect 519 4073 525 4107
rect 631 4073 637 4107
rect 519 4034 527 4073
rect 629 4034 637 4073
rect 519 4000 525 4034
rect 631 4000 637 4034
rect 519 3961 527 4000
rect 629 3961 637 4000
rect 519 3927 525 3961
rect 631 3927 637 3961
rect 519 3888 527 3927
rect 629 3888 637 3927
rect 519 3854 525 3888
rect 631 3854 637 3888
rect 519 3815 527 3854
rect 629 3815 637 3854
rect 519 3781 525 3815
rect 631 3781 637 3815
rect 519 3742 527 3781
rect 629 3742 637 3781
rect 519 3708 525 3742
rect 631 3708 637 3742
rect 519 3669 527 3708
rect 629 3669 637 3708
rect 519 3635 525 3669
rect 631 3635 637 3669
rect 519 3596 527 3635
rect 629 3596 637 3635
rect 519 3562 525 3596
rect 631 3562 637 3596
rect 519 3523 527 3562
rect 629 3523 637 3562
rect 519 3489 525 3523
rect 631 3489 637 3523
rect 519 3450 527 3489
rect 629 3450 637 3489
rect 519 3416 525 3450
rect 631 3416 637 3450
rect 519 3377 527 3416
rect 629 3377 637 3416
rect 519 3343 525 3377
rect 631 3343 637 3377
rect 519 3304 527 3343
rect 629 3304 637 3343
rect 519 3270 525 3304
rect 631 3270 637 3304
rect 519 3231 527 3270
rect 629 3231 637 3270
rect 519 3197 525 3231
rect 631 3197 637 3231
rect 519 3158 527 3197
rect 629 3158 637 3197
rect 519 3124 525 3158
rect 631 3124 637 3158
rect 519 3085 527 3124
rect 629 3085 637 3124
rect 519 3051 525 3085
rect 631 3051 637 3085
rect 519 3012 527 3051
rect 629 3012 637 3051
rect 2975 4016 2981 5162
rect 3087 4016 3093 5202
rect 2975 3977 2983 4016
rect 3085 3977 3093 4016
rect 2975 3943 2981 3977
rect 3087 3943 3093 3977
rect 2975 3904 2983 3943
rect 3085 3904 3093 3943
rect 2975 3870 2981 3904
rect 3087 3870 3093 3904
rect 2975 3831 2983 3870
rect 3085 3831 3093 3870
rect 2975 3797 2981 3831
rect 3087 3797 3093 3831
rect 2975 3758 2983 3797
rect 3085 3758 3093 3797
rect 2975 3724 2981 3758
rect 3087 3724 3093 3758
rect 2975 3685 2983 3724
rect 3085 3685 3093 3724
rect 2975 3651 2981 3685
rect 3087 3651 3093 3685
rect 2975 3612 2983 3651
rect 3085 3612 3093 3651
rect 2975 3578 2981 3612
rect 3087 3578 3093 3612
rect 2975 3539 2983 3578
rect 3085 3539 3093 3578
rect 2975 3505 2981 3539
rect 3087 3505 3093 3539
rect 2975 3466 2983 3505
rect 3085 3466 3093 3505
rect 2975 3432 2981 3466
rect 3087 3432 3093 3466
rect 2975 3393 2983 3432
rect 3085 3393 3093 3432
rect 2975 3359 2981 3393
rect 3087 3359 3093 3393
rect 2975 3320 2983 3359
rect 3085 3320 3093 3359
rect 2975 3286 2981 3320
rect 3087 3286 3093 3320
rect 2975 3247 2983 3286
rect 3085 3247 3093 3286
rect 2975 3213 2981 3247
rect 3087 3213 3093 3247
rect 2975 3174 2983 3213
rect 3085 3174 3093 3213
rect 2975 3140 2981 3174
rect 3087 3140 3093 3174
rect 2975 3101 2983 3140
rect 3085 3101 3093 3140
rect 2975 3067 2981 3101
rect 3087 3067 3093 3101
rect 519 2978 525 3012
rect 631 2978 637 3012
rect 742 3007 758 3041
rect 808 3007 827 3041
rect 881 3007 896 3041
rect 954 3007 965 3041
rect 1027 3007 1034 3041
rect 1100 3007 1103 3041
rect 1137 3007 1139 3041
rect 1206 3007 1211 3041
rect 1275 3007 1283 3041
rect 1344 3007 1355 3041
rect 1413 3007 1427 3041
rect 1482 3007 1499 3041
rect 1551 3007 1571 3041
rect 1620 3007 1643 3041
rect 1689 3007 1715 3041
rect 1758 3007 1787 3041
rect 1827 3007 1859 3041
rect 1896 3007 1931 3041
rect 1965 3007 2000 3041
rect 2037 3007 2069 3041
rect 2109 3007 2138 3041
rect 2181 3007 2207 3041
rect 2253 3007 2276 3041
rect 2325 3007 2344 3041
rect 2397 3007 2412 3041
rect 2469 3007 2480 3041
rect 2541 3007 2548 3041
rect 2613 3007 2616 3041
rect 2650 3007 2651 3041
rect 2718 3007 2723 3041
rect 2786 3007 2795 3041
rect 2854 3007 2870 3041
rect 2975 3028 2983 3067
rect 3085 3028 3093 3067
rect 519 2939 527 2978
rect 629 2939 637 2978
rect 519 2905 525 2939
rect 631 2905 637 2939
rect 2975 2994 2981 3028
rect 3087 2994 3093 3028
rect 2975 2955 2983 2994
rect 3085 2955 3093 2994
rect 2975 2921 2981 2955
rect 3087 2921 3093 2955
rect 519 2866 527 2905
rect 629 2866 637 2905
rect 742 2887 758 2921
rect 808 2887 827 2921
rect 881 2887 896 2921
rect 954 2887 965 2921
rect 1027 2887 1034 2921
rect 1100 2887 1103 2921
rect 1137 2887 1139 2921
rect 1206 2887 1211 2921
rect 1275 2887 1283 2921
rect 1344 2887 1355 2921
rect 1413 2887 1427 2921
rect 1482 2887 1499 2921
rect 1551 2887 1571 2921
rect 1620 2887 1643 2921
rect 1689 2887 1715 2921
rect 1758 2887 1787 2921
rect 1827 2887 1859 2921
rect 1896 2887 1931 2921
rect 1965 2887 2000 2921
rect 2037 2887 2069 2921
rect 2109 2887 2138 2921
rect 2181 2887 2207 2921
rect 2253 2887 2276 2921
rect 2325 2887 2344 2921
rect 2397 2887 2412 2921
rect 2469 2887 2480 2921
rect 2541 2887 2548 2921
rect 2613 2887 2616 2921
rect 2650 2887 2651 2921
rect 2718 2887 2723 2921
rect 2786 2887 2795 2921
rect 2854 2887 2870 2921
rect 519 2832 525 2866
rect 631 2832 637 2866
rect 519 2793 527 2832
rect 629 2793 637 2832
rect 519 2759 525 2793
rect 631 2759 637 2793
rect 519 2720 527 2759
rect 629 2720 637 2759
rect 519 2686 525 2720
rect 631 2686 637 2720
rect 519 2647 527 2686
rect 629 2647 637 2686
rect 519 2613 525 2647
rect 631 2613 637 2647
rect 519 2574 527 2613
rect 629 2574 637 2613
rect 519 2540 525 2574
rect 631 2540 637 2574
rect 519 2501 527 2540
rect 629 2501 637 2540
rect 519 2467 525 2501
rect 631 2467 637 2501
rect 519 2428 527 2467
rect 629 2428 637 2467
rect 519 2394 525 2428
rect 631 2394 637 2428
rect 519 2355 527 2394
rect 629 2355 637 2394
rect 519 2321 525 2355
rect 631 2321 637 2355
rect 519 2282 527 2321
rect 629 2282 637 2321
rect 519 2248 525 2282
rect 631 2248 637 2282
rect 519 2209 527 2248
rect 629 2209 637 2248
rect 519 2175 525 2209
rect 631 2175 637 2209
rect 519 2136 527 2175
rect 629 2136 637 2175
rect 519 2102 525 2136
rect 631 2102 637 2136
rect 519 2063 527 2102
rect 629 2063 637 2102
rect 519 2029 525 2063
rect 631 2029 637 2063
rect 519 1990 527 2029
rect 629 1990 637 2029
rect 519 1956 525 1990
rect 631 1956 637 1990
rect 519 1917 527 1956
rect 629 1917 637 1956
rect 519 731 525 1917
rect 631 771 637 1917
rect 2975 2882 2983 2921
rect 3085 2882 3093 2921
rect 2975 2848 2981 2882
rect 3087 2848 3093 2882
rect 2975 2809 2983 2848
rect 3085 2809 3093 2848
rect 2975 2775 2981 2809
rect 3087 2775 3093 2809
rect 2975 2736 2983 2775
rect 3085 2736 3093 2775
rect 2975 2702 2981 2736
rect 3087 2702 3093 2736
rect 2975 2663 2983 2702
rect 3085 2663 3093 2702
rect 2975 2629 2981 2663
rect 3087 2629 3093 2663
rect 2975 2590 2983 2629
rect 3085 2590 3093 2629
rect 2975 2556 2981 2590
rect 3087 2556 3093 2590
rect 2975 2517 2983 2556
rect 3085 2517 3093 2556
rect 2975 2483 2981 2517
rect 3087 2483 3093 2517
rect 2975 2444 2983 2483
rect 3085 2444 3093 2483
rect 2975 2410 2981 2444
rect 3087 2410 3093 2444
rect 2975 2371 2983 2410
rect 3085 2371 3093 2410
rect 2975 2337 2981 2371
rect 3087 2337 3093 2371
rect 2975 2298 2983 2337
rect 3085 2298 3093 2337
rect 2975 2264 2981 2298
rect 3087 2264 3093 2298
rect 2975 2225 2983 2264
rect 3085 2225 3093 2264
rect 2975 2191 2981 2225
rect 3087 2191 3093 2225
rect 2975 2152 2983 2191
rect 3085 2152 3093 2191
rect 2975 2118 2981 2152
rect 3087 2118 3093 2152
rect 2975 2079 2983 2118
rect 3085 2079 3093 2118
rect 2975 2045 2981 2079
rect 3087 2045 3093 2079
rect 2975 2006 2983 2045
rect 3085 2006 3093 2045
rect 2975 1972 2981 2006
rect 3087 1972 3093 2006
rect 2975 1933 2983 1972
rect 3085 1933 3093 1972
rect 2975 1899 2981 1933
rect 3087 1899 3093 1933
rect 2975 1860 2983 1899
rect 3085 1860 3093 1899
rect 2975 1826 2981 1860
rect 3087 1826 3093 1860
rect 2975 1787 2983 1826
rect 3085 1787 3093 1826
rect 2975 1753 2981 1787
rect 3087 1753 3093 1787
rect 2975 1714 2983 1753
rect 3085 1714 3093 1753
rect 2975 1680 2981 1714
rect 3087 1680 3093 1714
rect 2975 1641 2983 1680
rect 3085 1641 3093 1680
rect 2975 1607 2981 1641
rect 3087 1607 3093 1641
rect 2975 1568 2983 1607
rect 3085 1568 3093 1607
rect 2975 1534 2981 1568
rect 3087 1534 3093 1568
rect 2975 1495 2983 1534
rect 3085 1495 3093 1534
rect 2975 1461 2981 1495
rect 3087 1461 3093 1495
rect 2975 1422 2983 1461
rect 3085 1422 3093 1461
rect 2975 1388 2981 1422
rect 3087 1388 3093 1422
rect 2975 1349 2983 1388
rect 3085 1349 3093 1388
rect 2975 1315 2981 1349
rect 3087 1315 3093 1349
rect 2975 1276 2983 1315
rect 3085 1276 3093 1315
rect 2975 1242 2981 1276
rect 3087 1242 3093 1276
rect 2975 1203 2983 1242
rect 3085 1203 3093 1242
rect 2975 1169 2981 1203
rect 3087 1169 3093 1203
rect 2975 1130 2983 1169
rect 3085 1130 3093 1169
rect 2975 1096 2981 1130
rect 3087 1096 3093 1130
rect 2975 1057 2983 1096
rect 3085 1057 3093 1096
rect 2975 1023 2981 1057
rect 3087 1023 3093 1057
rect 2975 984 2983 1023
rect 3085 984 3093 1023
rect 2975 950 2981 984
rect 3087 950 3093 984
rect 2975 911 2983 950
rect 3085 911 3093 950
rect 2975 877 2981 911
rect 3087 877 3093 911
rect 2975 838 2983 877
rect 3085 838 3093 877
rect 2975 804 2981 838
rect 3087 804 3093 838
rect 2975 771 2983 804
rect 631 765 2983 771
rect 3085 765 3093 804
rect 519 663 595 731
rect 3087 731 3093 765
rect 519 659 597 663
rect 631 659 670 663
rect 704 659 743 663
rect 777 659 816 663
rect 850 659 889 663
rect 923 659 962 663
rect 996 659 1035 663
rect 1069 659 1108 663
rect 1142 659 1181 663
rect 3015 659 3093 731
rect 519 653 3093 659
rect 3247 5258 3293 5282
rect 3247 5248 3253 5258
rect 3247 5214 3252 5248
rect 3287 5224 3293 5258
rect 3286 5214 3293 5224
rect 3247 5186 3293 5214
rect 3247 5180 3253 5186
rect 3247 5146 3252 5180
rect 3287 5152 3293 5186
rect 3286 5146 3293 5152
rect 3247 5114 3293 5146
rect 3247 5112 3253 5114
rect 3247 5078 3252 5112
rect 3287 5080 3293 5114
rect 3286 5078 3293 5080
rect 3247 5044 3293 5078
rect 3247 5010 3252 5044
rect 3286 5042 3293 5044
rect 3247 5008 3253 5010
rect 3287 5008 3293 5042
rect 3247 4976 3293 5008
rect 3247 4942 3252 4976
rect 3286 4970 3293 4976
rect 3247 4936 3253 4942
rect 3287 4936 3293 4970
rect 3247 4908 3293 4936
rect 3247 4874 3252 4908
rect 3286 4898 3293 4908
rect 3247 4864 3253 4874
rect 3287 4864 3293 4898
rect 3247 4840 3293 4864
rect 3247 4806 3252 4840
rect 3286 4826 3293 4840
rect 3247 4792 3253 4806
rect 3287 4792 3293 4826
rect 3247 4772 3293 4792
rect 3247 4738 3252 4772
rect 3286 4754 3293 4772
rect 3247 4720 3253 4738
rect 3287 4720 3293 4754
rect 3247 4704 3293 4720
rect 3247 4670 3252 4704
rect 3286 4682 3293 4704
rect 3247 4648 3253 4670
rect 3287 4648 3293 4682
rect 3247 4636 3293 4648
rect 3247 4602 3252 4636
rect 3286 4610 3293 4636
rect 3247 4576 3253 4602
rect 3287 4576 3293 4610
rect 3247 4568 3293 4576
rect 3247 4534 3252 4568
rect 3286 4538 3293 4568
rect 3247 4504 3253 4534
rect 3287 4504 3293 4538
rect 3247 4500 3293 4504
rect 3247 4466 3252 4500
rect 3286 4466 3293 4500
rect 3247 4432 3253 4466
rect 3287 4432 3293 4466
rect 3247 4398 3252 4432
rect 3286 4398 3293 4432
rect 3247 4394 3293 4398
rect 3247 4364 3253 4394
rect 3247 4330 3252 4364
rect 3287 4360 3293 4394
rect 3286 4330 3293 4360
rect 3247 4322 3293 4330
rect 3247 4296 3253 4322
rect 3247 4262 3252 4296
rect 3287 4288 3293 4322
rect 3286 4262 3293 4288
rect 3247 4250 3293 4262
rect 3247 4228 3253 4250
rect 3247 4194 3252 4228
rect 3287 4216 3293 4250
rect 3286 4194 3293 4216
rect 3247 4178 3293 4194
rect 3247 4160 3253 4178
rect 3247 4126 3252 4160
rect 3287 4144 3293 4178
rect 3286 4126 3293 4144
rect 3247 4106 3293 4126
rect 3247 4092 3253 4106
rect 3247 4058 3252 4092
rect 3287 4072 3293 4106
rect 3286 4058 3293 4072
rect 3247 4034 3293 4058
rect 3247 4024 3253 4034
rect 3247 3990 3252 4024
rect 3287 4000 3293 4034
rect 3286 3990 3293 4000
rect 3247 3962 3293 3990
rect 3247 3956 3253 3962
rect 3247 3922 3252 3956
rect 3287 3928 3293 3962
rect 3286 3922 3293 3928
rect 3247 3890 3293 3922
rect 3247 3888 3253 3890
rect 3247 3854 3252 3888
rect 3287 3856 3293 3890
rect 3286 3854 3293 3856
rect 3247 3820 3293 3854
rect 3247 3786 3252 3820
rect 3286 3818 3293 3820
rect 3247 3784 3253 3786
rect 3287 3784 3293 3818
rect 3247 3752 3293 3784
rect 3247 3718 3252 3752
rect 3286 3746 3293 3752
rect 3247 3712 3253 3718
rect 3287 3712 3293 3746
rect 3247 3684 3293 3712
rect 3247 3650 3252 3684
rect 3286 3674 3293 3684
rect 3247 3640 3253 3650
rect 3287 3640 3293 3674
rect 3247 3616 3293 3640
rect 3247 3582 3252 3616
rect 3286 3602 3293 3616
rect 3247 3568 3253 3582
rect 3287 3568 3293 3602
rect 3247 3548 3293 3568
rect 3247 3514 3252 3548
rect 3286 3530 3293 3548
rect 3247 3496 3253 3514
rect 3287 3496 3293 3530
rect 3247 3480 3293 3496
rect 3247 3446 3252 3480
rect 3286 3458 3293 3480
rect 3247 3424 3253 3446
rect 3287 3424 3293 3458
rect 3247 3412 3293 3424
rect 3247 3378 3252 3412
rect 3286 3386 3293 3412
rect 3247 3352 3253 3378
rect 3287 3352 3293 3386
rect 3247 3344 3293 3352
rect 3247 3310 3252 3344
rect 3286 3314 3293 3344
rect 3247 3280 3253 3310
rect 3287 3280 3293 3314
rect 3247 3276 3293 3280
rect 3247 3242 3252 3276
rect 3286 3242 3293 3276
rect 3247 3208 3253 3242
rect 3287 3208 3293 3242
rect 3247 3174 3252 3208
rect 3286 3174 3293 3208
rect 3247 3170 3293 3174
rect 3247 3140 3253 3170
rect 3247 3106 3252 3140
rect 3287 3136 3293 3170
rect 3286 3106 3293 3136
rect 3247 3098 3293 3106
rect 3247 3072 3253 3098
rect 3247 3038 3252 3072
rect 3287 3064 3293 3098
rect 3286 3038 3293 3064
rect 3247 3026 3293 3038
rect 3247 3004 3253 3026
rect 3247 2970 3252 3004
rect 3287 2992 3293 3026
rect 3286 2970 3293 2992
rect 3247 2954 3293 2970
rect 3247 2936 3253 2954
rect 3247 2902 3252 2936
rect 3287 2920 3293 2954
rect 3286 2902 3293 2920
rect 3247 2882 3293 2902
rect 3247 2868 3253 2882
rect 3247 2834 3252 2868
rect 3287 2848 3293 2882
rect 3286 2834 3293 2848
rect 3247 2810 3293 2834
rect 3247 2800 3253 2810
rect 3247 2766 3252 2800
rect 3287 2776 3293 2810
rect 3286 2766 3293 2776
rect 3247 2738 3293 2766
rect 3247 2732 3253 2738
rect 3247 2698 3252 2732
rect 3287 2704 3293 2738
rect 3286 2698 3293 2704
rect 3247 2666 3293 2698
rect 3247 2664 3253 2666
rect 3247 2630 3252 2664
rect 3287 2632 3293 2666
rect 3286 2630 3293 2632
rect 3247 2596 3293 2630
rect 3247 2562 3252 2596
rect 3286 2594 3293 2596
rect 3247 2560 3253 2562
rect 3287 2560 3293 2594
rect 3247 2528 3293 2560
rect 3247 2494 3252 2528
rect 3286 2522 3293 2528
rect 3247 2488 3253 2494
rect 3287 2488 3293 2522
rect 3247 2460 3293 2488
rect 3247 2426 3252 2460
rect 3286 2450 3293 2460
rect 3247 2416 3253 2426
rect 3287 2416 3293 2450
rect 3247 2392 3293 2416
rect 3247 2358 3252 2392
rect 3286 2378 3293 2392
rect 3247 2344 3253 2358
rect 3287 2344 3293 2378
rect 3247 2324 3293 2344
rect 3247 2290 3252 2324
rect 3286 2306 3293 2324
rect 3247 2272 3253 2290
rect 3287 2272 3293 2306
rect 3247 2256 3293 2272
rect 3247 2222 3252 2256
rect 3286 2234 3293 2256
rect 3247 2200 3253 2222
rect 3287 2200 3293 2234
rect 3247 2188 3293 2200
rect 3247 2154 3252 2188
rect 3286 2162 3293 2188
rect 3247 2128 3253 2154
rect 3287 2128 3293 2162
rect 3247 2120 3293 2128
rect 3247 2086 3252 2120
rect 3286 2090 3293 2120
rect 3247 2056 3253 2086
rect 3287 2056 3293 2090
rect 3247 2052 3293 2056
rect 3247 2018 3252 2052
rect 3286 2018 3293 2052
rect 3247 1984 3253 2018
rect 3287 1984 3293 2018
rect 3247 1950 3252 1984
rect 3286 1950 3293 1984
rect 3247 1946 3293 1950
rect 3247 1916 3253 1946
rect 3247 1882 3252 1916
rect 3287 1912 3293 1946
rect 3286 1882 3293 1912
rect 3247 1874 3293 1882
rect 3247 1848 3253 1874
rect 3247 1814 3252 1848
rect 3287 1840 3293 1874
rect 3286 1814 3293 1840
rect 3247 1801 3293 1814
rect 3247 1780 3253 1801
rect 3247 1746 3252 1780
rect 3287 1767 3293 1801
rect 3286 1746 3293 1767
rect 3247 1728 3293 1746
rect 3247 1712 3253 1728
rect 3247 1678 3252 1712
rect 3287 1694 3293 1728
rect 3286 1678 3293 1694
rect 3247 1655 3293 1678
rect 3247 1644 3253 1655
rect 3247 1610 3252 1644
rect 3287 1621 3293 1655
rect 3286 1610 3293 1621
rect 3247 1582 3293 1610
rect 3247 1576 3253 1582
rect 3247 1542 3252 1576
rect 3287 1548 3293 1582
rect 3286 1542 3293 1548
rect 3247 1509 3293 1542
rect 3247 1508 3253 1509
rect 3247 1474 3252 1508
rect 3287 1475 3293 1509
rect 3286 1474 3293 1475
rect 3247 1440 3293 1474
rect 3247 1406 3252 1440
rect 3286 1436 3293 1440
rect 3247 1402 3253 1406
rect 3287 1402 3293 1436
rect 3247 1372 3293 1402
rect 3247 1338 3252 1372
rect 3286 1363 3293 1372
rect 3247 1329 3253 1338
rect 3287 1329 3293 1363
rect 3247 1304 3293 1329
rect 3247 1270 3252 1304
rect 3286 1290 3293 1304
rect 3247 1256 3253 1270
rect 3287 1256 3293 1290
rect 3247 1236 3293 1256
rect 3247 1202 3252 1236
rect 3286 1217 3293 1236
rect 3247 1183 3253 1202
rect 3287 1183 3293 1217
rect 3247 1168 3293 1183
rect 3247 1134 3252 1168
rect 3286 1144 3293 1168
rect 3247 1110 3253 1134
rect 3287 1110 3293 1144
rect 3247 1100 3293 1110
rect 3247 1066 3252 1100
rect 3286 1071 3293 1100
rect 3247 1037 3253 1066
rect 3287 1037 3293 1071
rect 3247 1032 3293 1037
rect 3247 998 3252 1032
rect 3286 998 3293 1032
rect 3247 964 3253 998
rect 3287 964 3293 998
rect 3247 930 3252 964
rect 3286 930 3293 964
rect 3247 925 3293 930
rect 3247 896 3253 925
rect 3247 862 3252 896
rect 3287 891 3293 925
rect 3286 862 3293 891
rect 3247 852 3293 862
rect 3247 828 3253 852
rect 3247 794 3252 828
rect 3287 818 3293 852
rect 3286 794 3293 818
rect 3247 779 3293 794
rect 3247 760 3253 779
rect 3247 726 3252 760
rect 3287 745 3293 779
rect 3286 726 3293 745
rect 3247 706 3293 726
rect 3247 692 3253 706
rect 3247 658 3252 692
rect 3287 672 3293 706
rect 3286 658 3293 672
rect 320 598 326 646
rect 360 598 366 646
rect 320 560 366 598
rect 320 526 326 560
rect 360 526 366 560
rect 320 494 366 526
rect 3247 633 3293 658
rect 3247 624 3253 633
rect 3247 590 3252 624
rect 3287 599 3293 633
rect 3286 590 3293 599
rect 3247 560 3293 590
rect 3247 556 3253 560
rect 3247 522 3252 556
rect 3287 526 3293 560
rect 3286 522 3293 526
rect 3247 494 3293 522
rect 320 488 3293 494
rect 320 454 394 488
rect 432 454 462 488
rect 506 454 530 488
rect 580 454 598 488
rect 654 454 666 488
rect 728 454 734 488
rect 836 454 842 488
rect 904 454 916 488
rect 972 454 990 488
rect 1040 454 1063 488
rect 1108 454 1136 488
rect 1176 454 1209 488
rect 1244 454 1278 488
rect 1316 454 1346 488
rect 1389 454 1414 488
rect 1462 454 1482 488
rect 1535 454 1550 488
rect 1608 454 1618 488
rect 1681 454 1686 488
rect 1788 454 1793 488
rect 1856 454 1866 488
rect 1924 454 1939 488
rect 1992 454 2012 488
rect 2060 454 2085 488
rect 2128 454 2158 488
rect 2196 454 2230 488
rect 2265 454 2298 488
rect 2338 454 2366 488
rect 2411 454 2434 488
rect 2484 454 2502 488
rect 2557 454 2570 488
rect 2630 454 2638 488
rect 2703 454 2706 488
rect 2740 454 2742 488
rect 2808 454 2815 488
rect 2876 454 2888 488
rect 2944 454 2961 488
rect 3012 454 3034 488
rect 3080 454 3107 488
rect 3148 454 3180 488
rect 3216 454 3293 488
rect 320 448 3293 454
rect 3463 5453 3473 5492
rect 3643 5453 3653 5492
rect 3463 5419 3469 5453
rect 3647 5419 3653 5453
rect 3463 5380 3473 5419
rect 3643 5380 3653 5419
rect 3463 5346 3469 5380
rect 3647 5346 3653 5380
rect 3463 5307 3473 5346
rect 3643 5307 3653 5346
rect 3463 5273 3469 5307
rect 3647 5273 3653 5307
rect 3463 5234 3473 5273
rect 3643 5234 3653 5273
rect 3463 5200 3469 5234
rect 3647 5200 3653 5234
rect 3463 5161 3473 5200
rect 3643 5161 3653 5200
rect 3463 5127 3469 5161
rect 3647 5127 3653 5161
rect 3463 5088 3473 5127
rect 3643 5088 3653 5127
rect 3463 5054 3469 5088
rect 3647 5054 3653 5088
rect 3463 5015 3473 5054
rect 3643 5015 3653 5054
rect 3463 4981 3469 5015
rect 3647 4981 3653 5015
rect 3463 4942 3473 4981
rect 3643 4942 3653 4981
rect 3463 4908 3469 4942
rect 3647 4908 3653 4942
rect 3463 4869 3473 4908
rect 3643 4869 3653 4908
rect 3463 4835 3469 4869
rect 3647 4835 3653 4869
rect 3463 4796 3473 4835
rect 3643 4796 3653 4835
rect 3463 4762 3469 4796
rect 3647 4762 3653 4796
rect 3463 4723 3473 4762
rect 3643 4723 3653 4762
rect 3463 4689 3469 4723
rect 3647 4689 3653 4723
rect 3463 4650 3473 4689
rect 3643 4650 3653 4689
rect 3463 4616 3469 4650
rect 3647 4616 3653 4650
rect 3463 4577 3473 4616
rect 3643 4577 3653 4616
rect 3463 4543 3469 4577
rect 3647 4543 3653 4577
rect 3463 4504 3473 4543
rect 3643 4504 3653 4543
rect 3463 4470 3469 4504
rect 3647 4470 3653 4504
rect 3463 4431 3473 4470
rect 3643 4431 3653 4470
rect 3463 4397 3469 4431
rect 3647 4397 3653 4431
rect 3463 4358 3473 4397
rect 3643 4358 3653 4397
rect 3463 4324 3469 4358
rect 3647 4324 3653 4358
rect 3463 4285 3473 4324
rect 3643 4285 3653 4324
rect 3463 4251 3469 4285
rect 3647 4251 3653 4285
rect 3463 4212 3473 4251
rect 3643 4212 3653 4251
rect 3463 4178 3469 4212
rect 3647 4178 3653 4212
rect 3463 4139 3473 4178
rect 3643 4139 3653 4178
rect 3463 4105 3469 4139
rect 3647 4105 3653 4139
rect 3463 4066 3473 4105
rect 3643 4066 3653 4105
rect 3463 4032 3469 4066
rect 3647 4032 3653 4066
rect 3463 3993 3473 4032
rect 3643 3993 3653 4032
rect 3463 3959 3469 3993
rect 3647 3959 3653 3993
rect 3463 3920 3473 3959
rect 3643 3920 3653 3959
rect 3463 3886 3469 3920
rect 3647 3886 3653 3920
rect 3463 3847 3473 3886
rect 3643 3847 3653 3886
rect 3463 3813 3469 3847
rect 3647 3813 3653 3847
rect 3463 3774 3473 3813
rect 3643 3774 3653 3813
rect 3463 3740 3469 3774
rect 3647 3740 3653 3774
rect 3463 3701 3473 3740
rect 3643 3701 3653 3740
rect 3463 3667 3469 3701
rect 3647 3667 3653 3701
rect 3463 3628 3473 3667
rect 3643 3628 3653 3667
rect 3463 3594 3469 3628
rect 3647 3594 3653 3628
rect 3463 3555 3473 3594
rect 3643 3555 3653 3594
rect 3463 3521 3469 3555
rect 3647 3521 3653 3555
rect 3463 3482 3473 3521
rect 3643 3482 3653 3521
rect 3463 3448 3469 3482
rect 3647 3448 3653 3482
rect 3463 3409 3473 3448
rect 3643 3409 3653 3448
rect 3463 3375 3469 3409
rect 3647 3375 3653 3409
rect 3463 3336 3473 3375
rect 3643 3336 3653 3375
rect 3463 3302 3469 3336
rect 3647 3302 3653 3336
rect 3463 3263 3473 3302
rect 3643 3263 3653 3302
rect 3463 3229 3469 3263
rect 3647 3229 3653 3263
rect 3463 3190 3473 3229
rect 3643 3190 3653 3229
rect 3463 3156 3469 3190
rect 3647 3156 3653 3190
rect 3463 3117 3473 3156
rect 3643 3117 3653 3156
rect 3463 3083 3469 3117
rect 3647 3083 3653 3117
rect 3463 3044 3473 3083
rect 3643 3044 3653 3083
rect 3463 3010 3469 3044
rect 3647 3010 3653 3044
rect 3463 2971 3473 3010
rect 3643 2971 3653 3010
rect 3463 2937 3469 2971
rect 3647 2937 3653 2971
rect 3463 2898 3473 2937
rect 3643 2898 3653 2937
rect 3463 2864 3469 2898
rect 3647 2864 3653 2898
rect 3463 2825 3473 2864
rect 3643 2825 3653 2864
rect 3463 2791 3469 2825
rect 3647 2791 3653 2825
rect 3463 2752 3473 2791
rect 3643 2752 3653 2791
rect 3463 2718 3469 2752
rect 3647 2718 3653 2752
rect 3463 2679 3473 2718
rect 3643 2679 3653 2718
rect 3463 2645 3469 2679
rect 3647 2645 3653 2679
rect 3463 2606 3473 2645
rect 3643 2606 3653 2645
rect 3463 2572 3469 2606
rect 3647 2572 3653 2606
rect 3463 2533 3473 2572
rect 3643 2533 3653 2572
rect 4586 5638 4592 5704
rect 4770 5704 10279 5710
rect 4770 5638 4776 5704
rect 4586 5599 4596 5638
rect 4766 5599 4776 5638
rect 4586 5565 4592 5599
rect 4770 5565 4776 5599
rect 4586 5526 4596 5565
rect 4766 5526 4776 5565
rect 4586 5492 4592 5526
rect 4770 5492 4776 5526
rect 4586 5453 4596 5492
rect 4766 5453 4776 5492
rect 10271 5671 10279 5704
rect 10381 5671 10389 5710
rect 10271 5637 10277 5671
rect 10383 5637 10389 5671
rect 10271 5598 10279 5637
rect 10381 5598 10389 5637
rect 10271 5564 10277 5598
rect 10383 5564 10389 5598
rect 10271 5525 10279 5564
rect 10381 5525 10389 5564
rect 10271 5491 10277 5525
rect 10383 5491 10389 5525
rect 4586 5419 4592 5453
rect 4770 5419 4776 5453
rect 4586 5380 4596 5419
rect 4766 5380 4776 5419
rect 4586 5346 4592 5380
rect 4770 5346 4776 5380
rect 4586 5307 4596 5346
rect 4766 5307 4776 5346
rect 4586 5273 4592 5307
rect 4770 5273 4776 5307
rect 4586 5234 4596 5273
rect 4766 5234 4776 5273
rect 4586 5200 4592 5234
rect 4770 5200 4776 5234
rect 4586 5161 4596 5200
rect 4766 5161 4776 5200
rect 4586 5127 4592 5161
rect 4770 5127 4776 5161
rect 4586 5088 4596 5127
rect 4766 5088 4776 5127
rect 4586 5054 4592 5088
rect 4770 5054 4776 5088
rect 4586 5015 4596 5054
rect 4766 5015 4776 5054
rect 4586 4981 4592 5015
rect 4770 4981 4776 5015
rect 4586 4942 4596 4981
rect 4766 4942 4776 4981
rect 4586 4908 4592 4942
rect 4770 4908 4776 4942
rect 4586 4869 4596 4908
rect 4766 4869 4776 4908
rect 4586 4835 4592 4869
rect 4770 4835 4776 4869
rect 4586 4796 4596 4835
rect 4766 4796 4776 4835
rect 4586 4762 4592 4796
rect 4770 4762 4776 4796
rect 4586 4723 4596 4762
rect 4766 4723 4776 4762
rect 4586 4689 4592 4723
rect 4770 4689 4776 4723
rect 4586 4650 4596 4689
rect 4766 4650 4776 4689
rect 4586 4616 4592 4650
rect 4770 4616 4776 4650
rect 4586 4577 4596 4616
rect 4766 4577 4776 4616
rect 4586 4543 4592 4577
rect 4770 4543 4776 4577
rect 4586 4504 4596 4543
rect 4766 4504 4776 4543
rect 4586 4470 4592 4504
rect 4770 4470 4776 4504
rect 4586 4431 4596 4470
rect 4766 4431 4776 4470
rect 4586 4397 4592 4431
rect 4770 4397 4776 4431
rect 4586 4358 4596 4397
rect 4766 4358 4776 4397
rect 4586 4324 4592 4358
rect 4770 4324 4776 4358
rect 4586 4285 4596 4324
rect 4766 4285 4776 4324
rect 4586 4251 4592 4285
rect 4770 4251 4776 4285
rect 4586 4212 4596 4251
rect 4766 4212 4776 4251
rect 4586 4178 4592 4212
rect 4770 4178 4776 4212
rect 4586 4139 4596 4178
rect 4766 4139 4776 4178
rect 4586 4105 4592 4139
rect 4770 4105 4776 4139
rect 4586 4066 4596 4105
rect 4766 4066 4776 4105
rect 4586 4032 4592 4066
rect 4770 4032 4776 4066
rect 4586 3993 4596 4032
rect 4766 3993 4776 4032
rect 4586 3959 4592 3993
rect 4770 3959 4776 3993
rect 4586 3920 4596 3959
rect 4766 3920 4776 3959
rect 4586 3886 4592 3920
rect 4770 3886 4776 3920
rect 4586 3847 4596 3886
rect 4766 3847 4776 3886
rect 4586 3813 4592 3847
rect 4770 3813 4776 3847
rect 4586 3774 4596 3813
rect 4766 3774 4776 3813
rect 4586 3740 4592 3774
rect 4770 3740 4776 3774
rect 4586 3701 4596 3740
rect 4766 3701 4776 3740
rect 4586 3667 4592 3701
rect 4770 3667 4776 3701
rect 4586 3628 4596 3667
rect 4766 3628 4776 3667
rect 4586 3594 4592 3628
rect 4770 3594 4776 3628
rect 4586 3555 4596 3594
rect 4766 3555 4776 3594
rect 4586 3521 4592 3555
rect 4770 3521 4776 3555
rect 4586 3482 4596 3521
rect 4766 3482 4776 3521
rect 4586 3448 4592 3482
rect 4770 3448 4776 3482
rect 4586 3409 4596 3448
rect 4766 3409 4776 3448
rect 4586 3375 4592 3409
rect 4770 3375 4776 3409
rect 4586 3336 4596 3375
rect 4766 3336 4776 3375
rect 4586 3302 4592 3336
rect 4770 3302 4776 3336
rect 4586 3263 4596 3302
rect 4766 3263 4776 3302
rect 4586 3229 4592 3263
rect 4770 3229 4776 3263
rect 4586 3190 4596 3229
rect 4766 3190 4776 3229
rect 4586 3156 4592 3190
rect 4770 3156 4776 3190
rect 4586 3117 4596 3156
rect 4766 3117 4776 3156
rect 4586 3083 4592 3117
rect 4770 3083 4776 3117
rect 4586 3044 4596 3083
rect 4766 3044 4776 3083
rect 4586 3010 4592 3044
rect 4770 3010 4776 3044
rect 4586 2971 4596 3010
rect 4766 2971 4776 3010
rect 4586 2937 4592 2971
rect 4770 2937 4776 2971
rect 4586 2898 4596 2937
rect 4766 2898 4776 2937
rect 4586 2864 4592 2898
rect 4770 2864 4776 2898
rect 4586 2825 4596 2864
rect 4766 2825 4776 2864
rect 4586 2791 4592 2825
rect 4770 2791 4776 2825
rect 4586 2752 4596 2791
rect 4766 2752 4776 2791
rect 4586 2718 4592 2752
rect 4770 2718 4776 2752
rect 4586 2679 4596 2718
rect 4766 2679 4776 2718
rect 4586 2645 4592 2679
rect 4770 2645 4776 2679
rect 4586 2606 4596 2645
rect 4766 2606 4776 2645
rect 4586 2572 4592 2606
rect 4770 2572 4776 2606
rect 3463 2499 3469 2533
rect 3647 2499 3653 2533
rect 3977 2530 3992 2564
rect 4027 2530 4084 2564
rect 4122 2530 4177 2564
rect 4217 2530 4233 2564
rect 4586 2533 4596 2572
rect 4766 2533 4776 2572
rect 3463 2460 3473 2499
rect 3643 2460 3653 2499
rect 4586 2499 4592 2533
rect 4770 2499 4776 2533
rect 3463 2426 3469 2460
rect 3647 2426 3653 2460
rect 3463 2387 3473 2426
rect 3643 2387 3653 2426
rect 3463 2353 3469 2387
rect 3647 2353 3653 2387
rect 3463 2314 3473 2353
rect 3643 2314 3653 2353
rect 3463 2280 3469 2314
rect 3647 2280 3653 2314
rect 3463 2241 3473 2280
rect 3643 2241 3653 2280
rect 3463 2207 3469 2241
rect 3647 2207 3653 2241
rect 3463 2168 3473 2207
rect 3643 2168 3653 2207
rect 3463 2134 3469 2168
rect 3647 2134 3653 2168
rect 3463 2095 3473 2134
rect 3643 2095 3653 2134
rect 3463 2061 3469 2095
rect 3647 2061 3653 2095
rect 3463 2022 3473 2061
rect 3643 2022 3653 2061
rect 3463 1988 3469 2022
rect 3647 1988 3653 2022
rect 3463 1949 3473 1988
rect 3643 1949 3653 1988
rect 3463 1915 3469 1949
rect 3647 1915 3653 1949
rect 3463 1876 3473 1915
rect 3643 1876 3653 1915
rect 3463 1842 3469 1876
rect 3647 1842 3653 1876
rect 3463 1803 3473 1842
rect 3643 1803 3653 1842
rect 3463 1769 3469 1803
rect 3647 1769 3653 1803
rect 3463 1730 3473 1769
rect 3643 1730 3653 1769
rect -30 403 -24 437
rect 82 403 88 437
rect -30 364 -22 403
rect 80 364 88 403
rect -30 330 -24 364
rect 82 330 88 364
rect -30 291 -22 330
rect 80 291 88 330
rect -30 257 -24 291
rect 82 257 88 291
rect -30 218 -22 257
rect 80 224 88 257
rect 3463 224 3469 1730
rect 80 218 3469 224
rect -30 184 -24 218
rect -30 182 -22 184
rect 3647 224 3653 1730
rect 3810 2480 3844 2492
rect 3810 2406 3844 2434
rect 3810 2331 3844 2361
rect 3810 2256 3844 2288
rect 3810 2181 3844 2216
rect 3810 2106 3844 2144
rect 3810 2034 3844 2072
rect 3810 1962 3844 1997
rect 3810 1890 3844 1922
rect 3810 1818 3844 1847
rect 3810 1746 3844 1772
rect 3810 1674 3844 1697
rect 3810 1602 3844 1622
rect 3810 1530 3844 1547
rect 4369 2480 4403 2492
rect 4369 2406 4403 2434
rect 4369 2331 4403 2361
rect 4369 2256 4403 2288
rect 4369 2181 4403 2216
rect 4369 2106 4403 2144
rect 4369 2034 4403 2072
rect 4369 1962 4403 1997
rect 4369 1890 4403 1922
rect 4369 1818 4403 1847
rect 4369 1746 4403 1772
rect 4369 1674 4403 1697
rect 4369 1602 4403 1622
rect 4369 1530 4403 1547
rect 4586 2460 4596 2499
rect 4766 2460 4776 2499
rect 4586 2426 4592 2460
rect 4770 2426 4776 2460
rect 4586 2387 4596 2426
rect 4766 2387 4776 2426
rect 4586 2353 4592 2387
rect 4770 2353 4776 2387
rect 4586 2314 4596 2353
rect 4766 2314 4776 2353
rect 4586 2280 4592 2314
rect 4770 2280 4776 2314
rect 4586 2241 4596 2280
rect 4766 2241 4776 2280
rect 4586 2207 4592 2241
rect 4770 2207 4776 2241
rect 4586 2168 4596 2207
rect 4766 2168 4776 2207
rect 4586 2134 4592 2168
rect 4770 2134 4776 2168
rect 4586 2095 4596 2134
rect 4766 2095 4776 2134
rect 4586 2061 4592 2095
rect 4770 2061 4776 2095
rect 4586 2022 4596 2061
rect 4766 2022 4776 2061
rect 4586 1988 4592 2022
rect 4770 1988 4776 2022
rect 4586 1949 4596 1988
rect 4766 1949 4776 1988
rect 4586 1915 4592 1949
rect 4770 1915 4776 1949
rect 4586 1876 4596 1915
rect 4766 1876 4776 1915
rect 4586 1842 4592 1876
rect 4770 1842 4776 1876
rect 4586 1803 4596 1842
rect 4766 1803 4776 1842
rect 4586 1769 4592 1803
rect 4770 1769 4776 1803
rect 4586 1730 4596 1769
rect 4766 1730 4776 1769
rect 3972 1346 4013 1380
rect 4047 1346 4088 1380
rect 4122 1346 4163 1380
rect 4197 1346 4238 1380
rect 3938 1308 4272 1346
rect 3972 1274 4013 1308
rect 4047 1274 4088 1308
rect 4122 1274 4163 1308
rect 4197 1274 4238 1308
rect 3945 506 3985 540
rect 4019 506 4059 540
rect 4093 506 4133 540
rect 4167 506 4207 540
rect 4241 506 4281 540
rect 3911 468 4315 506
rect 3945 434 3985 468
rect 4019 434 4059 468
rect 4093 434 4133 468
rect 4167 434 4207 468
rect 4241 434 4281 468
rect 4586 224 4592 1730
rect 3647 218 4592 224
rect 4770 224 4776 1730
rect 4925 5449 10035 5455
rect 4925 5448 5003 5449
rect 5037 5448 5076 5449
rect 5110 5448 5149 5449
rect 5183 5448 5222 5449
rect 5256 5448 5295 5449
rect 6049 5448 6125 5449
rect 6159 5448 6199 5449
rect 6233 5448 6272 5449
rect 6306 5448 6345 5449
rect 6379 5448 6418 5449
rect 6452 5448 6491 5449
rect 6525 5448 6564 5449
rect 6598 5448 6637 5449
rect 6671 5448 6710 5449
rect 6744 5448 6783 5449
rect 6817 5448 6856 5449
rect 6890 5448 6929 5449
rect 6963 5448 7002 5449
rect 7036 5448 7075 5449
rect 7109 5448 7148 5449
rect 7182 5448 7221 5449
rect 7255 5448 7294 5449
rect 7328 5448 7367 5449
rect 7401 5448 7440 5449
rect 7474 5448 7513 5449
rect 7547 5448 7586 5449
rect 7620 5448 7659 5449
rect 7693 5448 7732 5449
rect 7766 5448 7805 5449
rect 7839 5448 7878 5449
rect 7912 5448 7951 5449
rect 7985 5448 8024 5449
rect 8058 5448 8097 5449
rect 8131 5448 8170 5449
rect 8204 5448 8243 5449
rect 8277 5448 8316 5449
rect 8350 5448 8389 5449
rect 8423 5448 8462 5449
rect 8496 5448 8535 5449
rect 8569 5448 8608 5449
rect 8642 5448 8681 5449
rect 8715 5448 8754 5449
rect 8788 5448 8827 5449
rect 8861 5448 8900 5449
rect 8934 5448 8973 5449
rect 9007 5448 9046 5449
rect 9080 5448 9119 5449
rect 9153 5448 9192 5449
rect 9226 5448 9265 5449
rect 9299 5448 9338 5449
rect 9372 5448 9411 5449
rect 9445 5448 9484 5449
rect 9518 5448 9557 5449
rect 9591 5448 9630 5449
rect 9664 5448 9703 5449
rect 9737 5448 9776 5449
rect 9810 5448 9849 5449
rect 9883 5448 9922 5449
rect 4925 5377 5001 5448
rect 4925 3543 4931 5377
rect 9883 5415 9897 5448
rect 9956 5415 10035 5449
rect 9863 5414 9897 5415
rect 9931 5414 10035 5415
rect 9863 5380 10035 5414
rect 9863 5377 9925 5380
rect 10027 5377 10035 5380
rect 5037 5343 5076 5346
rect 5110 5343 5149 5346
rect 5183 5343 5222 5346
rect 5256 5343 5295 5346
rect 6049 5343 6125 5346
rect 6159 5343 6199 5346
rect 6233 5343 6272 5346
rect 6306 5343 6345 5346
rect 6379 5343 6418 5346
rect 6452 5343 6491 5346
rect 6525 5343 6564 5346
rect 6598 5343 6637 5346
rect 6671 5343 6710 5346
rect 6744 5343 6783 5346
rect 6817 5343 6856 5346
rect 6890 5343 6929 5346
rect 6963 5343 7002 5346
rect 7036 5343 7075 5346
rect 7109 5343 7148 5346
rect 7182 5343 7221 5346
rect 7255 5343 7294 5346
rect 7328 5343 7367 5346
rect 7401 5343 7440 5346
rect 7474 5343 7513 5346
rect 7547 5343 7586 5346
rect 7620 5343 7659 5346
rect 7693 5343 7732 5346
rect 7766 5343 7805 5346
rect 7839 5343 7878 5346
rect 7912 5343 7951 5346
rect 7985 5343 8024 5346
rect 8058 5343 8097 5346
rect 8131 5343 8170 5346
rect 8204 5343 8243 5346
rect 8277 5343 8316 5346
rect 8350 5343 8389 5346
rect 8423 5343 8462 5346
rect 8496 5343 8535 5346
rect 8569 5343 8608 5346
rect 8642 5343 8681 5346
rect 8715 5343 8754 5346
rect 8788 5343 8827 5346
rect 8861 5343 8900 5346
rect 8934 5343 8973 5346
rect 9007 5343 9046 5346
rect 9080 5343 9119 5346
rect 9153 5343 9192 5346
rect 9226 5343 9265 5346
rect 9299 5343 9338 5346
rect 9372 5343 9411 5346
rect 9445 5343 9484 5346
rect 9518 5343 9557 5346
rect 9591 5343 9630 5346
rect 9664 5343 9703 5346
rect 9737 5343 9776 5346
rect 9810 5343 9849 5346
rect 9883 5343 9923 5377
rect 10029 5343 10035 5377
rect 5037 5337 9925 5343
rect 5037 3543 5043 5337
rect 4925 3504 4933 3543
rect 5035 3504 5043 3543
rect 4925 3470 4931 3504
rect 5037 3470 5043 3504
rect 4925 3431 4933 3470
rect 5035 3431 5043 3470
rect 4925 3397 4931 3431
rect 5037 3397 5043 3431
rect 4925 3358 4933 3397
rect 5035 3358 5043 3397
rect 4925 3324 4931 3358
rect 5037 3324 5043 3358
rect 4925 3285 4933 3324
rect 5035 3285 5043 3324
rect 4925 3251 4931 3285
rect 5037 3251 5043 3285
rect 4925 3212 4933 3251
rect 5035 3212 5043 3251
rect 9917 5304 9925 5337
rect 10027 5304 10035 5343
rect 9917 5270 9923 5304
rect 10029 5270 10035 5304
rect 9917 5231 9925 5270
rect 10027 5231 10035 5270
rect 9917 5197 9923 5231
rect 10029 5197 10035 5231
rect 9917 5158 9925 5197
rect 10027 5158 10035 5197
rect 9917 5124 9923 5158
rect 10029 5124 10035 5158
rect 9917 5085 9925 5124
rect 10027 5085 10035 5124
rect 9917 5051 9923 5085
rect 10029 5051 10035 5085
rect 9917 5012 9925 5051
rect 10027 5012 10035 5051
rect 9917 4978 9923 5012
rect 10029 4978 10035 5012
rect 9917 4939 9925 4978
rect 10027 4939 10035 4978
rect 9917 4905 9923 4939
rect 10029 4905 10035 4939
rect 9917 4866 9925 4905
rect 10027 4866 10035 4905
rect 9917 4832 9923 4866
rect 10029 4832 10035 4866
rect 9917 4793 9925 4832
rect 10027 4793 10035 4832
rect 9917 4759 9923 4793
rect 10029 4759 10035 4793
rect 9917 4720 9925 4759
rect 10027 4720 10035 4759
rect 9917 4686 9923 4720
rect 10029 4686 10035 4720
rect 9917 4647 9925 4686
rect 10027 4647 10035 4686
rect 9917 4613 9923 4647
rect 10029 4613 10035 4647
rect 9917 4574 9925 4613
rect 10027 4574 10035 4613
rect 9917 4540 9923 4574
rect 10029 4540 10035 4574
rect 9917 4501 9925 4540
rect 10027 4501 10035 4540
rect 9917 4467 9923 4501
rect 10029 4467 10035 4501
rect 9917 4428 9925 4467
rect 10027 4428 10035 4467
rect 9917 4394 9923 4428
rect 10029 4394 10035 4428
rect 9917 4355 9925 4394
rect 10027 4355 10035 4394
rect 9917 4321 9923 4355
rect 10029 4321 10035 4355
rect 9917 4282 9925 4321
rect 10027 4282 10035 4321
rect 9917 4248 9923 4282
rect 10029 4248 10035 4282
rect 9917 4209 9925 4248
rect 10027 4209 10035 4248
rect 9917 4175 9923 4209
rect 10029 4175 10035 4209
rect 9917 4136 9925 4175
rect 10027 4136 10035 4175
rect 9917 4102 9923 4136
rect 10029 4102 10035 4136
rect 9917 4063 9925 4102
rect 10027 4063 10035 4102
rect 9917 4029 9923 4063
rect 10029 4029 10035 4063
rect 9917 3990 9925 4029
rect 10027 3990 10035 4029
rect 9917 3956 9923 3990
rect 10029 3956 10035 3990
rect 9917 3917 9925 3956
rect 10027 3917 10035 3956
rect 9917 3883 9923 3917
rect 10029 3883 10035 3917
rect 9917 3844 9925 3883
rect 10027 3844 10035 3883
rect 9917 3810 9923 3844
rect 10029 3810 10035 3844
rect 9917 3771 9925 3810
rect 10027 3771 10035 3810
rect 9917 3737 9923 3771
rect 10029 3737 10035 3771
rect 9917 3698 9925 3737
rect 10027 3698 10035 3737
rect 9917 3664 9923 3698
rect 10029 3664 10035 3698
rect 9917 3625 9925 3664
rect 10027 3625 10035 3664
rect 9917 3591 9923 3625
rect 10029 3591 10035 3625
rect 9917 3552 9925 3591
rect 10027 3552 10035 3591
rect 9917 3518 9923 3552
rect 10029 3518 10035 3552
rect 9917 3479 9925 3518
rect 10027 3479 10035 3518
rect 9917 3445 9923 3479
rect 10029 3445 10035 3479
rect 9917 3406 9925 3445
rect 10027 3406 10035 3445
rect 9917 3372 9923 3406
rect 10029 3372 10035 3406
rect 9917 3333 9925 3372
rect 10027 3333 10035 3372
rect 9917 3299 9923 3333
rect 10029 3299 10035 3333
rect 9917 3260 9925 3299
rect 10027 3260 10035 3299
rect 9917 3226 9923 3260
rect 10029 3226 10035 3260
rect 4925 3178 4931 3212
rect 5037 3178 5043 3212
rect 5168 3182 5184 3216
rect 5237 3182 5252 3216
rect 5309 3182 5320 3216
rect 5381 3182 5388 3216
rect 5453 3182 5456 3216
rect 5490 3182 5491 3216
rect 5558 3182 5563 3216
rect 5626 3182 5635 3216
rect 5694 3182 5707 3216
rect 5762 3182 5779 3216
rect 5830 3182 5851 3216
rect 5898 3182 5923 3216
rect 5966 3182 5995 3216
rect 6034 3182 6067 3216
rect 6102 3182 6136 3216
rect 6173 3182 6204 3216
rect 6245 3182 6272 3216
rect 6317 3182 6340 3216
rect 6389 3182 6408 3216
rect 6461 3182 6476 3216
rect 6533 3182 6544 3216
rect 6605 3182 6612 3216
rect 6677 3182 6680 3216
rect 6714 3182 6715 3216
rect 6782 3182 6787 3216
rect 6850 3182 6859 3216
rect 6918 3182 6931 3216
rect 6986 3182 7003 3216
rect 7054 3182 7075 3216
rect 7122 3182 7147 3216
rect 7190 3182 7219 3216
rect 7258 3182 7291 3216
rect 7326 3182 7360 3216
rect 7397 3182 7428 3216
rect 7469 3182 7496 3216
rect 7541 3182 7564 3216
rect 7613 3182 7632 3216
rect 7685 3182 7700 3216
rect 7757 3182 7768 3216
rect 7829 3182 7836 3216
rect 7901 3182 7904 3216
rect 7938 3182 7939 3216
rect 8006 3182 8011 3216
rect 8074 3182 8083 3216
rect 8142 3182 8155 3216
rect 8210 3182 8227 3216
rect 8278 3182 8299 3216
rect 8346 3182 8371 3216
rect 8414 3182 8443 3216
rect 8482 3182 8515 3216
rect 8550 3182 8584 3216
rect 8621 3182 8652 3216
rect 8693 3182 8720 3216
rect 8765 3182 8788 3216
rect 8837 3182 8856 3216
rect 8909 3182 8924 3216
rect 8981 3182 8992 3216
rect 9053 3182 9060 3216
rect 9125 3182 9128 3216
rect 9162 3182 9163 3216
rect 9230 3182 9235 3216
rect 9298 3182 9307 3216
rect 9366 3182 9379 3216
rect 9434 3182 9451 3216
rect 9502 3182 9523 3216
rect 9570 3182 9595 3216
rect 9638 3182 9667 3216
rect 9707 3182 9739 3216
rect 9776 3182 9792 3216
rect 9917 3187 9925 3226
rect 10027 3187 10035 3226
rect 4925 3139 4933 3178
rect 5035 3139 5043 3178
rect 4925 3105 4931 3139
rect 5037 3105 5043 3139
rect 4925 3066 4933 3105
rect 5035 3066 5043 3105
rect 4925 3032 4931 3066
rect 5037 3032 5043 3066
rect 4925 2993 4933 3032
rect 5035 3020 5043 3032
rect 9917 3153 9923 3187
rect 10029 3153 10035 3187
rect 9917 3114 9925 3153
rect 10027 3114 10035 3153
rect 9917 3080 9923 3114
rect 10029 3080 10035 3114
rect 9917 3041 9925 3080
rect 10027 3041 10035 3080
rect 9917 3020 9923 3041
rect 5035 3014 9923 3020
rect 5035 2993 5075 3014
rect 5109 3012 5148 3014
rect 5182 3012 5221 3014
rect 5255 3012 5294 3014
rect 5328 3012 5367 3014
rect 5401 3012 5440 3014
rect 5474 3012 5513 3014
rect 5547 3012 5586 3014
rect 5620 3012 5659 3014
rect 5693 3012 5732 3014
rect 5766 3012 5805 3014
rect 5839 3012 5878 3014
rect 5912 3012 5951 3014
rect 5985 3012 6024 3014
rect 6058 3012 6097 3014
rect 6131 3012 6170 3014
rect 6204 3012 6243 3014
rect 6277 3012 6316 3014
rect 6350 3012 6389 3014
rect 6423 3012 6462 3014
rect 6496 3012 6535 3014
rect 6569 3012 6608 3014
rect 6642 3012 6681 3014
rect 6715 3012 6754 3014
rect 6788 3012 6827 3014
rect 9885 3012 9923 3014
rect 4925 2959 4931 2993
rect 5037 2980 5075 2993
rect 5037 2959 5097 2980
rect 4925 2920 4933 2959
rect 5035 2942 5097 2959
rect 5035 2920 5075 2942
rect 4925 2886 4931 2920
rect 5037 2908 5075 2920
rect 10029 3007 10035 3041
rect 10027 2968 10035 3007
rect 9891 2934 9923 2966
rect 9957 2934 9995 2966
rect 10029 2934 10035 2968
rect 9891 2910 10035 2934
rect 5109 2908 5148 2910
rect 5182 2908 5221 2910
rect 5255 2908 5294 2910
rect 5328 2908 5367 2910
rect 5401 2908 5440 2910
rect 5474 2908 5513 2910
rect 5547 2908 5586 2910
rect 5620 2908 5659 2910
rect 5693 2908 5732 2910
rect 5766 2908 5805 2910
rect 5839 2908 5878 2910
rect 5912 2908 5951 2910
rect 5985 2908 6024 2910
rect 6058 2908 6097 2910
rect 6131 2908 6170 2910
rect 6204 2908 6243 2910
rect 6277 2908 6316 2910
rect 6350 2908 6389 2910
rect 6423 2908 6462 2910
rect 6496 2908 6535 2910
rect 6569 2908 6608 2910
rect 6642 2908 6681 2910
rect 6715 2908 6754 2910
rect 6788 2908 6827 2910
rect 9885 2908 10035 2910
rect 5037 2902 10035 2908
rect 5037 2886 5043 2902
rect 4925 2847 4933 2886
rect 5035 2847 5043 2886
rect 4925 2813 4931 2847
rect 5037 2813 5043 2847
rect 4925 2774 4933 2813
rect 5035 2774 5043 2813
rect 4925 2740 4931 2774
rect 5037 2740 5043 2774
rect 9917 2895 10035 2902
rect 9917 2861 9923 2895
rect 9957 2861 9995 2895
rect 10029 2861 10035 2895
rect 9917 2838 10035 2861
rect 9917 2822 9925 2838
rect 10027 2822 10035 2838
rect 9917 2788 9923 2822
rect 10029 2788 10035 2822
rect 9917 2749 9925 2788
rect 10027 2749 10035 2788
rect 4925 2701 4933 2740
rect 5035 2701 5043 2740
rect 5168 2712 5184 2746
rect 5237 2712 5252 2746
rect 5309 2712 5320 2746
rect 5381 2712 5388 2746
rect 5453 2712 5456 2746
rect 5490 2712 5491 2746
rect 5558 2712 5563 2746
rect 5626 2712 5635 2746
rect 5694 2712 5707 2746
rect 5762 2712 5779 2746
rect 5830 2712 5851 2746
rect 5898 2712 5923 2746
rect 5966 2712 5995 2746
rect 6034 2712 6067 2746
rect 6102 2712 6136 2746
rect 6173 2712 6204 2746
rect 6245 2712 6272 2746
rect 6317 2712 6340 2746
rect 6389 2712 6408 2746
rect 6461 2712 6476 2746
rect 6533 2712 6544 2746
rect 6605 2712 6612 2746
rect 6677 2712 6680 2746
rect 6714 2712 6715 2746
rect 6782 2712 6787 2746
rect 6850 2712 6859 2746
rect 6918 2712 6931 2746
rect 6986 2712 7003 2746
rect 7054 2712 7075 2746
rect 7122 2712 7147 2746
rect 7190 2712 7219 2746
rect 7258 2712 7291 2746
rect 7326 2712 7360 2746
rect 7397 2712 7428 2746
rect 7469 2712 7496 2746
rect 7541 2712 7564 2746
rect 7613 2712 7632 2746
rect 7685 2712 7700 2746
rect 7757 2712 7768 2746
rect 7829 2712 7836 2746
rect 7901 2712 7904 2746
rect 7938 2712 7939 2746
rect 8006 2712 8011 2746
rect 8074 2712 8083 2746
rect 8142 2712 8155 2746
rect 8210 2712 8227 2746
rect 8278 2712 8299 2746
rect 8346 2712 8371 2746
rect 8414 2712 8443 2746
rect 8482 2712 8515 2746
rect 8550 2712 8584 2746
rect 8621 2712 8652 2746
rect 8693 2712 8720 2746
rect 8765 2712 8788 2746
rect 8837 2712 8856 2746
rect 8909 2712 8924 2746
rect 8981 2712 8992 2746
rect 9053 2712 9060 2746
rect 9125 2712 9128 2746
rect 9162 2712 9163 2746
rect 9230 2712 9235 2746
rect 9298 2712 9307 2746
rect 9366 2712 9379 2746
rect 9434 2712 9451 2746
rect 9502 2712 9523 2746
rect 9570 2712 9595 2746
rect 9638 2712 9667 2746
rect 9707 2712 9739 2746
rect 9776 2712 9792 2746
rect 9917 2715 9923 2749
rect 10029 2715 10035 2749
rect 4925 2667 4931 2701
rect 5037 2667 5043 2701
rect 4925 2628 4933 2667
rect 5035 2628 5043 2667
rect 4925 2594 4931 2628
rect 5037 2594 5043 2628
rect 4925 2555 4933 2594
rect 5035 2555 5043 2594
rect 4925 2521 4931 2555
rect 5037 2521 5043 2555
rect 4925 2482 4933 2521
rect 5035 2482 5043 2521
rect 4925 2448 4931 2482
rect 5037 2448 5043 2482
rect 4925 2409 4933 2448
rect 5035 2409 5043 2448
rect 4925 2375 4931 2409
rect 5037 2375 5043 2409
rect 4925 2336 4933 2375
rect 5035 2336 5043 2375
rect 4925 2302 4931 2336
rect 5037 2302 5043 2336
rect 4925 2263 4933 2302
rect 5035 2263 5043 2302
rect 4925 2229 4931 2263
rect 5037 2229 5043 2263
rect 4925 2190 4933 2229
rect 5035 2190 5043 2229
rect 4925 2156 4931 2190
rect 5037 2156 5043 2190
rect 4925 2117 4933 2156
rect 5035 2117 5043 2156
rect 4925 2083 4931 2117
rect 5037 2083 5043 2117
rect 4925 2044 4933 2083
rect 5035 2044 5043 2083
rect 4925 2010 4931 2044
rect 5037 2010 5043 2044
rect 4925 1971 4933 2010
rect 5035 1971 5043 2010
rect 4925 1937 4931 1971
rect 5037 1937 5043 1971
rect 4925 1898 4933 1937
rect 5035 1898 5043 1937
rect 4925 1864 4931 1898
rect 5037 1864 5043 1898
rect 4925 1825 4933 1864
rect 5035 1825 5043 1864
rect 4925 1791 4931 1825
rect 5037 1791 5043 1825
rect 4925 1752 4933 1791
rect 5035 1752 5043 1791
rect 4925 1718 4931 1752
rect 5037 1718 5043 1752
rect 4925 1679 4933 1718
rect 5035 1679 5043 1718
rect 4925 1645 4931 1679
rect 5037 1645 5043 1679
rect 4925 1606 4933 1645
rect 5035 1606 5043 1645
rect 4925 1572 4931 1606
rect 5037 1572 5043 1606
rect 4925 1533 4933 1572
rect 5035 1533 5043 1572
rect 4925 1499 4931 1533
rect 5037 1499 5043 1533
rect 4925 1460 4933 1499
rect 5035 1460 5043 1499
rect 4925 1426 4931 1460
rect 5037 1426 5043 1460
rect 4925 1387 4933 1426
rect 5035 1387 5043 1426
rect 4925 1353 4931 1387
rect 5037 1353 5043 1387
rect 4925 1314 4933 1353
rect 5035 1314 5043 1353
rect 4925 1280 4931 1314
rect 5037 1280 5043 1314
rect 4925 1241 4933 1280
rect 5035 1241 5043 1280
rect 4925 1207 4931 1241
rect 5037 1207 5043 1241
rect 4925 1168 4933 1207
rect 5035 1168 5043 1207
rect 4925 1134 4931 1168
rect 5037 1134 5043 1168
rect 4925 1095 4933 1134
rect 5035 1095 5043 1134
rect 4925 1061 4931 1095
rect 5037 1061 5043 1095
rect 4925 1022 4933 1061
rect 5035 1022 5043 1061
rect 4925 988 4931 1022
rect 5037 988 5043 1022
rect 4925 949 4933 988
rect 5035 949 5043 988
rect 4925 915 4931 949
rect 5037 915 5043 949
rect 4925 876 4933 915
rect 5035 876 5043 915
rect 4925 842 4931 876
rect 5037 842 5043 876
rect 4925 803 4933 842
rect 5035 803 5043 842
rect 4925 769 4931 803
rect 5037 769 5043 803
rect 4925 730 4933 769
rect 5035 730 5043 769
rect 4925 696 4931 730
rect 5037 696 5043 730
rect 4925 657 4933 696
rect 5035 657 5043 696
rect 4925 623 4931 657
rect 5037 623 5043 657
rect 4925 584 4933 623
rect 5035 590 5043 623
rect 9917 2676 9925 2715
rect 10027 2676 10035 2715
rect 9917 2642 9923 2676
rect 10029 2642 10035 2676
rect 9917 2603 9925 2642
rect 10027 2603 10035 2642
rect 9917 2569 9923 2603
rect 10029 2569 10035 2603
rect 9917 2530 9925 2569
rect 10027 2530 10035 2569
rect 9917 2496 9923 2530
rect 10029 2496 10035 2530
rect 9917 2457 9925 2496
rect 10027 2457 10035 2496
rect 9917 2423 9923 2457
rect 10029 2423 10035 2457
rect 9917 2384 9925 2423
rect 10027 2384 10035 2423
rect 9917 590 9923 2384
rect 5035 584 9923 590
rect 4925 550 4931 584
rect 4925 548 4933 550
rect 8205 582 8244 584
rect 8278 582 8317 584
rect 8351 582 8390 584
rect 8424 582 8463 584
rect 8497 582 8536 584
rect 8570 582 8609 584
rect 8643 582 8682 584
rect 8716 582 8755 584
rect 8789 582 8828 584
rect 8862 582 8901 584
rect 8935 582 8974 584
rect 9008 582 9047 584
rect 9081 582 9120 584
rect 9154 582 9193 584
rect 9227 582 9266 584
rect 9300 582 9339 584
rect 9373 582 9412 584
rect 9446 582 9485 584
rect 9519 582 9558 584
rect 9592 582 9631 584
rect 9665 582 9704 584
rect 9738 582 9777 584
rect 9811 582 9850 584
rect 9884 582 9923 584
rect 4925 478 5003 548
rect 10029 550 10035 2384
rect 9959 480 10035 550
rect 8205 478 8244 480
rect 8278 478 8317 480
rect 8351 478 8390 480
rect 8424 478 8463 480
rect 8497 478 8536 480
rect 8570 478 8609 480
rect 8643 478 8682 480
rect 8716 478 8755 480
rect 8789 478 8828 480
rect 8862 478 8901 480
rect 8935 478 8974 480
rect 9008 478 9047 480
rect 9081 478 9120 480
rect 9154 478 9193 480
rect 9227 478 9266 480
rect 9300 478 9339 480
rect 9373 478 9412 480
rect 9446 478 9485 480
rect 9519 478 9558 480
rect 9592 478 9631 480
rect 9665 478 9704 480
rect 9738 478 9777 480
rect 9811 478 9850 480
rect 9884 478 9923 480
rect 9957 478 10035 480
rect 4925 472 10035 478
rect 10271 5452 10279 5491
rect 10381 5452 10389 5491
rect 10271 5418 10277 5452
rect 10383 5418 10389 5452
rect 10271 5379 10279 5418
rect 10381 5379 10389 5418
rect 10271 5345 10277 5379
rect 10383 5345 10389 5379
rect 10271 5306 10279 5345
rect 10381 5306 10389 5345
rect 10271 5272 10277 5306
rect 10383 5272 10389 5306
rect 10271 5233 10279 5272
rect 10381 5233 10389 5272
rect 10271 5199 10277 5233
rect 10383 5199 10389 5233
rect 10271 5160 10279 5199
rect 10381 5160 10389 5199
rect 10271 5126 10277 5160
rect 10383 5126 10389 5160
rect 10271 5087 10279 5126
rect 10381 5087 10389 5126
rect 10271 5053 10277 5087
rect 10383 5053 10389 5087
rect 10271 5014 10279 5053
rect 10381 5014 10389 5053
rect 10271 4980 10277 5014
rect 10383 4980 10389 5014
rect 10271 4941 10279 4980
rect 10381 4941 10389 4980
rect 10271 4907 10277 4941
rect 10383 4907 10389 4941
rect 10271 4868 10279 4907
rect 10381 4868 10389 4907
rect 10271 4834 10277 4868
rect 10383 4834 10389 4868
rect 10271 4795 10279 4834
rect 10381 4795 10389 4834
rect 10271 4761 10277 4795
rect 10383 4761 10389 4795
rect 10271 4722 10279 4761
rect 10381 4722 10389 4761
rect 10271 4688 10277 4722
rect 10383 4688 10389 4722
rect 10271 4649 10279 4688
rect 10381 4649 10389 4688
rect 10271 4615 10277 4649
rect 10383 4615 10389 4649
rect 10271 4576 10279 4615
rect 10381 4576 10389 4615
rect 10271 4542 10277 4576
rect 10383 4542 10389 4576
rect 10271 4503 10279 4542
rect 10381 4503 10389 4542
rect 10271 4469 10277 4503
rect 10383 4469 10389 4503
rect 10271 4430 10279 4469
rect 10381 4430 10389 4469
rect 10271 4396 10277 4430
rect 10383 4396 10389 4430
rect 10271 4357 10279 4396
rect 10381 4357 10389 4396
rect 10271 4323 10277 4357
rect 10383 4323 10389 4357
rect 10271 4284 10279 4323
rect 10381 4284 10389 4323
rect 10271 4250 10277 4284
rect 10383 4250 10389 4284
rect 10271 4211 10279 4250
rect 10381 4211 10389 4250
rect 10271 4177 10277 4211
rect 10383 4177 10389 4211
rect 10271 4138 10279 4177
rect 10381 4138 10389 4177
rect 10271 4104 10277 4138
rect 10383 4104 10389 4138
rect 10271 4065 10279 4104
rect 10381 4065 10389 4104
rect 10271 4031 10277 4065
rect 10383 4031 10389 4065
rect 10271 3992 10279 4031
rect 10381 3992 10389 4031
rect 10271 3958 10277 3992
rect 10383 3958 10389 3992
rect 10271 3919 10279 3958
rect 10381 3919 10389 3958
rect 10271 3885 10277 3919
rect 10383 3885 10389 3919
rect 10271 3846 10279 3885
rect 10381 3846 10389 3885
rect 10271 3812 10277 3846
rect 10383 3812 10389 3846
rect 10271 3773 10279 3812
rect 10381 3773 10389 3812
rect 10271 3739 10277 3773
rect 10383 3739 10389 3773
rect 10271 3700 10279 3739
rect 10381 3700 10389 3739
rect 10271 3666 10277 3700
rect 10383 3666 10389 3700
rect 10271 3627 10279 3666
rect 10381 3627 10389 3666
rect 10271 3593 10277 3627
rect 10383 3593 10389 3627
rect 10271 3554 10279 3593
rect 10381 3554 10389 3593
rect 10271 3520 10277 3554
rect 10383 3520 10389 3554
rect 10271 3481 10279 3520
rect 10381 3481 10389 3520
rect 10271 3447 10277 3481
rect 10383 3447 10389 3481
rect 10271 3408 10279 3447
rect 10381 3408 10389 3447
rect 10271 3374 10277 3408
rect 10383 3374 10389 3408
rect 10271 3335 10279 3374
rect 10381 3335 10389 3374
rect 10271 3301 10277 3335
rect 10383 3301 10389 3335
rect 10271 3262 10279 3301
rect 10381 3262 10389 3301
rect 10271 3228 10277 3262
rect 10383 3228 10389 3262
rect 10271 3189 10279 3228
rect 10381 3189 10389 3228
rect 10271 3155 10277 3189
rect 10383 3155 10389 3189
rect 10271 3116 10279 3155
rect 10381 3116 10389 3155
rect 10271 3082 10277 3116
rect 10383 3082 10389 3116
rect 10271 3043 10279 3082
rect 10381 3043 10389 3082
rect 10271 3009 10277 3043
rect 10383 3009 10389 3043
rect 10271 2970 10279 3009
rect 10381 2970 10389 3009
rect 10271 2936 10277 2970
rect 10383 2936 10389 2970
rect 10271 2897 10279 2936
rect 10381 2897 10389 2936
rect 10271 2863 10277 2897
rect 10383 2863 10389 2897
rect 10271 2824 10279 2863
rect 10381 2824 10389 2863
rect 10271 2790 10277 2824
rect 10383 2790 10389 2824
rect 10271 2751 10279 2790
rect 10381 2751 10389 2790
rect 10271 2717 10277 2751
rect 10383 2717 10389 2751
rect 10271 2678 10279 2717
rect 10381 2678 10389 2717
rect 10271 2644 10277 2678
rect 10383 2644 10389 2678
rect 10271 2605 10279 2644
rect 10381 2605 10389 2644
rect 10271 2571 10277 2605
rect 10383 2571 10389 2605
rect 10271 2532 10279 2571
rect 10381 2532 10389 2571
rect 10271 2498 10277 2532
rect 10383 2498 10389 2532
rect 10271 2459 10279 2498
rect 10381 2459 10389 2498
rect 10271 2425 10277 2459
rect 10383 2425 10389 2459
rect 10271 2386 10279 2425
rect 10381 2386 10389 2425
rect 10271 2352 10277 2386
rect 10383 2352 10389 2386
rect 10271 2313 10279 2352
rect 10381 2313 10389 2352
rect 10271 2279 10277 2313
rect 10383 2279 10389 2313
rect 10271 2240 10279 2279
rect 10381 2240 10389 2279
rect 10271 2206 10277 2240
rect 10383 2206 10389 2240
rect 10271 2167 10279 2206
rect 10381 2167 10389 2206
rect 10271 2133 10277 2167
rect 10383 2133 10389 2167
rect 10271 2094 10279 2133
rect 10381 2094 10389 2133
rect 10271 2060 10277 2094
rect 10383 2060 10389 2094
rect 10271 2021 10279 2060
rect 10381 2021 10389 2060
rect 10271 1987 10277 2021
rect 10383 1987 10389 2021
rect 10271 1948 10279 1987
rect 10381 1948 10389 1987
rect 10271 1914 10277 1948
rect 10383 1914 10389 1948
rect 10271 1875 10279 1914
rect 10381 1875 10389 1914
rect 10271 1841 10277 1875
rect 10383 1841 10389 1875
rect 10271 1802 10279 1841
rect 10381 1802 10389 1841
rect 10271 224 10277 1802
rect 4770 218 10277 224
rect 9946 216 9985 218
rect 10019 216 10058 218
rect 10092 216 10131 218
rect 10165 216 10204 218
rect 10238 216 10277 218
rect -30 112 48 182
rect 10383 184 10389 1802
rect 10313 114 10389 184
rect 9946 112 9985 114
rect 10019 112 10058 114
rect 10092 112 10131 114
rect 10165 112 10204 114
rect 10238 112 10277 114
rect 10311 112 10389 114
rect -30 106 10389 112
<< viali >>
rect 48 5814 82 5816
rect 121 5814 155 5816
rect 194 5814 228 5816
rect 267 5814 301 5816
rect 340 5814 374 5816
rect 413 5814 447 5816
rect 486 5814 520 5816
rect 559 5814 593 5816
rect 632 5814 666 5816
rect 705 5814 739 5816
rect 778 5814 812 5816
rect 851 5814 885 5816
rect 924 5814 958 5816
rect 997 5814 1031 5816
rect 1070 5814 1104 5816
rect 1143 5814 1177 5816
rect 1216 5814 9458 5816
rect 9534 5814 9568 5816
rect 9609 5814 9643 5816
rect 9683 5814 9717 5816
rect 9757 5814 9791 5816
rect 9831 5814 9865 5816
rect 9905 5814 9939 5816
rect 9979 5814 10013 5816
rect 10053 5814 10087 5816
rect 10127 5814 10161 5816
rect 10201 5814 10235 5816
rect 10275 5814 10309 5816
rect 48 5782 82 5814
rect 121 5782 155 5814
rect 194 5782 228 5814
rect 267 5782 301 5814
rect 340 5782 374 5814
rect 413 5782 447 5814
rect 486 5782 520 5814
rect 559 5782 593 5814
rect 632 5782 666 5814
rect 705 5782 739 5814
rect 778 5782 812 5814
rect 851 5782 885 5814
rect 924 5782 958 5814
rect 997 5782 1031 5814
rect 1070 5782 1104 5814
rect 1143 5782 1177 5814
rect -24 5724 46 5744
rect -24 5690 -22 5724
rect -22 5690 12 5724
rect 12 5712 46 5724
rect 46 5712 82 5744
rect 121 5712 155 5744
rect 194 5712 228 5744
rect 267 5712 301 5744
rect 340 5712 374 5744
rect 413 5712 447 5744
rect 486 5712 520 5744
rect 559 5712 593 5744
rect 632 5712 666 5744
rect 705 5712 739 5744
rect 778 5712 812 5744
rect 851 5712 885 5744
rect 924 5712 958 5744
rect 997 5712 1031 5744
rect 1070 5712 1104 5744
rect 1143 5712 1177 5744
rect 1216 5712 9458 5814
rect 9534 5782 9568 5814
rect 9609 5782 9643 5814
rect 9683 5782 9717 5814
rect 9757 5782 9791 5814
rect 9831 5782 9865 5814
rect 9905 5782 9939 5814
rect 9979 5782 10013 5814
rect 10053 5782 10087 5814
rect 10127 5782 10161 5814
rect 10201 5782 10212 5814
rect 10212 5782 10235 5814
rect 10275 5782 10280 5814
rect 10280 5782 10309 5814
rect 9534 5712 9568 5744
rect 9609 5712 9643 5744
rect 9683 5712 9717 5744
rect 9757 5712 9791 5744
rect 9831 5712 9865 5744
rect 9905 5712 9939 5744
rect 9979 5712 10013 5744
rect 10053 5712 10087 5744
rect 10127 5712 10161 5744
rect 10201 5712 10212 5744
rect 10212 5712 10235 5744
rect 12 5690 82 5712
rect 121 5710 155 5712
rect 194 5710 228 5712
rect 267 5710 301 5712
rect 340 5710 374 5712
rect 413 5710 447 5712
rect 486 5710 520 5712
rect 559 5710 593 5712
rect 632 5710 666 5712
rect 705 5710 739 5712
rect 778 5710 812 5712
rect 851 5710 885 5712
rect 924 5710 958 5712
rect 997 5710 1031 5712
rect 1070 5710 1104 5712
rect 1143 5710 1177 5712
rect 1216 5710 9458 5712
rect 9534 5710 9568 5712
rect 9609 5710 9643 5712
rect 9683 5710 9717 5712
rect 9757 5710 9791 5712
rect 9831 5710 9865 5712
rect 9905 5710 9939 5712
rect 9979 5710 10013 5712
rect 10053 5710 10087 5712
rect 10127 5710 10161 5712
rect 10201 5710 10235 5712
rect 10277 5710 10279 5744
rect 10279 5710 10311 5744
rect 10349 5710 10381 5744
rect 10381 5710 10383 5744
rect -24 5656 82 5690
rect -24 4126 -22 5656
rect -22 4126 80 5656
rect 80 4126 82 5656
rect 3469 5656 3647 5710
rect 3469 5638 3473 5656
rect 3473 5638 3643 5656
rect 3643 5638 3647 5656
rect 3469 5565 3473 5599
rect 3473 5565 3503 5599
rect 3541 5565 3575 5599
rect 3613 5565 3643 5599
rect 3643 5565 3647 5599
rect 3469 5492 3473 5526
rect 3473 5492 3503 5526
rect 3541 5492 3575 5526
rect 3613 5492 3643 5526
rect 3643 5492 3647 5526
rect -24 4053 -22 4087
rect -22 4053 10 4087
rect 48 4053 80 4087
rect 80 4053 82 4087
rect -24 3980 -22 4014
rect -22 3980 10 4014
rect 48 3980 80 4014
rect 80 3980 82 4014
rect -24 3907 -22 3941
rect -22 3907 10 3941
rect 48 3907 80 3941
rect 80 3907 82 3941
rect -24 3834 -22 3868
rect -22 3834 10 3868
rect 48 3834 80 3868
rect 80 3834 82 3868
rect -24 3761 -22 3795
rect -22 3761 10 3795
rect 48 3761 80 3795
rect 80 3761 82 3795
rect -24 3688 -22 3722
rect -22 3688 10 3722
rect 48 3688 80 3722
rect 80 3688 82 3722
rect -24 3615 -22 3649
rect -22 3615 10 3649
rect 48 3615 80 3649
rect 80 3615 82 3649
rect -24 3542 -22 3576
rect -22 3542 10 3576
rect 48 3542 80 3576
rect 80 3542 82 3576
rect -24 3469 -22 3503
rect -22 3469 10 3503
rect 48 3469 80 3503
rect 80 3469 82 3503
rect -24 3396 -22 3430
rect -22 3396 10 3430
rect 48 3396 80 3430
rect 80 3396 82 3430
rect -24 3323 -22 3357
rect -22 3323 10 3357
rect 48 3323 80 3357
rect 80 3323 82 3357
rect -24 3250 -22 3284
rect -22 3250 10 3284
rect 48 3250 80 3284
rect 80 3250 82 3284
rect -24 3177 -22 3211
rect -22 3177 10 3211
rect 48 3177 80 3211
rect 80 3177 82 3211
rect -24 3104 -22 3138
rect -22 3104 10 3138
rect 48 3104 80 3138
rect 80 3104 82 3138
rect -24 3031 -22 3065
rect -22 3031 10 3065
rect 48 3031 80 3065
rect 80 3031 82 3065
rect -24 2958 -22 2992
rect -22 2958 10 2992
rect 48 2958 80 2992
rect 80 2958 82 2992
rect -24 2885 -22 2919
rect -22 2885 10 2919
rect 48 2885 80 2919
rect 80 2885 82 2919
rect -24 2812 -22 2846
rect -22 2812 10 2846
rect 48 2812 80 2846
rect 80 2812 82 2846
rect -24 2739 -22 2773
rect -22 2739 10 2773
rect 48 2739 80 2773
rect 80 2739 82 2773
rect -24 2666 -22 2700
rect -22 2666 10 2700
rect 48 2666 80 2700
rect 80 2666 82 2700
rect -24 2593 -22 2627
rect -22 2593 10 2627
rect 48 2593 80 2627
rect 80 2593 82 2627
rect -24 2520 -22 2554
rect -22 2520 10 2554
rect 48 2520 80 2554
rect 80 2520 82 2554
rect -24 2447 -22 2481
rect -22 2447 10 2481
rect 48 2447 80 2481
rect 80 2447 82 2481
rect -24 2374 -22 2408
rect -22 2374 10 2408
rect 48 2374 80 2408
rect 80 2374 82 2408
rect -24 2301 -22 2335
rect -22 2301 10 2335
rect 48 2301 80 2335
rect 80 2301 82 2335
rect -24 2228 -22 2262
rect -22 2228 10 2262
rect 48 2228 80 2262
rect 80 2228 82 2262
rect -24 2155 -22 2189
rect -22 2155 10 2189
rect 48 2155 80 2189
rect 80 2155 82 2189
rect -24 2082 -22 2116
rect -22 2082 10 2116
rect 48 2082 80 2116
rect 80 2082 82 2116
rect -24 2009 -22 2043
rect -22 2009 10 2043
rect 48 2009 80 2043
rect 80 2009 82 2043
rect -24 1936 -22 1970
rect -22 1936 10 1970
rect 48 1936 80 1970
rect 80 1936 82 1970
rect -24 1863 -22 1897
rect -22 1863 10 1897
rect 48 1863 80 1897
rect 80 1863 82 1897
rect -24 1790 -22 1824
rect -22 1790 10 1824
rect 48 1790 80 1824
rect 80 1790 82 1824
rect -24 1717 -22 1751
rect -22 1717 10 1751
rect 48 1717 80 1751
rect 80 1717 82 1751
rect -24 1644 -22 1678
rect -22 1644 10 1678
rect 48 1644 80 1678
rect 80 1644 82 1678
rect -24 1571 -22 1605
rect -22 1571 10 1605
rect 48 1571 80 1605
rect 80 1571 82 1605
rect -24 1498 -22 1532
rect -22 1498 10 1532
rect 48 1498 80 1532
rect 80 1498 82 1532
rect -24 1425 -22 1459
rect -22 1425 10 1459
rect 48 1425 80 1459
rect 80 1425 82 1459
rect -24 1352 -22 1386
rect -22 1352 10 1386
rect 48 1352 80 1386
rect 80 1352 82 1386
rect -24 1279 -22 1313
rect -22 1279 10 1313
rect 48 1279 80 1313
rect 80 1279 82 1313
rect -24 1206 -22 1240
rect -22 1206 10 1240
rect 48 1206 80 1240
rect 80 1206 82 1240
rect -24 1133 -22 1167
rect -22 1133 10 1167
rect 48 1133 80 1167
rect 80 1133 82 1167
rect -24 1060 -22 1094
rect -22 1060 10 1094
rect 48 1060 80 1094
rect 80 1060 82 1094
rect -24 987 -22 1021
rect -22 987 10 1021
rect 48 987 80 1021
rect 80 987 82 1021
rect -24 914 -22 948
rect -22 914 10 948
rect 48 914 80 948
rect 80 914 82 948
rect -24 841 -22 875
rect -22 841 10 875
rect 48 841 80 875
rect 80 841 82 875
rect -24 768 -22 802
rect -22 768 10 802
rect 48 768 80 802
rect 80 768 82 802
rect -24 695 -22 729
rect -22 695 10 729
rect 48 695 80 729
rect 80 695 82 729
rect -24 622 -22 656
rect -22 622 10 656
rect 48 622 80 656
rect 80 622 82 656
rect -24 549 -22 583
rect -22 549 10 583
rect 48 549 80 583
rect 80 549 82 583
rect -24 476 -22 510
rect -22 476 10 510
rect 48 476 80 510
rect 80 476 82 510
rect 408 5440 430 5474
rect 430 5440 442 5474
rect 490 5440 498 5474
rect 498 5440 524 5474
rect 572 5440 600 5474
rect 600 5440 606 5474
rect 654 5440 668 5474
rect 668 5440 688 5474
rect 736 5440 770 5474
rect 819 5440 838 5474
rect 838 5440 853 5474
rect 929 5440 940 5474
rect 940 5440 963 5474
rect 1001 5440 1008 5474
rect 1008 5440 1035 5474
rect 1073 5440 1076 5474
rect 1076 5440 1107 5474
rect 1145 5440 1178 5474
rect 1178 5440 1179 5474
rect 1217 5440 1246 5474
rect 1246 5440 1251 5474
rect 1289 5440 1314 5474
rect 1314 5440 1323 5474
rect 1361 5440 1382 5474
rect 1382 5440 1395 5474
rect 1433 5440 1450 5474
rect 1450 5440 1467 5474
rect 1505 5440 1518 5474
rect 1518 5440 1539 5474
rect 1577 5440 1586 5474
rect 1586 5440 1611 5474
rect 1649 5440 1654 5474
rect 1654 5440 1683 5474
rect 1721 5440 1722 5474
rect 1722 5440 1755 5474
rect 1794 5440 1824 5474
rect 1824 5440 1828 5474
rect 1867 5440 1892 5474
rect 1892 5440 1901 5474
rect 1940 5440 1960 5474
rect 1960 5440 1974 5474
rect 2013 5440 2028 5474
rect 2028 5440 2047 5474
rect 2086 5440 2096 5474
rect 2096 5440 2120 5474
rect 2159 5440 2164 5474
rect 2164 5440 2193 5474
rect 2232 5440 2266 5474
rect 2305 5440 2334 5474
rect 2334 5440 2339 5474
rect 2378 5440 2402 5474
rect 2402 5440 2412 5474
rect 2451 5440 2470 5474
rect 2470 5440 2485 5474
rect 2524 5440 2538 5474
rect 2538 5440 2558 5474
rect 2597 5440 2606 5474
rect 2606 5440 2631 5474
rect 2670 5440 2674 5474
rect 2674 5440 2704 5474
rect 2743 5440 2776 5474
rect 2776 5440 2777 5474
rect 2816 5440 2844 5474
rect 2844 5440 2850 5474
rect 2889 5440 2912 5474
rect 2912 5440 2923 5474
rect 2962 5440 2980 5474
rect 2980 5440 2996 5474
rect 3035 5440 3048 5474
rect 3048 5440 3069 5474
rect 3108 5440 3116 5474
rect 3116 5440 3142 5474
rect 3181 5440 3184 5474
rect 3184 5440 3215 5474
rect 326 5372 360 5402
rect 326 5368 360 5372
rect 326 5304 360 5329
rect 326 5295 360 5304
rect 3253 5384 3287 5402
rect 3253 5368 3286 5384
rect 3286 5368 3287 5384
rect 3253 5316 3287 5330
rect 3253 5296 3286 5316
rect 3286 5296 3287 5316
rect 326 5236 360 5256
rect 326 5222 360 5236
rect 326 5168 360 5183
rect 326 5149 360 5168
rect 326 5100 360 5110
rect 326 5076 360 5100
rect 326 5032 360 5037
rect 326 5003 360 5032
rect 326 4930 360 4964
rect 326 4862 360 4891
rect 326 4857 360 4862
rect 326 4794 360 4818
rect 326 4784 360 4794
rect 326 4726 360 4745
rect 326 4711 360 4726
rect 326 4658 360 4672
rect 326 4638 360 4658
rect 326 4590 360 4599
rect 326 4565 360 4590
rect 326 4522 360 4526
rect 326 4492 360 4522
rect 326 4420 360 4453
rect 326 4419 360 4420
rect 326 4352 360 4380
rect 326 4346 360 4352
rect 326 4284 360 4307
rect 326 4273 360 4284
rect 326 4216 360 4234
rect 326 4200 360 4216
rect 326 4148 360 4161
rect 326 4127 360 4148
rect 326 4080 360 4088
rect 326 4054 360 4080
rect 326 4012 360 4016
rect 326 3982 360 4012
rect 326 3910 360 3944
rect 326 3842 360 3872
rect 326 3838 360 3842
rect 326 3774 360 3800
rect 326 3766 360 3774
rect 326 3706 360 3728
rect 326 3694 360 3706
rect 326 3638 360 3656
rect 326 3622 360 3638
rect 326 3570 360 3584
rect 326 3550 360 3570
rect 326 3502 360 3512
rect 326 3478 360 3502
rect 326 3434 360 3440
rect 326 3406 360 3434
rect 326 3366 360 3368
rect 326 3334 360 3366
rect 326 3264 360 3296
rect 326 3262 360 3264
rect 326 3196 360 3224
rect 326 3190 360 3196
rect 326 3128 360 3152
rect 326 3118 360 3128
rect 326 3060 360 3080
rect 326 3046 360 3060
rect 326 2992 360 3008
rect 326 2974 360 2992
rect 326 2924 360 2936
rect 326 2902 360 2924
rect 326 2856 360 2864
rect 326 2830 360 2856
rect 326 2788 360 2792
rect 326 2758 360 2788
rect 326 2686 360 2720
rect 326 2618 360 2648
rect 326 2614 360 2618
rect 326 2550 360 2576
rect 326 2542 360 2550
rect 326 2482 360 2504
rect 326 2470 360 2482
rect 326 2414 360 2432
rect 326 2398 360 2414
rect 326 2346 360 2360
rect 326 2326 360 2346
rect 326 2278 360 2288
rect 326 2254 360 2278
rect 326 2210 360 2216
rect 326 2182 360 2210
rect 326 2142 360 2144
rect 326 2110 360 2142
rect 326 2040 360 2072
rect 326 2038 360 2040
rect 326 1972 360 2000
rect 326 1966 360 1972
rect 326 1904 360 1928
rect 326 1894 360 1904
rect 326 1836 360 1856
rect 326 1822 360 1836
rect 326 1768 360 1784
rect 326 1750 360 1768
rect 326 1700 360 1712
rect 326 1678 360 1700
rect 326 1632 360 1640
rect 326 1606 360 1632
rect 326 1564 360 1568
rect 326 1534 360 1564
rect 326 1462 360 1496
rect 326 1394 360 1424
rect 326 1390 360 1394
rect 326 1326 360 1352
rect 326 1318 360 1326
rect 326 1258 360 1280
rect 326 1246 360 1258
rect 326 1190 360 1208
rect 326 1174 360 1190
rect 326 1122 360 1136
rect 326 1102 360 1122
rect 326 1054 360 1064
rect 326 1030 360 1054
rect 326 986 360 992
rect 326 958 360 986
rect 326 918 360 920
rect 326 886 360 918
rect 326 816 360 848
rect 326 814 360 816
rect 326 748 360 776
rect 326 742 360 748
rect 326 680 360 704
rect 326 670 360 680
rect 600 5265 634 5274
rect 675 5265 709 5274
rect 750 5265 784 5274
rect 825 5265 859 5274
rect 900 5265 934 5274
rect 976 5265 1010 5274
rect 1052 5265 1086 5274
rect 1128 5265 1162 5274
rect 1204 5265 1238 5274
rect 1280 5265 1314 5274
rect 1356 5265 1390 5274
rect 1432 5265 1466 5274
rect 1508 5265 1542 5274
rect 1584 5265 1618 5274
rect 1660 5265 1694 5274
rect 1736 5265 1770 5274
rect 1846 5265 1880 5274
rect 1921 5265 1955 5274
rect 1996 5265 2030 5274
rect 2071 5265 2105 5274
rect 2146 5265 2180 5274
rect 2221 5265 2255 5274
rect 2297 5265 2331 5274
rect 2373 5265 2407 5274
rect 2449 5265 2483 5274
rect 2525 5265 2559 5274
rect 2601 5265 2635 5274
rect 2677 5265 2711 5274
rect 2753 5265 2787 5274
rect 2829 5265 2863 5274
rect 2905 5265 2939 5274
rect 2981 5265 3015 5274
rect 600 5240 603 5265
rect 603 5240 634 5265
rect 675 5240 709 5265
rect 750 5240 784 5265
rect 825 5240 859 5265
rect 900 5240 934 5265
rect 976 5240 1010 5265
rect 1052 5240 1086 5265
rect 1128 5240 1162 5265
rect 1204 5240 1238 5265
rect 1280 5240 1314 5265
rect 1356 5240 1390 5265
rect 1432 5240 1466 5265
rect 1508 5240 1542 5265
rect 1584 5240 1618 5265
rect 1660 5240 1694 5265
rect 1736 5240 1770 5265
rect 1846 5240 1880 5265
rect 1921 5240 1955 5265
rect 1996 5240 2030 5265
rect 2071 5240 2105 5265
rect 2146 5240 2180 5265
rect 2221 5240 2255 5265
rect 2297 5240 2331 5265
rect 2373 5240 2407 5265
rect 2449 5240 2483 5265
rect 2525 5240 2559 5265
rect 2601 5240 2635 5265
rect 2677 5240 2711 5265
rect 2753 5240 2787 5265
rect 2829 5240 2863 5265
rect 2905 5240 2939 5265
rect 2981 5240 3015 5265
rect 525 5197 559 5202
rect 597 5197 631 5202
rect 525 5168 527 5197
rect 527 5168 559 5197
rect 597 5168 629 5197
rect 629 5168 631 5197
rect 675 5168 709 5202
rect 750 5168 784 5202
rect 825 5168 859 5202
rect 900 5168 934 5202
rect 976 5168 1010 5202
rect 1052 5168 1086 5202
rect 1128 5168 1162 5202
rect 1204 5168 1238 5202
rect 1280 5168 1314 5202
rect 1356 5168 1390 5202
rect 1432 5168 1466 5202
rect 1508 5168 1542 5202
rect 1584 5168 1618 5202
rect 1660 5168 1694 5202
rect 1736 5168 1770 5202
rect 1846 5168 1880 5202
rect 1921 5168 1955 5202
rect 1996 5168 2030 5202
rect 2071 5168 2105 5202
rect 2146 5168 2180 5202
rect 2221 5168 2255 5202
rect 2297 5168 2331 5202
rect 2373 5168 2407 5202
rect 2449 5168 2483 5202
rect 2525 5168 2559 5202
rect 2601 5168 2635 5202
rect 2677 5168 2711 5202
rect 2753 5168 2787 5202
rect 2829 5168 2863 5202
rect 2905 5168 2939 5202
rect 2981 5163 3017 5202
rect 3017 5185 3087 5202
rect 3017 5163 3051 5185
rect 525 5095 527 5129
rect 527 5095 559 5129
rect 597 5095 629 5129
rect 629 5095 631 5129
rect 525 5022 527 5056
rect 527 5022 559 5056
rect 597 5022 629 5056
rect 629 5022 631 5056
rect 525 4949 527 4983
rect 527 4949 559 4983
rect 597 4949 629 4983
rect 629 4949 631 4983
rect 525 4876 527 4910
rect 527 4876 559 4910
rect 597 4876 629 4910
rect 629 4876 631 4910
rect 525 4803 527 4837
rect 527 4803 559 4837
rect 597 4803 629 4837
rect 629 4803 631 4837
rect 525 4730 527 4764
rect 527 4730 559 4764
rect 597 4730 629 4764
rect 629 4730 631 4764
rect 525 4657 527 4691
rect 527 4657 559 4691
rect 597 4657 629 4691
rect 629 4657 631 4691
rect 525 4584 527 4618
rect 527 4584 559 4618
rect 597 4584 629 4618
rect 629 4584 631 4618
rect 525 4511 527 4545
rect 527 4511 559 4545
rect 597 4511 629 4545
rect 629 4511 631 4545
rect 525 4438 527 4472
rect 527 4438 559 4472
rect 597 4438 629 4472
rect 629 4438 631 4472
rect 525 4365 527 4399
rect 527 4365 559 4399
rect 597 4365 629 4399
rect 629 4365 631 4399
rect 525 4292 527 4326
rect 527 4292 559 4326
rect 597 4292 629 4326
rect 629 4292 631 4326
rect 525 4219 527 4253
rect 527 4219 559 4253
rect 597 4219 629 4253
rect 629 4219 631 4253
rect 525 4146 527 4180
rect 527 4146 559 4180
rect 597 4146 629 4180
rect 629 4146 631 4180
rect 525 4073 527 4107
rect 527 4073 559 4107
rect 597 4073 629 4107
rect 629 4073 631 4107
rect 525 4000 527 4034
rect 527 4000 559 4034
rect 597 4000 629 4034
rect 629 4000 631 4034
rect 525 3927 527 3961
rect 527 3927 559 3961
rect 597 3927 629 3961
rect 629 3927 631 3961
rect 525 3854 527 3888
rect 527 3854 559 3888
rect 597 3854 629 3888
rect 629 3854 631 3888
rect 525 3781 527 3815
rect 527 3781 559 3815
rect 597 3781 629 3815
rect 629 3781 631 3815
rect 525 3708 527 3742
rect 527 3708 559 3742
rect 597 3708 629 3742
rect 629 3708 631 3742
rect 525 3635 527 3669
rect 527 3635 559 3669
rect 597 3635 629 3669
rect 629 3635 631 3669
rect 525 3562 527 3596
rect 527 3562 559 3596
rect 597 3562 629 3596
rect 629 3562 631 3596
rect 525 3489 527 3523
rect 527 3489 559 3523
rect 597 3489 629 3523
rect 629 3489 631 3523
rect 525 3416 527 3450
rect 527 3416 559 3450
rect 597 3416 629 3450
rect 629 3416 631 3450
rect 525 3343 527 3377
rect 527 3343 559 3377
rect 597 3343 629 3377
rect 629 3343 631 3377
rect 525 3270 527 3304
rect 527 3270 559 3304
rect 597 3270 629 3304
rect 629 3270 631 3304
rect 525 3197 527 3231
rect 527 3197 559 3231
rect 597 3197 629 3231
rect 629 3197 631 3231
rect 525 3124 527 3158
rect 527 3124 559 3158
rect 597 3124 629 3158
rect 629 3124 631 3158
rect 525 3051 527 3085
rect 527 3051 559 3085
rect 597 3051 629 3085
rect 629 3051 631 3085
rect 2981 5151 3051 5163
rect 3051 5151 3085 5185
rect 3085 5151 3087 5185
rect 2981 5117 3087 5151
rect 2981 4016 2983 5117
rect 2983 4016 3085 5117
rect 3085 4016 3087 5117
rect 2981 3943 2983 3977
rect 2983 3943 3015 3977
rect 3053 3943 3085 3977
rect 3085 3943 3087 3977
rect 2981 3870 2983 3904
rect 2983 3870 3015 3904
rect 3053 3870 3085 3904
rect 3085 3870 3087 3904
rect 2981 3797 2983 3831
rect 2983 3797 3015 3831
rect 3053 3797 3085 3831
rect 3085 3797 3087 3831
rect 2981 3724 2983 3758
rect 2983 3724 3015 3758
rect 3053 3724 3085 3758
rect 3085 3724 3087 3758
rect 2981 3651 2983 3685
rect 2983 3651 3015 3685
rect 3053 3651 3085 3685
rect 3085 3651 3087 3685
rect 2981 3578 2983 3612
rect 2983 3578 3015 3612
rect 3053 3578 3085 3612
rect 3085 3578 3087 3612
rect 2981 3505 2983 3539
rect 2983 3505 3015 3539
rect 3053 3505 3085 3539
rect 3085 3505 3087 3539
rect 2981 3432 2983 3466
rect 2983 3432 3015 3466
rect 3053 3432 3085 3466
rect 3085 3432 3087 3466
rect 2981 3359 2983 3393
rect 2983 3359 3015 3393
rect 3053 3359 3085 3393
rect 3085 3359 3087 3393
rect 2981 3286 2983 3320
rect 2983 3286 3015 3320
rect 3053 3286 3085 3320
rect 3085 3286 3087 3320
rect 2981 3213 2983 3247
rect 2983 3213 3015 3247
rect 3053 3213 3085 3247
rect 3085 3213 3087 3247
rect 2981 3140 2983 3174
rect 2983 3140 3015 3174
rect 3053 3140 3085 3174
rect 3085 3140 3087 3174
rect 2981 3067 2983 3101
rect 2983 3067 3015 3101
rect 3053 3067 3085 3101
rect 3085 3067 3087 3101
rect 525 2978 527 3012
rect 527 2978 559 3012
rect 597 2978 629 3012
rect 629 2978 631 3012
rect 774 3007 792 3041
rect 792 3007 808 3041
rect 847 3007 861 3041
rect 861 3007 881 3041
rect 920 3007 930 3041
rect 930 3007 954 3041
rect 993 3007 999 3041
rect 999 3007 1027 3041
rect 1066 3007 1068 3041
rect 1068 3007 1100 3041
rect 1139 3007 1172 3041
rect 1172 3007 1173 3041
rect 1211 3007 1241 3041
rect 1241 3007 1245 3041
rect 1283 3007 1310 3041
rect 1310 3007 1317 3041
rect 1355 3007 1379 3041
rect 1379 3007 1389 3041
rect 1427 3007 1448 3041
rect 1448 3007 1461 3041
rect 1499 3007 1517 3041
rect 1517 3007 1533 3041
rect 1571 3007 1586 3041
rect 1586 3007 1605 3041
rect 1643 3007 1655 3041
rect 1655 3007 1677 3041
rect 1715 3007 1724 3041
rect 1724 3007 1749 3041
rect 1787 3007 1793 3041
rect 1793 3007 1821 3041
rect 1859 3007 1862 3041
rect 1862 3007 1893 3041
rect 1931 3007 1965 3041
rect 2003 3007 2034 3041
rect 2034 3007 2037 3041
rect 2075 3007 2103 3041
rect 2103 3007 2109 3041
rect 2147 3007 2172 3041
rect 2172 3007 2181 3041
rect 2219 3007 2241 3041
rect 2241 3007 2253 3041
rect 2291 3007 2310 3041
rect 2310 3007 2325 3041
rect 2363 3007 2378 3041
rect 2378 3007 2397 3041
rect 2435 3007 2446 3041
rect 2446 3007 2469 3041
rect 2507 3007 2514 3041
rect 2514 3007 2541 3041
rect 2579 3007 2582 3041
rect 2582 3007 2613 3041
rect 2651 3007 2684 3041
rect 2684 3007 2685 3041
rect 2723 3007 2752 3041
rect 2752 3007 2757 3041
rect 2795 3007 2820 3041
rect 2820 3007 2829 3041
rect 525 2905 527 2939
rect 527 2905 559 2939
rect 597 2905 629 2939
rect 629 2905 631 2939
rect 2981 2994 2983 3028
rect 2983 2994 3015 3028
rect 3053 2994 3085 3028
rect 3085 2994 3087 3028
rect 2981 2921 2983 2955
rect 2983 2921 3015 2955
rect 3053 2921 3085 2955
rect 3085 2921 3087 2955
rect 774 2887 792 2921
rect 792 2887 808 2921
rect 847 2887 861 2921
rect 861 2887 881 2921
rect 920 2887 930 2921
rect 930 2887 954 2921
rect 993 2887 999 2921
rect 999 2887 1027 2921
rect 1066 2887 1068 2921
rect 1068 2887 1100 2921
rect 1139 2887 1172 2921
rect 1172 2887 1173 2921
rect 1211 2887 1241 2921
rect 1241 2887 1245 2921
rect 1283 2887 1310 2921
rect 1310 2887 1317 2921
rect 1355 2887 1379 2921
rect 1379 2887 1389 2921
rect 1427 2887 1448 2921
rect 1448 2887 1461 2921
rect 1499 2887 1517 2921
rect 1517 2887 1533 2921
rect 1571 2887 1586 2921
rect 1586 2887 1605 2921
rect 1643 2887 1655 2921
rect 1655 2887 1677 2921
rect 1715 2887 1724 2921
rect 1724 2887 1749 2921
rect 1787 2887 1793 2921
rect 1793 2887 1821 2921
rect 1859 2887 1862 2921
rect 1862 2887 1893 2921
rect 1931 2887 1965 2921
rect 2003 2887 2034 2921
rect 2034 2887 2037 2921
rect 2075 2887 2103 2921
rect 2103 2887 2109 2921
rect 2147 2887 2172 2921
rect 2172 2887 2181 2921
rect 2219 2887 2241 2921
rect 2241 2887 2253 2921
rect 2291 2887 2310 2921
rect 2310 2887 2325 2921
rect 2363 2887 2378 2921
rect 2378 2887 2397 2921
rect 2435 2887 2446 2921
rect 2446 2887 2469 2921
rect 2507 2887 2514 2921
rect 2514 2887 2541 2921
rect 2579 2887 2582 2921
rect 2582 2887 2613 2921
rect 2651 2887 2684 2921
rect 2684 2887 2685 2921
rect 2723 2887 2752 2921
rect 2752 2887 2757 2921
rect 2795 2887 2820 2921
rect 2820 2887 2829 2921
rect 525 2832 527 2866
rect 527 2832 559 2866
rect 597 2832 629 2866
rect 629 2832 631 2866
rect 525 2759 527 2793
rect 527 2759 559 2793
rect 597 2759 629 2793
rect 629 2759 631 2793
rect 525 2686 527 2720
rect 527 2686 559 2720
rect 597 2686 629 2720
rect 629 2686 631 2720
rect 525 2613 527 2647
rect 527 2613 559 2647
rect 597 2613 629 2647
rect 629 2613 631 2647
rect 525 2540 527 2574
rect 527 2540 559 2574
rect 597 2540 629 2574
rect 629 2540 631 2574
rect 525 2467 527 2501
rect 527 2467 559 2501
rect 597 2467 629 2501
rect 629 2467 631 2501
rect 525 2394 527 2428
rect 527 2394 559 2428
rect 597 2394 629 2428
rect 629 2394 631 2428
rect 525 2321 527 2355
rect 527 2321 559 2355
rect 597 2321 629 2355
rect 629 2321 631 2355
rect 525 2248 527 2282
rect 527 2248 559 2282
rect 597 2248 629 2282
rect 629 2248 631 2282
rect 525 2175 527 2209
rect 527 2175 559 2209
rect 597 2175 629 2209
rect 629 2175 631 2209
rect 525 2102 527 2136
rect 527 2102 559 2136
rect 597 2102 629 2136
rect 629 2102 631 2136
rect 525 2029 527 2063
rect 527 2029 559 2063
rect 597 2029 629 2063
rect 629 2029 631 2063
rect 525 1956 527 1990
rect 527 1956 559 1990
rect 597 1956 629 1990
rect 629 1956 631 1990
rect 525 879 527 1917
rect 527 879 629 1917
rect 629 879 631 1917
rect 525 765 631 879
rect 2981 2848 2983 2882
rect 2983 2848 3015 2882
rect 3053 2848 3085 2882
rect 3085 2848 3087 2882
rect 2981 2775 2983 2809
rect 2983 2775 3015 2809
rect 3053 2775 3085 2809
rect 3085 2775 3087 2809
rect 2981 2702 2983 2736
rect 2983 2702 3015 2736
rect 3053 2702 3085 2736
rect 3085 2702 3087 2736
rect 2981 2629 2983 2663
rect 2983 2629 3015 2663
rect 3053 2629 3085 2663
rect 3085 2629 3087 2663
rect 2981 2556 2983 2590
rect 2983 2556 3015 2590
rect 3053 2556 3085 2590
rect 3085 2556 3087 2590
rect 2981 2483 2983 2517
rect 2983 2483 3015 2517
rect 3053 2483 3085 2517
rect 3085 2483 3087 2517
rect 2981 2410 2983 2444
rect 2983 2410 3015 2444
rect 3053 2410 3085 2444
rect 3085 2410 3087 2444
rect 2981 2337 2983 2371
rect 2983 2337 3015 2371
rect 3053 2337 3085 2371
rect 3085 2337 3087 2371
rect 2981 2264 2983 2298
rect 2983 2264 3015 2298
rect 3053 2264 3085 2298
rect 3085 2264 3087 2298
rect 2981 2191 2983 2225
rect 2983 2191 3015 2225
rect 3053 2191 3085 2225
rect 3085 2191 3087 2225
rect 2981 2118 2983 2152
rect 2983 2118 3015 2152
rect 3053 2118 3085 2152
rect 3085 2118 3087 2152
rect 2981 2045 2983 2079
rect 2983 2045 3015 2079
rect 3053 2045 3085 2079
rect 3085 2045 3087 2079
rect 2981 1972 2983 2006
rect 2983 1972 3015 2006
rect 3053 1972 3085 2006
rect 3085 1972 3087 2006
rect 2981 1899 2983 1933
rect 2983 1899 3015 1933
rect 3053 1899 3085 1933
rect 3085 1899 3087 1933
rect 2981 1826 2983 1860
rect 2983 1826 3015 1860
rect 3053 1826 3085 1860
rect 3085 1826 3087 1860
rect 2981 1753 2983 1787
rect 2983 1753 3015 1787
rect 3053 1753 3085 1787
rect 3085 1753 3087 1787
rect 2981 1680 2983 1714
rect 2983 1680 3015 1714
rect 3053 1680 3085 1714
rect 3085 1680 3087 1714
rect 2981 1607 2983 1641
rect 2983 1607 3015 1641
rect 3053 1607 3085 1641
rect 3085 1607 3087 1641
rect 2981 1534 2983 1568
rect 2983 1534 3015 1568
rect 3053 1534 3085 1568
rect 3085 1534 3087 1568
rect 2981 1461 2983 1495
rect 2983 1461 3015 1495
rect 3053 1461 3085 1495
rect 3085 1461 3087 1495
rect 2981 1388 2983 1422
rect 2983 1388 3015 1422
rect 3053 1388 3085 1422
rect 3085 1388 3087 1422
rect 2981 1315 2983 1349
rect 2983 1315 3015 1349
rect 3053 1315 3085 1349
rect 3085 1315 3087 1349
rect 2981 1242 2983 1276
rect 2983 1242 3015 1276
rect 3053 1242 3085 1276
rect 3085 1242 3087 1276
rect 2981 1169 2983 1203
rect 2983 1169 3015 1203
rect 3053 1169 3085 1203
rect 3085 1169 3087 1203
rect 2981 1096 2983 1130
rect 2983 1096 3015 1130
rect 3053 1096 3085 1130
rect 3085 1096 3087 1130
rect 2981 1023 2983 1057
rect 2983 1023 3015 1057
rect 3053 1023 3085 1057
rect 3085 1023 3087 1057
rect 2981 950 2983 984
rect 2983 950 3015 984
rect 3053 950 3085 984
rect 3085 950 3087 984
rect 2981 877 2983 911
rect 2983 877 3015 911
rect 3053 877 3085 911
rect 3085 877 3087 911
rect 2981 804 2983 838
rect 2983 804 3015 838
rect 3053 804 3085 838
rect 3085 804 3087 838
rect 525 731 595 765
rect 595 731 631 765
rect 670 731 704 765
rect 743 731 777 765
rect 816 731 850 765
rect 889 731 923 765
rect 962 731 996 765
rect 1035 731 1069 765
rect 1108 731 1142 765
rect 597 663 631 693
rect 670 663 704 693
rect 743 663 777 693
rect 816 663 850 693
rect 889 663 923 693
rect 962 663 996 693
rect 1035 663 1069 693
rect 1108 663 1142 693
rect 1181 663 2941 765
rect 2941 731 2983 765
rect 2983 731 3015 765
rect 3053 731 3085 765
rect 3085 731 3087 765
rect 2941 697 3015 731
rect 2941 663 2975 697
rect 2975 663 3009 697
rect 3009 663 3015 697
rect 597 659 631 663
rect 670 659 704 663
rect 743 659 777 663
rect 816 659 850 663
rect 889 659 923 663
rect 962 659 996 663
rect 1035 659 1069 663
rect 1108 659 1142 663
rect 1181 659 3015 663
rect 3253 5248 3287 5258
rect 3253 5224 3286 5248
rect 3286 5224 3287 5248
rect 3253 5180 3287 5186
rect 3253 5152 3286 5180
rect 3286 5152 3287 5180
rect 3253 5112 3287 5114
rect 3253 5080 3286 5112
rect 3286 5080 3287 5112
rect 3253 5010 3286 5042
rect 3286 5010 3287 5042
rect 3253 5008 3287 5010
rect 3253 4942 3286 4970
rect 3286 4942 3287 4970
rect 3253 4936 3287 4942
rect 3253 4874 3286 4898
rect 3286 4874 3287 4898
rect 3253 4864 3287 4874
rect 3253 4806 3286 4826
rect 3286 4806 3287 4826
rect 3253 4792 3287 4806
rect 3253 4738 3286 4754
rect 3286 4738 3287 4754
rect 3253 4720 3287 4738
rect 3253 4670 3286 4682
rect 3286 4670 3287 4682
rect 3253 4648 3287 4670
rect 3253 4602 3286 4610
rect 3286 4602 3287 4610
rect 3253 4576 3287 4602
rect 3253 4534 3286 4538
rect 3286 4534 3287 4538
rect 3253 4504 3287 4534
rect 3253 4432 3287 4466
rect 3253 4364 3287 4394
rect 3253 4360 3286 4364
rect 3286 4360 3287 4364
rect 3253 4296 3287 4322
rect 3253 4288 3286 4296
rect 3286 4288 3287 4296
rect 3253 4228 3287 4250
rect 3253 4216 3286 4228
rect 3286 4216 3287 4228
rect 3253 4160 3287 4178
rect 3253 4144 3286 4160
rect 3286 4144 3287 4160
rect 3253 4092 3287 4106
rect 3253 4072 3286 4092
rect 3286 4072 3287 4092
rect 3253 4024 3287 4034
rect 3253 4000 3286 4024
rect 3286 4000 3287 4024
rect 3253 3956 3287 3962
rect 3253 3928 3286 3956
rect 3286 3928 3287 3956
rect 3253 3888 3287 3890
rect 3253 3856 3286 3888
rect 3286 3856 3287 3888
rect 3253 3786 3286 3818
rect 3286 3786 3287 3818
rect 3253 3784 3287 3786
rect 3253 3718 3286 3746
rect 3286 3718 3287 3746
rect 3253 3712 3287 3718
rect 3253 3650 3286 3674
rect 3286 3650 3287 3674
rect 3253 3640 3287 3650
rect 3253 3582 3286 3602
rect 3286 3582 3287 3602
rect 3253 3568 3287 3582
rect 3253 3514 3286 3530
rect 3286 3514 3287 3530
rect 3253 3496 3287 3514
rect 3253 3446 3286 3458
rect 3286 3446 3287 3458
rect 3253 3424 3287 3446
rect 3253 3378 3286 3386
rect 3286 3378 3287 3386
rect 3253 3352 3287 3378
rect 3253 3310 3286 3314
rect 3286 3310 3287 3314
rect 3253 3280 3287 3310
rect 3253 3208 3287 3242
rect 3253 3140 3287 3170
rect 3253 3136 3286 3140
rect 3286 3136 3287 3140
rect 3253 3072 3287 3098
rect 3253 3064 3286 3072
rect 3286 3064 3287 3072
rect 3253 3004 3287 3026
rect 3253 2992 3286 3004
rect 3286 2992 3287 3004
rect 3253 2936 3287 2954
rect 3253 2920 3286 2936
rect 3286 2920 3287 2936
rect 3253 2868 3287 2882
rect 3253 2848 3286 2868
rect 3286 2848 3287 2868
rect 3253 2800 3287 2810
rect 3253 2776 3286 2800
rect 3286 2776 3287 2800
rect 3253 2732 3287 2738
rect 3253 2704 3286 2732
rect 3286 2704 3287 2732
rect 3253 2664 3287 2666
rect 3253 2632 3286 2664
rect 3286 2632 3287 2664
rect 3253 2562 3286 2594
rect 3286 2562 3287 2594
rect 3253 2560 3287 2562
rect 3253 2494 3286 2522
rect 3286 2494 3287 2522
rect 3253 2488 3287 2494
rect 3253 2426 3286 2450
rect 3286 2426 3287 2450
rect 3253 2416 3287 2426
rect 3253 2358 3286 2378
rect 3286 2358 3287 2378
rect 3253 2344 3287 2358
rect 3253 2290 3286 2306
rect 3286 2290 3287 2306
rect 3253 2272 3287 2290
rect 3253 2222 3286 2234
rect 3286 2222 3287 2234
rect 3253 2200 3287 2222
rect 3253 2154 3286 2162
rect 3286 2154 3287 2162
rect 3253 2128 3287 2154
rect 3253 2086 3286 2090
rect 3286 2086 3287 2090
rect 3253 2056 3287 2086
rect 3253 1984 3287 2018
rect 3253 1916 3287 1946
rect 3253 1912 3286 1916
rect 3286 1912 3287 1916
rect 3253 1848 3287 1874
rect 3253 1840 3286 1848
rect 3286 1840 3287 1848
rect 3253 1780 3287 1801
rect 3253 1767 3286 1780
rect 3286 1767 3287 1780
rect 3253 1712 3287 1728
rect 3253 1694 3286 1712
rect 3286 1694 3287 1712
rect 3253 1644 3287 1655
rect 3253 1621 3286 1644
rect 3286 1621 3287 1644
rect 3253 1576 3287 1582
rect 3253 1548 3286 1576
rect 3286 1548 3287 1576
rect 3253 1508 3287 1509
rect 3253 1475 3286 1508
rect 3286 1475 3287 1508
rect 3253 1406 3286 1436
rect 3286 1406 3287 1436
rect 3253 1402 3287 1406
rect 3253 1338 3286 1363
rect 3286 1338 3287 1363
rect 3253 1329 3287 1338
rect 3253 1270 3286 1290
rect 3286 1270 3287 1290
rect 3253 1256 3287 1270
rect 3253 1202 3286 1217
rect 3286 1202 3287 1217
rect 3253 1183 3287 1202
rect 3253 1134 3286 1144
rect 3286 1134 3287 1144
rect 3253 1110 3287 1134
rect 3253 1066 3286 1071
rect 3286 1066 3287 1071
rect 3253 1037 3287 1066
rect 3253 964 3287 998
rect 3253 896 3287 925
rect 3253 891 3286 896
rect 3286 891 3287 896
rect 3253 828 3287 852
rect 3253 818 3286 828
rect 3286 818 3287 828
rect 3253 760 3287 779
rect 3253 745 3286 760
rect 3286 745 3287 760
rect 3253 692 3287 706
rect 3253 672 3286 692
rect 3286 672 3287 692
rect 326 612 360 632
rect 326 598 360 612
rect 326 526 360 560
rect 3253 624 3287 633
rect 3253 599 3286 624
rect 3286 599 3287 624
rect 3253 556 3287 560
rect 3253 526 3286 556
rect 3286 526 3287 556
rect 398 454 428 488
rect 428 454 432 488
rect 472 454 496 488
rect 496 454 506 488
rect 546 454 564 488
rect 564 454 580 488
rect 620 454 632 488
rect 632 454 654 488
rect 694 454 700 488
rect 700 454 728 488
rect 768 454 802 488
rect 842 454 870 488
rect 870 454 876 488
rect 916 454 938 488
rect 938 454 950 488
rect 990 454 1006 488
rect 1006 454 1024 488
rect 1063 454 1074 488
rect 1074 454 1097 488
rect 1136 454 1142 488
rect 1142 454 1170 488
rect 1209 454 1210 488
rect 1210 454 1243 488
rect 1282 454 1312 488
rect 1312 454 1316 488
rect 1355 454 1380 488
rect 1380 454 1389 488
rect 1428 454 1448 488
rect 1448 454 1462 488
rect 1501 454 1516 488
rect 1516 454 1535 488
rect 1574 454 1584 488
rect 1584 454 1608 488
rect 1647 454 1652 488
rect 1652 454 1681 488
rect 1720 454 1754 488
rect 1793 454 1822 488
rect 1822 454 1827 488
rect 1866 454 1890 488
rect 1890 454 1900 488
rect 1939 454 1958 488
rect 1958 454 1973 488
rect 2012 454 2026 488
rect 2026 454 2046 488
rect 2085 454 2094 488
rect 2094 454 2119 488
rect 2158 454 2162 488
rect 2162 454 2192 488
rect 2231 454 2264 488
rect 2264 454 2265 488
rect 2304 454 2332 488
rect 2332 454 2338 488
rect 2377 454 2400 488
rect 2400 454 2411 488
rect 2450 454 2468 488
rect 2468 454 2484 488
rect 2523 454 2536 488
rect 2536 454 2557 488
rect 2596 454 2604 488
rect 2604 454 2630 488
rect 2669 454 2672 488
rect 2672 454 2703 488
rect 2742 454 2774 488
rect 2774 454 2776 488
rect 2815 454 2842 488
rect 2842 454 2849 488
rect 2888 454 2910 488
rect 2910 454 2922 488
rect 2961 454 2978 488
rect 2978 454 2995 488
rect 3034 454 3046 488
rect 3046 454 3068 488
rect 3107 454 3114 488
rect 3114 454 3141 488
rect 3180 454 3182 488
rect 3182 454 3214 488
rect 3469 5419 3473 5453
rect 3473 5419 3503 5453
rect 3541 5419 3575 5453
rect 3613 5419 3643 5453
rect 3643 5419 3647 5453
rect 3469 5346 3473 5380
rect 3473 5346 3503 5380
rect 3541 5346 3575 5380
rect 3613 5346 3643 5380
rect 3643 5346 3647 5380
rect 3469 5273 3473 5307
rect 3473 5273 3503 5307
rect 3541 5273 3575 5307
rect 3613 5273 3643 5307
rect 3643 5273 3647 5307
rect 3469 5200 3473 5234
rect 3473 5200 3503 5234
rect 3541 5200 3575 5234
rect 3613 5200 3643 5234
rect 3643 5200 3647 5234
rect 3469 5127 3473 5161
rect 3473 5127 3503 5161
rect 3541 5127 3575 5161
rect 3613 5127 3643 5161
rect 3643 5127 3647 5161
rect 3469 5054 3473 5088
rect 3473 5054 3503 5088
rect 3541 5054 3575 5088
rect 3613 5054 3643 5088
rect 3643 5054 3647 5088
rect 3469 4981 3473 5015
rect 3473 4981 3503 5015
rect 3541 4981 3575 5015
rect 3613 4981 3643 5015
rect 3643 4981 3647 5015
rect 3469 4908 3473 4942
rect 3473 4908 3503 4942
rect 3541 4908 3575 4942
rect 3613 4908 3643 4942
rect 3643 4908 3647 4942
rect 3469 4835 3473 4869
rect 3473 4835 3503 4869
rect 3541 4835 3575 4869
rect 3613 4835 3643 4869
rect 3643 4835 3647 4869
rect 3469 4762 3473 4796
rect 3473 4762 3503 4796
rect 3541 4762 3575 4796
rect 3613 4762 3643 4796
rect 3643 4762 3647 4796
rect 3469 4689 3473 4723
rect 3473 4689 3503 4723
rect 3541 4689 3575 4723
rect 3613 4689 3643 4723
rect 3643 4689 3647 4723
rect 3469 4616 3473 4650
rect 3473 4616 3503 4650
rect 3541 4616 3575 4650
rect 3613 4616 3643 4650
rect 3643 4616 3647 4650
rect 3469 4543 3473 4577
rect 3473 4543 3503 4577
rect 3541 4543 3575 4577
rect 3613 4543 3643 4577
rect 3643 4543 3647 4577
rect 3469 4470 3473 4504
rect 3473 4470 3503 4504
rect 3541 4470 3575 4504
rect 3613 4470 3643 4504
rect 3643 4470 3647 4504
rect 3469 4397 3473 4431
rect 3473 4397 3503 4431
rect 3541 4397 3575 4431
rect 3613 4397 3643 4431
rect 3643 4397 3647 4431
rect 3469 4324 3473 4358
rect 3473 4324 3503 4358
rect 3541 4324 3575 4358
rect 3613 4324 3643 4358
rect 3643 4324 3647 4358
rect 3469 4251 3473 4285
rect 3473 4251 3503 4285
rect 3541 4251 3575 4285
rect 3613 4251 3643 4285
rect 3643 4251 3647 4285
rect 3469 4178 3473 4212
rect 3473 4178 3503 4212
rect 3541 4178 3575 4212
rect 3613 4178 3643 4212
rect 3643 4178 3647 4212
rect 3469 4105 3473 4139
rect 3473 4105 3503 4139
rect 3541 4105 3575 4139
rect 3613 4105 3643 4139
rect 3643 4105 3647 4139
rect 3469 4032 3473 4066
rect 3473 4032 3503 4066
rect 3541 4032 3575 4066
rect 3613 4032 3643 4066
rect 3643 4032 3647 4066
rect 3469 3959 3473 3993
rect 3473 3959 3503 3993
rect 3541 3959 3575 3993
rect 3613 3959 3643 3993
rect 3643 3959 3647 3993
rect 3469 3886 3473 3920
rect 3473 3886 3503 3920
rect 3541 3886 3575 3920
rect 3613 3886 3643 3920
rect 3643 3886 3647 3920
rect 3469 3813 3473 3847
rect 3473 3813 3503 3847
rect 3541 3813 3575 3847
rect 3613 3813 3643 3847
rect 3643 3813 3647 3847
rect 3469 3740 3473 3774
rect 3473 3740 3503 3774
rect 3541 3740 3575 3774
rect 3613 3740 3643 3774
rect 3643 3740 3647 3774
rect 3469 3667 3473 3701
rect 3473 3667 3503 3701
rect 3541 3667 3575 3701
rect 3613 3667 3643 3701
rect 3643 3667 3647 3701
rect 3469 3594 3473 3628
rect 3473 3594 3503 3628
rect 3541 3594 3575 3628
rect 3613 3594 3643 3628
rect 3643 3594 3647 3628
rect 3469 3521 3473 3555
rect 3473 3521 3503 3555
rect 3541 3521 3575 3555
rect 3613 3521 3643 3555
rect 3643 3521 3647 3555
rect 3469 3448 3473 3482
rect 3473 3448 3503 3482
rect 3541 3448 3575 3482
rect 3613 3448 3643 3482
rect 3643 3448 3647 3482
rect 3469 3375 3473 3409
rect 3473 3375 3503 3409
rect 3541 3375 3575 3409
rect 3613 3375 3643 3409
rect 3643 3375 3647 3409
rect 3469 3302 3473 3336
rect 3473 3302 3503 3336
rect 3541 3302 3575 3336
rect 3613 3302 3643 3336
rect 3643 3302 3647 3336
rect 3469 3229 3473 3263
rect 3473 3229 3503 3263
rect 3541 3229 3575 3263
rect 3613 3229 3643 3263
rect 3643 3229 3647 3263
rect 3469 3156 3473 3190
rect 3473 3156 3503 3190
rect 3541 3156 3575 3190
rect 3613 3156 3643 3190
rect 3643 3156 3647 3190
rect 3469 3083 3473 3117
rect 3473 3083 3503 3117
rect 3541 3083 3575 3117
rect 3613 3083 3643 3117
rect 3643 3083 3647 3117
rect 3469 3010 3473 3044
rect 3473 3010 3503 3044
rect 3541 3010 3575 3044
rect 3613 3010 3643 3044
rect 3643 3010 3647 3044
rect 3469 2937 3473 2971
rect 3473 2937 3503 2971
rect 3541 2937 3575 2971
rect 3613 2937 3643 2971
rect 3643 2937 3647 2971
rect 3469 2864 3473 2898
rect 3473 2864 3503 2898
rect 3541 2864 3575 2898
rect 3613 2864 3643 2898
rect 3643 2864 3647 2898
rect 3469 2791 3473 2825
rect 3473 2791 3503 2825
rect 3541 2791 3575 2825
rect 3613 2791 3643 2825
rect 3643 2791 3647 2825
rect 3469 2718 3473 2752
rect 3473 2718 3503 2752
rect 3541 2718 3575 2752
rect 3613 2718 3643 2752
rect 3643 2718 3647 2752
rect 3469 2645 3473 2679
rect 3473 2645 3503 2679
rect 3541 2645 3575 2679
rect 3613 2645 3643 2679
rect 3643 2645 3647 2679
rect 3469 2572 3473 2606
rect 3473 2572 3503 2606
rect 3541 2572 3575 2606
rect 3613 2572 3643 2606
rect 3643 2572 3647 2606
rect 4592 5656 4770 5710
rect 4592 5638 4596 5656
rect 4596 5638 4766 5656
rect 4766 5638 4770 5656
rect 4592 5565 4596 5599
rect 4596 5565 4626 5599
rect 4664 5565 4698 5599
rect 4736 5565 4766 5599
rect 4766 5565 4770 5599
rect 4592 5492 4596 5526
rect 4596 5492 4626 5526
rect 4664 5492 4698 5526
rect 4736 5492 4766 5526
rect 4766 5492 4770 5526
rect 10277 5637 10279 5671
rect 10279 5637 10311 5671
rect 10349 5637 10381 5671
rect 10381 5637 10383 5671
rect 10277 5564 10279 5598
rect 10279 5564 10311 5598
rect 10349 5564 10381 5598
rect 10381 5564 10383 5598
rect 10277 5491 10279 5525
rect 10279 5491 10311 5525
rect 10349 5491 10381 5525
rect 10381 5491 10383 5525
rect 4592 5419 4596 5453
rect 4596 5419 4626 5453
rect 4664 5419 4698 5453
rect 4736 5419 4766 5453
rect 4766 5419 4770 5453
rect 4592 5346 4596 5380
rect 4596 5346 4626 5380
rect 4664 5346 4698 5380
rect 4736 5346 4766 5380
rect 4766 5346 4770 5380
rect 4592 5273 4596 5307
rect 4596 5273 4626 5307
rect 4664 5273 4698 5307
rect 4736 5273 4766 5307
rect 4766 5273 4770 5307
rect 4592 5200 4596 5234
rect 4596 5200 4626 5234
rect 4664 5200 4698 5234
rect 4736 5200 4766 5234
rect 4766 5200 4770 5234
rect 4592 5127 4596 5161
rect 4596 5127 4626 5161
rect 4664 5127 4698 5161
rect 4736 5127 4766 5161
rect 4766 5127 4770 5161
rect 4592 5054 4596 5088
rect 4596 5054 4626 5088
rect 4664 5054 4698 5088
rect 4736 5054 4766 5088
rect 4766 5054 4770 5088
rect 4592 4981 4596 5015
rect 4596 4981 4626 5015
rect 4664 4981 4698 5015
rect 4736 4981 4766 5015
rect 4766 4981 4770 5015
rect 4592 4908 4596 4942
rect 4596 4908 4626 4942
rect 4664 4908 4698 4942
rect 4736 4908 4766 4942
rect 4766 4908 4770 4942
rect 4592 4835 4596 4869
rect 4596 4835 4626 4869
rect 4664 4835 4698 4869
rect 4736 4835 4766 4869
rect 4766 4835 4770 4869
rect 4592 4762 4596 4796
rect 4596 4762 4626 4796
rect 4664 4762 4698 4796
rect 4736 4762 4766 4796
rect 4766 4762 4770 4796
rect 4592 4689 4596 4723
rect 4596 4689 4626 4723
rect 4664 4689 4698 4723
rect 4736 4689 4766 4723
rect 4766 4689 4770 4723
rect 4592 4616 4596 4650
rect 4596 4616 4626 4650
rect 4664 4616 4698 4650
rect 4736 4616 4766 4650
rect 4766 4616 4770 4650
rect 4592 4543 4596 4577
rect 4596 4543 4626 4577
rect 4664 4543 4698 4577
rect 4736 4543 4766 4577
rect 4766 4543 4770 4577
rect 4592 4470 4596 4504
rect 4596 4470 4626 4504
rect 4664 4470 4698 4504
rect 4736 4470 4766 4504
rect 4766 4470 4770 4504
rect 4592 4397 4596 4431
rect 4596 4397 4626 4431
rect 4664 4397 4698 4431
rect 4736 4397 4766 4431
rect 4766 4397 4770 4431
rect 4592 4324 4596 4358
rect 4596 4324 4626 4358
rect 4664 4324 4698 4358
rect 4736 4324 4766 4358
rect 4766 4324 4770 4358
rect 4592 4251 4596 4285
rect 4596 4251 4626 4285
rect 4664 4251 4698 4285
rect 4736 4251 4766 4285
rect 4766 4251 4770 4285
rect 4592 4178 4596 4212
rect 4596 4178 4626 4212
rect 4664 4178 4698 4212
rect 4736 4178 4766 4212
rect 4766 4178 4770 4212
rect 4592 4105 4596 4139
rect 4596 4105 4626 4139
rect 4664 4105 4698 4139
rect 4736 4105 4766 4139
rect 4766 4105 4770 4139
rect 4592 4032 4596 4066
rect 4596 4032 4626 4066
rect 4664 4032 4698 4066
rect 4736 4032 4766 4066
rect 4766 4032 4770 4066
rect 4592 3959 4596 3993
rect 4596 3959 4626 3993
rect 4664 3959 4698 3993
rect 4736 3959 4766 3993
rect 4766 3959 4770 3993
rect 4592 3886 4596 3920
rect 4596 3886 4626 3920
rect 4664 3886 4698 3920
rect 4736 3886 4766 3920
rect 4766 3886 4770 3920
rect 4592 3813 4596 3847
rect 4596 3813 4626 3847
rect 4664 3813 4698 3847
rect 4736 3813 4766 3847
rect 4766 3813 4770 3847
rect 4592 3740 4596 3774
rect 4596 3740 4626 3774
rect 4664 3740 4698 3774
rect 4736 3740 4766 3774
rect 4766 3740 4770 3774
rect 4592 3667 4596 3701
rect 4596 3667 4626 3701
rect 4664 3667 4698 3701
rect 4736 3667 4766 3701
rect 4766 3667 4770 3701
rect 4592 3594 4596 3628
rect 4596 3594 4626 3628
rect 4664 3594 4698 3628
rect 4736 3594 4766 3628
rect 4766 3594 4770 3628
rect 4592 3521 4596 3555
rect 4596 3521 4626 3555
rect 4664 3521 4698 3555
rect 4736 3521 4766 3555
rect 4766 3521 4770 3555
rect 4592 3448 4596 3482
rect 4596 3448 4626 3482
rect 4664 3448 4698 3482
rect 4736 3448 4766 3482
rect 4766 3448 4770 3482
rect 4592 3375 4596 3409
rect 4596 3375 4626 3409
rect 4664 3375 4698 3409
rect 4736 3375 4766 3409
rect 4766 3375 4770 3409
rect 4592 3302 4596 3336
rect 4596 3302 4626 3336
rect 4664 3302 4698 3336
rect 4736 3302 4766 3336
rect 4766 3302 4770 3336
rect 4592 3229 4596 3263
rect 4596 3229 4626 3263
rect 4664 3229 4698 3263
rect 4736 3229 4766 3263
rect 4766 3229 4770 3263
rect 4592 3156 4596 3190
rect 4596 3156 4626 3190
rect 4664 3156 4698 3190
rect 4736 3156 4766 3190
rect 4766 3156 4770 3190
rect 4592 3083 4596 3117
rect 4596 3083 4626 3117
rect 4664 3083 4698 3117
rect 4736 3083 4766 3117
rect 4766 3083 4770 3117
rect 4592 3010 4596 3044
rect 4596 3010 4626 3044
rect 4664 3010 4698 3044
rect 4736 3010 4766 3044
rect 4766 3010 4770 3044
rect 4592 2937 4596 2971
rect 4596 2937 4626 2971
rect 4664 2937 4698 2971
rect 4736 2937 4766 2971
rect 4766 2937 4770 2971
rect 4592 2864 4596 2898
rect 4596 2864 4626 2898
rect 4664 2864 4698 2898
rect 4736 2864 4766 2898
rect 4766 2864 4770 2898
rect 4592 2791 4596 2825
rect 4596 2791 4626 2825
rect 4664 2791 4698 2825
rect 4736 2791 4766 2825
rect 4766 2791 4770 2825
rect 4592 2718 4596 2752
rect 4596 2718 4626 2752
rect 4664 2718 4698 2752
rect 4736 2718 4766 2752
rect 4766 2718 4770 2752
rect 4592 2645 4596 2679
rect 4596 2645 4626 2679
rect 4664 2645 4698 2679
rect 4736 2645 4766 2679
rect 4766 2645 4770 2679
rect 4592 2572 4596 2606
rect 4596 2572 4626 2606
rect 4664 2572 4698 2606
rect 4736 2572 4766 2606
rect 4766 2572 4770 2606
rect 3469 2499 3473 2533
rect 3473 2499 3503 2533
rect 3541 2499 3575 2533
rect 3613 2499 3643 2533
rect 3643 2499 3647 2533
rect 3992 2530 3993 2564
rect 3993 2530 4026 2564
rect 4084 2530 4088 2564
rect 4088 2530 4118 2564
rect 4177 2530 4183 2564
rect 4183 2530 4211 2564
rect 4592 2499 4596 2533
rect 4596 2499 4626 2533
rect 4664 2499 4698 2533
rect 4736 2499 4766 2533
rect 4766 2499 4770 2533
rect 3469 2426 3473 2460
rect 3473 2426 3503 2460
rect 3541 2426 3575 2460
rect 3613 2426 3643 2460
rect 3643 2426 3647 2460
rect 3469 2353 3473 2387
rect 3473 2353 3503 2387
rect 3541 2353 3575 2387
rect 3613 2353 3643 2387
rect 3643 2353 3647 2387
rect 3469 2280 3473 2314
rect 3473 2280 3503 2314
rect 3541 2280 3575 2314
rect 3613 2280 3643 2314
rect 3643 2280 3647 2314
rect 3469 2207 3473 2241
rect 3473 2207 3503 2241
rect 3541 2207 3575 2241
rect 3613 2207 3643 2241
rect 3643 2207 3647 2241
rect 3469 2134 3473 2168
rect 3473 2134 3503 2168
rect 3541 2134 3575 2168
rect 3613 2134 3643 2168
rect 3643 2134 3647 2168
rect 3469 2061 3473 2095
rect 3473 2061 3503 2095
rect 3541 2061 3575 2095
rect 3613 2061 3643 2095
rect 3643 2061 3647 2095
rect 3469 1988 3473 2022
rect 3473 1988 3503 2022
rect 3541 1988 3575 2022
rect 3613 1988 3643 2022
rect 3643 1988 3647 2022
rect 3469 1915 3473 1949
rect 3473 1915 3503 1949
rect 3541 1915 3575 1949
rect 3613 1915 3643 1949
rect 3643 1915 3647 1949
rect 3469 1842 3473 1876
rect 3473 1842 3503 1876
rect 3541 1842 3575 1876
rect 3613 1842 3643 1876
rect 3643 1842 3647 1876
rect 3469 1769 3473 1803
rect 3473 1769 3503 1803
rect 3541 1769 3575 1803
rect 3613 1769 3643 1803
rect 3643 1769 3647 1803
rect -24 403 -22 437
rect -22 403 10 437
rect 48 403 80 437
rect 80 403 82 437
rect -24 330 -22 364
rect -22 330 10 364
rect 48 330 80 364
rect 80 330 82 364
rect -24 257 -22 291
rect -22 257 10 291
rect 48 257 80 291
rect 80 257 82 291
rect 3469 218 3473 1730
rect -24 184 -22 218
rect -22 184 10 218
rect 48 182 80 218
rect 80 216 3473 218
rect 3473 216 3643 1730
rect 3643 218 3647 1730
rect 3810 2468 3844 2480
rect 3810 2446 3844 2468
rect 3810 2395 3844 2406
rect 3810 2372 3844 2395
rect 3810 2322 3844 2331
rect 3810 2297 3844 2322
rect 3810 2250 3844 2256
rect 3810 2222 3844 2250
rect 3810 2178 3844 2181
rect 3810 2147 3844 2178
rect 3810 2072 3844 2106
rect 3810 2000 3844 2031
rect 3810 1997 3844 2000
rect 3810 1928 3844 1956
rect 3810 1922 3844 1928
rect 3810 1856 3844 1881
rect 3810 1847 3844 1856
rect 3810 1784 3844 1806
rect 3810 1772 3844 1784
rect 3810 1712 3844 1731
rect 3810 1697 3844 1712
rect 3810 1640 3844 1656
rect 3810 1622 3844 1640
rect 3810 1568 3844 1581
rect 3810 1547 3844 1568
rect 3810 1496 3844 1506
rect 3810 1472 3844 1496
rect 4369 2468 4403 2480
rect 4369 2446 4403 2468
rect 4369 2395 4403 2406
rect 4369 2372 4403 2395
rect 4369 2322 4403 2331
rect 4369 2297 4403 2322
rect 4369 2250 4403 2256
rect 4369 2222 4403 2250
rect 4369 2178 4403 2181
rect 4369 2147 4403 2178
rect 4369 2072 4403 2106
rect 4369 2000 4403 2031
rect 4369 1997 4403 2000
rect 4369 1928 4403 1956
rect 4369 1922 4403 1928
rect 4369 1856 4403 1881
rect 4369 1847 4403 1856
rect 4369 1784 4403 1806
rect 4369 1772 4403 1784
rect 4369 1712 4403 1731
rect 4369 1697 4403 1712
rect 4369 1640 4403 1656
rect 4369 1622 4403 1640
rect 4369 1568 4403 1581
rect 4369 1547 4403 1568
rect 4369 1496 4403 1506
rect 4369 1472 4403 1496
rect 4592 2426 4596 2460
rect 4596 2426 4626 2460
rect 4664 2426 4698 2460
rect 4736 2426 4766 2460
rect 4766 2426 4770 2460
rect 4592 2353 4596 2387
rect 4596 2353 4626 2387
rect 4664 2353 4698 2387
rect 4736 2353 4766 2387
rect 4766 2353 4770 2387
rect 4592 2280 4596 2314
rect 4596 2280 4626 2314
rect 4664 2280 4698 2314
rect 4736 2280 4766 2314
rect 4766 2280 4770 2314
rect 4592 2207 4596 2241
rect 4596 2207 4626 2241
rect 4664 2207 4698 2241
rect 4736 2207 4766 2241
rect 4766 2207 4770 2241
rect 4592 2134 4596 2168
rect 4596 2134 4626 2168
rect 4664 2134 4698 2168
rect 4736 2134 4766 2168
rect 4766 2134 4770 2168
rect 4592 2061 4596 2095
rect 4596 2061 4626 2095
rect 4664 2061 4698 2095
rect 4736 2061 4766 2095
rect 4766 2061 4770 2095
rect 4592 1988 4596 2022
rect 4596 1988 4626 2022
rect 4664 1988 4698 2022
rect 4736 1988 4766 2022
rect 4766 1988 4770 2022
rect 4592 1915 4596 1949
rect 4596 1915 4626 1949
rect 4664 1915 4698 1949
rect 4736 1915 4766 1949
rect 4766 1915 4770 1949
rect 4592 1842 4596 1876
rect 4596 1842 4626 1876
rect 4664 1842 4698 1876
rect 4736 1842 4766 1876
rect 4766 1842 4770 1876
rect 4592 1769 4596 1803
rect 4596 1769 4626 1803
rect 4664 1769 4698 1803
rect 4736 1769 4766 1803
rect 4766 1769 4770 1803
rect 3938 1346 3972 1380
rect 4013 1346 4047 1380
rect 4088 1346 4122 1380
rect 4163 1346 4197 1380
rect 4238 1346 4272 1380
rect 3938 1274 3972 1308
rect 4013 1274 4047 1308
rect 4088 1274 4122 1308
rect 4163 1274 4197 1308
rect 4238 1274 4272 1308
rect 3911 506 3945 540
rect 3985 506 4019 540
rect 4059 506 4093 540
rect 4133 506 4167 540
rect 4207 506 4241 540
rect 4281 506 4315 540
rect 3911 434 3945 468
rect 3985 434 4019 468
rect 4059 434 4093 468
rect 4133 434 4167 468
rect 4207 434 4241 468
rect 4281 434 4315 468
rect 4592 218 4596 1730
rect 3643 216 4596 218
rect 4596 216 4766 1730
rect 4766 218 4770 1730
rect 5003 5448 5037 5449
rect 5076 5448 5110 5449
rect 5149 5448 5183 5449
rect 5222 5448 5256 5449
rect 5295 5448 6049 5449
rect 6125 5448 6159 5449
rect 6199 5448 6233 5449
rect 6272 5448 6306 5449
rect 6345 5448 6379 5449
rect 6418 5448 6452 5449
rect 6491 5448 6525 5449
rect 6564 5448 6598 5449
rect 6637 5448 6671 5449
rect 6710 5448 6744 5449
rect 6783 5448 6817 5449
rect 6856 5448 6890 5449
rect 6929 5448 6963 5449
rect 7002 5448 7036 5449
rect 7075 5448 7109 5449
rect 7148 5448 7182 5449
rect 7221 5448 7255 5449
rect 7294 5448 7328 5449
rect 7367 5448 7401 5449
rect 7440 5448 7474 5449
rect 7513 5448 7547 5449
rect 7586 5448 7620 5449
rect 7659 5448 7693 5449
rect 7732 5448 7766 5449
rect 7805 5448 7839 5449
rect 7878 5448 7912 5449
rect 7951 5448 7985 5449
rect 8024 5448 8058 5449
rect 8097 5448 8131 5449
rect 8170 5448 8204 5449
rect 8243 5448 8277 5449
rect 8316 5448 8350 5449
rect 8389 5448 8423 5449
rect 8462 5448 8496 5449
rect 8535 5448 8569 5449
rect 8608 5448 8642 5449
rect 8681 5448 8715 5449
rect 8754 5448 8788 5449
rect 8827 5448 8861 5449
rect 8900 5448 8934 5449
rect 8973 5448 9007 5449
rect 9046 5448 9080 5449
rect 9119 5448 9153 5449
rect 9192 5448 9226 5449
rect 9265 5448 9299 5449
rect 9338 5448 9372 5449
rect 9411 5448 9445 5449
rect 9484 5448 9518 5449
rect 9557 5448 9591 5449
rect 9630 5448 9664 5449
rect 9703 5448 9737 5449
rect 9776 5448 9810 5449
rect 9849 5448 9883 5449
rect 9922 5448 9956 5449
rect 5003 5415 5037 5448
rect 5076 5415 5110 5448
rect 5149 5415 5183 5448
rect 5222 5415 5256 5448
rect 4931 5346 5001 5377
rect 5001 5346 5037 5377
rect 5076 5346 5110 5377
rect 5149 5346 5183 5377
rect 5222 5346 5256 5377
rect 5295 5346 6049 5448
rect 6125 5415 6159 5448
rect 6199 5415 6233 5448
rect 6272 5415 6306 5448
rect 6345 5415 6379 5448
rect 6418 5415 6452 5448
rect 6491 5415 6525 5448
rect 6564 5415 6598 5448
rect 6637 5415 6671 5448
rect 6710 5415 6744 5448
rect 6783 5415 6817 5448
rect 6856 5415 6890 5448
rect 6929 5415 6963 5448
rect 7002 5415 7036 5448
rect 7075 5415 7109 5448
rect 7148 5415 7182 5448
rect 7221 5415 7255 5448
rect 7294 5415 7328 5448
rect 7367 5415 7401 5448
rect 7440 5415 7474 5448
rect 7513 5415 7547 5448
rect 7586 5415 7620 5448
rect 7659 5415 7693 5448
rect 7732 5415 7766 5448
rect 7805 5415 7839 5448
rect 7878 5415 7912 5448
rect 7951 5415 7985 5448
rect 8024 5415 8058 5448
rect 8097 5415 8131 5448
rect 8170 5415 8204 5448
rect 8243 5415 8277 5448
rect 8316 5415 8350 5448
rect 8389 5415 8423 5448
rect 8462 5415 8496 5448
rect 8535 5415 8569 5448
rect 8608 5415 8642 5448
rect 8681 5415 8715 5448
rect 8754 5415 8788 5448
rect 8827 5415 8861 5448
rect 8900 5415 8934 5448
rect 8973 5415 9007 5448
rect 9046 5415 9080 5448
rect 9119 5415 9153 5448
rect 9192 5415 9226 5448
rect 9265 5415 9299 5448
rect 9338 5415 9372 5448
rect 9411 5415 9445 5448
rect 9484 5415 9518 5448
rect 9557 5415 9591 5448
rect 9630 5415 9664 5448
rect 9703 5415 9737 5448
rect 9776 5415 9810 5448
rect 9849 5415 9863 5448
rect 9863 5415 9883 5448
rect 9922 5415 9931 5448
rect 9931 5415 9956 5448
rect 6125 5346 6159 5377
rect 6199 5346 6233 5377
rect 6272 5346 6306 5377
rect 6345 5346 6379 5377
rect 6418 5346 6452 5377
rect 6491 5346 6525 5377
rect 6564 5346 6598 5377
rect 6637 5346 6671 5377
rect 6710 5346 6744 5377
rect 6783 5346 6817 5377
rect 6856 5346 6890 5377
rect 6929 5346 6963 5377
rect 7002 5346 7036 5377
rect 7075 5346 7109 5377
rect 7148 5346 7182 5377
rect 7221 5346 7255 5377
rect 7294 5346 7328 5377
rect 7367 5346 7401 5377
rect 7440 5346 7474 5377
rect 7513 5346 7547 5377
rect 7586 5346 7620 5377
rect 7659 5346 7693 5377
rect 7732 5346 7766 5377
rect 7805 5346 7839 5377
rect 7878 5346 7912 5377
rect 7951 5346 7985 5377
rect 8024 5346 8058 5377
rect 8097 5346 8131 5377
rect 8170 5346 8204 5377
rect 8243 5346 8277 5377
rect 8316 5346 8350 5377
rect 8389 5346 8423 5377
rect 8462 5346 8496 5377
rect 8535 5346 8569 5377
rect 8608 5346 8642 5377
rect 8681 5346 8715 5377
rect 8754 5346 8788 5377
rect 8827 5346 8861 5377
rect 8900 5346 8934 5377
rect 8973 5346 9007 5377
rect 9046 5346 9080 5377
rect 9119 5346 9153 5377
rect 9192 5346 9226 5377
rect 9265 5346 9299 5377
rect 9338 5346 9372 5377
rect 9411 5346 9445 5377
rect 9484 5346 9518 5377
rect 9557 5346 9591 5377
rect 9630 5346 9664 5377
rect 9703 5346 9737 5377
rect 9776 5346 9810 5377
rect 9849 5346 9863 5377
rect 9863 5346 9883 5377
rect 4931 5342 5037 5346
rect 5076 5343 5110 5346
rect 5149 5343 5183 5346
rect 5222 5343 5256 5346
rect 5295 5343 6049 5346
rect 6125 5343 6159 5346
rect 6199 5343 6233 5346
rect 6272 5343 6306 5346
rect 6345 5343 6379 5346
rect 6418 5343 6452 5346
rect 6491 5343 6525 5346
rect 6564 5343 6598 5346
rect 6637 5343 6671 5346
rect 6710 5343 6744 5346
rect 6783 5343 6817 5346
rect 6856 5343 6890 5346
rect 6929 5343 6963 5346
rect 7002 5343 7036 5346
rect 7075 5343 7109 5346
rect 7148 5343 7182 5346
rect 7221 5343 7255 5346
rect 7294 5343 7328 5346
rect 7367 5343 7401 5346
rect 7440 5343 7474 5346
rect 7513 5343 7547 5346
rect 7586 5343 7620 5346
rect 7659 5343 7693 5346
rect 7732 5343 7766 5346
rect 7805 5343 7839 5346
rect 7878 5343 7912 5346
rect 7951 5343 7985 5346
rect 8024 5343 8058 5346
rect 8097 5343 8131 5346
rect 8170 5343 8204 5346
rect 8243 5343 8277 5346
rect 8316 5343 8350 5346
rect 8389 5343 8423 5346
rect 8462 5343 8496 5346
rect 8535 5343 8569 5346
rect 8608 5343 8642 5346
rect 8681 5343 8715 5346
rect 8754 5343 8788 5346
rect 8827 5343 8861 5346
rect 8900 5343 8934 5346
rect 8973 5343 9007 5346
rect 9046 5343 9080 5346
rect 9119 5343 9153 5346
rect 9192 5343 9226 5346
rect 9265 5343 9299 5346
rect 9338 5343 9372 5346
rect 9411 5343 9445 5346
rect 9484 5343 9518 5346
rect 9557 5343 9591 5346
rect 9630 5343 9664 5346
rect 9703 5343 9737 5346
rect 9776 5343 9810 5346
rect 9849 5343 9883 5346
rect 9923 5343 9925 5377
rect 9925 5343 9957 5377
rect 9995 5343 10027 5377
rect 10027 5343 10029 5377
rect 4931 5308 4933 5342
rect 4933 5308 4967 5342
rect 4967 5308 5037 5342
rect 4931 5274 5037 5308
rect 4931 3543 4933 5274
rect 4933 3543 5035 5274
rect 5035 3543 5037 5274
rect 4931 3470 4933 3504
rect 4933 3470 4965 3504
rect 5003 3470 5035 3504
rect 5035 3470 5037 3504
rect 4931 3397 4933 3431
rect 4933 3397 4965 3431
rect 5003 3397 5035 3431
rect 5035 3397 5037 3431
rect 4931 3324 4933 3358
rect 4933 3324 4965 3358
rect 5003 3324 5035 3358
rect 5035 3324 5037 3358
rect 4931 3251 4933 3285
rect 4933 3251 4965 3285
rect 5003 3251 5035 3285
rect 5035 3251 5037 3285
rect 9923 5270 9925 5304
rect 9925 5270 9957 5304
rect 9995 5270 10027 5304
rect 10027 5270 10029 5304
rect 9923 5197 9925 5231
rect 9925 5197 9957 5231
rect 9995 5197 10027 5231
rect 10027 5197 10029 5231
rect 9923 5124 9925 5158
rect 9925 5124 9957 5158
rect 9995 5124 10027 5158
rect 10027 5124 10029 5158
rect 9923 5051 9925 5085
rect 9925 5051 9957 5085
rect 9995 5051 10027 5085
rect 10027 5051 10029 5085
rect 9923 4978 9925 5012
rect 9925 4978 9957 5012
rect 9995 4978 10027 5012
rect 10027 4978 10029 5012
rect 9923 4905 9925 4939
rect 9925 4905 9957 4939
rect 9995 4905 10027 4939
rect 10027 4905 10029 4939
rect 9923 4832 9925 4866
rect 9925 4832 9957 4866
rect 9995 4832 10027 4866
rect 10027 4832 10029 4866
rect 9923 4759 9925 4793
rect 9925 4759 9957 4793
rect 9995 4759 10027 4793
rect 10027 4759 10029 4793
rect 9923 4686 9925 4720
rect 9925 4686 9957 4720
rect 9995 4686 10027 4720
rect 10027 4686 10029 4720
rect 9923 4613 9925 4647
rect 9925 4613 9957 4647
rect 9995 4613 10027 4647
rect 10027 4613 10029 4647
rect 9923 4540 9925 4574
rect 9925 4540 9957 4574
rect 9995 4540 10027 4574
rect 10027 4540 10029 4574
rect 9923 4467 9925 4501
rect 9925 4467 9957 4501
rect 9995 4467 10027 4501
rect 10027 4467 10029 4501
rect 9923 4394 9925 4428
rect 9925 4394 9957 4428
rect 9995 4394 10027 4428
rect 10027 4394 10029 4428
rect 9923 4321 9925 4355
rect 9925 4321 9957 4355
rect 9995 4321 10027 4355
rect 10027 4321 10029 4355
rect 9923 4248 9925 4282
rect 9925 4248 9957 4282
rect 9995 4248 10027 4282
rect 10027 4248 10029 4282
rect 9923 4175 9925 4209
rect 9925 4175 9957 4209
rect 9995 4175 10027 4209
rect 10027 4175 10029 4209
rect 9923 4102 9925 4136
rect 9925 4102 9957 4136
rect 9995 4102 10027 4136
rect 10027 4102 10029 4136
rect 9923 4029 9925 4063
rect 9925 4029 9957 4063
rect 9995 4029 10027 4063
rect 10027 4029 10029 4063
rect 9923 3956 9925 3990
rect 9925 3956 9957 3990
rect 9995 3956 10027 3990
rect 10027 3956 10029 3990
rect 9923 3883 9925 3917
rect 9925 3883 9957 3917
rect 9995 3883 10027 3917
rect 10027 3883 10029 3917
rect 9923 3810 9925 3844
rect 9925 3810 9957 3844
rect 9995 3810 10027 3844
rect 10027 3810 10029 3844
rect 9923 3737 9925 3771
rect 9925 3737 9957 3771
rect 9995 3737 10027 3771
rect 10027 3737 10029 3771
rect 9923 3664 9925 3698
rect 9925 3664 9957 3698
rect 9995 3664 10027 3698
rect 10027 3664 10029 3698
rect 9923 3591 9925 3625
rect 9925 3591 9957 3625
rect 9995 3591 10027 3625
rect 10027 3591 10029 3625
rect 9923 3518 9925 3552
rect 9925 3518 9957 3552
rect 9995 3518 10027 3552
rect 10027 3518 10029 3552
rect 9923 3445 9925 3479
rect 9925 3445 9957 3479
rect 9995 3445 10027 3479
rect 10027 3445 10029 3479
rect 9923 3372 9925 3406
rect 9925 3372 9957 3406
rect 9995 3372 10027 3406
rect 10027 3372 10029 3406
rect 9923 3299 9925 3333
rect 9925 3299 9957 3333
rect 9995 3299 10027 3333
rect 10027 3299 10029 3333
rect 9923 3226 9925 3260
rect 9925 3226 9957 3260
rect 9995 3226 10027 3260
rect 10027 3226 10029 3260
rect 4931 3178 4933 3212
rect 4933 3178 4965 3212
rect 5003 3178 5035 3212
rect 5035 3178 5037 3212
rect 5203 3182 5218 3216
rect 5218 3182 5237 3216
rect 5275 3182 5286 3216
rect 5286 3182 5309 3216
rect 5347 3182 5354 3216
rect 5354 3182 5381 3216
rect 5419 3182 5422 3216
rect 5422 3182 5453 3216
rect 5491 3182 5524 3216
rect 5524 3182 5525 3216
rect 5563 3182 5592 3216
rect 5592 3182 5597 3216
rect 5635 3182 5660 3216
rect 5660 3182 5669 3216
rect 5707 3182 5728 3216
rect 5728 3182 5741 3216
rect 5779 3182 5796 3216
rect 5796 3182 5813 3216
rect 5851 3182 5864 3216
rect 5864 3182 5885 3216
rect 5923 3182 5932 3216
rect 5932 3182 5957 3216
rect 5995 3182 6000 3216
rect 6000 3182 6029 3216
rect 6067 3182 6068 3216
rect 6068 3182 6101 3216
rect 6139 3182 6170 3216
rect 6170 3182 6173 3216
rect 6211 3182 6238 3216
rect 6238 3182 6245 3216
rect 6283 3182 6306 3216
rect 6306 3182 6317 3216
rect 6355 3182 6374 3216
rect 6374 3182 6389 3216
rect 6427 3182 6442 3216
rect 6442 3182 6461 3216
rect 6499 3182 6510 3216
rect 6510 3182 6533 3216
rect 6571 3182 6578 3216
rect 6578 3182 6605 3216
rect 6643 3182 6646 3216
rect 6646 3182 6677 3216
rect 6715 3182 6748 3216
rect 6748 3182 6749 3216
rect 6787 3182 6816 3216
rect 6816 3182 6821 3216
rect 6859 3182 6884 3216
rect 6884 3182 6893 3216
rect 6931 3182 6952 3216
rect 6952 3182 6965 3216
rect 7003 3182 7020 3216
rect 7020 3182 7037 3216
rect 7075 3182 7088 3216
rect 7088 3182 7109 3216
rect 7147 3182 7156 3216
rect 7156 3182 7181 3216
rect 7219 3182 7224 3216
rect 7224 3182 7253 3216
rect 7291 3182 7292 3216
rect 7292 3182 7325 3216
rect 7363 3182 7394 3216
rect 7394 3182 7397 3216
rect 7435 3182 7462 3216
rect 7462 3182 7469 3216
rect 7507 3182 7530 3216
rect 7530 3182 7541 3216
rect 7579 3182 7598 3216
rect 7598 3182 7613 3216
rect 7651 3182 7666 3216
rect 7666 3182 7685 3216
rect 7723 3182 7734 3216
rect 7734 3182 7757 3216
rect 7795 3182 7802 3216
rect 7802 3182 7829 3216
rect 7867 3182 7870 3216
rect 7870 3182 7901 3216
rect 7939 3182 7972 3216
rect 7972 3182 7973 3216
rect 8011 3182 8040 3216
rect 8040 3182 8045 3216
rect 8083 3182 8108 3216
rect 8108 3182 8117 3216
rect 8155 3182 8176 3216
rect 8176 3182 8189 3216
rect 8227 3182 8244 3216
rect 8244 3182 8261 3216
rect 8299 3182 8312 3216
rect 8312 3182 8333 3216
rect 8371 3182 8380 3216
rect 8380 3182 8405 3216
rect 8443 3182 8448 3216
rect 8448 3182 8477 3216
rect 8515 3182 8516 3216
rect 8516 3182 8549 3216
rect 8587 3182 8618 3216
rect 8618 3182 8621 3216
rect 8659 3182 8686 3216
rect 8686 3182 8693 3216
rect 8731 3182 8754 3216
rect 8754 3182 8765 3216
rect 8803 3182 8822 3216
rect 8822 3182 8837 3216
rect 8875 3182 8890 3216
rect 8890 3182 8909 3216
rect 8947 3182 8958 3216
rect 8958 3182 8981 3216
rect 9019 3182 9026 3216
rect 9026 3182 9053 3216
rect 9091 3182 9094 3216
rect 9094 3182 9125 3216
rect 9163 3182 9196 3216
rect 9196 3182 9197 3216
rect 9235 3182 9264 3216
rect 9264 3182 9269 3216
rect 9307 3182 9332 3216
rect 9332 3182 9341 3216
rect 9379 3182 9400 3216
rect 9400 3182 9413 3216
rect 9451 3182 9468 3216
rect 9468 3182 9485 3216
rect 9523 3182 9536 3216
rect 9536 3182 9557 3216
rect 9595 3182 9604 3216
rect 9604 3182 9629 3216
rect 9667 3182 9673 3216
rect 9673 3182 9701 3216
rect 9739 3182 9742 3216
rect 9742 3182 9773 3216
rect 4931 3105 4933 3139
rect 4933 3105 4965 3139
rect 5003 3105 5035 3139
rect 5035 3105 5037 3139
rect 4931 3032 4933 3066
rect 4933 3032 4965 3066
rect 5003 3032 5035 3066
rect 5035 3032 5037 3066
rect 9923 3153 9925 3187
rect 9925 3153 9957 3187
rect 9995 3153 10027 3187
rect 10027 3153 10029 3187
rect 9923 3080 9925 3114
rect 9925 3080 9957 3114
rect 9995 3080 10027 3114
rect 10027 3080 10029 3114
rect 5075 3012 5109 3014
rect 5148 3012 5182 3014
rect 5221 3012 5255 3014
rect 5294 3012 5328 3014
rect 5367 3012 5401 3014
rect 5440 3012 5474 3014
rect 5513 3012 5547 3014
rect 5586 3012 5620 3014
rect 5659 3012 5693 3014
rect 5732 3012 5766 3014
rect 5805 3012 5839 3014
rect 5878 3012 5912 3014
rect 5951 3012 5985 3014
rect 6024 3012 6058 3014
rect 6097 3012 6131 3014
rect 6170 3012 6204 3014
rect 6243 3012 6277 3014
rect 6316 3012 6350 3014
rect 6389 3012 6423 3014
rect 6462 3012 6496 3014
rect 6535 3012 6569 3014
rect 6608 3012 6642 3014
rect 6681 3012 6715 3014
rect 6754 3012 6788 3014
rect 6827 3012 9885 3014
rect 9923 3012 9925 3041
rect 9925 3012 9957 3041
rect 4931 2959 4933 2993
rect 4933 2959 4965 2993
rect 5003 2959 5035 2993
rect 5035 2959 5037 2993
rect 5075 2980 5097 3012
rect 5097 2980 5109 3012
rect 5148 2980 5182 3012
rect 5221 2980 5255 3012
rect 5294 2980 5328 3012
rect 5367 2980 5401 3012
rect 5440 2980 5474 3012
rect 5513 2980 5547 3012
rect 5586 2980 5620 3012
rect 5659 2980 5693 3012
rect 5732 2980 5766 3012
rect 5805 2980 5839 3012
rect 5878 2980 5912 3012
rect 5951 2980 5985 3012
rect 6024 2980 6058 3012
rect 6097 2980 6131 3012
rect 6170 2980 6204 3012
rect 6243 2980 6277 3012
rect 6316 2980 6350 3012
rect 6389 2980 6423 3012
rect 6462 2980 6496 3012
rect 6535 2980 6569 3012
rect 6608 2980 6642 3012
rect 6681 2980 6715 3012
rect 6754 2980 6788 3012
rect 4931 2886 4933 2920
rect 4933 2886 4965 2920
rect 5003 2886 5035 2920
rect 5035 2886 5037 2920
rect 5075 2910 5097 2942
rect 5097 2910 5109 2942
rect 5148 2910 5182 2942
rect 5221 2910 5255 2942
rect 5294 2910 5328 2942
rect 5367 2910 5401 2942
rect 5440 2910 5474 2942
rect 5513 2910 5547 2942
rect 5586 2910 5620 2942
rect 5659 2910 5693 2942
rect 5732 2910 5766 2942
rect 5805 2910 5839 2942
rect 5878 2910 5912 2942
rect 5951 2910 5985 2942
rect 6024 2910 6058 2942
rect 6097 2910 6131 2942
rect 6170 2910 6204 2942
rect 6243 2910 6277 2942
rect 6316 2910 6350 2942
rect 6389 2910 6423 2942
rect 6462 2910 6496 2942
rect 6535 2910 6569 2942
rect 6608 2910 6642 2942
rect 6681 2910 6715 2942
rect 6754 2910 6788 2942
rect 6827 2910 9885 3012
rect 9923 3007 9957 3012
rect 9995 3007 10027 3041
rect 10027 3007 10029 3041
rect 9923 2966 9957 2968
rect 9995 2966 10027 2968
rect 10027 2966 10029 2968
rect 9923 2934 9957 2966
rect 9995 2934 10029 2966
rect 5075 2908 5109 2910
rect 5148 2908 5182 2910
rect 5221 2908 5255 2910
rect 5294 2908 5328 2910
rect 5367 2908 5401 2910
rect 5440 2908 5474 2910
rect 5513 2908 5547 2910
rect 5586 2908 5620 2910
rect 5659 2908 5693 2910
rect 5732 2908 5766 2910
rect 5805 2908 5839 2910
rect 5878 2908 5912 2910
rect 5951 2908 5985 2910
rect 6024 2908 6058 2910
rect 6097 2908 6131 2910
rect 6170 2908 6204 2910
rect 6243 2908 6277 2910
rect 6316 2908 6350 2910
rect 6389 2908 6423 2910
rect 6462 2908 6496 2910
rect 6535 2908 6569 2910
rect 6608 2908 6642 2910
rect 6681 2908 6715 2910
rect 6754 2908 6788 2910
rect 6827 2908 9885 2910
rect 4931 2813 4933 2847
rect 4933 2813 4965 2847
rect 5003 2813 5035 2847
rect 5035 2813 5037 2847
rect 4931 2740 4933 2774
rect 4933 2740 4965 2774
rect 5003 2740 5035 2774
rect 5035 2740 5037 2774
rect 9923 2861 9957 2895
rect 9995 2861 10029 2895
rect 9923 2788 9925 2822
rect 9925 2788 9957 2822
rect 9995 2788 10027 2822
rect 10027 2788 10029 2822
rect 5203 2712 5218 2746
rect 5218 2712 5237 2746
rect 5275 2712 5286 2746
rect 5286 2712 5309 2746
rect 5347 2712 5354 2746
rect 5354 2712 5381 2746
rect 5419 2712 5422 2746
rect 5422 2712 5453 2746
rect 5491 2712 5524 2746
rect 5524 2712 5525 2746
rect 5563 2712 5592 2746
rect 5592 2712 5597 2746
rect 5635 2712 5660 2746
rect 5660 2712 5669 2746
rect 5707 2712 5728 2746
rect 5728 2712 5741 2746
rect 5779 2712 5796 2746
rect 5796 2712 5813 2746
rect 5851 2712 5864 2746
rect 5864 2712 5885 2746
rect 5923 2712 5932 2746
rect 5932 2712 5957 2746
rect 5995 2712 6000 2746
rect 6000 2712 6029 2746
rect 6067 2712 6068 2746
rect 6068 2712 6101 2746
rect 6139 2712 6170 2746
rect 6170 2712 6173 2746
rect 6211 2712 6238 2746
rect 6238 2712 6245 2746
rect 6283 2712 6306 2746
rect 6306 2712 6317 2746
rect 6355 2712 6374 2746
rect 6374 2712 6389 2746
rect 6427 2712 6442 2746
rect 6442 2712 6461 2746
rect 6499 2712 6510 2746
rect 6510 2712 6533 2746
rect 6571 2712 6578 2746
rect 6578 2712 6605 2746
rect 6643 2712 6646 2746
rect 6646 2712 6677 2746
rect 6715 2712 6748 2746
rect 6748 2712 6749 2746
rect 6787 2712 6816 2746
rect 6816 2712 6821 2746
rect 6859 2712 6884 2746
rect 6884 2712 6893 2746
rect 6931 2712 6952 2746
rect 6952 2712 6965 2746
rect 7003 2712 7020 2746
rect 7020 2712 7037 2746
rect 7075 2712 7088 2746
rect 7088 2712 7109 2746
rect 7147 2712 7156 2746
rect 7156 2712 7181 2746
rect 7219 2712 7224 2746
rect 7224 2712 7253 2746
rect 7291 2712 7292 2746
rect 7292 2712 7325 2746
rect 7363 2712 7394 2746
rect 7394 2712 7397 2746
rect 7435 2712 7462 2746
rect 7462 2712 7469 2746
rect 7507 2712 7530 2746
rect 7530 2712 7541 2746
rect 7579 2712 7598 2746
rect 7598 2712 7613 2746
rect 7651 2712 7666 2746
rect 7666 2712 7685 2746
rect 7723 2712 7734 2746
rect 7734 2712 7757 2746
rect 7795 2712 7802 2746
rect 7802 2712 7829 2746
rect 7867 2712 7870 2746
rect 7870 2712 7901 2746
rect 7939 2712 7972 2746
rect 7972 2712 7973 2746
rect 8011 2712 8040 2746
rect 8040 2712 8045 2746
rect 8083 2712 8108 2746
rect 8108 2712 8117 2746
rect 8155 2712 8176 2746
rect 8176 2712 8189 2746
rect 8227 2712 8244 2746
rect 8244 2712 8261 2746
rect 8299 2712 8312 2746
rect 8312 2712 8333 2746
rect 8371 2712 8380 2746
rect 8380 2712 8405 2746
rect 8443 2712 8448 2746
rect 8448 2712 8477 2746
rect 8515 2712 8516 2746
rect 8516 2712 8549 2746
rect 8587 2712 8618 2746
rect 8618 2712 8621 2746
rect 8659 2712 8686 2746
rect 8686 2712 8693 2746
rect 8731 2712 8754 2746
rect 8754 2712 8765 2746
rect 8803 2712 8822 2746
rect 8822 2712 8837 2746
rect 8875 2712 8890 2746
rect 8890 2712 8909 2746
rect 8947 2712 8958 2746
rect 8958 2712 8981 2746
rect 9019 2712 9026 2746
rect 9026 2712 9053 2746
rect 9091 2712 9094 2746
rect 9094 2712 9125 2746
rect 9163 2712 9196 2746
rect 9196 2712 9197 2746
rect 9235 2712 9264 2746
rect 9264 2712 9269 2746
rect 9307 2712 9332 2746
rect 9332 2712 9341 2746
rect 9379 2712 9400 2746
rect 9400 2712 9413 2746
rect 9451 2712 9468 2746
rect 9468 2712 9485 2746
rect 9523 2712 9536 2746
rect 9536 2712 9557 2746
rect 9595 2712 9604 2746
rect 9604 2712 9629 2746
rect 9667 2712 9673 2746
rect 9673 2712 9701 2746
rect 9739 2712 9742 2746
rect 9742 2712 9773 2746
rect 9923 2715 9925 2749
rect 9925 2715 9957 2749
rect 9995 2715 10027 2749
rect 10027 2715 10029 2749
rect 4931 2667 4933 2701
rect 4933 2667 4965 2701
rect 5003 2667 5035 2701
rect 5035 2667 5037 2701
rect 4931 2594 4933 2628
rect 4933 2594 4965 2628
rect 5003 2594 5035 2628
rect 5035 2594 5037 2628
rect 4931 2521 4933 2555
rect 4933 2521 4965 2555
rect 5003 2521 5035 2555
rect 5035 2521 5037 2555
rect 4931 2448 4933 2482
rect 4933 2448 4965 2482
rect 5003 2448 5035 2482
rect 5035 2448 5037 2482
rect 4931 2375 4933 2409
rect 4933 2375 4965 2409
rect 5003 2375 5035 2409
rect 5035 2375 5037 2409
rect 4931 2302 4933 2336
rect 4933 2302 4965 2336
rect 5003 2302 5035 2336
rect 5035 2302 5037 2336
rect 4931 2229 4933 2263
rect 4933 2229 4965 2263
rect 5003 2229 5035 2263
rect 5035 2229 5037 2263
rect 4931 2156 4933 2190
rect 4933 2156 4965 2190
rect 5003 2156 5035 2190
rect 5035 2156 5037 2190
rect 4931 2083 4933 2117
rect 4933 2083 4965 2117
rect 5003 2083 5035 2117
rect 5035 2083 5037 2117
rect 4931 2010 4933 2044
rect 4933 2010 4965 2044
rect 5003 2010 5035 2044
rect 5035 2010 5037 2044
rect 4931 1937 4933 1971
rect 4933 1937 4965 1971
rect 5003 1937 5035 1971
rect 5035 1937 5037 1971
rect 4931 1864 4933 1898
rect 4933 1864 4965 1898
rect 5003 1864 5035 1898
rect 5035 1864 5037 1898
rect 4931 1791 4933 1825
rect 4933 1791 4965 1825
rect 5003 1791 5035 1825
rect 5035 1791 5037 1825
rect 4931 1718 4933 1752
rect 4933 1718 4965 1752
rect 5003 1718 5035 1752
rect 5035 1718 5037 1752
rect 4931 1645 4933 1679
rect 4933 1645 4965 1679
rect 5003 1645 5035 1679
rect 5035 1645 5037 1679
rect 4931 1572 4933 1606
rect 4933 1572 4965 1606
rect 5003 1572 5035 1606
rect 5035 1572 5037 1606
rect 4931 1499 4933 1533
rect 4933 1499 4965 1533
rect 5003 1499 5035 1533
rect 5035 1499 5037 1533
rect 4931 1426 4933 1460
rect 4933 1426 4965 1460
rect 5003 1426 5035 1460
rect 5035 1426 5037 1460
rect 4931 1353 4933 1387
rect 4933 1353 4965 1387
rect 5003 1353 5035 1387
rect 5035 1353 5037 1387
rect 4931 1280 4933 1314
rect 4933 1280 4965 1314
rect 5003 1280 5035 1314
rect 5035 1280 5037 1314
rect 4931 1207 4933 1241
rect 4933 1207 4965 1241
rect 5003 1207 5035 1241
rect 5035 1207 5037 1241
rect 4931 1134 4933 1168
rect 4933 1134 4965 1168
rect 5003 1134 5035 1168
rect 5035 1134 5037 1168
rect 4931 1061 4933 1095
rect 4933 1061 4965 1095
rect 5003 1061 5035 1095
rect 5035 1061 5037 1095
rect 4931 988 4933 1022
rect 4933 988 4965 1022
rect 5003 988 5035 1022
rect 5035 988 5037 1022
rect 4931 915 4933 949
rect 4933 915 4965 949
rect 5003 915 5035 949
rect 5035 915 5037 949
rect 4931 842 4933 876
rect 4933 842 4965 876
rect 5003 842 5035 876
rect 5035 842 5037 876
rect 4931 769 4933 803
rect 4933 769 4965 803
rect 5003 769 5035 803
rect 5035 769 5037 803
rect 4931 696 4933 730
rect 4933 696 4965 730
rect 5003 696 5035 730
rect 5035 696 5037 730
rect 4931 623 4933 657
rect 4933 623 4965 657
rect 5003 623 5035 657
rect 5035 623 5037 657
rect 9923 2642 9925 2676
rect 9925 2642 9957 2676
rect 9995 2642 10027 2676
rect 10027 2642 10029 2676
rect 9923 2569 9925 2603
rect 9925 2569 9957 2603
rect 9995 2569 10027 2603
rect 10027 2569 10029 2603
rect 9923 2496 9925 2530
rect 9925 2496 9957 2530
rect 9995 2496 10027 2530
rect 10027 2496 10029 2530
rect 9923 2423 9925 2457
rect 9925 2423 9957 2457
rect 9995 2423 10027 2457
rect 10027 2423 10029 2457
rect 9923 628 9925 2384
rect 9925 628 10027 2384
rect 10027 628 10029 2384
rect 9923 594 10029 628
rect 4931 550 4933 584
rect 4933 550 4965 584
rect 5003 548 5035 584
rect 5035 582 8205 584
rect 8244 582 8278 584
rect 8317 582 8351 584
rect 8390 582 8424 584
rect 8463 582 8497 584
rect 8536 582 8570 584
rect 8609 582 8643 584
rect 8682 582 8716 584
rect 8755 582 8789 584
rect 8828 582 8862 584
rect 8901 582 8935 584
rect 8974 582 9008 584
rect 9047 582 9081 584
rect 9120 582 9154 584
rect 9193 582 9227 584
rect 9266 582 9300 584
rect 9339 582 9373 584
rect 9412 582 9446 584
rect 9485 582 9519 584
rect 9558 582 9592 584
rect 9631 582 9665 584
rect 9704 582 9738 584
rect 9777 582 9811 584
rect 9850 582 9884 584
rect 9923 582 9993 594
rect 5035 548 5097 582
rect 5003 514 5097 548
rect 5003 480 5029 514
rect 5029 480 5063 514
rect 5063 480 5097 514
rect 5097 480 8205 582
rect 8244 550 8278 582
rect 8317 550 8351 582
rect 8390 550 8424 582
rect 8463 550 8497 582
rect 8536 550 8570 582
rect 8609 550 8643 582
rect 8682 550 8716 582
rect 8755 550 8789 582
rect 8828 550 8862 582
rect 8901 550 8935 582
rect 8974 550 9008 582
rect 9047 550 9081 582
rect 9120 550 9154 582
rect 9193 550 9227 582
rect 9266 550 9300 582
rect 9339 550 9373 582
rect 9412 550 9446 582
rect 9485 550 9519 582
rect 9558 550 9592 582
rect 9631 550 9665 582
rect 9704 550 9738 582
rect 9777 550 9811 582
rect 9850 550 9884 582
rect 9923 550 9959 582
rect 9959 560 9993 582
rect 9993 560 10027 594
rect 10027 560 10029 594
rect 9959 550 10029 560
rect 8244 480 8278 512
rect 8317 480 8351 512
rect 8390 480 8424 512
rect 8463 480 8497 512
rect 8536 480 8570 512
rect 8609 480 8643 512
rect 8682 480 8716 512
rect 8755 480 8789 512
rect 8828 480 8862 512
rect 8901 480 8935 512
rect 8974 480 9008 512
rect 9047 480 9081 512
rect 9120 480 9154 512
rect 9193 480 9227 512
rect 9266 480 9300 512
rect 9339 480 9373 512
rect 9412 480 9446 512
rect 9485 480 9519 512
rect 9558 480 9592 512
rect 9631 480 9665 512
rect 9704 480 9738 512
rect 9777 480 9811 512
rect 9850 480 9884 512
rect 9923 480 9957 512
rect 5003 478 8205 480
rect 8244 478 8278 480
rect 8317 478 8351 480
rect 8390 478 8424 480
rect 8463 478 8497 480
rect 8536 478 8570 480
rect 8609 478 8643 480
rect 8682 478 8716 480
rect 8755 478 8789 480
rect 8828 478 8862 480
rect 8901 478 8935 480
rect 8974 478 9008 480
rect 9047 478 9081 480
rect 9120 478 9154 480
rect 9193 478 9227 480
rect 9266 478 9300 480
rect 9339 478 9373 480
rect 9412 478 9446 480
rect 9485 478 9519 480
rect 9558 478 9592 480
rect 9631 478 9665 480
rect 9704 478 9738 480
rect 9777 478 9811 480
rect 9850 478 9884 480
rect 9923 478 9957 480
rect 10277 5418 10279 5452
rect 10279 5418 10311 5452
rect 10349 5418 10381 5452
rect 10381 5418 10383 5452
rect 10277 5345 10279 5379
rect 10279 5345 10311 5379
rect 10349 5345 10381 5379
rect 10381 5345 10383 5379
rect 10277 5272 10279 5306
rect 10279 5272 10311 5306
rect 10349 5272 10381 5306
rect 10381 5272 10383 5306
rect 10277 5199 10279 5233
rect 10279 5199 10311 5233
rect 10349 5199 10381 5233
rect 10381 5199 10383 5233
rect 10277 5126 10279 5160
rect 10279 5126 10311 5160
rect 10349 5126 10381 5160
rect 10381 5126 10383 5160
rect 10277 5053 10279 5087
rect 10279 5053 10311 5087
rect 10349 5053 10381 5087
rect 10381 5053 10383 5087
rect 10277 4980 10279 5014
rect 10279 4980 10311 5014
rect 10349 4980 10381 5014
rect 10381 4980 10383 5014
rect 10277 4907 10279 4941
rect 10279 4907 10311 4941
rect 10349 4907 10381 4941
rect 10381 4907 10383 4941
rect 10277 4834 10279 4868
rect 10279 4834 10311 4868
rect 10349 4834 10381 4868
rect 10381 4834 10383 4868
rect 10277 4761 10279 4795
rect 10279 4761 10311 4795
rect 10349 4761 10381 4795
rect 10381 4761 10383 4795
rect 10277 4688 10279 4722
rect 10279 4688 10311 4722
rect 10349 4688 10381 4722
rect 10381 4688 10383 4722
rect 10277 4615 10279 4649
rect 10279 4615 10311 4649
rect 10349 4615 10381 4649
rect 10381 4615 10383 4649
rect 10277 4542 10279 4576
rect 10279 4542 10311 4576
rect 10349 4542 10381 4576
rect 10381 4542 10383 4576
rect 10277 4469 10279 4503
rect 10279 4469 10311 4503
rect 10349 4469 10381 4503
rect 10381 4469 10383 4503
rect 10277 4396 10279 4430
rect 10279 4396 10311 4430
rect 10349 4396 10381 4430
rect 10381 4396 10383 4430
rect 10277 4323 10279 4357
rect 10279 4323 10311 4357
rect 10349 4323 10381 4357
rect 10381 4323 10383 4357
rect 10277 4250 10279 4284
rect 10279 4250 10311 4284
rect 10349 4250 10381 4284
rect 10381 4250 10383 4284
rect 10277 4177 10279 4211
rect 10279 4177 10311 4211
rect 10349 4177 10381 4211
rect 10381 4177 10383 4211
rect 10277 4104 10279 4138
rect 10279 4104 10311 4138
rect 10349 4104 10381 4138
rect 10381 4104 10383 4138
rect 10277 4031 10279 4065
rect 10279 4031 10311 4065
rect 10349 4031 10381 4065
rect 10381 4031 10383 4065
rect 10277 3958 10279 3992
rect 10279 3958 10311 3992
rect 10349 3958 10381 3992
rect 10381 3958 10383 3992
rect 10277 3885 10279 3919
rect 10279 3885 10311 3919
rect 10349 3885 10381 3919
rect 10381 3885 10383 3919
rect 10277 3812 10279 3846
rect 10279 3812 10311 3846
rect 10349 3812 10381 3846
rect 10381 3812 10383 3846
rect 10277 3739 10279 3773
rect 10279 3739 10311 3773
rect 10349 3739 10381 3773
rect 10381 3739 10383 3773
rect 10277 3666 10279 3700
rect 10279 3666 10311 3700
rect 10349 3666 10381 3700
rect 10381 3666 10383 3700
rect 10277 3593 10279 3627
rect 10279 3593 10311 3627
rect 10349 3593 10381 3627
rect 10381 3593 10383 3627
rect 10277 3520 10279 3554
rect 10279 3520 10311 3554
rect 10349 3520 10381 3554
rect 10381 3520 10383 3554
rect 10277 3447 10279 3481
rect 10279 3447 10311 3481
rect 10349 3447 10381 3481
rect 10381 3447 10383 3481
rect 10277 3374 10279 3408
rect 10279 3374 10311 3408
rect 10349 3374 10381 3408
rect 10381 3374 10383 3408
rect 10277 3301 10279 3335
rect 10279 3301 10311 3335
rect 10349 3301 10381 3335
rect 10381 3301 10383 3335
rect 10277 3228 10279 3262
rect 10279 3228 10311 3262
rect 10349 3228 10381 3262
rect 10381 3228 10383 3262
rect 10277 3155 10279 3189
rect 10279 3155 10311 3189
rect 10349 3155 10381 3189
rect 10381 3155 10383 3189
rect 10277 3082 10279 3116
rect 10279 3082 10311 3116
rect 10349 3082 10381 3116
rect 10381 3082 10383 3116
rect 10277 3009 10279 3043
rect 10279 3009 10311 3043
rect 10349 3009 10381 3043
rect 10381 3009 10383 3043
rect 10277 2936 10279 2970
rect 10279 2936 10311 2970
rect 10349 2936 10381 2970
rect 10381 2936 10383 2970
rect 10277 2863 10279 2897
rect 10279 2863 10311 2897
rect 10349 2863 10381 2897
rect 10381 2863 10383 2897
rect 10277 2790 10279 2824
rect 10279 2790 10311 2824
rect 10349 2790 10381 2824
rect 10381 2790 10383 2824
rect 10277 2717 10279 2751
rect 10279 2717 10311 2751
rect 10349 2717 10381 2751
rect 10381 2717 10383 2751
rect 10277 2644 10279 2678
rect 10279 2644 10311 2678
rect 10349 2644 10381 2678
rect 10381 2644 10383 2678
rect 10277 2571 10279 2605
rect 10279 2571 10311 2605
rect 10349 2571 10381 2605
rect 10381 2571 10383 2605
rect 10277 2498 10279 2532
rect 10279 2498 10311 2532
rect 10349 2498 10381 2532
rect 10381 2498 10383 2532
rect 10277 2425 10279 2459
rect 10279 2425 10311 2459
rect 10349 2425 10381 2459
rect 10381 2425 10383 2459
rect 10277 2352 10279 2386
rect 10279 2352 10311 2386
rect 10349 2352 10381 2386
rect 10381 2352 10383 2386
rect 10277 2279 10279 2313
rect 10279 2279 10311 2313
rect 10349 2279 10381 2313
rect 10381 2279 10383 2313
rect 10277 2206 10279 2240
rect 10279 2206 10311 2240
rect 10349 2206 10381 2240
rect 10381 2206 10383 2240
rect 10277 2133 10279 2167
rect 10279 2133 10311 2167
rect 10349 2133 10381 2167
rect 10381 2133 10383 2167
rect 10277 2060 10279 2094
rect 10279 2060 10311 2094
rect 10349 2060 10381 2094
rect 10381 2060 10383 2094
rect 10277 1987 10279 2021
rect 10279 1987 10311 2021
rect 10349 1987 10381 2021
rect 10381 1987 10383 2021
rect 10277 1914 10279 1948
rect 10279 1914 10311 1948
rect 10349 1914 10381 1948
rect 10381 1914 10383 1948
rect 10277 1841 10279 1875
rect 10279 1841 10311 1875
rect 10349 1841 10381 1875
rect 10381 1841 10383 1875
rect 10277 1496 10279 1802
rect 10279 1496 10381 1802
rect 10381 1496 10383 1802
rect 10277 1376 10383 1496
rect 10277 254 10279 1376
rect 10279 254 10381 1376
rect 10381 254 10383 1376
rect 10277 220 10383 254
rect 4766 216 9946 218
rect 9985 216 10019 218
rect 10058 216 10092 218
rect 10131 216 10165 218
rect 10204 216 10238 218
rect 10277 216 10347 220
rect 80 182 147 216
rect 48 148 147 182
rect 48 114 79 148
rect 79 114 113 148
rect 113 114 147 148
rect 147 114 9946 216
rect 9985 184 10019 216
rect 10058 184 10092 216
rect 10131 184 10165 216
rect 10204 184 10238 216
rect 10277 184 10313 216
rect 10313 186 10347 216
rect 10347 186 10381 220
rect 10381 186 10383 220
rect 10313 184 10383 186
rect 9985 114 10019 146
rect 10058 114 10092 146
rect 10131 114 10165 146
rect 10204 114 10238 146
rect 10277 114 10311 146
rect 48 112 9946 114
rect 9985 112 10019 114
rect 10058 112 10092 114
rect 10131 112 10165 114
rect 10204 112 10238 114
rect 10277 112 10311 114
<< metal1 >>
rect -30 5770 -16 5822
rect 36 5770 48 5822
rect 100 5770 112 5822
rect 164 5770 176 5822
rect 228 5770 240 5822
rect 292 5816 304 5822
rect 356 5816 368 5822
rect 420 5816 432 5822
rect 484 5816 496 5822
rect 548 5816 560 5822
rect 301 5782 304 5816
rect 484 5782 486 5816
rect 548 5782 559 5816
rect 292 5770 304 5782
rect 356 5770 368 5782
rect 420 5770 432 5782
rect 484 5770 496 5782
rect 548 5770 560 5782
rect 612 5770 624 5822
rect 676 5770 688 5822
rect 740 5770 752 5822
rect 804 5816 816 5822
rect 868 5816 880 5822
rect 932 5816 944 5822
rect 996 5816 1008 5822
rect 1060 5816 1072 5822
rect 812 5782 816 5816
rect 996 5782 997 5816
rect 1060 5782 1070 5816
rect 804 5770 816 5782
rect 868 5770 880 5782
rect 932 5770 944 5782
rect 996 5770 1008 5782
rect 1060 5770 1072 5782
rect 1124 5770 1136 5822
rect 1188 5770 1200 5822
rect 1252 5816 1264 5822
rect 1316 5816 1328 5822
rect 1380 5816 1392 5822
rect 1444 5816 1456 5822
rect 1508 5816 1520 5822
rect 1572 5816 1584 5822
rect 1636 5816 1648 5822
rect 1700 5816 1712 5822
rect 1764 5816 1776 5822
rect 1828 5816 1840 5822
rect 1892 5816 1904 5822
rect 1956 5816 1968 5822
rect 2020 5816 2032 5822
rect 2084 5816 2096 5822
rect 2148 5816 2160 5822
rect 2212 5816 2224 5822
rect 2276 5816 2288 5822
rect 2340 5816 2352 5822
rect 2404 5816 2416 5822
rect 2468 5816 2480 5822
rect 2532 5816 2544 5822
rect 2596 5816 2608 5822
rect 2660 5816 2672 5822
rect 2724 5816 2736 5822
rect 2788 5816 2800 5822
rect 2852 5816 2864 5822
rect 2916 5816 2928 5822
rect 2980 5816 2992 5822
rect 3044 5816 3056 5822
rect 3108 5816 3120 5822
rect 3172 5816 3184 5822
rect 3236 5816 3248 5822
rect 3300 5816 3312 5822
rect 3364 5816 3376 5822
rect 3428 5816 3440 5822
rect 3492 5816 3504 5822
rect 3556 5816 3568 5822
rect 3620 5816 3632 5822
rect 3684 5816 3696 5822
rect 3748 5816 3760 5822
rect 3812 5816 3824 5822
rect 3876 5816 3888 5822
rect 3940 5816 3952 5822
rect 4004 5816 4016 5822
rect 4068 5816 4080 5822
rect 4132 5816 4144 5822
rect 4196 5816 4208 5822
rect 4260 5816 4272 5822
rect 4324 5816 4336 5822
rect 4388 5816 4400 5822
rect 4452 5816 4464 5822
rect 4516 5816 4528 5822
rect 4580 5816 4592 5822
rect 4644 5816 4656 5822
rect 4708 5816 4720 5822
rect 4772 5816 4784 5822
rect 4836 5816 4848 5822
rect 4900 5816 4912 5822
rect 4964 5816 4976 5822
rect 5028 5816 5040 5822
rect 5092 5816 5104 5822
rect 5156 5816 5168 5822
rect 5220 5816 5232 5822
rect 5284 5816 5296 5822
rect 5348 5816 5360 5822
rect 5412 5816 5424 5822
rect 5476 5816 5488 5822
rect 5540 5816 5552 5822
rect 5604 5816 5616 5822
rect 5668 5816 5680 5822
rect 5732 5816 5744 5822
rect 5796 5816 5808 5822
rect 5860 5816 5872 5822
rect 5924 5816 5936 5822
rect 5988 5816 6000 5822
rect 6052 5816 6064 5822
rect 6116 5816 6128 5822
rect 6180 5816 6192 5822
rect 6244 5816 6256 5822
rect 6308 5816 6320 5822
rect 6372 5816 6384 5822
rect 6436 5816 6448 5822
rect 6500 5816 6512 5822
rect 6564 5816 6576 5822
rect 6628 5816 6640 5822
rect 6692 5816 6704 5822
rect 6756 5816 6768 5822
rect 6820 5816 6832 5822
rect 6884 5816 6896 5822
rect 6948 5816 6960 5822
rect 7012 5816 7024 5822
rect 7076 5816 7088 5822
rect 7140 5816 7152 5822
rect 7204 5816 7216 5822
rect 7268 5816 7280 5822
rect 7332 5816 7344 5822
rect 7396 5816 7408 5822
rect 7460 5816 7472 5822
rect 7524 5816 7536 5822
rect 7588 5816 7600 5822
rect 7652 5816 7664 5822
rect 7716 5816 7728 5822
rect 7780 5816 7792 5822
rect 7844 5816 7856 5822
rect 7908 5816 7920 5822
rect 7972 5816 7984 5822
rect 8036 5816 8048 5822
rect 8100 5816 8112 5822
rect 8164 5816 8176 5822
rect 8228 5816 8240 5822
rect 8292 5816 8304 5822
rect 8356 5816 8368 5822
rect 8420 5816 8432 5822
rect 8484 5816 8496 5822
rect 8548 5816 8560 5822
rect 8612 5816 8624 5822
rect 8676 5816 8688 5822
rect 8740 5816 8752 5822
rect 8804 5816 8816 5822
rect 8868 5816 8880 5822
rect 8932 5816 8944 5822
rect 8996 5816 9008 5822
rect 9060 5816 9072 5822
rect 9124 5816 9136 5822
rect 9188 5816 9200 5822
rect 9252 5816 9264 5822
rect 9316 5816 9329 5822
rect 9381 5816 9394 5822
rect 9446 5816 9459 5822
rect 9458 5770 9459 5816
rect 9511 5770 9524 5822
rect 9576 5770 9589 5822
rect 9641 5816 9654 5822
rect 9706 5816 9719 5822
rect 9771 5816 9784 5822
rect 9836 5816 9849 5822
rect 9901 5816 9914 5822
rect 9643 5782 9654 5816
rect 9717 5782 9719 5816
rect 9901 5782 9905 5816
rect 9641 5770 9654 5782
rect 9706 5770 9719 5782
rect 9771 5770 9784 5782
rect 9836 5770 9849 5782
rect 9901 5770 9914 5782
rect 9966 5770 9979 5822
rect 10031 5770 10044 5822
rect 10096 5770 10109 5822
rect 10161 5770 10174 5822
rect 10226 5816 10239 5822
rect 10291 5816 10389 5822
rect 10235 5782 10239 5816
rect 10309 5782 10389 5816
rect 10226 5770 10239 5782
rect 10291 5770 10389 5782
rect -30 5756 1216 5770
rect 9458 5756 10389 5770
rect -30 5744 -16 5756
rect 36 5744 48 5756
rect -30 4126 -24 5744
rect 100 5704 112 5756
rect 164 5704 176 5756
rect 228 5704 240 5756
rect 292 5744 304 5756
rect 356 5744 368 5756
rect 420 5744 432 5756
rect 484 5744 496 5756
rect 548 5744 560 5756
rect 301 5710 304 5744
rect 484 5710 486 5744
rect 548 5710 559 5744
rect 292 5704 304 5710
rect 356 5704 368 5710
rect 420 5704 432 5710
rect 484 5704 496 5710
rect 548 5704 560 5710
rect 612 5704 624 5756
rect 676 5704 688 5756
rect 740 5704 752 5756
rect 804 5744 816 5756
rect 868 5744 880 5756
rect 932 5744 944 5756
rect 996 5744 1008 5756
rect 1060 5744 1072 5756
rect 812 5710 816 5744
rect 996 5710 997 5744
rect 1060 5710 1070 5744
rect 804 5704 816 5710
rect 868 5704 880 5710
rect 932 5704 944 5710
rect 996 5704 1008 5710
rect 1060 5704 1072 5710
rect 1124 5704 1136 5756
rect 1188 5704 1200 5756
rect 1252 5704 1264 5710
rect 1316 5704 1328 5710
rect 1380 5704 1392 5710
rect 1444 5704 1456 5710
rect 1508 5704 1520 5710
rect 1572 5704 1584 5710
rect 1636 5704 1648 5710
rect 1700 5704 1712 5710
rect 1764 5704 1776 5710
rect 1828 5704 1840 5710
rect 1892 5704 1904 5710
rect 1956 5704 1968 5710
rect 2020 5704 2032 5710
rect 2084 5704 2096 5710
rect 2148 5704 2160 5710
rect 2212 5704 2224 5710
rect 2276 5704 2288 5710
rect 2340 5704 2352 5710
rect 2404 5704 2416 5710
rect 2468 5704 2480 5710
rect 2532 5704 2544 5710
rect 2596 5704 2608 5710
rect 2660 5704 2672 5710
rect 2724 5704 2736 5710
rect 2788 5704 2800 5710
rect 2852 5704 2864 5710
rect 2916 5704 2928 5710
rect 2980 5704 2992 5710
rect 3044 5704 3056 5710
rect 3108 5704 3120 5710
rect 3172 5704 3184 5710
rect 3236 5704 3248 5710
rect 3300 5704 3312 5710
rect 3364 5704 3376 5710
rect 3428 5704 3440 5710
rect 3684 5704 3696 5710
rect 3748 5704 3760 5710
rect 3812 5704 3824 5710
rect 3876 5704 3888 5710
rect 3940 5704 3952 5710
rect 4004 5704 4016 5710
rect 4068 5704 4080 5710
rect 4132 5704 4144 5710
rect 4196 5704 4208 5710
rect 4260 5704 4272 5710
rect 4324 5704 4336 5710
rect 4388 5704 4400 5710
rect 4452 5704 4464 5710
rect 4516 5704 4528 5710
rect 4580 5704 4592 5710
rect 9458 5710 9459 5756
rect 4772 5704 4784 5710
rect 4836 5704 4848 5710
rect 4900 5704 4912 5710
rect 4964 5704 4976 5710
rect 5028 5704 5040 5710
rect 5092 5704 5104 5710
rect 5156 5704 5168 5710
rect 5220 5704 5232 5710
rect 5284 5704 5296 5710
rect 5348 5704 5360 5710
rect 5412 5704 5424 5710
rect 5476 5704 5488 5710
rect 5540 5704 5552 5710
rect 5604 5704 5616 5710
rect 5668 5704 5680 5710
rect 5732 5704 5744 5710
rect 5796 5704 5808 5710
rect 5860 5704 5872 5710
rect 5924 5704 5936 5710
rect 5988 5704 6000 5710
rect 6052 5704 6064 5710
rect 6116 5704 6128 5710
rect 6180 5704 6192 5710
rect 6244 5704 6256 5710
rect 6308 5704 6320 5710
rect 6372 5704 6384 5710
rect 6436 5704 6448 5710
rect 6500 5704 6512 5710
rect 6564 5704 6576 5710
rect 6628 5704 6640 5710
rect 6692 5704 6704 5710
rect 6756 5704 6768 5710
rect 6820 5704 6832 5710
rect 6884 5704 6896 5710
rect 6948 5704 6960 5710
rect 7012 5704 7024 5710
rect 7076 5704 7088 5710
rect 7140 5704 7152 5710
rect 7204 5704 7216 5710
rect 7268 5704 7280 5710
rect 7332 5704 7344 5710
rect 7396 5704 7408 5710
rect 7460 5704 7472 5710
rect 7524 5704 7536 5710
rect 7588 5704 7600 5710
rect 7652 5704 7664 5710
rect 7716 5704 7728 5710
rect 7780 5704 7792 5710
rect 7844 5704 7856 5710
rect 7908 5704 7920 5710
rect 7972 5704 7984 5710
rect 8036 5704 8048 5710
rect 8100 5704 8112 5710
rect 8164 5704 8176 5710
rect 8228 5704 8240 5710
rect 8292 5704 8304 5710
rect 8356 5704 8368 5710
rect 8420 5704 8432 5710
rect 8484 5704 8496 5710
rect 8548 5704 8560 5710
rect 8612 5704 8624 5710
rect 8676 5704 8688 5710
rect 8740 5704 8752 5710
rect 8804 5704 8816 5710
rect 8868 5704 8880 5710
rect 8932 5704 8944 5710
rect 8996 5704 9008 5710
rect 9060 5704 9072 5710
rect 9124 5704 9136 5710
rect 9188 5704 9200 5710
rect 9252 5704 9264 5710
rect 9316 5704 9329 5710
rect 9381 5704 9394 5710
rect 9446 5704 9459 5710
rect 9511 5704 9524 5756
rect 9576 5704 9589 5756
rect 9641 5744 9654 5756
rect 9706 5744 9719 5756
rect 9771 5744 9784 5756
rect 9836 5744 9849 5756
rect 9901 5744 9914 5756
rect 9643 5710 9654 5744
rect 9717 5710 9719 5744
rect 9901 5710 9905 5744
rect 9641 5704 9654 5710
rect 9706 5704 9719 5710
rect 9771 5704 9784 5710
rect 9836 5704 9849 5710
rect 9901 5704 9914 5710
rect 9966 5704 9979 5756
rect 10031 5704 10044 5756
rect 10096 5704 10109 5756
rect 10161 5704 10174 5756
rect 10226 5744 10239 5756
rect 10291 5744 10389 5756
rect 10235 5710 10239 5744
rect 10311 5710 10349 5744
rect 10383 5710 10389 5744
rect 10226 5704 10239 5710
rect 10291 5704 10389 5710
rect 82 4126 88 5704
tri 88 5670 122 5704 nw
tri 3429 5670 3463 5704 ne
rect 3463 5638 3469 5704
rect 3647 5638 3653 5704
tri 3653 5670 3687 5704 nw
tri 4552 5670 4586 5704 ne
rect 3463 5599 3653 5638
rect 3463 5565 3469 5599
rect 3503 5565 3541 5599
rect 3575 5565 3613 5599
rect 3647 5565 3653 5599
rect 3463 5526 3653 5565
rect 3463 5492 3469 5526
rect 3503 5492 3541 5526
rect 3575 5492 3613 5526
rect 3647 5492 3653 5526
rect -30 4087 88 4126
rect -30 4053 -24 4087
rect 10 4053 48 4087
rect 82 4053 88 4087
rect -30 4014 88 4053
rect -30 3980 -24 4014
rect 10 3980 48 4014
rect 82 3980 88 4014
rect -30 3941 88 3980
rect -30 3907 -24 3941
rect 10 3907 48 3941
rect 82 3907 88 3941
rect -30 3868 88 3907
rect -30 3834 -24 3868
rect 10 3834 48 3868
rect 82 3834 88 3868
rect -30 3795 88 3834
rect -30 3761 -24 3795
rect 10 3761 48 3795
rect 82 3761 88 3795
rect -30 3722 88 3761
rect -30 3688 -24 3722
rect 10 3688 48 3722
rect 82 3688 88 3722
rect -30 3649 88 3688
rect -30 3615 -24 3649
rect 10 3615 48 3649
rect 82 3615 88 3649
rect -30 3576 88 3615
rect -30 3542 -24 3576
rect 10 3542 48 3576
rect 82 3542 88 3576
rect -30 3503 88 3542
rect -30 3469 -24 3503
rect 10 3469 48 3503
rect 82 3469 88 3503
rect -30 3430 88 3469
rect -30 3396 -24 3430
rect 10 3396 48 3430
rect 82 3396 88 3430
rect -30 3357 88 3396
rect -30 3323 -24 3357
rect 10 3323 48 3357
rect 82 3323 88 3357
rect -30 3284 88 3323
rect -30 3250 -24 3284
rect 10 3250 48 3284
rect 82 3250 88 3284
rect -30 3211 88 3250
rect -30 3177 -24 3211
rect 10 3177 48 3211
rect 82 3177 88 3211
rect -30 3138 88 3177
rect -30 3104 -24 3138
rect 10 3104 48 3138
rect 82 3104 88 3138
rect -30 3065 88 3104
rect -30 3031 -24 3065
rect 10 3031 48 3065
rect 82 3031 88 3065
rect -30 2992 88 3031
rect -30 2958 -24 2992
rect 10 2958 48 2992
rect 82 2958 88 2992
rect -30 2919 88 2958
rect -30 2885 -24 2919
rect 10 2885 48 2919
rect 82 2885 88 2919
rect -30 2846 88 2885
rect -30 2812 -24 2846
rect 10 2812 48 2846
rect 82 2812 88 2846
rect -30 2773 88 2812
rect -30 2739 -24 2773
rect 10 2739 48 2773
rect 82 2739 88 2773
rect -30 2700 88 2739
rect -30 2666 -24 2700
rect 10 2666 48 2700
rect 82 2666 88 2700
rect -30 2627 88 2666
rect -30 2593 -24 2627
rect 10 2593 48 2627
rect 82 2593 88 2627
rect -30 2554 88 2593
rect -30 2520 -24 2554
rect 10 2520 48 2554
rect 82 2520 88 2554
rect -30 2481 88 2520
rect -30 2447 -24 2481
rect 10 2447 48 2481
rect 82 2447 88 2481
rect -30 2408 88 2447
rect -30 2374 -24 2408
rect 10 2374 48 2408
rect 82 2374 88 2408
rect -30 2335 88 2374
rect -30 2301 -24 2335
rect 10 2301 48 2335
rect 82 2301 88 2335
rect -30 2262 88 2301
rect -30 2228 -24 2262
rect 10 2228 48 2262
rect 82 2228 88 2262
rect -30 2189 88 2228
rect -30 2155 -24 2189
rect 10 2155 48 2189
rect 82 2155 88 2189
rect -30 2116 88 2155
rect -30 2082 -24 2116
rect 10 2082 48 2116
rect 82 2082 88 2116
rect -30 2043 88 2082
rect -30 2009 -24 2043
rect 10 2009 48 2043
rect 82 2009 88 2043
rect -30 1970 88 2009
rect -30 1936 -24 1970
rect 10 1936 48 1970
rect 82 1936 88 1970
rect -30 1897 88 1936
rect -30 1863 -24 1897
rect 10 1863 48 1897
rect 82 1863 88 1897
rect -30 1824 88 1863
rect -30 1790 -24 1824
rect 10 1790 48 1824
rect 82 1790 88 1824
rect -30 1751 88 1790
rect -30 1717 -24 1751
rect 10 1717 48 1751
rect 82 1717 88 1751
rect -30 1678 88 1717
rect -30 1644 -24 1678
rect 10 1644 48 1678
rect 82 1644 88 1678
rect -30 1605 88 1644
rect -30 1571 -24 1605
rect 10 1571 48 1605
rect 82 1571 88 1605
rect -30 1532 88 1571
rect -30 1498 -24 1532
rect 10 1498 48 1532
rect 82 1498 88 1532
rect -30 1459 88 1498
rect -30 1425 -24 1459
rect 10 1425 48 1459
rect 82 1425 88 1459
rect -30 1386 88 1425
rect -30 1352 -24 1386
rect 10 1352 48 1386
rect 82 1352 88 1386
rect -30 1313 88 1352
rect -30 1279 -24 1313
rect 10 1279 48 1313
rect 82 1279 88 1313
rect -30 1240 88 1279
rect -30 1206 -24 1240
rect 10 1206 48 1240
rect 82 1206 88 1240
rect -30 1167 88 1206
rect -30 1133 -24 1167
rect 10 1133 48 1167
rect 82 1133 88 1167
rect -30 1094 88 1133
rect -30 1060 -24 1094
rect 10 1060 48 1094
rect 82 1060 88 1094
rect -30 1021 88 1060
rect -30 987 -24 1021
rect 10 987 48 1021
rect 82 987 88 1021
rect -30 948 88 987
rect -30 914 -24 948
rect 10 914 48 948
rect 82 914 88 948
rect -30 875 88 914
rect -30 841 -24 875
rect 10 841 48 875
rect 82 841 88 875
rect -30 802 88 841
rect -30 768 -24 802
rect 10 768 48 802
rect 82 768 88 802
rect -30 729 88 768
rect -30 695 -24 729
rect 10 695 48 729
rect 82 695 88 729
rect -30 656 88 695
rect -30 622 -24 656
rect 10 622 48 656
rect 82 622 88 656
rect -30 583 88 622
rect -30 549 -24 583
rect 10 549 48 583
rect 82 549 88 583
rect -30 510 88 549
rect -30 476 -24 510
rect 10 476 48 510
rect 82 476 88 510
rect -30 437 88 476
rect 320 5474 3293 5480
rect 320 5440 408 5474
rect 442 5440 490 5474
rect 524 5440 572 5474
rect 606 5440 654 5474
rect 688 5440 736 5474
rect 770 5440 819 5474
rect 853 5440 929 5474
rect 963 5440 1001 5474
rect 1035 5440 1073 5474
rect 1107 5440 1145 5474
rect 1179 5440 1217 5474
rect 1251 5440 1289 5474
rect 1323 5440 1361 5474
rect 1395 5440 1433 5474
rect 1467 5440 1505 5474
rect 1539 5440 1577 5474
rect 1611 5440 1649 5474
rect 1683 5440 1721 5474
rect 1755 5440 1794 5474
rect 1828 5440 1867 5474
rect 1901 5440 1940 5474
rect 1974 5440 2013 5474
rect 2047 5440 2086 5474
rect 2120 5440 2159 5474
rect 2193 5440 2232 5474
rect 2266 5440 2305 5474
rect 2339 5440 2378 5474
rect 2412 5440 2451 5474
rect 2485 5440 2524 5474
rect 2558 5440 2597 5474
rect 2631 5440 2670 5474
rect 2704 5440 2743 5474
rect 2777 5440 2816 5474
rect 2850 5440 2889 5474
rect 2923 5440 2962 5474
rect 2996 5440 3035 5474
rect 3069 5440 3108 5474
rect 3142 5440 3181 5474
rect 3215 5440 3293 5474
rect 320 5434 3293 5440
rect 320 5419 385 5434
tri 385 5419 400 5434 nw
tri 3213 5419 3228 5434 ne
rect 3228 5419 3293 5434
rect 320 5415 381 5419
tri 381 5415 385 5419 nw
tri 3228 5415 3232 5419 ne
rect 3232 5415 3293 5419
rect 320 5402 368 5415
tri 368 5402 381 5415 nw
tri 3232 5402 3245 5415 ne
rect 3245 5402 3293 5415
rect 320 5368 326 5402
rect 360 5368 366 5402
tri 366 5400 368 5402 nw
tri 3245 5400 3247 5402 ne
rect 320 5329 366 5368
rect 320 5295 326 5329
rect 360 5295 366 5329
rect 320 5256 366 5295
rect 3247 5368 3253 5402
rect 3287 5368 3293 5402
rect 3247 5330 3293 5368
rect 3247 5296 3253 5330
rect 3287 5296 3293 5330
rect 320 5222 326 5256
rect 360 5222 366 5256
rect 320 5183 366 5222
rect 320 5149 326 5183
rect 360 5149 366 5183
rect 320 5110 366 5149
rect 320 5076 326 5110
rect 360 5076 366 5110
rect 320 5037 366 5076
rect 320 5003 326 5037
rect 360 5003 366 5037
rect 320 4964 366 5003
rect 320 4930 326 4964
rect 360 4930 366 4964
rect 320 4891 366 4930
rect 320 4857 326 4891
rect 360 4857 366 4891
rect 320 4818 366 4857
rect 320 4784 326 4818
rect 360 4784 366 4818
rect 320 4745 366 4784
rect 320 4711 326 4745
rect 360 4711 366 4745
rect 320 4672 366 4711
rect 320 4638 326 4672
rect 360 4638 366 4672
rect 320 4599 366 4638
rect 320 4565 326 4599
rect 360 4565 366 4599
rect 320 4526 366 4565
rect 320 4492 326 4526
rect 360 4492 366 4526
rect 320 4453 366 4492
rect 320 4419 326 4453
rect 360 4419 366 4453
rect 320 4380 366 4419
rect 320 4346 326 4380
rect 360 4346 366 4380
rect 320 4307 366 4346
rect 320 4273 326 4307
rect 360 4273 366 4307
rect 320 4234 366 4273
rect 320 4200 326 4234
rect 360 4200 366 4234
rect 320 4161 366 4200
rect 320 4127 326 4161
rect 360 4127 366 4161
rect 320 4088 366 4127
rect 320 4054 326 4088
rect 360 4054 366 4088
rect 320 4016 366 4054
rect 320 3982 326 4016
rect 360 3982 366 4016
rect 320 3944 366 3982
rect 320 3910 326 3944
rect 360 3910 366 3944
rect 320 3872 366 3910
rect 320 3838 326 3872
rect 360 3838 366 3872
rect 320 3800 366 3838
rect 320 3766 326 3800
rect 360 3766 366 3800
rect 320 3728 366 3766
rect 320 3694 326 3728
rect 360 3694 366 3728
rect 320 3656 366 3694
rect 320 3622 326 3656
rect 360 3622 366 3656
rect 320 3584 366 3622
rect 320 3550 326 3584
rect 360 3550 366 3584
rect 320 3512 366 3550
rect 320 3478 326 3512
rect 360 3478 366 3512
rect 320 3440 366 3478
rect 320 3406 326 3440
rect 360 3406 366 3440
rect 320 3368 366 3406
rect 320 3334 326 3368
rect 360 3334 366 3368
rect 320 3296 366 3334
rect 320 3262 326 3296
rect 360 3262 366 3296
rect 320 3224 366 3262
rect 320 3190 326 3224
rect 360 3190 366 3224
rect 320 3152 366 3190
rect 320 3118 326 3152
rect 360 3118 366 3152
rect 320 3080 366 3118
rect 320 3046 326 3080
rect 360 3046 366 3080
rect 320 3008 366 3046
rect 320 2974 326 3008
rect 360 2974 366 3008
rect 320 2936 366 2974
rect 320 2902 326 2936
rect 360 2902 366 2936
rect 320 2864 366 2902
rect 320 2830 326 2864
rect 360 2830 366 2864
rect 320 2792 366 2830
rect 320 2758 326 2792
rect 360 2758 366 2792
rect 320 2720 366 2758
rect 320 2686 326 2720
rect 360 2686 366 2720
rect 320 2648 366 2686
rect 320 2614 326 2648
rect 360 2614 366 2648
rect 320 2576 366 2614
rect 320 2542 326 2576
rect 360 2542 366 2576
rect 320 2504 366 2542
rect 320 2470 326 2504
rect 360 2470 366 2504
rect 320 2432 366 2470
rect 320 2398 326 2432
rect 360 2398 366 2432
rect 320 2360 366 2398
rect 320 2326 326 2360
rect 360 2326 366 2360
rect 320 2288 366 2326
rect 320 2254 326 2288
rect 360 2254 366 2288
rect 320 2216 366 2254
rect 320 2182 326 2216
rect 360 2182 366 2216
rect 320 2144 366 2182
rect 320 2110 326 2144
rect 360 2110 366 2144
rect 320 2072 366 2110
rect 320 2038 326 2072
rect 360 2038 366 2072
rect 320 2000 366 2038
rect 320 1966 326 2000
rect 360 1966 366 2000
rect 320 1928 366 1966
rect 320 1894 326 1928
rect 360 1894 366 1928
rect 320 1856 366 1894
rect 320 1822 326 1856
rect 360 1822 366 1856
rect 320 1784 366 1822
rect 320 1750 326 1784
rect 360 1750 366 1784
rect 320 1712 366 1750
rect 320 1678 326 1712
rect 360 1678 366 1712
rect 320 1640 366 1678
rect 320 1606 326 1640
rect 360 1606 366 1640
rect 320 1568 366 1606
rect 320 1534 326 1568
rect 360 1534 366 1568
rect 320 1496 366 1534
rect 320 1462 326 1496
rect 360 1462 366 1496
rect 320 1424 366 1462
rect 320 1390 326 1424
rect 360 1390 366 1424
rect 320 1352 366 1390
rect 320 1318 326 1352
rect 360 1318 366 1352
rect 320 1280 366 1318
rect 320 1246 326 1280
rect 360 1246 366 1280
rect 320 1208 366 1246
rect 320 1174 326 1208
rect 360 1174 366 1208
rect 320 1136 366 1174
rect 320 1102 326 1136
rect 360 1102 366 1136
rect 320 1064 366 1102
rect 320 1030 326 1064
rect 360 1030 366 1064
rect 320 992 366 1030
rect 320 958 326 992
rect 360 958 366 992
rect 320 920 366 958
rect 320 886 326 920
rect 360 886 366 920
rect 320 848 366 886
rect 320 814 326 848
rect 360 814 366 848
rect 320 776 366 814
rect 320 742 326 776
rect 360 742 366 776
rect 320 704 366 742
rect 320 670 326 704
rect 360 670 366 704
rect 320 632 366 670
rect 519 5228 525 5280
rect 577 5274 658 5280
rect 710 5274 791 5280
rect 843 5274 923 5280
rect 975 5274 1055 5280
rect 1107 5274 1187 5280
rect 1239 5274 1319 5280
rect 1371 5274 1451 5280
rect 1503 5274 1583 5280
rect 1635 5274 1715 5280
rect 1767 5274 1847 5280
rect 1899 5274 1979 5280
rect 2031 5274 2111 5280
rect 2163 5274 2243 5280
rect 2295 5274 2375 5280
rect 2427 5274 2507 5280
rect 2559 5274 2639 5280
rect 2691 5274 2771 5280
rect 2823 5274 2903 5280
rect 2955 5274 3035 5280
rect 577 5240 600 5274
rect 634 5240 658 5274
rect 710 5240 750 5274
rect 784 5240 791 5274
rect 859 5240 900 5274
rect 975 5240 976 5274
rect 1010 5240 1052 5274
rect 1107 5240 1128 5274
rect 1162 5240 1187 5274
rect 1239 5240 1280 5274
rect 1314 5240 1319 5274
rect 1390 5240 1432 5274
rect 1503 5240 1508 5274
rect 1542 5240 1583 5274
rect 1635 5240 1660 5274
rect 1694 5240 1715 5274
rect 1770 5240 1846 5274
rect 1899 5240 1921 5274
rect 1955 5240 1979 5274
rect 2031 5240 2071 5274
rect 2105 5240 2111 5274
rect 2180 5240 2221 5274
rect 2295 5240 2297 5274
rect 2331 5240 2373 5274
rect 2427 5240 2449 5274
rect 2483 5240 2507 5274
rect 2559 5240 2601 5274
rect 2635 5240 2639 5274
rect 2711 5240 2753 5274
rect 2823 5240 2829 5274
rect 2863 5240 2903 5274
rect 2955 5240 2981 5274
rect 3015 5240 3035 5274
rect 577 5228 658 5240
rect 710 5228 791 5240
rect 843 5228 923 5240
rect 975 5228 1055 5240
rect 1107 5228 1187 5240
rect 1239 5228 1319 5240
rect 1371 5228 1451 5240
rect 1503 5228 1583 5240
rect 1635 5228 1715 5240
rect 1767 5228 1847 5240
rect 1899 5228 1979 5240
rect 2031 5228 2111 5240
rect 2163 5228 2243 5240
rect 2295 5228 2375 5240
rect 2427 5228 2507 5240
rect 2559 5228 2639 5240
rect 2691 5228 2771 5240
rect 2823 5228 2903 5240
rect 2955 5228 3035 5240
rect 3087 5228 3093 5280
rect 519 5214 3093 5228
rect 519 5162 525 5214
rect 577 5202 658 5214
rect 710 5202 791 5214
rect 843 5202 923 5214
rect 975 5202 1055 5214
rect 1107 5202 1187 5214
rect 1239 5202 1319 5214
rect 1371 5202 1451 5214
rect 1503 5202 1583 5214
rect 1635 5202 1715 5214
rect 1767 5202 1847 5214
rect 1899 5202 1979 5214
rect 2031 5202 2111 5214
rect 2163 5202 2243 5214
rect 2295 5202 2375 5214
rect 2427 5202 2507 5214
rect 2559 5202 2639 5214
rect 2691 5202 2771 5214
rect 2823 5202 2903 5214
rect 2955 5202 3035 5214
rect 577 5168 597 5202
rect 631 5168 658 5202
rect 710 5168 750 5202
rect 784 5168 791 5202
rect 859 5168 900 5202
rect 975 5168 976 5202
rect 1010 5168 1052 5202
rect 1107 5168 1128 5202
rect 1162 5168 1187 5202
rect 1239 5168 1280 5202
rect 1314 5168 1319 5202
rect 1390 5168 1432 5202
rect 1503 5168 1508 5202
rect 1542 5168 1583 5202
rect 1635 5168 1660 5202
rect 1694 5168 1715 5202
rect 1770 5168 1846 5202
rect 1899 5168 1921 5202
rect 1955 5168 1979 5202
rect 2031 5168 2071 5202
rect 2105 5168 2111 5202
rect 2180 5168 2221 5202
rect 2295 5168 2297 5202
rect 2331 5168 2373 5202
rect 2427 5168 2449 5202
rect 2483 5168 2507 5202
rect 2559 5168 2601 5202
rect 2635 5168 2639 5202
rect 2711 5168 2753 5202
rect 2823 5168 2829 5202
rect 2863 5168 2903 5202
rect 577 5162 658 5168
rect 710 5162 791 5168
rect 843 5162 923 5168
rect 975 5162 1055 5168
rect 1107 5162 1187 5168
rect 1239 5162 1319 5168
rect 1371 5162 1451 5168
rect 1503 5162 1583 5168
rect 1635 5162 1715 5168
rect 1767 5162 1847 5168
rect 1899 5162 1979 5168
rect 2031 5162 2111 5168
rect 2163 5162 2243 5168
rect 2295 5162 2375 5168
rect 2427 5162 2507 5168
rect 2559 5162 2639 5168
rect 2691 5162 2771 5168
rect 2823 5162 2903 5168
rect 2955 5162 2981 5202
rect 519 5129 637 5162
rect 519 5095 525 5129
rect 559 5095 597 5129
rect 631 5095 637 5129
tri 637 5128 671 5162 nw
tri 2941 5128 2975 5162 ne
rect 519 5056 637 5095
rect 519 5022 525 5056
rect 559 5022 597 5056
rect 631 5022 637 5056
rect 519 4983 637 5022
rect 519 4949 525 4983
rect 559 4949 597 4983
rect 631 4949 637 4983
rect 519 4910 637 4949
rect 519 4876 525 4910
rect 559 4876 597 4910
rect 631 4876 637 4910
rect 519 4837 637 4876
rect 519 4803 525 4837
rect 559 4803 597 4837
rect 631 4803 637 4837
rect 519 4764 637 4803
rect 519 4730 525 4764
rect 559 4730 597 4764
rect 631 4730 637 4764
rect 519 4691 637 4730
rect 519 4657 525 4691
rect 559 4657 597 4691
rect 631 4657 637 4691
rect 519 4618 637 4657
rect 519 4584 525 4618
rect 559 4584 597 4618
rect 631 4584 637 4618
rect 519 4545 637 4584
rect 519 4511 525 4545
rect 559 4511 597 4545
rect 631 4511 637 4545
rect 519 4472 637 4511
rect 519 4438 525 4472
rect 559 4438 597 4472
rect 631 4438 637 4472
rect 519 4399 637 4438
rect 519 4365 525 4399
rect 559 4365 597 4399
rect 631 4365 637 4399
rect 519 4326 637 4365
rect 519 4292 525 4326
rect 559 4292 597 4326
rect 631 4292 637 4326
rect 519 4253 637 4292
rect 519 4219 525 4253
rect 559 4219 597 4253
rect 631 4219 637 4253
rect 519 4180 637 4219
rect 519 4146 525 4180
rect 559 4146 597 4180
rect 631 4146 637 4180
rect 519 4107 637 4146
rect 519 4073 525 4107
rect 559 4073 597 4107
rect 631 4073 637 4107
rect 519 4034 637 4073
rect 519 4000 525 4034
rect 559 4000 597 4034
rect 631 4000 637 4034
rect 519 3961 637 4000
rect 519 3927 525 3961
rect 559 3927 597 3961
rect 631 3927 637 3961
rect 519 3888 637 3927
rect 519 3854 525 3888
rect 559 3854 597 3888
rect 631 3854 637 3888
rect 519 3815 637 3854
rect 519 3781 525 3815
rect 559 3781 597 3815
rect 631 3781 637 3815
rect 519 3742 637 3781
rect 519 3708 525 3742
rect 559 3708 597 3742
rect 631 3708 637 3742
rect 519 3669 637 3708
rect 519 3635 525 3669
rect 559 3635 597 3669
rect 631 3635 637 3669
rect 519 3596 637 3635
rect 519 3562 525 3596
rect 559 3562 597 3596
rect 631 3562 637 3596
rect 519 3523 637 3562
rect 519 3489 525 3523
rect 559 3489 597 3523
rect 631 3489 637 3523
rect 519 3450 637 3489
rect 519 3416 525 3450
rect 559 3416 597 3450
rect 631 3416 637 3450
rect 519 3377 637 3416
rect 519 3343 525 3377
rect 559 3343 597 3377
rect 631 3343 637 3377
rect 519 3304 637 3343
rect 519 3270 525 3304
rect 559 3270 597 3304
rect 631 3270 637 3304
rect 519 3231 637 3270
rect 519 3197 525 3231
rect 559 3197 597 3231
rect 631 3197 637 3231
rect 519 3158 637 3197
rect 519 3124 525 3158
rect 559 3124 597 3158
rect 631 3124 637 3158
rect 519 3085 637 3124
rect 688 4114 740 5105
rect 688 4047 740 4062
rect 688 3980 740 3995
rect 688 3913 740 3928
rect 688 3846 740 3861
rect 688 3779 740 3794
rect 688 3712 740 3727
rect 688 3645 740 3660
rect 688 3578 740 3593
rect 688 3103 740 3526
rect 844 4854 896 5105
rect 844 4787 896 4802
rect 844 4720 896 4735
rect 844 4653 896 4668
rect 844 4586 896 4601
rect 844 4519 896 4534
rect 844 4452 896 4467
rect 844 4385 896 4400
rect 844 4318 896 4333
rect 844 3103 896 4266
rect 1000 4114 1052 5105
rect 1000 4047 1052 4062
rect 1000 3980 1052 3995
rect 1000 3913 1052 3928
rect 1000 3846 1052 3861
rect 1000 3779 1052 3794
rect 1000 3712 1052 3727
rect 1000 3645 1052 3660
rect 1000 3578 1052 3593
rect 1000 3103 1052 3526
rect 1156 4854 1208 5105
rect 1156 4787 1208 4802
rect 1156 4720 1208 4735
rect 1156 4653 1208 4668
rect 1156 4586 1208 4601
rect 1156 4519 1208 4534
rect 1156 4452 1208 4467
rect 1156 4385 1208 4400
rect 1156 4318 1208 4333
rect 1156 3103 1208 4266
rect 1312 4114 1364 5105
rect 1312 4047 1364 4062
rect 1312 3980 1364 3995
rect 1312 3913 1364 3928
rect 1312 3846 1364 3861
rect 1312 3779 1364 3794
rect 1312 3712 1364 3727
rect 1312 3645 1364 3660
rect 1312 3578 1364 3593
rect 1312 3103 1364 3526
rect 1468 4854 1520 5105
rect 1468 4787 1520 4802
rect 1468 4720 1520 4735
rect 1468 4653 1520 4668
rect 1468 4586 1520 4601
rect 1468 4519 1520 4534
rect 1468 4452 1520 4467
rect 1468 4385 1520 4400
rect 1468 4318 1520 4333
rect 1468 3103 1520 4266
rect 1624 4114 1676 5105
rect 1624 4047 1676 4062
rect 1624 3980 1676 3995
rect 1624 3913 1676 3928
rect 1624 3846 1676 3861
rect 1624 3779 1676 3794
rect 1624 3712 1676 3727
rect 1624 3645 1676 3660
rect 1624 3578 1676 3593
rect 1624 3103 1676 3526
rect 1780 4854 1832 5105
rect 1780 4787 1832 4802
rect 1780 4720 1832 4735
rect 1780 4653 1832 4668
rect 1780 4586 1832 4601
rect 1780 4519 1832 4534
rect 1780 4452 1832 4467
rect 1780 4385 1832 4400
rect 1780 4318 1832 4333
rect 1780 3103 1832 4266
rect 1936 4114 1988 5105
rect 1936 4047 1988 4062
rect 1936 3980 1988 3995
rect 1936 3913 1988 3928
rect 1936 3846 1988 3861
rect 1936 3779 1988 3794
rect 1936 3712 1988 3727
rect 1936 3645 1988 3660
rect 1936 3578 1988 3593
rect 1936 3103 1988 3526
rect 2092 4854 2144 5105
rect 2092 4787 2144 4802
rect 2092 4720 2144 4735
rect 2092 4653 2144 4668
rect 2092 4586 2144 4601
rect 2092 4519 2144 4534
rect 2092 4452 2144 4467
rect 2092 4385 2144 4400
rect 2092 4318 2144 4333
rect 2092 3103 2144 4266
rect 2248 4114 2300 5105
rect 2248 4047 2300 4062
rect 2248 3980 2300 3995
rect 2248 3913 2300 3928
rect 2248 3846 2300 3861
rect 2248 3779 2300 3794
rect 2248 3712 2300 3727
rect 2248 3645 2300 3660
rect 2248 3578 2300 3593
rect 2248 3103 2300 3526
rect 2404 4854 2456 5105
rect 2404 4787 2456 4802
rect 2404 4720 2456 4735
rect 2404 4653 2456 4668
rect 2404 4586 2456 4601
rect 2404 4519 2456 4534
rect 2404 4452 2456 4467
rect 2404 4385 2456 4400
rect 2404 4318 2456 4333
rect 2404 3103 2456 4266
rect 2560 4114 2612 5105
rect 2560 4047 2612 4062
rect 2560 3980 2612 3995
rect 2560 3913 2612 3928
rect 2560 3846 2612 3861
rect 2560 3779 2612 3794
rect 2560 3712 2612 3727
rect 2560 3645 2612 3660
rect 2560 3578 2612 3593
rect 2560 3103 2612 3526
rect 2716 4854 2768 5105
rect 2716 4787 2768 4802
rect 2716 4720 2768 4735
rect 2716 4653 2768 4668
rect 2716 4586 2768 4601
rect 2716 4519 2768 4534
rect 2716 4452 2768 4467
rect 2716 4385 2768 4400
rect 2716 4318 2768 4333
rect 2716 3103 2768 4266
rect 2872 4114 2924 5105
rect 2872 4047 2924 4062
rect 2872 3980 2924 3995
rect 2872 3913 2924 3928
rect 2872 3846 2924 3861
rect 2872 3779 2924 3794
rect 2872 3712 2924 3727
rect 2872 3645 2924 3660
rect 2872 3578 2924 3593
rect 2872 3103 2924 3526
rect 2975 4016 2981 5162
rect 3087 4016 3093 5214
rect 3247 5258 3293 5296
rect 3247 5224 3253 5258
rect 3287 5224 3293 5258
rect 3247 5186 3293 5224
rect 3247 5152 3253 5186
rect 3287 5152 3293 5186
rect 3247 5114 3293 5152
rect 3247 5080 3253 5114
rect 3287 5080 3293 5114
rect 3247 5042 3293 5080
rect 3247 5008 3253 5042
rect 3287 5008 3293 5042
tri 3240 4970 3247 4977 se
rect 3247 4970 3293 5008
rect 3463 5453 3653 5492
rect 3463 5419 3469 5453
rect 3503 5419 3541 5453
rect 3575 5419 3613 5453
rect 3647 5419 3653 5453
rect 3463 5380 3653 5419
rect 3463 5346 3469 5380
rect 3503 5346 3541 5380
rect 3575 5346 3613 5380
rect 3647 5346 3653 5380
rect 3463 5307 3653 5346
rect 3463 5273 3469 5307
rect 3503 5273 3541 5307
rect 3575 5273 3613 5307
rect 3647 5273 3653 5307
rect 3463 5234 3653 5273
rect 3463 5200 3469 5234
rect 3503 5200 3541 5234
rect 3575 5200 3613 5234
rect 3647 5200 3653 5234
rect 3463 5161 3653 5200
rect 3463 5127 3469 5161
rect 3503 5127 3541 5161
rect 3575 5127 3613 5161
rect 3647 5127 3653 5161
rect 3463 5088 3653 5127
rect 3463 5054 3469 5088
rect 3503 5054 3541 5088
rect 3575 5054 3613 5088
rect 3647 5054 3653 5088
rect 3463 5015 3653 5054
rect 3463 4981 3469 5015
rect 3503 4981 3541 5015
rect 3575 4981 3613 5015
rect 3647 4981 3653 5015
tri 3213 4943 3240 4970 se
rect 3240 4943 3253 4970
rect 3287 4943 3293 4970
tri 3293 4943 3327 4977 sw
rect 3204 4891 3210 4943
rect 3262 4898 3274 4936
rect 3326 4891 3332 4943
rect 3463 4942 3653 4981
rect 3463 4908 3469 4942
rect 3503 4908 3541 4942
rect 3575 4908 3613 4942
rect 3647 4908 3653 4942
tri 3213 4864 3240 4891 ne
rect 3240 4864 3253 4891
rect 3287 4869 3305 4891
tri 3305 4869 3327 4891 nw
rect 3463 4869 3653 4908
rect 3287 4864 3293 4869
tri 3240 4857 3247 4864 ne
rect 3247 4826 3293 4864
tri 3293 4857 3305 4869 nw
rect 3247 4792 3253 4826
rect 3287 4792 3293 4826
rect 3247 4754 3293 4792
rect 3247 4720 3253 4754
rect 3287 4720 3293 4754
rect 3247 4682 3293 4720
rect 3247 4648 3253 4682
rect 3287 4648 3293 4682
rect 3247 4610 3293 4648
rect 3247 4576 3253 4610
rect 3287 4576 3293 4610
rect 3247 4538 3293 4576
rect 3247 4504 3253 4538
rect 3287 4504 3293 4538
rect 3247 4466 3293 4504
rect 3247 4432 3253 4466
rect 3287 4432 3293 4466
rect 3247 4394 3293 4432
rect 3247 4360 3253 4394
rect 3287 4360 3293 4394
rect 3247 4322 3293 4360
rect 3247 4288 3253 4322
rect 3287 4288 3293 4322
tri 3236 4251 3247 4262 se
rect 3247 4251 3293 4288
rect 3463 4835 3469 4869
rect 3503 4835 3541 4869
rect 3575 4835 3613 4869
rect 3647 4835 3653 4869
rect 3463 4796 3653 4835
rect 3463 4762 3469 4796
rect 3503 4762 3541 4796
rect 3575 4762 3613 4796
rect 3647 4762 3653 4796
rect 3463 4723 3653 4762
rect 3463 4689 3469 4723
rect 3503 4689 3541 4723
rect 3575 4689 3613 4723
rect 3647 4689 3653 4723
rect 3463 4650 3653 4689
rect 3463 4616 3469 4650
rect 3503 4616 3541 4650
rect 3575 4616 3613 4650
rect 3647 4616 3653 4650
rect 3463 4577 3653 4616
rect 3463 4543 3469 4577
rect 3503 4543 3541 4577
rect 3575 4543 3613 4577
rect 3647 4543 3653 4577
rect 3463 4504 3653 4543
rect 3463 4470 3469 4504
rect 3503 4470 3541 4504
rect 3575 4470 3613 4504
rect 3647 4470 3653 4504
rect 3463 4431 3653 4470
rect 3463 4397 3469 4431
rect 3503 4397 3541 4431
rect 3575 4397 3613 4431
rect 3647 4397 3653 4431
rect 3463 4358 3653 4397
rect 3463 4324 3469 4358
rect 3503 4324 3541 4358
rect 3575 4324 3613 4358
rect 3647 4324 3653 4358
rect 3463 4285 3653 4324
tri 3293 4251 3304 4262 sw
rect 3463 4251 3469 4285
rect 3503 4251 3541 4285
rect 3575 4251 3613 4285
rect 3647 4251 3653 4285
tri 3235 4250 3236 4251 se
rect 3236 4250 3304 4251
tri 3213 4228 3235 4250 se
rect 3235 4228 3253 4250
rect 3287 4228 3304 4250
tri 3304 4228 3327 4251 sw
rect 3204 4176 3210 4228
rect 3262 4178 3274 4216
rect 3326 4176 3332 4228
rect 3463 4212 3653 4251
rect 3463 4178 3469 4212
rect 3503 4178 3541 4212
rect 3575 4178 3613 4212
rect 3647 4178 3653 4212
tri 3213 4144 3245 4176 ne
rect 3245 4144 3253 4176
rect 3287 4144 3293 4176
tri 3245 4142 3247 4144 ne
rect 2975 3977 3093 4016
rect 2975 3943 2981 3977
rect 3015 3943 3053 3977
rect 3087 3943 3093 3977
rect 2975 3904 3093 3943
rect 2975 3870 2981 3904
rect 3015 3870 3053 3904
rect 3087 3870 3093 3904
rect 2975 3831 3093 3870
rect 2975 3797 2981 3831
rect 3015 3797 3053 3831
rect 3087 3797 3093 3831
rect 2975 3758 3093 3797
rect 2975 3724 2981 3758
rect 3015 3724 3053 3758
rect 3087 3724 3093 3758
rect 2975 3685 3093 3724
rect 2975 3651 2981 3685
rect 3015 3651 3053 3685
rect 3087 3651 3093 3685
rect 2975 3612 3093 3651
rect 2975 3578 2981 3612
rect 3015 3578 3053 3612
rect 3087 3578 3093 3612
rect 2975 3539 3093 3578
rect 2975 3505 2981 3539
rect 3015 3505 3053 3539
rect 3087 3505 3093 3539
rect 2975 3466 3093 3505
rect 2975 3432 2981 3466
rect 3015 3432 3053 3466
rect 3087 3432 3093 3466
rect 2975 3393 3093 3432
rect 2975 3359 2981 3393
rect 3015 3359 3053 3393
rect 3087 3359 3093 3393
rect 2975 3320 3093 3359
rect 2975 3286 2981 3320
rect 3015 3286 3053 3320
rect 3087 3286 3093 3320
rect 2975 3247 3093 3286
rect 2975 3213 2981 3247
rect 3015 3213 3053 3247
rect 3087 3213 3093 3247
rect 2975 3174 3093 3213
rect 2975 3140 2981 3174
rect 3015 3140 3053 3174
rect 3087 3140 3093 3174
rect 519 3051 525 3085
rect 559 3051 597 3085
rect 631 3051 637 3085
rect 519 3012 637 3051
rect 2975 3101 3093 3140
rect 2975 3067 2981 3101
rect 3015 3067 3053 3101
rect 3087 3067 3093 3101
rect 519 2978 525 3012
rect 559 2978 597 3012
rect 631 2978 637 3012
rect 762 3041 1335 3049
rect 1387 3041 1471 3049
rect 1523 3041 1607 3049
rect 1659 3041 1743 3049
rect 1795 3041 1879 3049
rect 1931 3041 2015 3049
rect 2067 3041 2151 3049
rect 2203 3041 2287 3049
rect 2339 3041 2423 3049
rect 2475 3041 2560 3049
rect 2612 3041 2697 3049
rect 2749 3041 2841 3049
rect 762 3007 774 3041
rect 808 3007 847 3041
rect 881 3007 920 3041
rect 954 3007 993 3041
rect 1027 3007 1066 3041
rect 1100 3007 1139 3041
rect 1173 3007 1211 3041
rect 1245 3007 1283 3041
rect 1317 3007 1335 3041
rect 1389 3007 1427 3041
rect 1461 3007 1471 3041
rect 1533 3007 1571 3041
rect 1605 3007 1607 3041
rect 1677 3007 1715 3041
rect 1821 3007 1859 3041
rect 1965 3007 2003 3041
rect 2067 3007 2075 3041
rect 2109 3007 2147 3041
rect 2203 3007 2219 3041
rect 2253 3007 2287 3041
rect 2339 3007 2363 3041
rect 2397 3007 2423 3041
rect 2475 3007 2507 3041
rect 2541 3007 2560 3041
rect 2613 3007 2651 3041
rect 2685 3007 2697 3041
rect 2757 3007 2795 3041
rect 2829 3007 2841 3041
rect 762 2997 1335 3007
rect 1387 2997 1471 3007
rect 1523 2997 1607 3007
rect 1659 2997 1743 3007
rect 1795 2997 1879 3007
rect 1931 2997 2015 3007
rect 2067 2997 2151 3007
rect 2203 2997 2287 3007
rect 2339 2997 2423 3007
rect 2475 2997 2560 3007
rect 2612 2997 2697 3007
rect 2749 2997 2841 3007
rect 2975 3028 3093 3067
rect 519 2939 637 2978
rect 519 2905 525 2939
rect 559 2905 597 2939
rect 631 2905 637 2939
rect 2975 2994 2981 3028
rect 3015 2994 3053 3028
rect 3087 2994 3093 3028
rect 2975 2955 3093 2994
rect 519 2866 637 2905
rect 762 2921 1335 2930
rect 1387 2921 1471 2930
rect 1523 2921 1607 2930
rect 1659 2921 1743 2930
rect 1795 2921 1879 2930
rect 1931 2921 2015 2930
rect 2067 2921 2151 2930
rect 2203 2921 2287 2930
rect 2339 2921 2423 2930
rect 2475 2921 2560 2930
rect 2612 2921 2697 2930
rect 2749 2921 2841 2930
rect 762 2887 774 2921
rect 808 2887 847 2921
rect 881 2887 920 2921
rect 954 2887 993 2921
rect 1027 2887 1066 2921
rect 1100 2887 1139 2921
rect 1173 2887 1211 2921
rect 1245 2887 1283 2921
rect 1317 2887 1335 2921
rect 1389 2887 1427 2921
rect 1461 2887 1471 2921
rect 1533 2887 1571 2921
rect 1605 2887 1607 2921
rect 1677 2887 1715 2921
rect 1821 2887 1859 2921
rect 1965 2887 2003 2921
rect 2067 2887 2075 2921
rect 2109 2887 2147 2921
rect 2203 2887 2219 2921
rect 2253 2887 2287 2921
rect 2339 2887 2363 2921
rect 2397 2887 2423 2921
rect 2475 2887 2507 2921
rect 2541 2887 2560 2921
rect 2613 2887 2651 2921
rect 2685 2887 2697 2921
rect 2757 2887 2795 2921
rect 2829 2887 2841 2921
rect 762 2878 1335 2887
rect 1387 2878 1471 2887
rect 1523 2878 1607 2887
rect 1659 2878 1743 2887
rect 1795 2878 1879 2887
rect 1931 2878 2015 2887
rect 2067 2878 2151 2887
rect 2203 2878 2287 2887
rect 2339 2878 2423 2887
rect 2475 2878 2560 2887
rect 2612 2878 2697 2887
rect 2749 2878 2841 2887
rect 2975 2921 2981 2955
rect 3015 2921 3053 2955
rect 3087 2921 3093 2955
rect 2975 2882 3093 2921
rect 519 2832 525 2866
rect 559 2832 597 2866
rect 631 2832 637 2866
rect 519 2793 637 2832
rect 2975 2848 2981 2882
rect 3015 2848 3053 2882
rect 3087 2848 3093 2882
rect 519 2759 525 2793
rect 559 2759 597 2793
rect 631 2759 637 2793
rect 519 2720 637 2759
rect 519 2686 525 2720
rect 559 2686 597 2720
rect 631 2686 637 2720
rect 519 2647 637 2686
rect 519 2613 525 2647
rect 559 2613 597 2647
rect 631 2613 637 2647
rect 519 2574 637 2613
rect 519 2540 525 2574
rect 559 2540 597 2574
rect 631 2540 637 2574
rect 519 2501 637 2540
rect 519 2467 525 2501
rect 559 2467 597 2501
rect 631 2467 637 2501
rect 519 2428 637 2467
rect 519 2394 525 2428
rect 559 2394 597 2428
rect 631 2394 637 2428
rect 519 2355 637 2394
rect 519 2321 525 2355
rect 559 2321 597 2355
rect 631 2321 637 2355
rect 519 2282 637 2321
rect 519 2248 525 2282
rect 559 2248 597 2282
rect 631 2248 637 2282
rect 519 2209 637 2248
rect 519 2175 525 2209
rect 559 2175 597 2209
rect 631 2175 637 2209
rect 519 2136 637 2175
rect 519 2102 525 2136
rect 559 2102 597 2136
rect 631 2102 637 2136
rect 519 2063 637 2102
rect 519 2029 525 2063
rect 559 2029 597 2063
rect 631 2029 637 2063
rect 519 1990 637 2029
rect 519 1956 525 1990
rect 559 1956 597 1990
rect 631 1956 637 1990
rect 519 1917 637 1956
rect 519 731 525 1917
rect 631 804 637 1917
rect 688 2564 740 2825
rect 688 2493 740 2512
rect 688 2422 740 2441
rect 688 2351 740 2370
rect 688 2280 740 2299
rect 688 2209 740 2228
rect 688 2138 740 2157
rect 688 2068 740 2086
rect 688 823 740 2016
rect 844 1865 896 2825
rect 844 1798 896 1813
rect 844 1731 896 1746
rect 844 1664 896 1679
rect 844 1597 896 1612
rect 844 1530 896 1545
rect 844 1463 896 1478
rect 844 1396 896 1411
rect 844 1329 896 1344
rect 844 823 896 1277
rect 1000 2604 1052 2825
rect 1000 2537 1052 2552
rect 1000 2470 1052 2485
rect 1000 2403 1052 2418
rect 1000 2336 1052 2351
rect 1000 2269 1052 2284
rect 1000 2202 1052 2217
rect 1000 2135 1052 2150
rect 1000 2068 1052 2083
rect 1000 823 1052 2016
rect 1156 1865 1208 2825
rect 1156 1798 1208 1813
rect 1156 1731 1208 1746
rect 1156 1664 1208 1679
rect 1156 1597 1208 1612
rect 1156 1530 1208 1545
rect 1156 1463 1208 1478
rect 1156 1396 1208 1411
rect 1156 1329 1208 1344
rect 1156 823 1208 1277
rect 1312 2604 1364 2825
rect 1312 2537 1364 2552
rect 1312 2470 1364 2485
rect 1312 2403 1364 2418
rect 1312 2336 1364 2351
rect 1312 2269 1364 2284
rect 1312 2202 1364 2217
rect 1312 2135 1364 2150
rect 1312 2068 1364 2083
rect 1312 823 1364 2016
rect 1468 1865 1520 2825
rect 1468 1798 1520 1813
rect 1468 1731 1520 1746
rect 1468 1664 1520 1679
rect 1468 1597 1520 1612
rect 1468 1530 1520 1545
rect 1468 1463 1520 1478
rect 1468 1396 1520 1411
rect 1468 1329 1520 1344
rect 1468 823 1520 1277
rect 1624 2604 1676 2825
rect 1624 2537 1676 2552
rect 1624 2470 1676 2485
rect 1624 2403 1676 2418
rect 1624 2336 1676 2351
rect 1624 2269 1676 2284
rect 1624 2202 1676 2217
rect 1624 2135 1676 2150
rect 1624 2068 1676 2083
rect 1624 823 1676 2016
rect 1780 1865 1832 2825
rect 1780 1798 1832 1813
rect 1780 1731 1832 1746
rect 1780 1664 1832 1679
rect 1780 1597 1832 1612
rect 1780 1530 1832 1545
rect 1780 1463 1832 1478
rect 1780 1396 1832 1411
rect 1780 1329 1832 1344
rect 1780 823 1832 1277
rect 1936 2604 1988 2825
rect 1936 2537 1988 2552
rect 1936 2470 1988 2485
rect 1936 2403 1988 2418
rect 1936 2336 1988 2351
rect 1936 2269 1988 2284
rect 1936 2202 1988 2217
rect 1936 2135 1988 2150
rect 1936 2068 1988 2083
rect 1936 823 1988 2016
rect 2092 1865 2144 2825
rect 2092 1798 2144 1813
rect 2092 1731 2144 1746
rect 2092 1664 2144 1679
rect 2092 1597 2144 1612
rect 2092 1530 2144 1545
rect 2092 1463 2144 1478
rect 2092 1396 2144 1411
rect 2092 1329 2144 1344
rect 2092 823 2144 1277
rect 2248 2604 2300 2825
rect 2248 2537 2300 2552
rect 2248 2470 2300 2485
rect 2248 2403 2300 2418
rect 2248 2336 2300 2351
rect 2248 2269 2300 2284
rect 2248 2202 2300 2217
rect 2248 2135 2300 2150
rect 2248 2068 2300 2083
rect 2248 823 2300 2016
rect 2404 1865 2456 2825
rect 2404 1798 2456 1813
rect 2404 1731 2456 1746
rect 2404 1664 2456 1679
rect 2404 1597 2456 1612
rect 2404 1530 2456 1545
rect 2404 1463 2456 1478
rect 2404 1396 2456 1411
rect 2404 1329 2456 1344
rect 2404 823 2456 1277
rect 2560 2604 2612 2825
rect 2560 2537 2612 2552
rect 2560 2470 2612 2485
rect 2560 2403 2612 2418
rect 2560 2336 2612 2351
rect 2560 2269 2612 2284
rect 2560 2202 2612 2217
rect 2560 2135 2612 2150
rect 2560 2068 2612 2083
rect 2560 823 2612 2016
rect 2716 1865 2768 2825
rect 2716 1798 2768 1813
rect 2716 1731 2768 1746
rect 2716 1664 2768 1679
rect 2716 1597 2768 1612
rect 2716 1530 2768 1545
rect 2716 1463 2768 1478
rect 2716 1396 2768 1411
rect 2716 1329 2768 1344
rect 2716 823 2768 1277
rect 2872 2604 2924 2825
rect 2872 2537 2924 2552
rect 2872 2470 2924 2485
rect 2872 2403 2924 2418
rect 2872 2336 2924 2351
rect 2872 2269 2924 2284
rect 2872 2202 2924 2217
rect 2872 2135 2924 2150
rect 2872 2068 2924 2083
rect 2872 823 2924 2016
rect 2975 2809 3093 2848
rect 2975 2775 2981 2809
rect 3015 2775 3053 2809
rect 3087 2775 3093 2809
rect 2975 2736 3093 2775
rect 2975 2702 2981 2736
rect 3015 2702 3053 2736
rect 3087 2702 3093 2736
rect 2975 2663 3093 2702
rect 2975 2629 2981 2663
rect 3015 2629 3053 2663
rect 3087 2629 3093 2663
rect 2975 2590 3093 2629
rect 2975 2556 2981 2590
rect 3015 2556 3053 2590
rect 3087 2556 3093 2590
rect 2975 2517 3093 2556
rect 2975 2483 2981 2517
rect 3015 2483 3053 2517
rect 3087 2483 3093 2517
rect 2975 2444 3093 2483
rect 2975 2410 2981 2444
rect 3015 2410 3053 2444
rect 3087 2410 3093 2444
rect 2975 2371 3093 2410
rect 2975 2337 2981 2371
rect 3015 2337 3053 2371
rect 3087 2337 3093 2371
rect 2975 2298 3093 2337
rect 2975 2264 2981 2298
rect 3015 2264 3053 2298
rect 3087 2264 3093 2298
rect 2975 2225 3093 2264
rect 2975 2191 2981 2225
rect 3015 2191 3053 2225
rect 3087 2191 3093 2225
rect 2975 2152 3093 2191
rect 2975 2118 2981 2152
rect 3015 2118 3053 2152
rect 3087 2118 3093 2152
rect 2975 2079 3093 2118
rect 2975 2045 2981 2079
rect 3015 2045 3053 2079
rect 3087 2045 3093 2079
rect 2975 2006 3093 2045
rect 2975 1972 2981 2006
rect 3015 1972 3053 2006
rect 3087 1972 3093 2006
rect 3247 4106 3293 4144
tri 3293 4142 3327 4176 nw
rect 3247 4072 3253 4106
rect 3287 4072 3293 4106
rect 3247 4034 3293 4072
rect 3247 4000 3253 4034
rect 3287 4000 3293 4034
rect 3247 3962 3293 4000
rect 3247 3928 3253 3962
rect 3287 3928 3293 3962
rect 3247 3890 3293 3928
rect 3247 3856 3253 3890
rect 3287 3856 3293 3890
rect 3247 3818 3293 3856
rect 3247 3784 3253 3818
rect 3287 3784 3293 3818
rect 3247 3746 3293 3784
rect 3247 3712 3253 3746
rect 3287 3712 3293 3746
rect 3247 3674 3293 3712
rect 3247 3640 3253 3674
rect 3287 3640 3293 3674
rect 3247 3602 3293 3640
rect 3247 3568 3253 3602
rect 3287 3568 3293 3602
rect 3247 3530 3293 3568
rect 3247 3496 3253 3530
rect 3287 3496 3293 3530
rect 3247 3458 3293 3496
rect 3247 3424 3253 3458
rect 3287 3424 3293 3458
rect 3247 3386 3293 3424
rect 3247 3352 3253 3386
rect 3287 3352 3293 3386
rect 3247 3314 3293 3352
rect 3247 3280 3253 3314
rect 3287 3280 3293 3314
rect 3247 3242 3293 3280
rect 3247 3208 3253 3242
rect 3287 3208 3293 3242
rect 3247 3170 3293 3208
rect 3247 3136 3253 3170
rect 3287 3136 3293 3170
rect 3247 3098 3293 3136
rect 3247 3064 3253 3098
rect 3287 3064 3293 3098
rect 3247 3026 3293 3064
rect 3247 2992 3253 3026
rect 3287 2992 3293 3026
rect 3247 2954 3293 2992
rect 3247 2920 3253 2954
rect 3287 2920 3293 2954
rect 3247 2882 3293 2920
rect 3247 2848 3253 2882
rect 3287 2848 3293 2882
rect 3247 2810 3293 2848
rect 3247 2776 3253 2810
rect 3287 2776 3293 2810
rect 3247 2738 3293 2776
rect 3247 2704 3253 2738
rect 3287 2704 3293 2738
rect 3247 2666 3293 2704
rect 3247 2632 3253 2666
rect 3287 2632 3293 2666
rect 3247 2594 3293 2632
rect 3247 2560 3253 2594
rect 3287 2560 3293 2594
rect 3247 2522 3293 2560
rect 3247 2488 3253 2522
rect 3287 2488 3293 2522
rect 3247 2450 3293 2488
rect 3247 2416 3253 2450
rect 3287 2416 3293 2450
rect 3247 2378 3293 2416
rect 3247 2344 3253 2378
rect 3287 2344 3293 2378
rect 3247 2306 3293 2344
rect 3247 2272 3253 2306
rect 3287 2272 3293 2306
rect 3247 2234 3293 2272
rect 3247 2200 3253 2234
rect 3287 2200 3293 2234
rect 3247 2162 3293 2200
rect 3247 2128 3253 2162
rect 3287 2128 3293 2162
rect 3247 2090 3293 2128
rect 3247 2056 3253 2090
rect 3287 2056 3293 2090
rect 3247 2018 3293 2056
tri 3243 1984 3247 1988 se
rect 3247 1984 3253 2018
rect 3287 1984 3293 2018
rect 3463 4139 3653 4178
rect 3463 4105 3469 4139
rect 3503 4105 3541 4139
rect 3575 4105 3613 4139
rect 3647 4105 3653 4139
rect 3463 4066 3653 4105
rect 3463 4032 3469 4066
rect 3503 4032 3541 4066
rect 3575 4032 3613 4066
rect 3647 4032 3653 4066
rect 3463 3993 3653 4032
rect 3463 3959 3469 3993
rect 3503 3959 3541 3993
rect 3575 3959 3613 3993
rect 3647 3959 3653 3993
rect 3463 3920 3653 3959
rect 3463 3886 3469 3920
rect 3503 3886 3541 3920
rect 3575 3886 3613 3920
rect 3647 3886 3653 3920
rect 3463 3847 3653 3886
rect 3463 3813 3469 3847
rect 3503 3813 3541 3847
rect 3575 3813 3613 3847
rect 3647 3813 3653 3847
rect 3463 3774 3653 3813
rect 3463 3740 3469 3774
rect 3503 3740 3541 3774
rect 3575 3740 3613 3774
rect 3647 3740 3653 3774
rect 3463 3701 3653 3740
rect 3463 3667 3469 3701
rect 3503 3667 3541 3701
rect 3575 3667 3613 3701
rect 3647 3667 3653 3701
rect 3463 3628 3653 3667
rect 3463 3594 3469 3628
rect 3503 3594 3541 3628
rect 3575 3594 3613 3628
rect 3647 3594 3653 3628
rect 3463 3555 3653 3594
rect 3463 3521 3469 3555
rect 3503 3521 3541 3555
rect 3575 3521 3613 3555
rect 3647 3521 3653 3555
rect 3463 3482 3653 3521
rect 3463 3448 3469 3482
rect 3503 3448 3541 3482
rect 3575 3448 3613 3482
rect 3647 3448 3653 3482
rect 3463 3409 3653 3448
rect 3463 3375 3469 3409
rect 3503 3375 3541 3409
rect 3575 3375 3613 3409
rect 3647 3375 3653 3409
rect 3463 3336 3653 3375
rect 3463 3302 3469 3336
rect 3503 3302 3541 3336
rect 3575 3302 3613 3336
rect 3647 3302 3653 3336
rect 3463 3263 3653 3302
rect 3463 3229 3469 3263
rect 3503 3229 3541 3263
rect 3575 3229 3613 3263
rect 3647 3229 3653 3263
rect 3463 3190 3653 3229
rect 3463 3156 3469 3190
rect 3503 3156 3541 3190
rect 3575 3156 3613 3190
rect 3647 3156 3653 3190
rect 3463 3117 3653 3156
rect 3463 3083 3469 3117
rect 3503 3083 3541 3117
rect 3575 3083 3613 3117
rect 3647 3083 3653 3117
rect 3463 3044 3653 3083
rect 3463 3010 3469 3044
rect 3503 3010 3541 3044
rect 3575 3010 3613 3044
rect 3647 3010 3653 3044
rect 3463 2971 3653 3010
rect 3463 2937 3469 2971
rect 3503 2937 3541 2971
rect 3575 2937 3613 2971
rect 3647 2937 3653 2971
rect 3463 2898 3653 2937
rect 3463 2864 3469 2898
rect 3503 2864 3541 2898
rect 3575 2864 3613 2898
rect 3647 2864 3653 2898
rect 3463 2825 3653 2864
rect 3463 2791 3469 2825
rect 3503 2791 3541 2825
rect 3575 2791 3613 2825
rect 3647 2791 3653 2825
rect 3463 2752 3653 2791
rect 4586 5638 4592 5704
rect 4770 5671 4777 5704
tri 4777 5671 4810 5704 nw
tri 10237 5671 10270 5704 ne
rect 10270 5671 10389 5704
rect 4770 5638 4776 5671
tri 4776 5670 4777 5671 nw
tri 10270 5670 10271 5671 ne
rect 4586 5599 4776 5638
rect 4586 5565 4592 5599
rect 4626 5565 4664 5599
rect 4698 5565 4736 5599
rect 4770 5565 4776 5599
rect 4586 5526 4776 5565
rect 4586 5492 4592 5526
rect 4626 5492 4664 5526
rect 4698 5492 4736 5526
rect 4770 5492 4776 5526
rect 4586 5453 4776 5492
rect 10271 5637 10277 5671
rect 10311 5637 10349 5671
rect 10383 5637 10389 5671
rect 10271 5598 10389 5637
rect 10271 5564 10277 5598
rect 10311 5564 10349 5598
rect 10383 5564 10389 5598
rect 10271 5525 10389 5564
rect 10271 5491 10277 5525
rect 10311 5491 10349 5525
rect 10383 5491 10389 5525
rect 4586 5419 4592 5453
rect 4626 5419 4664 5453
rect 4698 5419 4736 5453
rect 4770 5419 4776 5453
rect 4586 5380 4776 5419
rect 4586 5346 4592 5380
rect 4626 5346 4664 5380
rect 4698 5346 4736 5380
rect 4770 5346 4776 5380
rect 4586 5307 4776 5346
rect 4586 5273 4592 5307
rect 4626 5273 4664 5307
rect 4698 5273 4736 5307
rect 4770 5273 4776 5307
rect 4586 5234 4776 5273
rect 4586 5200 4592 5234
rect 4626 5200 4664 5234
rect 4698 5200 4736 5234
rect 4770 5200 4776 5234
rect 4586 5161 4776 5200
rect 4586 5127 4592 5161
rect 4626 5127 4664 5161
rect 4698 5127 4736 5161
rect 4770 5127 4776 5161
rect 4586 5088 4776 5127
rect 4586 5054 4592 5088
rect 4626 5054 4664 5088
rect 4698 5054 4736 5088
rect 4770 5054 4776 5088
rect 4586 5015 4776 5054
rect 4586 4981 4592 5015
rect 4626 4981 4664 5015
rect 4698 4981 4736 5015
rect 4770 4981 4776 5015
rect 4586 4942 4776 4981
rect 4586 4908 4592 4942
rect 4626 4908 4664 4942
rect 4698 4908 4736 4942
rect 4770 4908 4776 4942
rect 4586 4869 4776 4908
rect 4586 4835 4592 4869
rect 4626 4835 4664 4869
rect 4698 4835 4736 4869
rect 4770 4835 4776 4869
rect 4586 4796 4776 4835
rect 4586 4762 4592 4796
rect 4626 4762 4664 4796
rect 4698 4762 4736 4796
rect 4770 4762 4776 4796
rect 4586 4723 4776 4762
rect 4586 4689 4592 4723
rect 4626 4689 4664 4723
rect 4698 4689 4736 4723
rect 4770 4689 4776 4723
rect 4586 4650 4776 4689
rect 4586 4616 4592 4650
rect 4626 4616 4664 4650
rect 4698 4616 4736 4650
rect 4770 4616 4776 4650
rect 4586 4577 4776 4616
rect 4586 4543 4592 4577
rect 4626 4543 4664 4577
rect 4698 4543 4736 4577
rect 4770 4543 4776 4577
rect 4586 4504 4776 4543
rect 4586 4470 4592 4504
rect 4626 4470 4664 4504
rect 4698 4470 4736 4504
rect 4770 4470 4776 4504
rect 4586 4431 4776 4470
rect 4586 4397 4592 4431
rect 4626 4397 4664 4431
rect 4698 4397 4736 4431
rect 4770 4397 4776 4431
rect 4586 4358 4776 4397
rect 4586 4324 4592 4358
rect 4626 4324 4664 4358
rect 4698 4324 4736 4358
rect 4770 4324 4776 4358
rect 4586 4285 4776 4324
rect 4586 4251 4592 4285
rect 4626 4251 4664 4285
rect 4698 4251 4736 4285
rect 4770 4251 4776 4285
rect 4586 4212 4776 4251
rect 4586 4178 4592 4212
rect 4626 4178 4664 4212
rect 4698 4178 4736 4212
rect 4770 4178 4776 4212
rect 4586 4139 4776 4178
rect 4586 4105 4592 4139
rect 4626 4105 4664 4139
rect 4698 4105 4736 4139
rect 4770 4105 4776 4139
rect 4586 4066 4776 4105
rect 4586 4032 4592 4066
rect 4626 4032 4664 4066
rect 4698 4032 4736 4066
rect 4770 4032 4776 4066
rect 4586 3993 4776 4032
rect 4586 3959 4592 3993
rect 4626 3959 4664 3993
rect 4698 3959 4736 3993
rect 4770 3959 4776 3993
rect 4586 3920 4776 3959
rect 4586 3886 4592 3920
rect 4626 3886 4664 3920
rect 4698 3886 4736 3920
rect 4770 3886 4776 3920
rect 4586 3847 4776 3886
rect 4586 3813 4592 3847
rect 4626 3813 4664 3847
rect 4698 3813 4736 3847
rect 4770 3813 4776 3847
rect 4586 3774 4776 3813
rect 4586 3740 4592 3774
rect 4626 3740 4664 3774
rect 4698 3740 4736 3774
rect 4770 3740 4776 3774
rect 4586 3701 4776 3740
rect 4586 3667 4592 3701
rect 4626 3667 4664 3701
rect 4698 3667 4736 3701
rect 4770 3667 4776 3701
rect 4586 3628 4776 3667
rect 4586 3594 4592 3628
rect 4626 3594 4664 3628
rect 4698 3594 4736 3628
rect 4770 3594 4776 3628
rect 4586 3555 4776 3594
rect 4586 3521 4592 3555
rect 4626 3521 4664 3555
rect 4698 3521 4736 3555
rect 4770 3521 4776 3555
rect 4586 3482 4776 3521
rect 4586 3448 4592 3482
rect 4626 3448 4664 3482
rect 4698 3448 4736 3482
rect 4770 3448 4776 3482
rect 4586 3409 4776 3448
rect 4586 3375 4592 3409
rect 4626 3375 4664 3409
rect 4698 3375 4736 3409
rect 4770 3375 4776 3409
rect 4586 3336 4776 3375
rect 4586 3302 4592 3336
rect 4626 3302 4664 3336
rect 4698 3302 4736 3336
rect 4770 3302 4776 3336
rect 4586 3263 4776 3302
rect 4586 3229 4592 3263
rect 4626 3229 4664 3263
rect 4698 3229 4736 3263
rect 4770 3229 4776 3263
rect 4586 3190 4776 3229
rect 4586 3156 4592 3190
rect 4626 3156 4664 3190
rect 4698 3156 4736 3190
rect 4770 3156 4776 3190
rect 4586 3117 4776 3156
rect 4586 3083 4592 3117
rect 4626 3083 4664 3117
rect 4698 3083 4736 3117
rect 4770 3083 4776 3117
rect 4586 3044 4776 3083
rect 4586 3010 4592 3044
rect 4626 3010 4664 3044
rect 4698 3010 4736 3044
rect 4770 3010 4776 3044
rect 4586 2971 4776 3010
rect 4586 2937 4592 2971
rect 4626 2937 4664 2971
rect 4698 2937 4736 2971
rect 4770 2937 4776 2971
rect 4586 2898 4776 2937
rect 4586 2864 4592 2898
rect 4626 2864 4664 2898
rect 4698 2864 4736 2898
rect 4770 2864 4776 2898
rect 4586 2825 4776 2864
rect 4586 2791 4592 2825
rect 4626 2791 4664 2825
rect 4698 2791 4736 2825
rect 4770 2791 4776 2825
rect 3463 2718 3469 2752
rect 3503 2718 3541 2752
rect 3575 2718 3613 2752
rect 3647 2718 3653 2752
rect 3463 2679 3653 2718
rect 3463 2645 3469 2679
rect 3503 2645 3541 2679
rect 3575 2645 3613 2679
rect 3647 2645 3653 2679
rect 3463 2606 3653 2645
rect 3463 2572 3469 2606
rect 3503 2572 3541 2606
rect 3575 2572 3613 2606
rect 3647 2572 3653 2606
rect 3463 2533 3653 2572
rect 3463 2499 3469 2533
rect 3503 2499 3541 2533
rect 3575 2499 3613 2533
rect 3647 2499 3653 2533
rect 3979 2703 3985 2755
rect 4037 2703 4165 2755
rect 4217 2703 4223 2755
rect 3979 2564 4223 2703
rect 3979 2530 3992 2564
rect 4026 2530 4084 2564
rect 4118 2530 4177 2564
rect 4211 2530 4223 2564
rect 3979 2524 4223 2530
rect 4586 2752 4776 2791
rect 4586 2718 4592 2752
rect 4626 2718 4664 2752
rect 4698 2718 4736 2752
rect 4770 2718 4776 2752
rect 4586 2679 4776 2718
rect 4586 2645 4592 2679
rect 4626 2645 4664 2679
rect 4698 2645 4736 2679
rect 4770 2645 4776 2679
rect 4586 2606 4776 2645
rect 4586 2572 4592 2606
rect 4626 2572 4664 2606
rect 4698 2572 4736 2606
rect 4770 2572 4776 2606
rect 4586 2533 4776 2572
rect 3463 2460 3653 2499
rect 3463 2426 3469 2460
rect 3503 2426 3541 2460
rect 3575 2426 3613 2460
rect 3647 2426 3653 2460
rect 3463 2387 3653 2426
rect 3463 2353 3469 2387
rect 3503 2353 3541 2387
rect 3575 2353 3613 2387
rect 3647 2353 3653 2387
rect 3463 2314 3653 2353
rect 3463 2280 3469 2314
rect 3503 2280 3541 2314
rect 3575 2280 3613 2314
rect 3647 2280 3653 2314
rect 3463 2241 3653 2280
rect 3463 2207 3469 2241
rect 3503 2207 3541 2241
rect 3575 2207 3613 2241
rect 3647 2207 3653 2241
rect 3463 2168 3653 2207
rect 3463 2134 3469 2168
rect 3503 2134 3541 2168
rect 3575 2134 3613 2168
rect 3647 2134 3653 2168
rect 3463 2095 3653 2134
rect 3463 2061 3469 2095
rect 3503 2061 3541 2095
rect 3575 2061 3613 2095
rect 3647 2061 3653 2095
rect 3463 2022 3653 2061
rect 3463 1988 3469 2022
rect 3503 1988 3541 2022
rect 3575 1988 3613 2022
rect 3647 1988 3653 2022
rect 2975 1933 3093 1972
tri 3230 1971 3243 1984 se
rect 3243 1971 3293 1984
tri 3293 1971 3310 1988 sw
tri 3215 1956 3230 1971 se
rect 3230 1956 3310 1971
tri 3310 1956 3325 1971 sw
tri 3213 1954 3215 1956 se
rect 3215 1954 3325 1956
tri 3325 1954 3327 1956 sw
rect 2975 1899 2981 1933
rect 3015 1899 3053 1933
rect 3087 1899 3093 1933
rect 3204 1902 3210 1954
rect 3262 1946 3274 1954
rect 3262 1902 3274 1912
rect 3326 1902 3332 1954
rect 3463 1949 3653 1988
rect 3463 1915 3469 1949
rect 3503 1915 3541 1949
rect 3575 1915 3613 1949
rect 3647 1915 3653 1949
rect 2975 1860 3093 1899
tri 3213 1898 3217 1902 ne
rect 3217 1898 3323 1902
tri 3323 1898 3327 1902 nw
tri 3217 1881 3234 1898 ne
rect 3234 1881 3306 1898
tri 3306 1881 3323 1898 nw
tri 3234 1876 3239 1881 ne
rect 3239 1876 3301 1881
tri 3301 1876 3306 1881 nw
rect 3463 1876 3653 1915
tri 3239 1874 3241 1876 ne
rect 3241 1874 3293 1876
tri 3241 1868 3247 1874 ne
rect 2975 1826 2981 1860
rect 3015 1826 3053 1860
rect 3087 1826 3093 1860
rect 2975 1787 3093 1826
rect 2975 1753 2981 1787
rect 3015 1753 3053 1787
rect 3087 1753 3093 1787
rect 2975 1714 3093 1753
rect 2975 1680 2981 1714
rect 3015 1680 3053 1714
rect 3087 1680 3093 1714
rect 2975 1641 3093 1680
rect 2975 1607 2981 1641
rect 3015 1607 3053 1641
rect 3087 1607 3093 1641
rect 2975 1568 3093 1607
rect 2975 1534 2981 1568
rect 3015 1534 3053 1568
rect 3087 1534 3093 1568
rect 2975 1495 3093 1534
rect 2975 1461 2981 1495
rect 3015 1461 3053 1495
rect 3087 1461 3093 1495
rect 2975 1422 3093 1461
rect 2975 1388 2981 1422
rect 3015 1388 3053 1422
rect 3087 1388 3093 1422
rect 2975 1349 3093 1388
rect 2975 1315 2981 1349
rect 3015 1315 3053 1349
rect 3087 1315 3093 1349
rect 2975 1276 3093 1315
rect 2975 1242 2981 1276
rect 3015 1242 3053 1276
rect 3087 1242 3093 1276
rect 3247 1840 3253 1874
rect 3287 1840 3293 1874
tri 3293 1868 3301 1876 nw
rect 3247 1801 3293 1840
rect 3247 1767 3253 1801
rect 3287 1767 3293 1801
rect 3247 1728 3293 1767
rect 3247 1694 3253 1728
rect 3287 1694 3293 1728
rect 3247 1655 3293 1694
rect 3247 1621 3253 1655
rect 3287 1621 3293 1655
rect 3247 1582 3293 1621
rect 3247 1548 3253 1582
rect 3287 1548 3293 1582
rect 3247 1509 3293 1548
rect 3247 1475 3253 1509
rect 3287 1475 3293 1509
rect 3247 1436 3293 1475
rect 3247 1402 3253 1436
rect 3287 1402 3293 1436
rect 3247 1363 3293 1402
rect 3247 1329 3253 1363
rect 3287 1329 3293 1363
rect 3247 1290 3293 1329
tri 3230 1256 3247 1273 se
rect 3247 1256 3253 1290
rect 3287 1256 3293 1290
rect 3463 1842 3469 1876
rect 3503 1842 3541 1876
rect 3575 1842 3613 1876
rect 3647 1842 3653 1876
rect 3463 1803 3653 1842
rect 3463 1769 3469 1803
rect 3503 1769 3541 1803
rect 3575 1769 3613 1803
rect 3647 1769 3653 1803
rect 3463 1730 3653 1769
rect 2975 1203 3093 1242
tri 3213 1239 3230 1256 se
rect 3230 1239 3293 1256
tri 3293 1239 3327 1273 sw
rect 2975 1169 2981 1203
rect 3015 1169 3053 1203
rect 3087 1169 3093 1203
rect 3204 1187 3210 1239
rect 3262 1217 3274 1239
rect 3326 1187 3332 1239
tri 3213 1183 3217 1187 ne
rect 3217 1183 3253 1187
rect 3287 1183 3293 1187
rect 2975 1130 3093 1169
tri 3217 1153 3247 1183 ne
rect 2975 1096 2981 1130
rect 3015 1096 3053 1130
rect 3087 1096 3093 1130
rect 2975 1057 3093 1096
rect 2975 1023 2981 1057
rect 3015 1023 3053 1057
rect 3087 1023 3093 1057
rect 2975 984 3093 1023
rect 2975 950 2981 984
rect 3015 950 3053 984
rect 3087 950 3093 984
rect 2975 911 3093 950
rect 2975 877 2981 911
rect 3015 877 3053 911
rect 3087 877 3093 911
rect 2975 838 3093 877
tri 637 804 638 805 sw
tri 2974 804 2975 805 se
rect 2975 804 2981 838
rect 3015 804 3053 838
rect 3087 804 3093 838
rect 631 779 638 804
tri 638 779 663 804 sw
tri 2949 779 2974 804 se
rect 2974 779 3093 804
rect 631 771 663 779
tri 663 771 671 779 sw
tri 2941 771 2949 779 se
rect 2949 771 3093 779
rect 631 765 3093 771
rect 631 731 670 765
rect 704 731 743 765
rect 777 731 816 765
rect 850 731 889 765
rect 923 731 962 765
rect 996 731 1035 765
rect 1069 731 1108 765
rect 1142 731 1181 765
rect 519 693 1181 731
rect 519 659 597 693
rect 631 659 670 693
rect 704 659 743 693
rect 777 659 816 693
rect 850 659 889 693
rect 923 659 962 693
rect 996 659 1035 693
rect 1069 659 1108 693
rect 1142 659 1181 693
rect 3015 731 3053 765
rect 3087 731 3093 765
rect 3015 659 3093 731
rect 519 653 3093 659
rect 3247 1144 3293 1183
tri 3293 1153 3327 1187 nw
rect 3247 1110 3253 1144
rect 3287 1110 3293 1144
rect 3247 1071 3293 1110
rect 3247 1037 3253 1071
rect 3287 1037 3293 1071
rect 3247 998 3293 1037
rect 3247 964 3253 998
rect 3287 964 3293 998
rect 3247 925 3293 964
rect 3247 891 3253 925
rect 3287 891 3293 925
rect 3247 852 3293 891
rect 3247 818 3253 852
rect 3287 818 3293 852
rect 3247 779 3293 818
rect 3247 745 3253 779
rect 3287 745 3293 779
rect 3247 706 3293 745
rect 3247 672 3253 706
rect 3287 672 3293 706
rect 320 598 326 632
rect 360 598 366 632
rect 320 560 366 598
rect 320 526 326 560
rect 360 526 366 560
rect 3247 633 3293 672
rect 3247 599 3253 633
rect 3287 599 3293 633
rect 3247 560 3293 599
tri 366 526 371 531 sw
tri 3242 526 3247 531 se
rect 3247 526 3253 560
rect 3287 526 3293 560
rect 320 497 371 526
tri 371 497 400 526 sw
tri 3213 497 3242 526 se
rect 3242 497 3293 526
rect 320 445 326 497
rect 378 445 391 497
rect 443 445 456 497
rect 508 445 521 497
rect 573 488 586 497
rect 638 488 651 497
rect 703 488 716 497
rect 768 488 781 497
rect 833 488 846 497
rect 580 454 586 488
rect 833 454 842 488
rect 573 445 586 454
rect 638 445 651 454
rect 703 445 716 454
rect 768 445 781 454
rect 833 445 846 454
rect 898 445 911 497
rect 963 445 976 497
rect 1028 445 1041 497
rect 1093 488 1106 497
rect 1158 488 1171 497
rect 1223 488 1236 497
rect 1288 488 1301 497
rect 1353 488 1366 497
rect 1418 488 1431 497
rect 1097 454 1106 488
rect 1170 454 1171 488
rect 1353 454 1355 488
rect 1418 454 1428 488
rect 1093 445 1106 454
rect 1158 445 1171 454
rect 1223 445 1236 454
rect 1288 445 1301 454
rect 1353 445 1366 454
rect 1418 445 1431 454
rect 1483 445 1496 497
rect 1548 445 1561 497
rect 1613 445 1626 497
rect 1678 488 1691 497
rect 1743 488 1756 497
rect 1808 488 1821 497
rect 1873 488 1886 497
rect 1938 488 1951 497
rect 2003 488 2016 497
rect 1681 454 1691 488
rect 1754 454 1756 488
rect 1938 454 1939 488
rect 2003 454 2012 488
rect 1678 445 1691 454
rect 1743 445 1756 454
rect 1808 445 1821 454
rect 1873 445 1886 454
rect 1938 445 1951 454
rect 2003 445 2016 454
rect 2068 445 2081 497
rect 2133 445 2146 497
rect 2198 445 2211 497
rect 2263 488 2275 497
rect 2327 488 2339 497
rect 2391 488 2403 497
rect 2455 488 2467 497
rect 2519 488 2531 497
rect 2265 454 2275 488
rect 2338 454 2339 488
rect 2519 454 2523 488
rect 2263 445 2275 454
rect 2327 445 2339 454
rect 2391 445 2403 454
rect 2455 445 2467 454
rect 2519 445 2531 454
rect 2583 445 2595 497
rect 2647 445 2659 497
rect 2711 445 2723 497
rect 2775 488 2787 497
rect 2839 488 2851 497
rect 2903 488 2915 497
rect 2967 488 2979 497
rect 3031 488 3043 497
rect 2776 454 2787 488
rect 2849 454 2851 488
rect 3031 454 3034 488
rect 2775 445 2787 454
rect 2839 445 2851 454
rect 2903 445 2915 454
rect 2967 445 2979 454
rect 3031 445 3043 454
rect 3095 445 3107 497
rect 3159 445 3171 497
rect 3223 445 3235 497
rect 3287 445 3293 497
rect -30 403 -24 437
rect 10 403 48 437
rect 82 403 88 437
rect -30 364 88 403
rect -30 330 -24 364
rect 10 330 48 364
rect 82 330 88 364
rect -30 291 88 330
rect -30 257 -24 291
rect 10 257 48 291
rect 82 257 88 291
rect -30 224 88 257
tri 88 224 122 258 sw
tri 3429 224 3463 258 se
rect 3463 224 3469 1730
rect -30 218 3469 224
rect 3647 224 3653 1730
rect 3722 2480 3850 2518
rect 4363 2480 4491 2518
rect 3722 2446 3810 2480
rect 3844 2446 3850 2480
rect 3722 2406 3850 2446
rect 3722 2372 3810 2406
rect 3844 2372 3850 2406
rect 3722 2331 3850 2372
rect 3722 2297 3810 2331
rect 3844 2297 3850 2331
rect 3722 2256 3850 2297
rect 3722 2222 3810 2256
rect 3844 2222 3850 2256
rect 3722 2181 3850 2222
rect 3722 2147 3810 2181
rect 3844 2147 3850 2181
rect 3722 2106 3850 2147
rect 3722 2072 3810 2106
rect 3844 2072 3850 2106
rect 3722 2031 3850 2072
rect 3722 1997 3810 2031
rect 3844 1997 3850 2031
rect 3722 1956 3850 1997
rect 3722 1922 3810 1956
rect 3844 1922 3850 1956
rect 3722 1881 3850 1922
rect 3722 1847 3810 1881
rect 3844 1847 3850 1881
rect 3722 1806 3850 1847
rect 3722 1772 3810 1806
rect 3844 1772 3850 1806
rect 3722 1731 3850 1772
rect 3722 1697 3810 1731
rect 3844 1697 3850 1731
rect 3722 1656 3850 1697
rect 3722 1622 3810 1656
rect 3844 1622 3850 1656
rect 3722 1581 3850 1622
rect 3722 1547 3810 1581
rect 3844 1547 3850 1581
rect 3722 1506 3850 1547
rect 4079 2474 4131 2480
rect 4079 2401 4131 2422
rect 4079 2328 4131 2349
rect 4079 2255 4131 2276
rect 4079 2182 4131 2203
rect 4079 2108 4131 2130
rect 3722 1472 3810 1506
rect 3844 1472 3850 1506
rect 3722 546 3850 1472
rect 3926 1386 3972 1507
rect 4079 1466 4131 2056
rect 4363 2446 4369 2480
rect 4403 2446 4491 2480
rect 4363 2406 4491 2446
rect 4363 2372 4369 2406
rect 4403 2372 4491 2406
rect 4363 2331 4491 2372
rect 4363 2297 4369 2331
rect 4403 2297 4491 2331
rect 4363 2256 4491 2297
rect 4363 2222 4369 2256
rect 4403 2222 4491 2256
rect 4363 2181 4491 2222
rect 4363 2147 4369 2181
rect 4403 2147 4491 2181
rect 4363 2106 4491 2147
rect 4363 2072 4369 2106
rect 4403 2072 4491 2106
rect 4363 2031 4491 2072
rect 4363 1997 4369 2031
rect 4403 1997 4491 2031
rect 4363 1956 4491 1997
rect 4363 1922 4369 1956
rect 4403 1922 4491 1956
rect 4363 1881 4491 1922
rect 4363 1847 4369 1881
rect 4403 1847 4491 1881
rect 4363 1806 4491 1847
rect 4363 1772 4369 1806
rect 4403 1772 4491 1806
rect 4363 1731 4491 1772
rect 4363 1697 4369 1731
rect 4403 1697 4491 1731
rect 4363 1656 4491 1697
rect 4363 1622 4369 1656
rect 4403 1622 4491 1656
rect 4363 1581 4491 1622
rect 4363 1547 4369 1581
rect 4403 1547 4491 1581
tri 3972 1386 4006 1420 sw
tri 4204 1386 4238 1420 se
rect 4238 1386 4284 1507
rect 3926 1380 4284 1386
rect 3926 1346 3938 1380
rect 3972 1346 4013 1380
rect 4047 1346 4088 1380
rect 4122 1346 4163 1380
rect 4197 1346 4238 1380
rect 4272 1346 4284 1380
rect 3926 1308 4284 1346
rect 3926 1274 3938 1308
rect 3972 1274 4013 1308
rect 4047 1274 4088 1308
rect 4122 1274 4163 1308
rect 4197 1274 4238 1308
rect 4272 1274 4284 1308
rect 3926 1268 4284 1274
rect 4363 1506 4491 1547
rect 4363 1472 4369 1506
rect 4403 1472 4491 1506
tri 3850 546 3884 580 sw
tri 4329 546 4363 580 se
rect 4363 546 4491 1472
rect 3722 540 4491 546
rect 3722 506 3911 540
rect 3945 506 3985 540
rect 4019 506 4059 540
rect 4093 506 4133 540
rect 4167 506 4207 540
rect 4241 506 4281 540
rect 4315 506 4491 540
rect 3722 490 4491 506
rect 3722 438 3728 490
rect 3780 438 3828 490
rect 3880 468 3928 490
rect 3980 468 4029 490
rect 4081 468 4130 490
rect 4182 468 4231 490
rect 4283 468 4332 490
rect 3880 438 3911 468
rect 3980 438 3985 468
rect 3722 434 3911 438
rect 3945 434 3985 438
rect 4019 438 4029 468
rect 4093 438 4130 468
rect 4182 438 4207 468
rect 4315 438 4332 468
rect 4384 438 4433 490
rect 4485 438 4491 490
rect 4019 434 4059 438
rect 4093 434 4133 438
rect 4167 434 4207 438
rect 4241 434 4281 438
rect 4315 434 4491 438
rect 3722 428 4491 434
rect 4586 2499 4592 2533
rect 4626 2499 4664 2533
rect 4698 2499 4736 2533
rect 4770 2499 4776 2533
rect 4586 2460 4776 2499
rect 4586 2426 4592 2460
rect 4626 2426 4664 2460
rect 4698 2426 4736 2460
rect 4770 2426 4776 2460
rect 4586 2387 4776 2426
rect 4586 2353 4592 2387
rect 4626 2353 4664 2387
rect 4698 2353 4736 2387
rect 4770 2353 4776 2387
rect 4586 2314 4776 2353
rect 4586 2280 4592 2314
rect 4626 2280 4664 2314
rect 4698 2280 4736 2314
rect 4770 2280 4776 2314
rect 4586 2241 4776 2280
rect 4586 2207 4592 2241
rect 4626 2207 4664 2241
rect 4698 2207 4736 2241
rect 4770 2207 4776 2241
rect 4586 2168 4776 2207
rect 4586 2134 4592 2168
rect 4626 2134 4664 2168
rect 4698 2134 4736 2168
rect 4770 2134 4776 2168
rect 4586 2095 4776 2134
rect 4586 2061 4592 2095
rect 4626 2061 4664 2095
rect 4698 2061 4736 2095
rect 4770 2061 4776 2095
rect 4586 2022 4776 2061
rect 4586 1988 4592 2022
rect 4626 1988 4664 2022
rect 4698 1988 4736 2022
rect 4770 1988 4776 2022
rect 4586 1949 4776 1988
rect 4586 1915 4592 1949
rect 4626 1915 4664 1949
rect 4698 1915 4736 1949
rect 4770 1915 4776 1949
rect 4586 1876 4776 1915
rect 4586 1842 4592 1876
rect 4626 1842 4664 1876
rect 4698 1842 4736 1876
rect 4770 1842 4776 1876
rect 4586 1803 4776 1842
rect 4586 1769 4592 1803
rect 4626 1769 4664 1803
rect 4698 1769 4736 1803
rect 4770 1769 4776 1803
rect 4586 1730 4776 1769
tri 3653 224 3687 258 sw
tri 4552 224 4586 258 se
rect 4586 224 4592 1730
rect 3647 218 4592 224
rect 4770 224 4776 1730
rect 4925 5449 10035 5455
rect 4925 5415 5003 5449
rect 5037 5415 5076 5449
rect 5110 5415 5149 5449
rect 5183 5415 5222 5449
rect 5256 5415 5295 5449
rect 4925 5377 5295 5415
rect 4925 4114 4931 5377
rect 5037 5343 5076 5377
rect 5110 5343 5149 5377
rect 5183 5343 5222 5377
rect 5256 5343 5295 5377
rect 6049 5415 6125 5449
rect 6159 5415 6199 5449
rect 6233 5415 6272 5449
rect 6306 5415 6345 5449
rect 6379 5415 6418 5449
rect 6452 5415 6491 5449
rect 6525 5415 6564 5449
rect 6598 5415 6637 5449
rect 6671 5415 6710 5449
rect 6744 5415 6783 5449
rect 6817 5415 6856 5449
rect 6890 5415 6929 5449
rect 6963 5415 7002 5449
rect 7036 5415 7075 5449
rect 7109 5415 7148 5449
rect 7182 5415 7221 5449
rect 7255 5415 7294 5449
rect 7328 5415 7367 5449
rect 7401 5415 7440 5449
rect 7474 5415 7513 5449
rect 7547 5415 7586 5449
rect 7620 5415 7659 5449
rect 7693 5415 7732 5449
rect 7766 5415 7805 5449
rect 7839 5415 7878 5449
rect 7912 5415 7951 5449
rect 7985 5415 8024 5449
rect 8058 5415 8097 5449
rect 8131 5415 8170 5449
rect 8204 5415 8243 5449
rect 8277 5415 8316 5449
rect 8350 5415 8389 5449
rect 8423 5415 8462 5449
rect 8496 5415 8535 5449
rect 8569 5415 8608 5449
rect 8642 5415 8681 5449
rect 8715 5415 8754 5449
rect 8788 5415 8827 5449
rect 8861 5415 8900 5449
rect 8934 5415 8973 5449
rect 9007 5415 9046 5449
rect 9080 5415 9119 5449
rect 9153 5415 9192 5449
rect 9226 5415 9265 5449
rect 9299 5415 9338 5449
rect 9372 5415 9411 5449
rect 9445 5415 9484 5449
rect 9518 5415 9557 5449
rect 9591 5415 9630 5449
rect 9664 5415 9703 5449
rect 9737 5415 9776 5449
rect 9810 5415 9849 5449
rect 9883 5415 9922 5449
rect 9956 5415 10035 5449
rect 6049 5377 10035 5415
rect 6049 5343 6125 5377
rect 6159 5343 6199 5377
rect 6233 5343 6272 5377
rect 6306 5343 6345 5377
rect 6379 5343 6418 5377
rect 6452 5343 6491 5377
rect 6525 5343 6564 5377
rect 6598 5343 6637 5377
rect 6671 5343 6710 5377
rect 6744 5343 6783 5377
rect 6817 5343 6856 5377
rect 6890 5343 6929 5377
rect 6963 5343 7002 5377
rect 7036 5343 7075 5377
rect 7109 5343 7148 5377
rect 7182 5343 7221 5377
rect 7255 5343 7294 5377
rect 7328 5343 7367 5377
rect 7401 5343 7440 5377
rect 7474 5343 7513 5377
rect 7547 5343 7586 5377
rect 7620 5343 7659 5377
rect 7693 5343 7732 5377
rect 7766 5343 7805 5377
rect 7839 5343 7878 5377
rect 7912 5343 7951 5377
rect 7985 5343 8024 5377
rect 8058 5343 8097 5377
rect 8131 5343 8170 5377
rect 8204 5343 8243 5377
rect 8277 5343 8316 5377
rect 8350 5343 8389 5377
rect 8423 5343 8462 5377
rect 8496 5343 8535 5377
rect 8569 5343 8608 5377
rect 8642 5343 8681 5377
rect 8715 5343 8754 5377
rect 8788 5343 8827 5377
rect 8861 5343 8900 5377
rect 8934 5343 8973 5377
rect 9007 5343 9046 5377
rect 9080 5343 9119 5377
rect 9153 5343 9192 5377
rect 9226 5343 9265 5377
rect 9299 5343 9338 5377
rect 9372 5343 9411 5377
rect 9445 5343 9484 5377
rect 9518 5343 9557 5377
rect 9591 5343 9630 5377
rect 9664 5343 9703 5377
rect 9737 5343 9776 5377
rect 9810 5343 9849 5377
rect 9883 5343 9923 5377
rect 9957 5343 9995 5377
rect 10029 5343 10035 5377
rect 5037 5337 10035 5343
rect 5037 5306 5046 5337
tri 5046 5306 5077 5337 nw
tri 9883 5306 9914 5337 ne
rect 9914 5306 10035 5337
rect 5037 5304 5044 5306
tri 5044 5304 5046 5306 nw
tri 9914 5304 9916 5306 ne
rect 9916 5304 10035 5306
rect 5037 4114 5043 5304
tri 5043 5303 5044 5304 nw
tri 9916 5303 9917 5304 ne
rect 4925 4025 4931 4062
rect 5037 4025 5043 4062
rect 4925 3936 4931 3973
rect 5037 3936 5043 3973
rect 4925 3847 4931 3884
rect 5037 3847 5043 3884
rect 4925 3758 4931 3795
rect 5037 3758 5043 3795
rect 4925 3668 4931 3706
rect 5037 3668 5043 3706
rect 4925 3578 4931 3616
rect 5037 3578 5043 3616
rect 4977 3526 4991 3543
rect 4925 3504 5043 3526
rect 4925 3470 4931 3504
rect 4965 3470 5003 3504
rect 5037 3470 5043 3504
rect 4925 3431 5043 3470
rect 4925 3397 4931 3431
rect 4965 3397 5003 3431
rect 5037 3397 5043 3431
rect 4925 3358 5043 3397
rect 4925 3324 4931 3358
rect 4965 3324 5003 3358
rect 5037 3324 5043 3358
rect 4925 3285 5043 3324
rect 4925 3251 4931 3285
rect 4965 3251 5003 3285
rect 5037 3251 5043 3285
rect 5114 4114 5166 5280
rect 5114 4047 5166 4062
rect 5114 3980 5166 3995
rect 5114 3913 5166 3928
rect 5114 3846 5166 3861
rect 5114 3779 5166 3794
rect 5114 3712 5166 3727
rect 5114 3645 5166 3660
rect 5114 3578 5166 3593
rect 5114 3278 5166 3526
rect 5270 4854 5322 5280
rect 5270 4787 5322 4802
rect 5270 4720 5322 4735
rect 5270 4653 5322 4668
rect 5270 4586 5322 4601
rect 5270 4519 5322 4534
rect 5270 4452 5322 4467
rect 5270 4385 5322 4400
rect 5270 4318 5322 4333
rect 5270 3278 5322 4266
rect 5426 4114 5478 5280
rect 5426 4047 5478 4062
rect 5426 3980 5478 3995
rect 5426 3913 5478 3928
rect 5426 3846 5478 3861
rect 5426 3779 5478 3794
rect 5426 3712 5478 3727
rect 5426 3645 5478 3660
rect 5426 3578 5478 3593
rect 5426 3278 5478 3526
rect 5582 4854 5634 5280
rect 5582 4787 5634 4802
rect 5582 4720 5634 4735
rect 5582 4653 5634 4668
rect 5582 4586 5634 4601
rect 5582 4519 5634 4534
rect 5582 4452 5634 4467
rect 5582 4385 5634 4400
rect 5582 4318 5634 4333
rect 5582 3278 5634 4266
rect 5738 4114 5790 5280
rect 5738 4047 5790 4062
rect 5738 3980 5790 3995
rect 5738 3913 5790 3928
rect 5738 3846 5790 3861
rect 5738 3779 5790 3794
rect 5738 3712 5790 3727
rect 5738 3645 5790 3660
rect 5738 3578 5790 3593
rect 5738 3278 5790 3526
rect 5894 4854 5946 5280
rect 5894 4787 5946 4802
rect 5894 4720 5946 4735
rect 5894 4653 5946 4668
rect 5894 4586 5946 4601
rect 5894 4519 5946 4534
rect 5894 4452 5946 4467
rect 5894 4385 5946 4400
rect 5894 4318 5946 4333
rect 5894 3278 5946 4266
rect 6050 4114 6102 5280
rect 6050 4047 6102 4062
rect 6050 3980 6102 3995
rect 6050 3913 6102 3928
rect 6050 3846 6102 3861
rect 6050 3779 6102 3794
rect 6050 3712 6102 3727
rect 6050 3645 6102 3660
rect 6050 3578 6102 3593
rect 6050 3278 6102 3526
rect 6205 4854 6257 5280
rect 6205 4787 6257 4802
rect 6205 4720 6257 4735
rect 6205 4653 6257 4668
rect 6205 4586 6257 4601
rect 6205 4519 6257 4534
rect 6205 4452 6257 4467
rect 6205 4385 6257 4400
rect 6205 4318 6257 4333
rect 6205 3278 6257 4266
rect 6361 4114 6413 5280
rect 6361 4047 6413 4062
rect 6361 3980 6413 3995
rect 6361 3913 6413 3928
rect 6361 3846 6413 3861
rect 6361 3779 6413 3794
rect 6361 3712 6413 3727
rect 6361 3645 6413 3660
rect 6361 3578 6413 3593
rect 6361 3278 6413 3526
rect 6517 4854 6569 5280
rect 6517 4787 6569 4802
rect 6517 4720 6569 4735
rect 6517 4653 6569 4668
rect 6517 4586 6569 4601
rect 6517 4519 6569 4534
rect 6517 4452 6569 4467
rect 6517 4385 6569 4400
rect 6517 4318 6569 4333
rect 6517 3278 6569 4266
rect 6673 4114 6725 5280
rect 6673 4047 6725 4062
rect 6673 3980 6725 3995
rect 6673 3913 6725 3928
rect 6673 3846 6725 3861
rect 6673 3779 6725 3794
rect 6673 3712 6725 3727
rect 6673 3645 6725 3660
rect 6673 3578 6725 3593
rect 6673 3278 6725 3526
rect 6830 4854 6882 5280
rect 6830 4787 6882 4802
rect 6830 4720 6882 4735
rect 6830 4653 6882 4668
rect 6830 4586 6882 4601
rect 6830 4519 6882 4534
rect 6830 4452 6882 4467
rect 6830 4385 6882 4400
rect 6830 4318 6882 4333
rect 6830 3278 6882 4266
rect 6986 4114 7038 5280
rect 6986 4047 7038 4062
rect 6986 3980 7038 3995
rect 6986 3913 7038 3928
rect 6986 3846 7038 3861
rect 6986 3779 7038 3794
rect 6986 3712 7038 3727
rect 6986 3645 7038 3660
rect 6986 3578 7038 3593
rect 6986 3278 7038 3526
rect 7142 4854 7194 5280
rect 7142 4787 7194 4802
rect 7142 4720 7194 4735
rect 7142 4653 7194 4668
rect 7142 4586 7194 4601
rect 7142 4519 7194 4534
rect 7142 4452 7194 4467
rect 7142 4385 7194 4400
rect 7142 4318 7194 4333
rect 7142 3278 7194 4266
rect 7298 4114 7350 5280
rect 7298 4047 7350 4062
rect 7298 3980 7350 3995
rect 7298 3913 7350 3928
rect 7298 3846 7350 3861
rect 7298 3779 7350 3794
rect 7298 3712 7350 3727
rect 7298 3645 7350 3660
rect 7298 3578 7350 3593
rect 7298 3278 7350 3526
rect 7454 4854 7506 5280
rect 7454 4787 7506 4802
rect 7454 4720 7506 4735
rect 7454 4653 7506 4668
rect 7454 4586 7506 4601
rect 7454 4519 7506 4534
rect 7454 4452 7506 4467
rect 7454 4385 7506 4400
rect 7454 4318 7506 4333
rect 7454 3278 7506 4266
rect 7610 4114 7662 5280
rect 7610 4047 7662 4062
rect 7610 3980 7662 3995
rect 7610 3913 7662 3928
rect 7610 3846 7662 3861
rect 7610 3779 7662 3794
rect 7610 3712 7662 3727
rect 7610 3645 7662 3660
rect 7610 3578 7662 3593
rect 7610 3278 7662 3526
rect 7766 4854 7818 5280
rect 7766 4787 7818 4802
rect 7766 4720 7818 4735
rect 7766 4653 7818 4668
rect 7766 4586 7818 4601
rect 7766 4519 7818 4534
rect 7766 4452 7818 4467
rect 7766 4385 7818 4400
rect 7766 4318 7818 4333
rect 7766 3278 7818 4266
rect 7922 4114 7974 5280
rect 7922 4047 7974 4062
rect 7922 3980 7974 3995
rect 7922 3913 7974 3928
rect 7922 3846 7974 3861
rect 7922 3779 7974 3794
rect 7922 3712 7974 3727
rect 7922 3645 7974 3660
rect 7922 3578 7974 3593
rect 7922 3278 7974 3526
rect 8078 4854 8130 5280
rect 8078 4787 8130 4802
rect 8078 4720 8130 4735
rect 8078 4653 8130 4668
rect 8078 4586 8130 4601
rect 8078 4519 8130 4534
rect 8078 4452 8130 4467
rect 8078 4385 8130 4400
rect 8078 4318 8130 4333
rect 8078 3278 8130 4266
rect 8234 4114 8286 5280
rect 8234 4047 8286 4062
rect 8234 3980 8286 3995
rect 8234 3913 8286 3928
rect 8234 3846 8286 3861
rect 8234 3779 8286 3794
rect 8234 3712 8286 3727
rect 8234 3645 8286 3660
rect 8234 3578 8286 3593
rect 8234 3278 8286 3526
rect 8390 4854 8442 5280
rect 8390 4787 8442 4802
rect 8390 4720 8442 4735
rect 8390 4653 8442 4668
rect 8390 4586 8442 4601
rect 8390 4519 8442 4534
rect 8390 4452 8442 4467
rect 8390 4385 8442 4400
rect 8390 4318 8442 4333
rect 8390 3278 8442 4266
rect 8546 4114 8598 5280
rect 8546 4047 8598 4062
rect 8546 3980 8598 3995
rect 8546 3913 8598 3928
rect 8546 3846 8598 3861
rect 8546 3779 8598 3794
rect 8546 3712 8598 3727
rect 8546 3645 8598 3660
rect 8546 3578 8598 3593
rect 8546 3278 8598 3526
rect 8702 4854 8754 5280
rect 8702 4787 8754 4802
rect 8702 4720 8754 4735
rect 8702 4653 8754 4668
rect 8702 4586 8754 4601
rect 8702 4519 8754 4534
rect 8702 4452 8754 4467
rect 8702 4385 8754 4400
rect 8702 4318 8754 4333
rect 8702 3278 8754 4266
rect 8858 4114 8910 5280
rect 8858 4047 8910 4062
rect 8858 3980 8910 3995
rect 8858 3913 8910 3928
rect 8858 3846 8910 3861
rect 8858 3779 8910 3794
rect 8858 3712 8910 3727
rect 8858 3645 8910 3660
rect 8858 3578 8910 3593
rect 8858 3278 8910 3526
rect 9014 4854 9066 5280
rect 9014 4787 9066 4802
rect 9014 4720 9066 4735
rect 9014 4653 9066 4668
rect 9014 4586 9066 4601
rect 9014 4519 9066 4534
rect 9014 4452 9066 4467
rect 9014 4385 9066 4400
rect 9014 4318 9066 4333
rect 9014 3278 9066 4266
rect 9170 4114 9222 5280
rect 9170 4047 9222 4062
rect 9170 3980 9222 3995
rect 9170 3913 9222 3928
rect 9170 3846 9222 3861
rect 9170 3779 9222 3794
rect 9170 3712 9222 3727
rect 9170 3645 9222 3660
rect 9170 3578 9222 3593
rect 9170 3278 9222 3526
rect 9326 4854 9378 5280
rect 9326 4787 9378 4802
rect 9326 4720 9378 4735
rect 9326 4653 9378 4668
rect 9326 4586 9378 4601
rect 9326 4519 9378 4534
rect 9326 4452 9378 4467
rect 9326 4385 9378 4400
rect 9326 4318 9378 4333
rect 9326 3278 9378 4266
rect 9482 4114 9534 5280
rect 9482 4047 9534 4062
rect 9482 3980 9534 3995
rect 9482 3913 9534 3928
rect 9482 3846 9534 3861
rect 9482 3779 9534 3794
rect 9482 3712 9534 3727
rect 9482 3645 9534 3660
rect 9482 3578 9534 3593
rect 9482 3278 9534 3526
rect 9638 4854 9690 5280
rect 9638 4787 9690 4802
rect 9638 4720 9690 4735
rect 9638 4653 9690 4668
rect 9638 4586 9690 4601
rect 9638 4519 9690 4534
rect 9638 4452 9690 4467
rect 9638 4385 9690 4400
rect 9638 4318 9690 4333
rect 9638 3278 9690 4266
rect 9794 4114 9846 5280
rect 9794 4047 9846 4062
rect 9794 3980 9846 3995
rect 9794 3913 9846 3928
rect 9794 3846 9846 3861
rect 9794 3779 9846 3794
rect 9794 3712 9846 3727
rect 9794 3645 9846 3660
rect 9794 3578 9846 3593
rect 9794 3278 9846 3526
rect 9917 5270 9923 5304
rect 9957 5270 9995 5304
rect 10029 5270 10035 5304
rect 9917 5231 10035 5270
rect 9917 5197 9923 5231
rect 9957 5197 9995 5231
rect 10029 5197 10035 5231
rect 9917 5158 10035 5197
rect 9917 5124 9923 5158
rect 9957 5124 9995 5158
rect 10029 5124 10035 5158
rect 9917 5085 10035 5124
rect 9917 5051 9923 5085
rect 9957 5051 9995 5085
rect 10029 5051 10035 5085
rect 9917 5012 10035 5051
rect 9917 4978 9923 5012
rect 9957 4978 9995 5012
rect 10029 4978 10035 5012
rect 9917 4939 10035 4978
rect 9917 4905 9923 4939
rect 9957 4905 9995 4939
rect 10029 4905 10035 4939
rect 9917 4866 10035 4905
rect 9917 4832 9923 4866
rect 9957 4832 9995 4866
rect 10029 4832 10035 4866
rect 9917 4793 10035 4832
rect 9917 4759 9923 4793
rect 9957 4759 9995 4793
rect 10029 4759 10035 4793
rect 9917 4720 10035 4759
rect 9917 4686 9923 4720
rect 9957 4686 9995 4720
rect 10029 4686 10035 4720
rect 9917 4647 10035 4686
rect 9917 4613 9923 4647
rect 9957 4613 9995 4647
rect 10029 4613 10035 4647
rect 9917 4574 10035 4613
rect 9917 4540 9923 4574
rect 9957 4540 9995 4574
rect 10029 4540 10035 4574
rect 9917 4501 10035 4540
rect 9917 4467 9923 4501
rect 9957 4467 9995 4501
rect 10029 4467 10035 4501
rect 9917 4428 10035 4467
rect 9917 4394 9923 4428
rect 9957 4394 9995 4428
rect 10029 4394 10035 4428
rect 9917 4355 10035 4394
rect 9917 4321 9923 4355
rect 9957 4321 9995 4355
rect 10029 4321 10035 4355
rect 9917 4282 10035 4321
rect 9917 4248 9923 4282
rect 9957 4248 9995 4282
rect 10029 4248 10035 4282
rect 9917 4209 10035 4248
rect 9917 4175 9923 4209
rect 9957 4175 9995 4209
rect 10029 4175 10035 4209
rect 9917 4136 10035 4175
rect 9917 4114 9923 4136
rect 9957 4114 9995 4136
rect 10029 4114 10035 4136
rect 9969 4062 9983 4114
rect 9917 4029 9923 4062
rect 9957 4029 9995 4062
rect 10029 4029 10035 4062
rect 9917 4025 10035 4029
rect 9969 3973 9983 4025
rect 9917 3956 9923 3973
rect 9957 3956 9995 3973
rect 10029 3956 10035 3973
rect 9917 3936 10035 3956
rect 9969 3884 9983 3936
rect 9917 3883 9923 3884
rect 9957 3883 9995 3884
rect 10029 3883 10035 3884
rect 9917 3847 10035 3883
rect 9969 3795 9983 3847
rect 9917 3771 10035 3795
rect 9917 3758 9923 3771
rect 9957 3758 9995 3771
rect 10029 3758 10035 3771
rect 9969 3706 9983 3758
rect 9917 3698 10035 3706
rect 9917 3668 9923 3698
rect 9957 3668 9995 3698
rect 10029 3668 10035 3698
rect 9969 3616 9983 3668
rect 9917 3591 9923 3616
rect 9957 3591 9995 3616
rect 10029 3591 10035 3616
rect 9917 3578 10035 3591
rect 9969 3526 9983 3578
rect 9917 3518 9923 3526
rect 9957 3518 9995 3526
rect 10029 3518 10035 3526
rect 9917 3479 10035 3518
rect 9917 3445 9923 3479
rect 9957 3445 9995 3479
rect 10029 3445 10035 3479
rect 9917 3406 10035 3445
rect 9917 3372 9923 3406
rect 9957 3372 9995 3406
rect 10029 3372 10035 3406
rect 9917 3333 10035 3372
rect 9917 3299 9923 3333
rect 9957 3299 9995 3333
rect 10029 3299 10035 3333
rect 4925 3212 5043 3251
rect 9917 3260 10035 3299
rect 9917 3226 9923 3260
rect 9957 3226 9995 3260
rect 10029 3226 10035 3260
rect 4925 3178 4931 3212
rect 4965 3178 5003 3212
rect 5037 3178 5043 3212
rect 4925 3139 5043 3178
rect 5191 3216 5303 3225
rect 5355 3216 5367 3225
rect 5419 3216 5431 3225
rect 5483 3216 5495 3225
rect 5191 3182 5203 3216
rect 5237 3182 5275 3216
rect 5483 3182 5491 3216
rect 5191 3173 5303 3182
rect 5355 3173 5367 3182
rect 5419 3173 5431 3182
rect 5483 3173 5495 3182
rect 5547 3173 5559 3225
rect 5611 3173 5623 3225
rect 5675 3173 5687 3225
rect 5739 3216 5751 3225
rect 5803 3216 5815 3225
rect 5867 3216 5879 3225
rect 5931 3216 5943 3225
rect 5995 3216 6007 3225
rect 6059 3216 6071 3225
rect 5741 3182 5751 3216
rect 5813 3182 5815 3216
rect 6059 3182 6067 3216
rect 5739 3173 5751 3182
rect 5803 3173 5815 3182
rect 5867 3173 5879 3182
rect 5931 3173 5943 3182
rect 5995 3173 6007 3182
rect 6059 3173 6071 3182
rect 6123 3173 6135 3225
rect 6187 3173 6199 3225
rect 6251 3173 6263 3225
rect 6315 3216 6327 3225
rect 6379 3216 6391 3225
rect 6443 3216 6456 3225
rect 6508 3216 6521 3225
rect 6573 3216 6586 3225
rect 6638 3216 6651 3225
rect 6703 3216 6716 3225
rect 6317 3182 6327 3216
rect 6389 3182 6391 3216
rect 6638 3182 6643 3216
rect 6703 3182 6715 3216
rect 6315 3173 6327 3182
rect 6379 3173 6391 3182
rect 6443 3173 6456 3182
rect 6508 3173 6521 3182
rect 6573 3173 6586 3182
rect 6638 3173 6651 3182
rect 6703 3173 6716 3182
rect 6768 3173 6781 3225
rect 6833 3173 6846 3225
rect 6898 3173 6911 3225
rect 6963 3216 6976 3225
rect 7028 3216 7041 3225
rect 7093 3216 7106 3225
rect 7158 3216 7171 3225
rect 7223 3216 7236 3225
rect 7288 3216 7301 3225
rect 7353 3216 7366 3225
rect 6965 3182 6976 3216
rect 7037 3182 7041 3216
rect 7288 3182 7291 3216
rect 7353 3182 7363 3216
rect 6963 3173 6976 3182
rect 7028 3173 7041 3182
rect 7093 3173 7106 3182
rect 7158 3173 7171 3182
rect 7223 3173 7236 3182
rect 7288 3173 7301 3182
rect 7353 3173 7366 3182
rect 7418 3173 7431 3225
rect 7483 3173 7496 3225
rect 7548 3173 7561 3225
rect 7613 3173 7626 3225
rect 7678 3216 7691 3225
rect 7743 3216 7756 3225
rect 7808 3216 7821 3225
rect 7873 3216 7886 3225
rect 7938 3216 7951 3225
rect 8003 3216 8016 3225
rect 7685 3182 7691 3216
rect 7938 3182 7939 3216
rect 8003 3182 8011 3216
rect 7678 3173 7691 3182
rect 7743 3173 7756 3182
rect 7808 3173 7821 3182
rect 7873 3173 7886 3182
rect 7938 3173 7951 3182
rect 8003 3173 8016 3182
rect 8068 3173 8081 3225
rect 8133 3173 8146 3225
rect 8198 3173 8211 3225
rect 8263 3173 8276 3225
rect 8328 3216 8341 3225
rect 8393 3216 8406 3225
rect 8458 3216 8471 3225
rect 8523 3216 8536 3225
rect 8588 3216 8601 3225
rect 8653 3216 8666 3225
rect 8333 3182 8341 3216
rect 8405 3182 8406 3216
rect 8653 3182 8659 3216
rect 8328 3173 8341 3182
rect 8393 3173 8406 3182
rect 8458 3173 8471 3182
rect 8523 3173 8536 3182
rect 8588 3173 8601 3182
rect 8653 3173 8666 3182
rect 8718 3173 8731 3225
rect 8783 3173 8796 3225
rect 8848 3173 8861 3225
rect 8913 3173 8926 3225
rect 8978 3216 8991 3225
rect 9043 3216 9056 3225
rect 9108 3216 9121 3225
rect 9173 3216 9186 3225
rect 9238 3216 9251 3225
rect 9303 3216 9316 3225
rect 9368 3216 9381 3225
rect 8981 3182 8991 3216
rect 9053 3182 9056 3216
rect 9303 3182 9307 3216
rect 9368 3182 9379 3216
rect 8978 3173 8991 3182
rect 9043 3173 9056 3182
rect 9108 3173 9121 3182
rect 9173 3173 9186 3182
rect 9238 3173 9251 3182
rect 9303 3173 9316 3182
rect 9368 3173 9381 3182
rect 9433 3173 9446 3225
rect 9498 3216 9785 3225
rect 9498 3182 9523 3216
rect 9557 3182 9595 3216
rect 9629 3182 9667 3216
rect 9701 3182 9739 3216
rect 9773 3182 9785 3216
rect 9498 3173 9785 3182
rect 9917 3187 10035 3226
rect 4925 3105 4931 3139
rect 4965 3105 5003 3139
rect 5037 3105 5043 3139
rect 4925 3066 5043 3105
rect 4925 3032 4931 3066
rect 4965 3032 5003 3066
rect 5037 3043 5043 3066
rect 9917 3153 9923 3187
rect 9957 3153 9995 3187
rect 10029 3153 10035 3187
rect 9917 3114 10035 3153
rect 9917 3080 9923 3114
rect 9957 3080 9995 3114
rect 10029 3080 10035 3114
tri 5043 3043 5054 3054 sw
tri 9906 3043 9917 3054 se
rect 9917 3043 10035 3080
rect 5037 3041 5054 3043
tri 5054 3041 5056 3043 sw
tri 9904 3041 9906 3043 se
rect 9906 3041 10035 3043
rect 5037 3032 5056 3041
rect 4925 3020 5056 3032
tri 5056 3020 5077 3041 sw
tri 9883 3020 9904 3041 se
rect 9904 3020 9923 3041
rect 4925 3014 9923 3020
rect 4925 2993 5075 3014
rect 4925 2959 4931 2993
rect 4965 2959 5003 2993
rect 5037 2980 5075 2993
rect 5109 2980 5148 3014
rect 5182 2980 5221 3014
rect 5255 2980 5294 3014
rect 5328 2980 5367 3014
rect 5401 2980 5440 3014
rect 5474 2980 5513 3014
rect 5547 2980 5586 3014
rect 5620 2980 5659 3014
rect 5693 2980 5732 3014
rect 5766 2980 5805 3014
rect 5839 2980 5878 3014
rect 5912 2980 5951 3014
rect 5985 2980 6024 3014
rect 6058 2980 6097 3014
rect 6131 2980 6170 3014
rect 6204 2980 6243 3014
rect 6277 2980 6316 3014
rect 6350 2980 6389 3014
rect 6423 2980 6462 3014
rect 6496 2980 6535 3014
rect 6569 2980 6608 3014
rect 6642 2980 6681 3014
rect 6715 2980 6754 3014
rect 6788 2980 6827 3014
rect 5037 2959 6827 2980
rect 4925 2942 6827 2959
rect 4925 2920 5075 2942
rect 4925 2886 4931 2920
rect 4965 2886 5003 2920
rect 5037 2908 5075 2920
rect 5109 2908 5148 2942
rect 5182 2908 5221 2942
rect 5255 2908 5294 2942
rect 5328 2908 5367 2942
rect 5401 2908 5440 2942
rect 5474 2908 5513 2942
rect 5547 2908 5586 2942
rect 5620 2908 5659 2942
rect 5693 2908 5732 2942
rect 5766 2908 5805 2942
rect 5839 2908 5878 2942
rect 5912 2908 5951 2942
rect 5985 2908 6024 2942
rect 6058 2908 6097 2942
rect 6131 2908 6170 2942
rect 6204 2908 6243 2942
rect 6277 2908 6316 2942
rect 6350 2908 6389 2942
rect 6423 2908 6462 2942
rect 6496 2908 6535 2942
rect 6569 2908 6608 2942
rect 6642 2908 6681 2942
rect 6715 2908 6754 2942
rect 6788 2908 6827 2942
rect 9885 3007 9923 3014
rect 9957 3007 9995 3041
rect 10029 3007 10035 3041
rect 9885 2968 10035 3007
rect 9885 2934 9923 2968
rect 9957 2934 9995 2968
rect 10029 2934 10035 2968
rect 9885 2908 10035 2934
rect 5037 2902 10035 2908
rect 5037 2897 5072 2902
tri 5072 2897 5077 2902 nw
tri 9883 2897 9888 2902 ne
rect 9888 2897 10035 2902
rect 5037 2895 5070 2897
tri 5070 2895 5072 2897 nw
tri 9888 2895 9890 2897 ne
rect 9890 2895 10035 2897
rect 5037 2886 5043 2895
rect 4925 2847 5043 2886
tri 5043 2868 5070 2895 nw
tri 9890 2868 9917 2895 ne
rect 4925 2813 4931 2847
rect 4965 2813 5003 2847
rect 5037 2813 5043 2847
rect 4925 2774 5043 2813
rect 4925 2740 4931 2774
rect 4965 2740 5003 2774
rect 5037 2740 5043 2774
rect 9917 2861 9923 2895
rect 9957 2861 9995 2895
rect 10029 2861 10035 2895
rect 9917 2822 10035 2861
rect 9917 2788 9923 2822
rect 9957 2788 9995 2822
rect 10029 2788 10035 2822
rect 4925 2701 5043 2740
rect 5191 2746 5303 2755
rect 5355 2746 5367 2755
rect 5419 2746 5431 2755
rect 5483 2746 5495 2755
rect 5191 2712 5203 2746
rect 5237 2712 5275 2746
rect 5483 2712 5491 2746
rect 5191 2703 5303 2712
rect 5355 2703 5367 2712
rect 5419 2703 5431 2712
rect 5483 2703 5495 2712
rect 5547 2703 5559 2755
rect 5611 2703 5623 2755
rect 5675 2703 5687 2755
rect 5739 2746 5751 2755
rect 5803 2746 5815 2755
rect 5867 2746 5879 2755
rect 5931 2746 5943 2755
rect 5995 2746 6007 2755
rect 6059 2746 6071 2755
rect 5741 2712 5751 2746
rect 5813 2712 5815 2746
rect 6059 2712 6067 2746
rect 5739 2703 5751 2712
rect 5803 2703 5815 2712
rect 5867 2703 5879 2712
rect 5931 2703 5943 2712
rect 5995 2703 6007 2712
rect 6059 2703 6071 2712
rect 6123 2703 6135 2755
rect 6187 2703 6199 2755
rect 6251 2703 6263 2755
rect 6315 2746 6327 2755
rect 6379 2746 6391 2755
rect 6443 2746 6456 2755
rect 6508 2746 6521 2755
rect 6573 2746 6586 2755
rect 6638 2746 6651 2755
rect 6703 2746 6716 2755
rect 6317 2712 6327 2746
rect 6389 2712 6391 2746
rect 6638 2712 6643 2746
rect 6703 2712 6715 2746
rect 6315 2703 6327 2712
rect 6379 2703 6391 2712
rect 6443 2703 6456 2712
rect 6508 2703 6521 2712
rect 6573 2703 6586 2712
rect 6638 2703 6651 2712
rect 6703 2703 6716 2712
rect 6768 2703 6781 2755
rect 6833 2703 6846 2755
rect 6898 2703 6911 2755
rect 6963 2746 6976 2755
rect 7028 2746 7041 2755
rect 7093 2746 7106 2755
rect 7158 2746 7171 2755
rect 7223 2746 7236 2755
rect 7288 2746 7301 2755
rect 7353 2746 7366 2755
rect 6965 2712 6976 2746
rect 7037 2712 7041 2746
rect 7288 2712 7291 2746
rect 7353 2712 7363 2746
rect 6963 2703 6976 2712
rect 7028 2703 7041 2712
rect 7093 2703 7106 2712
rect 7158 2703 7171 2712
rect 7223 2703 7236 2712
rect 7288 2703 7301 2712
rect 7353 2703 7366 2712
rect 7418 2703 7431 2755
rect 7483 2703 7496 2755
rect 7548 2703 7561 2755
rect 7613 2703 7626 2755
rect 7678 2746 7691 2755
rect 7743 2746 7756 2755
rect 7808 2746 7821 2755
rect 7873 2746 7886 2755
rect 7938 2746 7951 2755
rect 8003 2746 8016 2755
rect 7685 2712 7691 2746
rect 7938 2712 7939 2746
rect 8003 2712 8011 2746
rect 7678 2703 7691 2712
rect 7743 2703 7756 2712
rect 7808 2703 7821 2712
rect 7873 2703 7886 2712
rect 7938 2703 7951 2712
rect 8003 2703 8016 2712
rect 8068 2703 8081 2755
rect 8133 2703 8146 2755
rect 8198 2703 8211 2755
rect 8263 2703 8276 2755
rect 8328 2746 8341 2755
rect 8393 2746 8406 2755
rect 8458 2746 8471 2755
rect 8523 2746 8536 2755
rect 8588 2746 8601 2755
rect 8653 2746 8666 2755
rect 8333 2712 8341 2746
rect 8405 2712 8406 2746
rect 8653 2712 8659 2746
rect 8328 2703 8341 2712
rect 8393 2703 8406 2712
rect 8458 2703 8471 2712
rect 8523 2703 8536 2712
rect 8588 2703 8601 2712
rect 8653 2703 8666 2712
rect 8718 2703 8731 2755
rect 8783 2703 8796 2755
rect 8848 2703 8861 2755
rect 8913 2703 8926 2755
rect 8978 2746 8991 2755
rect 9043 2746 9056 2755
rect 9108 2746 9121 2755
rect 9173 2746 9186 2755
rect 9238 2746 9251 2755
rect 9303 2746 9316 2755
rect 9368 2746 9381 2755
rect 8981 2712 8991 2746
rect 9053 2712 9056 2746
rect 9303 2712 9307 2746
rect 9368 2712 9379 2746
rect 8978 2703 8991 2712
rect 9043 2703 9056 2712
rect 9108 2703 9121 2712
rect 9173 2703 9186 2712
rect 9238 2703 9251 2712
rect 9303 2703 9316 2712
rect 9368 2703 9381 2712
rect 9433 2703 9446 2755
rect 9498 2746 9785 2755
rect 9498 2712 9523 2746
rect 9557 2712 9595 2746
rect 9629 2712 9667 2746
rect 9701 2712 9739 2746
rect 9773 2712 9785 2746
rect 9498 2703 9785 2712
rect 9917 2749 10035 2788
rect 9917 2715 9923 2749
rect 9957 2715 9995 2749
rect 10029 2715 10035 2749
rect 4925 2667 4931 2701
rect 4965 2667 5003 2701
rect 5037 2667 5043 2701
rect 4925 2628 5043 2667
rect 9917 2676 10035 2715
rect 4925 2604 4931 2628
rect 4965 2604 5003 2628
rect 5037 2604 5043 2628
rect 4977 2552 4991 2604
rect 4925 2522 4931 2552
rect 4965 2522 5003 2552
rect 5037 2522 5043 2552
rect 4977 2470 4991 2522
rect 4925 2448 4931 2470
rect 4965 2448 5003 2470
rect 5037 2448 5043 2470
rect 4925 2440 5043 2448
rect 4977 2388 4991 2440
rect 4925 2375 4931 2388
rect 4965 2375 5003 2388
rect 5037 2375 5043 2388
rect 4925 2357 5043 2375
rect 4977 2305 4991 2357
rect 4925 2302 4931 2305
rect 4965 2302 5003 2305
rect 5037 2302 5043 2305
rect 4925 2274 5043 2302
rect 4977 2222 4991 2274
rect 4925 2191 5043 2222
rect 4977 2139 4991 2191
rect 4925 2117 5043 2139
rect 4925 2108 4931 2117
rect 4965 2108 5003 2117
rect 5037 2108 5043 2117
rect 4977 2056 4991 2108
rect 4925 2044 5043 2056
rect 4925 2010 4931 2044
rect 4965 2010 5003 2044
rect 5037 2010 5043 2044
rect 4925 1971 5043 2010
rect 4925 1937 4931 1971
rect 4965 1937 5003 1971
rect 5037 1937 5043 1971
rect 4925 1898 5043 1937
rect 4925 1864 4931 1898
rect 4965 1864 5003 1898
rect 5037 1864 5043 1898
rect 4925 1825 5043 1864
rect 4925 1791 4931 1825
rect 4965 1791 5003 1825
rect 5037 1791 5043 1825
rect 4925 1752 5043 1791
rect 4925 1718 4931 1752
rect 4965 1718 5003 1752
rect 5037 1718 5043 1752
rect 4925 1679 5043 1718
rect 4925 1645 4931 1679
rect 4965 1645 5003 1679
rect 5037 1645 5043 1679
rect 4925 1606 5043 1645
rect 4925 1572 4931 1606
rect 4965 1572 5003 1606
rect 5037 1572 5043 1606
rect 4925 1533 5043 1572
rect 4925 1499 4931 1533
rect 4965 1499 5003 1533
rect 5037 1499 5043 1533
rect 4925 1460 5043 1499
rect 4925 1426 4931 1460
rect 4965 1426 5003 1460
rect 5037 1426 5043 1460
rect 4925 1387 5043 1426
rect 4925 1353 4931 1387
rect 4965 1353 5003 1387
rect 5037 1353 5043 1387
rect 4925 1314 5043 1353
rect 4925 1280 4931 1314
rect 4965 1280 5003 1314
rect 5037 1280 5043 1314
rect 4925 1241 5043 1280
rect 4925 1207 4931 1241
rect 4965 1207 5003 1241
rect 5037 1207 5043 1241
rect 4925 1168 5043 1207
rect 4925 1134 4931 1168
rect 4965 1134 5003 1168
rect 5037 1134 5043 1168
rect 4925 1095 5043 1134
rect 4925 1061 4931 1095
rect 4965 1061 5003 1095
rect 5037 1061 5043 1095
rect 4925 1022 5043 1061
rect 4925 988 4931 1022
rect 4965 988 5003 1022
rect 5037 988 5043 1022
rect 4925 949 5043 988
rect 4925 915 4931 949
rect 4965 915 5003 949
rect 5037 915 5043 949
rect 4925 876 5043 915
rect 4925 842 4931 876
rect 4965 842 5003 876
rect 5037 842 5043 876
rect 4925 803 5043 842
rect 4925 769 4931 803
rect 4965 769 5003 803
rect 5037 769 5043 803
rect 4925 730 5043 769
rect 4925 696 4931 730
rect 4965 696 5003 730
rect 5037 696 5043 730
rect 4925 657 5043 696
rect 4925 623 4931 657
rect 4965 623 5003 657
rect 5037 623 5043 657
rect 5114 2604 5166 2650
rect 5114 2537 5166 2552
rect 5114 2470 5166 2485
rect 5114 2403 5166 2418
rect 5114 2336 5166 2351
rect 5114 2269 5166 2284
rect 5114 2202 5166 2217
rect 5114 2135 5166 2150
rect 5114 2068 5166 2083
rect 5114 648 5166 2016
rect 5270 1865 5322 2650
rect 5270 1798 5322 1813
rect 5270 1731 5322 1746
rect 5270 1664 5322 1679
rect 5270 1597 5322 1612
rect 5270 1530 5322 1545
rect 5270 1463 5322 1478
rect 5270 1396 5322 1411
rect 5270 1329 5322 1344
rect 5270 648 5322 1277
rect 5426 2604 5478 2650
rect 5426 2537 5478 2552
rect 5426 2470 5478 2485
rect 5426 2403 5478 2418
rect 5426 2336 5478 2351
rect 5426 2269 5478 2284
rect 5426 2202 5478 2217
rect 5426 2135 5478 2150
rect 5426 2068 5478 2083
rect 5426 648 5478 2016
rect 5582 1865 5634 2650
rect 5582 1798 5634 1813
rect 5582 1731 5634 1746
rect 5582 1664 5634 1679
rect 5582 1597 5634 1612
rect 5582 1530 5634 1545
rect 5582 1463 5634 1478
rect 5582 1396 5634 1411
rect 5582 1329 5634 1344
rect 5582 648 5634 1277
rect 5738 2604 5790 2650
rect 5738 2537 5790 2552
rect 5738 2470 5790 2485
rect 5738 2403 5790 2418
rect 5738 2336 5790 2351
rect 5738 2269 5790 2284
rect 5738 2202 5790 2217
rect 5738 2135 5790 2150
rect 5738 2068 5790 2083
rect 5738 648 5790 2016
rect 5894 1865 5946 2650
rect 5894 1798 5946 1813
rect 5894 1731 5946 1746
rect 5894 1664 5946 1679
rect 5894 1597 5946 1612
rect 5894 1530 5946 1545
rect 5894 1463 5946 1478
rect 5894 1396 5946 1411
rect 5894 1329 5946 1344
rect 5894 648 5946 1277
rect 6050 2604 6102 2650
rect 6050 2537 6102 2552
rect 6050 2470 6102 2485
rect 6050 2403 6102 2418
rect 6050 2336 6102 2351
rect 6050 2269 6102 2284
rect 6050 2202 6102 2217
rect 6050 2135 6102 2150
rect 6050 2068 6102 2083
rect 6050 648 6102 2016
rect 6205 1865 6257 2650
rect 6205 1798 6257 1813
rect 6205 1731 6257 1746
rect 6205 1664 6257 1679
rect 6205 1597 6257 1612
rect 6205 1530 6257 1545
rect 6205 1463 6257 1478
rect 6205 1396 6257 1411
rect 6205 1329 6257 1344
rect 6205 648 6257 1277
rect 6361 2604 6413 2650
rect 6361 2537 6413 2552
rect 6361 2470 6413 2485
rect 6361 2403 6413 2418
rect 6361 2336 6413 2351
rect 6361 2269 6413 2284
rect 6361 2202 6413 2217
rect 6361 2135 6413 2150
rect 6361 2068 6413 2083
rect 6361 648 6413 2016
rect 6517 1865 6569 2650
rect 6517 1798 6569 1813
rect 6517 1731 6569 1746
rect 6517 1664 6569 1679
rect 6517 1597 6569 1612
rect 6517 1530 6569 1545
rect 6517 1463 6569 1478
rect 6517 1396 6569 1411
rect 6517 1329 6569 1344
rect 6517 648 6569 1277
rect 6673 2604 6725 2650
rect 6673 2537 6725 2552
rect 6673 2470 6725 2485
rect 6673 2403 6725 2418
rect 6673 2336 6725 2351
rect 6673 2269 6725 2284
rect 6673 2202 6725 2217
rect 6673 2135 6725 2150
rect 6673 2068 6725 2083
rect 6673 648 6725 2016
rect 6830 1865 6882 2650
rect 6830 1798 6882 1813
rect 6830 1731 6882 1746
rect 6830 1664 6882 1679
rect 6830 1597 6882 1612
rect 6830 1530 6882 1545
rect 6830 1463 6882 1478
rect 6830 1396 6882 1411
rect 6830 1329 6882 1344
rect 6830 648 6882 1277
rect 6986 2604 7038 2650
rect 6986 2537 7038 2552
rect 6986 2470 7038 2485
rect 6986 2403 7038 2418
rect 6986 2336 7038 2351
rect 6986 2269 7038 2284
rect 6986 2202 7038 2217
rect 6986 2135 7038 2150
rect 6986 2068 7038 2083
rect 6986 648 7038 2016
rect 7142 1865 7194 2650
rect 7142 1798 7194 1813
rect 7142 1731 7194 1746
rect 7142 1664 7194 1679
rect 7142 1597 7194 1612
rect 7142 1530 7194 1545
rect 7142 1463 7194 1478
rect 7142 1396 7194 1411
rect 7142 1329 7194 1344
rect 7142 648 7194 1277
rect 7298 2604 7350 2650
rect 7298 2537 7350 2552
rect 7298 2470 7350 2485
rect 7298 2403 7350 2418
rect 7298 2336 7350 2351
rect 7298 2269 7350 2284
rect 7298 2202 7350 2217
rect 7298 2135 7350 2150
rect 7298 2068 7350 2083
rect 7298 648 7350 2016
rect 7454 1865 7506 2650
rect 7454 1798 7506 1813
rect 7454 1731 7506 1746
rect 7454 1664 7506 1679
rect 7454 1597 7506 1612
rect 7454 1530 7506 1545
rect 7454 1463 7506 1478
rect 7454 1396 7506 1411
rect 7454 1329 7506 1344
rect 7454 648 7506 1277
rect 7610 2604 7662 2650
rect 7610 2537 7662 2552
rect 7610 2470 7662 2485
rect 7610 2403 7662 2418
rect 7610 2336 7662 2351
rect 7610 2269 7662 2284
rect 7610 2202 7662 2217
rect 7610 2135 7662 2150
rect 7610 2068 7662 2083
rect 7610 648 7662 2016
rect 7766 1865 7818 2650
rect 7766 1798 7818 1813
rect 7766 1731 7818 1746
rect 7766 1664 7818 1679
rect 7766 1597 7818 1612
rect 7766 1530 7818 1545
rect 7766 1463 7818 1478
rect 7766 1396 7818 1411
rect 7766 1329 7818 1344
rect 7766 648 7818 1277
rect 7922 2604 7974 2650
rect 7922 2537 7974 2552
rect 7922 2470 7974 2485
rect 7922 2403 7974 2418
rect 7922 2336 7974 2351
rect 7922 2269 7974 2284
rect 7922 2202 7974 2217
rect 7922 2135 7974 2150
rect 7922 2068 7974 2083
rect 7922 648 7974 2016
rect 8078 1865 8130 2650
rect 8078 1798 8130 1813
rect 8078 1731 8130 1746
rect 8078 1664 8130 1679
rect 8078 1597 8130 1612
rect 8078 1530 8130 1545
rect 8078 1463 8130 1478
rect 8078 1396 8130 1411
rect 8078 1329 8130 1344
rect 8078 648 8130 1277
rect 8234 2604 8286 2650
rect 8234 2537 8286 2552
rect 8234 2470 8286 2485
rect 8234 2403 8286 2418
rect 8234 2336 8286 2351
rect 8234 2269 8286 2284
rect 8234 2202 8286 2217
rect 8234 2135 8286 2150
rect 8234 2068 8286 2083
rect 8234 648 8286 2016
rect 8390 1865 8442 2650
rect 8390 1798 8442 1813
rect 8390 1731 8442 1746
rect 8390 1664 8442 1679
rect 8390 1597 8442 1612
rect 8390 1530 8442 1545
rect 8390 1463 8442 1478
rect 8390 1396 8442 1411
rect 8390 1329 8442 1344
rect 8390 648 8442 1277
rect 8546 2604 8598 2650
rect 8546 2537 8598 2552
rect 8546 2470 8598 2485
rect 8546 2403 8598 2418
rect 8546 2336 8598 2351
rect 8546 2269 8598 2284
rect 8546 2202 8598 2217
rect 8546 2135 8598 2150
rect 8546 2068 8598 2083
rect 8546 648 8598 2016
rect 8702 1865 8754 2650
rect 8702 1798 8754 1813
rect 8702 1731 8754 1746
rect 8702 1664 8754 1679
rect 8702 1597 8754 1612
rect 8702 1530 8754 1545
rect 8702 1463 8754 1478
rect 8702 1396 8754 1411
rect 8702 1329 8754 1344
rect 8702 648 8754 1277
rect 8858 2604 8910 2650
rect 8858 2537 8910 2552
rect 8858 2470 8910 2485
rect 8858 2403 8910 2418
rect 8858 2336 8910 2351
rect 8858 2269 8910 2284
rect 8858 2202 8910 2217
rect 8858 2135 8910 2150
rect 8858 2068 8910 2083
rect 8858 648 8910 2016
rect 9014 1865 9066 2650
rect 9014 1798 9066 1813
rect 9014 1731 9066 1746
rect 9014 1664 9066 1679
rect 9014 1597 9066 1612
rect 9014 1530 9066 1545
rect 9014 1463 9066 1478
rect 9014 1396 9066 1411
rect 9014 1329 9066 1344
rect 9014 648 9066 1277
rect 9170 2604 9222 2650
rect 9170 2537 9222 2552
rect 9170 2470 9222 2485
rect 9170 2403 9222 2418
rect 9170 2336 9222 2351
rect 9170 2269 9222 2284
rect 9170 2202 9222 2217
rect 9170 2135 9222 2150
rect 9170 2068 9222 2083
rect 9170 648 9222 2016
rect 9326 1865 9378 2650
rect 9326 1798 9378 1813
rect 9326 1731 9378 1746
rect 9326 1664 9378 1679
rect 9326 1597 9378 1612
rect 9326 1530 9378 1545
rect 9326 1463 9378 1478
rect 9326 1396 9378 1411
rect 9326 1329 9378 1344
rect 9326 648 9378 1277
rect 9482 2604 9534 2650
rect 9482 2537 9534 2552
rect 9482 2470 9534 2485
rect 9482 2403 9534 2418
rect 9482 2336 9534 2351
rect 9482 2269 9534 2284
rect 9482 2202 9534 2217
rect 9482 2135 9534 2150
rect 9482 2068 9534 2083
rect 9482 648 9534 2016
rect 9638 1865 9690 2650
rect 9638 1798 9690 1813
rect 9638 1731 9690 1746
rect 9638 1664 9690 1679
rect 9638 1597 9690 1612
rect 9638 1530 9690 1545
rect 9638 1463 9690 1478
rect 9638 1396 9690 1411
rect 9638 1329 9690 1344
rect 9638 648 9690 1277
rect 9794 2604 9846 2650
rect 9794 2537 9846 2552
rect 9794 2470 9846 2485
rect 9794 2403 9846 2418
rect 9794 2336 9846 2351
rect 9794 2269 9846 2284
rect 9794 2202 9846 2217
rect 9794 2135 9846 2150
rect 9794 2068 9846 2083
rect 9794 648 9846 2016
rect 9917 2642 9923 2676
rect 9957 2642 9995 2676
rect 10029 2642 10035 2676
rect 9917 2604 10035 2642
rect 9969 2552 9983 2604
rect 9917 2530 10035 2552
rect 9917 2522 9923 2530
rect 9957 2522 9995 2530
rect 10029 2522 10035 2530
rect 9969 2470 9983 2522
rect 9917 2457 10035 2470
rect 9917 2440 9923 2457
rect 9957 2440 9995 2457
rect 10029 2440 10035 2457
rect 9969 2388 9983 2440
rect 9917 2384 10035 2388
rect 9917 2357 9923 2384
rect 10029 2357 10035 2384
rect 9917 2274 9923 2305
rect 10029 2274 10035 2305
rect 9917 2191 9923 2222
rect 10029 2191 10035 2222
rect 9917 2108 9923 2139
rect 10029 2108 10035 2139
rect 4925 590 5043 623
tri 5043 590 5077 624 sw
tri 9883 590 9917 624 se
rect 9917 590 9923 2056
rect 4925 584 9923 590
rect 4925 550 4931 584
rect 4965 550 5003 584
rect 4925 478 5003 550
rect 8205 550 8244 584
rect 8278 550 8317 584
rect 8351 550 8390 584
rect 8424 550 8463 584
rect 8497 550 8536 584
rect 8570 550 8609 584
rect 8643 550 8682 584
rect 8716 550 8755 584
rect 8789 550 8828 584
rect 8862 550 8901 584
rect 8935 550 8974 584
rect 9008 550 9047 584
rect 9081 550 9120 584
rect 9154 550 9193 584
rect 9227 550 9266 584
rect 9300 550 9339 584
rect 9373 550 9412 584
rect 9446 550 9485 584
rect 9519 550 9558 584
rect 9592 550 9631 584
rect 9665 550 9704 584
rect 9738 550 9777 584
rect 9811 550 9850 584
rect 9884 550 9923 584
rect 10029 550 10035 2056
rect 8205 512 10035 550
rect 8205 478 8244 512
rect 8278 478 8317 512
rect 8351 478 8390 512
rect 8424 478 8463 512
rect 8497 478 8536 512
rect 8570 478 8609 512
rect 8643 478 8682 512
rect 8716 478 8755 512
rect 8789 478 8828 512
rect 8862 478 8901 512
rect 8935 478 8974 512
rect 9008 478 9047 512
rect 9081 478 9120 512
rect 9154 478 9193 512
rect 9227 478 9266 512
rect 9300 478 9339 512
rect 9373 478 9412 512
rect 9446 478 9485 512
rect 9519 478 9558 512
rect 9592 478 9631 512
rect 9665 478 9704 512
rect 9738 478 9777 512
rect 9811 478 9850 512
rect 9884 478 9923 512
rect 9957 478 10035 512
rect 4925 472 10035 478
rect 10271 5452 10389 5491
rect 10271 5418 10277 5452
rect 10311 5418 10349 5452
rect 10383 5418 10389 5452
rect 10271 5379 10389 5418
rect 10271 5345 10277 5379
rect 10311 5345 10349 5379
rect 10383 5345 10389 5379
rect 10271 5306 10389 5345
rect 10271 5272 10277 5306
rect 10311 5272 10349 5306
rect 10383 5272 10389 5306
rect 10271 5233 10389 5272
rect 10271 5199 10277 5233
rect 10311 5199 10349 5233
rect 10383 5199 10389 5233
rect 10271 5160 10389 5199
rect 10271 5126 10277 5160
rect 10311 5126 10349 5160
rect 10383 5126 10389 5160
rect 10271 5087 10389 5126
rect 10271 5053 10277 5087
rect 10311 5053 10349 5087
rect 10383 5053 10389 5087
rect 10271 5014 10389 5053
rect 10271 4980 10277 5014
rect 10311 4980 10349 5014
rect 10383 4980 10389 5014
rect 10271 4941 10389 4980
rect 10271 4907 10277 4941
rect 10311 4907 10349 4941
rect 10383 4907 10389 4941
rect 10271 4868 10389 4907
rect 10271 4834 10277 4868
rect 10311 4834 10349 4868
rect 10383 4834 10389 4868
rect 10271 4795 10389 4834
rect 10271 4761 10277 4795
rect 10311 4761 10349 4795
rect 10383 4761 10389 4795
rect 10271 4722 10389 4761
rect 10271 4688 10277 4722
rect 10311 4688 10349 4722
rect 10383 4688 10389 4722
rect 10271 4649 10389 4688
rect 10271 4615 10277 4649
rect 10311 4615 10349 4649
rect 10383 4615 10389 4649
rect 10271 4576 10389 4615
rect 10271 4542 10277 4576
rect 10311 4542 10349 4576
rect 10383 4542 10389 4576
rect 10271 4503 10389 4542
rect 10271 4469 10277 4503
rect 10311 4469 10349 4503
rect 10383 4469 10389 4503
rect 10271 4430 10389 4469
rect 10271 4396 10277 4430
rect 10311 4396 10349 4430
rect 10383 4396 10389 4430
rect 10271 4357 10389 4396
rect 10271 4323 10277 4357
rect 10311 4323 10349 4357
rect 10383 4323 10389 4357
rect 10271 4284 10389 4323
rect 10271 4250 10277 4284
rect 10311 4250 10349 4284
rect 10383 4250 10389 4284
rect 10271 4211 10389 4250
rect 10271 4177 10277 4211
rect 10311 4177 10349 4211
rect 10383 4177 10389 4211
rect 10271 4138 10389 4177
rect 10271 4104 10277 4138
rect 10311 4104 10349 4138
rect 10383 4104 10389 4138
rect 10271 4065 10389 4104
rect 10271 4031 10277 4065
rect 10311 4031 10349 4065
rect 10383 4031 10389 4065
rect 10271 3992 10389 4031
rect 10271 3958 10277 3992
rect 10311 3958 10349 3992
rect 10383 3958 10389 3992
rect 10271 3919 10389 3958
rect 10271 3885 10277 3919
rect 10311 3885 10349 3919
rect 10383 3885 10389 3919
rect 10271 3846 10389 3885
rect 10271 3812 10277 3846
rect 10311 3812 10349 3846
rect 10383 3812 10389 3846
rect 10271 3773 10389 3812
rect 10271 3739 10277 3773
rect 10311 3739 10349 3773
rect 10383 3739 10389 3773
rect 10271 3700 10389 3739
rect 10271 3666 10277 3700
rect 10311 3666 10349 3700
rect 10383 3666 10389 3700
rect 10271 3627 10389 3666
rect 10271 3593 10277 3627
rect 10311 3593 10349 3627
rect 10383 3593 10389 3627
rect 10271 3554 10389 3593
rect 10271 3520 10277 3554
rect 10311 3520 10349 3554
rect 10383 3520 10389 3554
rect 10271 3481 10389 3520
rect 10271 3447 10277 3481
rect 10311 3447 10349 3481
rect 10383 3447 10389 3481
rect 10271 3408 10389 3447
rect 10271 3374 10277 3408
rect 10311 3374 10349 3408
rect 10383 3374 10389 3408
rect 10271 3335 10389 3374
rect 10271 3301 10277 3335
rect 10311 3301 10349 3335
rect 10383 3301 10389 3335
rect 10271 3262 10389 3301
rect 10271 3228 10277 3262
rect 10311 3228 10349 3262
rect 10383 3228 10389 3262
rect 10271 3189 10389 3228
rect 10271 3155 10277 3189
rect 10311 3155 10349 3189
rect 10383 3155 10389 3189
rect 10271 3116 10389 3155
rect 10271 3082 10277 3116
rect 10311 3082 10349 3116
rect 10383 3082 10389 3116
rect 10271 3043 10389 3082
rect 10271 3009 10277 3043
rect 10311 3009 10349 3043
rect 10383 3009 10389 3043
rect 10271 2970 10389 3009
rect 10271 2936 10277 2970
rect 10311 2936 10349 2970
rect 10383 2936 10389 2970
rect 10271 2897 10389 2936
rect 10271 2863 10277 2897
rect 10311 2863 10349 2897
rect 10383 2863 10389 2897
rect 10271 2824 10389 2863
rect 10271 2790 10277 2824
rect 10311 2790 10349 2824
rect 10383 2790 10389 2824
rect 10271 2751 10389 2790
rect 10271 2717 10277 2751
rect 10311 2717 10349 2751
rect 10383 2717 10389 2751
rect 10271 2678 10389 2717
rect 10271 2644 10277 2678
rect 10311 2644 10349 2678
rect 10383 2644 10389 2678
rect 10271 2605 10389 2644
rect 10271 2571 10277 2605
rect 10311 2571 10349 2605
rect 10383 2571 10389 2605
rect 10271 2532 10389 2571
rect 10271 2498 10277 2532
rect 10311 2498 10349 2532
rect 10383 2498 10389 2532
rect 10271 2459 10389 2498
rect 10271 2425 10277 2459
rect 10311 2425 10349 2459
rect 10383 2425 10389 2459
rect 10271 2386 10389 2425
rect 10271 2352 10277 2386
rect 10311 2352 10349 2386
rect 10383 2352 10389 2386
rect 10271 2313 10389 2352
rect 10271 2279 10277 2313
rect 10311 2279 10349 2313
rect 10383 2279 10389 2313
rect 10271 2240 10389 2279
rect 10271 2206 10277 2240
rect 10311 2206 10349 2240
rect 10383 2206 10389 2240
rect 10271 2167 10389 2206
rect 10271 2133 10277 2167
rect 10311 2133 10349 2167
rect 10383 2133 10389 2167
rect 10271 2094 10389 2133
rect 10271 2060 10277 2094
rect 10311 2060 10349 2094
rect 10383 2060 10389 2094
rect 10271 2021 10389 2060
rect 10271 1987 10277 2021
rect 10311 1987 10349 2021
rect 10383 1987 10389 2021
rect 10271 1948 10389 1987
rect 10271 1914 10277 1948
rect 10311 1914 10349 1948
rect 10383 1914 10389 1948
rect 10271 1875 10389 1914
rect 10271 1841 10277 1875
rect 10311 1841 10349 1875
rect 10383 1841 10389 1875
rect 10271 1802 10389 1841
tri 4776 224 4810 258 sw
tri 10237 224 10271 258 se
rect 10271 224 10277 1802
rect 4770 218 10277 224
rect -30 184 -24 218
rect 10 184 48 218
rect -30 112 48 184
rect 9946 184 9985 218
rect 10019 184 10058 218
rect 10092 184 10131 218
rect 10165 184 10204 218
rect 10238 184 10277 218
rect 10383 184 10389 1802
rect 9946 146 10389 184
rect 9946 112 9985 146
rect 10019 112 10058 146
rect 10092 112 10131 146
rect 10165 112 10204 146
rect 10238 112 10277 146
rect 10311 112 10389 146
rect -30 106 10389 112
<< via1 >>
rect -16 5770 36 5822
rect 48 5816 100 5822
rect 48 5782 82 5816
rect 82 5782 100 5816
rect 48 5770 100 5782
rect 112 5816 164 5822
rect 112 5782 121 5816
rect 121 5782 155 5816
rect 155 5782 164 5816
rect 112 5770 164 5782
rect 176 5816 228 5822
rect 176 5782 194 5816
rect 194 5782 228 5816
rect 176 5770 228 5782
rect 240 5816 292 5822
rect 304 5816 356 5822
rect 368 5816 420 5822
rect 432 5816 484 5822
rect 496 5816 548 5822
rect 560 5816 612 5822
rect 240 5782 267 5816
rect 267 5782 292 5816
rect 304 5782 340 5816
rect 340 5782 356 5816
rect 368 5782 374 5816
rect 374 5782 413 5816
rect 413 5782 420 5816
rect 432 5782 447 5816
rect 447 5782 484 5816
rect 496 5782 520 5816
rect 520 5782 548 5816
rect 560 5782 593 5816
rect 593 5782 612 5816
rect 240 5770 292 5782
rect 304 5770 356 5782
rect 368 5770 420 5782
rect 432 5770 484 5782
rect 496 5770 548 5782
rect 560 5770 612 5782
rect 624 5816 676 5822
rect 624 5782 632 5816
rect 632 5782 666 5816
rect 666 5782 676 5816
rect 624 5770 676 5782
rect 688 5816 740 5822
rect 688 5782 705 5816
rect 705 5782 739 5816
rect 739 5782 740 5816
rect 688 5770 740 5782
rect 752 5816 804 5822
rect 816 5816 868 5822
rect 880 5816 932 5822
rect 944 5816 996 5822
rect 1008 5816 1060 5822
rect 1072 5816 1124 5822
rect 752 5782 778 5816
rect 778 5782 804 5816
rect 816 5782 851 5816
rect 851 5782 868 5816
rect 880 5782 885 5816
rect 885 5782 924 5816
rect 924 5782 932 5816
rect 944 5782 958 5816
rect 958 5782 996 5816
rect 1008 5782 1031 5816
rect 1031 5782 1060 5816
rect 1072 5782 1104 5816
rect 1104 5782 1124 5816
rect 752 5770 804 5782
rect 816 5770 868 5782
rect 880 5770 932 5782
rect 944 5770 996 5782
rect 1008 5770 1060 5782
rect 1072 5770 1124 5782
rect 1136 5816 1188 5822
rect 1136 5782 1143 5816
rect 1143 5782 1177 5816
rect 1177 5782 1188 5816
rect 1136 5770 1188 5782
rect 1200 5816 1252 5822
rect 1264 5816 1316 5822
rect 1328 5816 1380 5822
rect 1392 5816 1444 5822
rect 1456 5816 1508 5822
rect 1520 5816 1572 5822
rect 1584 5816 1636 5822
rect 1648 5816 1700 5822
rect 1712 5816 1764 5822
rect 1776 5816 1828 5822
rect 1840 5816 1892 5822
rect 1904 5816 1956 5822
rect 1968 5816 2020 5822
rect 2032 5816 2084 5822
rect 2096 5816 2148 5822
rect 2160 5816 2212 5822
rect 2224 5816 2276 5822
rect 2288 5816 2340 5822
rect 2352 5816 2404 5822
rect 2416 5816 2468 5822
rect 2480 5816 2532 5822
rect 2544 5816 2596 5822
rect 2608 5816 2660 5822
rect 2672 5816 2724 5822
rect 2736 5816 2788 5822
rect 2800 5816 2852 5822
rect 2864 5816 2916 5822
rect 2928 5816 2980 5822
rect 2992 5816 3044 5822
rect 3056 5816 3108 5822
rect 3120 5816 3172 5822
rect 3184 5816 3236 5822
rect 3248 5816 3300 5822
rect 3312 5816 3364 5822
rect 3376 5816 3428 5822
rect 3440 5816 3492 5822
rect 3504 5816 3556 5822
rect 3568 5816 3620 5822
rect 3632 5816 3684 5822
rect 3696 5816 3748 5822
rect 3760 5816 3812 5822
rect 3824 5816 3876 5822
rect 3888 5816 3940 5822
rect 3952 5816 4004 5822
rect 4016 5816 4068 5822
rect 4080 5816 4132 5822
rect 4144 5816 4196 5822
rect 4208 5816 4260 5822
rect 4272 5816 4324 5822
rect 4336 5816 4388 5822
rect 4400 5816 4452 5822
rect 4464 5816 4516 5822
rect 4528 5816 4580 5822
rect 4592 5816 4644 5822
rect 4656 5816 4708 5822
rect 4720 5816 4772 5822
rect 4784 5816 4836 5822
rect 4848 5816 4900 5822
rect 4912 5816 4964 5822
rect 4976 5816 5028 5822
rect 5040 5816 5092 5822
rect 5104 5816 5156 5822
rect 5168 5816 5220 5822
rect 5232 5816 5284 5822
rect 5296 5816 5348 5822
rect 5360 5816 5412 5822
rect 5424 5816 5476 5822
rect 5488 5816 5540 5822
rect 5552 5816 5604 5822
rect 5616 5816 5668 5822
rect 5680 5816 5732 5822
rect 5744 5816 5796 5822
rect 5808 5816 5860 5822
rect 5872 5816 5924 5822
rect 5936 5816 5988 5822
rect 6000 5816 6052 5822
rect 6064 5816 6116 5822
rect 6128 5816 6180 5822
rect 6192 5816 6244 5822
rect 6256 5816 6308 5822
rect 6320 5816 6372 5822
rect 6384 5816 6436 5822
rect 6448 5816 6500 5822
rect 6512 5816 6564 5822
rect 6576 5816 6628 5822
rect 6640 5816 6692 5822
rect 6704 5816 6756 5822
rect 6768 5816 6820 5822
rect 6832 5816 6884 5822
rect 6896 5816 6948 5822
rect 6960 5816 7012 5822
rect 7024 5816 7076 5822
rect 7088 5816 7140 5822
rect 7152 5816 7204 5822
rect 7216 5816 7268 5822
rect 7280 5816 7332 5822
rect 7344 5816 7396 5822
rect 7408 5816 7460 5822
rect 7472 5816 7524 5822
rect 7536 5816 7588 5822
rect 7600 5816 7652 5822
rect 7664 5816 7716 5822
rect 7728 5816 7780 5822
rect 7792 5816 7844 5822
rect 7856 5816 7908 5822
rect 7920 5816 7972 5822
rect 7984 5816 8036 5822
rect 8048 5816 8100 5822
rect 8112 5816 8164 5822
rect 8176 5816 8228 5822
rect 8240 5816 8292 5822
rect 8304 5816 8356 5822
rect 8368 5816 8420 5822
rect 8432 5816 8484 5822
rect 8496 5816 8548 5822
rect 8560 5816 8612 5822
rect 8624 5816 8676 5822
rect 8688 5816 8740 5822
rect 8752 5816 8804 5822
rect 8816 5816 8868 5822
rect 8880 5816 8932 5822
rect 8944 5816 8996 5822
rect 9008 5816 9060 5822
rect 9072 5816 9124 5822
rect 9136 5816 9188 5822
rect 9200 5816 9252 5822
rect 9264 5816 9316 5822
rect 9329 5816 9381 5822
rect 9394 5816 9446 5822
rect 1200 5770 1216 5816
rect 1216 5770 1252 5816
rect 1264 5770 1316 5816
rect 1328 5770 1380 5816
rect 1392 5770 1444 5816
rect 1456 5770 1508 5816
rect 1520 5770 1572 5816
rect 1584 5770 1636 5816
rect 1648 5770 1700 5816
rect 1712 5770 1764 5816
rect 1776 5770 1828 5816
rect 1840 5770 1892 5816
rect 1904 5770 1956 5816
rect 1968 5770 2020 5816
rect 2032 5770 2084 5816
rect 2096 5770 2148 5816
rect 2160 5770 2212 5816
rect 2224 5770 2276 5816
rect 2288 5770 2340 5816
rect 2352 5770 2404 5816
rect 2416 5770 2468 5816
rect 2480 5770 2532 5816
rect 2544 5770 2596 5816
rect 2608 5770 2660 5816
rect 2672 5770 2724 5816
rect 2736 5770 2788 5816
rect 2800 5770 2852 5816
rect 2864 5770 2916 5816
rect 2928 5770 2980 5816
rect 2992 5770 3044 5816
rect 3056 5770 3108 5816
rect 3120 5770 3172 5816
rect 3184 5770 3236 5816
rect 3248 5770 3300 5816
rect 3312 5770 3364 5816
rect 3376 5770 3428 5816
rect 3440 5770 3492 5816
rect 3504 5770 3556 5816
rect 3568 5770 3620 5816
rect 3632 5770 3684 5816
rect 3696 5770 3748 5816
rect 3760 5770 3812 5816
rect 3824 5770 3876 5816
rect 3888 5770 3940 5816
rect 3952 5770 4004 5816
rect 4016 5770 4068 5816
rect 4080 5770 4132 5816
rect 4144 5770 4196 5816
rect 4208 5770 4260 5816
rect 4272 5770 4324 5816
rect 4336 5770 4388 5816
rect 4400 5770 4452 5816
rect 4464 5770 4516 5816
rect 4528 5770 4580 5816
rect 4592 5770 4644 5816
rect 4656 5770 4708 5816
rect 4720 5770 4772 5816
rect 4784 5770 4836 5816
rect 4848 5770 4900 5816
rect 4912 5770 4964 5816
rect 4976 5770 5028 5816
rect 5040 5770 5092 5816
rect 5104 5770 5156 5816
rect 5168 5770 5220 5816
rect 5232 5770 5284 5816
rect 5296 5770 5348 5816
rect 5360 5770 5412 5816
rect 5424 5770 5476 5816
rect 5488 5770 5540 5816
rect 5552 5770 5604 5816
rect 5616 5770 5668 5816
rect 5680 5770 5732 5816
rect 5744 5770 5796 5816
rect 5808 5770 5860 5816
rect 5872 5770 5924 5816
rect 5936 5770 5988 5816
rect 6000 5770 6052 5816
rect 6064 5770 6116 5816
rect 6128 5770 6180 5816
rect 6192 5770 6244 5816
rect 6256 5770 6308 5816
rect 6320 5770 6372 5816
rect 6384 5770 6436 5816
rect 6448 5770 6500 5816
rect 6512 5770 6564 5816
rect 6576 5770 6628 5816
rect 6640 5770 6692 5816
rect 6704 5770 6756 5816
rect 6768 5770 6820 5816
rect 6832 5770 6884 5816
rect 6896 5770 6948 5816
rect 6960 5770 7012 5816
rect 7024 5770 7076 5816
rect 7088 5770 7140 5816
rect 7152 5770 7204 5816
rect 7216 5770 7268 5816
rect 7280 5770 7332 5816
rect 7344 5770 7396 5816
rect 7408 5770 7460 5816
rect 7472 5770 7524 5816
rect 7536 5770 7588 5816
rect 7600 5770 7652 5816
rect 7664 5770 7716 5816
rect 7728 5770 7780 5816
rect 7792 5770 7844 5816
rect 7856 5770 7908 5816
rect 7920 5770 7972 5816
rect 7984 5770 8036 5816
rect 8048 5770 8100 5816
rect 8112 5770 8164 5816
rect 8176 5770 8228 5816
rect 8240 5770 8292 5816
rect 8304 5770 8356 5816
rect 8368 5770 8420 5816
rect 8432 5770 8484 5816
rect 8496 5770 8548 5816
rect 8560 5770 8612 5816
rect 8624 5770 8676 5816
rect 8688 5770 8740 5816
rect 8752 5770 8804 5816
rect 8816 5770 8868 5816
rect 8880 5770 8932 5816
rect 8944 5770 8996 5816
rect 9008 5770 9060 5816
rect 9072 5770 9124 5816
rect 9136 5770 9188 5816
rect 9200 5770 9252 5816
rect 9264 5770 9316 5816
rect 9329 5770 9381 5816
rect 9394 5770 9446 5816
rect 9459 5770 9511 5822
rect 9524 5816 9576 5822
rect 9524 5782 9534 5816
rect 9534 5782 9568 5816
rect 9568 5782 9576 5816
rect 9524 5770 9576 5782
rect 9589 5816 9641 5822
rect 9654 5816 9706 5822
rect 9719 5816 9771 5822
rect 9784 5816 9836 5822
rect 9849 5816 9901 5822
rect 9914 5816 9966 5822
rect 9589 5782 9609 5816
rect 9609 5782 9641 5816
rect 9654 5782 9683 5816
rect 9683 5782 9706 5816
rect 9719 5782 9757 5816
rect 9757 5782 9771 5816
rect 9784 5782 9791 5816
rect 9791 5782 9831 5816
rect 9831 5782 9836 5816
rect 9849 5782 9865 5816
rect 9865 5782 9901 5816
rect 9914 5782 9939 5816
rect 9939 5782 9966 5816
rect 9589 5770 9641 5782
rect 9654 5770 9706 5782
rect 9719 5770 9771 5782
rect 9784 5770 9836 5782
rect 9849 5770 9901 5782
rect 9914 5770 9966 5782
rect 9979 5816 10031 5822
rect 9979 5782 10013 5816
rect 10013 5782 10031 5816
rect 9979 5770 10031 5782
rect 10044 5816 10096 5822
rect 10044 5782 10053 5816
rect 10053 5782 10087 5816
rect 10087 5782 10096 5816
rect 10044 5770 10096 5782
rect 10109 5816 10161 5822
rect 10109 5782 10127 5816
rect 10127 5782 10161 5816
rect 10109 5770 10161 5782
rect 10174 5816 10226 5822
rect 10239 5816 10291 5822
rect 10174 5782 10201 5816
rect 10201 5782 10226 5816
rect 10239 5782 10275 5816
rect 10275 5782 10291 5816
rect 10174 5770 10226 5782
rect 10239 5770 10291 5782
rect -16 5744 36 5756
rect 48 5744 100 5756
rect -16 5704 36 5744
rect 48 5704 82 5744
rect 82 5704 100 5744
rect 112 5744 164 5756
rect 112 5710 121 5744
rect 121 5710 155 5744
rect 155 5710 164 5744
rect 112 5704 164 5710
rect 176 5744 228 5756
rect 176 5710 194 5744
rect 194 5710 228 5744
rect 176 5704 228 5710
rect 240 5744 292 5756
rect 304 5744 356 5756
rect 368 5744 420 5756
rect 432 5744 484 5756
rect 496 5744 548 5756
rect 560 5744 612 5756
rect 240 5710 267 5744
rect 267 5710 292 5744
rect 304 5710 340 5744
rect 340 5710 356 5744
rect 368 5710 374 5744
rect 374 5710 413 5744
rect 413 5710 420 5744
rect 432 5710 447 5744
rect 447 5710 484 5744
rect 496 5710 520 5744
rect 520 5710 548 5744
rect 560 5710 593 5744
rect 593 5710 612 5744
rect 240 5704 292 5710
rect 304 5704 356 5710
rect 368 5704 420 5710
rect 432 5704 484 5710
rect 496 5704 548 5710
rect 560 5704 612 5710
rect 624 5744 676 5756
rect 624 5710 632 5744
rect 632 5710 666 5744
rect 666 5710 676 5744
rect 624 5704 676 5710
rect 688 5744 740 5756
rect 688 5710 705 5744
rect 705 5710 739 5744
rect 739 5710 740 5744
rect 688 5704 740 5710
rect 752 5744 804 5756
rect 816 5744 868 5756
rect 880 5744 932 5756
rect 944 5744 996 5756
rect 1008 5744 1060 5756
rect 1072 5744 1124 5756
rect 752 5710 778 5744
rect 778 5710 804 5744
rect 816 5710 851 5744
rect 851 5710 868 5744
rect 880 5710 885 5744
rect 885 5710 924 5744
rect 924 5710 932 5744
rect 944 5710 958 5744
rect 958 5710 996 5744
rect 1008 5710 1031 5744
rect 1031 5710 1060 5744
rect 1072 5710 1104 5744
rect 1104 5710 1124 5744
rect 752 5704 804 5710
rect 816 5704 868 5710
rect 880 5704 932 5710
rect 944 5704 996 5710
rect 1008 5704 1060 5710
rect 1072 5704 1124 5710
rect 1136 5744 1188 5756
rect 1136 5710 1143 5744
rect 1143 5710 1177 5744
rect 1177 5710 1188 5744
rect 1136 5704 1188 5710
rect 1200 5710 1216 5756
rect 1216 5710 1252 5756
rect 1264 5710 1316 5756
rect 1328 5710 1380 5756
rect 1392 5710 1444 5756
rect 1456 5710 1508 5756
rect 1520 5710 1572 5756
rect 1584 5710 1636 5756
rect 1648 5710 1700 5756
rect 1712 5710 1764 5756
rect 1776 5710 1828 5756
rect 1840 5710 1892 5756
rect 1904 5710 1956 5756
rect 1968 5710 2020 5756
rect 2032 5710 2084 5756
rect 2096 5710 2148 5756
rect 2160 5710 2212 5756
rect 2224 5710 2276 5756
rect 2288 5710 2340 5756
rect 2352 5710 2404 5756
rect 2416 5710 2468 5756
rect 2480 5710 2532 5756
rect 2544 5710 2596 5756
rect 2608 5710 2660 5756
rect 2672 5710 2724 5756
rect 2736 5710 2788 5756
rect 2800 5710 2852 5756
rect 2864 5710 2916 5756
rect 2928 5710 2980 5756
rect 2992 5710 3044 5756
rect 3056 5710 3108 5756
rect 3120 5710 3172 5756
rect 3184 5710 3236 5756
rect 3248 5710 3300 5756
rect 3312 5710 3364 5756
rect 3376 5710 3428 5756
rect 3440 5710 3492 5756
rect 1200 5704 1252 5710
rect 1264 5704 1316 5710
rect 1328 5704 1380 5710
rect 1392 5704 1444 5710
rect 1456 5704 1508 5710
rect 1520 5704 1572 5710
rect 1584 5704 1636 5710
rect 1648 5704 1700 5710
rect 1712 5704 1764 5710
rect 1776 5704 1828 5710
rect 1840 5704 1892 5710
rect 1904 5704 1956 5710
rect 1968 5704 2020 5710
rect 2032 5704 2084 5710
rect 2096 5704 2148 5710
rect 2160 5704 2212 5710
rect 2224 5704 2276 5710
rect 2288 5704 2340 5710
rect 2352 5704 2404 5710
rect 2416 5704 2468 5710
rect 2480 5704 2532 5710
rect 2544 5704 2596 5710
rect 2608 5704 2660 5710
rect 2672 5704 2724 5710
rect 2736 5704 2788 5710
rect 2800 5704 2852 5710
rect 2864 5704 2916 5710
rect 2928 5704 2980 5710
rect 2992 5704 3044 5710
rect 3056 5704 3108 5710
rect 3120 5704 3172 5710
rect 3184 5704 3236 5710
rect 3248 5704 3300 5710
rect 3312 5704 3364 5710
rect 3376 5704 3428 5710
rect 3440 5704 3469 5710
rect 3469 5704 3492 5710
rect 3504 5704 3556 5756
rect 3568 5704 3620 5756
rect 3632 5710 3684 5756
rect 3696 5710 3748 5756
rect 3760 5710 3812 5756
rect 3824 5710 3876 5756
rect 3888 5710 3940 5756
rect 3952 5710 4004 5756
rect 4016 5710 4068 5756
rect 4080 5710 4132 5756
rect 4144 5710 4196 5756
rect 4208 5710 4260 5756
rect 4272 5710 4324 5756
rect 4336 5710 4388 5756
rect 4400 5710 4452 5756
rect 4464 5710 4516 5756
rect 4528 5710 4580 5756
rect 3632 5704 3647 5710
rect 3647 5704 3684 5710
rect 3696 5704 3748 5710
rect 3760 5704 3812 5710
rect 3824 5704 3876 5710
rect 3888 5704 3940 5710
rect 3952 5704 4004 5710
rect 4016 5704 4068 5710
rect 4080 5704 4132 5710
rect 4144 5704 4196 5710
rect 4208 5704 4260 5710
rect 4272 5704 4324 5710
rect 4336 5704 4388 5710
rect 4400 5704 4452 5710
rect 4464 5704 4516 5710
rect 4528 5704 4580 5710
rect 4592 5704 4644 5756
rect 4656 5704 4708 5756
rect 4720 5710 4772 5756
rect 4784 5710 4836 5756
rect 4848 5710 4900 5756
rect 4912 5710 4964 5756
rect 4976 5710 5028 5756
rect 5040 5710 5092 5756
rect 5104 5710 5156 5756
rect 5168 5710 5220 5756
rect 5232 5710 5284 5756
rect 5296 5710 5348 5756
rect 5360 5710 5412 5756
rect 5424 5710 5476 5756
rect 5488 5710 5540 5756
rect 5552 5710 5604 5756
rect 5616 5710 5668 5756
rect 5680 5710 5732 5756
rect 5744 5710 5796 5756
rect 5808 5710 5860 5756
rect 5872 5710 5924 5756
rect 5936 5710 5988 5756
rect 6000 5710 6052 5756
rect 6064 5710 6116 5756
rect 6128 5710 6180 5756
rect 6192 5710 6244 5756
rect 6256 5710 6308 5756
rect 6320 5710 6372 5756
rect 6384 5710 6436 5756
rect 6448 5710 6500 5756
rect 6512 5710 6564 5756
rect 6576 5710 6628 5756
rect 6640 5710 6692 5756
rect 6704 5710 6756 5756
rect 6768 5710 6820 5756
rect 6832 5710 6884 5756
rect 6896 5710 6948 5756
rect 6960 5710 7012 5756
rect 7024 5710 7076 5756
rect 7088 5710 7140 5756
rect 7152 5710 7204 5756
rect 7216 5710 7268 5756
rect 7280 5710 7332 5756
rect 7344 5710 7396 5756
rect 7408 5710 7460 5756
rect 7472 5710 7524 5756
rect 7536 5710 7588 5756
rect 7600 5710 7652 5756
rect 7664 5710 7716 5756
rect 7728 5710 7780 5756
rect 7792 5710 7844 5756
rect 7856 5710 7908 5756
rect 7920 5710 7972 5756
rect 7984 5710 8036 5756
rect 8048 5710 8100 5756
rect 8112 5710 8164 5756
rect 8176 5710 8228 5756
rect 8240 5710 8292 5756
rect 8304 5710 8356 5756
rect 8368 5710 8420 5756
rect 8432 5710 8484 5756
rect 8496 5710 8548 5756
rect 8560 5710 8612 5756
rect 8624 5710 8676 5756
rect 8688 5710 8740 5756
rect 8752 5710 8804 5756
rect 8816 5710 8868 5756
rect 8880 5710 8932 5756
rect 8944 5710 8996 5756
rect 9008 5710 9060 5756
rect 9072 5710 9124 5756
rect 9136 5710 9188 5756
rect 9200 5710 9252 5756
rect 9264 5710 9316 5756
rect 9329 5710 9381 5756
rect 9394 5710 9446 5756
rect 4720 5704 4770 5710
rect 4770 5704 4772 5710
rect 4784 5704 4836 5710
rect 4848 5704 4900 5710
rect 4912 5704 4964 5710
rect 4976 5704 5028 5710
rect 5040 5704 5092 5710
rect 5104 5704 5156 5710
rect 5168 5704 5220 5710
rect 5232 5704 5284 5710
rect 5296 5704 5348 5710
rect 5360 5704 5412 5710
rect 5424 5704 5476 5710
rect 5488 5704 5540 5710
rect 5552 5704 5604 5710
rect 5616 5704 5668 5710
rect 5680 5704 5732 5710
rect 5744 5704 5796 5710
rect 5808 5704 5860 5710
rect 5872 5704 5924 5710
rect 5936 5704 5988 5710
rect 6000 5704 6052 5710
rect 6064 5704 6116 5710
rect 6128 5704 6180 5710
rect 6192 5704 6244 5710
rect 6256 5704 6308 5710
rect 6320 5704 6372 5710
rect 6384 5704 6436 5710
rect 6448 5704 6500 5710
rect 6512 5704 6564 5710
rect 6576 5704 6628 5710
rect 6640 5704 6692 5710
rect 6704 5704 6756 5710
rect 6768 5704 6820 5710
rect 6832 5704 6884 5710
rect 6896 5704 6948 5710
rect 6960 5704 7012 5710
rect 7024 5704 7076 5710
rect 7088 5704 7140 5710
rect 7152 5704 7204 5710
rect 7216 5704 7268 5710
rect 7280 5704 7332 5710
rect 7344 5704 7396 5710
rect 7408 5704 7460 5710
rect 7472 5704 7524 5710
rect 7536 5704 7588 5710
rect 7600 5704 7652 5710
rect 7664 5704 7716 5710
rect 7728 5704 7780 5710
rect 7792 5704 7844 5710
rect 7856 5704 7908 5710
rect 7920 5704 7972 5710
rect 7984 5704 8036 5710
rect 8048 5704 8100 5710
rect 8112 5704 8164 5710
rect 8176 5704 8228 5710
rect 8240 5704 8292 5710
rect 8304 5704 8356 5710
rect 8368 5704 8420 5710
rect 8432 5704 8484 5710
rect 8496 5704 8548 5710
rect 8560 5704 8612 5710
rect 8624 5704 8676 5710
rect 8688 5704 8740 5710
rect 8752 5704 8804 5710
rect 8816 5704 8868 5710
rect 8880 5704 8932 5710
rect 8944 5704 8996 5710
rect 9008 5704 9060 5710
rect 9072 5704 9124 5710
rect 9136 5704 9188 5710
rect 9200 5704 9252 5710
rect 9264 5704 9316 5710
rect 9329 5704 9381 5710
rect 9394 5704 9446 5710
rect 9459 5704 9511 5756
rect 9524 5744 9576 5756
rect 9524 5710 9534 5744
rect 9534 5710 9568 5744
rect 9568 5710 9576 5744
rect 9524 5704 9576 5710
rect 9589 5744 9641 5756
rect 9654 5744 9706 5756
rect 9719 5744 9771 5756
rect 9784 5744 9836 5756
rect 9849 5744 9901 5756
rect 9914 5744 9966 5756
rect 9589 5710 9609 5744
rect 9609 5710 9641 5744
rect 9654 5710 9683 5744
rect 9683 5710 9706 5744
rect 9719 5710 9757 5744
rect 9757 5710 9771 5744
rect 9784 5710 9791 5744
rect 9791 5710 9831 5744
rect 9831 5710 9836 5744
rect 9849 5710 9865 5744
rect 9865 5710 9901 5744
rect 9914 5710 9939 5744
rect 9939 5710 9966 5744
rect 9589 5704 9641 5710
rect 9654 5704 9706 5710
rect 9719 5704 9771 5710
rect 9784 5704 9836 5710
rect 9849 5704 9901 5710
rect 9914 5704 9966 5710
rect 9979 5744 10031 5756
rect 9979 5710 10013 5744
rect 10013 5710 10031 5744
rect 9979 5704 10031 5710
rect 10044 5744 10096 5756
rect 10044 5710 10053 5744
rect 10053 5710 10087 5744
rect 10087 5710 10096 5744
rect 10044 5704 10096 5710
rect 10109 5744 10161 5756
rect 10109 5710 10127 5744
rect 10127 5710 10161 5744
rect 10109 5704 10161 5710
rect 10174 5744 10226 5756
rect 10239 5744 10291 5756
rect 10174 5710 10201 5744
rect 10201 5710 10226 5744
rect 10239 5710 10277 5744
rect 10277 5710 10291 5744
rect 10174 5704 10226 5710
rect 10239 5704 10291 5710
rect 525 5228 577 5280
rect 658 5274 710 5280
rect 791 5274 843 5280
rect 923 5274 975 5280
rect 1055 5274 1107 5280
rect 1187 5274 1239 5280
rect 1319 5274 1371 5280
rect 1451 5274 1503 5280
rect 1583 5274 1635 5280
rect 1715 5274 1767 5280
rect 1847 5274 1899 5280
rect 1979 5274 2031 5280
rect 2111 5274 2163 5280
rect 2243 5274 2295 5280
rect 2375 5274 2427 5280
rect 2507 5274 2559 5280
rect 2639 5274 2691 5280
rect 2771 5274 2823 5280
rect 2903 5274 2955 5280
rect 658 5240 675 5274
rect 675 5240 709 5274
rect 709 5240 710 5274
rect 791 5240 825 5274
rect 825 5240 843 5274
rect 923 5240 934 5274
rect 934 5240 975 5274
rect 1055 5240 1086 5274
rect 1086 5240 1107 5274
rect 1187 5240 1204 5274
rect 1204 5240 1238 5274
rect 1238 5240 1239 5274
rect 1319 5240 1356 5274
rect 1356 5240 1371 5274
rect 1451 5240 1466 5274
rect 1466 5240 1503 5274
rect 1583 5240 1584 5274
rect 1584 5240 1618 5274
rect 1618 5240 1635 5274
rect 1715 5240 1736 5274
rect 1736 5240 1767 5274
rect 1847 5240 1880 5274
rect 1880 5240 1899 5274
rect 1979 5240 1996 5274
rect 1996 5240 2030 5274
rect 2030 5240 2031 5274
rect 2111 5240 2146 5274
rect 2146 5240 2163 5274
rect 2243 5240 2255 5274
rect 2255 5240 2295 5274
rect 2375 5240 2407 5274
rect 2407 5240 2427 5274
rect 2507 5240 2525 5274
rect 2525 5240 2559 5274
rect 2639 5240 2677 5274
rect 2677 5240 2691 5274
rect 2771 5240 2787 5274
rect 2787 5240 2823 5274
rect 2903 5240 2905 5274
rect 2905 5240 2939 5274
rect 2939 5240 2955 5274
rect 658 5228 710 5240
rect 791 5228 843 5240
rect 923 5228 975 5240
rect 1055 5228 1107 5240
rect 1187 5228 1239 5240
rect 1319 5228 1371 5240
rect 1451 5228 1503 5240
rect 1583 5228 1635 5240
rect 1715 5228 1767 5240
rect 1847 5228 1899 5240
rect 1979 5228 2031 5240
rect 2111 5228 2163 5240
rect 2243 5228 2295 5240
rect 2375 5228 2427 5240
rect 2507 5228 2559 5240
rect 2639 5228 2691 5240
rect 2771 5228 2823 5240
rect 2903 5228 2955 5240
rect 3035 5228 3087 5280
rect 525 5202 577 5214
rect 658 5202 710 5214
rect 791 5202 843 5214
rect 923 5202 975 5214
rect 1055 5202 1107 5214
rect 1187 5202 1239 5214
rect 1319 5202 1371 5214
rect 1451 5202 1503 5214
rect 1583 5202 1635 5214
rect 1715 5202 1767 5214
rect 1847 5202 1899 5214
rect 1979 5202 2031 5214
rect 2111 5202 2163 5214
rect 2243 5202 2295 5214
rect 2375 5202 2427 5214
rect 2507 5202 2559 5214
rect 2639 5202 2691 5214
rect 2771 5202 2823 5214
rect 2903 5202 2955 5214
rect 3035 5202 3087 5214
rect 525 5168 559 5202
rect 559 5168 577 5202
rect 658 5168 675 5202
rect 675 5168 709 5202
rect 709 5168 710 5202
rect 791 5168 825 5202
rect 825 5168 843 5202
rect 923 5168 934 5202
rect 934 5168 975 5202
rect 1055 5168 1086 5202
rect 1086 5168 1107 5202
rect 1187 5168 1204 5202
rect 1204 5168 1238 5202
rect 1238 5168 1239 5202
rect 1319 5168 1356 5202
rect 1356 5168 1371 5202
rect 1451 5168 1466 5202
rect 1466 5168 1503 5202
rect 1583 5168 1584 5202
rect 1584 5168 1618 5202
rect 1618 5168 1635 5202
rect 1715 5168 1736 5202
rect 1736 5168 1767 5202
rect 1847 5168 1880 5202
rect 1880 5168 1899 5202
rect 1979 5168 1996 5202
rect 1996 5168 2030 5202
rect 2030 5168 2031 5202
rect 2111 5168 2146 5202
rect 2146 5168 2163 5202
rect 2243 5168 2255 5202
rect 2255 5168 2295 5202
rect 2375 5168 2407 5202
rect 2407 5168 2427 5202
rect 2507 5168 2525 5202
rect 2525 5168 2559 5202
rect 2639 5168 2677 5202
rect 2677 5168 2691 5202
rect 2771 5168 2787 5202
rect 2787 5168 2823 5202
rect 2903 5168 2905 5202
rect 2905 5168 2939 5202
rect 2939 5168 2955 5202
rect 525 5162 577 5168
rect 658 5162 710 5168
rect 791 5162 843 5168
rect 923 5162 975 5168
rect 1055 5162 1107 5168
rect 1187 5162 1239 5168
rect 1319 5162 1371 5168
rect 1451 5162 1503 5168
rect 1583 5162 1635 5168
rect 1715 5162 1767 5168
rect 1847 5162 1899 5168
rect 1979 5162 2031 5168
rect 2111 5162 2163 5168
rect 2243 5162 2295 5168
rect 2375 5162 2427 5168
rect 2507 5162 2559 5168
rect 2639 5162 2691 5168
rect 2771 5162 2823 5168
rect 2903 5162 2955 5168
rect 3035 5162 3087 5202
rect 688 4062 740 4114
rect 688 3995 740 4047
rect 688 3928 740 3980
rect 688 3861 740 3913
rect 688 3794 740 3846
rect 688 3727 740 3779
rect 688 3660 740 3712
rect 688 3593 740 3645
rect 688 3526 740 3578
rect 844 4802 896 4854
rect 844 4735 896 4787
rect 844 4668 896 4720
rect 844 4601 896 4653
rect 844 4534 896 4586
rect 844 4467 896 4519
rect 844 4400 896 4452
rect 844 4333 896 4385
rect 844 4266 896 4318
rect 1000 4062 1052 4114
rect 1000 3995 1052 4047
rect 1000 3928 1052 3980
rect 1000 3861 1052 3913
rect 1000 3794 1052 3846
rect 1000 3727 1052 3779
rect 1000 3660 1052 3712
rect 1000 3593 1052 3645
rect 1000 3526 1052 3578
rect 1156 4802 1208 4854
rect 1156 4735 1208 4787
rect 1156 4668 1208 4720
rect 1156 4601 1208 4653
rect 1156 4534 1208 4586
rect 1156 4467 1208 4519
rect 1156 4400 1208 4452
rect 1156 4333 1208 4385
rect 1156 4266 1208 4318
rect 1312 4062 1364 4114
rect 1312 3995 1364 4047
rect 1312 3928 1364 3980
rect 1312 3861 1364 3913
rect 1312 3794 1364 3846
rect 1312 3727 1364 3779
rect 1312 3660 1364 3712
rect 1312 3593 1364 3645
rect 1312 3526 1364 3578
rect 1468 4802 1520 4854
rect 1468 4735 1520 4787
rect 1468 4668 1520 4720
rect 1468 4601 1520 4653
rect 1468 4534 1520 4586
rect 1468 4467 1520 4519
rect 1468 4400 1520 4452
rect 1468 4333 1520 4385
rect 1468 4266 1520 4318
rect 1624 4062 1676 4114
rect 1624 3995 1676 4047
rect 1624 3928 1676 3980
rect 1624 3861 1676 3913
rect 1624 3794 1676 3846
rect 1624 3727 1676 3779
rect 1624 3660 1676 3712
rect 1624 3593 1676 3645
rect 1624 3526 1676 3578
rect 1780 4802 1832 4854
rect 1780 4735 1832 4787
rect 1780 4668 1832 4720
rect 1780 4601 1832 4653
rect 1780 4534 1832 4586
rect 1780 4467 1832 4519
rect 1780 4400 1832 4452
rect 1780 4333 1832 4385
rect 1780 4266 1832 4318
rect 1936 4062 1988 4114
rect 1936 3995 1988 4047
rect 1936 3928 1988 3980
rect 1936 3861 1988 3913
rect 1936 3794 1988 3846
rect 1936 3727 1988 3779
rect 1936 3660 1988 3712
rect 1936 3593 1988 3645
rect 1936 3526 1988 3578
rect 2092 4802 2144 4854
rect 2092 4735 2144 4787
rect 2092 4668 2144 4720
rect 2092 4601 2144 4653
rect 2092 4534 2144 4586
rect 2092 4467 2144 4519
rect 2092 4400 2144 4452
rect 2092 4333 2144 4385
rect 2092 4266 2144 4318
rect 2248 4062 2300 4114
rect 2248 3995 2300 4047
rect 2248 3928 2300 3980
rect 2248 3861 2300 3913
rect 2248 3794 2300 3846
rect 2248 3727 2300 3779
rect 2248 3660 2300 3712
rect 2248 3593 2300 3645
rect 2248 3526 2300 3578
rect 2404 4802 2456 4854
rect 2404 4735 2456 4787
rect 2404 4668 2456 4720
rect 2404 4601 2456 4653
rect 2404 4534 2456 4586
rect 2404 4467 2456 4519
rect 2404 4400 2456 4452
rect 2404 4333 2456 4385
rect 2404 4266 2456 4318
rect 2560 4062 2612 4114
rect 2560 3995 2612 4047
rect 2560 3928 2612 3980
rect 2560 3861 2612 3913
rect 2560 3794 2612 3846
rect 2560 3727 2612 3779
rect 2560 3660 2612 3712
rect 2560 3593 2612 3645
rect 2560 3526 2612 3578
rect 2716 4802 2768 4854
rect 2716 4735 2768 4787
rect 2716 4668 2768 4720
rect 2716 4601 2768 4653
rect 2716 4534 2768 4586
rect 2716 4467 2768 4519
rect 2716 4400 2768 4452
rect 2716 4333 2768 4385
rect 2716 4266 2768 4318
rect 2872 4062 2924 4114
rect 2872 3995 2924 4047
rect 2872 3928 2924 3980
rect 2872 3861 2924 3913
rect 2872 3794 2924 3846
rect 2872 3727 2924 3779
rect 2872 3660 2924 3712
rect 2872 3593 2924 3645
rect 2872 3526 2924 3578
rect 3210 4936 3253 4943
rect 3253 4936 3262 4943
rect 3274 4936 3287 4943
rect 3287 4936 3326 4943
rect 3210 4898 3262 4936
rect 3274 4898 3326 4936
rect 3210 4891 3253 4898
rect 3253 4891 3262 4898
rect 3274 4891 3287 4898
rect 3287 4891 3326 4898
rect 3210 4216 3253 4228
rect 3253 4216 3262 4228
rect 3274 4216 3287 4228
rect 3287 4216 3326 4228
rect 3210 4178 3262 4216
rect 3274 4178 3326 4216
rect 3210 4176 3253 4178
rect 3253 4176 3262 4178
rect 3274 4176 3287 4178
rect 3287 4176 3326 4178
rect 1335 3041 1387 3049
rect 1471 3041 1523 3049
rect 1607 3041 1659 3049
rect 1743 3041 1795 3049
rect 1879 3041 1931 3049
rect 2015 3041 2067 3049
rect 2151 3041 2203 3049
rect 2287 3041 2339 3049
rect 2423 3041 2475 3049
rect 2560 3041 2612 3049
rect 2697 3041 2749 3049
rect 1335 3007 1355 3041
rect 1355 3007 1387 3041
rect 1471 3007 1499 3041
rect 1499 3007 1523 3041
rect 1607 3007 1643 3041
rect 1643 3007 1659 3041
rect 1743 3007 1749 3041
rect 1749 3007 1787 3041
rect 1787 3007 1795 3041
rect 1879 3007 1893 3041
rect 1893 3007 1931 3041
rect 2015 3007 2037 3041
rect 2037 3007 2067 3041
rect 2151 3007 2181 3041
rect 2181 3007 2203 3041
rect 2287 3007 2291 3041
rect 2291 3007 2325 3041
rect 2325 3007 2339 3041
rect 2423 3007 2435 3041
rect 2435 3007 2469 3041
rect 2469 3007 2475 3041
rect 2560 3007 2579 3041
rect 2579 3007 2612 3041
rect 2697 3007 2723 3041
rect 2723 3007 2749 3041
rect 1335 2997 1387 3007
rect 1471 2997 1523 3007
rect 1607 2997 1659 3007
rect 1743 2997 1795 3007
rect 1879 2997 1931 3007
rect 2015 2997 2067 3007
rect 2151 2997 2203 3007
rect 2287 2997 2339 3007
rect 2423 2997 2475 3007
rect 2560 2997 2612 3007
rect 2697 2997 2749 3007
rect 1335 2921 1387 2930
rect 1471 2921 1523 2930
rect 1607 2921 1659 2930
rect 1743 2921 1795 2930
rect 1879 2921 1931 2930
rect 2015 2921 2067 2930
rect 2151 2921 2203 2930
rect 2287 2921 2339 2930
rect 2423 2921 2475 2930
rect 2560 2921 2612 2930
rect 2697 2921 2749 2930
rect 1335 2887 1355 2921
rect 1355 2887 1387 2921
rect 1471 2887 1499 2921
rect 1499 2887 1523 2921
rect 1607 2887 1643 2921
rect 1643 2887 1659 2921
rect 1743 2887 1749 2921
rect 1749 2887 1787 2921
rect 1787 2887 1795 2921
rect 1879 2887 1893 2921
rect 1893 2887 1931 2921
rect 2015 2887 2037 2921
rect 2037 2887 2067 2921
rect 2151 2887 2181 2921
rect 2181 2887 2203 2921
rect 2287 2887 2291 2921
rect 2291 2887 2325 2921
rect 2325 2887 2339 2921
rect 2423 2887 2435 2921
rect 2435 2887 2469 2921
rect 2469 2887 2475 2921
rect 2560 2887 2579 2921
rect 2579 2887 2612 2921
rect 2697 2887 2723 2921
rect 2723 2887 2749 2921
rect 1335 2878 1387 2887
rect 1471 2878 1523 2887
rect 1607 2878 1659 2887
rect 1743 2878 1795 2887
rect 1879 2878 1931 2887
rect 2015 2878 2067 2887
rect 2151 2878 2203 2887
rect 2287 2878 2339 2887
rect 2423 2878 2475 2887
rect 2560 2878 2612 2887
rect 2697 2878 2749 2887
rect 688 2512 740 2564
rect 688 2441 740 2493
rect 688 2370 740 2422
rect 688 2299 740 2351
rect 688 2228 740 2280
rect 688 2157 740 2209
rect 688 2086 740 2138
rect 688 2016 740 2068
rect 844 1813 896 1865
rect 844 1746 896 1798
rect 844 1679 896 1731
rect 844 1612 896 1664
rect 844 1545 896 1597
rect 844 1478 896 1530
rect 844 1411 896 1463
rect 844 1344 896 1396
rect 844 1277 896 1329
rect 1000 2552 1052 2604
rect 1000 2485 1052 2537
rect 1000 2418 1052 2470
rect 1000 2351 1052 2403
rect 1000 2284 1052 2336
rect 1000 2217 1052 2269
rect 1000 2150 1052 2202
rect 1000 2083 1052 2135
rect 1000 2016 1052 2068
rect 1156 1813 1208 1865
rect 1156 1746 1208 1798
rect 1156 1679 1208 1731
rect 1156 1612 1208 1664
rect 1156 1545 1208 1597
rect 1156 1478 1208 1530
rect 1156 1411 1208 1463
rect 1156 1344 1208 1396
rect 1156 1277 1208 1329
rect 1312 2552 1364 2604
rect 1312 2485 1364 2537
rect 1312 2418 1364 2470
rect 1312 2351 1364 2403
rect 1312 2284 1364 2336
rect 1312 2217 1364 2269
rect 1312 2150 1364 2202
rect 1312 2083 1364 2135
rect 1312 2016 1364 2068
rect 1468 1813 1520 1865
rect 1468 1746 1520 1798
rect 1468 1679 1520 1731
rect 1468 1612 1520 1664
rect 1468 1545 1520 1597
rect 1468 1478 1520 1530
rect 1468 1411 1520 1463
rect 1468 1344 1520 1396
rect 1468 1277 1520 1329
rect 1624 2552 1676 2604
rect 1624 2485 1676 2537
rect 1624 2418 1676 2470
rect 1624 2351 1676 2403
rect 1624 2284 1676 2336
rect 1624 2217 1676 2269
rect 1624 2150 1676 2202
rect 1624 2083 1676 2135
rect 1624 2016 1676 2068
rect 1780 1813 1832 1865
rect 1780 1746 1832 1798
rect 1780 1679 1832 1731
rect 1780 1612 1832 1664
rect 1780 1545 1832 1597
rect 1780 1478 1832 1530
rect 1780 1411 1832 1463
rect 1780 1344 1832 1396
rect 1780 1277 1832 1329
rect 1936 2552 1988 2604
rect 1936 2485 1988 2537
rect 1936 2418 1988 2470
rect 1936 2351 1988 2403
rect 1936 2284 1988 2336
rect 1936 2217 1988 2269
rect 1936 2150 1988 2202
rect 1936 2083 1988 2135
rect 1936 2016 1988 2068
rect 2092 1813 2144 1865
rect 2092 1746 2144 1798
rect 2092 1679 2144 1731
rect 2092 1612 2144 1664
rect 2092 1545 2144 1597
rect 2092 1478 2144 1530
rect 2092 1411 2144 1463
rect 2092 1344 2144 1396
rect 2092 1277 2144 1329
rect 2248 2552 2300 2604
rect 2248 2485 2300 2537
rect 2248 2418 2300 2470
rect 2248 2351 2300 2403
rect 2248 2284 2300 2336
rect 2248 2217 2300 2269
rect 2248 2150 2300 2202
rect 2248 2083 2300 2135
rect 2248 2016 2300 2068
rect 2404 1813 2456 1865
rect 2404 1746 2456 1798
rect 2404 1679 2456 1731
rect 2404 1612 2456 1664
rect 2404 1545 2456 1597
rect 2404 1478 2456 1530
rect 2404 1411 2456 1463
rect 2404 1344 2456 1396
rect 2404 1277 2456 1329
rect 2560 2552 2612 2604
rect 2560 2485 2612 2537
rect 2560 2418 2612 2470
rect 2560 2351 2612 2403
rect 2560 2284 2612 2336
rect 2560 2217 2612 2269
rect 2560 2150 2612 2202
rect 2560 2083 2612 2135
rect 2560 2016 2612 2068
rect 2716 1813 2768 1865
rect 2716 1746 2768 1798
rect 2716 1679 2768 1731
rect 2716 1612 2768 1664
rect 2716 1545 2768 1597
rect 2716 1478 2768 1530
rect 2716 1411 2768 1463
rect 2716 1344 2768 1396
rect 2716 1277 2768 1329
rect 2872 2552 2924 2604
rect 2872 2485 2924 2537
rect 2872 2418 2924 2470
rect 2872 2351 2924 2403
rect 2872 2284 2924 2336
rect 2872 2217 2924 2269
rect 2872 2150 2924 2202
rect 2872 2083 2924 2135
rect 2872 2016 2924 2068
rect 3985 2703 4037 2755
rect 4165 2703 4217 2755
rect 3210 1946 3262 1954
rect 3274 1946 3326 1954
rect 3210 1912 3253 1946
rect 3253 1912 3262 1946
rect 3274 1912 3287 1946
rect 3287 1912 3326 1946
rect 3210 1902 3262 1912
rect 3274 1902 3326 1912
rect 3210 1217 3262 1239
rect 3274 1217 3326 1239
rect 3210 1187 3253 1217
rect 3253 1187 3262 1217
rect 3274 1187 3287 1217
rect 3287 1187 3326 1217
rect 326 445 378 497
rect 391 488 443 497
rect 391 454 398 488
rect 398 454 432 488
rect 432 454 443 488
rect 391 445 443 454
rect 456 488 508 497
rect 456 454 472 488
rect 472 454 506 488
rect 506 454 508 488
rect 456 445 508 454
rect 521 488 573 497
rect 586 488 638 497
rect 651 488 703 497
rect 716 488 768 497
rect 781 488 833 497
rect 846 488 898 497
rect 521 454 546 488
rect 546 454 573 488
rect 586 454 620 488
rect 620 454 638 488
rect 651 454 654 488
rect 654 454 694 488
rect 694 454 703 488
rect 716 454 728 488
rect 728 454 768 488
rect 781 454 802 488
rect 802 454 833 488
rect 846 454 876 488
rect 876 454 898 488
rect 521 445 573 454
rect 586 445 638 454
rect 651 445 703 454
rect 716 445 768 454
rect 781 445 833 454
rect 846 445 898 454
rect 911 488 963 497
rect 911 454 916 488
rect 916 454 950 488
rect 950 454 963 488
rect 911 445 963 454
rect 976 488 1028 497
rect 976 454 990 488
rect 990 454 1024 488
rect 1024 454 1028 488
rect 976 445 1028 454
rect 1041 488 1093 497
rect 1106 488 1158 497
rect 1171 488 1223 497
rect 1236 488 1288 497
rect 1301 488 1353 497
rect 1366 488 1418 497
rect 1431 488 1483 497
rect 1041 454 1063 488
rect 1063 454 1093 488
rect 1106 454 1136 488
rect 1136 454 1158 488
rect 1171 454 1209 488
rect 1209 454 1223 488
rect 1236 454 1243 488
rect 1243 454 1282 488
rect 1282 454 1288 488
rect 1301 454 1316 488
rect 1316 454 1353 488
rect 1366 454 1389 488
rect 1389 454 1418 488
rect 1431 454 1462 488
rect 1462 454 1483 488
rect 1041 445 1093 454
rect 1106 445 1158 454
rect 1171 445 1223 454
rect 1236 445 1288 454
rect 1301 445 1353 454
rect 1366 445 1418 454
rect 1431 445 1483 454
rect 1496 488 1548 497
rect 1496 454 1501 488
rect 1501 454 1535 488
rect 1535 454 1548 488
rect 1496 445 1548 454
rect 1561 488 1613 497
rect 1561 454 1574 488
rect 1574 454 1608 488
rect 1608 454 1613 488
rect 1561 445 1613 454
rect 1626 488 1678 497
rect 1691 488 1743 497
rect 1756 488 1808 497
rect 1821 488 1873 497
rect 1886 488 1938 497
rect 1951 488 2003 497
rect 2016 488 2068 497
rect 1626 454 1647 488
rect 1647 454 1678 488
rect 1691 454 1720 488
rect 1720 454 1743 488
rect 1756 454 1793 488
rect 1793 454 1808 488
rect 1821 454 1827 488
rect 1827 454 1866 488
rect 1866 454 1873 488
rect 1886 454 1900 488
rect 1900 454 1938 488
rect 1951 454 1973 488
rect 1973 454 2003 488
rect 2016 454 2046 488
rect 2046 454 2068 488
rect 1626 445 1678 454
rect 1691 445 1743 454
rect 1756 445 1808 454
rect 1821 445 1873 454
rect 1886 445 1938 454
rect 1951 445 2003 454
rect 2016 445 2068 454
rect 2081 488 2133 497
rect 2081 454 2085 488
rect 2085 454 2119 488
rect 2119 454 2133 488
rect 2081 445 2133 454
rect 2146 488 2198 497
rect 2146 454 2158 488
rect 2158 454 2192 488
rect 2192 454 2198 488
rect 2146 445 2198 454
rect 2211 488 2263 497
rect 2275 488 2327 497
rect 2339 488 2391 497
rect 2403 488 2455 497
rect 2467 488 2519 497
rect 2531 488 2583 497
rect 2211 454 2231 488
rect 2231 454 2263 488
rect 2275 454 2304 488
rect 2304 454 2327 488
rect 2339 454 2377 488
rect 2377 454 2391 488
rect 2403 454 2411 488
rect 2411 454 2450 488
rect 2450 454 2455 488
rect 2467 454 2484 488
rect 2484 454 2519 488
rect 2531 454 2557 488
rect 2557 454 2583 488
rect 2211 445 2263 454
rect 2275 445 2327 454
rect 2339 445 2391 454
rect 2403 445 2455 454
rect 2467 445 2519 454
rect 2531 445 2583 454
rect 2595 488 2647 497
rect 2595 454 2596 488
rect 2596 454 2630 488
rect 2630 454 2647 488
rect 2595 445 2647 454
rect 2659 488 2711 497
rect 2659 454 2669 488
rect 2669 454 2703 488
rect 2703 454 2711 488
rect 2659 445 2711 454
rect 2723 488 2775 497
rect 2787 488 2839 497
rect 2851 488 2903 497
rect 2915 488 2967 497
rect 2979 488 3031 497
rect 3043 488 3095 497
rect 2723 454 2742 488
rect 2742 454 2775 488
rect 2787 454 2815 488
rect 2815 454 2839 488
rect 2851 454 2888 488
rect 2888 454 2903 488
rect 2915 454 2922 488
rect 2922 454 2961 488
rect 2961 454 2967 488
rect 2979 454 2995 488
rect 2995 454 3031 488
rect 3043 454 3068 488
rect 3068 454 3095 488
rect 2723 445 2775 454
rect 2787 445 2839 454
rect 2851 445 2903 454
rect 2915 445 2967 454
rect 2979 445 3031 454
rect 3043 445 3095 454
rect 3107 488 3159 497
rect 3107 454 3141 488
rect 3141 454 3159 488
rect 3107 445 3159 454
rect 3171 488 3223 497
rect 3171 454 3180 488
rect 3180 454 3214 488
rect 3214 454 3223 488
rect 3171 445 3223 454
rect 3235 445 3287 497
rect 4079 2422 4131 2474
rect 4079 2349 4131 2401
rect 4079 2276 4131 2328
rect 4079 2203 4131 2255
rect 4079 2130 4131 2182
rect 4079 2056 4131 2108
rect 3728 438 3780 490
rect 3828 438 3880 490
rect 3928 468 3980 490
rect 4029 468 4081 490
rect 4130 468 4182 490
rect 4231 468 4283 490
rect 3928 438 3945 468
rect 3945 438 3980 468
rect 4029 438 4059 468
rect 4059 438 4081 468
rect 4130 438 4133 468
rect 4133 438 4167 468
rect 4167 438 4182 468
rect 4231 438 4241 468
rect 4241 438 4281 468
rect 4281 438 4283 468
rect 4332 438 4384 490
rect 4433 438 4485 490
rect 4925 4062 4931 4114
rect 4931 4062 4977 4114
rect 4991 4062 5037 4114
rect 5037 4062 5043 4114
rect 4925 3973 4931 4025
rect 4931 3973 4977 4025
rect 4991 3973 5037 4025
rect 5037 3973 5043 4025
rect 4925 3884 4931 3936
rect 4931 3884 4977 3936
rect 4991 3884 5037 3936
rect 5037 3884 5043 3936
rect 4925 3795 4931 3847
rect 4931 3795 4977 3847
rect 4991 3795 5037 3847
rect 5037 3795 5043 3847
rect 4925 3706 4931 3758
rect 4931 3706 4977 3758
rect 4991 3706 5037 3758
rect 5037 3706 5043 3758
rect 4925 3616 4931 3668
rect 4931 3616 4977 3668
rect 4991 3616 5037 3668
rect 5037 3616 5043 3668
rect 4925 3543 4931 3578
rect 4931 3543 4977 3578
rect 4991 3543 5037 3578
rect 5037 3543 5043 3578
rect 4925 3526 4977 3543
rect 4991 3526 5043 3543
rect 5114 4062 5166 4114
rect 5114 3995 5166 4047
rect 5114 3928 5166 3980
rect 5114 3861 5166 3913
rect 5114 3794 5166 3846
rect 5114 3727 5166 3779
rect 5114 3660 5166 3712
rect 5114 3593 5166 3645
rect 5114 3526 5166 3578
rect 5270 4802 5322 4854
rect 5270 4735 5322 4787
rect 5270 4668 5322 4720
rect 5270 4601 5322 4653
rect 5270 4534 5322 4586
rect 5270 4467 5322 4519
rect 5270 4400 5322 4452
rect 5270 4333 5322 4385
rect 5270 4266 5322 4318
rect 5426 4062 5478 4114
rect 5426 3995 5478 4047
rect 5426 3928 5478 3980
rect 5426 3861 5478 3913
rect 5426 3794 5478 3846
rect 5426 3727 5478 3779
rect 5426 3660 5478 3712
rect 5426 3593 5478 3645
rect 5426 3526 5478 3578
rect 5582 4802 5634 4854
rect 5582 4735 5634 4787
rect 5582 4668 5634 4720
rect 5582 4601 5634 4653
rect 5582 4534 5634 4586
rect 5582 4467 5634 4519
rect 5582 4400 5634 4452
rect 5582 4333 5634 4385
rect 5582 4266 5634 4318
rect 5738 4062 5790 4114
rect 5738 3995 5790 4047
rect 5738 3928 5790 3980
rect 5738 3861 5790 3913
rect 5738 3794 5790 3846
rect 5738 3727 5790 3779
rect 5738 3660 5790 3712
rect 5738 3593 5790 3645
rect 5738 3526 5790 3578
rect 5894 4802 5946 4854
rect 5894 4735 5946 4787
rect 5894 4668 5946 4720
rect 5894 4601 5946 4653
rect 5894 4534 5946 4586
rect 5894 4467 5946 4519
rect 5894 4400 5946 4452
rect 5894 4333 5946 4385
rect 5894 4266 5946 4318
rect 6050 4062 6102 4114
rect 6050 3995 6102 4047
rect 6050 3928 6102 3980
rect 6050 3861 6102 3913
rect 6050 3794 6102 3846
rect 6050 3727 6102 3779
rect 6050 3660 6102 3712
rect 6050 3593 6102 3645
rect 6050 3526 6102 3578
rect 6205 4802 6257 4854
rect 6205 4735 6257 4787
rect 6205 4668 6257 4720
rect 6205 4601 6257 4653
rect 6205 4534 6257 4586
rect 6205 4467 6257 4519
rect 6205 4400 6257 4452
rect 6205 4333 6257 4385
rect 6205 4266 6257 4318
rect 6361 4062 6413 4114
rect 6361 3995 6413 4047
rect 6361 3928 6413 3980
rect 6361 3861 6413 3913
rect 6361 3794 6413 3846
rect 6361 3727 6413 3779
rect 6361 3660 6413 3712
rect 6361 3593 6413 3645
rect 6361 3526 6413 3578
rect 6517 4802 6569 4854
rect 6517 4735 6569 4787
rect 6517 4668 6569 4720
rect 6517 4601 6569 4653
rect 6517 4534 6569 4586
rect 6517 4467 6569 4519
rect 6517 4400 6569 4452
rect 6517 4333 6569 4385
rect 6517 4266 6569 4318
rect 6673 4062 6725 4114
rect 6673 3995 6725 4047
rect 6673 3928 6725 3980
rect 6673 3861 6725 3913
rect 6673 3794 6725 3846
rect 6673 3727 6725 3779
rect 6673 3660 6725 3712
rect 6673 3593 6725 3645
rect 6673 3526 6725 3578
rect 6830 4802 6882 4854
rect 6830 4735 6882 4787
rect 6830 4668 6882 4720
rect 6830 4601 6882 4653
rect 6830 4534 6882 4586
rect 6830 4467 6882 4519
rect 6830 4400 6882 4452
rect 6830 4333 6882 4385
rect 6830 4266 6882 4318
rect 6986 4062 7038 4114
rect 6986 3995 7038 4047
rect 6986 3928 7038 3980
rect 6986 3861 7038 3913
rect 6986 3794 7038 3846
rect 6986 3727 7038 3779
rect 6986 3660 7038 3712
rect 6986 3593 7038 3645
rect 6986 3526 7038 3578
rect 7142 4802 7194 4854
rect 7142 4735 7194 4787
rect 7142 4668 7194 4720
rect 7142 4601 7194 4653
rect 7142 4534 7194 4586
rect 7142 4467 7194 4519
rect 7142 4400 7194 4452
rect 7142 4333 7194 4385
rect 7142 4266 7194 4318
rect 7298 4062 7350 4114
rect 7298 3995 7350 4047
rect 7298 3928 7350 3980
rect 7298 3861 7350 3913
rect 7298 3794 7350 3846
rect 7298 3727 7350 3779
rect 7298 3660 7350 3712
rect 7298 3593 7350 3645
rect 7298 3526 7350 3578
rect 7454 4802 7506 4854
rect 7454 4735 7506 4787
rect 7454 4668 7506 4720
rect 7454 4601 7506 4653
rect 7454 4534 7506 4586
rect 7454 4467 7506 4519
rect 7454 4400 7506 4452
rect 7454 4333 7506 4385
rect 7454 4266 7506 4318
rect 7610 4062 7662 4114
rect 7610 3995 7662 4047
rect 7610 3928 7662 3980
rect 7610 3861 7662 3913
rect 7610 3794 7662 3846
rect 7610 3727 7662 3779
rect 7610 3660 7662 3712
rect 7610 3593 7662 3645
rect 7610 3526 7662 3578
rect 7766 4802 7818 4854
rect 7766 4735 7818 4787
rect 7766 4668 7818 4720
rect 7766 4601 7818 4653
rect 7766 4534 7818 4586
rect 7766 4467 7818 4519
rect 7766 4400 7818 4452
rect 7766 4333 7818 4385
rect 7766 4266 7818 4318
rect 7922 4062 7974 4114
rect 7922 3995 7974 4047
rect 7922 3928 7974 3980
rect 7922 3861 7974 3913
rect 7922 3794 7974 3846
rect 7922 3727 7974 3779
rect 7922 3660 7974 3712
rect 7922 3593 7974 3645
rect 7922 3526 7974 3578
rect 8078 4802 8130 4854
rect 8078 4735 8130 4787
rect 8078 4668 8130 4720
rect 8078 4601 8130 4653
rect 8078 4534 8130 4586
rect 8078 4467 8130 4519
rect 8078 4400 8130 4452
rect 8078 4333 8130 4385
rect 8078 4266 8130 4318
rect 8234 4062 8286 4114
rect 8234 3995 8286 4047
rect 8234 3928 8286 3980
rect 8234 3861 8286 3913
rect 8234 3794 8286 3846
rect 8234 3727 8286 3779
rect 8234 3660 8286 3712
rect 8234 3593 8286 3645
rect 8234 3526 8286 3578
rect 8390 4802 8442 4854
rect 8390 4735 8442 4787
rect 8390 4668 8442 4720
rect 8390 4601 8442 4653
rect 8390 4534 8442 4586
rect 8390 4467 8442 4519
rect 8390 4400 8442 4452
rect 8390 4333 8442 4385
rect 8390 4266 8442 4318
rect 8546 4062 8598 4114
rect 8546 3995 8598 4047
rect 8546 3928 8598 3980
rect 8546 3861 8598 3913
rect 8546 3794 8598 3846
rect 8546 3727 8598 3779
rect 8546 3660 8598 3712
rect 8546 3593 8598 3645
rect 8546 3526 8598 3578
rect 8702 4802 8754 4854
rect 8702 4735 8754 4787
rect 8702 4668 8754 4720
rect 8702 4601 8754 4653
rect 8702 4534 8754 4586
rect 8702 4467 8754 4519
rect 8702 4400 8754 4452
rect 8702 4333 8754 4385
rect 8702 4266 8754 4318
rect 8858 4062 8910 4114
rect 8858 3995 8910 4047
rect 8858 3928 8910 3980
rect 8858 3861 8910 3913
rect 8858 3794 8910 3846
rect 8858 3727 8910 3779
rect 8858 3660 8910 3712
rect 8858 3593 8910 3645
rect 8858 3526 8910 3578
rect 9014 4802 9066 4854
rect 9014 4735 9066 4787
rect 9014 4668 9066 4720
rect 9014 4601 9066 4653
rect 9014 4534 9066 4586
rect 9014 4467 9066 4519
rect 9014 4400 9066 4452
rect 9014 4333 9066 4385
rect 9014 4266 9066 4318
rect 9170 4062 9222 4114
rect 9170 3995 9222 4047
rect 9170 3928 9222 3980
rect 9170 3861 9222 3913
rect 9170 3794 9222 3846
rect 9170 3727 9222 3779
rect 9170 3660 9222 3712
rect 9170 3593 9222 3645
rect 9170 3526 9222 3578
rect 9326 4802 9378 4854
rect 9326 4735 9378 4787
rect 9326 4668 9378 4720
rect 9326 4601 9378 4653
rect 9326 4534 9378 4586
rect 9326 4467 9378 4519
rect 9326 4400 9378 4452
rect 9326 4333 9378 4385
rect 9326 4266 9378 4318
rect 9482 4062 9534 4114
rect 9482 3995 9534 4047
rect 9482 3928 9534 3980
rect 9482 3861 9534 3913
rect 9482 3794 9534 3846
rect 9482 3727 9534 3779
rect 9482 3660 9534 3712
rect 9482 3593 9534 3645
rect 9482 3526 9534 3578
rect 9638 4802 9690 4854
rect 9638 4735 9690 4787
rect 9638 4668 9690 4720
rect 9638 4601 9690 4653
rect 9638 4534 9690 4586
rect 9638 4467 9690 4519
rect 9638 4400 9690 4452
rect 9638 4333 9690 4385
rect 9638 4266 9690 4318
rect 9794 4062 9846 4114
rect 9794 3995 9846 4047
rect 9794 3928 9846 3980
rect 9794 3861 9846 3913
rect 9794 3794 9846 3846
rect 9794 3727 9846 3779
rect 9794 3660 9846 3712
rect 9794 3593 9846 3645
rect 9794 3526 9846 3578
rect 9917 4102 9923 4114
rect 9923 4102 9957 4114
rect 9957 4102 9969 4114
rect 9917 4063 9969 4102
rect 9917 4062 9923 4063
rect 9923 4062 9957 4063
rect 9957 4062 9969 4063
rect 9983 4102 9995 4114
rect 9995 4102 10029 4114
rect 10029 4102 10035 4114
rect 9983 4063 10035 4102
rect 9983 4062 9995 4063
rect 9995 4062 10029 4063
rect 10029 4062 10035 4063
rect 9917 3990 9969 4025
rect 9917 3973 9923 3990
rect 9923 3973 9957 3990
rect 9957 3973 9969 3990
rect 9983 3990 10035 4025
rect 9983 3973 9995 3990
rect 9995 3973 10029 3990
rect 10029 3973 10035 3990
rect 9917 3917 9969 3936
rect 9917 3884 9923 3917
rect 9923 3884 9957 3917
rect 9957 3884 9969 3917
rect 9983 3917 10035 3936
rect 9983 3884 9995 3917
rect 9995 3884 10029 3917
rect 10029 3884 10035 3917
rect 9917 3844 9969 3847
rect 9917 3810 9923 3844
rect 9923 3810 9957 3844
rect 9957 3810 9969 3844
rect 9917 3795 9969 3810
rect 9983 3844 10035 3847
rect 9983 3810 9995 3844
rect 9995 3810 10029 3844
rect 10029 3810 10035 3844
rect 9983 3795 10035 3810
rect 9917 3737 9923 3758
rect 9923 3737 9957 3758
rect 9957 3737 9969 3758
rect 9917 3706 9969 3737
rect 9983 3737 9995 3758
rect 9995 3737 10029 3758
rect 10029 3737 10035 3758
rect 9983 3706 10035 3737
rect 9917 3664 9923 3668
rect 9923 3664 9957 3668
rect 9957 3664 9969 3668
rect 9917 3625 9969 3664
rect 9917 3616 9923 3625
rect 9923 3616 9957 3625
rect 9957 3616 9969 3625
rect 9983 3664 9995 3668
rect 9995 3664 10029 3668
rect 10029 3664 10035 3668
rect 9983 3625 10035 3664
rect 9983 3616 9995 3625
rect 9995 3616 10029 3625
rect 10029 3616 10035 3625
rect 9917 3552 9969 3578
rect 9917 3526 9923 3552
rect 9923 3526 9957 3552
rect 9957 3526 9969 3552
rect 9983 3552 10035 3578
rect 9983 3526 9995 3552
rect 9995 3526 10029 3552
rect 10029 3526 10035 3552
rect 5303 3216 5355 3225
rect 5367 3216 5419 3225
rect 5431 3216 5483 3225
rect 5495 3216 5547 3225
rect 5303 3182 5309 3216
rect 5309 3182 5347 3216
rect 5347 3182 5355 3216
rect 5367 3182 5381 3216
rect 5381 3182 5419 3216
rect 5431 3182 5453 3216
rect 5453 3182 5483 3216
rect 5495 3182 5525 3216
rect 5525 3182 5547 3216
rect 5303 3173 5355 3182
rect 5367 3173 5419 3182
rect 5431 3173 5483 3182
rect 5495 3173 5547 3182
rect 5559 3216 5611 3225
rect 5559 3182 5563 3216
rect 5563 3182 5597 3216
rect 5597 3182 5611 3216
rect 5559 3173 5611 3182
rect 5623 3216 5675 3225
rect 5623 3182 5635 3216
rect 5635 3182 5669 3216
rect 5669 3182 5675 3216
rect 5623 3173 5675 3182
rect 5687 3216 5739 3225
rect 5751 3216 5803 3225
rect 5815 3216 5867 3225
rect 5879 3216 5931 3225
rect 5943 3216 5995 3225
rect 6007 3216 6059 3225
rect 6071 3216 6123 3225
rect 5687 3182 5707 3216
rect 5707 3182 5739 3216
rect 5751 3182 5779 3216
rect 5779 3182 5803 3216
rect 5815 3182 5851 3216
rect 5851 3182 5867 3216
rect 5879 3182 5885 3216
rect 5885 3182 5923 3216
rect 5923 3182 5931 3216
rect 5943 3182 5957 3216
rect 5957 3182 5995 3216
rect 6007 3182 6029 3216
rect 6029 3182 6059 3216
rect 6071 3182 6101 3216
rect 6101 3182 6123 3216
rect 5687 3173 5739 3182
rect 5751 3173 5803 3182
rect 5815 3173 5867 3182
rect 5879 3173 5931 3182
rect 5943 3173 5995 3182
rect 6007 3173 6059 3182
rect 6071 3173 6123 3182
rect 6135 3216 6187 3225
rect 6135 3182 6139 3216
rect 6139 3182 6173 3216
rect 6173 3182 6187 3216
rect 6135 3173 6187 3182
rect 6199 3216 6251 3225
rect 6199 3182 6211 3216
rect 6211 3182 6245 3216
rect 6245 3182 6251 3216
rect 6199 3173 6251 3182
rect 6263 3216 6315 3225
rect 6327 3216 6379 3225
rect 6391 3216 6443 3225
rect 6456 3216 6508 3225
rect 6521 3216 6573 3225
rect 6586 3216 6638 3225
rect 6651 3216 6703 3225
rect 6716 3216 6768 3225
rect 6263 3182 6283 3216
rect 6283 3182 6315 3216
rect 6327 3182 6355 3216
rect 6355 3182 6379 3216
rect 6391 3182 6427 3216
rect 6427 3182 6443 3216
rect 6456 3182 6461 3216
rect 6461 3182 6499 3216
rect 6499 3182 6508 3216
rect 6521 3182 6533 3216
rect 6533 3182 6571 3216
rect 6571 3182 6573 3216
rect 6586 3182 6605 3216
rect 6605 3182 6638 3216
rect 6651 3182 6677 3216
rect 6677 3182 6703 3216
rect 6716 3182 6749 3216
rect 6749 3182 6768 3216
rect 6263 3173 6315 3182
rect 6327 3173 6379 3182
rect 6391 3173 6443 3182
rect 6456 3173 6508 3182
rect 6521 3173 6573 3182
rect 6586 3173 6638 3182
rect 6651 3173 6703 3182
rect 6716 3173 6768 3182
rect 6781 3216 6833 3225
rect 6781 3182 6787 3216
rect 6787 3182 6821 3216
rect 6821 3182 6833 3216
rect 6781 3173 6833 3182
rect 6846 3216 6898 3225
rect 6846 3182 6859 3216
rect 6859 3182 6893 3216
rect 6893 3182 6898 3216
rect 6846 3173 6898 3182
rect 6911 3216 6963 3225
rect 6976 3216 7028 3225
rect 7041 3216 7093 3225
rect 7106 3216 7158 3225
rect 7171 3216 7223 3225
rect 7236 3216 7288 3225
rect 7301 3216 7353 3225
rect 7366 3216 7418 3225
rect 6911 3182 6931 3216
rect 6931 3182 6963 3216
rect 6976 3182 7003 3216
rect 7003 3182 7028 3216
rect 7041 3182 7075 3216
rect 7075 3182 7093 3216
rect 7106 3182 7109 3216
rect 7109 3182 7147 3216
rect 7147 3182 7158 3216
rect 7171 3182 7181 3216
rect 7181 3182 7219 3216
rect 7219 3182 7223 3216
rect 7236 3182 7253 3216
rect 7253 3182 7288 3216
rect 7301 3182 7325 3216
rect 7325 3182 7353 3216
rect 7366 3182 7397 3216
rect 7397 3182 7418 3216
rect 6911 3173 6963 3182
rect 6976 3173 7028 3182
rect 7041 3173 7093 3182
rect 7106 3173 7158 3182
rect 7171 3173 7223 3182
rect 7236 3173 7288 3182
rect 7301 3173 7353 3182
rect 7366 3173 7418 3182
rect 7431 3216 7483 3225
rect 7431 3182 7435 3216
rect 7435 3182 7469 3216
rect 7469 3182 7483 3216
rect 7431 3173 7483 3182
rect 7496 3216 7548 3225
rect 7496 3182 7507 3216
rect 7507 3182 7541 3216
rect 7541 3182 7548 3216
rect 7496 3173 7548 3182
rect 7561 3216 7613 3225
rect 7561 3182 7579 3216
rect 7579 3182 7613 3216
rect 7561 3173 7613 3182
rect 7626 3216 7678 3225
rect 7691 3216 7743 3225
rect 7756 3216 7808 3225
rect 7821 3216 7873 3225
rect 7886 3216 7938 3225
rect 7951 3216 8003 3225
rect 8016 3216 8068 3225
rect 7626 3182 7651 3216
rect 7651 3182 7678 3216
rect 7691 3182 7723 3216
rect 7723 3182 7743 3216
rect 7756 3182 7757 3216
rect 7757 3182 7795 3216
rect 7795 3182 7808 3216
rect 7821 3182 7829 3216
rect 7829 3182 7867 3216
rect 7867 3182 7873 3216
rect 7886 3182 7901 3216
rect 7901 3182 7938 3216
rect 7951 3182 7973 3216
rect 7973 3182 8003 3216
rect 8016 3182 8045 3216
rect 8045 3182 8068 3216
rect 7626 3173 7678 3182
rect 7691 3173 7743 3182
rect 7756 3173 7808 3182
rect 7821 3173 7873 3182
rect 7886 3173 7938 3182
rect 7951 3173 8003 3182
rect 8016 3173 8068 3182
rect 8081 3216 8133 3225
rect 8081 3182 8083 3216
rect 8083 3182 8117 3216
rect 8117 3182 8133 3216
rect 8081 3173 8133 3182
rect 8146 3216 8198 3225
rect 8146 3182 8155 3216
rect 8155 3182 8189 3216
rect 8189 3182 8198 3216
rect 8146 3173 8198 3182
rect 8211 3216 8263 3225
rect 8211 3182 8227 3216
rect 8227 3182 8261 3216
rect 8261 3182 8263 3216
rect 8211 3173 8263 3182
rect 8276 3216 8328 3225
rect 8341 3216 8393 3225
rect 8406 3216 8458 3225
rect 8471 3216 8523 3225
rect 8536 3216 8588 3225
rect 8601 3216 8653 3225
rect 8666 3216 8718 3225
rect 8276 3182 8299 3216
rect 8299 3182 8328 3216
rect 8341 3182 8371 3216
rect 8371 3182 8393 3216
rect 8406 3182 8443 3216
rect 8443 3182 8458 3216
rect 8471 3182 8477 3216
rect 8477 3182 8515 3216
rect 8515 3182 8523 3216
rect 8536 3182 8549 3216
rect 8549 3182 8587 3216
rect 8587 3182 8588 3216
rect 8601 3182 8621 3216
rect 8621 3182 8653 3216
rect 8666 3182 8693 3216
rect 8693 3182 8718 3216
rect 8276 3173 8328 3182
rect 8341 3173 8393 3182
rect 8406 3173 8458 3182
rect 8471 3173 8523 3182
rect 8536 3173 8588 3182
rect 8601 3173 8653 3182
rect 8666 3173 8718 3182
rect 8731 3216 8783 3225
rect 8731 3182 8765 3216
rect 8765 3182 8783 3216
rect 8731 3173 8783 3182
rect 8796 3216 8848 3225
rect 8796 3182 8803 3216
rect 8803 3182 8837 3216
rect 8837 3182 8848 3216
rect 8796 3173 8848 3182
rect 8861 3216 8913 3225
rect 8861 3182 8875 3216
rect 8875 3182 8909 3216
rect 8909 3182 8913 3216
rect 8861 3173 8913 3182
rect 8926 3216 8978 3225
rect 8991 3216 9043 3225
rect 9056 3216 9108 3225
rect 9121 3216 9173 3225
rect 9186 3216 9238 3225
rect 9251 3216 9303 3225
rect 9316 3216 9368 3225
rect 9381 3216 9433 3225
rect 8926 3182 8947 3216
rect 8947 3182 8978 3216
rect 8991 3182 9019 3216
rect 9019 3182 9043 3216
rect 9056 3182 9091 3216
rect 9091 3182 9108 3216
rect 9121 3182 9125 3216
rect 9125 3182 9163 3216
rect 9163 3182 9173 3216
rect 9186 3182 9197 3216
rect 9197 3182 9235 3216
rect 9235 3182 9238 3216
rect 9251 3182 9269 3216
rect 9269 3182 9303 3216
rect 9316 3182 9341 3216
rect 9341 3182 9368 3216
rect 9381 3182 9413 3216
rect 9413 3182 9433 3216
rect 8926 3173 8978 3182
rect 8991 3173 9043 3182
rect 9056 3173 9108 3182
rect 9121 3173 9173 3182
rect 9186 3173 9238 3182
rect 9251 3173 9303 3182
rect 9316 3173 9368 3182
rect 9381 3173 9433 3182
rect 9446 3216 9498 3225
rect 9446 3182 9451 3216
rect 9451 3182 9485 3216
rect 9485 3182 9498 3216
rect 9446 3173 9498 3182
rect 5303 2746 5355 2755
rect 5367 2746 5419 2755
rect 5431 2746 5483 2755
rect 5495 2746 5547 2755
rect 5303 2712 5309 2746
rect 5309 2712 5347 2746
rect 5347 2712 5355 2746
rect 5367 2712 5381 2746
rect 5381 2712 5419 2746
rect 5431 2712 5453 2746
rect 5453 2712 5483 2746
rect 5495 2712 5525 2746
rect 5525 2712 5547 2746
rect 5303 2703 5355 2712
rect 5367 2703 5419 2712
rect 5431 2703 5483 2712
rect 5495 2703 5547 2712
rect 5559 2746 5611 2755
rect 5559 2712 5563 2746
rect 5563 2712 5597 2746
rect 5597 2712 5611 2746
rect 5559 2703 5611 2712
rect 5623 2746 5675 2755
rect 5623 2712 5635 2746
rect 5635 2712 5669 2746
rect 5669 2712 5675 2746
rect 5623 2703 5675 2712
rect 5687 2746 5739 2755
rect 5751 2746 5803 2755
rect 5815 2746 5867 2755
rect 5879 2746 5931 2755
rect 5943 2746 5995 2755
rect 6007 2746 6059 2755
rect 6071 2746 6123 2755
rect 5687 2712 5707 2746
rect 5707 2712 5739 2746
rect 5751 2712 5779 2746
rect 5779 2712 5803 2746
rect 5815 2712 5851 2746
rect 5851 2712 5867 2746
rect 5879 2712 5885 2746
rect 5885 2712 5923 2746
rect 5923 2712 5931 2746
rect 5943 2712 5957 2746
rect 5957 2712 5995 2746
rect 6007 2712 6029 2746
rect 6029 2712 6059 2746
rect 6071 2712 6101 2746
rect 6101 2712 6123 2746
rect 5687 2703 5739 2712
rect 5751 2703 5803 2712
rect 5815 2703 5867 2712
rect 5879 2703 5931 2712
rect 5943 2703 5995 2712
rect 6007 2703 6059 2712
rect 6071 2703 6123 2712
rect 6135 2746 6187 2755
rect 6135 2712 6139 2746
rect 6139 2712 6173 2746
rect 6173 2712 6187 2746
rect 6135 2703 6187 2712
rect 6199 2746 6251 2755
rect 6199 2712 6211 2746
rect 6211 2712 6245 2746
rect 6245 2712 6251 2746
rect 6199 2703 6251 2712
rect 6263 2746 6315 2755
rect 6327 2746 6379 2755
rect 6391 2746 6443 2755
rect 6456 2746 6508 2755
rect 6521 2746 6573 2755
rect 6586 2746 6638 2755
rect 6651 2746 6703 2755
rect 6716 2746 6768 2755
rect 6263 2712 6283 2746
rect 6283 2712 6315 2746
rect 6327 2712 6355 2746
rect 6355 2712 6379 2746
rect 6391 2712 6427 2746
rect 6427 2712 6443 2746
rect 6456 2712 6461 2746
rect 6461 2712 6499 2746
rect 6499 2712 6508 2746
rect 6521 2712 6533 2746
rect 6533 2712 6571 2746
rect 6571 2712 6573 2746
rect 6586 2712 6605 2746
rect 6605 2712 6638 2746
rect 6651 2712 6677 2746
rect 6677 2712 6703 2746
rect 6716 2712 6749 2746
rect 6749 2712 6768 2746
rect 6263 2703 6315 2712
rect 6327 2703 6379 2712
rect 6391 2703 6443 2712
rect 6456 2703 6508 2712
rect 6521 2703 6573 2712
rect 6586 2703 6638 2712
rect 6651 2703 6703 2712
rect 6716 2703 6768 2712
rect 6781 2746 6833 2755
rect 6781 2712 6787 2746
rect 6787 2712 6821 2746
rect 6821 2712 6833 2746
rect 6781 2703 6833 2712
rect 6846 2746 6898 2755
rect 6846 2712 6859 2746
rect 6859 2712 6893 2746
rect 6893 2712 6898 2746
rect 6846 2703 6898 2712
rect 6911 2746 6963 2755
rect 6976 2746 7028 2755
rect 7041 2746 7093 2755
rect 7106 2746 7158 2755
rect 7171 2746 7223 2755
rect 7236 2746 7288 2755
rect 7301 2746 7353 2755
rect 7366 2746 7418 2755
rect 6911 2712 6931 2746
rect 6931 2712 6963 2746
rect 6976 2712 7003 2746
rect 7003 2712 7028 2746
rect 7041 2712 7075 2746
rect 7075 2712 7093 2746
rect 7106 2712 7109 2746
rect 7109 2712 7147 2746
rect 7147 2712 7158 2746
rect 7171 2712 7181 2746
rect 7181 2712 7219 2746
rect 7219 2712 7223 2746
rect 7236 2712 7253 2746
rect 7253 2712 7288 2746
rect 7301 2712 7325 2746
rect 7325 2712 7353 2746
rect 7366 2712 7397 2746
rect 7397 2712 7418 2746
rect 6911 2703 6963 2712
rect 6976 2703 7028 2712
rect 7041 2703 7093 2712
rect 7106 2703 7158 2712
rect 7171 2703 7223 2712
rect 7236 2703 7288 2712
rect 7301 2703 7353 2712
rect 7366 2703 7418 2712
rect 7431 2746 7483 2755
rect 7431 2712 7435 2746
rect 7435 2712 7469 2746
rect 7469 2712 7483 2746
rect 7431 2703 7483 2712
rect 7496 2746 7548 2755
rect 7496 2712 7507 2746
rect 7507 2712 7541 2746
rect 7541 2712 7548 2746
rect 7496 2703 7548 2712
rect 7561 2746 7613 2755
rect 7561 2712 7579 2746
rect 7579 2712 7613 2746
rect 7561 2703 7613 2712
rect 7626 2746 7678 2755
rect 7691 2746 7743 2755
rect 7756 2746 7808 2755
rect 7821 2746 7873 2755
rect 7886 2746 7938 2755
rect 7951 2746 8003 2755
rect 8016 2746 8068 2755
rect 7626 2712 7651 2746
rect 7651 2712 7678 2746
rect 7691 2712 7723 2746
rect 7723 2712 7743 2746
rect 7756 2712 7757 2746
rect 7757 2712 7795 2746
rect 7795 2712 7808 2746
rect 7821 2712 7829 2746
rect 7829 2712 7867 2746
rect 7867 2712 7873 2746
rect 7886 2712 7901 2746
rect 7901 2712 7938 2746
rect 7951 2712 7973 2746
rect 7973 2712 8003 2746
rect 8016 2712 8045 2746
rect 8045 2712 8068 2746
rect 7626 2703 7678 2712
rect 7691 2703 7743 2712
rect 7756 2703 7808 2712
rect 7821 2703 7873 2712
rect 7886 2703 7938 2712
rect 7951 2703 8003 2712
rect 8016 2703 8068 2712
rect 8081 2746 8133 2755
rect 8081 2712 8083 2746
rect 8083 2712 8117 2746
rect 8117 2712 8133 2746
rect 8081 2703 8133 2712
rect 8146 2746 8198 2755
rect 8146 2712 8155 2746
rect 8155 2712 8189 2746
rect 8189 2712 8198 2746
rect 8146 2703 8198 2712
rect 8211 2746 8263 2755
rect 8211 2712 8227 2746
rect 8227 2712 8261 2746
rect 8261 2712 8263 2746
rect 8211 2703 8263 2712
rect 8276 2746 8328 2755
rect 8341 2746 8393 2755
rect 8406 2746 8458 2755
rect 8471 2746 8523 2755
rect 8536 2746 8588 2755
rect 8601 2746 8653 2755
rect 8666 2746 8718 2755
rect 8276 2712 8299 2746
rect 8299 2712 8328 2746
rect 8341 2712 8371 2746
rect 8371 2712 8393 2746
rect 8406 2712 8443 2746
rect 8443 2712 8458 2746
rect 8471 2712 8477 2746
rect 8477 2712 8515 2746
rect 8515 2712 8523 2746
rect 8536 2712 8549 2746
rect 8549 2712 8587 2746
rect 8587 2712 8588 2746
rect 8601 2712 8621 2746
rect 8621 2712 8653 2746
rect 8666 2712 8693 2746
rect 8693 2712 8718 2746
rect 8276 2703 8328 2712
rect 8341 2703 8393 2712
rect 8406 2703 8458 2712
rect 8471 2703 8523 2712
rect 8536 2703 8588 2712
rect 8601 2703 8653 2712
rect 8666 2703 8718 2712
rect 8731 2746 8783 2755
rect 8731 2712 8765 2746
rect 8765 2712 8783 2746
rect 8731 2703 8783 2712
rect 8796 2746 8848 2755
rect 8796 2712 8803 2746
rect 8803 2712 8837 2746
rect 8837 2712 8848 2746
rect 8796 2703 8848 2712
rect 8861 2746 8913 2755
rect 8861 2712 8875 2746
rect 8875 2712 8909 2746
rect 8909 2712 8913 2746
rect 8861 2703 8913 2712
rect 8926 2746 8978 2755
rect 8991 2746 9043 2755
rect 9056 2746 9108 2755
rect 9121 2746 9173 2755
rect 9186 2746 9238 2755
rect 9251 2746 9303 2755
rect 9316 2746 9368 2755
rect 9381 2746 9433 2755
rect 8926 2712 8947 2746
rect 8947 2712 8978 2746
rect 8991 2712 9019 2746
rect 9019 2712 9043 2746
rect 9056 2712 9091 2746
rect 9091 2712 9108 2746
rect 9121 2712 9125 2746
rect 9125 2712 9163 2746
rect 9163 2712 9173 2746
rect 9186 2712 9197 2746
rect 9197 2712 9235 2746
rect 9235 2712 9238 2746
rect 9251 2712 9269 2746
rect 9269 2712 9303 2746
rect 9316 2712 9341 2746
rect 9341 2712 9368 2746
rect 9381 2712 9413 2746
rect 9413 2712 9433 2746
rect 8926 2703 8978 2712
rect 8991 2703 9043 2712
rect 9056 2703 9108 2712
rect 9121 2703 9173 2712
rect 9186 2703 9238 2712
rect 9251 2703 9303 2712
rect 9316 2703 9368 2712
rect 9381 2703 9433 2712
rect 9446 2746 9498 2755
rect 9446 2712 9451 2746
rect 9451 2712 9485 2746
rect 9485 2712 9498 2746
rect 9446 2703 9498 2712
rect 4925 2594 4931 2604
rect 4931 2594 4965 2604
rect 4965 2594 4977 2604
rect 4925 2555 4977 2594
rect 4925 2552 4931 2555
rect 4931 2552 4965 2555
rect 4965 2552 4977 2555
rect 4991 2594 5003 2604
rect 5003 2594 5037 2604
rect 5037 2594 5043 2604
rect 4991 2555 5043 2594
rect 4991 2552 5003 2555
rect 5003 2552 5037 2555
rect 5037 2552 5043 2555
rect 4925 2521 4931 2522
rect 4931 2521 4965 2522
rect 4965 2521 4977 2522
rect 4925 2482 4977 2521
rect 4925 2470 4931 2482
rect 4931 2470 4965 2482
rect 4965 2470 4977 2482
rect 4991 2521 5003 2522
rect 5003 2521 5037 2522
rect 5037 2521 5043 2522
rect 4991 2482 5043 2521
rect 4991 2470 5003 2482
rect 5003 2470 5037 2482
rect 5037 2470 5043 2482
rect 4925 2409 4977 2440
rect 4925 2388 4931 2409
rect 4931 2388 4965 2409
rect 4965 2388 4977 2409
rect 4991 2409 5043 2440
rect 4991 2388 5003 2409
rect 5003 2388 5037 2409
rect 5037 2388 5043 2409
rect 4925 2336 4977 2357
rect 4925 2305 4931 2336
rect 4931 2305 4965 2336
rect 4965 2305 4977 2336
rect 4991 2336 5043 2357
rect 4991 2305 5003 2336
rect 5003 2305 5037 2336
rect 5037 2305 5043 2336
rect 4925 2263 4977 2274
rect 4925 2229 4931 2263
rect 4931 2229 4965 2263
rect 4965 2229 4977 2263
rect 4925 2222 4977 2229
rect 4991 2263 5043 2274
rect 4991 2229 5003 2263
rect 5003 2229 5037 2263
rect 5037 2229 5043 2263
rect 4991 2222 5043 2229
rect 4925 2190 4977 2191
rect 4925 2156 4931 2190
rect 4931 2156 4965 2190
rect 4965 2156 4977 2190
rect 4925 2139 4977 2156
rect 4991 2190 5043 2191
rect 4991 2156 5003 2190
rect 5003 2156 5037 2190
rect 5037 2156 5043 2190
rect 4991 2139 5043 2156
rect 4925 2083 4931 2108
rect 4931 2083 4965 2108
rect 4965 2083 4977 2108
rect 4925 2056 4977 2083
rect 4991 2083 5003 2108
rect 5003 2083 5037 2108
rect 5037 2083 5043 2108
rect 4991 2056 5043 2083
rect 5114 2552 5166 2604
rect 5114 2485 5166 2537
rect 5114 2418 5166 2470
rect 5114 2351 5166 2403
rect 5114 2284 5166 2336
rect 5114 2217 5166 2269
rect 5114 2150 5166 2202
rect 5114 2083 5166 2135
rect 5114 2016 5166 2068
rect 5270 1813 5322 1865
rect 5270 1746 5322 1798
rect 5270 1679 5322 1731
rect 5270 1612 5322 1664
rect 5270 1545 5322 1597
rect 5270 1478 5322 1530
rect 5270 1411 5322 1463
rect 5270 1344 5322 1396
rect 5270 1277 5322 1329
rect 5426 2552 5478 2604
rect 5426 2485 5478 2537
rect 5426 2418 5478 2470
rect 5426 2351 5478 2403
rect 5426 2284 5478 2336
rect 5426 2217 5478 2269
rect 5426 2150 5478 2202
rect 5426 2083 5478 2135
rect 5426 2016 5478 2068
rect 5582 1813 5634 1865
rect 5582 1746 5634 1798
rect 5582 1679 5634 1731
rect 5582 1612 5634 1664
rect 5582 1545 5634 1597
rect 5582 1478 5634 1530
rect 5582 1411 5634 1463
rect 5582 1344 5634 1396
rect 5582 1277 5634 1329
rect 5738 2552 5790 2604
rect 5738 2485 5790 2537
rect 5738 2418 5790 2470
rect 5738 2351 5790 2403
rect 5738 2284 5790 2336
rect 5738 2217 5790 2269
rect 5738 2150 5790 2202
rect 5738 2083 5790 2135
rect 5738 2016 5790 2068
rect 5894 1813 5946 1865
rect 5894 1746 5946 1798
rect 5894 1679 5946 1731
rect 5894 1612 5946 1664
rect 5894 1545 5946 1597
rect 5894 1478 5946 1530
rect 5894 1411 5946 1463
rect 5894 1344 5946 1396
rect 5894 1277 5946 1329
rect 6050 2552 6102 2604
rect 6050 2485 6102 2537
rect 6050 2418 6102 2470
rect 6050 2351 6102 2403
rect 6050 2284 6102 2336
rect 6050 2217 6102 2269
rect 6050 2150 6102 2202
rect 6050 2083 6102 2135
rect 6050 2016 6102 2068
rect 6205 1813 6257 1865
rect 6205 1746 6257 1798
rect 6205 1679 6257 1731
rect 6205 1612 6257 1664
rect 6205 1545 6257 1597
rect 6205 1478 6257 1530
rect 6205 1411 6257 1463
rect 6205 1344 6257 1396
rect 6205 1277 6257 1329
rect 6361 2552 6413 2604
rect 6361 2485 6413 2537
rect 6361 2418 6413 2470
rect 6361 2351 6413 2403
rect 6361 2284 6413 2336
rect 6361 2217 6413 2269
rect 6361 2150 6413 2202
rect 6361 2083 6413 2135
rect 6361 2016 6413 2068
rect 6517 1813 6569 1865
rect 6517 1746 6569 1798
rect 6517 1679 6569 1731
rect 6517 1612 6569 1664
rect 6517 1545 6569 1597
rect 6517 1478 6569 1530
rect 6517 1411 6569 1463
rect 6517 1344 6569 1396
rect 6517 1277 6569 1329
rect 6673 2552 6725 2604
rect 6673 2485 6725 2537
rect 6673 2418 6725 2470
rect 6673 2351 6725 2403
rect 6673 2284 6725 2336
rect 6673 2217 6725 2269
rect 6673 2150 6725 2202
rect 6673 2083 6725 2135
rect 6673 2016 6725 2068
rect 6830 1813 6882 1865
rect 6830 1746 6882 1798
rect 6830 1679 6882 1731
rect 6830 1612 6882 1664
rect 6830 1545 6882 1597
rect 6830 1478 6882 1530
rect 6830 1411 6882 1463
rect 6830 1344 6882 1396
rect 6830 1277 6882 1329
rect 6986 2552 7038 2604
rect 6986 2485 7038 2537
rect 6986 2418 7038 2470
rect 6986 2351 7038 2403
rect 6986 2284 7038 2336
rect 6986 2217 7038 2269
rect 6986 2150 7038 2202
rect 6986 2083 7038 2135
rect 6986 2016 7038 2068
rect 7142 1813 7194 1865
rect 7142 1746 7194 1798
rect 7142 1679 7194 1731
rect 7142 1612 7194 1664
rect 7142 1545 7194 1597
rect 7142 1478 7194 1530
rect 7142 1411 7194 1463
rect 7142 1344 7194 1396
rect 7142 1277 7194 1329
rect 7298 2552 7350 2604
rect 7298 2485 7350 2537
rect 7298 2418 7350 2470
rect 7298 2351 7350 2403
rect 7298 2284 7350 2336
rect 7298 2217 7350 2269
rect 7298 2150 7350 2202
rect 7298 2083 7350 2135
rect 7298 2016 7350 2068
rect 7454 1813 7506 1865
rect 7454 1746 7506 1798
rect 7454 1679 7506 1731
rect 7454 1612 7506 1664
rect 7454 1545 7506 1597
rect 7454 1478 7506 1530
rect 7454 1411 7506 1463
rect 7454 1344 7506 1396
rect 7454 1277 7506 1329
rect 7610 2552 7662 2604
rect 7610 2485 7662 2537
rect 7610 2418 7662 2470
rect 7610 2351 7662 2403
rect 7610 2284 7662 2336
rect 7610 2217 7662 2269
rect 7610 2150 7662 2202
rect 7610 2083 7662 2135
rect 7610 2016 7662 2068
rect 7766 1813 7818 1865
rect 7766 1746 7818 1798
rect 7766 1679 7818 1731
rect 7766 1612 7818 1664
rect 7766 1545 7818 1597
rect 7766 1478 7818 1530
rect 7766 1411 7818 1463
rect 7766 1344 7818 1396
rect 7766 1277 7818 1329
rect 7922 2552 7974 2604
rect 7922 2485 7974 2537
rect 7922 2418 7974 2470
rect 7922 2351 7974 2403
rect 7922 2284 7974 2336
rect 7922 2217 7974 2269
rect 7922 2150 7974 2202
rect 7922 2083 7974 2135
rect 7922 2016 7974 2068
rect 8078 1813 8130 1865
rect 8078 1746 8130 1798
rect 8078 1679 8130 1731
rect 8078 1612 8130 1664
rect 8078 1545 8130 1597
rect 8078 1478 8130 1530
rect 8078 1411 8130 1463
rect 8078 1344 8130 1396
rect 8078 1277 8130 1329
rect 8234 2552 8286 2604
rect 8234 2485 8286 2537
rect 8234 2418 8286 2470
rect 8234 2351 8286 2403
rect 8234 2284 8286 2336
rect 8234 2217 8286 2269
rect 8234 2150 8286 2202
rect 8234 2083 8286 2135
rect 8234 2016 8286 2068
rect 8390 1813 8442 1865
rect 8390 1746 8442 1798
rect 8390 1679 8442 1731
rect 8390 1612 8442 1664
rect 8390 1545 8442 1597
rect 8390 1478 8442 1530
rect 8390 1411 8442 1463
rect 8390 1344 8442 1396
rect 8390 1277 8442 1329
rect 8546 2552 8598 2604
rect 8546 2485 8598 2537
rect 8546 2418 8598 2470
rect 8546 2351 8598 2403
rect 8546 2284 8598 2336
rect 8546 2217 8598 2269
rect 8546 2150 8598 2202
rect 8546 2083 8598 2135
rect 8546 2016 8598 2068
rect 8702 1813 8754 1865
rect 8702 1746 8754 1798
rect 8702 1679 8754 1731
rect 8702 1612 8754 1664
rect 8702 1545 8754 1597
rect 8702 1478 8754 1530
rect 8702 1411 8754 1463
rect 8702 1344 8754 1396
rect 8702 1277 8754 1329
rect 8858 2552 8910 2604
rect 8858 2485 8910 2537
rect 8858 2418 8910 2470
rect 8858 2351 8910 2403
rect 8858 2284 8910 2336
rect 8858 2217 8910 2269
rect 8858 2150 8910 2202
rect 8858 2083 8910 2135
rect 8858 2016 8910 2068
rect 9014 1813 9066 1865
rect 9014 1746 9066 1798
rect 9014 1679 9066 1731
rect 9014 1612 9066 1664
rect 9014 1545 9066 1597
rect 9014 1478 9066 1530
rect 9014 1411 9066 1463
rect 9014 1344 9066 1396
rect 9014 1277 9066 1329
rect 9170 2552 9222 2604
rect 9170 2485 9222 2537
rect 9170 2418 9222 2470
rect 9170 2351 9222 2403
rect 9170 2284 9222 2336
rect 9170 2217 9222 2269
rect 9170 2150 9222 2202
rect 9170 2083 9222 2135
rect 9170 2016 9222 2068
rect 9326 1813 9378 1865
rect 9326 1746 9378 1798
rect 9326 1679 9378 1731
rect 9326 1612 9378 1664
rect 9326 1545 9378 1597
rect 9326 1478 9378 1530
rect 9326 1411 9378 1463
rect 9326 1344 9378 1396
rect 9326 1277 9378 1329
rect 9482 2552 9534 2604
rect 9482 2485 9534 2537
rect 9482 2418 9534 2470
rect 9482 2351 9534 2403
rect 9482 2284 9534 2336
rect 9482 2217 9534 2269
rect 9482 2150 9534 2202
rect 9482 2083 9534 2135
rect 9482 2016 9534 2068
rect 9638 1813 9690 1865
rect 9638 1746 9690 1798
rect 9638 1679 9690 1731
rect 9638 1612 9690 1664
rect 9638 1545 9690 1597
rect 9638 1478 9690 1530
rect 9638 1411 9690 1463
rect 9638 1344 9690 1396
rect 9638 1277 9690 1329
rect 9794 2552 9846 2604
rect 9794 2485 9846 2537
rect 9794 2418 9846 2470
rect 9794 2351 9846 2403
rect 9794 2284 9846 2336
rect 9794 2217 9846 2269
rect 9794 2150 9846 2202
rect 9794 2083 9846 2135
rect 9794 2016 9846 2068
rect 9917 2603 9969 2604
rect 9917 2569 9923 2603
rect 9923 2569 9957 2603
rect 9957 2569 9969 2603
rect 9917 2552 9969 2569
rect 9983 2603 10035 2604
rect 9983 2569 9995 2603
rect 9995 2569 10029 2603
rect 10029 2569 10035 2603
rect 9983 2552 10035 2569
rect 9917 2496 9923 2522
rect 9923 2496 9957 2522
rect 9957 2496 9969 2522
rect 9917 2470 9969 2496
rect 9983 2496 9995 2522
rect 9995 2496 10029 2522
rect 10029 2496 10035 2522
rect 9983 2470 10035 2496
rect 9917 2423 9923 2440
rect 9923 2423 9957 2440
rect 9957 2423 9969 2440
rect 9917 2388 9969 2423
rect 9983 2423 9995 2440
rect 9995 2423 10029 2440
rect 10029 2423 10035 2440
rect 9983 2388 10035 2423
rect 9917 2305 9923 2357
rect 9923 2305 9969 2357
rect 9983 2305 10029 2357
rect 10029 2305 10035 2357
rect 9917 2222 9923 2274
rect 9923 2222 9969 2274
rect 9983 2222 10029 2274
rect 10029 2222 10035 2274
rect 9917 2139 9923 2191
rect 9923 2139 9969 2191
rect 9983 2139 10029 2191
rect 10029 2139 10035 2191
rect 9917 2056 9923 2108
rect 9923 2056 9969 2108
rect 9983 2056 10029 2108
rect 10029 2056 10035 2108
<< metal2 >>
rect -22 5770 -16 5822
rect 36 5770 48 5822
rect 100 5770 112 5822
rect 164 5770 176 5822
rect 228 5770 240 5822
rect 292 5770 304 5822
rect 356 5770 368 5822
rect 420 5770 432 5822
rect 484 5770 496 5822
rect 548 5770 560 5822
rect 612 5770 624 5822
rect 676 5770 688 5822
rect 740 5770 752 5822
rect 804 5770 816 5822
rect 868 5770 880 5822
rect 932 5770 944 5822
rect 996 5770 1008 5822
rect 1060 5770 1072 5822
rect 1124 5770 1136 5822
rect 1188 5770 1200 5822
rect 1252 5770 1264 5822
rect 1316 5770 1328 5822
rect 1380 5770 1392 5822
rect 1444 5770 1456 5822
rect 1508 5770 1520 5822
rect 1572 5770 1584 5822
rect 1636 5770 1648 5822
rect 1700 5770 1712 5822
rect 1764 5770 1776 5822
rect 1828 5770 1840 5822
rect 1892 5770 1904 5822
rect 1956 5770 1968 5822
rect 2020 5770 2032 5822
rect 2084 5770 2096 5822
rect 2148 5770 2160 5822
rect 2212 5770 2224 5822
rect 2276 5770 2288 5822
rect 2340 5770 2352 5822
rect 2404 5770 2416 5822
rect 2468 5770 2480 5822
rect 2532 5770 2544 5822
rect 2596 5770 2608 5822
rect 2660 5770 2672 5822
rect 2724 5770 2736 5822
rect 2788 5770 2800 5822
rect 2852 5770 2864 5822
rect 2916 5770 2928 5822
rect 2980 5770 2992 5822
rect 3044 5770 3056 5822
rect 3108 5770 3120 5822
rect 3172 5770 3184 5822
rect 3236 5770 3248 5822
rect 3300 5770 3312 5822
rect 3364 5770 3376 5822
rect 3428 5770 3440 5822
rect 3492 5770 3504 5822
rect 3556 5770 3568 5822
rect 3620 5770 3632 5822
rect 3684 5770 3696 5822
rect 3748 5770 3760 5822
rect 3812 5770 3824 5822
rect 3876 5770 3888 5822
rect 3940 5770 3952 5822
rect 4004 5770 4016 5822
rect 4068 5770 4080 5822
rect 4132 5770 4144 5822
rect 4196 5770 4208 5822
rect 4260 5770 4272 5822
rect 4324 5770 4336 5822
rect 4388 5770 4400 5822
rect 4452 5770 4464 5822
rect 4516 5770 4528 5822
rect 4580 5770 4592 5822
rect 4644 5770 4656 5822
rect 4708 5770 4720 5822
rect 4772 5770 4784 5822
rect 4836 5770 4848 5822
rect 4900 5770 4912 5822
rect 4964 5770 4976 5822
rect 5028 5770 5040 5822
rect 5092 5770 5104 5822
rect 5156 5770 5168 5822
rect 5220 5770 5232 5822
rect 5284 5770 5296 5822
rect 5348 5770 5360 5822
rect 5412 5770 5424 5822
rect 5476 5770 5488 5822
rect 5540 5770 5552 5822
rect 5604 5770 5616 5822
rect 5668 5770 5680 5822
rect 5732 5770 5744 5822
rect 5796 5770 5808 5822
rect 5860 5770 5872 5822
rect 5924 5770 5936 5822
rect 5988 5770 6000 5822
rect 6052 5770 6064 5822
rect 6116 5770 6128 5822
rect 6180 5770 6192 5822
rect 6244 5770 6256 5822
rect 6308 5770 6320 5822
rect 6372 5770 6384 5822
rect 6436 5770 6448 5822
rect 6500 5770 6512 5822
rect 6564 5770 6576 5822
rect 6628 5770 6640 5822
rect 6692 5770 6704 5822
rect 6756 5770 6768 5822
rect 6820 5770 6832 5822
rect 6884 5770 6896 5822
rect 6948 5770 6960 5822
rect 7012 5770 7024 5822
rect 7076 5770 7088 5822
rect 7140 5770 7152 5822
rect 7204 5770 7216 5822
rect 7268 5770 7280 5822
rect 7332 5770 7344 5822
rect 7396 5770 7408 5822
rect 7460 5770 7472 5822
rect 7524 5770 7536 5822
rect 7588 5770 7600 5822
rect 7652 5770 7664 5822
rect 7716 5770 7728 5822
rect 7780 5770 7792 5822
rect 7844 5770 7856 5822
rect 7908 5770 7920 5822
rect 7972 5770 7984 5822
rect 8036 5770 8048 5822
rect 8100 5770 8112 5822
rect 8164 5770 8176 5822
rect 8228 5770 8240 5822
rect 8292 5770 8304 5822
rect 8356 5770 8368 5822
rect 8420 5770 8432 5822
rect 8484 5770 8496 5822
rect 8548 5770 8560 5822
rect 8612 5770 8624 5822
rect 8676 5770 8688 5822
rect 8740 5770 8752 5822
rect 8804 5770 8816 5822
rect 8868 5770 8880 5822
rect 8932 5770 8944 5822
rect 8996 5770 9008 5822
rect 9060 5770 9072 5822
rect 9124 5770 9136 5822
rect 9188 5770 9200 5822
rect 9252 5770 9264 5822
rect 9316 5770 9329 5822
rect 9381 5770 9394 5822
rect 9446 5770 9459 5822
rect 9511 5770 9524 5822
rect 9576 5770 9589 5822
rect 9641 5770 9654 5822
rect 9706 5770 9719 5822
rect 9771 5770 9784 5822
rect 9836 5770 9849 5822
rect 9901 5770 9914 5822
rect 9966 5770 9979 5822
rect 10031 5770 10044 5822
rect 10096 5770 10109 5822
rect 10161 5770 10174 5822
rect 10226 5770 10239 5822
rect 10291 5770 10499 5822
rect -22 5756 10499 5770
rect -22 5704 -16 5756
rect 36 5704 48 5756
rect 100 5704 112 5756
rect 164 5704 176 5756
rect 228 5704 240 5756
rect 292 5704 304 5756
rect 356 5704 368 5756
rect 420 5704 432 5756
rect 484 5704 496 5756
rect 548 5704 560 5756
rect 612 5704 624 5756
rect 676 5704 688 5756
rect 740 5704 752 5756
rect 804 5704 816 5756
rect 868 5704 880 5756
rect 932 5704 944 5756
rect 996 5704 1008 5756
rect 1060 5704 1072 5756
rect 1124 5704 1136 5756
rect 1188 5704 1200 5756
rect 1252 5704 1264 5756
rect 1316 5704 1328 5756
rect 1380 5704 1392 5756
rect 1444 5704 1456 5756
rect 1508 5704 1520 5756
rect 1572 5704 1584 5756
rect 1636 5704 1648 5756
rect 1700 5704 1712 5756
rect 1764 5704 1776 5756
rect 1828 5704 1840 5756
rect 1892 5704 1904 5756
rect 1956 5704 1968 5756
rect 2020 5704 2032 5756
rect 2084 5704 2096 5756
rect 2148 5704 2160 5756
rect 2212 5704 2224 5756
rect 2276 5704 2288 5756
rect 2340 5704 2352 5756
rect 2404 5704 2416 5756
rect 2468 5704 2480 5756
rect 2532 5704 2544 5756
rect 2596 5704 2608 5756
rect 2660 5704 2672 5756
rect 2724 5704 2736 5756
rect 2788 5704 2800 5756
rect 2852 5704 2864 5756
rect 2916 5704 2928 5756
rect 2980 5704 2992 5756
rect 3044 5704 3056 5756
rect 3108 5704 3120 5756
rect 3172 5704 3184 5756
rect 3236 5704 3248 5756
rect 3300 5704 3312 5756
rect 3364 5704 3376 5756
rect 3428 5704 3440 5756
rect 3492 5704 3504 5756
rect 3556 5704 3568 5756
rect 3620 5704 3632 5756
rect 3684 5704 3696 5756
rect 3748 5704 3760 5756
rect 3812 5704 3824 5756
rect 3876 5704 3888 5756
rect 3940 5704 3952 5756
rect 4004 5704 4016 5756
rect 4068 5704 4080 5756
rect 4132 5704 4144 5756
rect 4196 5704 4208 5756
rect 4260 5704 4272 5756
rect 4324 5704 4336 5756
rect 4388 5704 4400 5756
rect 4452 5704 4464 5756
rect 4516 5704 4528 5756
rect 4580 5704 4592 5756
rect 4644 5704 4656 5756
rect 4708 5704 4720 5756
rect 4772 5704 4784 5756
rect 4836 5704 4848 5756
rect 4900 5704 4912 5756
rect 4964 5704 4976 5756
rect 5028 5704 5040 5756
rect 5092 5704 5104 5756
rect 5156 5704 5168 5756
rect 5220 5704 5232 5756
rect 5284 5704 5296 5756
rect 5348 5704 5360 5756
rect 5412 5704 5424 5756
rect 5476 5704 5488 5756
rect 5540 5704 5552 5756
rect 5604 5704 5616 5756
rect 5668 5704 5680 5756
rect 5732 5704 5744 5756
rect 5796 5704 5808 5756
rect 5860 5704 5872 5756
rect 5924 5704 5936 5756
rect 5988 5704 6000 5756
rect 6052 5704 6064 5756
rect 6116 5704 6128 5756
rect 6180 5704 6192 5756
rect 6244 5704 6256 5756
rect 6308 5704 6320 5756
rect 6372 5704 6384 5756
rect 6436 5704 6448 5756
rect 6500 5704 6512 5756
rect 6564 5704 6576 5756
rect 6628 5704 6640 5756
rect 6692 5704 6704 5756
rect 6756 5704 6768 5756
rect 6820 5704 6832 5756
rect 6884 5704 6896 5756
rect 6948 5704 6960 5756
rect 7012 5704 7024 5756
rect 7076 5704 7088 5756
rect 7140 5704 7152 5756
rect 7204 5704 7216 5756
rect 7268 5704 7280 5756
rect 7332 5704 7344 5756
rect 7396 5704 7408 5756
rect 7460 5704 7472 5756
rect 7524 5704 7536 5756
rect 7588 5704 7600 5756
rect 7652 5704 7664 5756
rect 7716 5704 7728 5756
rect 7780 5704 7792 5756
rect 7844 5704 7856 5756
rect 7908 5704 7920 5756
rect 7972 5704 7984 5756
rect 8036 5704 8048 5756
rect 8100 5704 8112 5756
rect 8164 5704 8176 5756
rect 8228 5704 8240 5756
rect 8292 5704 8304 5756
rect 8356 5704 8368 5756
rect 8420 5704 8432 5756
rect 8484 5704 8496 5756
rect 8548 5704 8560 5756
rect 8612 5704 8624 5756
rect 8676 5704 8688 5756
rect 8740 5704 8752 5756
rect 8804 5704 8816 5756
rect 8868 5704 8880 5756
rect 8932 5704 8944 5756
rect 8996 5704 9008 5756
rect 9060 5704 9072 5756
rect 9124 5704 9136 5756
rect 9188 5704 9200 5756
rect 9252 5704 9264 5756
rect 9316 5704 9329 5756
rect 9381 5704 9394 5756
rect 9446 5704 9459 5756
rect 9511 5704 9524 5756
rect 9576 5704 9589 5756
rect 9641 5704 9654 5756
rect 9706 5704 9719 5756
rect 9771 5704 9784 5756
rect 9836 5704 9849 5756
rect 9901 5704 9914 5756
rect 9966 5704 9979 5756
rect 10031 5704 10044 5756
rect 10096 5704 10109 5756
rect 10161 5704 10174 5756
rect 10226 5704 10239 5756
rect 10291 5704 10499 5756
rect -22 5280 10499 5704
rect -22 5228 525 5280
rect 577 5228 658 5280
rect 710 5228 791 5280
rect 843 5228 923 5280
rect 975 5228 1055 5280
rect 1107 5228 1187 5280
rect 1239 5228 1319 5280
rect 1371 5228 1451 5280
rect 1503 5228 1583 5280
rect 1635 5228 1715 5280
rect 1767 5228 1847 5280
rect 1899 5228 1979 5280
rect 2031 5228 2111 5280
rect 2163 5228 2243 5280
rect 2295 5228 2375 5280
rect 2427 5228 2507 5280
rect 2559 5228 2639 5280
rect 2691 5228 2771 5280
rect 2823 5228 2903 5280
rect 2955 5228 3035 5280
rect 3087 5228 10499 5280
rect -22 5214 10499 5228
rect -22 5162 525 5214
rect 577 5162 658 5214
rect 710 5162 791 5214
rect 843 5162 923 5214
rect 975 5162 1055 5214
rect 1107 5162 1187 5214
rect 1239 5162 1319 5214
rect 1371 5162 1451 5214
rect 1503 5162 1583 5214
rect 1635 5162 1715 5214
rect 1767 5162 1847 5214
rect 1899 5162 1979 5214
rect 2031 5162 2111 5214
rect 2163 5162 2243 5214
rect 2295 5162 2375 5214
rect 2427 5162 2507 5214
rect 2559 5162 2639 5214
rect 2691 5162 2771 5214
rect 2823 5162 2903 5214
rect 2955 5162 3035 5214
rect 3087 5162 10499 5214
rect 686 4891 3210 4943
rect 3262 4891 3274 4943
rect 3326 4891 9848 4943
rect 686 4854 9848 4860
rect 686 4802 844 4854
rect 896 4802 1156 4854
rect 1208 4802 1468 4854
rect 1520 4802 1780 4854
rect 1832 4802 2092 4854
rect 2144 4802 2404 4854
rect 2456 4802 2716 4854
rect 2768 4802 5270 4854
rect 5322 4802 5582 4854
rect 5634 4802 5894 4854
rect 5946 4802 6205 4854
rect 6257 4802 6517 4854
rect 6569 4802 6830 4854
rect 6882 4802 7142 4854
rect 7194 4802 7454 4854
rect 7506 4802 7766 4854
rect 7818 4802 8078 4854
rect 8130 4802 8390 4854
rect 8442 4802 8702 4854
rect 8754 4802 9014 4854
rect 9066 4802 9326 4854
rect 9378 4802 9638 4854
rect 9690 4802 9848 4854
rect 686 4787 9848 4802
rect 686 4735 844 4787
rect 896 4735 1156 4787
rect 1208 4735 1468 4787
rect 1520 4735 1780 4787
rect 1832 4735 2092 4787
rect 2144 4735 2404 4787
rect 2456 4735 2716 4787
rect 2768 4735 5270 4787
rect 5322 4735 5582 4787
rect 5634 4735 5894 4787
rect 5946 4735 6205 4787
rect 6257 4735 6517 4787
rect 6569 4735 6830 4787
rect 6882 4735 7142 4787
rect 7194 4735 7454 4787
rect 7506 4735 7766 4787
rect 7818 4735 8078 4787
rect 8130 4735 8390 4787
rect 8442 4735 8702 4787
rect 8754 4735 9014 4787
rect 9066 4735 9326 4787
rect 9378 4735 9638 4787
rect 9690 4735 9848 4787
rect 686 4720 9848 4735
rect 686 4668 844 4720
rect 896 4668 1156 4720
rect 1208 4668 1468 4720
rect 1520 4668 1780 4720
rect 1832 4668 2092 4720
rect 2144 4668 2404 4720
rect 2456 4668 2716 4720
rect 2768 4668 5270 4720
rect 5322 4668 5582 4720
rect 5634 4668 5894 4720
rect 5946 4668 6205 4720
rect 6257 4668 6517 4720
rect 6569 4668 6830 4720
rect 6882 4668 7142 4720
rect 7194 4668 7454 4720
rect 7506 4668 7766 4720
rect 7818 4668 8078 4720
rect 8130 4668 8390 4720
rect 8442 4668 8702 4720
rect 8754 4668 9014 4720
rect 9066 4668 9326 4720
rect 9378 4668 9638 4720
rect 9690 4668 9848 4720
rect 686 4653 9848 4668
rect 686 4601 844 4653
rect 896 4601 1156 4653
rect 1208 4601 1468 4653
rect 1520 4601 1780 4653
rect 1832 4601 2092 4653
rect 2144 4601 2404 4653
rect 2456 4601 2716 4653
rect 2768 4601 5270 4653
rect 5322 4601 5582 4653
rect 5634 4601 5894 4653
rect 5946 4601 6205 4653
rect 6257 4601 6517 4653
rect 6569 4601 6830 4653
rect 6882 4601 7142 4653
rect 7194 4601 7454 4653
rect 7506 4601 7766 4653
rect 7818 4601 8078 4653
rect 8130 4601 8390 4653
rect 8442 4601 8702 4653
rect 8754 4601 9014 4653
rect 9066 4601 9326 4653
rect 9378 4601 9638 4653
rect 9690 4601 9848 4653
rect 686 4586 9848 4601
rect 686 4534 844 4586
rect 896 4534 1156 4586
rect 1208 4534 1468 4586
rect 1520 4534 1780 4586
rect 1832 4534 2092 4586
rect 2144 4534 2404 4586
rect 2456 4534 2716 4586
rect 2768 4534 5270 4586
rect 5322 4534 5582 4586
rect 5634 4534 5894 4586
rect 5946 4534 6205 4586
rect 6257 4534 6517 4586
rect 6569 4534 6830 4586
rect 6882 4534 7142 4586
rect 7194 4534 7454 4586
rect 7506 4534 7766 4586
rect 7818 4534 8078 4586
rect 8130 4534 8390 4586
rect 8442 4534 8702 4586
rect 8754 4534 9014 4586
rect 9066 4534 9326 4586
rect 9378 4534 9638 4586
rect 9690 4534 9848 4586
rect 686 4519 9848 4534
rect 686 4467 844 4519
rect 896 4467 1156 4519
rect 1208 4467 1468 4519
rect 1520 4467 1780 4519
rect 1832 4467 2092 4519
rect 2144 4467 2404 4519
rect 2456 4467 2716 4519
rect 2768 4467 5270 4519
rect 5322 4467 5582 4519
rect 5634 4467 5894 4519
rect 5946 4467 6205 4519
rect 6257 4467 6517 4519
rect 6569 4467 6830 4519
rect 6882 4467 7142 4519
rect 7194 4467 7454 4519
rect 7506 4467 7766 4519
rect 7818 4467 8078 4519
rect 8130 4467 8390 4519
rect 8442 4467 8702 4519
rect 8754 4467 9014 4519
rect 9066 4467 9326 4519
rect 9378 4467 9638 4519
rect 9690 4467 9848 4519
rect 686 4452 9848 4467
rect 686 4400 844 4452
rect 896 4400 1156 4452
rect 1208 4400 1468 4452
rect 1520 4400 1780 4452
rect 1832 4400 2092 4452
rect 2144 4400 2404 4452
rect 2456 4400 2716 4452
rect 2768 4400 5270 4452
rect 5322 4400 5582 4452
rect 5634 4400 5894 4452
rect 5946 4400 6205 4452
rect 6257 4400 6517 4452
rect 6569 4400 6830 4452
rect 6882 4400 7142 4452
rect 7194 4400 7454 4452
rect 7506 4400 7766 4452
rect 7818 4400 8078 4452
rect 8130 4400 8390 4452
rect 8442 4400 8702 4452
rect 8754 4400 9014 4452
rect 9066 4400 9326 4452
rect 9378 4400 9638 4452
rect 9690 4400 9848 4452
rect 686 4385 9848 4400
rect 686 4333 844 4385
rect 896 4333 1156 4385
rect 1208 4333 1468 4385
rect 1520 4333 1780 4385
rect 1832 4333 2092 4385
rect 2144 4333 2404 4385
rect 2456 4333 2716 4385
rect 2768 4333 5270 4385
rect 5322 4333 5582 4385
rect 5634 4333 5894 4385
rect 5946 4333 6205 4385
rect 6257 4333 6517 4385
rect 6569 4333 6830 4385
rect 6882 4333 7142 4385
rect 7194 4333 7454 4385
rect 7506 4333 7766 4385
rect 7818 4333 8078 4385
rect 8130 4333 8390 4385
rect 8442 4333 8702 4385
rect 8754 4333 9014 4385
rect 9066 4333 9326 4385
rect 9378 4333 9638 4385
rect 9690 4333 9848 4385
rect 686 4318 9848 4333
rect 686 4266 844 4318
rect 896 4266 1156 4318
rect 1208 4266 1468 4318
rect 1520 4266 1780 4318
rect 1832 4266 2092 4318
rect 2144 4266 2404 4318
rect 2456 4266 2716 4318
rect 2768 4266 5270 4318
rect 5322 4266 5582 4318
rect 5634 4266 5894 4318
rect 5946 4266 6205 4318
rect 6257 4266 6517 4318
rect 6569 4266 6830 4318
rect 6882 4266 7142 4318
rect 7194 4266 7454 4318
rect 7506 4266 7766 4318
rect 7818 4266 8078 4318
rect 8130 4266 8390 4318
rect 8442 4266 8702 4318
rect 8754 4266 9014 4318
rect 9066 4266 9326 4318
rect 9378 4266 9638 4318
rect 9690 4266 9848 4318
rect 686 4260 9848 4266
rect 686 4176 3210 4228
rect 3262 4176 3274 4228
rect 3326 4176 9848 4228
rect 144 4114 10035 4120
rect 144 4062 688 4114
rect 740 4062 1000 4114
rect 1052 4062 1312 4114
rect 1364 4062 1624 4114
rect 1676 4062 1936 4114
rect 1988 4062 2248 4114
rect 2300 4062 2560 4114
rect 2612 4062 2872 4114
rect 2924 4062 4925 4114
rect 4977 4062 4991 4114
rect 5043 4062 5114 4114
rect 5166 4062 5426 4114
rect 5478 4062 5738 4114
rect 5790 4062 6050 4114
rect 6102 4062 6361 4114
rect 6413 4062 6673 4114
rect 6725 4062 6986 4114
rect 7038 4062 7298 4114
rect 7350 4062 7610 4114
rect 7662 4062 7922 4114
rect 7974 4062 8234 4114
rect 8286 4062 8546 4114
rect 8598 4062 8858 4114
rect 8910 4062 9170 4114
rect 9222 4062 9482 4114
rect 9534 4062 9794 4114
rect 9846 4062 9917 4114
rect 9969 4062 9983 4114
rect 144 4047 10035 4062
rect 144 3995 688 4047
rect 740 3995 1000 4047
rect 1052 3995 1312 4047
rect 1364 3995 1624 4047
rect 1676 3995 1936 4047
rect 1988 3995 2248 4047
rect 2300 3995 2560 4047
rect 2612 3995 2872 4047
rect 2924 4025 5114 4047
rect 2924 3995 4925 4025
rect 144 3980 4925 3995
rect 144 3928 688 3980
rect 740 3928 1000 3980
rect 1052 3928 1312 3980
rect 1364 3928 1624 3980
rect 1676 3928 1936 3980
rect 1988 3928 2248 3980
rect 2300 3928 2560 3980
rect 2612 3928 2872 3980
rect 2924 3973 4925 3980
rect 4977 3973 4991 4025
rect 5043 3995 5114 4025
rect 5166 3995 5426 4047
rect 5478 3995 5738 4047
rect 5790 3995 6050 4047
rect 6102 3995 6361 4047
rect 6413 3995 6673 4047
rect 6725 3995 6986 4047
rect 7038 3995 7298 4047
rect 7350 3995 7610 4047
rect 7662 3995 7922 4047
rect 7974 3995 8234 4047
rect 8286 3995 8546 4047
rect 8598 3995 8858 4047
rect 8910 3995 9170 4047
rect 9222 3995 9482 4047
rect 9534 3995 9794 4047
rect 9846 4025 10035 4047
rect 9846 3995 9917 4025
rect 5043 3980 9917 3995
rect 5043 3973 5114 3980
rect 2924 3936 5114 3973
rect 2924 3928 4925 3936
rect 144 3913 4925 3928
rect 144 3861 688 3913
rect 740 3861 1000 3913
rect 1052 3861 1312 3913
rect 1364 3861 1624 3913
rect 1676 3861 1936 3913
rect 1988 3861 2248 3913
rect 2300 3861 2560 3913
rect 2612 3861 2872 3913
rect 2924 3884 4925 3913
rect 4977 3884 4991 3936
rect 5043 3928 5114 3936
rect 5166 3928 5426 3980
rect 5478 3928 5738 3980
rect 5790 3928 6050 3980
rect 6102 3928 6361 3980
rect 6413 3928 6673 3980
rect 6725 3928 6986 3980
rect 7038 3928 7298 3980
rect 7350 3928 7610 3980
rect 7662 3928 7922 3980
rect 7974 3928 8234 3980
rect 8286 3928 8546 3980
rect 8598 3928 8858 3980
rect 8910 3928 9170 3980
rect 9222 3928 9482 3980
rect 9534 3928 9794 3980
rect 9846 3973 9917 3980
rect 9969 3973 9983 4025
rect 9846 3936 10035 3973
rect 9846 3928 9917 3936
rect 5043 3913 9917 3928
rect 5043 3884 5114 3913
rect 2924 3861 5114 3884
rect 5166 3861 5426 3913
rect 5478 3861 5738 3913
rect 5790 3861 6050 3913
rect 6102 3861 6361 3913
rect 6413 3861 6673 3913
rect 6725 3861 6986 3913
rect 7038 3861 7298 3913
rect 7350 3861 7610 3913
rect 7662 3861 7922 3913
rect 7974 3861 8234 3913
rect 8286 3861 8546 3913
rect 8598 3861 8858 3913
rect 8910 3861 9170 3913
rect 9222 3861 9482 3913
rect 9534 3861 9794 3913
rect 9846 3884 9917 3913
rect 9969 3884 9983 3936
rect 9846 3861 10035 3884
rect 144 3847 10035 3861
rect 144 3846 4925 3847
rect 144 3794 688 3846
rect 740 3794 1000 3846
rect 1052 3794 1312 3846
rect 1364 3794 1624 3846
rect 1676 3794 1936 3846
rect 1988 3794 2248 3846
rect 2300 3794 2560 3846
rect 2612 3794 2872 3846
rect 2924 3795 4925 3846
rect 4977 3795 4991 3847
rect 5043 3846 9917 3847
rect 5043 3795 5114 3846
rect 2924 3794 5114 3795
rect 5166 3794 5426 3846
rect 5478 3794 5738 3846
rect 5790 3794 6050 3846
rect 6102 3794 6361 3846
rect 6413 3794 6673 3846
rect 6725 3794 6986 3846
rect 7038 3794 7298 3846
rect 7350 3794 7610 3846
rect 7662 3794 7922 3846
rect 7974 3794 8234 3846
rect 8286 3794 8546 3846
rect 8598 3794 8858 3846
rect 8910 3794 9170 3846
rect 9222 3794 9482 3846
rect 9534 3794 9794 3846
rect 9846 3795 9917 3846
rect 9969 3795 9983 3847
rect 9846 3794 10035 3795
rect 144 3779 10035 3794
rect 144 3727 688 3779
rect 740 3727 1000 3779
rect 1052 3727 1312 3779
rect 1364 3727 1624 3779
rect 1676 3727 1936 3779
rect 1988 3727 2248 3779
rect 2300 3727 2560 3779
rect 2612 3727 2872 3779
rect 2924 3758 5114 3779
rect 2924 3727 4925 3758
rect 144 3712 4925 3727
rect 144 3660 688 3712
rect 740 3660 1000 3712
rect 1052 3660 1312 3712
rect 1364 3660 1624 3712
rect 1676 3660 1936 3712
rect 1988 3660 2248 3712
rect 2300 3660 2560 3712
rect 2612 3660 2872 3712
rect 2924 3706 4925 3712
rect 4977 3706 4991 3758
rect 5043 3727 5114 3758
rect 5166 3727 5426 3779
rect 5478 3727 5738 3779
rect 5790 3727 6050 3779
rect 6102 3727 6361 3779
rect 6413 3727 6673 3779
rect 6725 3727 6986 3779
rect 7038 3727 7298 3779
rect 7350 3727 7610 3779
rect 7662 3727 7922 3779
rect 7974 3727 8234 3779
rect 8286 3727 8546 3779
rect 8598 3727 8858 3779
rect 8910 3727 9170 3779
rect 9222 3727 9482 3779
rect 9534 3727 9794 3779
rect 9846 3758 10035 3779
rect 9846 3727 9917 3758
rect 5043 3712 9917 3727
rect 5043 3706 5114 3712
rect 2924 3668 5114 3706
rect 2924 3660 4925 3668
rect 144 3645 4925 3660
rect 144 3593 688 3645
rect 740 3593 1000 3645
rect 1052 3593 1312 3645
rect 1364 3593 1624 3645
rect 1676 3593 1936 3645
rect 1988 3593 2248 3645
rect 2300 3593 2560 3645
rect 2612 3593 2872 3645
rect 2924 3616 4925 3645
rect 4977 3616 4991 3668
rect 5043 3660 5114 3668
rect 5166 3660 5426 3712
rect 5478 3660 5738 3712
rect 5790 3660 6050 3712
rect 6102 3660 6361 3712
rect 6413 3660 6673 3712
rect 6725 3660 6986 3712
rect 7038 3660 7298 3712
rect 7350 3660 7610 3712
rect 7662 3660 7922 3712
rect 7974 3660 8234 3712
rect 8286 3660 8546 3712
rect 8598 3660 8858 3712
rect 8910 3660 9170 3712
rect 9222 3660 9482 3712
rect 9534 3660 9794 3712
rect 9846 3706 9917 3712
rect 9969 3706 9983 3758
rect 9846 3668 10035 3706
rect 9846 3660 9917 3668
rect 5043 3645 9917 3660
rect 5043 3616 5114 3645
rect 2924 3593 5114 3616
rect 5166 3593 5426 3645
rect 5478 3593 5738 3645
rect 5790 3593 6050 3645
rect 6102 3593 6361 3645
rect 6413 3593 6673 3645
rect 6725 3593 6986 3645
rect 7038 3593 7298 3645
rect 7350 3593 7610 3645
rect 7662 3593 7922 3645
rect 7974 3593 8234 3645
rect 8286 3593 8546 3645
rect 8598 3593 8858 3645
rect 8910 3593 9170 3645
rect 9222 3593 9482 3645
rect 9534 3593 9794 3645
rect 9846 3616 9917 3645
rect 9969 3616 9983 3668
rect 9846 3593 10035 3616
rect 144 3578 10035 3593
rect 144 3526 688 3578
rect 740 3526 1000 3578
rect 1052 3526 1312 3578
rect 1364 3526 1624 3578
rect 1676 3526 1936 3578
rect 1988 3526 2248 3578
rect 2300 3526 2560 3578
rect 2612 3526 2872 3578
rect 2924 3526 4925 3578
rect 4977 3526 4991 3578
rect 5043 3526 5114 3578
rect 5166 3526 5426 3578
rect 5478 3526 5738 3578
rect 5790 3526 6050 3578
rect 6102 3526 6361 3578
rect 6413 3526 6673 3578
rect 6725 3526 6986 3578
rect 7038 3526 7298 3578
rect 7350 3526 7610 3578
rect 7662 3526 7922 3578
rect 7974 3526 8234 3578
rect 8286 3526 8546 3578
rect 8598 3526 8858 3578
rect 8910 3526 9170 3578
rect 9222 3526 9482 3578
rect 9534 3526 9794 3578
rect 9846 3526 9917 3578
rect 9969 3526 9983 3578
rect 144 3520 10035 3526
rect 144 2755 694 3520
tri 694 3282 932 3520 nw
rect 5297 3173 5303 3225
rect 5355 3173 5367 3225
rect 5419 3173 5431 3225
rect 5483 3173 5495 3225
rect 5547 3173 5559 3225
rect 5611 3173 5623 3225
rect 5675 3173 5687 3225
rect 5739 3173 5751 3225
rect 5803 3173 5815 3225
rect 5867 3173 5879 3225
rect 5931 3173 5943 3225
rect 5995 3173 6007 3225
rect 6059 3173 6071 3225
rect 6123 3173 6135 3225
rect 6187 3173 6199 3225
rect 6251 3173 6263 3225
rect 6315 3173 6327 3225
rect 6379 3173 6391 3225
rect 6443 3173 6456 3225
rect 6508 3173 6521 3225
rect 6573 3173 6586 3225
rect 6638 3173 6651 3225
rect 6703 3173 6716 3225
rect 6768 3173 6781 3225
rect 6833 3173 6846 3225
rect 6898 3173 6911 3225
rect 6963 3173 6976 3225
rect 7028 3173 7041 3225
rect 7093 3173 7106 3225
rect 7158 3173 7171 3225
rect 7223 3173 7236 3225
rect 7288 3173 7301 3225
rect 7353 3173 7366 3225
rect 7418 3173 7431 3225
rect 7483 3173 7496 3225
rect 7548 3173 7561 3225
rect 7613 3173 7626 3225
rect 7678 3173 7691 3225
rect 7743 3173 7756 3225
rect 7808 3173 7821 3225
rect 7873 3173 7886 3225
rect 7938 3173 7951 3225
rect 8003 3173 8016 3225
rect 8068 3173 8081 3225
rect 8133 3173 8146 3225
rect 8198 3173 8211 3225
rect 8263 3173 8276 3225
rect 8328 3173 8341 3225
rect 8393 3173 8406 3225
rect 8458 3173 8471 3225
rect 8523 3173 8536 3225
rect 8588 3173 8601 3225
rect 8653 3173 8666 3225
rect 8718 3173 8731 3225
rect 8783 3173 8796 3225
rect 8848 3173 8861 3225
rect 8913 3173 8926 3225
rect 8978 3173 8991 3225
rect 9043 3173 9056 3225
rect 9108 3173 9121 3225
rect 9173 3173 9186 3225
rect 9238 3173 9251 3225
rect 9303 3173 9316 3225
rect 9368 3173 9381 3225
rect 9433 3173 9446 3225
rect 9498 3173 9504 3225
rect 1329 2997 1335 3049
rect 1387 2997 1471 3049
rect 1523 2997 1607 3049
rect 1659 2997 1743 3049
rect 1795 2997 1879 3049
rect 1931 2997 2015 3049
rect 2067 2997 2151 3049
rect 2203 2997 2287 3049
rect 2339 2997 2423 3049
rect 2475 2997 2560 3049
rect 2612 2997 2697 3049
rect 2749 2997 2755 3049
rect 1329 2878 1335 2930
rect 1387 2878 1471 2930
rect 1523 2878 1607 2930
rect 1659 2878 1743 2930
rect 1795 2878 1879 2930
rect 1931 2878 2015 2930
rect 2067 2878 2151 2930
rect 2203 2878 2287 2930
rect 2339 2878 2423 2930
rect 2475 2878 2560 2930
rect 2612 2878 2697 2930
rect 2749 2878 2755 2930
tri 694 2755 787 2848 sw
rect 144 2703 787 2755
tri 787 2703 839 2755 sw
rect 3979 2703 3985 2755
rect 4037 2703 4165 2755
rect 4217 2703 4223 2755
rect 5297 2703 5303 2755
rect 5355 2703 5367 2755
rect 5419 2703 5431 2755
rect 5483 2703 5495 2755
rect 5547 2703 5559 2755
rect 5611 2703 5623 2755
rect 5675 2703 5687 2755
rect 5739 2703 5751 2755
rect 5803 2703 5815 2755
rect 5867 2703 5879 2755
rect 5931 2703 5943 2755
rect 5995 2703 6007 2755
rect 6059 2703 6071 2755
rect 6123 2703 6135 2755
rect 6187 2703 6199 2755
rect 6251 2703 6263 2755
rect 6315 2703 6327 2755
rect 6379 2703 6391 2755
rect 6443 2703 6456 2755
rect 6508 2703 6521 2755
rect 6573 2703 6586 2755
rect 6638 2703 6651 2755
rect 6703 2703 6716 2755
rect 6768 2703 6781 2755
rect 6833 2703 6846 2755
rect 6898 2703 6911 2755
rect 6963 2703 6976 2755
rect 7028 2703 7041 2755
rect 7093 2703 7106 2755
rect 7158 2703 7171 2755
rect 7223 2703 7236 2755
rect 7288 2703 7301 2755
rect 7353 2703 7366 2755
rect 7418 2703 7431 2755
rect 7483 2703 7496 2755
rect 7548 2703 7561 2755
rect 7613 2703 7626 2755
rect 7678 2703 7691 2755
rect 7743 2703 7756 2755
rect 7808 2703 7821 2755
rect 7873 2703 7886 2755
rect 7938 2703 7951 2755
rect 8003 2703 8016 2755
rect 8068 2703 8081 2755
rect 8133 2703 8146 2755
rect 8198 2703 8211 2755
rect 8263 2703 8276 2755
rect 8328 2703 8341 2755
rect 8393 2703 8406 2755
rect 8458 2703 8471 2755
rect 8523 2703 8536 2755
rect 8588 2703 8601 2755
rect 8653 2703 8666 2755
rect 8718 2703 8731 2755
rect 8783 2703 8796 2755
rect 8848 2703 8861 2755
rect 8913 2703 8926 2755
rect 8978 2703 8991 2755
rect 9043 2703 9056 2755
rect 9108 2703 9121 2755
rect 9173 2703 9186 2755
rect 9238 2703 9251 2755
rect 9303 2703 9316 2755
rect 9368 2703 9381 2755
rect 9433 2703 9446 2755
rect 9498 2703 9504 2755
rect 144 2610 839 2703
tri 839 2610 932 2703 sw
rect 144 2604 10035 2610
rect 144 2564 1000 2604
rect 144 2512 688 2564
rect 740 2552 1000 2564
rect 1052 2552 1312 2604
rect 1364 2552 1624 2604
rect 1676 2552 1936 2604
rect 1988 2552 2248 2604
rect 2300 2552 2560 2604
rect 2612 2552 2872 2604
rect 2924 2552 4925 2604
rect 4977 2552 4991 2604
rect 5043 2552 5114 2604
rect 5166 2552 5426 2604
rect 5478 2552 5738 2604
rect 5790 2552 6050 2604
rect 6102 2552 6361 2604
rect 6413 2552 6673 2604
rect 6725 2552 6986 2604
rect 7038 2552 7298 2604
rect 7350 2552 7610 2604
rect 7662 2552 7922 2604
rect 7974 2552 8234 2604
rect 8286 2552 8546 2604
rect 8598 2552 8858 2604
rect 8910 2552 9170 2604
rect 9222 2552 9482 2604
rect 9534 2552 9794 2604
rect 9846 2552 9917 2604
rect 9969 2552 9983 2604
rect 740 2537 10035 2552
rect 740 2512 1000 2537
rect 144 2493 1000 2512
rect 144 2441 688 2493
rect 740 2485 1000 2493
rect 1052 2485 1312 2537
rect 1364 2485 1624 2537
rect 1676 2485 1936 2537
rect 1988 2485 2248 2537
rect 2300 2485 2560 2537
rect 2612 2485 2872 2537
rect 2924 2522 5114 2537
rect 2924 2485 4925 2522
rect 740 2474 4925 2485
rect 740 2470 4079 2474
rect 740 2441 1000 2470
rect 144 2422 1000 2441
rect 144 2370 688 2422
rect 740 2418 1000 2422
rect 1052 2418 1312 2470
rect 1364 2418 1624 2470
rect 1676 2418 1936 2470
rect 1988 2418 2248 2470
rect 2300 2418 2560 2470
rect 2612 2418 2872 2470
rect 2924 2422 4079 2470
rect 4131 2470 4925 2474
rect 4977 2470 4991 2522
rect 5043 2485 5114 2522
rect 5166 2485 5426 2537
rect 5478 2485 5738 2537
rect 5790 2485 6050 2537
rect 6102 2485 6361 2537
rect 6413 2485 6673 2537
rect 6725 2485 6986 2537
rect 7038 2485 7298 2537
rect 7350 2485 7610 2537
rect 7662 2485 7922 2537
rect 7974 2485 8234 2537
rect 8286 2485 8546 2537
rect 8598 2485 8858 2537
rect 8910 2485 9170 2537
rect 9222 2485 9482 2537
rect 9534 2485 9794 2537
rect 9846 2522 10035 2537
rect 9846 2485 9917 2522
rect 5043 2470 9917 2485
rect 9969 2470 9983 2522
rect 4131 2440 5114 2470
rect 4131 2422 4925 2440
rect 2924 2418 4925 2422
rect 740 2403 4925 2418
rect 740 2370 1000 2403
rect 144 2351 1000 2370
rect 1052 2351 1312 2403
rect 1364 2351 1624 2403
rect 1676 2351 1936 2403
rect 1988 2351 2248 2403
rect 2300 2351 2560 2403
rect 2612 2351 2872 2403
rect 2924 2401 4925 2403
rect 2924 2351 4079 2401
rect 144 2299 688 2351
rect 740 2349 4079 2351
rect 4131 2388 4925 2401
rect 4977 2388 4991 2440
rect 5043 2418 5114 2440
rect 5166 2418 5426 2470
rect 5478 2418 5738 2470
rect 5790 2418 6050 2470
rect 6102 2418 6361 2470
rect 6413 2418 6673 2470
rect 6725 2418 6986 2470
rect 7038 2418 7298 2470
rect 7350 2418 7610 2470
rect 7662 2418 7922 2470
rect 7974 2418 8234 2470
rect 8286 2418 8546 2470
rect 8598 2418 8858 2470
rect 8910 2418 9170 2470
rect 9222 2418 9482 2470
rect 9534 2418 9794 2470
rect 9846 2440 10035 2470
rect 9846 2418 9917 2440
rect 5043 2403 9917 2418
rect 5043 2388 5114 2403
rect 4131 2357 5114 2388
rect 4131 2349 4925 2357
rect 740 2336 4925 2349
rect 740 2299 1000 2336
rect 144 2284 1000 2299
rect 1052 2284 1312 2336
rect 1364 2284 1624 2336
rect 1676 2284 1936 2336
rect 1988 2284 2248 2336
rect 2300 2284 2560 2336
rect 2612 2284 2872 2336
rect 2924 2328 4925 2336
rect 2924 2284 4079 2328
rect 144 2280 4079 2284
rect 144 2228 688 2280
rect 740 2276 4079 2280
rect 4131 2305 4925 2328
rect 4977 2305 4991 2357
rect 5043 2351 5114 2357
rect 5166 2351 5426 2403
rect 5478 2351 5738 2403
rect 5790 2351 6050 2403
rect 6102 2351 6361 2403
rect 6413 2351 6673 2403
rect 6725 2351 6986 2403
rect 7038 2351 7298 2403
rect 7350 2351 7610 2403
rect 7662 2351 7922 2403
rect 7974 2351 8234 2403
rect 8286 2351 8546 2403
rect 8598 2351 8858 2403
rect 8910 2351 9170 2403
rect 9222 2351 9482 2403
rect 9534 2351 9794 2403
rect 9846 2388 9917 2403
rect 9969 2388 9983 2440
rect 9846 2357 10035 2388
rect 9846 2351 9917 2357
rect 5043 2336 9917 2351
rect 5043 2305 5114 2336
rect 4131 2284 5114 2305
rect 5166 2284 5426 2336
rect 5478 2284 5738 2336
rect 5790 2284 6050 2336
rect 6102 2284 6361 2336
rect 6413 2284 6673 2336
rect 6725 2284 6986 2336
rect 7038 2284 7298 2336
rect 7350 2284 7610 2336
rect 7662 2284 7922 2336
rect 7974 2284 8234 2336
rect 8286 2284 8546 2336
rect 8598 2284 8858 2336
rect 8910 2284 9170 2336
rect 9222 2284 9482 2336
rect 9534 2284 9794 2336
rect 9846 2305 9917 2336
rect 9969 2305 9983 2357
rect 9846 2284 10035 2305
rect 4131 2276 10035 2284
rect 740 2274 10035 2276
rect 740 2269 4925 2274
rect 740 2228 1000 2269
rect 144 2217 1000 2228
rect 1052 2217 1312 2269
rect 1364 2217 1624 2269
rect 1676 2217 1936 2269
rect 1988 2217 2248 2269
rect 2300 2217 2560 2269
rect 2612 2217 2872 2269
rect 2924 2255 4925 2269
rect 2924 2217 4079 2255
rect 144 2209 4079 2217
rect 144 2157 688 2209
rect 740 2203 4079 2209
rect 4131 2222 4925 2255
rect 4977 2222 4991 2274
rect 5043 2269 9917 2274
rect 5043 2222 5114 2269
rect 4131 2217 5114 2222
rect 5166 2217 5426 2269
rect 5478 2217 5738 2269
rect 5790 2217 6050 2269
rect 6102 2217 6361 2269
rect 6413 2217 6673 2269
rect 6725 2217 6986 2269
rect 7038 2217 7298 2269
rect 7350 2217 7610 2269
rect 7662 2217 7922 2269
rect 7974 2217 8234 2269
rect 8286 2217 8546 2269
rect 8598 2217 8858 2269
rect 8910 2217 9170 2269
rect 9222 2217 9482 2269
rect 9534 2217 9794 2269
rect 9846 2222 9917 2269
rect 9969 2222 9983 2274
rect 9846 2217 10035 2222
rect 4131 2203 10035 2217
rect 740 2202 10035 2203
rect 740 2157 1000 2202
rect 144 2150 1000 2157
rect 1052 2150 1312 2202
rect 1364 2150 1624 2202
rect 1676 2150 1936 2202
rect 1988 2150 2248 2202
rect 2300 2150 2560 2202
rect 2612 2150 2872 2202
rect 2924 2191 5114 2202
rect 2924 2182 4925 2191
rect 2924 2150 4079 2182
rect 144 2138 4079 2150
rect 144 2086 688 2138
rect 740 2135 4079 2138
rect 740 2086 1000 2135
rect 144 2083 1000 2086
rect 1052 2083 1312 2135
rect 1364 2083 1624 2135
rect 1676 2083 1936 2135
rect 1988 2083 2248 2135
rect 2300 2083 2560 2135
rect 2612 2083 2872 2135
rect 2924 2130 4079 2135
rect 4131 2139 4925 2182
rect 4977 2139 4991 2191
rect 5043 2150 5114 2191
rect 5166 2150 5426 2202
rect 5478 2150 5738 2202
rect 5790 2150 6050 2202
rect 6102 2150 6361 2202
rect 6413 2150 6673 2202
rect 6725 2150 6986 2202
rect 7038 2150 7298 2202
rect 7350 2150 7610 2202
rect 7662 2150 7922 2202
rect 7974 2150 8234 2202
rect 8286 2150 8546 2202
rect 8598 2150 8858 2202
rect 8910 2150 9170 2202
rect 9222 2150 9482 2202
rect 9534 2150 9794 2202
rect 9846 2191 10035 2202
rect 9846 2150 9917 2191
rect 5043 2139 9917 2150
rect 9969 2139 9983 2191
rect 4131 2135 10035 2139
rect 4131 2130 5114 2135
rect 2924 2108 5114 2130
rect 2924 2083 4079 2108
rect 144 2068 4079 2083
rect 144 2016 688 2068
rect 740 2016 1000 2068
rect 1052 2016 1312 2068
rect 1364 2016 1624 2068
rect 1676 2016 1936 2068
rect 1988 2016 2248 2068
rect 2300 2016 2560 2068
rect 2612 2016 2872 2068
rect 2924 2056 4079 2068
rect 4131 2056 4925 2108
rect 4977 2056 4991 2108
rect 5043 2083 5114 2108
rect 5166 2083 5426 2135
rect 5478 2083 5738 2135
rect 5790 2083 6050 2135
rect 6102 2083 6361 2135
rect 6413 2083 6673 2135
rect 6725 2083 6986 2135
rect 7038 2083 7298 2135
rect 7350 2083 7610 2135
rect 7662 2083 7922 2135
rect 7974 2083 8234 2135
rect 8286 2083 8546 2135
rect 8598 2083 8858 2135
rect 8910 2083 9170 2135
rect 9222 2083 9482 2135
rect 9534 2083 9794 2135
rect 9846 2108 10035 2135
rect 9846 2083 9917 2108
rect 5043 2068 9917 2083
rect 5043 2056 5114 2068
rect 2924 2016 5114 2056
rect 5166 2016 5426 2068
rect 5478 2016 5738 2068
rect 5790 2016 6050 2068
rect 6102 2016 6361 2068
rect 6413 2016 6673 2068
rect 6725 2016 6986 2068
rect 7038 2016 7298 2068
rect 7350 2016 7610 2068
rect 7662 2016 7922 2068
rect 7974 2016 8234 2068
rect 8286 2016 8546 2068
rect 8598 2016 8858 2068
rect 8910 2016 9170 2068
rect 9222 2016 9482 2068
rect 9534 2016 9794 2068
rect 9846 2056 9917 2068
rect 9969 2056 9983 2108
rect 9846 2016 10035 2056
rect 144 2010 10035 2016
rect 686 1902 3210 1954
rect 3262 1902 3274 1954
rect 3326 1902 9848 1954
rect 686 1865 9848 1871
rect 686 1813 844 1865
rect 896 1813 1156 1865
rect 1208 1813 1468 1865
rect 1520 1813 1780 1865
rect 1832 1813 2092 1865
rect 2144 1813 2404 1865
rect 2456 1813 2716 1865
rect 2768 1813 5270 1865
rect 5322 1813 5582 1865
rect 5634 1813 5894 1865
rect 5946 1813 6205 1865
rect 6257 1813 6517 1865
rect 6569 1813 6830 1865
rect 6882 1813 7142 1865
rect 7194 1813 7454 1865
rect 7506 1813 7766 1865
rect 7818 1813 8078 1865
rect 8130 1813 8390 1865
rect 8442 1813 8702 1865
rect 8754 1813 9014 1865
rect 9066 1813 9326 1865
rect 9378 1813 9638 1865
rect 9690 1813 9848 1865
rect 686 1798 9848 1813
rect 686 1746 844 1798
rect 896 1746 1156 1798
rect 1208 1746 1468 1798
rect 1520 1746 1780 1798
rect 1832 1746 2092 1798
rect 2144 1746 2404 1798
rect 2456 1746 2716 1798
rect 2768 1746 5270 1798
rect 5322 1746 5582 1798
rect 5634 1746 5894 1798
rect 5946 1746 6205 1798
rect 6257 1746 6517 1798
rect 6569 1746 6830 1798
rect 6882 1746 7142 1798
rect 7194 1746 7454 1798
rect 7506 1746 7766 1798
rect 7818 1746 8078 1798
rect 8130 1746 8390 1798
rect 8442 1746 8702 1798
rect 8754 1746 9014 1798
rect 9066 1746 9326 1798
rect 9378 1746 9638 1798
rect 9690 1746 9848 1798
rect 686 1731 9848 1746
rect 686 1679 844 1731
rect 896 1679 1156 1731
rect 1208 1679 1468 1731
rect 1520 1679 1780 1731
rect 1832 1679 2092 1731
rect 2144 1679 2404 1731
rect 2456 1679 2716 1731
rect 2768 1679 5270 1731
rect 5322 1679 5582 1731
rect 5634 1679 5894 1731
rect 5946 1679 6205 1731
rect 6257 1679 6517 1731
rect 6569 1679 6830 1731
rect 6882 1679 7142 1731
rect 7194 1679 7454 1731
rect 7506 1679 7766 1731
rect 7818 1679 8078 1731
rect 8130 1679 8390 1731
rect 8442 1679 8702 1731
rect 8754 1679 9014 1731
rect 9066 1679 9326 1731
rect 9378 1679 9638 1731
rect 9690 1679 9848 1731
rect 686 1664 9848 1679
rect 686 1612 844 1664
rect 896 1612 1156 1664
rect 1208 1612 1468 1664
rect 1520 1612 1780 1664
rect 1832 1612 2092 1664
rect 2144 1612 2404 1664
rect 2456 1612 2716 1664
rect 2768 1612 5270 1664
rect 5322 1612 5582 1664
rect 5634 1612 5894 1664
rect 5946 1612 6205 1664
rect 6257 1612 6517 1664
rect 6569 1612 6830 1664
rect 6882 1612 7142 1664
rect 7194 1612 7454 1664
rect 7506 1612 7766 1664
rect 7818 1612 8078 1664
rect 8130 1612 8390 1664
rect 8442 1612 8702 1664
rect 8754 1612 9014 1664
rect 9066 1612 9326 1664
rect 9378 1612 9638 1664
rect 9690 1612 9848 1664
rect 686 1597 9848 1612
rect 686 1545 844 1597
rect 896 1545 1156 1597
rect 1208 1545 1468 1597
rect 1520 1545 1780 1597
rect 1832 1545 2092 1597
rect 2144 1545 2404 1597
rect 2456 1545 2716 1597
rect 2768 1545 5270 1597
rect 5322 1545 5582 1597
rect 5634 1545 5894 1597
rect 5946 1545 6205 1597
rect 6257 1545 6517 1597
rect 6569 1545 6830 1597
rect 6882 1545 7142 1597
rect 7194 1545 7454 1597
rect 7506 1545 7766 1597
rect 7818 1545 8078 1597
rect 8130 1545 8390 1597
rect 8442 1545 8702 1597
rect 8754 1545 9014 1597
rect 9066 1545 9326 1597
rect 9378 1545 9638 1597
rect 9690 1545 9848 1597
rect 686 1530 9848 1545
rect 686 1478 844 1530
rect 896 1478 1156 1530
rect 1208 1478 1468 1530
rect 1520 1478 1780 1530
rect 1832 1478 2092 1530
rect 2144 1478 2404 1530
rect 2456 1478 2716 1530
rect 2768 1478 5270 1530
rect 5322 1478 5582 1530
rect 5634 1478 5894 1530
rect 5946 1478 6205 1530
rect 6257 1478 6517 1530
rect 6569 1478 6830 1530
rect 6882 1478 7142 1530
rect 7194 1478 7454 1530
rect 7506 1478 7766 1530
rect 7818 1478 8078 1530
rect 8130 1478 8390 1530
rect 8442 1478 8702 1530
rect 8754 1478 9014 1530
rect 9066 1478 9326 1530
rect 9378 1478 9638 1530
rect 9690 1478 9848 1530
rect 686 1463 9848 1478
rect 686 1411 844 1463
rect 896 1411 1156 1463
rect 1208 1411 1468 1463
rect 1520 1411 1780 1463
rect 1832 1411 2092 1463
rect 2144 1411 2404 1463
rect 2456 1411 2716 1463
rect 2768 1411 5270 1463
rect 5322 1411 5582 1463
rect 5634 1411 5894 1463
rect 5946 1411 6205 1463
rect 6257 1411 6517 1463
rect 6569 1411 6830 1463
rect 6882 1411 7142 1463
rect 7194 1411 7454 1463
rect 7506 1411 7766 1463
rect 7818 1411 8078 1463
rect 8130 1411 8390 1463
rect 8442 1411 8702 1463
rect 8754 1411 9014 1463
rect 9066 1411 9326 1463
rect 9378 1411 9638 1463
rect 9690 1411 9848 1463
rect 686 1396 9848 1411
rect 686 1344 844 1396
rect 896 1344 1156 1396
rect 1208 1344 1468 1396
rect 1520 1344 1780 1396
rect 1832 1344 2092 1396
rect 2144 1344 2404 1396
rect 2456 1344 2716 1396
rect 2768 1344 5270 1396
rect 5322 1344 5582 1396
rect 5634 1344 5894 1396
rect 5946 1344 6205 1396
rect 6257 1344 6517 1396
rect 6569 1344 6830 1396
rect 6882 1344 7142 1396
rect 7194 1344 7454 1396
rect 7506 1344 7766 1396
rect 7818 1344 8078 1396
rect 8130 1344 8390 1396
rect 8442 1344 8702 1396
rect 8754 1344 9014 1396
rect 9066 1344 9326 1396
rect 9378 1344 9638 1396
rect 9690 1344 9848 1396
rect 686 1329 9848 1344
rect 686 1277 844 1329
rect 896 1277 1156 1329
rect 1208 1277 1468 1329
rect 1520 1277 1780 1329
rect 1832 1277 2092 1329
rect 2144 1277 2404 1329
rect 2456 1277 2716 1329
rect 2768 1277 5270 1329
rect 5322 1277 5582 1329
rect 5634 1277 5894 1329
rect 5946 1277 6205 1329
rect 6257 1277 6517 1329
rect 6569 1277 6830 1329
rect 6882 1277 7142 1329
rect 7194 1277 7454 1329
rect 7506 1277 7766 1329
rect 7818 1277 8078 1329
rect 8130 1277 8390 1329
rect 8442 1277 8702 1329
rect 8754 1277 9014 1329
rect 9066 1277 9326 1329
rect 9378 1277 9638 1329
rect 9690 1277 9848 1329
rect 686 1271 9848 1277
rect 686 1187 3210 1239
rect 3262 1187 3274 1239
rect 3326 1187 9848 1239
rect -30 497 10507 870
rect -30 445 326 497
rect 378 445 391 497
rect 443 445 456 497
rect 508 445 521 497
rect 573 445 586 497
rect 638 445 651 497
rect 703 445 716 497
rect 768 445 781 497
rect 833 445 846 497
rect 898 445 911 497
rect 963 445 976 497
rect 1028 445 1041 497
rect 1093 445 1106 497
rect 1158 445 1171 497
rect 1223 445 1236 497
rect 1288 445 1301 497
rect 1353 445 1366 497
rect 1418 445 1431 497
rect 1483 445 1496 497
rect 1548 445 1561 497
rect 1613 445 1626 497
rect 1678 445 1691 497
rect 1743 445 1756 497
rect 1808 445 1821 497
rect 1873 445 1886 497
rect 1938 445 1951 497
rect 2003 445 2016 497
rect 2068 445 2081 497
rect 2133 445 2146 497
rect 2198 445 2211 497
rect 2263 445 2275 497
rect 2327 445 2339 497
rect 2391 445 2403 497
rect 2455 445 2467 497
rect 2519 445 2531 497
rect 2583 445 2595 497
rect 2647 445 2659 497
rect 2711 445 2723 497
rect 2775 445 2787 497
rect 2839 445 2851 497
rect 2903 445 2915 497
rect 2967 445 2979 497
rect 3031 445 3043 497
rect 3095 445 3107 497
rect 3159 445 3171 497
rect 3223 445 3235 497
rect 3287 490 10507 497
rect 3287 445 3728 490
rect -30 438 3728 445
rect 3780 438 3828 490
rect 3880 438 3928 490
rect 3980 438 4029 490
rect 4081 438 4130 490
rect 4182 438 4231 490
rect 4283 438 4332 490
rect 4384 438 4433 490
rect 4485 438 10507 490
rect -30 232 10507 438
use nfet_CDNS_5595914180826  nfet_CDNS_5595914180826_0
timestamp 1701704242
transform -1 0 4233 0 1 1482
box -82 -32 338 1032
use nfet_CDNS_5595914180828  nfet_CDNS_5595914180828_0
timestamp 1701704242
transform 1 0 5168 0 -1 5264
box -82 -32 4706 2032
use nfet_CDNS_5595914180828  nfet_CDNS_5595914180828_1
timestamp 1701704242
transform -1 0 9792 0 1 664
box -82 -32 4706 2032
use pfet_CDNS_5595914180830  pfet_CDNS_5595914180830_0
timestamp 1701704242
transform -1 0 2870 0 1 839
box -122 -66 2250 2066
use pfet_CDNS_5595914180830  pfet_CDNS_5595914180830_1
timestamp 1701704242
transform -1 0 2870 0 -1 5089
box -122 -66 2250 2066
use s8_esd_res75only_small  s8_esd_res75only_small_0
timestamp 1701704242
transform 0 1 3911 1 0 474
box 0 0 882 404
<< labels >>
flabel metal1 s 1451 3002 1632 3043 3 FreeSans 520 0 0 0 pgate_sl_h_n
port 1 nsew
flabel metal1 s 1733 2885 1929 2922 3 FreeSans 520 0 0 0 pgate_sr_h_n
port 2 nsew
flabel metal1 s 7996 3186 8259 3214 3 FreeSans 520 180 0 0 ngate_sl_h
port 3 nsew
flabel metal1 s 7984 2713 8161 2744 3 FreeSans 520 180 0 0 ngate_sr_h
port 4 nsew
flabel metal1 s 4046 2538 4160 2563 3 FreeSans 520 180 0 0 nmid_h
port 5 nsew
flabel metal2 s 915 4260 1148 4860 3 FreeSans 520 0 0 0 amuxbus_l
port 6 nsew
flabel metal2 s 760 1271 980 1871 3 FreeSans 520 0 0 0 amuxbus_r
port 7 nsew
flabel metal2 s 221 5252 474 5715 3 FreeSans 520 0 0 0 vdda
port 8 nsew
flabel metal2 s 418 513 891 724 3 FreeSans 520 180 0 0 vssa
port 9 nsew
flabel comment s 1225 392 1225 392 0 FreeSans 600 180 0 0 condiode
flabel comment s 5715 5538 5715 5538 0 FreeSans 600 180 0 0 condiode
flabel comment s 4059 421 4059 421 0 FreeSans 600 180 0 0 condiode
<< properties >>
string GDS_END 540200
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 42628
<< end >>
