magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< metal2 >>
rect 0 465 216 474
rect 0 0 216 9
<< via2 >>
rect 0 9 216 465
<< metal3 >>
rect -5 465 221 470
rect -5 9 0 465
rect 216 9 221 465
rect -5 4 221 9
<< properties >>
string GDS_END 89697512
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 89696228
<< end >>
