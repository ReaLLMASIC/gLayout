magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< metal2 >>
rect 0 1745 536 1754
rect 0 0 536 9
<< via2 >>
rect 0 9 536 1745
<< metal3 >>
rect -5 1745 541 1750
rect -5 9 0 1745
rect 536 9 541 1745
rect -5 4 541 9
<< properties >>
string GDS_END 93372738
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 93362750
<< end >>
