magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< pwell >>
rect -82 -26 282 110
<< mvnmos >>
rect 0 0 200 84
<< mvndiff >>
rect -56 46 0 84
rect -56 12 -45 46
rect -11 12 0 46
rect -56 0 0 12
rect 200 46 256 84
rect 200 12 211 46
rect 245 12 256 46
rect 200 0 256 12
<< mvndiffc >>
rect -45 12 -11 46
rect 211 12 245 46
<< poly >>
rect 0 84 200 116
rect 0 -32 200 0
<< locali >>
rect -45 46 -11 62
rect -45 -4 -11 12
rect 211 46 245 62
rect 211 -4 245 12
use hvDFL1sd2_CDNS_52468879185681  hvDFL1sd2_CDNS_52468879185681_0
timestamp 1701704242
transform -1 0 0 0 1 0
box 0 0 1 1
use hvDFL1sd2_CDNS_52468879185681  hvDFL1sd2_CDNS_52468879185681_1
timestamp 1701704242
transform 1 0 200 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s -28 29 -28 29 0 FreeSans 300 0 0 0 S
flabel comment s 228 29 228 29 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 85637356
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85636462
<< end >>
