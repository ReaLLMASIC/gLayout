magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -119 -66 1623 666
<< mvpmos >>
rect 0 0 100 600
rect 156 0 256 600
rect 312 0 412 600
rect 468 0 568 600
rect 624 0 724 600
rect 780 0 880 600
rect 936 0 1036 600
rect 1092 0 1192 600
rect 1248 0 1348 600
rect 1404 0 1504 600
<< mvpdiff >>
rect -50 0 0 600
rect 1504 0 1554 600
<< poly >>
rect 0 600 100 632
rect 0 -32 100 0
rect 156 600 256 632
rect 156 -32 256 0
rect 312 600 412 632
rect 312 -32 412 0
rect 468 600 568 632
rect 468 -32 568 0
rect 624 600 724 632
rect 624 -32 724 0
rect 780 600 880 632
rect 780 -32 880 0
rect 936 600 1036 632
rect 936 -32 1036 0
rect 1092 600 1192 632
rect 1092 -32 1192 0
rect 1248 600 1348 632
rect 1248 -32 1348 0
rect 1404 600 1504 632
rect 1404 -32 1504 0
<< locali >>
rect -45 -4 -11 538
rect 111 -4 145 538
rect 267 -4 301 538
rect 423 -4 457 538
rect 579 -4 613 538
rect 735 -4 769 538
rect 891 -4 925 538
rect 1047 -4 1081 538
rect 1203 -4 1237 538
rect 1359 -4 1393 538
rect 1515 -4 1549 538
use DFL1sd2_CDNS_5246887918535  DFL1sd2_CDNS_5246887918535_0
timestamp 1701704242
transform 1 0 1348 0 1 0
box -36 -36 92 636
use DFL1sd2_CDNS_5246887918535  DFL1sd2_CDNS_5246887918535_1
timestamp 1701704242
transform 1 0 1192 0 1 0
box -36 -36 92 636
use DFL1sd2_CDNS_5246887918535  DFL1sd2_CDNS_5246887918535_2
timestamp 1701704242
transform 1 0 1036 0 1 0
box -36 -36 92 636
use DFL1sd2_CDNS_5246887918535  DFL1sd2_CDNS_5246887918535_3
timestamp 1701704242
transform 1 0 880 0 1 0
box -36 -36 92 636
use DFL1sd2_CDNS_5246887918535  DFL1sd2_CDNS_5246887918535_4
timestamp 1701704242
transform 1 0 724 0 1 0
box -36 -36 92 636
use DFL1sd2_CDNS_5246887918535  DFL1sd2_CDNS_5246887918535_5
timestamp 1701704242
transform 1 0 568 0 1 0
box -36 -36 92 636
use DFL1sd2_CDNS_5246887918535  DFL1sd2_CDNS_5246887918535_6
timestamp 1701704242
transform 1 0 412 0 1 0
box -36 -36 92 636
use DFL1sd2_CDNS_5246887918535  DFL1sd2_CDNS_5246887918535_7
timestamp 1701704242
transform 1 0 256 0 1 0
box -36 -36 92 636
use DFL1sd2_CDNS_5246887918535  DFL1sd2_CDNS_5246887918535_8
timestamp 1701704242
transform 1 0 100 0 1 0
box -36 -36 92 636
use DFL1sd_CDNS_5246887918534  DFL1sd_CDNS_5246887918534_0
timestamp 1701704242
transform -1 0 0 0 1 0
box -36 -36 89 636
use DFL1sd_CDNS_5246887918534  DFL1sd_CDNS_5246887918534_1
timestamp 1701704242
transform 1 0 1504 0 1 0
box -36 -36 89 636
<< labels >>
flabel comment s -28 267 -28 267 0 FreeSans 300 0 0 0 S
flabel comment s 128 267 128 267 0 FreeSans 300 0 0 0 D
flabel comment s 284 267 284 267 0 FreeSans 300 0 0 0 S
flabel comment s 440 267 440 267 0 FreeSans 300 0 0 0 D
flabel comment s 596 267 596 267 0 FreeSans 300 0 0 0 S
flabel comment s 752 267 752 267 0 FreeSans 300 0 0 0 D
flabel comment s 908 267 908 267 0 FreeSans 300 0 0 0 S
flabel comment s 1064 267 1064 267 0 FreeSans 300 0 0 0 D
flabel comment s 1220 267 1220 267 0 FreeSans 300 0 0 0 S
flabel comment s 1376 267 1376 267 0 FreeSans 300 0 0 0 D
flabel comment s 1532 267 1532 267 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 24802994
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 24797516
<< end >>
