magic
tech sky130B
magscale 1 2
timestamp 1701704242
use sky130_fd_pr__hvdfl1sd__example_55959141808102  sky130_fd_pr__hvdfl1sd__example_55959141808102_0
timestamp 1701704242
transform -1 0 0 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 20907636
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 20906716
<< end >>
